

module b22_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P3_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, 
        P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN, 
        P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN, 
        P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN, 
        P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN, 
        P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN, 
        P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN, 
        P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN, 
        P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN, 
        P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN, 
        P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN,
         P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN,
         P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN,
         P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN,
         P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN,
         P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN,
         P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN,
         P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN,
         P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN,
         P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN,
         P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN,
         P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN,
         P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN,
         P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN,
         P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN,
         P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN,
         P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN,
         P3_ADDR_REG_3__SCAN_IN, P3_ADDR_REG_4__SCAN_IN,
         P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN,
         P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN,
         P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN,
         P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN,
         P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN,
         P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN,
         P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN,
         P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN,
         P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN,
         P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN,
         P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN,
         P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN,
         P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN,
         P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN,
         P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN,
         P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN,
         P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN,
         P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN,
         P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN,
         P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN,
         P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN,
         P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN,
         P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN,
         P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN,
         P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN,
         P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN,
         P3_REG0_REG_3__SCAN_IN, P3_REG0_REG_4__SCAN_IN,
         P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN,
         P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN,
         P3_REG0_REG_9__SCAN_IN, P3_REG0_REG_10__SCAN_IN,
         P3_REG0_REG_11__SCAN_IN, P3_REG0_REG_12__SCAN_IN,
         P3_REG0_REG_13__SCAN_IN, P3_REG0_REG_14__SCAN_IN,
         P3_REG0_REG_15__SCAN_IN, P3_REG0_REG_16__SCAN_IN,
         P3_REG0_REG_17__SCAN_IN, P3_REG0_REG_18__SCAN_IN,
         P3_REG0_REG_19__SCAN_IN, P3_REG0_REG_20__SCAN_IN,
         P3_REG0_REG_21__SCAN_IN, P3_REG0_REG_22__SCAN_IN,
         P3_REG0_REG_23__SCAN_IN, P3_REG0_REG_24__SCAN_IN,
         P3_REG0_REG_25__SCAN_IN, P3_REG0_REG_26__SCAN_IN,
         P3_REG0_REG_27__SCAN_IN, P3_REG0_REG_28__SCAN_IN,
         P3_REG0_REG_29__SCAN_IN, P3_REG0_REG_30__SCAN_IN,
         P3_REG0_REG_31__SCAN_IN, P3_REG1_REG_0__SCAN_IN,
         P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN,
         P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN,
         P3_REG1_REG_5__SCAN_IN, P3_REG1_REG_6__SCAN_IN,
         P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN,
         P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN,
         P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN,
         P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN,
         P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN,
         P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN,
         P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN,
         P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN,
         P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN,
         P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN,
         P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN,
         P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN,
         P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN,
         P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN,
         P3_REG2_REG_3__SCAN_IN, P3_REG2_REG_4__SCAN_IN,
         P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN,
         P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN,
         P3_REG2_REG_9__SCAN_IN, P3_REG2_REG_10__SCAN_IN,
         P3_REG2_REG_11__SCAN_IN, P3_REG2_REG_12__SCAN_IN,
         P3_REG2_REG_13__SCAN_IN, P3_REG2_REG_14__SCAN_IN,
         P3_REG2_REG_15__SCAN_IN, P3_REG2_REG_16__SCAN_IN,
         P3_REG2_REG_17__SCAN_IN, P3_REG2_REG_18__SCAN_IN,
         P3_REG2_REG_19__SCAN_IN, P3_REG2_REG_20__SCAN_IN,
         P3_REG2_REG_21__SCAN_IN, P3_REG2_REG_22__SCAN_IN,
         P3_REG2_REG_23__SCAN_IN, P3_REG2_REG_24__SCAN_IN,
         P3_REG2_REG_25__SCAN_IN, P3_REG2_REG_26__SCAN_IN,
         P3_REG2_REG_27__SCAN_IN, P3_REG2_REG_28__SCAN_IN,
         P3_REG2_REG_29__SCAN_IN, P3_REG2_REG_30__SCAN_IN,
         P3_REG2_REG_31__SCAN_IN, P3_ADDR_REG_19__SCAN_IN,
         P3_ADDR_REG_18__SCAN_IN, P3_ADDR_REG_17__SCAN_IN,
         P3_ADDR_REG_16__SCAN_IN, P3_ADDR_REG_15__SCAN_IN,
         P3_ADDR_REG_14__SCAN_IN, P3_ADDR_REG_13__SCAN_IN,
         P3_ADDR_REG_12__SCAN_IN, P3_ADDR_REG_11__SCAN_IN,
         P3_ADDR_REG_10__SCAN_IN;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16058;

  AOI211_X1 U7255 ( .C1(n13198), .C2(n13197), .A(n13196), .B(n13195), .ZN(
        n13199) );
  AND2_X1 U7256 ( .A1(n9117), .A2(n9116), .ZN(n12348) );
  AOI21_X1 U7257 ( .B1(n7766), .B2(n7189), .A(n7765), .ZN(n9027) );
  NOR2_X1 U7258 ( .A1(n12968), .A2(n7632), .ZN(n7631) );
  INV_X1 U7259 ( .A(n14586), .ZN(n14522) );
  CLKBUF_X1 U7260 ( .A(n12728), .Z(n12871) );
  CLKBUF_X2 U7261 ( .A(n12510), .Z(n7158) );
  NAND2_X1 U7262 ( .A1(n8924), .A2(n8923), .ZN(n11218) );
  INV_X4 U7263 ( .A(n8883), .ZN(n9362) );
  INV_X2 U7264 ( .A(n10335), .ZN(n9987) );
  NAND2_X2 U7265 ( .A1(n7194), .A2(n8797), .ZN(n13932) );
  NAND2_X1 U7266 ( .A1(n8686), .A2(n8685), .ZN(n12262) );
  NAND2_X1 U7267 ( .A1(n8685), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8152) );
  OAI21_X1 U7268 ( .B1(n8709), .B2(P3_IR_REG_24__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8682) );
  INV_X1 U7269 ( .A(n9145), .ZN(n8786) );
  XNOR2_X1 U7270 ( .A(n7961), .B(n9605), .ZN(n15429) );
  NAND2_X1 U7271 ( .A1(n8768), .A2(n8767), .ZN(n9525) );
  AND4_X1 U7272 ( .A1(n9212), .A2(n8751), .A3(n9162), .A4(n9526), .ZN(n8754)
         );
  INV_X1 U7274 ( .A(n16058), .ZN(n7155) );
  AND4_X1 U7275 ( .A1(n8767), .A2(n8773), .A3(n8764), .A4(n8750), .ZN(n8755)
         );
  INV_X1 U7276 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8773) );
  INV_X1 U7277 ( .A(n13361), .ZN(n12686) );
  INV_X1 U7278 ( .A(n15443), .ZN(n10051) );
  AOI21_X1 U7279 ( .B1(n9660), .B2(n9659), .A(n7233), .ZN(n15870) );
  INV_X1 U7281 ( .A(n8215), .ZN(n8495) );
  INV_X1 U7282 ( .A(n12635), .ZN(n12641) );
  INV_X1 U7283 ( .A(n12509), .ZN(n12496) );
  INV_X1 U7284 ( .A(n9040), .ZN(n8897) );
  INV_X1 U7285 ( .A(n8794), .ZN(n9474) );
  INV_X2 U7286 ( .A(n14282), .ZN(n14348) );
  AND2_X1 U7287 ( .A1(n9094), .A2(n9093), .ZN(n15997) );
  AND2_X1 U7288 ( .A1(n8970), .A2(n8969), .ZN(n11643) );
  INV_X1 U7289 ( .A(n11965), .ZN(n11867) );
  AND3_X1 U7290 ( .A1(n8253), .A2(n8252), .A3(n8251), .ZN(n11846) );
  XNOR2_X1 U7291 ( .A(n8183), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8186) );
  MUX2_X1 U7292 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8684), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n8686) );
  INV_X1 U7293 ( .A(n8098), .ZN(n14151) );
  INV_X1 U7294 ( .A(n15997), .ZN(n12141) );
  AOI211_X1 U7295 ( .C1(n14347), .C2(n14305), .A(n14304), .B(n14303), .ZN(
        n14306) );
  NAND2_X1 U7296 ( .A1(n9688), .A2(n9687), .ZN(n12738) );
  NAND2_X1 U7297 ( .A1(n9678), .A2(n9677), .ZN(n12729) );
  NAND3_X1 U7298 ( .A1(n7196), .A2(n8225), .A3(n8227), .ZN(n7349) );
  XNOR2_X1 U7299 ( .A(n8185), .B(n8184), .ZN(n13725) );
  NAND2_X1 U7300 ( .A1(n9031), .A2(n9011), .ZN(n10471) );
  AND4_X1 U7301 ( .A1(n8278), .A2(n8140), .A3(n8282), .A4(n8297), .ZN(n7156)
         );
  BUF_X1 U7302 ( .A(n8229), .Z(n12510) );
  AND2_X2 U7303 ( .A1(n7717), .A2(n7342), .ZN(n7715) );
  OAI21_X2 U7304 ( .B1(n15011), .B2(n7906), .A(n7904), .ZN(n14977) );
  AND2_X2 U7305 ( .A1(n7466), .A2(n7156), .ZN(n8324) );
  AND4_X2 U7306 ( .A1(n8145), .A2(n8144), .A3(n8143), .A4(n8142), .ZN(n8096)
         );
  INV_X1 U7307 ( .A(n13929), .ZN(n10758) );
  OAI21_X2 U7308 ( .B1(n11041), .B2(n10016), .A(n10017), .ZN(n11448) );
  OAI21_X2 U7309 ( .B1(n14677), .B2(n7800), .A(n7798), .ZN(n7797) );
  NAND2_X2 U7310 ( .A1(n14634), .A2(n14638), .ZN(n14677) );
  NAND2_X2 U7311 ( .A1(n12001), .A2(n12000), .ZN(n12228) );
  NAND2_X2 U7312 ( .A1(n11999), .A2(n11998), .ZN(n12001) );
  AOI21_X1 U7313 ( .B1(n10618), .B2(n10617), .A(n10616), .ZN(n10626) );
  NAND2_X2 U7314 ( .A1(n14635), .A2(n14636), .ZN(n14634) );
  OR2_X2 U7315 ( .A1(n13521), .A2(n13522), .ZN(n13519) );
  INV_X4 U7316 ( .A(n8806), .ZN(n10276) );
  NAND2_X2 U7317 ( .A1(n8161), .A2(n8160), .ZN(n8806) );
  XNOR2_X2 U7318 ( .A(n8780), .B(n12960), .ZN(n12484) );
  NAND2_X2 U7319 ( .A1(n12959), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8780) );
  NAND2_X2 U7320 ( .A1(n12389), .A2(n12388), .ZN(n14437) );
  AND2_X2 U7321 ( .A1(n14355), .A2(n14227), .ZN(n14216) );
  NOR2_X2 U7322 ( .A1(n15115), .A2(n14964), .ZN(n14953) );
  AOI21_X2 U7323 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(n15656), .A(n15655), .ZN(
        n15659) );
  INV_X2 U7324 ( .A(n14585), .ZN(n14492) );
  AND2_X4 U7325 ( .A1(n10583), .A2(n11221), .ZN(n14533) );
  BUF_X4 U7326 ( .A(n10240), .Z(n13773) );
  NAND2_X2 U7327 ( .A1(n8664), .A2(n8663), .ZN(n7157) );
  NAND2_X2 U7328 ( .A1(n8664), .A2(n8663), .ZN(n10850) );
  INV_X4 U7329 ( .A(n12695), .ZN(n13728) );
  AND3_X4 U7330 ( .A1(n9530), .A2(n12085), .A3(n9563), .ZN(n16024) );
  INV_X1 U7331 ( .A(n12085), .ZN(n14076) );
  BUF_X4 U7332 ( .A(n8098), .Z(n14282) );
  AND2_X2 U7333 ( .A1(n7642), .A2(n8236), .ZN(n11326) );
  NAND2_X2 U7334 ( .A1(n7308), .A2(n11310), .ZN(n11312) );
  AOI21_X1 U7335 ( .B1(n8983), .B2(n8982), .A(n7177), .ZN(n7766) );
  AOI21_X1 U7336 ( .B1(n8918), .B2(n8917), .A(n8916), .ZN(n8935) );
  AND2_X2 U7337 ( .A1(n8948), .A2(n8947), .ZN(n11546) );
  NAND2_X1 U7338 ( .A1(n11408), .A2(n15860), .ZN(n15867) );
  NOR2_X1 U7339 ( .A1(n10758), .A2(n14348), .ZN(n10247) );
  INV_X1 U7340 ( .A(n7349), .ZN(n11316) );
  CLKBUF_X2 U7341 ( .A(n8242), .Z(n12503) );
  INV_X1 U7342 ( .A(n12704), .ZN(n10633) );
  INV_X2 U7343 ( .A(n9395), .ZN(n9467) );
  INV_X1 U7344 ( .A(n13725), .ZN(n8187) );
  AND2_X1 U7345 ( .A1(n7506), .A2(n7339), .ZN(n10216) );
  AND3_X1 U7346 ( .A1(n15073), .A2(n15072), .A3(n15071), .ZN(n15384) );
  NOR2_X1 U7347 ( .A1(n7411), .A2(n7410), .ZN(n12701) );
  AND2_X1 U7348 ( .A1(n10044), .A2(n14876), .ZN(n14862) );
  NAND2_X1 U7349 ( .A1(n8072), .A2(n8071), .ZN(n14115) );
  OR2_X1 U7350 ( .A1(n14144), .A2(n14127), .ZN(n8072) );
  NAND2_X1 U7351 ( .A1(n13784), .A2(n13759), .ZN(n13846) );
  NAND2_X1 U7352 ( .A1(n14145), .A2(n7200), .ZN(n14144) );
  NAND2_X1 U7353 ( .A1(n14927), .A2(n14926), .ZN(n14925) );
  OR2_X1 U7354 ( .A1(n9195), .A2(n9196), .ZN(n9197) );
  AND2_X1 U7355 ( .A1(n14068), .A2(n14067), .ZN(n14304) );
  NAND2_X1 U7356 ( .A1(n14163), .A2(n14164), .ZN(n14166) );
  NAND2_X1 U7357 ( .A1(n13011), .A2(n13010), .ZN(n13144) );
  AND2_X1 U7358 ( .A1(n14945), .A2(n10036), .ZN(n14932) );
  XNOR2_X1 U7359 ( .A(n9385), .B(n9384), .ZN(n12861) );
  NAND2_X1 U7360 ( .A1(n9448), .A2(n9447), .ZN(n14309) );
  NAND2_X1 U7361 ( .A1(n9971), .A2(n9970), .ZN(n14599) );
  NAND2_X1 U7362 ( .A1(n12369), .A2(n7657), .ZN(n14268) );
  AND2_X1 U7363 ( .A1(n9337), .A2(n9336), .ZN(n14134) );
  NAND2_X1 U7364 ( .A1(n15444), .A2(n10323), .ZN(n15108) );
  NAND2_X1 U7365 ( .A1(n13303), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n13323) );
  NAND2_X1 U7366 ( .A1(n10123), .A2(n10122), .ZN(n12218) );
  XNOR2_X1 U7367 ( .A(n13322), .B(n13332), .ZN(n13303) );
  NAND2_X1 U7368 ( .A1(n13220), .A2(n12988), .ZN(n13120) );
  NAND2_X1 U7369 ( .A1(n13539), .A2(n13538), .ZN(n13537) );
  OAI21_X2 U7370 ( .B1(n11975), .B2(n9395), .A(n9216), .ZN(n14228) );
  NAND2_X1 U7371 ( .A1(n11729), .A2(n11730), .ZN(n10121) );
  AND2_X1 U7372 ( .A1(n7609), .A2(n15687), .ZN(n15694) );
  AND2_X1 U7373 ( .A1(n9183), .A2(n9182), .ZN(n16030) );
  OAI22_X1 U7374 ( .A1(n12185), .A2(n12184), .B1(n12183), .B2(n12182), .ZN(
        n12186) );
  AOI21_X1 U7375 ( .B1(n7721), .B2(n7204), .A(n7719), .ZN(n8981) );
  NAND2_X1 U7376 ( .A1(n9817), .A2(n9816), .ZN(n14561) );
  INV_X1 U7377 ( .A(n8935), .ZN(n7721) );
  INV_X1 U7378 ( .A(n10154), .ZN(n8022) );
  NAND2_X1 U7379 ( .A1(n9744), .A2(n9743), .ZN(n12760) );
  OAI21_X1 U7380 ( .B1(n9134), .B2(n7520), .A(n7517), .ZN(n9204) );
  OAI22_X1 U7381 ( .A1(n15791), .A2(n15790), .B1(n11798), .B2(n11830), .ZN(
        n15812) );
  NAND2_X1 U7382 ( .A1(n9773), .A2(n9772), .ZN(n12773) );
  AOI22_X1 U7383 ( .A1(n15770), .A2(n15769), .B1(n15780), .B2(n11796), .ZN(
        n15791) );
  NAND2_X1 U7384 ( .A1(n9758), .A2(n9757), .ZN(n12764) );
  NAND2_X1 U7385 ( .A1(n9086), .A2(n8077), .ZN(n9112) );
  NAND2_X1 U7386 ( .A1(n7340), .A2(n11794), .ZN(n15770) );
  INV_X1 U7387 ( .A(n10783), .ZN(n10256) );
  NAND2_X1 U7388 ( .A1(n9731), .A2(n9730), .ZN(n12753) );
  NAND2_X1 U7389 ( .A1(n9010), .A2(n9009), .ZN(n9031) );
  AOI21_X2 U7390 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(n15646), .A(n15645), .ZN(
        n15653) );
  NAND2_X1 U7391 ( .A1(n9702), .A2(n9701), .ZN(n12741) );
  AND2_X2 U7392 ( .A1(n8902), .A2(n8901), .ZN(n11535) );
  OR2_X1 U7393 ( .A1(n8863), .A2(n8864), .ZN(n7774) );
  XNOR2_X1 U7394 ( .A(n12723), .B(n14741), .ZN(n12876) );
  AND2_X1 U7395 ( .A1(n15627), .A2(n15626), .ZN(n15628) );
  NAND2_X1 U7396 ( .A1(n9664), .A2(n9663), .ZN(n12723) );
  CLKBUF_X3 U7397 ( .A(n12986), .Z(n13053) );
  NAND2_X2 U7398 ( .A1(n14837), .A2(n15051), .ZN(n15054) );
  XNOR2_X1 U7399 ( .A(n14743), .B(n15835), .ZN(n11151) );
  OR2_X1 U7400 ( .A1(n15608), .A2(n15607), .ZN(n7613) );
  CLKBUF_X2 U7401 ( .A(n10784), .Z(n13805) );
  NAND2_X1 U7402 ( .A1(n9651), .A2(n9650), .ZN(n15835) );
  NAND2_X1 U7403 ( .A1(n8862), .A2(n8861), .ZN(n13929) );
  INV_X1 U7404 ( .A(n14742), .ZN(n7903) );
  AND2_X1 U7405 ( .A1(n7614), .A2(n7254), .ZN(n15608) );
  OR2_X1 U7406 ( .A1(n15598), .A2(n15599), .ZN(n7614) );
  NAND2_X1 U7407 ( .A1(n9639), .A2(n9638), .ZN(n14743) );
  OAI211_X1 U7408 ( .C1(n9665), .C2(n10574), .A(n7240), .B(n9656), .ZN(n10632)
         );
  BUF_X2 U7409 ( .A(n8897), .Z(n9468) );
  NAND2_X2 U7410 ( .A1(n8187), .A2(n13721), .ZN(n8240) );
  INV_X1 U7411 ( .A(n9899), .ZN(n9988) );
  AND2_X1 U7412 ( .A1(n8777), .A2(n10183), .ZN(n11242) );
  XNOR2_X1 U7413 ( .A(n8682), .B(n8681), .ZN(n12194) );
  INV_X1 U7414 ( .A(n9653), .ZN(n9899) );
  INV_X2 U7415 ( .A(n9665), .ZN(n10336) );
  INV_X1 U7416 ( .A(n8186), .ZN(n13721) );
  NAND2_X1 U7417 ( .A1(n7436), .A2(n7431), .ZN(n15443) );
  NAND2_X1 U7418 ( .A1(n10004), .A2(n10084), .ZN(n12704) );
  NAND2_X1 U7419 ( .A1(n8488), .A2(n8598), .ZN(n13361) );
  INV_X1 U7420 ( .A(n12484), .ZN(n7544) );
  XNOR2_X1 U7421 ( .A(n8611), .B(n8610), .ZN(n11367) );
  XNOR2_X1 U7422 ( .A(n10008), .B(n10007), .ZN(n15827) );
  MUX2_X1 U7423 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10003), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n10004) );
  AND2_X2 U7424 ( .A1(n9610), .A2(n12957), .ZN(n9985) );
  NAND2_X1 U7425 ( .A1(n9525), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8778) );
  NAND2_X1 U7426 ( .A1(n7503), .A2(n7501), .ZN(n8785) );
  NAND2_X1 U7427 ( .A1(n8759), .A2(n8760), .ZN(n10443) );
  NAND2_X1 U7428 ( .A1(n7300), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8185) );
  NAND2_X1 U7429 ( .A1(n7360), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8150) );
  NAND2_X1 U7430 ( .A1(n7963), .A2(n7962), .ZN(n15432) );
  NAND2_X2 U7431 ( .A1(n10297), .A2(P1_U3086), .ZN(n15435) );
  NAND2_X2 U7432 ( .A1(n10297), .A2(P3_U3151), .ZN(n13723) );
  AND2_X1 U7433 ( .A1(n9998), .A2(n8093), .ZN(n10005) );
  NOR2_X1 U7434 ( .A1(n8471), .A2(n7716), .ZN(n7524) );
  OAI21_X1 U7435 ( .B1(n10060), .B2(P1_IR_REG_18__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9881) );
  NAND2_X1 U7436 ( .A1(n8761), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8762) );
  NAND2_X1 U7437 ( .A1(n9826), .A2(n7175), .ZN(n10060) );
  AND2_X1 U7438 ( .A1(n8004), .A2(n7266), .ZN(n7558) );
  AND2_X1 U7439 ( .A1(n9826), .A2(n9598), .ZN(n9998) );
  INV_X1 U7440 ( .A(n8005), .ZN(n8004) );
  AND2_X1 U7441 ( .A1(n8095), .A2(n8748), .ZN(n7593) );
  XNOR2_X1 U7442 ( .A(n8235), .B(n8234), .ZN(n11274) );
  AND3_X1 U7443 ( .A1(n8874), .A2(n8745), .A3(n8744), .ZN(n8095) );
  AND4_X1 U7444 ( .A1(n8377), .A2(n8440), .A3(n8427), .A4(n8345), .ZN(n8145)
         );
  NAND2_X1 U7445 ( .A1(n8757), .A2(n7592), .ZN(n8013) );
  AND2_X1 U7446 ( .A1(n8210), .A2(n7467), .ZN(n7466) );
  AND4_X1 U7447 ( .A1(n9593), .A2(n9592), .A3(n9591), .A4(n9590), .ZN(n9594)
         );
  AND3_X1 U7448 ( .A1(n9585), .A2(n9584), .A3(n9583), .ZN(n10061) );
  INV_X1 U7449 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9526) );
  NOR2_X1 U7450 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n9584) );
  NOR2_X1 U7451 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n9585) );
  INV_X1 U7452 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8377) );
  NOR2_X1 U7453 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n9583) );
  INV_X1 U7454 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8140) );
  INV_X1 U7455 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8297) );
  INV_X1 U7456 ( .A(P1_RD_REG_SCAN_IN), .ZN(n8154) );
  INV_X1 U7457 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8278) );
  INV_X1 U7458 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8282) );
  NOR2_X2 U7459 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n8210) );
  INV_X4 U7460 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7461 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8345) );
  NOR2_X1 U7462 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n9588) );
  NOR2_X1 U7463 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n7416) );
  NOR2_X1 U7464 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n7467) );
  INV_X1 U7465 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8678) );
  INV_X1 U7466 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8767) );
  INV_X1 U7467 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8764) );
  INV_X1 U7468 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8427) );
  INV_X1 U7469 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8607) );
  INV_X1 U7470 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8440) );
  INV_X1 U7471 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8610) );
  INV_X4 U7472 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X1 U7473 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8743) );
  INV_X1 U7474 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8602) );
  NOR2_X1 U7475 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n8741) );
  NOR2_X1 U7476 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n8742) );
  NAND2_X1 U7477 ( .A1(n10702), .A2(n10110), .ZN(n10743) );
  NAND2_X1 U7478 ( .A1(n10704), .A2(n10703), .ZN(n10702) );
  NAND2_X2 U7479 ( .A1(n7643), .A2(n10118), .ZN(n11587) );
  NAND2_X1 U7480 ( .A1(n11403), .A2(n8025), .ZN(n7643) );
  NAND3_X2 U7481 ( .A1(n14666), .A2(n14664), .A3(n14665), .ZN(n14663) );
  INV_X1 U7482 ( .A(n8664), .ZN(n12695) );
  NOR2_X2 U7483 ( .A1(n13863), .A2(n13756), .ZN(n13757) );
  NOR2_X2 U7484 ( .A1(n12966), .A2(n7278), .ZN(n13198) );
  NOR2_X2 U7485 ( .A1(n12427), .A2(n12428), .ZN(n12966) );
  AND3_X2 U7486 ( .A1(n8798), .A2(n8795), .A3(n8796), .ZN(n7194) );
  NOR2_X2 U7487 ( .A1(n14117), .A2(n14314), .ZN(n14102) );
  NAND2_X1 U7488 ( .A1(n9611), .A2(n9612), .ZN(n9653) );
  INV_X1 U7489 ( .A(n9266), .ZN(n7756) );
  NAND2_X1 U7490 ( .A1(n7756), .A2(n7757), .ZN(n7753) );
  NAND2_X1 U7491 ( .A1(n9112), .A2(n7223), .ZN(n9134) );
  INV_X1 U7492 ( .A(n9129), .ZN(n8079) );
  AND2_X1 U7493 ( .A1(n8186), .A2(n13725), .ZN(n8215) );
  NAND2_X1 U7494 ( .A1(n13725), .A2(n13721), .ZN(n8242) );
  INV_X1 U7495 ( .A(n8126), .ZN(n7691) );
  INV_X1 U7496 ( .A(n7690), .ZN(n7689) );
  OAI21_X1 U7497 ( .B1(n8412), .B2(n7691), .A(n8425), .ZN(n7690) );
  OAI21_X1 U7498 ( .B1(n9367), .B2(n9366), .A(n9368), .ZN(n9441) );
  INV_X1 U7499 ( .A(n8224), .ZN(n8597) );
  INV_X1 U7500 ( .A(n8240), .ZN(n8665) );
  NAND2_X1 U7501 ( .A1(n8785), .A2(n12484), .ZN(n9145) );
  AND2_X1 U7502 ( .A1(n14309), .A2(n13912), .ZN(n7644) );
  NAND2_X1 U7503 ( .A1(n14203), .A2(n7556), .ZN(n7653) );
  NOR2_X1 U7504 ( .A1(n7161), .A2(n7557), .ZN(n7556) );
  INV_X1 U7505 ( .A(n14206), .ZN(n7557) );
  INV_X1 U7506 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9590) );
  NAND2_X1 U7507 ( .A1(n7510), .A2(n7508), .ZN(n9086) );
  AOI21_X1 U7508 ( .B1(n7511), .B2(n7512), .A(n7509), .ZN(n7508) );
  INV_X1 U7509 ( .A(n9081), .ZN(n7509) );
  AOI21_X1 U7510 ( .B1(n7426), .B2(n12799), .A(n7427), .ZN(n7425) );
  INV_X1 U7511 ( .A(n12798), .ZN(n7427) );
  INV_X1 U7512 ( .A(n7868), .ZN(n7426) );
  NAND2_X1 U7513 ( .A1(n7534), .A2(n13558), .ZN(n7533) );
  NAND2_X1 U7514 ( .A1(n12597), .A2(n12596), .ZN(n7534) );
  AND2_X1 U7515 ( .A1(n7752), .A2(n7755), .ZN(n7751) );
  NAND2_X1 U7516 ( .A1(n7754), .A2(n7753), .ZN(n7752) );
  OR2_X1 U7517 ( .A1(n7747), .A2(n7201), .ZN(n7746) );
  NAND2_X1 U7518 ( .A1(n8085), .A2(n9176), .ZN(n8084) );
  INV_X1 U7519 ( .A(n9199), .ZN(n8085) );
  NAND2_X1 U7520 ( .A1(n7349), .A2(n11326), .ZN(n12533) );
  NAND2_X1 U7521 ( .A1(n7591), .A2(n8004), .ZN(n7590) );
  AND4_X1 U7522 ( .A1(n8746), .A2(n7593), .A3(n8749), .A4(n7592), .ZN(n7591)
         );
  NOR2_X1 U7523 ( .A1(n9061), .A2(n7514), .ZN(n7513) );
  INV_X1 U7524 ( .A(n9030), .ZN(n7514) );
  NAND2_X1 U7525 ( .A1(n12991), .A2(n13524), .ZN(n7884) );
  NOR2_X1 U7526 ( .A1(n12119), .A2(n12118), .ZN(n12120) );
  OR2_X1 U7527 ( .A1(n13514), .A2(n13525), .ZN(n12621) );
  OR2_X1 U7528 ( .A1(n13636), .A2(n13536), .ZN(n12611) );
  INV_X1 U7529 ( .A(n11367), .ZN(n12536) );
  NAND2_X1 U7530 ( .A1(n13518), .A2(n13522), .ZN(n7636) );
  AOI21_X1 U7531 ( .B1(n7631), .B2(n12576), .A(n7243), .ZN(n7629) );
  INV_X1 U7532 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8146) );
  INV_X1 U7533 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7894) );
  NAND2_X1 U7534 ( .A1(n7679), .A2(n7677), .ZN(n8122) );
  NAND2_X1 U7535 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n7678), .ZN(n7677) );
  NAND2_X1 U7536 ( .A1(n8389), .A2(n8388), .ZN(n7679) );
  INV_X1 U7537 ( .A(n8116), .ZN(n7560) );
  INV_X1 U7538 ( .A(n11383), .ZN(n8002) );
  NOR2_X1 U7540 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n9179) );
  NOR2_X1 U7541 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n8771) );
  OR2_X1 U7542 ( .A1(n14305), .A2(n13778), .ZN(n10179) );
  INV_X1 U7543 ( .A(n7200), .ZN(n8032) );
  AOI21_X1 U7544 ( .B1(n10167), .B2(n8010), .A(n8008), .ZN(n14207) );
  AND2_X1 U7545 ( .A1(n10169), .A2(n7197), .ZN(n8010) );
  OAI21_X1 U7546 ( .B1(n8009), .B2(n7166), .A(n7239), .ZN(n8008) );
  OR2_X1 U7547 ( .A1(n12200), .A2(n12144), .ZN(n10159) );
  NAND2_X1 U7548 ( .A1(n7491), .A2(n7490), .ZN(n8006) );
  INV_X1 U7549 ( .A(n11731), .ZN(n7491) );
  INV_X1 U7550 ( .A(n7497), .ZN(n7496) );
  OAI21_X1 U7551 ( .B1(n7184), .B2(n10150), .A(n10152), .ZN(n7497) );
  OAI21_X1 U7552 ( .B1(n10204), .B2(n10203), .A(n15450), .ZN(n10259) );
  OR2_X1 U7553 ( .A1(n9525), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n9534) );
  AND2_X1 U7554 ( .A1(n10622), .A2(n7786), .ZN(n10624) );
  NOR2_X1 U7555 ( .A1(n12710), .A2(n7785), .ZN(n7784) );
  NAND2_X1 U7556 ( .A1(n7430), .A2(n7429), .ZN(n7428) );
  INV_X1 U7557 ( .A(n12705), .ZN(n7430) );
  INV_X1 U7558 ( .A(n10039), .ZN(n7955) );
  NOR2_X1 U7559 ( .A1(n15100), .A2(n7670), .ZN(n7669) );
  INV_X1 U7560 ( .A(n15108), .ZN(n7670) );
  INV_X1 U7561 ( .A(n14961), .ZN(n9905) );
  NAND2_X1 U7562 ( .A1(n15443), .A2(n14816), .ZN(n12702) );
  NAND2_X1 U7563 ( .A1(n9349), .A2(n9348), .ZN(n9367) );
  NAND2_X1 U7564 ( .A1(n9228), .A2(n9227), .ZN(n9253) );
  AOI22_X1 U7565 ( .A1(n15663), .A2(n15662), .B1(P1_ADDR_REG_11__SCAN_IN), 
        .B2(n15661), .ZN(n15666) );
  INV_X1 U7566 ( .A(n11430), .ZN(n12986) );
  AND2_X1 U7567 ( .A1(n12645), .A2(n12644), .ZN(n12682) );
  INV_X1 U7568 ( .A(n8242), .ZN(n8506) );
  AND2_X1 U7569 ( .A1(n13401), .A2(n8661), .ZN(n9569) );
  AND2_X1 U7570 ( .A1(n8572), .A2(n8571), .ZN(n13437) );
  AOI21_X1 U7571 ( .B1(n7169), .B2(n7708), .A(n7271), .ZN(n7705) );
  OAI22_X1 U7572 ( .A1(n13533), .A2(n13538), .B1(n13524), .B2(n13700), .ZN(
        n13521) );
  NAND2_X1 U7573 ( .A1(n13537), .A2(n12609), .ZN(n13518) );
  AND2_X1 U7574 ( .A1(n12611), .A2(n12608), .ZN(n13522) );
  NAND2_X1 U7575 ( .A1(n7469), .A2(n7468), .ZN(n13583) );
  AOI21_X1 U7576 ( .B1(n7471), .B2(n7473), .A(n7179), .ZN(n7468) );
  INV_X1 U7577 ( .A(n7626), .ZN(n7473) );
  AOI21_X1 U7578 ( .B1(n12661), .B2(n7459), .A(n7458), .ZN(n7457) );
  INV_X1 U7579 ( .A(n12556), .ZN(n7459) );
  INV_X1 U7580 ( .A(n12560), .ZN(n7458) );
  AND2_X1 U7581 ( .A1(n11852), .A2(n8625), .ZN(n11905) );
  OR2_X1 U7582 ( .A1(n8289), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8304) );
  NAND2_X1 U7583 ( .A1(n10850), .A2(n10297), .ZN(n8229) );
  AND4_X1 U7584 ( .A1(n8207), .A2(n8206), .A3(n8205), .A4(n8204), .ZN(n11334)
         );
  OR2_X1 U7585 ( .A1(n8495), .A2(n10884), .ZN(n8206) );
  NAND3_X1 U7586 ( .A1(n10850), .A2(n10868), .A3(n12641), .ZN(n13582) );
  INV_X1 U7587 ( .A(n12510), .ZN(n8490) );
  INV_X1 U7588 ( .A(n10850), .ZN(n8489) );
  OR3_X1 U7589 ( .A1(n13709), .A2(n13711), .A3(n8732), .ZN(n11111) );
  AND2_X1 U7590 ( .A1(n11092), .A2(n13710), .ZN(n11109) );
  INV_X1 U7591 ( .A(n15846), .ZN(n13580) );
  NAND2_X1 U7592 ( .A1(n13715), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8183) );
  NAND2_X1 U7593 ( .A1(n7367), .A2(n8135), .ZN(n8194) );
  NAND2_X1 U7594 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n8134), .ZN(n8135) );
  NAND2_X1 U7595 ( .A1(n8576), .A2(n8574), .ZN(n7367) );
  OAI21_X1 U7596 ( .B1(P2_DATAO_REG_21__SCAN_IN), .B2(n12359), .A(n8132), .ZN(
        n8521) );
  NAND2_X1 U7597 ( .A1(n8512), .A2(n8510), .ZN(n8132) );
  NAND2_X1 U7598 ( .A1(n7559), .A2(n7696), .ZN(n8486) );
  NAND2_X1 U7599 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n7697), .ZN(n7696) );
  NAND2_X1 U7600 ( .A1(n8470), .A2(n8468), .ZN(n7559) );
  INV_X1 U7601 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7697) );
  INV_X1 U7602 ( .A(n7409), .ZN(n7408) );
  OAI21_X1 U7603 ( .B1(n7686), .B2(n7288), .A(n8127), .ZN(n7409) );
  INV_X1 U7604 ( .A(n13738), .ZN(n7971) );
  OAI21_X1 U7605 ( .B1(n7972), .B2(n7193), .A(n12057), .ZN(n12058) );
  OR2_X1 U7606 ( .A1(n9355), .A2(n13830), .ZN(n9471) );
  AND2_X1 U7607 ( .A1(n9521), .A2(n7734), .ZN(n7733) );
  NAND2_X1 U7608 ( .A1(n9494), .A2(n7735), .ZN(n7734) );
  OR2_X1 U7609 ( .A1(n9520), .A2(n9519), .ZN(n9521) );
  OAI22_X1 U7610 ( .A1(n9488), .A2(n9487), .B1(n9363), .B2(n9364), .ZN(n7735)
         );
  INV_X1 U7611 ( .A(n8786), .ZN(n9478) );
  INV_X1 U7612 ( .A(n13911), .ZN(n13778) );
  OR2_X1 U7613 ( .A1(n7482), .A2(n7489), .ZN(n7478) );
  AND2_X1 U7614 ( .A1(n7481), .A2(n14071), .ZN(n7480) );
  NOR2_X1 U7615 ( .A1(n14331), .A2(n13868), .ZN(n8035) );
  AND2_X1 U7616 ( .A1(n7652), .A2(n7654), .ZN(n7651) );
  INV_X1 U7617 ( .A(n14175), .ZN(n7652) );
  NAND2_X1 U7618 ( .A1(n14269), .A2(n14270), .ZN(n10167) );
  NOR2_X1 U7619 ( .A1(n14270), .A2(n7658), .ZN(n7657) );
  INV_X1 U7620 ( .A(n10127), .ZN(n7658) );
  NAND2_X1 U7621 ( .A1(n10712), .A2(n10109), .ZN(n10704) );
  NAND2_X1 U7622 ( .A1(n8802), .A2(n10276), .ZN(n9040) );
  OR2_X1 U7623 ( .A1(n13911), .A2(n14305), .ZN(n7366) );
  BUF_X1 U7624 ( .A(n8849), .Z(n9229) );
  INV_X1 U7625 ( .A(n8802), .ZN(n8849) );
  OR2_X1 U7626 ( .A1(n8758), .A2(n7504), .ZN(n7503) );
  NAND2_X1 U7627 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n7505), .ZN(n7504) );
  AND2_X1 U7628 ( .A1(n10727), .A2(n10730), .ZN(n7820) );
  INV_X1 U7629 ( .A(n11765), .ZN(n7808) );
  NAND2_X1 U7630 ( .A1(n7160), .A2(n7781), .ZN(n7780) );
  INV_X1 U7631 ( .A(n12299), .ZN(n7781) );
  AOI21_X1 U7632 ( .B1(n7802), .B2(n7804), .A(n7245), .ZN(n7801) );
  INV_X1 U7633 ( .A(n14678), .ZN(n7802) );
  NAND2_X1 U7634 ( .A1(n12957), .A2(n9612), .ZN(n9679) );
  AOI21_X1 U7635 ( .B1(n7960), .B2(n12902), .A(n7958), .ZN(n7957) );
  INV_X1 U7636 ( .A(n7960), .ZN(n7959) );
  OR2_X1 U7637 ( .A1(n14892), .A2(n15079), .ZN(n14878) );
  NAND2_X1 U7638 ( .A1(n14958), .A2(n10034), .ZN(n14946) );
  INV_X1 U7639 ( .A(n11163), .ZN(n9659) );
  OR2_X1 U7640 ( .A1(n9392), .A2(n9391), .ZN(n9394) );
  AND2_X1 U7641 ( .A1(n9597), .A2(n9596), .ZN(n9599) );
  INV_X1 U7642 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9609) );
  NAND2_X1 U7643 ( .A1(n9207), .A2(n9208), .ZN(n9228) );
  NOR2_X1 U7644 ( .A1(n9088), .A2(n8078), .ZN(n8077) );
  INV_X1 U7645 ( .A(n9085), .ZN(n8078) );
  AND2_X1 U7646 ( .A1(n9589), .A2(n9671), .ZN(n7417) );
  OR2_X1 U7647 ( .A1(n11997), .A2(n12242), .ZN(n11998) );
  AOI21_X1 U7648 ( .B1(n13388), .B2(n8597), .A(n8596), .ZN(n13397) );
  NAND2_X1 U7649 ( .A1(n13827), .A2(n13826), .ZN(n13825) );
  INV_X1 U7650 ( .A(n15407), .ZN(n14686) );
  OR2_X1 U7651 ( .A1(n8933), .A2(n8934), .ZN(n7728) );
  AND2_X1 U7652 ( .A1(n7728), .A2(n8957), .ZN(n7726) );
  OAI22_X1 U7653 ( .A1(n7852), .A2(n7851), .B1(n12751), .B2(n7850), .ZN(n12757) );
  INV_X1 U7654 ( .A(n12750), .ZN(n7850) );
  NOR2_X1 U7655 ( .A1(n12752), .A2(n12750), .ZN(n7851) );
  AOI22_X1 U7656 ( .A1(n7724), .A2(n7723), .B1(n7727), .B2(n7722), .ZN(n7720)
         );
  INV_X1 U7657 ( .A(n7728), .ZN(n7722) );
  INV_X1 U7658 ( .A(n7726), .ZN(n7723) );
  OR2_X1 U7659 ( .A1(n12757), .A2(n12756), .ZN(n12758) );
  INV_X1 U7660 ( .A(n9004), .ZN(n7768) );
  OAI21_X1 U7661 ( .B1(n7539), .B2(n12573), .A(n12572), .ZN(n7538) );
  AOI21_X1 U7662 ( .B1(n12564), .B2(n12563), .A(n12562), .ZN(n7539) );
  AND2_X1 U7663 ( .A1(n7632), .A2(n12641), .ZN(n7535) );
  INV_X1 U7664 ( .A(n9127), .ZN(n7772) );
  INV_X1 U7665 ( .A(n9128), .ZN(n7771) );
  NAND2_X1 U7666 ( .A1(n12801), .A2(n12803), .ZN(n7871) );
  NOR2_X1 U7667 ( .A1(n7224), .A2(n7425), .ZN(n7424) );
  INV_X1 U7668 ( .A(n9173), .ZN(n7763) );
  NOR2_X1 U7669 ( .A1(n7440), .A2(n7222), .ZN(n7439) );
  INV_X1 U7670 ( .A(n9196), .ZN(n7760) );
  NAND2_X1 U7671 ( .A1(n7763), .A2(n7764), .ZN(n7761) );
  NOR2_X1 U7672 ( .A1(n7763), .A2(n7764), .ZN(n7762) );
  OAI21_X1 U7673 ( .B1(n7533), .B2(n7529), .A(n7528), .ZN(n7527) );
  INV_X1 U7674 ( .A(n12600), .ZN(n7529) );
  NOR2_X1 U7675 ( .A1(n12599), .A2(n12641), .ZN(n7528) );
  OAI21_X1 U7676 ( .B1(n7533), .B2(n7532), .A(n7531), .ZN(n7530) );
  INV_X1 U7677 ( .A(n12603), .ZN(n7532) );
  NOR2_X1 U7678 ( .A1(n12602), .A2(n12635), .ZN(n7531) );
  NOR2_X1 U7679 ( .A1(n12613), .A2(n12607), .ZN(n7526) );
  INV_X1 U7680 ( .A(n12822), .ZN(n7862) );
  NOR2_X1 U7681 ( .A1(n7756), .A2(n7757), .ZN(n7754) );
  AOI21_X1 U7682 ( .B1(n7751), .B2(n7749), .A(n7748), .ZN(n7747) );
  INV_X1 U7683 ( .A(n9282), .ZN(n7748) );
  INV_X1 U7684 ( .A(n7753), .ZN(n7749) );
  INV_X1 U7685 ( .A(n7751), .ZN(n7750) );
  NAND2_X1 U7686 ( .A1(n12841), .A2(n7847), .ZN(n7846) );
  INV_X1 U7687 ( .A(n12840), .ZN(n7847) );
  NAND2_X1 U7688 ( .A1(n7404), .A2(n7403), .ZN(n7402) );
  NOR2_X1 U7689 ( .A1(n12529), .A2(n12641), .ZN(n7403) );
  NAND2_X1 U7690 ( .A1(n12531), .A2(n12641), .ZN(n7685) );
  NOR2_X1 U7691 ( .A1(n13422), .A2(n8586), .ZN(n7573) );
  NAND2_X1 U7692 ( .A1(n14423), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7680) );
  NAND2_X1 U7693 ( .A1(n12703), .A2(n12702), .ZN(n12705) );
  NAND2_X1 U7694 ( .A1(n7281), .A2(n9251), .ZN(n8055) );
  NOR2_X1 U7695 ( .A1(n8084), .A2(n7522), .ZN(n7521) );
  INV_X1 U7696 ( .A(n9154), .ZN(n7522) );
  OAI21_X1 U7697 ( .B1(n8086), .B2(n8084), .A(n9203), .ZN(n8083) );
  NAND2_X1 U7698 ( .A1(n7521), .A2(n7519), .ZN(n7518) );
  INV_X1 U7699 ( .A(n9133), .ZN(n7519) );
  INV_X1 U7700 ( .A(n12986), .ZN(n13050) );
  AND2_X1 U7701 ( .A1(n13004), .A2(n13002), .ZN(n7853) );
  NAND2_X1 U7702 ( .A1(n12686), .A2(n11367), .ZN(n11309) );
  NOR2_X1 U7703 ( .A1(n15797), .A2(n7297), .ZN(n11831) );
  AND2_X1 U7704 ( .A1(n11830), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7297) );
  NAND2_X1 U7705 ( .A1(n12123), .A2(n12124), .ZN(n12173) );
  NAND2_X1 U7706 ( .A1(n13258), .A2(n13257), .ZN(n13286) );
  NAND2_X1 U7707 ( .A1(n13301), .A2(n13302), .ZN(n13322) );
  OR2_X1 U7708 ( .A1(n8515), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8524) );
  AND2_X1 U7709 ( .A1(n8214), .A2(n7354), .ZN(n11311) );
  OR2_X1 U7710 ( .A1(n8229), .A2(SI_2_), .ZN(n8214) );
  AND2_X1 U7711 ( .A1(n8213), .A2(n8212), .ZN(n7354) );
  NAND2_X1 U7712 ( .A1(n7635), .A2(n7634), .ZN(n7633) );
  INV_X1 U7713 ( .A(n12283), .ZN(n7635) );
  OAI21_X1 U7714 ( .B1(n7396), .B2(n7182), .A(P1_DATAO_REG_24__SCAN_IN), .ZN(
        n7390) );
  NOR2_X1 U7715 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n8144) );
  NOR2_X1 U7716 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), .ZN(
        n8143) );
  INV_X1 U7717 ( .A(n7375), .ZN(n7374) );
  OAI21_X1 U7718 ( .B1(n8361), .B2(n7185), .A(n8375), .ZN(n7375) );
  INV_X1 U7719 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n8120) );
  NAND2_X1 U7720 ( .A1(n7374), .A2(n7185), .ZN(n7372) );
  NOR2_X1 U7721 ( .A1(n7401), .A2(n7562), .ZN(n7400) );
  NOR2_X1 U7722 ( .A1(n7164), .A2(n7698), .ZN(n7401) );
  INV_X1 U7723 ( .A(n8210), .ZN(n10864) );
  NOR2_X1 U7724 ( .A1(n9290), .A2(n13869), .ZN(n7328) );
  NAND2_X1 U7725 ( .A1(n10236), .A2(n10235), .ZN(n10784) );
  NOR2_X1 U7726 ( .A1(n9233), .A2(n9232), .ZN(n7329) );
  AND2_X1 U7727 ( .A1(n8793), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8782) );
  NAND2_X1 U7728 ( .A1(n7488), .A2(n7487), .ZN(n7486) );
  AND2_X1 U7729 ( .A1(n14197), .A2(n10170), .ZN(n8042) );
  AOI21_X1 U7730 ( .B1(n10151), .B2(n7496), .A(n7494), .ZN(n7493) );
  NAND2_X1 U7731 ( .A1(n7495), .A2(n10153), .ZN(n7494) );
  NAND2_X1 U7732 ( .A1(n7496), .A2(n7184), .ZN(n7495) );
  AOI21_X1 U7733 ( .B1(n10153), .B2(n8025), .A(n8022), .ZN(n8021) );
  INV_X1 U7734 ( .A(n10746), .ZN(n10142) );
  INV_X1 U7735 ( .A(n14384), .ZN(n14119) );
  NAND2_X1 U7736 ( .A1(n7476), .A2(n10145), .ZN(n10966) );
  MUX2_X1 U7737 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8756), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n8760) );
  AND4_X1 U7738 ( .A1(n9179), .A2(n8771), .A3(n8773), .A4(n8764), .ZN(n8765)
         );
  NOR2_X2 U7739 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n9012) );
  INV_X1 U7740 ( .A(n7801), .ZN(n7799) );
  OR2_X1 U7741 ( .A1(n12899), .A2(n7923), .ZN(n7922) );
  INV_X1 U7742 ( .A(n9938), .ZN(n7923) );
  NOR2_X1 U7743 ( .A1(n12897), .A2(n7925), .ZN(n7924) );
  INV_X1 U7744 ( .A(n9928), .ZN(n7925) );
  NOR2_X1 U7745 ( .A1(n7913), .A2(n7911), .ZN(n7910) );
  INV_X1 U7746 ( .A(n9796), .ZN(n7911) );
  INV_X1 U7747 ( .A(n7914), .ZN(n7913) );
  NOR2_X1 U7748 ( .A1(n12071), .A2(n7915), .ZN(n7914) );
  INV_X1 U7749 ( .A(n9811), .ZN(n7915) );
  NOR2_X1 U7750 ( .A1(n15413), .A2(n7675), .ZN(n7674) );
  INV_X1 U7751 ( .A(n7676), .ZN(n7675) );
  INV_X1 U7752 ( .A(n12888), .ZN(n7929) );
  XNOR2_X1 U7753 ( .A(n12738), .B(n14739), .ZN(n12879) );
  NAND2_X1 U7754 ( .A1(n15888), .A2(n7903), .ZN(n10010) );
  AOI21_X2 U7755 ( .B1(n10021), .B2(n8104), .A(n8103), .ZN(n11510) );
  OR2_X1 U7756 ( .A1(n10064), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n10066) );
  INV_X1 U7757 ( .A(n8055), .ZN(n8053) );
  INV_X1 U7758 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9996) );
  OR2_X1 U7759 ( .A1(n9253), .A2(n9252), .ZN(n8060) );
  AND2_X1 U7760 ( .A1(n9598), .A2(n9996), .ZN(n7825) );
  NAND2_X1 U7761 ( .A1(n9087), .A2(SI_13_), .ZN(n9111) );
  AOI21_X1 U7762 ( .B1(n7513), .B2(n9008), .A(n7242), .ZN(n7511) );
  INV_X1 U7763 ( .A(n7513), .ZN(n7512) );
  NOR2_X1 U7764 ( .A1(n8936), .A2(n8893), .ZN(n8067) );
  INV_X1 U7765 ( .A(n8939), .ZN(n8069) );
  INV_X1 U7766 ( .A(n8825), .ZN(n7316) );
  NAND2_X1 U7767 ( .A1(n8046), .A2(n8809), .ZN(n8045) );
  NAND2_X1 U7768 ( .A1(n8806), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8803) );
  NOR2_X1 U7769 ( .A1(n15624), .A2(n15623), .ZN(n15634) );
  AOI21_X1 U7770 ( .B1(n7832), .B2(n7834), .A(n7830), .ZN(n7829) );
  INV_X1 U7771 ( .A(n13040), .ZN(n7830) );
  INV_X1 U7772 ( .A(n13121), .ZN(n7882) );
  INV_X1 U7773 ( .A(n13145), .ZN(n7841) );
  OR2_X1 U7774 ( .A1(n8493), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8504) );
  XNOR2_X1 U7775 ( .A(n11312), .B(n11326), .ZN(n11315) );
  NAND2_X1 U7776 ( .A1(n12992), .A2(n7881), .ZN(n7880) );
  INV_X1 U7777 ( .A(n12990), .ZN(n7881) );
  OR2_X1 U7778 ( .A1(n8461), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8477) );
  NAND2_X1 U7779 ( .A1(n11720), .A2(n11856), .ZN(n7307) );
  NAND2_X1 U7780 ( .A1(n7415), .A2(n7413), .ZN(n12646) );
  OAI21_X1 U7781 ( .B1(n12638), .B2(n7414), .A(n7229), .ZN(n7413) );
  NAND2_X1 U7782 ( .A1(n12642), .A2(n12635), .ZN(n7415) );
  INV_X1 U7783 ( .A(n12640), .ZN(n7414) );
  OR3_X1 U7784 ( .A1(n12194), .A2(n8690), .A3(n12262), .ZN(n11092) );
  AOI22_X1 U7785 ( .A1(n10879), .A2(n10863), .B1(n7331), .B2(
        P3_REG2_REG_0__SCAN_IN), .ZN(n11261) );
  NAND2_X1 U7786 ( .A1(n11261), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n11260) );
  NAND2_X1 U7787 ( .A1(n11024), .A2(n11023), .ZN(n11022) );
  INV_X1 U7788 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n15356) );
  AND2_X1 U7789 ( .A1(n7299), .A2(n7298), .ZN(n15797) );
  INV_X1 U7790 ( .A(n15798), .ZN(n7298) );
  NAND2_X1 U7791 ( .A1(n11818), .A2(n11817), .ZN(n12123) );
  OR2_X1 U7792 ( .A1(n7585), .A2(n12182), .ZN(n7584) );
  NAND2_X1 U7793 ( .A1(n7584), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7583) );
  NOR2_X1 U7794 ( .A1(n12120), .A2(n12131), .ZN(n12169) );
  NAND2_X1 U7795 ( .A1(n12176), .A2(n12177), .ZN(n13257) );
  NAND2_X1 U7796 ( .A1(n13259), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n13287) );
  NAND2_X1 U7797 ( .A1(n13291), .A2(n13290), .ZN(n13301) );
  OR2_X1 U7798 ( .A1(n13299), .A2(n7292), .ZN(n7578) );
  OR2_X1 U7799 ( .A1(n8580), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8592) );
  NAND2_X1 U7800 ( .A1(n9573), .A2(n7543), .ZN(n9574) );
  NOR2_X1 U7801 ( .A1(n13413), .A2(n12520), .ZN(n7624) );
  INV_X1 U7802 ( .A(n8651), .ZN(n7714) );
  AOI21_X1 U7803 ( .B1(n13434), .B2(n13435), .A(n8559), .ZN(n13428) );
  NAND2_X1 U7804 ( .A1(n13428), .A2(n13427), .ZN(n13426) );
  NAND2_X1 U7805 ( .A1(n13486), .A2(n13489), .ZN(n13488) );
  AND2_X1 U7806 ( .A1(n8090), .A2(n8644), .ZN(n7718) );
  AND3_X1 U7807 ( .A1(n8509), .A2(n8508), .A3(n8507), .ZN(n13505) );
  AND4_X1 U7808 ( .A1(n8451), .A2(n8450), .A3(n8449), .A4(n8448), .ZN(n13535)
         );
  NAND2_X1 U7809 ( .A1(n8173), .A2(n12179), .ZN(n8431) );
  AND2_X1 U7810 ( .A1(n13583), .A2(n12595), .ZN(n13569) );
  AND2_X1 U7811 ( .A1(n12594), .A2(n12595), .ZN(n13575) );
  INV_X1 U7812 ( .A(n13575), .ZN(n13586) );
  INV_X1 U7813 ( .A(n7472), .ZN(n7471) );
  OAI21_X1 U7814 ( .B1(n7474), .B2(n7473), .A(n13056), .ZN(n7472) );
  OR2_X1 U7815 ( .A1(n8381), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8405) );
  NOR2_X1 U7816 ( .A1(n7628), .A2(n12574), .ZN(n7474) );
  INV_X1 U7817 ( .A(n7629), .ZN(n7628) );
  AOI21_X1 U7818 ( .B1(n7629), .B2(n7630), .A(n7627), .ZN(n7626) );
  INV_X1 U7819 ( .A(n13054), .ZN(n7627) );
  NOR2_X1 U7820 ( .A1(n12575), .A2(n7638), .ZN(n7637) );
  INV_X1 U7821 ( .A(n8330), .ZN(n7638) );
  AND4_X1 U7822 ( .A1(n8410), .A2(n8409), .A3(n8408), .A4(n8407), .ZN(n13581)
         );
  AND3_X1 U7823 ( .A1(n8368), .A2(n8367), .A3(n8366), .ZN(n12422) );
  NAND2_X1 U7824 ( .A1(n8352), .A2(n12251), .ZN(n12283) );
  AND3_X1 U7825 ( .A1(n8351), .A2(n8350), .A3(n8349), .ZN(n12225) );
  OR2_X1 U7826 ( .A1(n8333), .A2(n8168), .ZN(n8354) );
  AND4_X1 U7827 ( .A1(n8360), .A2(n8359), .A3(n8358), .A4(n8357), .ZN(n12423)
         );
  NOR2_X1 U7828 ( .A1(n12664), .A2(n7712), .ZN(n7711) );
  INV_X1 U7829 ( .A(n8628), .ZN(n7712) );
  NAND2_X1 U7830 ( .A1(n12244), .A2(n12664), .ZN(n12243) );
  NAND2_X1 U7831 ( .A1(n11989), .A2(n12562), .ZN(n11988) );
  NAND2_X1 U7832 ( .A1(n7457), .A2(n8626), .ZN(n7456) );
  NOR2_X1 U7833 ( .A1(n12662), .A2(n7710), .ZN(n7709) );
  INV_X1 U7834 ( .A(n8624), .ZN(n7710) );
  NAND2_X1 U7835 ( .A1(n11665), .A2(n11664), .ZN(n11663) );
  AND4_X1 U7836 ( .A1(n8246), .A2(n8245), .A3(n8244), .A4(n8243), .ZN(n11662)
         );
  AND2_X1 U7837 ( .A1(n8712), .A2(n8616), .ZN(n15855) );
  AND2_X1 U7838 ( .A1(n8711), .A2(n8710), .ZN(n11189) );
  NAND2_X1 U7839 ( .A1(n12261), .A2(n12496), .ZN(n7565) );
  NAND2_X1 U7840 ( .A1(n8564), .A2(n8563), .ZN(n13105) );
  NAND2_X1 U7841 ( .A1(n8503), .A2(n8502), .ZN(n12999) );
  NAND2_X1 U7842 ( .A1(n7636), .A2(n7218), .ZN(n13631) );
  AND2_X1 U7843 ( .A1(n8380), .A2(n8379), .ZN(n13191) );
  CLKBUF_X1 U7844 ( .A(n8692), .Z(n8693) );
  OAI21_X1 U7845 ( .B1(P2_DATAO_REG_28__SCAN_IN), .B2(n14409), .A(n8137), .ZN(
        n12489) );
  INV_X1 U7846 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8184) );
  NOR2_X1 U7847 ( .A1(n7716), .A2(P3_IR_REG_27__SCAN_IN), .ZN(n7342) );
  INV_X1 U7848 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8149) );
  NAND2_X1 U7849 ( .A1(n8133), .A2(n7368), .ZN(n8576) );
  NAND2_X1 U7850 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n7369), .ZN(n7368) );
  INV_X1 U7851 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8681) );
  NAND2_X1 U7852 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n7682), .ZN(n7681) );
  CLKBUF_X1 U7853 ( .A(n8677), .Z(n8604) );
  AND2_X1 U7854 ( .A1(n7893), .A2(n8607), .ZN(n7891) );
  NAND2_X1 U7855 ( .A1(n7383), .A2(n8131), .ZN(n8512) );
  NAND2_X1 U7856 ( .A1(n7695), .A2(n7693), .ZN(n8130) );
  NAND2_X1 U7857 ( .A1(n7382), .A2(n7692), .ZN(n7381) );
  INV_X1 U7858 ( .A(n7693), .ZN(n7382) );
  NAND2_X1 U7859 ( .A1(n8486), .A2(n8484), .ZN(n7695) );
  NAND2_X1 U7860 ( .A1(n8129), .A2(n8128), .ZN(n8470) );
  AOI21_X1 U7861 ( .B1(n7408), .B2(n7288), .A(n7407), .ZN(n7406) );
  AOI21_X1 U7862 ( .B1(n7689), .B2(n7691), .A(n7279), .ZN(n7686) );
  OR2_X1 U7863 ( .A1(n8415), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n8439) );
  NAND2_X1 U7864 ( .A1(n8124), .A2(n8123), .ZN(n8413) );
  XNOR2_X1 U7865 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n8326) );
  XNOR2_X1 U7866 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n8311) );
  NAND2_X1 U7867 ( .A1(n7701), .A2(n8116), .ZN(n8313) );
  NAND2_X1 U7868 ( .A1(n7700), .A2(n7698), .ZN(n7701) );
  NAND2_X1 U7869 ( .A1(n7156), .A2(n8141), .ZN(n8314) );
  NAND2_X1 U7870 ( .A1(n8276), .A2(n8275), .ZN(n7700) );
  XNOR2_X1 U7871 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n8275) );
  AND2_X1 U7872 ( .A1(n8284), .A2(n8296), .ZN(n10978) );
  XNOR2_X1 U7873 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n8260) );
  XNOR2_X1 U7874 ( .A(n8262), .B(P3_IR_REG_4__SCAN_IN), .ZN(n10985) );
  XNOR2_X1 U7875 ( .A(n11938), .B(n13805), .ZN(n11946) );
  NAND2_X1 U7876 ( .A1(n11877), .A2(n11876), .ZN(n11878) );
  NAND2_X1 U7877 ( .A1(n11650), .A2(n11641), .ZN(n8001) );
  NAND2_X1 U7878 ( .A1(n8003), .A2(n8002), .ZN(n11642) );
  NAND2_X1 U7879 ( .A1(n7329), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n9275) );
  NAND2_X1 U7880 ( .A1(n12449), .A2(n12450), .ZN(n13732) );
  AND2_X1 U7881 ( .A1(n10783), .A2(n10782), .ZN(n10787) );
  OAI21_X1 U7882 ( .B1(n11382), .B2(n7999), .A(n7998), .ZN(n11743) );
  NAND2_X1 U7883 ( .A1(n8001), .A2(n11649), .ZN(n7998) );
  NAND2_X1 U7884 ( .A1(n11649), .A2(n8002), .ZN(n7999) );
  NAND2_X1 U7885 ( .A1(n7970), .A2(n13743), .ZN(n7523) );
  AOI21_X1 U7886 ( .B1(n7969), .B2(n7968), .A(n7967), .ZN(n7966) );
  INV_X1 U7887 ( .A(n13837), .ZN(n7968) );
  NAND2_X1 U7888 ( .A1(n13732), .A2(n13731), .ZN(n13836) );
  NAND2_X1 U7889 ( .A1(n10787), .A2(n10786), .ZN(n10823) );
  OR2_X1 U7890 ( .A1(n10825), .A2(n7982), .ZN(n7981) );
  INV_X1 U7891 ( .A(n11058), .ZN(n7982) );
  CLKBUF_X1 U7892 ( .A(n10823), .Z(n7335) );
  NAND2_X1 U7893 ( .A1(n12410), .A2(n7989), .ZN(n7988) );
  NAND2_X1 U7894 ( .A1(n9494), .A2(n7737), .ZN(n7736) );
  NAND2_X1 U7895 ( .A1(n9363), .A2(n9364), .ZN(n7737) );
  AND2_X1 U7896 ( .A1(n9361), .A2(n9360), .ZN(n13898) );
  AND3_X1 U7897 ( .A1(n9172), .A2(n9171), .A3(n9170), .ZN(n12441) );
  AND4_X1 U7898 ( .A1(n8956), .A2(n8955), .A3(n8954), .A4(n8953), .ZN(n11391)
         );
  NAND2_X1 U7899 ( .A1(n10179), .A2(n9546), .ZN(n14078) );
  OAI22_X1 U7900 ( .A1(n7327), .A2(n7485), .B1(n7486), .B2(n7483), .ZN(n7482)
         );
  INV_X1 U7901 ( .A(n7487), .ZN(n7485) );
  INV_X1 U7902 ( .A(n7486), .ZN(n7484) );
  INV_X1 U7903 ( .A(n14086), .ZN(n7327) );
  NAND2_X1 U7904 ( .A1(n14314), .A2(n13829), .ZN(n7488) );
  INV_X1 U7905 ( .A(n8028), .ZN(n8027) );
  OAI21_X1 U7906 ( .B1(n8032), .B2(n8030), .A(n8088), .ZN(n8028) );
  AOI21_X1 U7907 ( .B1(n8074), .B2(n8034), .A(n7232), .ZN(n8073) );
  INV_X1 U7908 ( .A(n10135), .ZN(n8074) );
  NAND2_X1 U7909 ( .A1(n8033), .A2(n8032), .ZN(n8029) );
  INV_X1 U7910 ( .A(n14141), .ZN(n8033) );
  NAND2_X1 U7911 ( .A1(n14166), .A2(n10134), .ZN(n14145) );
  INV_X1 U7912 ( .A(n8029), .ZN(n14140) );
  INV_X1 U7913 ( .A(n7655), .ZN(n7654) );
  OAI21_X1 U7914 ( .B1(n7161), .B2(n10131), .A(n10132), .ZN(n7655) );
  AND2_X1 U7915 ( .A1(n14175), .A2(n7205), .ZN(n8040) );
  NAND2_X1 U7916 ( .A1(n10171), .A2(n8042), .ZN(n8041) );
  NAND2_X1 U7917 ( .A1(n14207), .A2(n7498), .ZN(n10171) );
  NAND2_X1 U7918 ( .A1(n14220), .A2(n14238), .ZN(n7498) );
  NAND2_X1 U7919 ( .A1(n14225), .A2(n10130), .ZN(n14203) );
  NAND2_X1 U7920 ( .A1(n14203), .A2(n14206), .ZN(n14205) );
  INV_X1 U7921 ( .A(n10168), .ZN(n8011) );
  NAND2_X1 U7922 ( .A1(n10167), .A2(n7197), .ZN(n8007) );
  NAND2_X1 U7923 ( .A1(n14226), .A2(n14233), .ZN(n14225) );
  INV_X1 U7924 ( .A(n14403), .ZN(n14284) );
  NAND2_X1 U7925 ( .A1(n8020), .A2(n8019), .ZN(n14269) );
  NAND2_X1 U7926 ( .A1(n16020), .A2(n14273), .ZN(n8019) );
  NOR2_X1 U7927 ( .A1(n10165), .A2(n8015), .ZN(n8014) );
  NAND2_X1 U7928 ( .A1(n7554), .A2(n7553), .ZN(n12369) );
  INV_X1 U7929 ( .A(n12372), .ZN(n7553) );
  AND4_X1 U7930 ( .A1(n9101), .A2(n9100), .A3(n9099), .A4(n9098), .ZN(n12216)
         );
  AOI21_X1 U7931 ( .B1(n12012), .B2(n7649), .A(n7231), .ZN(n7648) );
  INV_X1 U7932 ( .A(n10120), .ZN(n7649) );
  NAND2_X1 U7933 ( .A1(n12015), .A2(n10159), .ZN(n12143) );
  INV_X1 U7934 ( .A(n7330), .ZN(n9067) );
  AND2_X1 U7935 ( .A1(n7546), .A2(n7255), .ZN(n7545) );
  OAI21_X1 U7936 ( .B1(n7492), .B2(n11779), .A(n10158), .ZN(n11731) );
  INV_X1 U7937 ( .A(n11778), .ZN(n7492) );
  AND4_X1 U7938 ( .A1(n8977), .A2(n8976), .A3(n8975), .A4(n8974), .ZN(n11644)
         );
  INV_X1 U7939 ( .A(n14275), .ZN(n14237) );
  INV_X1 U7940 ( .A(n14274), .ZN(n14235) );
  NAND2_X1 U7941 ( .A1(n11211), .A2(n7555), .ZN(n11340) );
  AND2_X1 U7942 ( .A1(n11346), .A2(n10116), .ZN(n7555) );
  NAND2_X1 U7943 ( .A1(n11212), .A2(n11214), .ZN(n11211) );
  NAND2_X1 U7944 ( .A1(n10742), .A2(n10111), .ZN(n10752) );
  XNOR2_X1 U7945 ( .A(n11415), .B(n13929), .ZN(n10746) );
  NAND2_X1 U7946 ( .A1(n10743), .A2(n10746), .ZN(n10742) );
  INV_X1 U7947 ( .A(n10305), .ZN(n7991) );
  INV_X1 U7948 ( .A(n14134), .ZN(n14326) );
  AND2_X1 U7949 ( .A1(n9231), .A2(n9230), .ZN(n14355) );
  OR2_X1 U7950 ( .A1(n10764), .A2(n9395), .ZN(n9094) );
  AND3_X1 U7951 ( .A1(n10259), .A2(n15448), .A3(n10207), .ZN(n10215) );
  NAND2_X1 U7952 ( .A1(n9537), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9541) );
  NAND2_X1 U7953 ( .A1(n9541), .A2(n9540), .ZN(n9543) );
  NAND3_X1 U7954 ( .A1(n10092), .A2(n10091), .A3(n10083), .ZN(n10583) );
  OR2_X1 U7955 ( .A1(n10624), .A2(n10623), .ZN(n10625) );
  INV_X1 U7956 ( .A(n12304), .ZN(n7782) );
  AND2_X1 U7957 ( .A1(n7791), .A2(n14615), .ZN(n7790) );
  OR2_X1 U7958 ( .A1(n7794), .A2(n7162), .ZN(n7791) );
  NAND2_X1 U7959 ( .A1(n14508), .A2(n7795), .ZN(n7793) );
  OAI21_X1 U7960 ( .B1(n10646), .B2(n7819), .A(n7818), .ZN(n10915) );
  AND2_X1 U7961 ( .A1(n7816), .A2(n10911), .ZN(n7818) );
  INV_X1 U7962 ( .A(n7807), .ZN(n7805) );
  AND2_X1 U7963 ( .A1(n11301), .A2(n11296), .ZN(n7823) );
  OAI21_X1 U7964 ( .B1(n14437), .B2(n7812), .A(n7809), .ZN(n14456) );
  AOI21_X1 U7965 ( .B1(n7813), .B2(n7811), .A(n7810), .ZN(n7809) );
  INV_X1 U7966 ( .A(n7813), .ZN(n7812) );
  INV_X1 U7967 ( .A(n14453), .ZN(n7810) );
  INV_X1 U7968 ( .A(n12851), .ZN(n7420) );
  NAND2_X1 U7969 ( .A1(n12942), .A2(n12916), .ZN(n12937) );
  INV_X1 U7970 ( .A(n12915), .ZN(n12916) );
  OAI21_X1 U7971 ( .B1(n12914), .B2(n12917), .A(n12941), .ZN(n12915) );
  CLKBUF_X1 U7972 ( .A(n9620), .Z(n10057) );
  NOR2_X1 U7973 ( .A1(n9665), .A2(n9632), .ZN(n9636) );
  OR2_X1 U7974 ( .A1(n10562), .A2(n10561), .ZN(n10601) );
  INV_X1 U7975 ( .A(n10043), .ZN(n14877) );
  NAND2_X1 U7976 ( .A1(n14925), .A2(n7924), .ZN(n14910) );
  AND2_X1 U7977 ( .A1(n14935), .A2(n9918), .ZN(n14927) );
  NAND2_X1 U7978 ( .A1(n14931), .A2(n10037), .ZN(n14916) );
  OR2_X1 U7979 ( .A1(n7934), .A2(n9917), .ZN(n7932) );
  AND2_X1 U7980 ( .A1(n14943), .A2(n9906), .ZN(n7934) );
  AND2_X1 U7981 ( .A1(n12896), .A2(n7935), .ZN(n7933) );
  NAND2_X1 U7982 ( .A1(n9905), .A2(n12896), .ZN(n14963) );
  INV_X1 U7983 ( .A(n7905), .ZN(n7904) );
  OAI21_X1 U7984 ( .B1(n7191), .B2(n7906), .A(n14978), .ZN(n7905) );
  INV_X1 U7985 ( .A(n9880), .ZN(n7906) );
  NAND2_X1 U7986 ( .A1(n15134), .A2(n7950), .ZN(n14974) );
  NOR2_X1 U7987 ( .A1(n14978), .A2(n7951), .ZN(n7950) );
  INV_X1 U7988 ( .A(n10031), .ZN(n7951) );
  NAND2_X1 U7989 ( .A1(n15011), .A2(n7191), .ZN(n14992) );
  NOR2_X1 U7990 ( .A1(n15142), .A2(n15035), .ZN(n15015) );
  AOI21_X1 U7991 ( .B1(n7949), .B2(n15042), .A(n7214), .ZN(n7947) );
  INV_X1 U7992 ( .A(n7949), .ZN(n7948) );
  NAND2_X1 U7993 ( .A1(n11865), .A2(n9796), .ZN(n11964) );
  NAND2_X1 U7994 ( .A1(n11964), .A2(n12891), .ZN(n11963) );
  AND2_X1 U7995 ( .A1(n12888), .A2(n10022), .ZN(n7946) );
  XNOR2_X1 U7996 ( .A(n12773), .B(n14733), .ZN(n12888) );
  NAND2_X1 U7997 ( .A1(n11509), .A2(n11511), .ZN(n11508) );
  NAND2_X1 U7998 ( .A1(n11499), .A2(n10810), .ZN(n11456) );
  AND2_X1 U7999 ( .A1(n7661), .A2(n12742), .ZN(n10810) );
  NAND2_X1 U8000 ( .A1(n10686), .A2(n10011), .ZN(n7942) );
  AOI21_X1 U8001 ( .B1(n9670), .B2(n7898), .A(n7228), .ZN(n7896) );
  INV_X1 U8002 ( .A(n7902), .ZN(n7898) );
  NAND2_X1 U8003 ( .A1(n7903), .A2(n15880), .ZN(n7902) );
  NAND2_X1 U8004 ( .A1(n9965), .A2(n9964), .ZN(n14870) );
  NAND2_X1 U8005 ( .A1(n9950), .A2(n9949), .ZN(n15079) );
  NAND2_X1 U8006 ( .A1(n9920), .A2(n9919), .ZN(n15100) );
  NAND2_X1 U8007 ( .A1(n9895), .A2(n9894), .ZN(n14967) );
  NAND2_X1 U8008 ( .A1(n9785), .A2(n9784), .ZN(n12777) );
  NAND2_X1 U8009 ( .A1(n11510), .A2(n12886), .ZN(n11559) );
  INV_X1 U8010 ( .A(n16013), .ZN(n15987) );
  NAND2_X1 U8011 ( .A1(n10583), .A2(n10586), .ZN(n15415) );
  NAND2_X1 U8012 ( .A1(n9375), .A2(n9374), .ZN(n9425) );
  OR2_X1 U8013 ( .A1(n9441), .A2(n9369), .ZN(n9375) );
  OR2_X1 U8014 ( .A1(n9604), .A2(n9603), .ZN(n7964) );
  NAND2_X1 U8015 ( .A1(n8050), .A2(n8051), .ZN(n9328) );
  AND2_X1 U8016 ( .A1(n8052), .A2(n8056), .ZN(n8051) );
  NAND2_X1 U8017 ( .A1(n9253), .A2(n8054), .ZN(n8050) );
  AOI21_X1 U8018 ( .B1(n8058), .B2(n9285), .A(n7181), .ZN(n8056) );
  OR2_X1 U8019 ( .A1(n9581), .A2(n9301), .ZN(n9303) );
  INV_X1 U8020 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9999) );
  INV_X1 U8021 ( .A(n10002), .ZN(n10001) );
  INV_X1 U8022 ( .A(n7433), .ZN(n7432) );
  OAI21_X1 U8023 ( .B1(n7435), .B2(P1_IR_REG_22__SCAN_IN), .A(n7434), .ZN(
        n7433) );
  NAND2_X1 U8024 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n7434) );
  NOR2_X1 U8025 ( .A1(n9999), .A2(n15420), .ZN(n7435) );
  XNOR2_X1 U8026 ( .A(n9328), .B(SI_22_), .ZN(n9581) );
  NAND2_X1 U8027 ( .A1(n10005), .A2(n10007), .ZN(n10002) );
  AND2_X1 U8028 ( .A1(n9227), .A2(n9206), .ZN(n9207) );
  NAND2_X1 U8029 ( .A1(n8081), .A2(n9176), .ZN(n9200) );
  NAND2_X1 U8030 ( .A1(n9826), .A2(n7825), .ZN(n10068) );
  NAND2_X1 U8031 ( .A1(n8061), .A2(n8063), .ZN(n9010) );
  AOI21_X1 U8032 ( .B1(n8988), .B2(n8065), .A(n8064), .ZN(n8063) );
  INV_X1 U8033 ( .A(n9005), .ZN(n8064) );
  NAND2_X1 U8034 ( .A1(n8985), .A2(n8984), .ZN(n8989) );
  NAND2_X1 U8035 ( .A1(n8960), .A2(n8959), .ZN(n8964) );
  INV_X1 U8036 ( .A(n8045), .ZN(n8044) );
  NAND2_X1 U8037 ( .A1(n8805), .A2(SI_1_), .ZN(n8822) );
  INV_X1 U8038 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n15604) );
  AOI21_X1 U8039 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(n15614), .A(n15734), .ZN(
        n15625) );
  OAI21_X1 U8040 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n15642), .A(n15641), .ZN(
        n15649) );
  NAND2_X1 U8041 ( .A1(n7616), .A2(n15660), .ZN(n15670) );
  OAI21_X1 U8042 ( .B1(n15659), .B2(n15658), .A(n7617), .ZN(n7616) );
  OAI21_X1 U8043 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n15669), .A(n15668), .ZN(
        n15680) );
  OAI21_X1 U8044 ( .B1(n15686), .B2(n15685), .A(n7610), .ZN(n7609) );
  AND4_X1 U8045 ( .A1(n8295), .A2(n8294), .A3(n8293), .A4(n8292), .ZN(n11918)
         );
  INV_X1 U8046 ( .A(n13247), .ZN(n12568) );
  NAND2_X1 U8047 ( .A1(n8535), .A2(n8534), .ZN(n13073) );
  AND4_X1 U8048 ( .A1(n8483), .A2(n8482), .A3(n8481), .A4(n8480), .ZN(n13536)
         );
  NAND2_X1 U8049 ( .A1(n8591), .A2(n8590), .ZN(n13033) );
  OR2_X1 U8050 ( .A1(n11329), .A2(n7449), .ZN(n7448) );
  AND2_X1 U8051 ( .A1(n13215), .A2(n7450), .ZN(n7449) );
  OR2_X1 U8052 ( .A1(n12987), .A2(n13551), .ZN(n12988) );
  INV_X1 U8053 ( .A(n13683), .ZN(n13186) );
  AND2_X1 U8054 ( .A1(n11318), .A2(n15848), .ZN(n13215) );
  AND4_X1 U8055 ( .A1(n8274), .A2(n8273), .A3(n8272), .A4(n8271), .ZN(n11724)
         );
  AND4_X1 U8056 ( .A1(n8310), .A2(n8309), .A3(n8308), .A4(n8307), .ZN(n12242)
         );
  NAND2_X1 U8057 ( .A1(n11108), .A2(n15860), .ZN(n13190) );
  NAND2_X1 U8058 ( .A1(n13211), .A2(n13213), .ZN(n13212) );
  AND2_X1 U8059 ( .A1(n11104), .A2(n11109), .ZN(n13223) );
  NAND2_X1 U8060 ( .A1(n12652), .A2(n7210), .ZN(n7410) );
  INV_X1 U8061 ( .A(n13505), .ZN(n13473) );
  INV_X1 U8062 ( .A(n12242), .ZN(n13248) );
  OR2_X1 U8063 ( .A1(n8240), .A2(n10877), .ZN(n8227) );
  NAND2_X1 U8064 ( .A1(n10944), .A2(n10896), .ZN(n10898) );
  INV_X1 U8065 ( .A(n7338), .ZN(n13255) );
  NAND2_X1 U8066 ( .A1(n7338), .A2(n7580), .ZN(n7579) );
  AND3_X1 U8067 ( .A1(n7579), .A2(P3_REG1_REG_15__SCAN_IN), .A3(n13273), .ZN(
        n13274) );
  NAND2_X1 U8068 ( .A1(n7577), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n13339) );
  INV_X1 U8069 ( .A(n13300), .ZN(n7577) );
  XNOR2_X1 U8070 ( .A(n7578), .B(n13318), .ZN(n13300) );
  OR2_X1 U8071 ( .A1(n10869), .A2(n12695), .ZN(n15800) );
  NOR2_X1 U8072 ( .A1(n8674), .A2(n8673), .ZN(n8675) );
  NOR2_X1 U8073 ( .A1(n13397), .A2(n13582), .ZN(n8674) );
  AND2_X1 U8074 ( .A1(n9572), .A2(n9571), .ZN(n13393) );
  OAI211_X1 U8075 ( .C1(n9569), .C2(n12678), .A(n9568), .B(n15851), .ZN(n9572)
         );
  AOI21_X1 U8076 ( .B1(n13599), .B2(n15977), .A(n7572), .ZN(n13404) );
  OR2_X1 U8077 ( .A1(n13402), .A2(n13403), .ZN(n7572) );
  AND2_X1 U8078 ( .A1(n11308), .A2(n12686), .ZN(n15861) );
  NAND2_X1 U8079 ( .A1(n16039), .A2(n15907), .ZN(n13656) );
  NOR2_X1 U8080 ( .A1(n13380), .A2(n7344), .ZN(n8739) );
  NOR2_X1 U8081 ( .A1(n7345), .A2(n13639), .ZN(n7344) );
  INV_X1 U8082 ( .A(n13385), .ZN(n7345) );
  INV_X1 U8083 ( .A(n13033), .ZN(n13597) );
  AND2_X1 U8084 ( .A1(n13404), .A2(n7571), .ZN(n13662) );
  NAND2_X1 U8085 ( .A1(n13599), .A2(n15857), .ZN(n7571) );
  NAND2_X1 U8086 ( .A1(n8460), .A2(n8459), .ZN(n13700) );
  INV_X1 U8087 ( .A(SI_12_), .ZN(n15172) );
  NAND2_X1 U8088 ( .A1(n7516), .A2(n7515), .ZN(n13777) );
  NAND2_X1 U8089 ( .A1(n7159), .A2(n7992), .ZN(n7515) );
  NAND2_X1 U8090 ( .A1(n12343), .A2(n12342), .ZN(n12344) );
  NOR2_X1 U8091 ( .A1(n12341), .A2(n7997), .ZN(n7996) );
  INV_X1 U8092 ( .A(n12100), .ZN(n7997) );
  XNOR2_X1 U8093 ( .A(n13757), .B(n8089), .ZN(n13786) );
  NAND2_X1 U8094 ( .A1(n13786), .A2(n13785), .ZN(n13784) );
  XNOR2_X1 U8095 ( .A(n10238), .B(n10237), .ZN(n10543) );
  AOI21_X1 U8096 ( .B1(n13853), .B2(n13750), .A(n13749), .ZN(n13816) );
  NAND2_X1 U8097 ( .A1(n13844), .A2(n13763), .ZN(n13827) );
  AND2_X1 U8098 ( .A1(n9192), .A2(n9191), .ZN(n14236) );
  INV_X1 U8099 ( .A(n7731), .ZN(n7730) );
  OAI21_X1 U8100 ( .B1(n7733), .B2(n10264), .A(n7172), .ZN(n7731) );
  NAND2_X1 U8101 ( .A1(n9436), .A2(n9435), .ZN(n13911) );
  NAND2_X1 U8102 ( .A1(n9459), .A2(n9458), .ZN(n13912) );
  INV_X1 U8103 ( .A(n12441), .ZN(n14249) );
  OR2_X1 U8104 ( .A1(n8794), .A2(n10456), .ZN(n8797) );
  NAND2_X1 U8105 ( .A1(n14418), .A2(n9467), .ZN(n8080) );
  NAND2_X1 U8106 ( .A1(n9273), .A2(n9272), .ZN(n14182) );
  NAND2_X1 U8107 ( .A1(n9387), .A2(n9386), .ZN(n14295) );
  NAND2_X1 U8108 ( .A1(n9397), .A2(n9396), .ZN(n14299) );
  NOR2_X1 U8109 ( .A1(n14056), .A2(n14062), .ZN(n7339) );
  AND2_X1 U8110 ( .A1(n10438), .A2(n9544), .ZN(n15455) );
  INV_X1 U8111 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n12960) );
  INV_X1 U8112 ( .A(n8013), .ZN(n8012) );
  NAND2_X1 U8113 ( .A1(n12154), .A2(n12153), .ZN(n12300) );
  NAND2_X1 U8114 ( .A1(n9884), .A2(n9883), .ZN(n14980) );
  AOI21_X1 U8115 ( .B1(n9646), .B2(n9645), .A(n9644), .ZN(n9651) );
  NAND2_X1 U8116 ( .A1(n9801), .A2(n9800), .ZN(n15983) );
  OR2_X1 U8117 ( .A1(n10764), .A2(n12853), .ZN(n9801) );
  INV_X1 U8118 ( .A(n14711), .ZN(n14690) );
  NAND4_X1 U8119 ( .A1(n9669), .A2(n9668), .A3(n9667), .A4(n9666), .ZN(n14741)
         );
  NAND4_X1 U8120 ( .A1(n9625), .A2(n9624), .A3(n9623), .A4(n9622), .ZN(n14742)
         );
  NAND2_X1 U8121 ( .A1(n12865), .A2(n12864), .ZN(n15064) );
  AND2_X1 U8122 ( .A1(n9984), .A2(n9983), .ZN(n14842) );
  NAND2_X1 U8123 ( .A1(n9908), .A2(n9907), .ZN(n15115) );
  AND2_X1 U8124 ( .A1(n7666), .A2(n7665), .ZN(n15160) );
  AOI21_X1 U8125 ( .B1(n15064), .B2(n15982), .A(n15063), .ZN(n7665) );
  OR2_X1 U8126 ( .A1(n16017), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n7663) );
  NAND2_X1 U8127 ( .A1(n12855), .A2(n12854), .ZN(n15382) );
  OR2_X1 U8128 ( .A1(n15427), .A2(n12853), .ZN(n12855) );
  INV_X1 U8129 ( .A(n14842), .ZN(n10099) );
  AND2_X1 U8130 ( .A1(n10226), .A2(n7918), .ZN(n10231) );
  AND2_X1 U8131 ( .A1(n10227), .A2(n7919), .ZN(n7918) );
  INV_X1 U8132 ( .A(n14848), .ZN(n10226) );
  NAND2_X1 U8133 ( .A1(n9871), .A2(n9870), .ZN(n15407) );
  AND2_X1 U8134 ( .A1(n9605), .A2(n9609), .ZN(n7889) );
  NAND2_X1 U8135 ( .A1(n15587), .A2(n15586), .ZN(n15596) );
  NAND2_X1 U8136 ( .A1(n7603), .A2(n7602), .ZN(n15633) );
  INV_X1 U8137 ( .A(n15629), .ZN(n7602) );
  INV_X1 U8138 ( .A(n15628), .ZN(n7603) );
  NOR2_X1 U8139 ( .A1(n15644), .A2(n15643), .ZN(n15645) );
  NAND2_X1 U8140 ( .A1(n7309), .A2(n15712), .ZN(n15713) );
  INV_X1 U8141 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7604) );
  NOR2_X1 U8142 ( .A1(n15714), .A2(n15713), .ZN(n15716) );
  INV_X1 U8143 ( .A(n12713), .ZN(n12714) );
  AOI21_X1 U8144 ( .B1(n12712), .B2(n12874), .A(n12711), .ZN(n12713) );
  OAI21_X1 U8145 ( .B1(n12710), .B2(n15835), .A(n12716), .ZN(n12711) );
  AND2_X1 U8146 ( .A1(n12718), .A2(n12717), .ZN(n12719) );
  NAND2_X1 U8147 ( .A1(n7828), .A2(n7827), .ZN(n12718) );
  AND2_X1 U8148 ( .A1(n10010), .A2(n10009), .ZN(n7828) );
  OR2_X1 U8149 ( .A1(n7856), .A2(n12740), .ZN(n7857) );
  NAND2_X1 U8150 ( .A1(n12740), .A2(n7856), .ZN(n7855) );
  INV_X1 U8151 ( .A(n8958), .ZN(n7725) );
  NOR2_X1 U8152 ( .A1(n7227), .A2(n8957), .ZN(n7727) );
  NAND2_X1 U8153 ( .A1(n12761), .A2(n12763), .ZN(n7859) );
  NOR2_X1 U8154 ( .A1(n7768), .A2(n7767), .ZN(n7765) );
  NAND2_X1 U8155 ( .A1(n12774), .A2(n12776), .ZN(n7873) );
  NAND2_X1 U8156 ( .A1(n7887), .A2(n12786), .ZN(n7886) );
  NAND2_X1 U8157 ( .A1(n12796), .A2(n7869), .ZN(n7868) );
  NOR2_X1 U8158 ( .A1(n7423), .A2(n7238), .ZN(n7422) );
  AND2_X1 U8159 ( .A1(n7425), .A2(n12800), .ZN(n7423) );
  AOI21_X1 U8160 ( .B1(n7537), .B2(n7536), .A(n7226), .ZN(n12585) );
  NOR2_X1 U8161 ( .A1(n12577), .A2(n12576), .ZN(n7536) );
  NAND2_X1 U8162 ( .A1(n7538), .A2(n12578), .ZN(n7537) );
  NAND2_X1 U8163 ( .A1(n7772), .A2(n7771), .ZN(n7770) );
  NOR2_X1 U8164 ( .A1(n7439), .A2(n7438), .ZN(n7437) );
  NOR2_X1 U8165 ( .A1(n7222), .A2(n12815), .ZN(n7438) );
  AOI21_X1 U8166 ( .B1(n7865), .B2(n12818), .A(n7864), .ZN(n7863) );
  AND2_X1 U8167 ( .A1(n12816), .A2(n7867), .ZN(n7866) );
  INV_X1 U8168 ( .A(n12818), .ZN(n7867) );
  INV_X1 U8169 ( .A(n9225), .ZN(n7740) );
  AOI21_X1 U8170 ( .B1(n7762), .B2(n7761), .A(n7760), .ZN(n7759) );
  AND3_X1 U8171 ( .A1(n7530), .A2(n7527), .A3(n7526), .ZN(n12617) );
  NAND2_X1 U8172 ( .A1(n12831), .A2(n7443), .ZN(n7442) );
  AND2_X1 U8173 ( .A1(n12631), .A2(n12632), .ZN(n7541) );
  NAND2_X1 U8174 ( .A1(n12633), .A2(n12530), .ZN(n7404) );
  NOR2_X1 U8175 ( .A1(n7837), .A2(n7836), .ZN(n7835) );
  INV_X1 U8176 ( .A(n8691), .ZN(n7837) );
  INV_X1 U8177 ( .A(n7681), .ZN(n7567) );
  NOR2_X1 U8178 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n8142) );
  AOI21_X1 U8179 ( .B1(n7747), .B2(n7750), .A(n7745), .ZN(n7744) );
  AND2_X1 U8180 ( .A1(n7201), .A2(n7754), .ZN(n7745) );
  NAND2_X1 U8181 ( .A1(n14397), .A2(n14250), .ZN(n10169) );
  INV_X1 U8182 ( .A(n10169), .ZN(n8009) );
  OAI21_X1 U8183 ( .B1(n8022), .B2(n7551), .A(n11779), .ZN(n7550) );
  AND2_X1 U8184 ( .A1(n12138), .A2(n15997), .ZN(n12137) );
  NAND2_X1 U8185 ( .A1(n7849), .A2(n12840), .ZN(n7848) );
  NOR2_X1 U8186 ( .A1(n9789), .A2(n9788), .ZN(n9787) );
  AND2_X1 U8187 ( .A1(n12879), .A2(n10011), .ZN(n7940) );
  INV_X1 U8188 ( .A(n10012), .ZN(n7941) );
  NAND2_X1 U8189 ( .A1(n8045), .A2(n8822), .ZN(n8824) );
  INV_X1 U8190 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n8158) );
  OAI21_X1 U8191 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(n15585), .A(n15584), .ZN(
        n15588) );
  NOR2_X1 U8192 ( .A1(n13197), .A2(n7306), .ZN(n7305) );
  INV_X1 U8193 ( .A(n12970), .ZN(n7306) );
  INV_X1 U8194 ( .A(n7453), .ZN(n7452) );
  OAI21_X1 U8195 ( .B1(n7543), .B2(n7454), .A(n12637), .ZN(n7453) );
  INV_X1 U8196 ( .A(n12656), .ZN(n12636) );
  NAND2_X1 U8197 ( .A1(n7684), .A2(n7683), .ZN(n12638) );
  NOR2_X1 U8198 ( .A1(n12656), .A2(n7206), .ZN(n7683) );
  NAND2_X1 U8199 ( .A1(n7685), .A2(n7170), .ZN(n7684) );
  CLKBUF_X1 U8200 ( .A(n8210), .Z(n7331) );
  NAND2_X1 U8201 ( .A1(n7331), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10855) );
  OR2_X1 U8202 ( .A1(n11263), .A2(n15743), .ZN(n11030) );
  OAI21_X1 U8203 ( .B1(n10985), .B2(n11670), .A(n10971), .ZN(n10972) );
  NAND2_X1 U8204 ( .A1(n15792), .A2(n11813), .ZN(n11815) );
  NAND2_X1 U8205 ( .A1(n8178), .A2(n8177), .ZN(n8536) );
  INV_X1 U8206 ( .A(n8524), .ZN(n8178) );
  INV_X1 U8207 ( .A(n8647), .ZN(n7708) );
  OR2_X1 U8208 ( .A1(n12674), .A2(n7708), .ZN(n7707) );
  AOI21_X1 U8209 ( .B1(n7463), .B2(n7465), .A(n7462), .ZN(n7461) );
  OR2_X1 U8210 ( .A1(n13700), .A2(n13552), .ZN(n12609) );
  INV_X1 U8211 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n15264) );
  OR2_X1 U8212 ( .A1(n13243), .A2(n15971), .ZN(n13054) );
  NAND2_X1 U8213 ( .A1(n12547), .A2(n12546), .ZN(n8621) );
  NAND2_X1 U8214 ( .A1(n13252), .A2(n15845), .ZN(n12542) );
  NAND2_X1 U8215 ( .A1(n8239), .A2(n8238), .ZN(n15842) );
  NAND2_X1 U8216 ( .A1(n7450), .A2(n11314), .ZN(n11015) );
  NAND2_X1 U8217 ( .A1(n12521), .A2(n7623), .ZN(n7622) );
  NAND2_X1 U8218 ( .A1(n13428), .A2(n7573), .ZN(n7621) );
  INV_X1 U8219 ( .A(n7624), .ZN(n7623) );
  AND2_X1 U8220 ( .A1(n12525), .A2(n12524), .ZN(n13398) );
  OR2_X1 U8221 ( .A1(n7293), .A2(n7393), .ZN(n7386) );
  AND2_X1 U8222 ( .A1(n7182), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7393) );
  AND2_X1 U8223 ( .A1(n7396), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7392) );
  NAND2_X1 U8224 ( .A1(n7566), .A2(n7395), .ZN(n7388) );
  NAND2_X1 U8225 ( .A1(n7891), .A2(n8610), .ZN(n7890) );
  NAND2_X1 U8226 ( .A1(n7695), .A2(n7378), .ZN(n7376) );
  NOR2_X1 U8227 ( .A1(n7379), .A2(n7287), .ZN(n7378) );
  INV_X1 U8228 ( .A(n7381), .ZN(n7379) );
  NAND2_X1 U8229 ( .A1(n7381), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7380) );
  NAND2_X1 U8230 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n7694), .ZN(n7693) );
  INV_X1 U8231 ( .A(n8453), .ZN(n7407) );
  CLKBUF_X1 U8232 ( .A(n8471), .Z(n8472) );
  NOR2_X1 U8233 ( .A1(n8115), .A2(n7699), .ZN(n7698) );
  AND2_X1 U8234 ( .A1(n10318), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8115) );
  INV_X1 U8235 ( .A(n8114), .ZN(n7699) );
  INV_X1 U8236 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8139) );
  NOR2_X1 U8237 ( .A1(n9471), .A2(n13901), .ZN(n9449) );
  AND2_X1 U8238 ( .A1(n9449), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n9428) );
  OR2_X1 U8239 ( .A1(n7482), .A2(n7484), .ZN(n7481) );
  NAND2_X1 U8240 ( .A1(n14309), .A2(n10178), .ZN(n7487) );
  AND2_X1 U8241 ( .A1(n8042), .A2(n10172), .ZN(n8039) );
  NOR2_X1 U8242 ( .A1(n14182), .A2(n14346), .ZN(n7588) );
  INV_X1 U8243 ( .A(n7329), .ZN(n9258) );
  AND2_X1 U8244 ( .A1(n12379), .A2(n16020), .ZN(n12378) );
  INV_X1 U8245 ( .A(n10164), .ZN(n8015) );
  NAND2_X1 U8246 ( .A1(n10162), .A2(n8017), .ZN(n8016) );
  NOR2_X1 U8247 ( .A1(n10163), .A2(n8018), .ZN(n8017) );
  INV_X1 U8248 ( .A(n10161), .ZN(n8018) );
  INV_X1 U8249 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9118) );
  NOR2_X1 U8250 ( .A1(n9044), .A2(n9043), .ZN(n7330) );
  INV_X1 U8251 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9043) );
  INV_X1 U8252 ( .A(n7550), .ZN(n7548) );
  NOR2_X1 U8253 ( .A1(n11398), .A2(n11742), .ZN(n7598) );
  XNOR2_X1 U8254 ( .A(n11242), .B(n9530), .ZN(n10137) );
  AND2_X1 U8255 ( .A1(n12348), .A2(n12137), .ZN(n12379) );
  INV_X1 U8256 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8745) );
  NOR2_X1 U8257 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n7505), .ZN(n7502) );
  INV_X1 U8258 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8874) );
  INV_X1 U8259 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9788) );
  INV_X1 U8260 ( .A(n14645), .ZN(n7795) );
  AND2_X1 U8261 ( .A1(n14564), .A2(n14565), .ZN(n7796) );
  INV_X1 U8262 ( .A(n7820), .ZN(n7819) );
  NOR2_X1 U8263 ( .A1(n9748), .A2(n9747), .ZN(n9746) );
  INV_X1 U8264 ( .A(n14436), .ZN(n7811) );
  AND2_X1 U8265 ( .A1(n14861), .A2(n10044), .ZN(n7960) );
  INV_X1 U8266 ( .A(n10222), .ZN(n7958) );
  AND2_X1 U8267 ( .A1(n15030), .A2(n10027), .ZN(n7949) );
  INV_X1 U8268 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9818) );
  NOR2_X1 U8269 ( .A1(n15983), .A2(n14561), .ZN(n7676) );
  NAND2_X1 U8270 ( .A1(n11152), .A2(n11151), .ZN(n7827) );
  OR2_X1 U8271 ( .A1(n10632), .A2(n10634), .ZN(n12707) );
  NOR2_X1 U8272 ( .A1(n14980), .A2(n14997), .ZN(n14983) );
  INV_X1 U8273 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9596) );
  INV_X1 U8274 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9597) );
  NAND2_X1 U8275 ( .A1(n9334), .A2(n9333), .ZN(n9346) );
  NAND2_X1 U8276 ( .A1(n9328), .A2(n9327), .ZN(n9334) );
  NAND2_X1 U8277 ( .A1(n8054), .A2(n9252), .ZN(n8052) );
  INV_X1 U8278 ( .A(n7521), .ZN(n7520) );
  AND2_X1 U8279 ( .A1(n7518), .A2(n8082), .ZN(n7517) );
  INV_X1 U8280 ( .A(n8083), .ZN(n8082) );
  NAND2_X1 U8281 ( .A1(n9160), .A2(SI_16_), .ZN(n9176) );
  NOR2_X1 U8282 ( .A1(n9177), .A2(n8087), .ZN(n8086) );
  INV_X1 U8283 ( .A(n9158), .ZN(n8087) );
  NAND2_X1 U8284 ( .A1(n9155), .A2(n9154), .ZN(n9159) );
  NAND2_X1 U8285 ( .A1(n9134), .A2(n9133), .ZN(n9155) );
  NOR2_X1 U8286 ( .A1(n8987), .A2(n8962), .ZN(n8062) );
  INV_X1 U8287 ( .A(n8984), .ZN(n8065) );
  OR2_X1 U8288 ( .A1(n9699), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n9712) );
  NOR2_X2 U8289 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n9626) );
  OAI22_X1 U8290 ( .A1(n15617), .A2(n15616), .B1(P3_ADDR_REG_6__SCAN_IN), .B2(
        n15615), .ZN(n15620) );
  INV_X1 U8291 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n15615) );
  AOI21_X1 U8292 ( .B1(n13213), .B2(n7833), .A(n13022), .ZN(n7832) );
  INV_X1 U8293 ( .A(n13020), .ZN(n7833) );
  INV_X1 U8294 ( .A(n13213), .ZN(n7834) );
  NAND2_X1 U8295 ( .A1(n8180), .A2(n15162), .ZN(n8580) );
  INV_X1 U8296 ( .A(n13010), .ZN(n7346) );
  AND2_X1 U8297 ( .A1(n13020), .A2(n13018), .ZN(n13109) );
  AND2_X1 U8298 ( .A1(n13108), .A2(n13015), .ZN(n13145) );
  OR2_X1 U8299 ( .A1(n8536), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8551) );
  INV_X1 U8300 ( .A(n8504), .ZN(n8176) );
  INV_X1 U8301 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n15261) );
  INV_X1 U8302 ( .A(n13008), .ZN(n7355) );
  INV_X1 U8303 ( .A(n8477), .ZN(n8175) );
  AND2_X1 U8304 ( .A1(n12536), .A2(n8729), .ZN(n12685) );
  OR2_X1 U8305 ( .A1(n8242), .A2(n8222), .ZN(n8226) );
  NAND2_X1 U8306 ( .A1(n11260), .A2(n7219), .ZN(n11026) );
  NAND2_X1 U8307 ( .A1(n11027), .A2(n11026), .ZN(n11025) );
  AND2_X1 U8308 ( .A1(n10856), .A2(n10891), .ZN(n7574) );
  OR2_X1 U8309 ( .A1(n10867), .A2(n10866), .ZN(n10971) );
  NAND2_X1 U8310 ( .A1(n7575), .A2(n10949), .ZN(n10859) );
  OR2_X1 U8311 ( .A1(n11201), .A2(n8267), .ZN(n11203) );
  OAI21_X1 U8312 ( .B1(n11181), .B2(n8288), .A(n11171), .ZN(n11806) );
  NAND2_X1 U8313 ( .A1(n10984), .A2(n10983), .ZN(n11787) );
  NAND2_X1 U8314 ( .A1(n15793), .A2(n15794), .ZN(n15792) );
  NAND2_X1 U8315 ( .A1(n11827), .A2(n11828), .ZN(n7586) );
  AND2_X1 U8316 ( .A1(n11831), .A2(n15807), .ZN(n7587) );
  NAND2_X1 U8317 ( .A1(n12174), .A2(n12175), .ZN(n12176) );
  NOR2_X1 U8318 ( .A1(n13254), .A2(n13253), .ZN(n7338) );
  AOI21_X1 U8319 ( .B1(n13264), .B2(n13263), .A(n13262), .ZN(n13279) );
  NAND2_X1 U8320 ( .A1(n13287), .A2(n13288), .ZN(n13291) );
  INV_X1 U8321 ( .A(n7578), .ZN(n13333) );
  NAND2_X1 U8322 ( .A1(n13323), .A2(n7216), .ZN(n13357) );
  AOI21_X1 U8323 ( .B1(n13319), .B2(n13318), .A(n13317), .ZN(n13351) );
  OAI21_X1 U8324 ( .B1(n13357), .B2(n13356), .A(n13355), .ZN(n13360) );
  OR2_X1 U8325 ( .A1(n13374), .A2(n13373), .ZN(n16038) );
  AOI21_X1 U8326 ( .B1(n13405), .B2(n8597), .A(n8200), .ZN(n13412) );
  NAND2_X1 U8327 ( .A1(n8652), .A2(n8651), .ZN(n13436) );
  AND2_X1 U8328 ( .A1(n12528), .A2(n12530), .ZN(n13435) );
  NAND2_X1 U8329 ( .A1(n7706), .A2(n8647), .ZN(n13472) );
  NAND2_X1 U8330 ( .A1(n13490), .A2(n12674), .ZN(n7706) );
  NOR2_X1 U8331 ( .A1(n7269), .A2(n8097), .ZN(n8642) );
  NAND2_X1 U8332 ( .A1(n8174), .A2(n15264), .ZN(n8461) );
  INV_X1 U8333 ( .A(n8445), .ZN(n8174) );
  OR2_X1 U8334 ( .A1(n8431), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8445) );
  NAND2_X1 U8335 ( .A1(n8172), .A2(n8171), .ZN(n8419) );
  INV_X1 U8336 ( .A(n8405), .ZN(n8172) );
  OR2_X1 U8337 ( .A1(n8369), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8381) );
  NAND2_X1 U8338 ( .A1(n8170), .A2(n8169), .ZN(n8369) );
  INV_X1 U8339 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n8169) );
  INV_X1 U8340 ( .A(n8354), .ZN(n8170) );
  OAI21_X1 U8341 ( .B1(n12253), .B2(n8631), .A(n7343), .ZN(n12284) );
  OR2_X1 U8342 ( .A1(n15929), .A2(n12285), .ZN(n7343) );
  INV_X1 U8343 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n15269) );
  NAND2_X1 U8344 ( .A1(n8167), .A2(n8166), .ZN(n8333) );
  INV_X1 U8345 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n8166) );
  INV_X1 U8346 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8164) );
  NAND2_X1 U8347 ( .A1(n15842), .A2(n12543), .ZN(n7444) );
  INV_X1 U8348 ( .A(n8621), .ZN(n12658) );
  AND2_X1 U8349 ( .A1(n8671), .A2(n12641), .ZN(n15846) );
  AND4_X1 U8350 ( .A1(n8220), .A2(n8219), .A3(n8217), .A4(n8218), .ZN(n11016)
         );
  OR2_X1 U8351 ( .A1(n8495), .A2(n11411), .ZN(n8218) );
  INV_X1 U8352 ( .A(n7702), .ZN(n12657) );
  INV_X1 U8353 ( .A(n13578), .ZN(n15851) );
  NAND2_X1 U8354 ( .A1(n7636), .A2(n12608), .ZN(n13510) );
  NAND2_X1 U8355 ( .A1(n12283), .A2(n7631), .ZN(n7625) );
  NAND2_X1 U8356 ( .A1(n7633), .A2(n12532), .ZN(n12363) );
  OAI21_X1 U8357 ( .B1(P2_DATAO_REG_27__SCAN_IN), .B2(n14413), .A(n8136), .ZN(
        n8589) );
  NAND2_X1 U8358 ( .A1(n7385), .A2(n7384), .ZN(n8562) );
  NOR2_X1 U8359 ( .A1(n7387), .A2(n7392), .ZN(n7384) );
  NAND2_X1 U8360 ( .A1(n8521), .A2(n7386), .ZN(n7385) );
  AND2_X1 U8361 ( .A1(n7388), .A2(n7394), .ZN(n7387) );
  XNOR2_X1 U8362 ( .A(n8679), .B(n8678), .ZN(n8689) );
  OR2_X1 U8363 ( .A1(n8680), .A2(n8344), .ZN(n8679) );
  NAND2_X1 U8364 ( .A1(n7391), .A2(n7389), .ZN(n8545) );
  INV_X1 U8365 ( .A(n7390), .ZN(n7389) );
  OR2_X1 U8366 ( .A1(n8521), .A2(n7396), .ZN(n7391) );
  AOI21_X1 U8367 ( .B1(n8521), .B2(n7182), .A(n7388), .ZN(n8547) );
  NAND2_X1 U8368 ( .A1(n8709), .A2(n8708), .ZN(n10849) );
  AND2_X1 U8369 ( .A1(n8397), .A2(n8396), .ZN(n8401) );
  XNOR2_X1 U8370 ( .A(n8122), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8395) );
  NOR2_X1 U8371 ( .A1(n8390), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n8397) );
  INV_X1 U8372 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8396) );
  AOI21_X1 U8373 ( .B1(n8362), .B2(n7374), .A(n7371), .ZN(n7370) );
  NAND2_X1 U8374 ( .A1(n7372), .A2(n8121), .ZN(n7371) );
  OR2_X1 U8375 ( .A1(n8364), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n8390) );
  OAI21_X1 U8376 ( .B1(n7399), .B2(n7398), .A(n7397), .ZN(n8341) );
  INV_X1 U8377 ( .A(n7400), .ZN(n7398) );
  AOI21_X1 U8378 ( .B1(n7400), .B2(n7164), .A(n7244), .ZN(n7397) );
  XNOR2_X1 U8379 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n8339) );
  XNOR2_X1 U8380 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8232) );
  NOR2_X1 U8381 ( .A1(n8808), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8231) );
  AOI21_X1 U8382 ( .B1(n7994), .B2(n7993), .A(n8094), .ZN(n7992) );
  INV_X1 U8383 ( .A(n13826), .ZN(n7993) );
  INV_X1 U8384 ( .A(n7328), .ZN(n9307) );
  NAND2_X1 U8385 ( .A1(n7328), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n9339) );
  INV_X1 U8386 ( .A(n10257), .ZN(n10255) );
  NAND2_X1 U8387 ( .A1(n7324), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8972) );
  INV_X1 U8388 ( .A(n8951), .ZN(n7324) );
  INV_X1 U8389 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8971) );
  NAND2_X1 U8390 ( .A1(n9274), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n9290) );
  INV_X1 U8391 ( .A(n7987), .ZN(n7986) );
  OAI21_X1 U8392 ( .B1(n7988), .B2(n12407), .A(n12447), .ZN(n7987) );
  OR2_X1 U8393 ( .A1(n9168), .A2(n9167), .ZN(n9186) );
  NAND2_X1 U8394 ( .A1(n12058), .A2(n12059), .ZN(n12101) );
  INV_X1 U8395 ( .A(n11944), .ZN(n7977) );
  AOI21_X1 U8396 ( .B1(n7976), .B2(n11944), .A(n7975), .ZN(n7974) );
  NOR2_X1 U8397 ( .A1(n11946), .A2(n7334), .ZN(n7975) );
  INV_X1 U8398 ( .A(n11947), .ZN(n7334) );
  OR2_X1 U8399 ( .A1(n9218), .A2(n9217), .ZN(n9233) );
  XNOR2_X1 U8400 ( .A(n14228), .B(n13773), .ZN(n13739) );
  NAND2_X1 U8401 ( .A1(n13836), .A2(n13837), .ZN(n13835) );
  AND2_X1 U8402 ( .A1(n9398), .A2(n10183), .ZN(n10439) );
  NOR2_X1 U8403 ( .A1(n9560), .A2(n7325), .ZN(n9561) );
  AND4_X1 U8405 ( .A1(n8911), .A2(n8910), .A3(n8909), .A4(n8908), .ZN(n11067)
         );
  AND4_X1 U8406 ( .A1(n8882), .A2(n8881), .A3(n8880), .A4(n8879), .ZN(n10785)
         );
  AND4_X1 U8407 ( .A1(n8835), .A2(n8834), .A3(n8833), .A4(n8832), .ZN(n10241)
         );
  NAND2_X1 U8408 ( .A1(n8786), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8833) );
  OR2_X1 U8409 ( .A1(n8856), .A2(n10545), .ZN(n8795) );
  OR2_X1 U8410 ( .A1(n8856), .A2(n8784), .ZN(n8788) );
  INV_X1 U8411 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n9162) );
  INV_X1 U8412 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n9212) );
  OAI21_X2 U8413 ( .B1(n9135), .B2(n8772), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8779) );
  INV_X1 U8414 ( .A(n7595), .ZN(n14067) );
  NAND2_X1 U8415 ( .A1(n14314), .A2(n13913), .ZN(n7645) );
  OR2_X1 U8416 ( .A1(n14130), .A2(n14119), .ZN(n14117) );
  AND2_X1 U8417 ( .A1(n9471), .A2(n9356), .ZN(n14120) );
  AND2_X1 U8418 ( .A1(n8073), .A2(n14116), .ZN(n8071) );
  NAND3_X1 U8419 ( .A1(n14216), .A2(n14149), .A3(n7165), .ZN(n14152) );
  OR2_X1 U8420 ( .A1(n14152), .A2(n14326), .ZN(n14130) );
  NAND2_X1 U8421 ( .A1(n8038), .A2(n8036), .ZN(n14157) );
  OR2_X1 U8422 ( .A1(n8040), .A2(n8037), .ZN(n8036) );
  NAND2_X1 U8423 ( .A1(n10171), .A2(n8039), .ZN(n8038) );
  INV_X1 U8424 ( .A(n10172), .ZN(n8037) );
  NAND2_X1 U8425 ( .A1(n14216), .A2(n14195), .ZN(n14191) );
  NOR2_X1 U8426 ( .A1(n14254), .A2(n14228), .ZN(n14227) );
  OR2_X1 U8427 ( .A1(n9119), .A2(n9118), .ZN(n9140) );
  NAND2_X1 U8428 ( .A1(n8016), .A2(n10164), .ZN(n12373) );
  INV_X1 U8429 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9095) );
  OR2_X1 U8430 ( .A1(n9096), .A2(n9095), .ZN(n9119) );
  INV_X1 U8431 ( .A(n12012), .ZN(n7650) );
  AND4_X1 U8432 ( .A1(n9072), .A2(n9071), .A3(n9070), .A4(n9069), .ZN(n12144)
         );
  AND4_X1 U8433 ( .A1(n9126), .A2(n9125), .A3(n9124), .A4(n9123), .ZN(n12334)
         );
  NAND2_X1 U8434 ( .A1(n7330), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9096) );
  NAND2_X1 U8435 ( .A1(n8006), .A2(n7215), .ZN(n12015) );
  AND2_X1 U8436 ( .A1(n12007), .A2(n12203), .ZN(n12138) );
  NOR2_X1 U8437 ( .A1(n7596), .A2(n11737), .ZN(n12007) );
  INV_X1 U8438 ( .A(n8006), .ZN(n12014) );
  NAND2_X1 U8439 ( .A1(n9017), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9044) );
  INV_X1 U8440 ( .A(n9019), .ZN(n9017) );
  NAND2_X1 U8441 ( .A1(n10156), .A2(n10155), .ZN(n11778) );
  INV_X1 U8442 ( .A(n7596), .ZN(n11773) );
  INV_X1 U8443 ( .A(n7598), .ZN(n11774) );
  INV_X1 U8444 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8996) );
  OR2_X1 U8445 ( .A1(n8997), .A2(n8996), .ZN(n9019) );
  OR2_X1 U8446 ( .A1(n8972), .A2(n8971), .ZN(n8997) );
  CLKBUF_X1 U8447 ( .A(n10236), .Z(n14279) );
  NAND2_X1 U8448 ( .A1(n8024), .A2(n10153), .ZN(n11590) );
  OR2_X1 U8449 ( .A1(n11390), .A2(n8025), .ZN(n8024) );
  OAI21_X1 U8450 ( .B1(n10151), .B2(n7184), .A(n7496), .ZN(n11390) );
  AND2_X1 U8451 ( .A1(n11344), .A2(n11546), .ZN(n11397) );
  NAND2_X1 U8452 ( .A1(n10963), .A2(n11535), .ZN(n11213) );
  AND2_X1 U8453 ( .A1(n10753), .A2(n11524), .ZN(n10963) );
  NAND2_X1 U8454 ( .A1(n10144), .A2(n10143), .ZN(n10757) );
  AND2_X1 U8455 ( .A1(n11415), .A2(n10744), .ZN(n10753) );
  XNOR2_X1 U8456 ( .A(n11374), .B(n13931), .ZN(n10703) );
  NAND2_X1 U8457 ( .A1(n10108), .A2(n11250), .ZN(n10718) );
  AOI22_X1 U8458 ( .A1(n13931), .A2(n14275), .B1(n9548), .B2(n14274), .ZN(
        n10719) );
  AOI21_X1 U8459 ( .B1(n10610), .B2(n9467), .A(n9041), .ZN(n15965) );
  NAND2_X1 U8460 ( .A1(n10151), .A2(n10150), .ZN(n11347) );
  INV_X1 U8461 ( .A(n16033), .ZN(n14353) );
  INV_X1 U8462 ( .A(n16029), .ZN(n14347) );
  INV_X1 U8463 ( .A(n10209), .ZN(n15450) );
  XNOR2_X1 U8464 ( .A(n9527), .B(n9526), .ZN(n10438) );
  INV_X1 U8465 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8757) );
  INV_X1 U8466 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9540) );
  OAI21_X1 U8467 ( .B1(n9534), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9536) );
  INV_X1 U8468 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9535) );
  NAND2_X1 U8469 ( .A1(n8766), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8770) );
  INV_X1 U8470 ( .A(n8766), .ZN(n8768) );
  OR3_X1 U8471 ( .A1(n9014), .A2(P2_IR_REG_9__SCAN_IN), .A3(n9013), .ZN(n9032)
         );
  OR2_X1 U8472 ( .A1(n8899), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n9114) );
  NOR2_X1 U8473 ( .A1(n14556), .A2(n7814), .ZN(n7813) );
  INV_X1 U8474 ( .A(n14441), .ZN(n7814) );
  NAND2_X1 U8475 ( .A1(n14437), .A2(n14436), .ZN(n7815) );
  INV_X1 U8476 ( .A(n9922), .ZN(n9923) );
  NAND2_X1 U8477 ( .A1(n10583), .A2(n12706), .ZN(n14585) );
  OR2_X1 U8478 ( .A1(n9718), .A2(n9717), .ZN(n9733) );
  NAND2_X1 U8479 ( .A1(n14655), .A2(n7804), .ZN(n7800) );
  AOI21_X1 U8480 ( .B1(n7799), .B2(n14655), .A(n7806), .ZN(n7798) );
  AOI22_X1 U8481 ( .A1(n14700), .A2(n14699), .B1(n14457), .B2(n14458), .ZN(
        n14627) );
  INV_X1 U8482 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9691) );
  AND2_X1 U8483 ( .A1(n7796), .A2(n7795), .ZN(n7794) );
  NAND2_X1 U8484 ( .A1(n14663), .A2(n7796), .ZN(n14647) );
  OR2_X1 U8485 ( .A1(n9733), .A2(n9732), .ZN(n9748) );
  INV_X1 U8486 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9747) );
  NAND2_X1 U8487 ( .A1(n7783), .A2(n7160), .ZN(n12324) );
  NAND2_X1 U8488 ( .A1(n12300), .A2(n12299), .ZN(n7783) );
  OR2_X1 U8489 ( .A1(n12868), .A2(n10353), .ZN(n14607) );
  OR2_X1 U8490 ( .A1(n9872), .A2(n14681), .ZN(n9886) );
  NAND2_X1 U8491 ( .A1(n14677), .A2(n14678), .ZN(n14676) );
  OR2_X1 U8492 ( .A1(n11295), .A2(n11294), .ZN(n7824) );
  AOI21_X1 U8493 ( .B1(n7790), .B2(n7162), .A(n7788), .ZN(n7787) );
  INV_X1 U8494 ( .A(n14531), .ZN(n7788) );
  OR2_X1 U8495 ( .A1(n9819), .A2(n9818), .ZN(n9832) );
  MUX2_X1 U8496 ( .A(n12909), .B(n12908), .S(n12871), .Z(n12938) );
  INV_X1 U8497 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n15642) );
  AND2_X1 U8498 ( .A1(n10601), .A2(n10600), .ZN(n10602) );
  INV_X1 U8499 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10596) );
  INV_X1 U8500 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n14705) );
  NOR2_X1 U8501 ( .A1(n14826), .A2(n15382), .ZN(n14829) );
  NOR2_X1 U8502 ( .A1(n14865), .A2(n14599), .ZN(n10220) );
  OR2_X1 U8503 ( .A1(n14878), .A2(n14870), .ZN(n14865) );
  OAI21_X1 U8504 ( .B1(n14925), .B2(n7922), .A(n7920), .ZN(n14886) );
  INV_X1 U8505 ( .A(n7921), .ZN(n7920) );
  OAI21_X1 U8506 ( .B1(n7924), .B2(n7922), .A(n9948), .ZN(n7921) );
  AND2_X1 U8507 ( .A1(n7176), .A2(n15392), .ZN(n7667) );
  INV_X1 U8508 ( .A(n7954), .ZN(n7953) );
  OAI21_X1 U8509 ( .B1(n14915), .B2(n7192), .A(n10041), .ZN(n7954) );
  NAND2_X1 U8510 ( .A1(n14953), .A2(n7669), .ZN(n14917) );
  NAND2_X1 U8511 ( .A1(n14953), .A2(n15108), .ZN(n14939) );
  AND2_X1 U8512 ( .A1(n7932), .A2(n7864), .ZN(n7930) );
  NAND2_X1 U8513 ( .A1(n14974), .A2(n7220), .ZN(n14958) );
  AND2_X1 U8514 ( .A1(n7674), .A2(n7673), .ZN(n7672) );
  NAND2_X1 U8515 ( .A1(n15044), .A2(n7949), .ZN(n15029) );
  AOI21_X1 U8516 ( .B1(n7914), .B2(n11961), .A(n7199), .ZN(n7912) );
  NAND2_X1 U8517 ( .A1(n15046), .A2(n15045), .ZN(n15044) );
  NAND2_X1 U8518 ( .A1(n11867), .A2(n7674), .ZN(n15049) );
  NAND2_X1 U8519 ( .A1(n11867), .A2(n11970), .ZN(n12072) );
  OR2_X1 U8520 ( .A1(n7946), .A2(n7945), .ZN(n7944) );
  INV_X1 U8521 ( .A(n10023), .ZN(n7945) );
  AOI21_X1 U8522 ( .B1(n7927), .B2(n12886), .A(n7211), .ZN(n7926) );
  NAND2_X1 U8523 ( .A1(n11866), .A2(n12890), .ZN(n11865) );
  NAND2_X1 U8524 ( .A1(n11455), .A2(n7168), .ZN(n11578) );
  NAND2_X1 U8525 ( .A1(n7660), .A2(n7659), .ZN(n11701) );
  INV_X1 U8526 ( .A(n11456), .ZN(n7660) );
  NAND2_X1 U8527 ( .A1(n11455), .A2(n15943), .ZN(n11699) );
  AND2_X1 U8528 ( .A1(n15880), .A2(n15879), .ZN(n15881) );
  NAND2_X1 U8529 ( .A1(n7827), .A2(n10009), .ZN(n15872) );
  CLKBUF_X1 U8530 ( .A(n11151), .Z(n12874) );
  NAND2_X1 U8531 ( .A1(n7350), .A2(n15878), .ZN(n7666) );
  XNOR2_X1 U8532 ( .A(n14829), .B(n15064), .ZN(n7350) );
  INV_X1 U8533 ( .A(n9893), .ZN(n12863) );
  OR2_X1 U8534 ( .A1(n14858), .A2(n15884), .ZN(n7919) );
  OR2_X1 U8535 ( .A1(n12703), .A2(n7429), .ZN(n15884) );
  NAND2_X1 U8536 ( .A1(n15878), .A2(n10000), .ZN(n10581) );
  XNOR2_X1 U8537 ( .A(n9446), .B(n9445), .ZN(n14410) );
  NAND2_X1 U8538 ( .A1(n9443), .A2(n9442), .ZN(n9446) );
  XNOR2_X1 U8539 ( .A(n10069), .B(P1_IR_REG_26__SCAN_IN), .ZN(n10091) );
  XNOR2_X1 U8540 ( .A(n9466), .B(n9465), .ZN(n14414) );
  XNOR2_X1 U8541 ( .A(n10063), .B(P1_IR_REG_25__SCAN_IN), .ZN(n10092) );
  NAND2_X1 U8542 ( .A1(n10066), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10063) );
  AND2_X1 U8543 ( .A1(n10067), .A2(n10066), .ZN(n10083) );
  XNOR2_X1 U8544 ( .A(n10085), .B(P1_IR_REG_23__SCAN_IN), .ZN(n10324) );
  OAI21_X1 U8545 ( .B1(n10084), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10085) );
  NAND2_X1 U8546 ( .A1(n10001), .A2(n9999), .ZN(n10084) );
  NAND2_X1 U8547 ( .A1(n8060), .A2(n8053), .ZN(n8059) );
  INV_X1 U8548 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9997) );
  INV_X1 U8549 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n10007) );
  NAND2_X1 U8550 ( .A1(n8060), .A2(n9251), .ZN(n9271) );
  NAND2_X1 U8551 ( .A1(n9112), .A2(n9111), .ZN(n9130) );
  NAND2_X1 U8552 ( .A1(n7507), .A2(n7511), .ZN(n9082) );
  OR2_X1 U8553 ( .A1(n9010), .A2(n7512), .ZN(n7507) );
  XNOR2_X1 U8554 ( .A(n9062), .B(n9061), .ZN(n10610) );
  NAND2_X1 U8555 ( .A1(n9031), .A2(n9030), .ZN(n9062) );
  AOI21_X1 U8556 ( .B1(n8937), .B2(n8070), .A(n8069), .ZN(n8068) );
  INV_X1 U8557 ( .A(n8919), .ZN(n8070) );
  NAND2_X1 U8558 ( .A1(n7323), .A2(n8893), .ZN(n8896) );
  AND2_X1 U8559 ( .A1(n8866), .A2(n8848), .ZN(n10302) );
  XNOR2_X1 U8560 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n15573) );
  AND2_X1 U8561 ( .A1(n7607), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n15574) );
  AOI22_X1 U8562 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n15612), .B1(n15611), .B2(
        n15610), .ZN(n15616) );
  OR2_X1 U8563 ( .A1(n15612), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n15610) );
  INV_X1 U8564 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n15612) );
  OAI21_X1 U8565 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n15637), .A(n15636), .ZN(
        n15639) );
  AOI21_X1 U8566 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n15651), .A(n15650), .ZN(
        n15663) );
  NOR2_X1 U8567 ( .A1(n15649), .A2(n15648), .ZN(n15650) );
  CLKBUF_X1 U8568 ( .A(n13068), .Z(n13069) );
  INV_X1 U8569 ( .A(n13244), .ZN(n13048) );
  OAI22_X1 U8570 ( .A1(n11433), .A2(n11434), .B1(n11432), .B2(n13252), .ZN(
        n11435) );
  NAND2_X1 U8571 ( .A1(n7303), .A2(n13002), .ZN(n13087) );
  NAND2_X1 U8572 ( .A1(n8514), .A2(n8513), .ZN(n13480) );
  AND2_X1 U8573 ( .A1(n8557), .A2(n8556), .ZN(n13450) );
  CLKBUF_X1 U8574 ( .A(n13106), .Z(n13107) );
  NAND2_X1 U8575 ( .A1(n12228), .A2(n7183), .ZN(n12231) );
  CLKBUF_X1 U8576 ( .A(n13163), .Z(n7303) );
  AND4_X1 U8577 ( .A1(n8387), .A2(n8386), .A3(n8385), .A4(n8384), .ZN(n13193)
         );
  INV_X1 U8578 ( .A(n7877), .ZN(n7876) );
  OAI21_X1 U8579 ( .B1(n7167), .B2(n7878), .A(n13204), .ZN(n7877) );
  NAND2_X1 U8580 ( .A1(n7875), .A2(n7879), .ZN(n13205) );
  NAND2_X1 U8581 ( .A1(n7883), .A2(n7167), .ZN(n7875) );
  OAI21_X1 U8582 ( .B1(n12653), .B2(n8728), .A(n7412), .ZN(n7411) );
  NAND2_X1 U8583 ( .A1(n12653), .A2(n15861), .ZN(n7412) );
  INV_X1 U8584 ( .A(n13437), .ZN(n13238) );
  INV_X1 U8585 ( .A(n13450), .ZN(n13423) );
  OR2_X1 U8586 ( .A1(n11092), .A2(n10234), .ZN(n13240) );
  INV_X1 U8587 ( .A(n13193), .ZN(n13243) );
  INV_X1 U8588 ( .A(n12423), .ZN(n13245) );
  INV_X1 U8589 ( .A(n11918), .ZN(n13249) );
  INV_X1 U8590 ( .A(n11724), .ZN(n13250) );
  INV_X1 U8591 ( .A(n11662), .ZN(n15847) );
  INV_X1 U8592 ( .A(n11334), .ZN(n13252) );
  INV_X1 U8593 ( .A(n11016), .ZN(n7450) );
  INV_X1 U8594 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n15749) );
  INV_X1 U8595 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n15576) );
  NAND3_X1 U8596 ( .A1(n10859), .A2(n7576), .A3(P3_REG1_REG_3__SCAN_IN), .ZN(
        n10934) );
  NAND2_X1 U8597 ( .A1(n10976), .A2(n10975), .ZN(n11199) );
  OR2_X1 U8598 ( .A1(n11169), .A2(n11168), .ZN(n11171) );
  NOR2_X1 U8599 ( .A1(n8348), .A2(n8347), .ZN(n15780) );
  NOR2_X1 U8600 ( .A1(n7583), .A2(n12169), .ZN(n12168) );
  AND2_X1 U8601 ( .A1(n7583), .A2(n7581), .ZN(n12172) );
  NOR2_X1 U8602 ( .A1(n13274), .A2(n13275), .ZN(n13278) );
  AOI21_X1 U8603 ( .B1(n13339), .B2(n13338), .A(n13337), .ZN(n13346) );
  INV_X1 U8604 ( .A(n15742), .ZN(n15815) );
  AND2_X1 U8605 ( .A1(n12498), .A2(n12497), .ZN(n13376) );
  NAND2_X1 U8606 ( .A1(n9574), .A2(n12634), .ZN(n12487) );
  AND2_X1 U8607 ( .A1(n7221), .A2(n13415), .ZN(n13602) );
  NAND2_X1 U8608 ( .A1(n13426), .A2(n12519), .ZN(n13414) );
  NAND2_X1 U8609 ( .A1(n13488), .A2(n12619), .ZN(n13476) );
  NAND2_X1 U8610 ( .A1(n13519), .A2(n8644), .ZN(n13503) );
  NAND2_X1 U8611 ( .A1(n8492), .A2(n8491), .ZN(n13514) );
  NAND2_X1 U8612 ( .A1(n8476), .A2(n8475), .ZN(n13636) );
  NAND2_X1 U8613 ( .A1(n8639), .A2(n8638), .ZN(n13576) );
  NAND2_X1 U8614 ( .A1(n8411), .A2(n12588), .ZN(n13585) );
  NAND2_X1 U8615 ( .A1(n7470), .A2(n7626), .ZN(n12474) );
  NAND2_X1 U8616 ( .A1(n8352), .A2(n7474), .ZN(n7470) );
  INV_X1 U8617 ( .A(n12225), .ZN(n15929) );
  NAND2_X1 U8618 ( .A1(n12243), .A2(n8330), .ZN(n12252) );
  NAND2_X1 U8619 ( .A1(n11988), .A2(n8628), .ZN(n12240) );
  OAI21_X1 U8620 ( .B1(n11850), .B2(n8626), .A(n7457), .ZN(n11987) );
  NAND2_X1 U8621 ( .A1(n11903), .A2(n12661), .ZN(n11902) );
  NAND2_X1 U8622 ( .A1(n11850), .A2(n12556), .ZN(n11903) );
  NAND2_X1 U8623 ( .A1(n11663), .A2(n8624), .ZN(n11854) );
  AND2_X1 U8624 ( .A1(n15867), .A2(n11842), .ZN(n13592) );
  INV_X1 U8625 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n15169) );
  INV_X2 U8626 ( .A(n15867), .ZN(n15869) );
  NAND2_X1 U8627 ( .A1(n11109), .A2(n11107), .ZN(n15860) );
  AND2_X1 U8628 ( .A1(n15867), .A2(n15866), .ZN(n13500) );
  INV_X1 U8629 ( .A(n15860), .ZN(n13541) );
  AND3_X1 U8630 ( .A1(n8318), .A2(n8317), .A3(n8316), .ZN(n11994) );
  AND3_X1 U8631 ( .A1(n8287), .A2(n8286), .A3(n8285), .ZN(n13129) );
  INV_X1 U8632 ( .A(n15970), .ZN(n15907) );
  INV_X1 U8633 ( .A(n13376), .ZN(n16050) );
  NAND2_X1 U8634 ( .A1(n12512), .A2(n12511), .ZN(n16041) );
  INV_X1 U8635 ( .A(n13105), .ZN(n13671) );
  NAND2_X1 U8636 ( .A1(n13036), .A2(n7157), .ZN(n13675) );
  AND2_X1 U8637 ( .A1(n8523), .A2(n8522), .ZN(n13683) );
  INV_X1 U8638 ( .A(n12999), .ZN(n13691) );
  NAND2_X1 U8639 ( .A1(n8418), .A2(n8417), .ZN(n13706) );
  INV_X1 U8640 ( .A(n13191), .ZN(n12471) );
  AND3_X1 U8641 ( .A1(n8265), .A2(n8264), .A3(n8263), .ZN(n15906) );
  AND2_X1 U8642 ( .A1(n8695), .A2(n8694), .ZN(n13709) );
  AND2_X1 U8643 ( .A1(n10849), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13710) );
  AND2_X1 U8644 ( .A1(n8149), .A2(n8184), .ZN(n7475) );
  NAND2_X1 U8645 ( .A1(n7715), .A2(n7892), .ZN(n7360) );
  XNOR2_X1 U8646 ( .A(n8194), .B(n8193), .ZN(n13727) );
  XNOR2_X1 U8647 ( .A(n8576), .B(n8575), .ZN(n12261) );
  CLKBUF_X1 U8648 ( .A(n8689), .Z(n8690) );
  NAND2_X1 U8649 ( .A1(n7568), .A2(n7681), .ZN(n8532) );
  NAND2_X1 U8650 ( .A1(n8521), .A2(n8519), .ZN(n7568) );
  NOR2_X1 U8651 ( .A1(n8606), .A2(n8605), .ZN(n12697) );
  NAND2_X1 U8652 ( .A1(n7892), .A2(n7891), .ZN(n7895) );
  XNOR2_X1 U8653 ( .A(n8608), .B(n8607), .ZN(n11308) );
  OAI211_X1 U8654 ( .C1(n7695), .C2(P1_DATAO_REG_20__SCAN_IN), .A(n7377), .B(
        n7381), .ZN(n8501) );
  NAND2_X1 U8655 ( .A1(n7695), .A2(n7287), .ZN(n7377) );
  INV_X1 U8656 ( .A(SI_20_), .ZN(n15191) );
  INV_X1 U8657 ( .A(SI_18_), .ZN(n15300) );
  INV_X1 U8658 ( .A(SI_17_), .ZN(n15301) );
  OAI21_X1 U8659 ( .B1(n7687), .B2(n7288), .A(n7408), .ZN(n8454) );
  NAND2_X1 U8660 ( .A1(n7687), .A2(n7686), .ZN(n8438) );
  INV_X1 U8661 ( .A(SI_15_), .ZN(n15313) );
  NAND2_X1 U8662 ( .A1(n7688), .A2(n8126), .ZN(n8426) );
  NAND2_X1 U8663 ( .A1(n8413), .A2(n8412), .ZN(n7688) );
  INV_X1 U8664 ( .A(SI_11_), .ZN(n15275) );
  INV_X1 U8665 ( .A(n7373), .ZN(n8376) );
  AOI21_X1 U8666 ( .B1(n8362), .B2(n8361), .A(n7185), .ZN(n7373) );
  INV_X1 U8667 ( .A(n7561), .ZN(n8327) );
  AOI21_X1 U8668 ( .B1(n8313), .B2(n8311), .A(n7186), .ZN(n7561) );
  NAND2_X1 U8669 ( .A1(n7700), .A2(n8114), .ZN(n8300) );
  INV_X1 U8670 ( .A(n10978), .ZN(n11206) );
  AND4_X1 U8671 ( .A1(n9049), .A2(n9048), .A3(n9047), .A4(n9046), .ZN(n11948)
         );
  XNOR2_X1 U8672 ( .A(n11946), .B(n11947), .ZN(n11944) );
  NAND2_X1 U8673 ( .A1(n11879), .A2(n11878), .ZN(n11945) );
  NAND2_X1 U8674 ( .A1(n13877), .A2(n10245), .ZN(n10258) );
  AND2_X1 U8675 ( .A1(n10544), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13856) );
  AND2_X1 U8676 ( .A1(n9265), .A2(n9264), .ZN(n14210) );
  NAND2_X1 U8677 ( .A1(n7965), .A2(n7966), .ZN(n13793) );
  OR2_X1 U8678 ( .A1(n13836), .A2(n7970), .ZN(n7965) );
  INV_X1 U8679 ( .A(n8001), .ZN(n8000) );
  AND2_X1 U8680 ( .A1(n11642), .A2(n11641), .ZN(n11652) );
  NAND2_X1 U8681 ( .A1(n7337), .A2(n7336), .ZN(n10540) );
  INV_X1 U8682 ( .A(n10542), .ZN(n7336) );
  INV_X1 U8683 ( .A(n10543), .ZN(n7337) );
  NAND2_X1 U8684 ( .A1(n10825), .A2(n10824), .ZN(n11059) );
  NAND2_X1 U8685 ( .A1(n7335), .A2(n10822), .ZN(n10824) );
  INV_X1 U8686 ( .A(n13757), .ZN(n13758) );
  NAND2_X1 U8687 ( .A1(n7523), .A2(n13794), .ZN(n7358) );
  NAND2_X1 U8688 ( .A1(n12101), .A2(n12100), .ZN(n12340) );
  NAND2_X1 U8689 ( .A1(n13835), .A2(n13738), .ZN(n13886) );
  NAND2_X1 U8690 ( .A1(n7981), .A2(n7984), .ZN(n7979) );
  NAND2_X1 U8691 ( .A1(n7978), .A2(n7981), .ZN(n11066) );
  NAND2_X1 U8692 ( .A1(n7335), .A2(n7983), .ZN(n7978) );
  NAND2_X1 U8693 ( .A1(n13825), .A2(n13768), .ZN(n13896) );
  NAND2_X1 U8694 ( .A1(n10266), .A2(n14255), .ZN(n13905) );
  INV_X1 U8695 ( .A(n13856), .ZN(n13902) );
  INV_X1 U8696 ( .A(n7985), .ZN(n12448) );
  NAND2_X1 U8697 ( .A1(n12408), .A2(n12407), .ZN(n12409) );
  AOI21_X1 U8698 ( .B1(n12344), .B2(n12407), .A(n7988), .ZN(n7985) );
  INV_X1 U8699 ( .A(n13907), .ZN(n13881) );
  INV_X1 U8700 ( .A(n13905), .ZN(n13889) );
  INV_X1 U8701 ( .A(n13898), .ZN(n13914) );
  INV_X1 U8702 ( .A(n11644), .ZN(n13924) );
  AND2_X1 U8703 ( .A1(n8860), .A2(n8859), .ZN(n8861) );
  INV_X1 U8704 ( .A(n10241), .ZN(n13931) );
  NAND2_X1 U8705 ( .A1(n10192), .A2(n10191), .ZN(n14056) );
  NAND2_X1 U8706 ( .A1(n10186), .A2(n14271), .ZN(n10192) );
  INV_X1 U8707 ( .A(n7479), .ZN(n14072) );
  AOI21_X1 U8708 ( .B1(n14098), .B2(n7484), .A(n7482), .ZN(n7479) );
  NAND2_X1 U8709 ( .A1(n9427), .A2(n9426), .ZN(n14305) );
  INV_X1 U8710 ( .A(n14309), .ZN(n14093) );
  NAND2_X1 U8711 ( .A1(n7198), .A2(n7488), .ZN(n14083) );
  NAND2_X1 U8712 ( .A1(n14136), .A2(n8034), .ZN(n14135) );
  NAND2_X1 U8713 ( .A1(n14144), .A2(n10135), .ZN(n14136) );
  NAND2_X1 U8714 ( .A1(n8029), .A2(n8031), .ZN(n14126) );
  NAND2_X1 U8715 ( .A1(n7653), .A2(n7654), .ZN(n14174) );
  NAND2_X1 U8716 ( .A1(n8041), .A2(n8040), .ZN(n14170) );
  AND2_X1 U8717 ( .A1(n8041), .A2(n7205), .ZN(n14171) );
  NAND2_X1 U8718 ( .A1(n14205), .A2(n10131), .ZN(n14196) );
  AND2_X1 U8719 ( .A1(n10171), .A2(n10170), .ZN(n14187) );
  NAND2_X1 U8720 ( .A1(n8007), .A2(n7166), .ZN(n14234) );
  NAND2_X1 U8721 ( .A1(n10167), .A2(n10166), .ZN(n14248) );
  NAND2_X1 U8722 ( .A1(n14268), .A2(n10128), .ZN(n14253) );
  NAND2_X1 U8723 ( .A1(n12369), .A2(n10127), .ZN(n14266) );
  NAND2_X1 U8724 ( .A1(n10162), .A2(n10161), .ZN(n12214) );
  NAND2_X1 U8725 ( .A1(n11587), .A2(n8022), .ZN(n7549) );
  NAND2_X1 U8726 ( .A1(n11211), .A2(n10116), .ZN(n11342) );
  AND2_X1 U8727 ( .A1(n14280), .A2(n11249), .ZN(n14258) );
  INV_X1 U8728 ( .A(n12348), .ZN(n12279) );
  INV_X1 U8729 ( .A(n12203), .ZN(n12200) );
  INV_X1 U8730 ( .A(n11643), .ZN(n11657) );
  INV_X1 U8731 ( .A(n11546), .ZN(n11387) );
  INV_X1 U8732 ( .A(n11415), .ZN(n10750) );
  NAND2_X1 U8733 ( .A1(n7237), .A2(n8802), .ZN(n8812) );
  INV_X1 U8734 ( .A(n14369), .ZN(n14300) );
  INV_X1 U8735 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n7313) );
  NAND2_X1 U8736 ( .A1(n14294), .A2(n14296), .ZN(n14372) );
  AND2_X1 U8737 ( .A1(n9354), .A2(n9353), .ZN(n14384) );
  INV_X1 U8738 ( .A(n14182), .ZN(n14391) );
  INV_X1 U8739 ( .A(n14228), .ZN(n14397) );
  AND2_X1 U8740 ( .A1(n9166), .A2(n9165), .ZN(n14403) );
  NOR2_X1 U8741 ( .A1(n10260), .A2(n15452), .ZN(n15448) );
  INV_X1 U8742 ( .A(n15455), .ZN(n15452) );
  INV_X1 U8743 ( .A(n8785), .ZN(n14405) );
  XNOR2_X1 U8744 ( .A(n9539), .B(n9538), .ZN(n14417) );
  NAND2_X1 U8745 ( .A1(n9543), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9539) );
  NAND2_X1 U8746 ( .A1(n9543), .A2(n9542), .ZN(n12480) );
  OR2_X1 U8747 ( .A1(n9541), .A2(n9540), .ZN(n9542) );
  XNOR2_X1 U8748 ( .A(n9536), .B(n9535), .ZN(n12459) );
  INV_X1 U8749 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n14423) );
  INV_X1 U8750 ( .A(n9398), .ZN(n9530) );
  INV_X1 U8751 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n12359) );
  INV_X1 U8752 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10318) );
  INV_X1 U8753 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10298) );
  AOI21_X1 U8754 ( .B1(n7823), .B2(n11294), .A(n7213), .ZN(n7821) );
  NAND2_X1 U8755 ( .A1(n7815), .A2(n14441), .ZN(n14555) );
  NAND2_X1 U8756 ( .A1(n14676), .A2(n7807), .ZN(n14576) );
  NAND2_X1 U8757 ( .A1(n11762), .A2(n11761), .ZN(n11764) );
  NAND2_X1 U8758 ( .A1(n10625), .A2(n10644), .ZN(n7777) );
  AND2_X1 U8759 ( .A1(n7780), .A2(n12323), .ZN(n7779) );
  NAND2_X1 U8760 ( .A1(n7333), .A2(n7160), .ZN(n7778) );
  OAI21_X1 U8761 ( .B1(n14663), .B2(n7162), .A(n7790), .ZN(n14614) );
  NAND2_X1 U8762 ( .A1(n7792), .A2(n7793), .ZN(n14649) );
  NAND2_X1 U8763 ( .A1(n14663), .A2(n7794), .ZN(n7792) );
  OAI21_X1 U8764 ( .B1(n14677), .B2(n7803), .A(n7801), .ZN(n14656) );
  NAND2_X1 U8765 ( .A1(n7783), .A2(n12304), .ZN(n12306) );
  NAND2_X1 U8766 ( .A1(n7824), .A2(n7823), .ZN(n11485) );
  XNOR2_X1 U8767 ( .A(n14456), .B(n14457), .ZN(n14700) );
  OR2_X1 U8768 ( .A1(n10578), .A2(n10569), .ZN(n14711) );
  NAND2_X1 U8769 ( .A1(n7418), .A2(n7174), .ZN(n12950) );
  AOI21_X1 U8770 ( .B1(n7421), .B2(n12850), .A(n7420), .ZN(n7419) );
  AND2_X1 U8771 ( .A1(n12935), .A2(n8100), .ZN(n12936) );
  OAI21_X1 U8772 ( .B1(n14950), .B2(n9988), .A(n9916), .ZN(n14722) );
  NOR2_X1 U8773 ( .A1(n9636), .A2(n9635), .ZN(n9639) );
  AND2_X1 U8774 ( .A1(n9742), .A2(n9768), .ZN(n10432) );
  OR2_X1 U8775 ( .A1(n10355), .A2(n10353), .ZN(n15564) );
  INV_X1 U8776 ( .A(n7666), .ZN(n15062) );
  OR2_X1 U8777 ( .A1(n15415), .A2(n10581), .ZN(n15051) );
  NAND2_X1 U8778 ( .A1(n10225), .A2(n7321), .ZN(n14848) );
  INV_X1 U8779 ( .A(n7322), .ZN(n7321) );
  OAI21_X1 U8780 ( .B1(n14858), .B2(n15874), .A(n14596), .ZN(n7322) );
  NAND2_X1 U8781 ( .A1(n14910), .A2(n9938), .ZN(n14889) );
  NAND2_X1 U8782 ( .A1(n7956), .A2(n10039), .ZN(n14902) );
  NAND2_X1 U8783 ( .A1(n14916), .A2(n14915), .ZN(n7956) );
  AND2_X1 U8784 ( .A1(n14963), .A2(n9906), .ZN(n14944) );
  NAND2_X1 U8785 ( .A1(n14992), .A2(n9880), .ZN(n14979) );
  NAND2_X1 U8786 ( .A1(n15134), .A2(n10031), .ZN(n14976) );
  NOR2_X1 U8787 ( .A1(n7908), .A2(n7907), .ZN(n14993) );
  INV_X1 U8788 ( .A(n9867), .ZN(n7907) );
  NAND2_X1 U8789 ( .A1(n9856), .A2(n9855), .ZN(n15142) );
  NAND2_X1 U8790 ( .A1(n9842), .A2(n9841), .ZN(n15150) );
  NAND2_X1 U8791 ( .A1(n11963), .A2(n9811), .ZN(n12069) );
  AND2_X1 U8792 ( .A1(n11559), .A2(n10022), .ZN(n11575) );
  NAND2_X1 U8793 ( .A1(n11559), .A2(n7946), .ZN(n11574) );
  NAND2_X1 U8794 ( .A1(n7927), .A2(n11508), .ZN(n11584) );
  NAND2_X1 U8795 ( .A1(n11508), .A2(n9767), .ZN(n11582) );
  INV_X1 U8796 ( .A(n10810), .ZN(n11047) );
  NAND2_X1 U8797 ( .A1(n7942), .A2(n10012), .ZN(n11080) );
  NAND2_X1 U8798 ( .A1(n7896), .A2(n7897), .ZN(n10687) );
  NAND2_X1 U8799 ( .A1(n7901), .A2(n7902), .ZN(n11220) );
  INV_X1 U8800 ( .A(n15942), .ZN(n15887) );
  INV_X1 U8801 ( .A(n15057), .ZN(n15935) );
  INV_X1 U8802 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n7353) );
  INV_X1 U8803 ( .A(n14967), .ZN(n15403) );
  INV_X1 U8804 ( .A(n12760), .ZN(n15943) );
  INV_X1 U8805 ( .A(n12749), .ZN(n11499) );
  NAND2_X1 U8806 ( .A1(n9394), .A2(n9382), .ZN(n9385) );
  NAND2_X1 U8807 ( .A1(n9394), .A2(n9393), .ZN(n15427) );
  INV_X1 U8808 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9608) );
  NAND2_X1 U8809 ( .A1(n15421), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7937) );
  NAND2_X1 U8810 ( .A1(n7315), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7936) );
  NAND2_X1 U8811 ( .A1(n9607), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7961) );
  XNOR2_X1 U8812 ( .A(n9425), .B(n9424), .ZN(n15428) );
  NAND2_X1 U8813 ( .A1(n10068), .A2(n9595), .ZN(n7962) );
  AND2_X1 U8814 ( .A1(n7964), .A2(n9607), .ZN(n7963) );
  INV_X1 U8815 ( .A(n10091), .ZN(n15438) );
  INV_X1 U8816 ( .A(n10083), .ZN(n12458) );
  NAND2_X1 U8817 ( .A1(n9303), .A2(n9302), .ZN(n9305) );
  OR3_X1 U8818 ( .A1(n10001), .A2(P1_IR_REG_22__SCAN_IN), .A3(n15420), .ZN(
        n7436) );
  XNOR2_X1 U8819 ( .A(n9582), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15444) );
  NAND2_X1 U8820 ( .A1(n9211), .A2(n9228), .ZN(n11975) );
  INV_X1 U8821 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11572) );
  INV_X1 U8822 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11424) );
  INV_X1 U8823 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11293) );
  NAND2_X1 U8824 ( .A1(n9112), .A2(n9090), .ZN(n10764) );
  NAND2_X1 U8825 ( .A1(n9086), .A2(n9085), .ZN(n9089) );
  OR2_X1 U8826 ( .A1(n9010), .A2(n9009), .ZN(n9011) );
  INV_X1 U8827 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10434) );
  NAND2_X1 U8828 ( .A1(n8989), .A2(n8988), .ZN(n9006) );
  INV_X1 U8829 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10370) );
  OR2_X1 U8830 ( .A1(n8964), .A2(n8963), .ZN(n8965) );
  INV_X1 U8831 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10322) );
  INV_X1 U8832 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10315) );
  NAND2_X1 U8833 ( .A1(n8044), .A2(n8822), .ZN(n8823) );
  NAND2_X1 U8834 ( .A1(n8046), .A2(n8822), .ZN(n8810) );
  NOR2_X1 U8835 ( .A1(n15574), .A2(n7606), .ZN(n15571) );
  AND2_X1 U8836 ( .A1(n15749), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n7606) );
  XNOR2_X1 U8837 ( .A(n7608), .B(n15574), .ZN(n15740) );
  INV_X1 U8838 ( .A(n15573), .ZN(n7608) );
  OR2_X1 U8839 ( .A1(n15571), .A2(n7605), .ZN(n15739) );
  INV_X1 U8840 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n7605) );
  NOR2_X1 U8841 ( .A1(n15740), .A2(n15739), .ZN(n15738) );
  XNOR2_X1 U8842 ( .A(n7310), .B(n15595), .ZN(n15587) );
  INV_X1 U8843 ( .A(n15594), .ZN(n7310) );
  AND2_X1 U8844 ( .A1(n7613), .A2(n7611), .ZN(n15736) );
  NAND2_X1 U8845 ( .A1(n15632), .A2(n15633), .ZN(n15644) );
  NAND2_X1 U8846 ( .A1(n15659), .A2(n15658), .ZN(n15660) );
  XNOR2_X1 U8847 ( .A(n15670), .B(n7615), .ZN(n15665) );
  INV_X1 U8848 ( .A(n15671), .ZN(n7615) );
  OAI21_X1 U8849 ( .B1(n15678), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n15677), .ZN(
        n15686) );
  NAND2_X1 U8850 ( .A1(n15686), .A2(n15685), .ZN(n15687) );
  NOR2_X1 U8851 ( .A1(n15694), .A2(n15693), .ZN(n15695) );
  NAND2_X1 U8852 ( .A1(n15699), .A2(n15698), .ZN(n15711) );
  NOR2_X1 U8853 ( .A1(n15717), .A2(n15716), .ZN(n15726) );
  NOR2_X1 U8854 ( .A1(n11328), .A2(n7448), .ZN(n11330) );
  CLKBUF_X1 U8855 ( .A(n11323), .Z(n11324) );
  CLKBUF_X1 U8856 ( .A(n11433), .Z(n11317) );
  AND2_X1 U8857 ( .A1(n13219), .A2(n7275), .ZN(n7363) );
  NAND2_X1 U8858 ( .A1(n7446), .A2(n7445), .ZN(P3_U3491) );
  NAND2_X1 U8859 ( .A1(P3_U3897), .A2(n7450), .ZN(n7445) );
  OR2_X1 U8860 ( .A1(P3_U3897), .A2(n7447), .ZN(n7446) );
  INV_X1 U8861 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n7447) );
  INV_X1 U8862 ( .A(n13339), .ZN(n13331) );
  INV_X1 U8863 ( .A(n13404), .ZN(n13598) );
  NOR2_X1 U8864 ( .A1(n8725), .A2(n8724), .ZN(n8726) );
  NOR2_X1 U8865 ( .A1(n13383), .A2(n13656), .ZN(n8725) );
  OAI21_X1 U8866 ( .B1(n13595), .B2(n8727), .A(n7301), .ZN(n13596) );
  NAND2_X1 U8867 ( .A1(n8727), .A2(n7302), .ZN(n7301) );
  INV_X1 U8868 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n7302) );
  OAI21_X1 U8869 ( .B1(n13662), .B2(n8727), .A(n7640), .ZN(P3_U3486) );
  INV_X1 U8870 ( .A(n7641), .ZN(n7640) );
  OAI22_X1 U8871 ( .A1(n13664), .A2(n13656), .B1(n16039), .B2(n13600), .ZN(
        n7641) );
  OAI21_X1 U8872 ( .B1(n9580), .B2(n16048), .A(n9579), .ZN(P3_U3455) );
  INV_X1 U8873 ( .A(n9578), .ZN(n9579) );
  OAI22_X1 U8874 ( .A1(n13597), .A2(n13707), .B1(n9577), .B2(n16042), .ZN(
        n9578) );
  OAI21_X1 U8875 ( .B1(n13662), .B2(n16048), .A(n7569), .ZN(P3_U3454) );
  AOI21_X1 U8876 ( .B1(n8660), .B2(n16049), .A(n7570), .ZN(n7569) );
  NOR2_X1 U8877 ( .A1(n16042), .A2(n13663), .ZN(n7570) );
  OAI21_X1 U8878 ( .B1(n9365), .B2(n7178), .A(n7730), .ZN(n7729) );
  NAND2_X1 U8879 ( .A1(n7500), .A2(n7499), .ZN(P2_U3531) );
  NAND2_X1 U8880 ( .A1(P2_U3947), .A2(n9548), .ZN(n7499) );
  OR2_X1 U8881 ( .A1(P2_U3947), .A2(n8808), .ZN(n7500) );
  NAND2_X1 U8882 ( .A1(n7601), .A2(n7599), .ZN(P2_U3530) );
  AOI21_X1 U8883 ( .B1(n14295), .B2(n14300), .A(n7600), .ZN(n7599) );
  NAND2_X1 U8884 ( .A1(n14372), .A2(n16035), .ZN(n7601) );
  NOR2_X1 U8885 ( .A1(n16035), .A2(n9390), .ZN(n7600) );
  NOR2_X1 U8886 ( .A1(n8076), .A2(n7277), .ZN(n8075) );
  NOR2_X1 U8887 ( .A1(n16035), .A2(n10217), .ZN(n8076) );
  NAND2_X1 U8888 ( .A1(n7314), .A2(n7311), .ZN(P2_U3498) );
  INV_X1 U8889 ( .A(n7312), .ZN(n7311) );
  NAND2_X1 U8890 ( .A1(n14372), .A2(n14371), .ZN(n7314) );
  OAI22_X1 U8891 ( .A1(n14373), .A2(n14402), .B1(n14371), .B2(n7313), .ZN(
        n7312) );
  AND2_X1 U8892 ( .A1(n10728), .A2(n10727), .ZN(n10729) );
  NAND2_X1 U8893 ( .A1(n10099), .A2(n10229), .ZN(n10100) );
  OR2_X1 U8894 ( .A1(n16014), .A2(n10228), .ZN(n7361) );
  NAND2_X1 U8895 ( .A1(n14599), .A2(n10229), .ZN(n10230) );
  NAND2_X1 U8896 ( .A1(n7664), .A2(n7663), .ZN(n7662) );
  NAND2_X1 U8897 ( .A1(n7917), .A2(n7353), .ZN(n7352) );
  NAND2_X1 U8898 ( .A1(n7917), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7916) );
  INV_X1 U8899 ( .A(n7614), .ZN(n15601) );
  INV_X1 U8900 ( .A(n7613), .ZN(n15609) );
  INV_X1 U8901 ( .A(n15633), .ZN(n15630) );
  XNOR2_X1 U8902 ( .A(n7620), .B(n7618), .ZN(SUB_1596_U4) );
  XNOR2_X1 U8903 ( .A(n15733), .B(n7619), .ZN(n7618) );
  AOI21_X1 U8904 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n15728), .A(n15727), .ZN(
        n7620) );
  XNOR2_X1 U8905 ( .A(n7296), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n7619) );
  INV_X2 U8906 ( .A(n14590), .ZN(n14442) );
  INV_X2 U8907 ( .A(n14590), .ZN(n14509) );
  OR2_X1 U8908 ( .A1(n7995), .A2(n13762), .ZN(n7159) );
  AND2_X1 U8909 ( .A1(n9289), .A2(n9288), .ZN(n14162) );
  INV_X1 U8910 ( .A(n14162), .ZN(n14336) );
  CLKBUF_X3 U8911 ( .A(n8816), .Z(n8883) );
  NOR2_X1 U8912 ( .A1(n12307), .A2(n7782), .ZN(n7160) );
  CLKBUF_X1 U8913 ( .A(n9419), .Z(n9484) );
  INV_X2 U8914 ( .A(n8883), .ZN(n9489) );
  NOR2_X1 U8915 ( .A1(n14195), .A2(n14210), .ZN(n7161) );
  AND2_X2 U8916 ( .A1(n12484), .A2(n14405), .ZN(n8793) );
  INV_X1 U8917 ( .A(n14097), .ZN(n7483) );
  NAND2_X1 U8918 ( .A1(n7793), .A2(n14519), .ZN(n7162) );
  INV_X1 U8919 ( .A(n11312), .ZN(n11430) );
  AND2_X1 U8920 ( .A1(n11960), .A2(n10025), .ZN(n7163) );
  OR2_X1 U8921 ( .A1(n7186), .A2(n7560), .ZN(n7164) );
  AND2_X1 U8922 ( .A1(n7588), .A2(n14162), .ZN(n7165) );
  OR2_X1 U8923 ( .A1(n14252), .A2(n8011), .ZN(n7166) );
  AND2_X1 U8924 ( .A1(n7884), .A2(n7882), .ZN(n7167) );
  AND2_X1 U8925 ( .A1(n15943), .A2(n7671), .ZN(n7168) );
  AND2_X1 U8926 ( .A1(n13006), .A2(n7707), .ZN(n7169) );
  INV_X1 U8927 ( .A(n11250), .ZN(n10642) );
  AND3_X1 U8928 ( .A1(n7540), .A2(n7543), .A3(n7402), .ZN(n7170) );
  INV_X1 U8929 ( .A(n14355), .ZN(n14220) );
  AND3_X1 U8930 ( .A1(n12811), .A2(n12810), .A3(n7257), .ZN(n7171) );
  NOR3_X1 U8931 ( .A1(n9562), .A2(n10183), .A3(n14420), .ZN(n7172) );
  AND3_X1 U8932 ( .A1(n12795), .A2(n12794), .A3(n7258), .ZN(n7173) );
  INV_X1 U8933 ( .A(n11856), .ZN(n13251) );
  AND4_X1 U8934 ( .A1(n8259), .A2(n8258), .A3(n8257), .A4(n8256), .ZN(n11856)
         );
  OR2_X1 U8935 ( .A1(n7421), .A2(n12850), .ZN(n7174) );
  AND2_X1 U8936 ( .A1(n8146), .A2(n7894), .ZN(n7893) );
  INV_X1 U8937 ( .A(n7893), .ZN(n7716) );
  AND2_X1 U8938 ( .A1(n7825), .A2(n9868), .ZN(n7175) );
  INV_X1 U8939 ( .A(n7995), .ZN(n7994) );
  OR2_X1 U8940 ( .A1(n13897), .A2(n13767), .ZN(n7995) );
  AND2_X1 U8941 ( .A1(n7669), .A2(n7668), .ZN(n7176) );
  INV_X1 U8942 ( .A(n16020), .ZN(n12382) );
  AND2_X1 U8943 ( .A1(n7767), .A2(n7768), .ZN(n7177) );
  OR2_X1 U8944 ( .A1(n7736), .A2(n10264), .ZN(n7178) );
  OR2_X1 U8945 ( .A1(n13586), .A2(n7639), .ZN(n7179) );
  INV_X1 U8946 ( .A(n12797), .ZN(n7869) );
  AND2_X1 U8947 ( .A1(n8585), .A2(n8584), .ZN(n13396) );
  INV_X1 U8948 ( .A(n13396), .ZN(n7563) );
  OR2_X1 U8949 ( .A1(n13480), .A2(n13461), .ZN(n13003) );
  INV_X1 U8950 ( .A(n13003), .ZN(n7462) );
  INV_X1 U8951 ( .A(n12816), .ZN(n7865) );
  INV_X1 U8952 ( .A(n12896), .ZN(n7952) );
  AND2_X1 U8953 ( .A1(n14216), .A2(n7165), .ZN(n7180) );
  AND2_X1 U8954 ( .A1(n8542), .A2(n8541), .ZN(n13462) );
  AND2_X1 U8955 ( .A1(n9287), .A2(SI_21_), .ZN(n7181) );
  INV_X1 U8956 ( .A(n11730), .ZN(n7490) );
  AND2_X1 U8957 ( .A1(n8519), .A2(n7680), .ZN(n7182) );
  OR2_X1 U8958 ( .A1(n12227), .A2(n12568), .ZN(n7183) );
  AND2_X1 U8959 ( .A1(n11546), .A2(n13925), .ZN(n7184) );
  AND2_X1 U8960 ( .A1(n8119), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7185) );
  AND2_X1 U8961 ( .A1(n10322), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7186) );
  AND2_X1 U8962 ( .A1(n7842), .A2(n13462), .ZN(n7187) );
  AOI21_X1 U8963 ( .B1(n14111), .B2(n10177), .A(n10176), .ZN(n14098) );
  AND2_X1 U8964 ( .A1(n14953), .A2(n7176), .ZN(n7188) );
  NOR2_X2 U8965 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8800) );
  NAND2_X1 U8966 ( .A1(n8981), .A2(n8980), .ZN(n7189) );
  OR2_X1 U8967 ( .A1(n10218), .A2(n9981), .ZN(n7190) );
  INV_X1 U8968 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7505) );
  AND2_X1 U8969 ( .A1(n12560), .A2(n12561), .ZN(n12661) );
  AND2_X1 U8970 ( .A1(n14994), .A2(n9867), .ZN(n7191) );
  OR2_X1 U8971 ( .A1(n7955), .A2(n10040), .ZN(n7192) );
  OAI21_X1 U8972 ( .B1(n8311), .B2(n7186), .A(n8326), .ZN(n7562) );
  AND2_X1 U8973 ( .A1(n11879), .A2(n7974), .ZN(n7193) );
  AND2_X1 U8974 ( .A1(n9626), .A2(n9589), .ZN(n9628) );
  OR2_X1 U8975 ( .A1(n8472), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n7195) );
  AND2_X1 U8976 ( .A1(n8226), .A2(n8228), .ZN(n7196) );
  INV_X1 U8977 ( .A(n12634), .ZN(n7454) );
  INV_X1 U8978 ( .A(n7524), .ZN(n8598) );
  AND2_X1 U8979 ( .A1(n10168), .A2(n10166), .ZN(n7197) );
  NAND2_X1 U8980 ( .A1(n8749), .A2(n8748), .ZN(n8852) );
  NAND2_X1 U8981 ( .A1(n8059), .A2(n8057), .ZN(n9286) );
  INV_X1 U8982 ( .A(n7970), .ZN(n7969) );
  OR2_X1 U8983 ( .A1(n13885), .A2(n7971), .ZN(n7970) );
  INV_X1 U8984 ( .A(n11938), .ZN(n7597) );
  OR2_X1 U8985 ( .A1(n14098), .A2(n14097), .ZN(n7198) );
  INV_X1 U8986 ( .A(n12532), .ZN(n7632) );
  AND2_X1 U8987 ( .A1(n14561), .A2(n14730), .ZN(n7199) );
  XOR2_X1 U8988 ( .A(n14331), .B(n13916), .Z(n7200) );
  AND2_X1 U8989 ( .A1(n7753), .A2(n9283), .ZN(n7201) );
  AND3_X1 U8990 ( .A1(n10180), .A2(n7327), .A3(n7326), .ZN(n7202) );
  AND4_X1 U8991 ( .A1(n8678), .A2(n8607), .A3(n8610), .A4(n8602), .ZN(n7203)
         );
  OR2_X1 U8992 ( .A1(n7724), .A2(n7727), .ZN(n7204) );
  OR2_X1 U8993 ( .A1(n14195), .A2(n13918), .ZN(n7205) );
  AND2_X1 U8994 ( .A1(n7454), .A2(n12635), .ZN(n7206) );
  AND2_X1 U8995 ( .A1(n9256), .A2(n9255), .ZN(n14195) );
  OR2_X1 U8996 ( .A1(n9299), .A2(n9298), .ZN(n7207) );
  OR2_X1 U8997 ( .A1(n9152), .A2(n9151), .ZN(n7208) );
  OR2_X1 U8998 ( .A1(n12729), .A2(n14740), .ZN(n7209) );
  AND2_X1 U8999 ( .A1(n12694), .A2(n12655), .ZN(n7210) );
  AND2_X1 U9000 ( .A1(n12773), .A2(n14733), .ZN(n7211) );
  NAND2_X1 U9001 ( .A1(n9830), .A2(n9829), .ZN(n15413) );
  INV_X1 U9002 ( .A(n12902), .ZN(n14885) );
  INV_X1 U9003 ( .A(n8047), .ZN(n8809) );
  NOR2_X1 U9004 ( .A1(n14140), .A2(n8035), .ZN(n7212) );
  AND2_X1 U9005 ( .A1(n11484), .A2(n11483), .ZN(n7213) );
  INV_X1 U9006 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9605) );
  AND2_X1 U9007 ( .A1(n15150), .A2(n10028), .ZN(n7214) );
  INV_X1 U9008 ( .A(n13868), .ZN(n13916) );
  NOR2_X1 U9009 ( .A1(n12012), .A2(n12013), .ZN(n7215) );
  INV_X1 U9010 ( .A(n7804), .ZN(n7803) );
  NOR2_X1 U9011 ( .A1(n14486), .A2(n7805), .ZN(n7804) );
  OR2_X1 U9012 ( .A1(n13324), .A2(n13332), .ZN(n7216) );
  AND2_X1 U9013 ( .A1(n8072), .A2(n8073), .ZN(n7217) );
  INV_X1 U9014 ( .A(n15880), .ZN(n15888) );
  AND2_X1 U9015 ( .A1(n8500), .A2(n12608), .ZN(n7218) );
  INV_X1 U9016 ( .A(n12787), .ZN(n7887) );
  OR2_X1 U9017 ( .A1(n10864), .A2(n11411), .ZN(n7219) );
  INV_X1 U9018 ( .A(n12813), .ZN(n7888) );
  AND2_X1 U9019 ( .A1(n7952), .A2(n10033), .ZN(n7220) );
  NAND2_X1 U9020 ( .A1(n13426), .A2(n7624), .ZN(n7221) );
  AND2_X1 U9021 ( .A1(n7888), .A2(n12812), .ZN(n7222) );
  AND2_X1 U9022 ( .A1(n8079), .A2(n9111), .ZN(n7223) );
  AND2_X1 U9023 ( .A1(n12556), .A2(n12557), .ZN(n12662) );
  AND2_X1 U9024 ( .A1(n12800), .A2(n7868), .ZN(n7224) );
  NOR2_X1 U9025 ( .A1(n7482), .A2(n14116), .ZN(n7225) );
  INV_X1 U9026 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7592) );
  OR2_X1 U9027 ( .A1(n12968), .A2(n7535), .ZN(n7226) );
  NAND2_X1 U9028 ( .A1(n12542), .A2(n12543), .ZN(n15849) );
  INV_X1 U9029 ( .A(n15849), .ZN(n8239) );
  AND2_X1 U9030 ( .A1(n8933), .A2(n8934), .ZN(n7227) );
  AND2_X1 U9031 ( .A1(n15898), .A2(n12721), .ZN(n7228) );
  NOR2_X1 U9032 ( .A1(n12639), .A2(n12635), .ZN(n7229) );
  AND2_X1 U9033 ( .A1(n7713), .A2(n8654), .ZN(n7230) );
  INV_X1 U9034 ( .A(n7984), .ZN(n7983) );
  NAND2_X1 U9035 ( .A1(n11058), .A2(n10822), .ZN(n7984) );
  NOR2_X1 U9036 ( .A1(n12203), .A2(n12144), .ZN(n7231) );
  NOR2_X1 U9037 ( .A1(n14134), .A2(n13828), .ZN(n7232) );
  NOR2_X1 U9038 ( .A1(n14743), .A2(n15835), .ZN(n7233) );
  AND2_X1 U9039 ( .A1(n14974), .A2(n10033), .ZN(n7234) );
  INV_X1 U9040 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8950) );
  OR2_X1 U9041 ( .A1(n8598), .A2(n8148), .ZN(n7235) );
  INV_X1 U9042 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9868) );
  NAND2_X1 U9043 ( .A1(n7565), .A2(n8577), .ZN(n12518) );
  INV_X1 U9044 ( .A(n12518), .ZN(n7564) );
  INV_X1 U9045 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8344) );
  AND2_X1 U9046 ( .A1(n12824), .A2(n12823), .ZN(n7236) );
  AND2_X1 U9047 ( .A1(n7991), .A2(n10297), .ZN(n7237) );
  NOR2_X1 U9048 ( .A1(n12801), .A2(n12803), .ZN(n7238) );
  NAND2_X1 U9049 ( .A1(n14228), .A2(n14209), .ZN(n7239) );
  AND2_X1 U9050 ( .A1(n9654), .A2(n9655), .ZN(n7240) );
  AND2_X1 U9051 ( .A1(n7931), .A2(n7932), .ZN(n7241) );
  INV_X1 U9052 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8151) );
  AND2_X1 U9053 ( .A1(n10139), .A2(n14049), .ZN(n14062) );
  INV_X1 U9054 ( .A(n14331), .ZN(n14149) );
  NAND2_X1 U9055 ( .A1(n8080), .A2(n9306), .ZN(n14331) );
  AND2_X1 U9056 ( .A1(n9060), .A2(n15275), .ZN(n7242) );
  OR2_X1 U9057 ( .A1(n12580), .A2(n8394), .ZN(n7243) );
  AND2_X1 U9058 ( .A1(n10370), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7244) );
  INV_X1 U9059 ( .A(n12588), .ZN(n7639) );
  AND2_X1 U9060 ( .A1(n12519), .A2(n8573), .ZN(n13427) );
  NOR2_X1 U9061 ( .A1(n14485), .A2(n14484), .ZN(n7245) );
  NAND2_X1 U9062 ( .A1(n7564), .A2(n7563), .ZN(n12521) );
  INV_X1 U9063 ( .A(n13743), .ZN(n7967) );
  INV_X1 U9064 ( .A(n12739), .ZN(n7856) );
  INV_X1 U9065 ( .A(n12841), .ZN(n7849) );
  INV_X1 U9066 ( .A(n9003), .ZN(n7767) );
  NAND2_X1 U9067 ( .A1(n12640), .A2(n12634), .ZN(n12678) );
  INV_X1 U9068 ( .A(n12678), .ZN(n7543) );
  AND2_X1 U9069 ( .A1(n10023), .A2(n12886), .ZN(n7246) );
  INV_X1 U9070 ( .A(n12892), .ZN(n12071) );
  AND2_X1 U9071 ( .A1(n11721), .A2(n11724), .ZN(n7247) );
  AND2_X1 U9072 ( .A1(n12738), .A2(n10013), .ZN(n7248) );
  AND2_X1 U9073 ( .A1(n7992), .A2(n13845), .ZN(n7249) );
  AND2_X1 U9074 ( .A1(n12981), .A2(n12980), .ZN(n7250) );
  NOR2_X1 U9075 ( .A1(n8653), .A2(n7714), .ZN(n7251) );
  INV_X1 U9076 ( .A(n10119), .ZN(n7551) );
  AND2_X1 U9077 ( .A1(n14925), .A2(n9928), .ZN(n7252) );
  AND2_X1 U9078 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(n9999), .ZN(n7253) );
  NAND2_X1 U9079 ( .A1(n15600), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n7254) );
  NAND2_X1 U9080 ( .A1(n11938), .A2(n13922), .ZN(n7255) );
  OR2_X1 U9081 ( .A1(n7887), .A2(n12786), .ZN(n7256) );
  OR2_X1 U9082 ( .A1(n7888), .A2(n12812), .ZN(n7257) );
  OR2_X1 U9083 ( .A1(n7869), .A2(n12796), .ZN(n7258) );
  AND2_X1 U9084 ( .A1(n7808), .A2(n11761), .ZN(n7259) );
  AND2_X1 U9085 ( .A1(n13422), .A2(n8654), .ZN(n7260) );
  OR2_X1 U9086 ( .A1(n12761), .A2(n12763), .ZN(n7261) );
  OR2_X1 U9087 ( .A1(n12774), .A2(n12776), .ZN(n7262) );
  AND2_X1 U9088 ( .A1(n7456), .A2(n12659), .ZN(n7263) );
  AND2_X1 U9089 ( .A1(n12229), .A2(n7183), .ZN(n7264) );
  AND2_X1 U9090 ( .A1(n8659), .A2(n8657), .ZN(n7265) );
  AND2_X1 U9091 ( .A1(n8012), .A2(n7505), .ZN(n7266) );
  INV_X1 U9092 ( .A(n14897), .ZN(n15392) );
  NAND2_X1 U9093 ( .A1(n9940), .A2(n9939), .ZN(n14897) );
  INV_X1 U9094 ( .A(n7464), .ZN(n7463) );
  OAI21_X1 U9095 ( .B1(n13489), .B2(n7465), .A(n13005), .ZN(n7464) );
  INV_X1 U9096 ( .A(n7879), .ZN(n7878) );
  NAND2_X1 U9097 ( .A1(n7880), .A2(n7884), .ZN(n7879) );
  NAND2_X1 U9098 ( .A1(n8863), .A2(n8864), .ZN(n7267) );
  OR2_X1 U9099 ( .A1(n7772), .A2(n7771), .ZN(n7268) );
  INV_X1 U9100 ( .A(n10176), .ZN(n7489) );
  INV_X1 U9101 ( .A(n7928), .ZN(n7927) );
  NAND2_X1 U9102 ( .A1(n7929), .A2(n9767), .ZN(n7928) );
  INV_X1 U9103 ( .A(n14127), .ZN(n8034) );
  NAND2_X1 U9104 ( .A1(n9930), .A2(n9929), .ZN(n14905) );
  INV_X1 U9105 ( .A(n14905), .ZN(n7668) );
  INV_X1 U9106 ( .A(n12576), .ZN(n7634) );
  NAND2_X1 U9107 ( .A1(n7633), .A2(n7631), .ZN(n12362) );
  NAND2_X1 U9108 ( .A1(n9413), .A2(n9412), .ZN(n14060) );
  INV_X1 U9109 ( .A(n14060), .ZN(n7594) );
  NOR2_X1 U9110 ( .A1(n13644), .A2(n13565), .ZN(n7269) );
  AND2_X1 U9111 ( .A1(n11867), .A2(n7676), .ZN(n7270) );
  OAI21_X1 U9112 ( .B1(n10121), .B2(n7650), .A(n7648), .ZN(n12134) );
  NAND2_X1 U9113 ( .A1(n7549), .A2(n10119), .ZN(n11772) );
  NAND2_X1 U9114 ( .A1(n10121), .A2(n10120), .ZN(n12006) );
  INV_X1 U9115 ( .A(n13549), .ZN(n13558) );
  AND2_X1 U9116 ( .A1(n13480), .A2(n13493), .ZN(n7271) );
  INV_X1 U9117 ( .A(n12619), .ZN(n7465) );
  AND2_X1 U9118 ( .A1(n7883), .A2(n7882), .ZN(n7272) );
  AND2_X1 U9119 ( .A1(n7625), .A2(n7629), .ZN(n7273) );
  INV_X1 U9120 ( .A(n13913), .ZN(n13829) );
  AND3_X1 U9121 ( .A1(n9148), .A2(n9147), .A3(n9146), .ZN(n12401) );
  INV_X1 U9122 ( .A(n12401), .ZN(n14273) );
  NAND2_X1 U9123 ( .A1(n9866), .A2(n9865), .ZN(n15011) );
  INV_X1 U9124 ( .A(n15011), .ZN(n7908) );
  INV_X1 U9125 ( .A(n14238), .ZN(n14188) );
  AND2_X1 U9126 ( .A1(n9239), .A2(n9238), .ZN(n14238) );
  AND2_X1 U9127 ( .A1(n15044), .A2(n10027), .ZN(n7274) );
  NAND2_X1 U9128 ( .A1(n14216), .A2(n7588), .ZN(n7589) );
  OR2_X1 U9129 ( .A1(n7564), .A2(n13234), .ZN(n7275) );
  NOR2_X1 U9130 ( .A1(n9284), .A2(n8055), .ZN(n8054) );
  INV_X1 U9131 ( .A(n8031), .ZN(n8030) );
  NOR2_X1 U9132 ( .A1(n8035), .A2(n8034), .ZN(n8031) );
  AND2_X1 U9133 ( .A1(n7815), .A2(n7813), .ZN(n7276) );
  NOR2_X1 U9134 ( .A1(n7594), .A2(n14369), .ZN(n7277) );
  INV_X1 U9135 ( .A(n7990), .ZN(n12408) );
  NOR2_X1 U9136 ( .A1(n12344), .A2(n12345), .ZN(n7990) );
  AND2_X1 U9137 ( .A1(n12967), .A2(n13245), .ZN(n7278) );
  INV_X1 U9138 ( .A(n8660), .ZN(n13664) );
  NAND2_X1 U9139 ( .A1(n8196), .A2(n8195), .ZN(n8660) );
  AND2_X1 U9140 ( .A1(n11293), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7279) );
  INV_X1 U9141 ( .A(n8058), .ZN(n8057) );
  NOR2_X1 U9142 ( .A1(n9270), .A2(n15191), .ZN(n8058) );
  OR2_X1 U9143 ( .A1(n15387), .A2(n15402), .ZN(n7280) );
  OR2_X1 U9144 ( .A1(n9269), .A2(SI_20_), .ZN(n7281) );
  INV_X1 U9145 ( .A(n9226), .ZN(n7742) );
  OR2_X1 U9146 ( .A1(n13597), .A2(n13397), .ZN(n7282) );
  OR2_X1 U9147 ( .A1(n15387), .A2(n15125), .ZN(n7283) );
  INV_X1 U9148 ( .A(n13449), .ZN(n13474) );
  AND2_X1 U9149 ( .A1(n8530), .A2(n8529), .ZN(n13449) );
  INV_X1 U9150 ( .A(n13462), .ZN(n13239) );
  AND2_X1 U9151 ( .A1(n13586), .A2(n8638), .ZN(n7284) );
  AND2_X1 U9152 ( .A1(n10232), .A2(n7916), .ZN(n7285) );
  AND2_X1 U9153 ( .A1(n10230), .A2(n7361), .ZN(n7286) );
  INV_X1 U9154 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7369) );
  NAND2_X1 U9155 ( .A1(n16042), .A2(n15907), .ZN(n13707) );
  NAND2_X1 U9156 ( .A1(n7838), .A2(n8691), .ZN(n11307) );
  INV_X1 U9157 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7694) );
  AND2_X1 U9158 ( .A1(n7693), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7287) );
  XOR2_X1 U9159 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .Z(n7288) );
  INV_X1 U9160 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7692) );
  OAI21_X1 U9161 ( .B1(n11879), .B2(n7977), .A(n7974), .ZN(n12056) );
  INV_X1 U9162 ( .A(n15150), .ZN(n7673) );
  INV_X1 U9163 ( .A(n7631), .ZN(n7630) );
  XNOR2_X1 U9164 ( .A(n9305), .B(n9304), .ZN(n14418) );
  NAND2_X1 U9165 ( .A1(n7289), .A2(n7680), .ZN(n7566) );
  OR2_X1 U9166 ( .A1(n8533), .A2(n7567), .ZN(n7289) );
  INV_X1 U9167 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7682) );
  NAND2_X1 U9168 ( .A1(n10210), .A2(n10183), .ZN(n7290) );
  AND2_X1 U9169 ( .A1(n11642), .A2(n8000), .ZN(n7291) );
  AND2_X1 U9170 ( .A1(n13309), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n7292) );
  INV_X1 U9171 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11976) );
  INV_X1 U9172 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12463) );
  INV_X1 U9173 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n12067) );
  AND2_X1 U9174 ( .A1(n7182), .A2(n7394), .ZN(n7293) );
  AND2_X1 U9175 ( .A1(n7824), .A2(n11296), .ZN(n7294) );
  AND2_X2 U9176 ( .A1(n10103), .A2(n10102), .ZN(n16017) );
  INV_X1 U9177 ( .A(n16017), .ZN(n7917) );
  INV_X1 U9178 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7394) );
  INV_X1 U9179 ( .A(n15827), .ZN(n7429) );
  INV_X1 U9180 ( .A(n12764), .ZN(n7671) );
  INV_X1 U9181 ( .A(n12753), .ZN(n7659) );
  NAND2_X1 U9182 ( .A1(n12697), .A2(n12536), .ZN(n12635) );
  NAND2_X1 U9183 ( .A1(n15855), .A2(n15972), .ZN(n13658) );
  AND2_X2 U9184 ( .A1(n10215), .A2(n10251), .ZN(n16035) );
  INV_X1 U9185 ( .A(n11077), .ZN(n7661) );
  INV_X1 U9186 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12481) );
  AND2_X1 U9187 ( .A1(n10859), .A2(n7576), .ZN(n7295) );
  XOR2_X1 U9188 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n7296) );
  INV_X1 U9189 ( .A(SI_2_), .ZN(n7319) );
  INV_X1 U9190 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7678) );
  INV_X1 U9191 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8807) );
  INV_X1 U9192 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7617) );
  INV_X1 U9193 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7610) );
  INV_X1 U9194 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7607) );
  NAND2_X1 U9195 ( .A1(n7362), .A2(n9989), .ZN(n7351) );
  XOR2_X1 U9196 ( .A(n13285), .B(n13286), .Z(n13259) );
  NAND2_X1 U9197 ( .A1(n13255), .A2(n13285), .ZN(n13273) );
  INV_X1 U9198 ( .A(n13285), .ZN(n7580) );
  NAND2_X1 U9199 ( .A1(n10864), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8211) );
  INV_X1 U9200 ( .A(n7299), .ZN(n15799) );
  NAND2_X1 U9201 ( .A1(n15778), .A2(n7586), .ZN(n7299) );
  NAND2_X1 U9202 ( .A1(n15809), .A2(n11816), .ZN(n11818) );
  NAND2_X1 U9203 ( .A1(n15772), .A2(n11812), .ZN(n15793) );
  NAND2_X1 U9204 ( .A1(n11022), .A2(n10856), .ZN(n7575) );
  AOI21_X1 U9205 ( .B1(n15817), .B2(P3_REG1_REG_11__SCAN_IN), .A(n11832), .ZN(
        n11833) );
  NAND2_X1 U9206 ( .A1(n13447), .A2(n13452), .ZN(n8652) );
  NAND2_X1 U9207 ( .A1(n11905), .A2(n8626), .ZN(n11904) );
  NAND2_X1 U9208 ( .A1(n12538), .A2(n12533), .ZN(n7702) );
  NAND2_X1 U9209 ( .A1(n13519), .A2(n7718), .ZN(n8646) );
  NAND3_X1 U9210 ( .A1(n7715), .A2(n7892), .A3(n8149), .ZN(n7300) );
  NAND2_X1 U9211 ( .A1(n8622), .A2(n8621), .ZN(n11336) );
  OAI21_X1 U9212 ( .B1(n12360), .B2(n8635), .A(n8634), .ZN(n12433) );
  XNOR2_X1 U9213 ( .A(n7332), .B(n12656), .ZN(n8676) );
  NAND2_X1 U9214 ( .A1(n11471), .A2(n11316), .ZN(n12538) );
  NAND2_X1 U9215 ( .A1(n8646), .A2(n8645), .ZN(n13490) );
  NAND2_X1 U9216 ( .A1(n11988), .A2(n7711), .ZN(n12238) );
  NAND2_X1 U9217 ( .A1(n9568), .A2(n7282), .ZN(n7332) );
  NAND2_X1 U9218 ( .A1(n8636), .A2(n13055), .ZN(n12472) );
  NAND2_X1 U9219 ( .A1(n8618), .A2(n8617), .ZN(n15850) );
  INV_X1 U9220 ( .A(n7525), .ZN(n7642) );
  NAND2_X1 U9221 ( .A1(n8658), .A2(n7265), .ZN(n13401) );
  NAND2_X1 U9222 ( .A1(n7704), .A2(n7705), .ZN(n13459) );
  NAND2_X1 U9223 ( .A1(n8652), .A2(n7251), .ZN(n7713) );
  NAND2_X1 U9224 ( .A1(n8633), .A2(n8632), .ZN(n12360) );
  INV_X1 U9225 ( .A(n7419), .ZN(n7418) );
  AOI21_X1 U9226 ( .B1(n7863), .B2(n7866), .A(n7862), .ZN(n7861) );
  NAND2_X1 U9227 ( .A1(n9205), .A2(SI_18_), .ZN(n9227) );
  NAND2_X1 U9228 ( .A1(n12849), .A2(n12848), .ZN(n7421) );
  INV_X1 U9229 ( .A(n12950), .ZN(n12953) );
  INV_X1 U9230 ( .A(n14934), .ZN(n7864) );
  XNOR2_X1 U9231 ( .A(n10755), .B(n13928), .ZN(n10756) );
  NAND2_X1 U9232 ( .A1(n14077), .A2(n7366), .ZN(n7365) );
  NAND2_X1 U9233 ( .A1(n10114), .A2(n10113), .ZN(n10962) );
  NAND2_X1 U9234 ( .A1(n7341), .A2(n8987), .ZN(n8990) );
  NAND2_X1 U9235 ( .A1(n14079), .A2(n14078), .ZN(n14077) );
  NAND2_X1 U9236 ( .A1(n14268), .A2(n7656), .ZN(n7552) );
  AOI21_X1 U9237 ( .B1(n13126), .B2(n13125), .A(n7247), .ZN(n11723) );
  AOI21_X2 U9238 ( .B1(n15847), .B2(n11719), .A(n11718), .ZN(n13154) );
  NAND2_X2 U9239 ( .A1(n13019), .A2(n13109), .ZN(n13111) );
  NAND2_X1 U9240 ( .A1(n13165), .A2(n13164), .ZN(n13163) );
  NAND2_X1 U9241 ( .A1(n7356), .A2(n7355), .ZN(n7843) );
  NOR2_X1 U9242 ( .A1(n11435), .A2(n11436), .ZN(n11718) );
  AOI21_X1 U9243 ( .B1(n11323), .B2(n11325), .A(n7357), .ZN(n11433) );
  NAND2_X1 U9244 ( .A1(n11917), .A2(n11916), .ZN(n11999) );
  NAND2_X1 U9245 ( .A1(n13076), .A2(n12998), .ZN(n13165) );
  NAND2_X1 U9246 ( .A1(n13153), .A2(n7307), .ZN(n13126) );
  NAND2_X1 U9247 ( .A1(n12426), .A2(n12425), .ZN(n12427) );
  NAND2_X1 U9248 ( .A1(n7304), .A2(n7250), .ZN(n7826) );
  NAND2_X1 U9249 ( .A1(n13198), .A2(n7305), .ZN(n7304) );
  NAND2_X1 U9250 ( .A1(n13154), .A2(n13155), .ZN(n13153) );
  NAND2_X1 U9251 ( .A1(n10572), .A2(n10573), .ZN(n10618) );
  NAND2_X1 U9252 ( .A1(n14602), .A2(n14603), .ZN(n14666) );
  NAND2_X1 U9253 ( .A1(n10916), .A2(n10953), .ZN(n11295) );
  INV_X1 U9254 ( .A(n12300), .ZN(n7333) );
  NAND2_X1 U9255 ( .A1(n11762), .A2(n7259), .ZN(n12030) );
  NAND2_X1 U9256 ( .A1(n7822), .A2(n7821), .ZN(n11492) );
  AOI21_X2 U9257 ( .B1(n13896), .B2(n13897), .A(n13895), .ZN(n13908) );
  NAND2_X1 U9258 ( .A1(n13816), .A2(n13815), .ZN(n13814) );
  AOI21_X1 U9259 ( .B1(n13855), .B2(n13748), .A(n13852), .ZN(n13749) );
  NAND2_X1 U9260 ( .A1(n12345), .A2(n12407), .ZN(n7989) );
  NAND2_X1 U9261 ( .A1(n13203), .A2(n12995), .ZN(n13078) );
  NAND2_X1 U9262 ( .A1(n7826), .A2(n13058), .ZN(n13059) );
  NAND2_X1 U9263 ( .A1(n7874), .A2(n7876), .ZN(n13203) );
  NAND2_X1 U9264 ( .A1(n7838), .A2(n7835), .ZN(n7308) );
  NAND2_X1 U9265 ( .A1(n14061), .A2(n16033), .ZN(n7506) );
  NAND2_X1 U9266 ( .A1(n8891), .A2(n8890), .ZN(n8895) );
  OAI21_X2 U9267 ( .B1(n7359), .B2(n7358), .A(n13747), .ZN(n13855) );
  NAND2_X1 U9268 ( .A1(n15631), .A2(n13993), .ZN(n15632) );
  OAI21_X1 U9269 ( .B1(n15711), .B2(n15710), .A(n7604), .ZN(n7309) );
  NAND2_X1 U9270 ( .A1(n15608), .A2(n15607), .ZN(n7612) );
  NAND2_X1 U9271 ( .A1(n7612), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n7611) );
  NAND2_X1 U9272 ( .A1(n14281), .A2(n16030), .ZN(n14254) );
  NAND2_X1 U9273 ( .A1(n7598), .A2(n7597), .ZN(n7596) );
  NAND2_X1 U9274 ( .A1(n7595), .A2(n7594), .ZN(n14049) );
  NAND2_X1 U9275 ( .A1(n14102), .A2(n14093), .ZN(n14089) );
  NAND2_X4 U9276 ( .A1(n8802), .A2(n10297), .ZN(n9395) );
  AND3_X2 U9277 ( .A1(n8746), .A2(n7593), .A3(n8749), .ZN(n8763) );
  AND2_X2 U9278 ( .A1(n10010), .A2(n12716), .ZN(n15873) );
  AOI21_X2 U9279 ( .B1(n15010), .B2(n15013), .A(n10030), .ZN(n14999) );
  NAND2_X1 U9280 ( .A1(n14946), .A2(n14947), .ZN(n14945) );
  INV_X4 U9281 ( .A(n10323), .ZN(n9882) );
  NAND2_X1 U9282 ( .A1(n15872), .A2(n15873), .ZN(n15871) );
  NAND2_X1 U9283 ( .A1(n11224), .A2(n12876), .ZN(n11223) );
  NAND2_X1 U9284 ( .A1(n7163), .A2(n12071), .ZN(n12070) );
  NAND3_X1 U9285 ( .A1(n9826), .A2(n9605), .A3(n9602), .ZN(n7315) );
  OAI21_X1 U9286 ( .B1(n14862), .B2(n14861), .A(n14860), .ZN(n14864) );
  NAND2_X1 U9287 ( .A1(n15075), .A2(n7283), .ZN(P1_U3555) );
  NAND2_X1 U9288 ( .A1(n15386), .A2(n7280), .ZN(P1_U3523) );
  NAND2_X1 U9289 ( .A1(n10308), .A2(n12860), .ZN(n9688) );
  NAND2_X1 U9290 ( .A1(n11863), .A2(n11862), .ZN(n11861) );
  NAND2_X1 U9291 ( .A1(n7939), .A2(n7938), .ZN(n10803) );
  NAND2_X1 U9292 ( .A1(n7318), .A2(n8841), .ZN(n8826) );
  NAND2_X1 U9293 ( .A1(n7317), .A2(n7316), .ZN(n8842) );
  INV_X1 U9294 ( .A(n8826), .ZN(n7317) );
  NAND2_X1 U9295 ( .A1(n7320), .A2(n7319), .ZN(n7318) );
  INV_X1 U9296 ( .A(n8824), .ZN(n7320) );
  INV_X1 U9297 ( .A(n8895), .ZN(n7323) );
  AND2_X2 U9298 ( .A1(n12070), .A2(n10026), .ZN(n15046) );
  NAND2_X1 U9299 ( .A1(n14876), .A2(n7960), .ZN(n14860) );
  OAI21_X1 U9300 ( .B1(n10231), .B2(n7362), .A(n7286), .ZN(P1_U3556) );
  OAI21_X1 U9301 ( .B1(n10231), .B2(n7917), .A(n7285), .ZN(P1_U3524) );
  NAND3_X1 U9302 ( .A1(n7477), .A2(n7480), .A3(n7478), .ZN(n14070) );
  NAND2_X1 U9303 ( .A1(n9138), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9168) );
  NAND2_X1 U9304 ( .A1(n9184), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9218) );
  NAND3_X1 U9305 ( .A1(n9558), .A2(n9559), .A3(n7202), .ZN(n7325) );
  NOR2_X1 U9306 ( .A1(n14097), .A2(n7200), .ZN(n7326) );
  AND2_X1 U9307 ( .A1(n8896), .A2(n8920), .ZN(n10308) );
  NAND2_X1 U9308 ( .A1(n7347), .A2(n7346), .ZN(n13012) );
  INV_X1 U9309 ( .A(n12692), .ZN(n7836) );
  NAND3_X1 U9310 ( .A1(n7843), .A2(n7844), .A3(n13449), .ZN(n13181) );
  OAI22_X1 U9311 ( .A1(n8229), .A2(n8049), .B1(n7157), .B2(n11274), .ZN(n7525)
         );
  OAI21_X1 U9312 ( .B1(n8739), .B2(n16048), .A(n8738), .ZN(P3_U3456) );
  NAND2_X1 U9313 ( .A1(n10728), .A2(n7820), .ZN(n10912) );
  INV_X1 U9314 ( .A(n7797), .ZN(n14602) );
  NAND2_X1 U9315 ( .A1(n7789), .A2(n7787), .ZN(n14688) );
  OAI21_X4 U9316 ( .B1(n10471), .B2(n9395), .A(n9016), .ZN(n11938) );
  INV_X1 U9317 ( .A(n10784), .ZN(n10240) );
  NOR2_X1 U9318 ( .A1(n11315), .A2(n7349), .ZN(n7357) );
  NAND2_X1 U9319 ( .A1(n15775), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n15778) );
  INV_X1 U9320 ( .A(n12120), .ZN(n7585) );
  NOR2_X1 U9321 ( .A1(n11832), .A2(n7587), .ZN(n15817) );
  INV_X1 U9322 ( .A(n8989), .ZN(n7341) );
  OAI21_X4 U9323 ( .B1(n10433), .B2(n9395), .A(n8995), .ZN(n11742) );
  NAND2_X1 U9324 ( .A1(n8845), .A2(n8844), .ZN(n8866) );
  NAND2_X1 U9325 ( .A1(n10895), .A2(n10942), .ZN(n10944) );
  NAND2_X1 U9326 ( .A1(n15750), .A2(n15751), .ZN(n7340) );
  NAND2_X1 U9327 ( .A1(n8842), .A2(n8841), .ZN(n8845) );
  NAND2_X1 U9328 ( .A1(n10717), .A2(n10713), .ZN(n10712) );
  NAND2_X1 U9329 ( .A1(n8920), .A2(n8919), .ZN(n8938) );
  AOI21_X1 U9330 ( .B1(n7726), .B2(n7227), .A(n7725), .ZN(n7724) );
  OAI21_X2 U9331 ( .B1(n9365), .B2(n7736), .A(n7733), .ZN(n9564) );
  NAND2_X1 U9332 ( .A1(n9529), .A2(n9533), .ZN(n9567) );
  INV_X1 U9333 ( .A(n7720), .ZN(n7719) );
  NAND2_X1 U9334 ( .A1(n8092), .A2(n7203), .ZN(n8148) );
  NAND2_X1 U9335 ( .A1(n12472), .A2(n8637), .ZN(n8639) );
  NAND2_X1 U9336 ( .A1(n11336), .A2(n8623), .ZN(n11665) );
  NAND2_X1 U9337 ( .A1(n11904), .A2(n8627), .ZN(n11989) );
  NAND2_X1 U9338 ( .A1(n13421), .A2(n8655), .ZN(n13410) );
  NOR2_X2 U9339 ( .A1(n8148), .A2(P3_IR_REG_26__SCAN_IN), .ZN(n7717) );
  NAND2_X1 U9340 ( .A1(n7713), .A2(n7260), .ZN(n13421) );
  INV_X1 U9341 ( .A(n11326), .ZN(n11471) );
  INV_X1 U9342 ( .A(n13011), .ZN(n7347) );
  AOI21_X1 U9343 ( .B1(n10935), .B2(P3_REG2_REG_3__SCAN_IN), .A(n7348), .ZN(
        n10867) );
  AND2_X1 U9344 ( .A1(n10865), .A2(n10949), .ZN(n7348) );
  NAND2_X1 U9345 ( .A1(n15160), .A2(n16017), .ZN(n7664) );
  NAND3_X1 U9346 ( .A1(n7168), .A2(n11930), .A3(n11455), .ZN(n11868) );
  XNOR2_X1 U9347 ( .A(n7662), .B(n15379), .ZN(P1_U3527) );
  NAND2_X1 U9348 ( .A1(n10015), .A2(n10014), .ZN(n11041) );
  NAND2_X1 U9349 ( .A1(n11448), .A2(n11447), .ZN(n10019) );
  OAI21_X1 U9350 ( .B1(n10104), .B2(n7362), .A(n7351), .ZN(n10101) );
  OAI21_X1 U9351 ( .B1(n10104), .B2(n7917), .A(n7352), .ZN(n10107) );
  XNOR2_X1 U9352 ( .A(n13755), .B(n8101), .ZN(n13865) );
  INV_X1 U9353 ( .A(n11878), .ZN(n7976) );
  AND2_X2 U9354 ( .A1(n7966), .A2(n13836), .ZN(n7359) );
  XNOR2_X1 U9355 ( .A(n11312), .B(n11311), .ZN(n11431) );
  NAND2_X1 U9356 ( .A1(n11723), .A2(n11722), .ZN(n11915) );
  NAND2_X1 U9357 ( .A1(n7831), .A2(n7829), .ZN(n13039) );
  INV_X1 U9358 ( .A(n13009), .ZN(n7356) );
  XNOR2_X1 U9359 ( .A(n8689), .B(P3_B_REG_SCAN_IN), .ZN(n8683) );
  NAND2_X1 U9360 ( .A1(n7524), .A2(n7717), .ZN(n8685) );
  INV_X1 U9361 ( .A(n7981), .ZN(n7980) );
  NAND2_X1 U9362 ( .A1(n11743), .A2(n11744), .ZN(n11879) );
  NAND2_X1 U9363 ( .A1(n13221), .A2(n13222), .ZN(n13220) );
  NAND2_X1 U9364 ( .A1(n7931), .A2(n7930), .ZN(n14935) );
  INV_X2 U9365 ( .A(n16014), .ZN(n7362) );
  NAND2_X1 U9366 ( .A1(n7364), .A2(n7363), .ZN(P3_U3180) );
  NAND2_X1 U9367 ( .A1(n13214), .A2(n13223), .ZN(n7364) );
  NAND2_X1 U9368 ( .A1(n8043), .A2(n8049), .ZN(n8046) );
  NAND2_X1 U9369 ( .A1(n7974), .A2(n7977), .ZN(n7973) );
  XNOR2_X2 U9370 ( .A(n7365), .B(n10181), .ZN(n14061) );
  NAND2_X1 U9371 ( .A1(n7552), .A2(n10129), .ZN(n14226) );
  NAND2_X1 U9372 ( .A1(n7653), .A2(n7651), .ZN(n14177) );
  INV_X1 U9373 ( .A(n12371), .ZN(n7554) );
  OAI21_X1 U9374 ( .B1(n10216), .B2(n16034), .A(n8075), .ZN(P2_U3528) );
  OAI21_X1 U9375 ( .B1(n10216), .B2(n16001), .A(n10214), .ZN(P2_U3496) );
  OAI21_X2 U9376 ( .B1(n12344), .B2(n7988), .A(n7986), .ZN(n12449) );
  NAND2_X1 U9377 ( .A1(n7973), .A2(n12055), .ZN(n7972) );
  INV_X4 U9378 ( .A(n10276), .ZN(n9648) );
  INV_X1 U9379 ( .A(n7370), .ZN(n8389) );
  OAI211_X1 U9380 ( .C1(n7695), .C2(n7380), .A(n7376), .B(n12273), .ZN(n7383)
         );
  INV_X1 U9381 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7395) );
  INV_X1 U9382 ( .A(n7566), .ZN(n7396) );
  INV_X1 U9383 ( .A(n7700), .ZN(n7399) );
  NAND2_X1 U9384 ( .A1(n7687), .A2(n7408), .ZN(n7405) );
  NAND2_X1 U9385 ( .A1(n7405), .A2(n7406), .ZN(n8129) );
  AND2_X4 U9386 ( .A1(n9725), .A2(n9594), .ZN(n9826) );
  AND4_X2 U9387 ( .A1(n7417), .A2(n9588), .A3(n9626), .A4(n7416), .ZN(n9725)
         );
  OAI21_X1 U9388 ( .B1(n7173), .B2(n7424), .A(n7422), .ZN(n7870) );
  INV_X4 U9389 ( .A(n12728), .ZN(n12873) );
  NAND2_X2 U9390 ( .A1(n12858), .A2(n7428), .ZN(n12728) );
  AOI21_X1 U9391 ( .B1(n10001), .B2(n7253), .A(n7432), .ZN(n7431) );
  OAI22_X1 U9392 ( .A1(n7171), .A2(n7437), .B1(n12815), .B2(n7440), .ZN(n12817) );
  INV_X1 U9393 ( .A(n12814), .ZN(n7440) );
  OAI22_X1 U9394 ( .A1(n7441), .A2(n7236), .B1(n7443), .B2(n12831), .ZN(n12834) );
  NAND2_X1 U9395 ( .A1(n12829), .A2(n7442), .ZN(n7441) );
  INV_X1 U9396 ( .A(n12830), .ZN(n7443) );
  NAND2_X1 U9397 ( .A1(n12658), .A2(n7444), .ZN(n11332) );
  OAI21_X1 U9398 ( .B1(n12658), .B2(n7444), .A(n11332), .ZN(n11843) );
  OR2_X1 U9399 ( .A1(n9573), .A2(n7454), .ZN(n7451) );
  NAND2_X1 U9400 ( .A1(n7451), .A2(n7452), .ZN(n12690) );
  INV_X1 U9401 ( .A(n12690), .ZN(n12515) );
  NAND2_X1 U9402 ( .A1(n11850), .A2(n7457), .ZN(n7455) );
  NAND2_X1 U9403 ( .A1(n7455), .A2(n7263), .ZN(n11986) );
  INV_X1 U9404 ( .A(n13486), .ZN(n7460) );
  OAI21_X1 U9405 ( .B1(n7460), .B2(n7464), .A(n7461), .ZN(n13458) );
  AND2_X1 U9406 ( .A1(n8210), .A2(n8139), .ZN(n8141) );
  NAND2_X1 U9407 ( .A1(n8352), .A2(n7471), .ZN(n7469) );
  OAI21_X1 U9408 ( .B1(n8352), .B2(n7473), .A(n7471), .ZN(n8411) );
  NAND3_X1 U9409 ( .A1(n7892), .A2(n7475), .A3(n7715), .ZN(n13715) );
  NAND2_X1 U9410 ( .A1(n10966), .A2(n10146), .ZN(n10148) );
  NAND2_X1 U9411 ( .A1(n10757), .A2(n10756), .ZN(n7476) );
  NAND2_X1 U9412 ( .A1(n7225), .A2(n14111), .ZN(n7477) );
  INV_X1 U9413 ( .A(n7493), .ZN(n8023) );
  AOI21_X1 U9414 ( .B1(n8758), .B2(P2_IR_REG_29__SCAN_IN), .A(n7502), .ZN(
        n7501) );
  NAND2_X1 U9415 ( .A1(n9010), .A2(n7511), .ZN(n7510) );
  NAND2_X1 U9416 ( .A1(n13846), .A2(n13845), .ZN(n13844) );
  NAND2_X1 U9417 ( .A1(n13846), .A2(n7249), .ZN(n7516) );
  INV_X1 U9418 ( .A(n9204), .ZN(n9205) );
  INV_X1 U9419 ( .A(n8141), .ZN(n8249) );
  INV_X2 U9420 ( .A(n8471), .ZN(n7892) );
  NAND4_X1 U9421 ( .A1(n7542), .A2(n12633), .A3(n13435), .A4(n7541), .ZN(n7540) );
  NAND3_X1 U9422 ( .A1(n12630), .A2(n12629), .A3(n12675), .ZN(n7542) );
  NAND2_X1 U9423 ( .A1(n10112), .A2(n10752), .ZN(n10114) );
  NAND2_X2 U9424 ( .A1(n7544), .A2(n14405), .ZN(n8794) );
  NAND2_X2 U9425 ( .A1(n8785), .A2(n7544), .ZN(n8856) );
  NAND2_X1 U9426 ( .A1(n11587), .A2(n7548), .ZN(n7547) );
  NAND2_X1 U9427 ( .A1(n7547), .A2(n7545), .ZN(n11729) );
  OR2_X1 U9428 ( .A1(n7550), .A2(n10119), .ZN(n7546) );
  NAND2_X1 U9429 ( .A1(n11340), .A2(n10117), .ZN(n11403) );
  XNOR2_X2 U9430 ( .A(n13932), .B(n11503), .ZN(n10717) );
  AOI21_X2 U9431 ( .B1(n14087), .B2(n14086), .A(n7644), .ZN(n14079) );
  NAND2_X2 U9432 ( .A1(n14316), .A2(n7645), .ZN(n14087) );
  OR2_X2 U9433 ( .A1(n14108), .A2(n7483), .ZN(n14316) );
  NAND2_X1 U9434 ( .A1(n7558), .A2(n8763), .ZN(n12959) );
  NAND2_X1 U9435 ( .A1(n8763), .A2(n8004), .ZN(n8761) );
  NAND2_X1 U9436 ( .A1(n11022), .A2(n7574), .ZN(n7576) );
  NAND2_X1 U9437 ( .A1(n13273), .A2(n7579), .ZN(n13256) );
  INV_X1 U9438 ( .A(n12169), .ZN(n7581) );
  OR2_X1 U9439 ( .A1(n7582), .A2(n12169), .ZN(n12122) );
  INV_X1 U9440 ( .A(n7584), .ZN(n7582) );
  INV_X1 U9441 ( .A(n7589), .ZN(n14178) );
  NAND2_X1 U9442 ( .A1(n7590), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8756) );
  AND2_X2 U9443 ( .A1(n12378), .A2(n14403), .ZN(n14281) );
  NOR2_X2 U9444 ( .A1(n14089), .A2(n14305), .ZN(n7595) );
  NOR2_X2 U9445 ( .A1(n11213), .A2(n11218), .ZN(n11344) );
  NAND2_X1 U9446 ( .A1(n7621), .A2(n7622), .ZN(n13395) );
  NAND2_X1 U9447 ( .A1(n12243), .A2(n7637), .ZN(n8352) );
  NAND2_X1 U9448 ( .A1(n10121), .A2(n7648), .ZN(n7647) );
  NAND2_X1 U9449 ( .A1(n7647), .A2(n7646), .ZN(n10123) );
  AOI21_X1 U9450 ( .B1(n7648), .B2(n7650), .A(n10160), .ZN(n7646) );
  NAND2_X2 U9451 ( .A1(n10443), .A2(n14411), .ZN(n8802) );
  XNOR2_X2 U9452 ( .A(n8762), .B(n7592), .ZN(n14411) );
  NOR2_X2 U9453 ( .A1(n8761), .A2(n8013), .ZN(n8758) );
  AND2_X1 U9454 ( .A1(n14247), .A2(n10128), .ZN(n7656) );
  NAND2_X1 U9455 ( .A1(n14953), .A2(n7667), .ZN(n14892) );
  NAND2_X1 U9456 ( .A1(n11867), .A2(n7672), .ZN(n15035) );
  NAND2_X1 U9457 ( .A1(n8413), .A2(n7689), .ZN(n7687) );
  NAND2_X1 U9458 ( .A1(n7702), .A2(n11015), .ZN(n8618) );
  XNOR2_X1 U9459 ( .A(n12657), .B(n7703), .ZN(n11018) );
  INV_X1 U9460 ( .A(n11015), .ZN(n7703) );
  XNOR2_X1 U9461 ( .A(n11313), .B(n12657), .ZN(n11020) );
  NAND2_X1 U9462 ( .A1(n13490), .A2(n7169), .ZN(n7704) );
  NAND2_X1 U9463 ( .A1(n11663), .A2(n7709), .ZN(n11852) );
  NAND2_X1 U9464 ( .A1(n8639), .A2(n7284), .ZN(n13547) );
  NAND2_X1 U9465 ( .A1(n13547), .A2(n8641), .ZN(n8643) );
  NAND2_X1 U9466 ( .A1(n8658), .A2(n8657), .ZN(n13399) );
  NAND2_X2 U9467 ( .A1(n8324), .A2(n8096), .ZN(n8471) );
  OAI21_X1 U9468 ( .B1(n8676), .B2(n13578), .A(n8675), .ZN(n13380) );
  NAND2_X1 U9469 ( .A1(n7738), .A2(n7741), .ZN(n9243) );
  NAND3_X1 U9470 ( .A1(n9198), .A2(n7739), .A3(n9197), .ZN(n7738) );
  NAND2_X1 U9471 ( .A1(n7742), .A2(n7740), .ZN(n7739) );
  NAND2_X1 U9472 ( .A1(n9226), .A2(n9225), .ZN(n7741) );
  NAND2_X1 U9473 ( .A1(n9268), .A2(n7746), .ZN(n7743) );
  NAND2_X1 U9474 ( .A1(n7743), .A2(n7744), .ZN(n9299) );
  INV_X1 U9475 ( .A(n9283), .ZN(n7755) );
  INV_X1 U9476 ( .A(n9267), .ZN(n7757) );
  OAI21_X1 U9477 ( .B1(n9175), .B2(n7762), .A(n7761), .ZN(n9195) );
  NAND2_X1 U9478 ( .A1(n7758), .A2(n7759), .ZN(n9194) );
  NAND2_X1 U9479 ( .A1(n9175), .A2(n7761), .ZN(n7758) );
  INV_X1 U9480 ( .A(n9174), .ZN(n7764) );
  NAND3_X1 U9481 ( .A1(n9110), .A2(n7268), .A3(n9109), .ZN(n7769) );
  NAND2_X1 U9482 ( .A1(n7769), .A2(n7770), .ZN(n9152) );
  AOI21_X1 U9483 ( .B1(n9152), .B2(n9151), .A(n9149), .ZN(n9150) );
  NAND2_X1 U9484 ( .A1(n7773), .A2(n7774), .ZN(n8884) );
  NAND3_X1 U9485 ( .A1(n8840), .A2(n8839), .A3(n7267), .ZN(n7773) );
  NAND3_X1 U9486 ( .A1(n10625), .A2(n10644), .A3(n10626), .ZN(n10645) );
  NAND2_X1 U9487 ( .A1(n10645), .A2(n7775), .ZN(n10627) );
  NAND2_X1 U9488 ( .A1(n7776), .A2(n7777), .ZN(n7775) );
  INV_X1 U9489 ( .A(n10626), .ZN(n7776) );
  NAND2_X1 U9490 ( .A1(n7778), .A2(n7779), .ZN(n12389) );
  NAND2_X4 U9491 ( .A1(n14492), .A2(n15036), .ZN(n14588) );
  NAND2_X1 U9492 ( .A1(n14492), .A2(n7784), .ZN(n7786) );
  INV_X1 U9493 ( .A(n15036), .ZN(n7785) );
  NAND2_X1 U9494 ( .A1(n14663), .A2(n7790), .ZN(n7789) );
  AND2_X1 U9495 ( .A1(n14490), .A2(n14491), .ZN(n7806) );
  OR2_X1 U9496 ( .A1(n14477), .A2(n14478), .ZN(n7807) );
  NAND2_X1 U9497 ( .A1(n12030), .A2(n12029), .ZN(n12150) );
  XNOR2_X1 U9498 ( .A(n12150), .B(n12151), .ZN(n12037) );
  NAND3_X1 U9499 ( .A1(n10730), .A2(n10727), .A3(n7817), .ZN(n7816) );
  INV_X1 U9500 ( .A(n10647), .ZN(n7817) );
  NAND2_X1 U9501 ( .A1(n10646), .A2(n10647), .ZN(n10728) );
  NAND2_X1 U9502 ( .A1(n11295), .A2(n7823), .ZN(n7822) );
  NAND2_X1 U9503 ( .A1(n9985), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9638) );
  INV_X1 U9504 ( .A(n12707), .ZN(n11152) );
  OAI21_X1 U9505 ( .B1(n13111), .B2(n7834), .A(n7832), .ZN(n13038) );
  NAND2_X1 U9506 ( .A1(n13111), .A2(n7832), .ZN(n7831) );
  NAND2_X1 U9507 ( .A1(n13111), .A2(n13020), .ZN(n13211) );
  OR2_X2 U9508 ( .A1(n8692), .A2(P3_D_REG_0__SCAN_IN), .ZN(n7838) );
  NAND2_X1 U9509 ( .A1(n7840), .A2(n7839), .ZN(n13106) );
  AOI21_X1 U9510 ( .B1(n13144), .B2(n13239), .A(n7841), .ZN(n7839) );
  NAND2_X1 U9511 ( .A1(n13068), .A2(n13144), .ZN(n7840) );
  INV_X1 U9512 ( .A(n13069), .ZN(n7842) );
  NAND2_X1 U9513 ( .A1(n13009), .A2(n13008), .ZN(n7844) );
  NAND2_X1 U9514 ( .A1(n7843), .A2(n7844), .ZN(n13180) );
  NAND2_X1 U9515 ( .A1(n13181), .A2(n7844), .ZN(n13011) );
  NAND2_X1 U9516 ( .A1(n12228), .A2(n7264), .ZN(n12426) );
  NAND2_X1 U9517 ( .A1(n7845), .A2(n7848), .ZN(n12844) );
  NAND3_X1 U9518 ( .A1(n12839), .A2(n7846), .A3(n12838), .ZN(n7845) );
  OR2_X1 U9519 ( .A1(n12748), .A2(n12747), .ZN(n7852) );
  NAND2_X1 U9520 ( .A1(n13163), .A2(n7853), .ZN(n13007) );
  NAND2_X1 U9521 ( .A1(n7854), .A2(n7857), .ZN(n12746) );
  NAND3_X1 U9522 ( .A1(n12737), .A2(n7855), .A3(n12736), .ZN(n7854) );
  NAND2_X1 U9523 ( .A1(n7858), .A2(n7859), .ZN(n12767) );
  NAND3_X1 U9524 ( .A1(n12758), .A2(n12759), .A3(n7261), .ZN(n7858) );
  NAND2_X1 U9525 ( .A1(n12817), .A2(n7863), .ZN(n7860) );
  NAND2_X1 U9526 ( .A1(n7860), .A2(n7861), .ZN(n12825) );
  NAND2_X1 U9527 ( .A1(n7870), .A2(n7871), .ZN(n12806) );
  NAND3_X1 U9528 ( .A1(n12772), .A2(n12771), .A3(n7262), .ZN(n7872) );
  NAND2_X1 U9529 ( .A1(n7872), .A2(n7873), .ZN(n12780) );
  INV_X1 U9530 ( .A(n13120), .ZN(n7883) );
  NAND2_X1 U9531 ( .A1(n13120), .A2(n7879), .ZN(n7874) );
  NOR2_X1 U9532 ( .A1(n7272), .A2(n12990), .ZN(n13138) );
  NAND2_X1 U9533 ( .A1(n7885), .A2(n7886), .ZN(n12790) );
  NAND3_X1 U9534 ( .A1(n12785), .A2(n12784), .A3(n7256), .ZN(n7885) );
  NAND3_X1 U9535 ( .A1(n9826), .A2(n7889), .A3(n9602), .ZN(n15421) );
  NAND2_X1 U9536 ( .A1(n9826), .A2(n9602), .ZN(n9607) );
  NOR2_X2 U9537 ( .A1(n8471), .A2(n7890), .ZN(n8603) );
  NAND3_X1 U9538 ( .A1(n7896), .A2(n7897), .A3(n7209), .ZN(n9685) );
  NAND3_X1 U9539 ( .A1(n7900), .A2(n7899), .A3(n9670), .ZN(n7897) );
  INV_X1 U9540 ( .A(n15873), .ZN(n7899) );
  INV_X1 U9541 ( .A(n15870), .ZN(n7900) );
  OR2_X1 U9542 ( .A1(n15870), .A2(n15873), .ZN(n7901) );
  NAND2_X1 U9543 ( .A1(n11865), .A2(n7910), .ZN(n7909) );
  NAND2_X1 U9544 ( .A1(n7909), .A2(n7912), .ZN(n15043) );
  OAI21_X1 U9545 ( .B1(n11509), .B2(n7928), .A(n7926), .ZN(n9781) );
  NAND2_X1 U9546 ( .A1(n9905), .A2(n7933), .ZN(n7931) );
  INV_X1 U9547 ( .A(n9917), .ZN(n7935) );
  XNOR2_X2 U9548 ( .A(n7936), .B(n9609), .ZN(n12957) );
  XNOR2_X2 U9549 ( .A(n7937), .B(n9608), .ZN(n9610) );
  AOI21_X1 U9550 ( .B1(n7941), .B2(n12879), .A(n7248), .ZN(n7938) );
  NAND2_X1 U9551 ( .A1(n10686), .A2(n7940), .ZN(n7939) );
  NAND2_X1 U9552 ( .A1(n7943), .A2(n7944), .ZN(n11863) );
  NAND2_X1 U9553 ( .A1(n11510), .A2(n7246), .ZN(n7943) );
  OAI21_X2 U9554 ( .B1(n15046), .B2(n7948), .A(n7947), .ZN(n15010) );
  OAI21_X2 U9555 ( .B1(n14916), .B2(n7192), .A(n7953), .ZN(n14891) );
  OAI21_X1 U9556 ( .B1(n14877), .B2(n7959), .A(n7957), .ZN(n10046) );
  NAND2_X1 U9557 ( .A1(n14877), .A2(n14885), .ZN(n14876) );
  NAND2_X2 U9558 ( .A1(n15432), .A2(n15429), .ZN(n10323) );
  OAI211_X2 U9559 ( .C1(n7980), .C2(n10823), .A(n11065), .B(n7979), .ZN(n11380) );
  AND2_X2 U9560 ( .A1(n13825), .A2(n7994), .ZN(n13895) );
  NAND2_X1 U9561 ( .A1(n12101), .A2(n7996), .ZN(n12343) );
  INV_X1 U9562 ( .A(n11382), .ZN(n8003) );
  NAND3_X1 U9563 ( .A1(n13877), .A2(n10245), .A3(n10255), .ZN(n10783) );
  NAND4_X1 U9564 ( .A1(n8754), .A2(n8755), .A3(n8752), .A4(n8753), .ZN(n8005)
         );
  NAND2_X1 U9565 ( .A1(n8016), .A2(n8014), .ZN(n8020) );
  NAND2_X1 U9566 ( .A1(n8023), .A2(n8021), .ZN(n10156) );
  INV_X1 U9567 ( .A(n11402), .ZN(n8025) );
  NAND2_X1 U9568 ( .A1(n14141), .A2(n8031), .ZN(n8026) );
  NAND2_X1 U9569 ( .A1(n8026), .A2(n8027), .ZN(n14111) );
  INV_X1 U9570 ( .A(n8805), .ZN(n8043) );
  OAI211_X1 U9571 ( .C1(n8806), .C2(P2_DATAO_REG_0__SCAN_IN), .A(n8048), .B(
        SI_0_), .ZN(n8047) );
  NAND2_X1 U9572 ( .A1(n8806), .A2(n8807), .ZN(n8048) );
  INV_X1 U9573 ( .A(SI_1_), .ZN(n8049) );
  NAND2_X1 U9574 ( .A1(n8964), .A2(n8963), .ZN(n8985) );
  NAND2_X1 U9575 ( .A1(n8964), .A2(n8062), .ZN(n8061) );
  NAND2_X1 U9576 ( .A1(n8895), .A2(n8067), .ZN(n8066) );
  NAND2_X1 U9577 ( .A1(n8895), .A2(n8894), .ZN(n8920) );
  NAND2_X1 U9578 ( .A1(n8066), .A2(n8068), .ZN(n8943) );
  NAND2_X1 U9579 ( .A1(n9159), .A2(n8086), .ZN(n8081) );
  NAND2_X1 U9580 ( .A1(n9159), .A2(n9158), .ZN(n9178) );
  OR2_X1 U9581 ( .A1(n14069), .A2(n8856), .ZN(n9436) );
  INV_X1 U9582 ( .A(n8856), .ZN(n9452) );
  OR2_X1 U9583 ( .A1(n9573), .A2(n7543), .ZN(n9575) );
  NAND2_X1 U9584 ( .A1(n10062), .A2(n10061), .ZN(n10064) );
  INV_X1 U9585 ( .A(n10060), .ZN(n10062) );
  INV_X1 U9586 ( .A(n11333), .ZN(n8622) );
  INV_X1 U9587 ( .A(n9985), .ZN(n9620) );
  NOR2_X1 U9588 ( .A1(n9564), .A2(n9532), .ZN(n9566) );
  INV_X1 U9590 ( .A(n9053), .ZN(n9056) );
  NAND2_X1 U9591 ( .A1(n9153), .A2(n7208), .ZN(n9175) );
  CLKBUF_X1 U9592 ( .A(n11743), .Z(n11745) );
  INV_X1 U9593 ( .A(n9826), .ZN(n9827) );
  INV_X1 U9594 ( .A(n11151), .ZN(n9660) );
  INV_X1 U9595 ( .A(n9998), .ZN(n9838) );
  OAI21_X1 U9596 ( .B1(n8838), .B2(n8837), .A(n8836), .ZN(n8840) );
  AND2_X1 U9597 ( .A1(n8872), .A2(n8891), .ZN(n10296) );
  NAND2_X4 U9598 ( .A1(n12702), .A2(n12706), .ZN(n14586) );
  INV_X1 U9599 ( .A(n14588), .ZN(n14537) );
  AND2_X1 U9600 ( .A1(n10439), .A2(n10443), .ZN(n14275) );
  OR2_X1 U9601 ( .A1(n9581), .A2(n10297), .ZN(n9582) );
  INV_X1 U9602 ( .A(n9610), .ZN(n9612) );
  NAND2_X1 U9603 ( .A1(n8643), .A2(n8642), .ZN(n13533) );
  MUX2_X1 U9604 ( .A(P2_IR_REG_0__SCAN_IN), .B(n14424), .S(n8802), .Z(n11250)
         );
  NAND2_X1 U9605 ( .A1(n10059), .A2(n10058), .ZN(n10104) );
  XNOR2_X1 U9606 ( .A(n10240), .B(n10721), .ZN(n10238) );
  NAND2_X2 U9607 ( .A1(n9610), .A2(n9611), .ZN(n9665) );
  NAND2_X2 U9608 ( .A1(n8186), .A2(n8187), .ZN(n8224) );
  OR2_X1 U9609 ( .A1(n14134), .A2(n13915), .ZN(n8088) );
  XOR2_X1 U9610 ( .A(n14149), .B(n13764), .Z(n8089) );
  INV_X1 U9611 ( .A(n16001), .ZN(n14371) );
  AND2_X1 U9612 ( .A1(n10215), .A2(n15454), .ZN(n14398) );
  INV_X1 U9613 ( .A(n14398), .ZN(n16001) );
  NAND2_X2 U9614 ( .A1(n11247), .A2(n14255), .ZN(n14280) );
  AND2_X1 U9615 ( .A1(n10185), .A2(n10184), .ZN(n14243) );
  OR2_X1 U9616 ( .A1(n13514), .A2(n13492), .ZN(n8090) );
  NOR2_X1 U9617 ( .A1(n13383), .A2(n13707), .ZN(n8091) );
  INV_X1 U9618 ( .A(n16042), .ZN(n16048) );
  INV_X1 U9619 ( .A(n16039), .ZN(n8727) );
  INV_X1 U9620 ( .A(n12664), .ZN(n8629) );
  AND2_X1 U9621 ( .A1(n8147), .A2(n8681), .ZN(n8092) );
  AND4_X1 U9622 ( .A1(n9997), .A2(n9996), .A3(n9868), .A4(n9995), .ZN(n8093)
         );
  INV_X1 U9623 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14415) );
  AND2_X1 U9624 ( .A1(n13772), .A2(n13771), .ZN(n8094) );
  INV_X1 U9625 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n15420) );
  NOR2_X1 U9626 ( .A1(n13558), .A2(n13548), .ZN(n8097) );
  INV_X1 U9627 ( .A(n14250), .ZN(n14209) );
  INV_X1 U9628 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n8804) );
  INV_X1 U9629 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8155) );
  NAND2_X1 U9630 ( .A1(n10834), .A2(n9563), .ZN(n8098) );
  INV_X1 U9631 ( .A(n13567), .ZN(n8437) );
  AND2_X1 U9632 ( .A1(n12937), .A2(n12936), .ZN(n8099) );
  OR2_X1 U9633 ( .A1(n12934), .A2(n12951), .ZN(n8100) );
  XOR2_X1 U9634 ( .A(n14162), .B(n13805), .Z(n8101) );
  NAND3_X1 U9635 ( .A1(n14834), .A2(n14836), .A3(n14838), .ZN(n8102) );
  INV_X1 U9636 ( .A(n14599), .ZN(n14849) );
  OAI22_X1 U9637 ( .A1(n9425), .A2(n9424), .B1(SI_28_), .B2(n9376), .ZN(n9410)
         );
  INV_X1 U9638 ( .A(n8816), .ZN(n9419) );
  NAND2_X1 U9639 ( .A1(n16017), .A2(n15982), .ZN(n15402) );
  INV_X1 U9640 ( .A(n15402), .ZN(n10105) );
  INV_X1 U9641 ( .A(n15125), .ZN(n10229) );
  AND2_X1 U9642 ( .A1(n12760), .A2(n10020), .ZN(n8103) );
  OR2_X1 U9643 ( .A1(n12760), .A2(n10020), .ZN(n8104) );
  INV_X1 U9644 ( .A(n12751), .ZN(n12752) );
  NOR2_X1 U9645 ( .A1(n8792), .A2(n8791), .ZN(n8815) );
  AOI22_X1 U9646 ( .A1(n13932), .A2(n8883), .B1(n10721), .B2(n9484), .ZN(n8820) );
  OAI22_X1 U9647 ( .A1(n11524), .A2(n9489), .B1(n10785), .B2(n9315), .ZN(n8885) );
  OAI22_X1 U9648 ( .A1(n11524), .A2(n9315), .B1(n10785), .B2(n9362), .ZN(n8888) );
  AND2_X1 U9649 ( .A1(n8915), .A2(n8914), .ZN(n8916) );
  OAI22_X1 U9650 ( .A1(n15965), .A2(n9482), .B1(n11948), .B2(n9489), .ZN(n9054) );
  INV_X1 U9651 ( .A(n9054), .ZN(n9055) );
  OAI22_X1 U9652 ( .A1(n12203), .A2(n9362), .B1(n12144), .B2(n9315), .ZN(n9076) );
  OAI22_X1 U9653 ( .A1(n16030), .A2(n9362), .B1(n14236), .B2(n9315), .ZN(n9193) );
  NAND2_X1 U9654 ( .A1(n9246), .A2(n9245), .ZN(n9247) );
  INV_X1 U9655 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8744) );
  INV_X1 U9656 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8147) );
  INV_X1 U9657 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8747) );
  INV_X1 U9658 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9995) );
  OR2_X1 U9659 ( .A1(n12979), .A2(n12978), .ZN(n12980) );
  INV_X1 U9660 ( .A(n13398), .ZN(n8659) );
  INV_X1 U9661 ( .A(n12674), .ZN(n13489) );
  INV_X1 U9662 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n12179) );
  INV_X1 U9663 ( .A(n12661), .ZN(n8626) );
  INV_X1 U9664 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8134) );
  INV_X1 U9665 ( .A(n9186), .ZN(n9184) );
  NAND2_X1 U9666 ( .A1(n13751), .A2(n13753), .ZN(n13754) );
  INV_X1 U9667 ( .A(n11242), .ZN(n10235) );
  INV_X1 U9668 ( .A(n9275), .ZN(n9274) );
  INV_X1 U9669 ( .A(n10180), .ZN(n10181) );
  INV_X1 U9670 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8748) );
  INV_X1 U9671 ( .A(n14585), .ZN(n14532) );
  NOR2_X1 U9672 ( .A1(n9832), .A2(n14705), .ZN(n9831) );
  INV_X1 U9673 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9717) );
  INV_X1 U9674 ( .A(n15013), .ZN(n9865) );
  INV_X1 U9675 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9732) );
  INV_X1 U9676 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n15360) );
  INV_X1 U9677 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9589) );
  INV_X1 U9678 ( .A(n12232), .ZN(n12229) );
  OR2_X1 U9679 ( .A1(n8722), .A2(n13031), .ZN(n12637) );
  OR2_X1 U9680 ( .A1(n8693), .A2(n8706), .ZN(n8731) );
  INV_X1 U9681 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n8119) );
  NAND2_X1 U9682 ( .A1(n9338), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n9355) );
  AND2_X1 U9683 ( .A1(n14119), .A2(n13898), .ZN(n10176) );
  NOR2_X1 U9684 ( .A1(n10617), .A2(n14586), .ZN(n10616) );
  AND2_X1 U9685 ( .A1(n9831), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9843) );
  NAND2_X1 U9686 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(n9923), .ZN(n9932) );
  NOR2_X1 U9687 ( .A1(n9896), .A2(n14658), .ZN(n9909) );
  NAND2_X1 U9688 ( .A1(n9843), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9872) );
  OR2_X1 U9689 ( .A1(n15043), .A2(n15045), .ZN(n9837) );
  OR2_X1 U9690 ( .A1(n9775), .A2(n10596), .ZN(n9789) );
  INV_X1 U9691 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n15253) );
  AOI21_X1 U9692 ( .B1(n14845), .B2(n16013), .A(n8102), .ZN(n10058) );
  INV_X1 U9693 ( .A(n12860), .ZN(n12853) );
  AND2_X1 U9694 ( .A1(n10088), .A2(n10353), .ZN(n14702) );
  INV_X1 U9695 ( .A(n14607), .ZN(n14704) );
  NAND2_X1 U9696 ( .A1(n9346), .A2(n9345), .ZN(n9349) );
  INV_X1 U9697 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9598) );
  OR2_X1 U9698 ( .A1(n9782), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n9783) );
  INV_X1 U9699 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9671) );
  XNOR2_X1 U9700 ( .A(n11315), .B(n11316), .ZN(n11323) );
  NAND2_X1 U9701 ( .A1(n8179), .A2(n15267), .ZN(n8578) );
  OR2_X1 U9702 ( .A1(n8551), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8565) );
  NAND2_X1 U9703 ( .A1(n8176), .A2(n15261), .ZN(n8515) );
  NAND2_X1 U9704 ( .A1(n8175), .A2(n15253), .ZN(n8493) );
  NAND2_X1 U9705 ( .A1(n11318), .A2(n15846), .ZN(n13217) );
  OR2_X1 U9706 ( .A1(n8240), .A2(n8201), .ZN(n8207) );
  INV_X1 U9707 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15691) );
  INV_X1 U9708 ( .A(n13492), .ZN(n13525) );
  AND2_X1 U9709 ( .A1(n12609), .A2(n12612), .ZN(n13538) );
  AND2_X1 U9710 ( .A1(n13547), .A2(n13546), .ZN(n13563) );
  AND2_X1 U9711 ( .A1(n8731), .A2(n11109), .ZN(n8710) );
  OAI21_X1 U9712 ( .B1(n13395), .B2(n13398), .A(n13394), .ZN(n13599) );
  INV_X1 U9713 ( .A(n12697), .ZN(n8714) );
  INV_X1 U9714 ( .A(n8601), .ZN(n8606) );
  NAND2_X1 U9715 ( .A1(n13758), .A2(n8089), .ZN(n13759) );
  NAND2_X1 U9716 ( .A1(n13878), .A2(n13879), .ZN(n13877) );
  AND2_X1 U9717 ( .A1(n9451), .A2(n9450), .ZN(n14090) );
  AND2_X1 U9718 ( .A1(n8858), .A2(n8857), .ZN(n8859) );
  AND2_X1 U9719 ( .A1(n15505), .A2(n11133), .ZN(n14025) );
  INV_X1 U9720 ( .A(n10190), .ZN(n10191) );
  OR2_X1 U9721 ( .A1(n10265), .A2(n15452), .ZN(n14255) );
  INV_X1 U9722 ( .A(n14258), .ZN(n14288) );
  OR2_X1 U9723 ( .A1(n14371), .A2(n10211), .ZN(n10212) );
  INV_X1 U9724 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n14681) );
  AND2_X1 U9725 ( .A1(n10732), .A2(n15440), .ZN(n14701) );
  NAND2_X1 U9726 ( .A1(n12952), .A2(n12946), .ZN(n12947) );
  AND2_X1 U9727 ( .A1(n9909), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9911) );
  OR2_X1 U9728 ( .A1(n9886), .A2(n9885), .ZN(n9896) );
  INV_X1 U9729 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n15589) );
  INV_X1 U9730 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n15637) );
  OR2_X1 U9731 ( .A1(n10417), .A2(n10418), .ZN(n10415) );
  OR2_X1 U9732 ( .A1(n11004), .A2(n11003), .ZN(n11626) );
  INV_X1 U9733 ( .A(n12897), .ZN(n14911) );
  OR2_X1 U9734 ( .A1(n10799), .A2(n10000), .ZN(n15874) );
  INV_X1 U9735 ( .A(n15878), .ZN(n15985) );
  OR2_X1 U9736 ( .A1(n9741), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n9768) );
  OAI22_X1 U9737 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n15604), .B1(n15603), .B2(
        n15602), .ZN(n15611) );
  NAND2_X1 U9738 ( .A1(n11100), .A2(n11099), .ZN(n13230) );
  OR2_X1 U9739 ( .A1(n13371), .A2(n8224), .ZN(n12506) );
  INV_X1 U9740 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n15585) );
  INV_X1 U9741 ( .A(n13362), .ZN(n15808) );
  INV_X1 U9742 ( .A(n15800), .ZN(n15819) );
  INV_X1 U9743 ( .A(n13582), .ZN(n15848) );
  NAND2_X1 U9744 ( .A1(n11189), .A2(n11188), .ZN(n11408) );
  NAND2_X1 U9745 ( .A1(n8714), .A2(n11367), .ZN(n15970) );
  NOR3_X1 U9746 ( .A1(n12459), .A2(n14417), .A3(n12480), .ZN(n10233) );
  NAND2_X1 U9747 ( .A1(n11380), .A2(n11379), .ZN(n11382) );
  INV_X1 U9748 ( .A(n14195), .ZN(n14346) );
  INV_X1 U9749 ( .A(n13900), .ZN(n13872) );
  NAND2_X1 U9750 ( .A1(n9564), .A2(n9524), .ZN(n9529) );
  AND2_X1 U9751 ( .A1(n9314), .A2(n9313), .ZN(n13868) );
  OR2_X1 U9752 ( .A1(n15504), .A2(n15503), .ZN(n15505) );
  INV_X1 U9753 ( .A(n15502), .ZN(n15523) );
  AND2_X1 U9754 ( .A1(n15460), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15521) );
  AND2_X1 U9755 ( .A1(n10439), .A2(n10444), .ZN(n14274) );
  INV_X1 U9756 ( .A(n14243), .ZN(n14271) );
  AND2_X1 U9757 ( .A1(n11248), .A2(n14076), .ZN(n14290) );
  AND2_X1 U9758 ( .A1(n14280), .A2(n11370), .ZN(n14263) );
  NAND2_X1 U9759 ( .A1(n14279), .A2(n10138), .ZN(n16033) );
  OR2_X1 U9760 ( .A1(n14417), .A2(n10202), .ZN(n10209) );
  INV_X1 U9761 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n9538) );
  INV_X4 U9762 ( .A(n10276), .ZN(n10297) );
  INV_X1 U9763 ( .A(n12358), .ZN(n14419) );
  AND2_X1 U9764 ( .A1(n9898), .A2(n9897), .ZN(n14968) );
  INV_X1 U9765 ( .A(n14706), .ZN(n14671) );
  NAND2_X1 U9766 ( .A1(n10579), .A2(n15051), .ZN(n14709) );
  AND2_X1 U9767 ( .A1(n9618), .A2(n9617), .ZN(n14608) );
  AND2_X1 U9768 ( .A1(n10330), .A2(n15432), .ZN(n15566) );
  AND2_X1 U9769 ( .A1(n14963), .A2(n14962), .ZN(n15122) );
  AND2_X1 U9770 ( .A1(n15054), .A2(n16013), .ZN(n15000) );
  INV_X1 U9771 ( .A(n15061), .ZN(n15022) );
  NAND2_X1 U9772 ( .A1(n10098), .A2(n10811), .ZN(n15982) );
  NAND2_X1 U9773 ( .A1(n10050), .A2(n10049), .ZN(n16013) );
  NAND2_X1 U9774 ( .A1(n15874), .A2(n15884), .ZN(n15992) );
  INV_X1 U9775 ( .A(n15884), .ZN(n15926) );
  AND2_X1 U9776 ( .A1(n10872), .A2(n10871), .ZN(n15806) );
  INV_X1 U9777 ( .A(n13223), .ZN(n13196) );
  INV_X1 U9778 ( .A(n13230), .ZN(n13175) );
  AND2_X1 U9779 ( .A1(n12506), .A2(n8191), .ZN(n13031) );
  OR2_X1 U9780 ( .A1(n10869), .A2(n10868), .ZN(n15742) );
  INV_X1 U9781 ( .A(n15814), .ZN(n15763) );
  INV_X1 U9782 ( .A(n13500), .ZN(n12292) );
  AND2_X2 U9783 ( .A1(n11189), .A2(n8721), .ZN(n16039) );
  NOR2_X1 U9784 ( .A1(n8091), .A2(n8737), .ZN(n8738) );
  INV_X1 U9785 ( .A(n13073), .ZN(n13679) );
  AND2_X2 U9786 ( .A1(n8735), .A2(n11109), .ZN(n16042) );
  NAND2_X1 U9787 ( .A1(n8693), .A2(n13710), .ZN(n10638) );
  INV_X1 U9788 ( .A(SI_14_), .ZN(n15315) );
  NAND2_X1 U9789 ( .A1(n10268), .A2(n10254), .ZN(n13907) );
  INV_X1 U9790 ( .A(n14210), .ZN(n13918) );
  INV_X1 U9791 ( .A(n12334), .ZN(n13919) );
  INV_X1 U9792 ( .A(n10785), .ZN(n13928) );
  OR2_X1 U9793 ( .A1(n10455), .A2(P2_U3088), .ZN(n15534) );
  INV_X1 U9794 ( .A(n14290), .ZN(n14261) );
  AND3_X1 U9795 ( .A1(n14214), .A2(n14213), .A3(n14212), .ZN(n14359) );
  INV_X1 U9796 ( .A(n14263), .ZN(n14198) );
  INV_X2 U9797 ( .A(n16035), .ZN(n16034) );
  INV_X1 U9798 ( .A(n14295), .ZN(n14373) );
  NAND2_X1 U9799 ( .A1(n14371), .A2(n14347), .ZN(n14402) );
  OR2_X1 U9800 ( .A1(n15452), .A2(n15450), .ZN(n15451) );
  OAI21_X1 U9801 ( .B1(n10209), .B2(P2_D_REG_0__SCAN_IN), .A(n10208), .ZN(
        n15454) );
  INV_X1 U9802 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14413) );
  INV_X1 U9803 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10741) );
  AND2_X1 U9804 ( .A1(n10086), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10586) );
  INV_X1 U9805 ( .A(n12872), .ZN(n14714) );
  INV_X1 U9806 ( .A(n14608), .ZN(n14721) );
  INV_X1 U9807 ( .A(n15566), .ZN(n11897) );
  INV_X1 U9808 ( .A(n15544), .ZN(n15570) );
  NAND2_X1 U9809 ( .A1(n15054), .A2(n10812), .ZN(n15942) );
  NAND2_X1 U9810 ( .A1(n15054), .A2(n14816), .ZN(n15057) );
  NAND2_X1 U9811 ( .A1(n15054), .A2(n11558), .ZN(n15061) );
  AND2_X2 U9812 ( .A1(n10103), .A2(n10096), .ZN(n16014) );
  INV_X1 U9813 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n12273) );
  INV_X1 U9814 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10765) );
  INV_X2 U9815 ( .A(n13240), .ZN(P3_U3897) );
  OAI21_X1 U9816 ( .B1(n8739), .B2(n8727), .A(n8726), .ZN(P3_U3488) );
  AND2_X1 U9817 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10437), .ZN(P2_U3947) );
  AND2_X2 U9818 ( .A1(n10570), .A2(n10586), .ZN(P1_U4016) );
  INV_X1 U9819 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n14409) );
  INV_X1 U9820 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n15431) );
  AOI22_X1 U9821 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n14409), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n15431), .ZN(n8587) );
  INV_X1 U9822 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15434) );
  AOI22_X1 U9823 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n14413), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n15434), .ZN(n8192) );
  AOI22_X1 U9824 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n12481), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n7369), .ZN(n8560) );
  INV_X1 U9825 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n15442) );
  AOI22_X1 U9826 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(P1_DATAO_REG_23__SCAN_IN), .B1(n14423), .B2(n15442), .ZN(n8533) );
  AOI22_X1 U9827 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n12463), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n7682), .ZN(n8519) );
  INV_X1 U9828 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12355) );
  AOI22_X1 U9829 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n12359), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n12355), .ZN(n8510) );
  AOI22_X1 U9830 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n12067), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n7694), .ZN(n8484) );
  XNOR2_X1 U9831 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .ZN(n8468) );
  XNOR2_X1 U9832 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n8388) );
  NAND2_X1 U9833 ( .A1(n8232), .A2(n8231), .ZN(n8230) );
  INV_X1 U9834 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10304) );
  NAND2_X1 U9835 ( .A1(n10304), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8105) );
  NAND2_X1 U9836 ( .A1(n8230), .A2(n8105), .ZN(n8209) );
  XNOR2_X1 U9837 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8208) );
  NAND2_X1 U9838 ( .A1(n8209), .A2(n8208), .ZN(n8107) );
  INV_X1 U9839 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10310) );
  NAND2_X1 U9840 ( .A1(n10310), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8106) );
  NAND2_X1 U9841 ( .A1(n8107), .A2(n8106), .ZN(n8248) );
  XNOR2_X1 U9842 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8247) );
  NAND2_X1 U9843 ( .A1(n8248), .A2(n8247), .ZN(n8110) );
  INV_X1 U9844 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n8108) );
  NAND2_X1 U9845 ( .A1(n8108), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8109) );
  NAND2_X1 U9846 ( .A1(n8110), .A2(n8109), .ZN(n8261) );
  NAND2_X1 U9847 ( .A1(n8261), .A2(n8260), .ZN(n8112) );
  NAND2_X1 U9848 ( .A1(n10298), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8111) );
  NAND2_X1 U9849 ( .A1(n8112), .A2(n8111), .ZN(n8276) );
  INV_X1 U9850 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n8113) );
  NAND2_X1 U9851 ( .A1(n8113), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8114) );
  NAND2_X1 U9852 ( .A1(n10315), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8116) );
  NAND2_X1 U9853 ( .A1(n8341), .A2(n8339), .ZN(n8118) );
  NAND2_X1 U9854 ( .A1(n10434), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8117) );
  NAND2_X1 U9855 ( .A1(n8118), .A2(n8117), .ZN(n8362) );
  XNOR2_X1 U9856 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n8361) );
  XNOR2_X1 U9857 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8375) );
  NAND2_X1 U9858 ( .A1(n8120), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8121) );
  NAND2_X1 U9859 ( .A1(n8395), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8124) );
  NAND2_X1 U9860 ( .A1(n10765), .A2(n8122), .ZN(n8123) );
  XNOR2_X1 U9861 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8412) );
  INV_X1 U9862 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n8125) );
  NAND2_X1 U9863 ( .A1(n8125), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8126) );
  XNOR2_X1 U9864 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n8425) );
  NAND2_X1 U9865 ( .A1(n11424), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8127) );
  XNOR2_X1 U9866 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .ZN(n8453) );
  NAND2_X1 U9867 ( .A1(n11572), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8128) );
  NAND2_X1 U9868 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n8130), .ZN(n8131) );
  NAND2_X1 U9869 ( .A1(n8560), .A2(n8562), .ZN(n8133) );
  AOI22_X1 U9870 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n14415), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n8134), .ZN(n8574) );
  NAND2_X1 U9871 ( .A1(n8192), .A2(n8194), .ZN(n8136) );
  NAND2_X1 U9872 ( .A1(n8587), .A2(n8589), .ZN(n8137) );
  INV_X1 U9873 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n12958) );
  INV_X1 U9874 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14404) );
  OAI22_X1 U9875 ( .A1(n12958), .A2(n14404), .B1(P1_DATAO_REG_29__SCAN_IN), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12488) );
  INV_X1 U9876 ( .A(n12488), .ZN(n8138) );
  XNOR2_X1 U9877 ( .A(n12489), .B(n8138), .ZN(n13722) );
  XNOR2_X2 U9878 ( .A(n8150), .B(n8149), .ZN(n8663) );
  XNOR2_X2 U9879 ( .A(n8152), .B(n8151), .ZN(n8664) );
  INV_X1 U9880 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8153) );
  NAND3_X1 U9881 ( .A1(n8155), .A2(n8154), .A3(n8153), .ZN(n8156) );
  NAND2_X1 U9882 ( .A1(n8156), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n8161) );
  INV_X1 U9883 ( .A(P2_RD_REG_SCAN_IN), .ZN(n8157) );
  NAND3_X1 U9884 ( .A1(n8157), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n8159) );
  NAND2_X1 U9885 ( .A1(n8159), .A2(n8158), .ZN(n8160) );
  NAND2_X2 U9886 ( .A1(n7157), .A2(n10276), .ZN(n12509) );
  NAND2_X1 U9887 ( .A1(n13722), .A2(n12496), .ZN(n8163) );
  INV_X1 U9888 ( .A(SI_29_), .ZN(n13724) );
  OR2_X1 U9889 ( .A1(n7158), .A2(n13724), .ZN(n8162) );
  NAND2_X1 U9890 ( .A1(n8163), .A2(n8162), .ZN(n8722) );
  NAND2_X1 U9891 ( .A1(n15356), .A2(n15169), .ZN(n8268) );
  INV_X1 U9892 ( .A(n8268), .ZN(n8165) );
  NAND2_X1 U9893 ( .A1(n8165), .A2(n8164), .ZN(n8289) );
  INV_X1 U9894 ( .A(n8304), .ZN(n8167) );
  NAND2_X1 U9895 ( .A1(n15360), .A2(n15269), .ZN(n8168) );
  INV_X1 U9896 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8171) );
  INV_X1 U9897 ( .A(n8419), .ZN(n8173) );
  INV_X1 U9898 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n8177) );
  INV_X1 U9899 ( .A(n8565), .ZN(n8179) );
  INV_X1 U9900 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n15267) );
  INV_X1 U9901 ( .A(n8578), .ZN(n8180) );
  INV_X1 U9902 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n15162) );
  INV_X1 U9903 ( .A(n8592), .ZN(n8182) );
  INV_X1 U9904 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n8181) );
  NAND2_X1 U9905 ( .A1(n8182), .A2(n8181), .ZN(n13371) );
  INV_X1 U9906 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8736) );
  NAND2_X1 U9907 ( .A1(n8567), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8189) );
  NAND2_X1 U9908 ( .A1(n8665), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8188) );
  OAI211_X1 U9909 ( .C1(n12503), .C2(n8736), .A(n8189), .B(n8188), .ZN(n8190)
         );
  INV_X1 U9910 ( .A(n8190), .ZN(n8191) );
  NAND2_X1 U9911 ( .A1(n8722), .A2(n13031), .ZN(n12687) );
  NAND2_X1 U9912 ( .A1(n12637), .A2(n12687), .ZN(n12656) );
  INV_X1 U9913 ( .A(n8192), .ZN(n8193) );
  NAND2_X1 U9914 ( .A1(n13727), .A2(n12496), .ZN(n8196) );
  INV_X1 U9915 ( .A(SI_27_), .ZN(n15289) );
  OR2_X1 U9916 ( .A1(n7158), .A2(n15289), .ZN(n8195) );
  NAND2_X1 U9917 ( .A1(n8580), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8197) );
  NAND2_X1 U9918 ( .A1(n8592), .A2(n8197), .ZN(n13405) );
  INV_X1 U9919 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13663) );
  NAND2_X1 U9920 ( .A1(n8665), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8199) );
  NAND2_X1 U9921 ( .A1(n8567), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8198) );
  OAI211_X1 U9922 ( .C1(n13663), .C2(n12503), .A(n8199), .B(n8198), .ZN(n8200)
         );
  OR2_X1 U9923 ( .A1(n8660), .A2(n13412), .ZN(n12525) );
  NAND2_X1 U9924 ( .A1(n8660), .A2(n13412), .ZN(n12524) );
  INV_X1 U9925 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n8201) );
  INV_X1 U9926 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10884) );
  INV_X1 U9927 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n8202) );
  OR2_X1 U9928 ( .A1(n8242), .A2(n8202), .ZN(n8205) );
  INV_X1 U9929 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n8203) );
  OR2_X1 U9930 ( .A1(n8224), .A2(n8203), .ZN(n8204) );
  XNOR2_X1 U9931 ( .A(n8209), .B(n8208), .ZN(n10286) );
  OR2_X1 U9932 ( .A1(n12509), .A2(n10286), .ZN(n8213) );
  XNOR2_X1 U9933 ( .A(n8211), .B(P3_IR_REG_2__SCAN_IN), .ZN(n10885) );
  OR2_X1 U9934 ( .A1(n10850), .A2(n10885), .ZN(n8212) );
  INV_X1 U9935 ( .A(n11311), .ZN(n15845) );
  NAND2_X1 U9936 ( .A1(n11334), .A2(n11311), .ZN(n12543) );
  NAND2_X1 U9937 ( .A1(n8506), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8220) );
  INV_X1 U9938 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10883) );
  OR2_X1 U9939 ( .A1(n8240), .A2(n10883), .ZN(n8219) );
  INV_X1 U9940 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11411) );
  INV_X1 U9941 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n8216) );
  OR2_X1 U9942 ( .A1(n8224), .A2(n8216), .ZN(n8217) );
  INV_X1 U9943 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8808) );
  XNOR2_X1 U9944 ( .A(n8808), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8221) );
  MUX2_X1 U9945 ( .A(n8221), .B(SI_0_), .S(n10297), .Z(n10272) );
  MUX2_X1 U9946 ( .A(P3_IR_REG_0__SCAN_IN), .B(n10272), .S(n10850), .Z(n11314)
         );
  NAND2_X1 U9947 ( .A1(n11016), .A2(n11314), .ZN(n11313) );
  NAND2_X1 U9948 ( .A1(n8215), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8228) );
  INV_X1 U9949 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10877) );
  INV_X1 U9950 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n8222) );
  INV_X1 U9951 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n8223) );
  OR2_X1 U9952 ( .A1(n8224), .A2(n8223), .ZN(n8225) );
  OAI21_X1 U9953 ( .B1(n8232), .B2(n8231), .A(n8230), .ZN(n8233) );
  INV_X1 U9954 ( .A(n8233), .ZN(n10274) );
  OR2_X1 U9955 ( .A1(n12509), .A2(n10274), .ZN(n8236) );
  INV_X1 U9956 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n8235) );
  NAND2_X1 U9957 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n8234) );
  NAND2_X1 U9958 ( .A1(n11313), .A2(n12538), .ZN(n8237) );
  NAND2_X1 U9959 ( .A1(n8237), .A2(n12533), .ZN(n15844) );
  INV_X1 U9960 ( .A(n15844), .ZN(n8238) );
  NAND2_X1 U9961 ( .A1(n8567), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8246) );
  INV_X1 U9962 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10890) );
  OR2_X1 U9963 ( .A1(n8240), .A2(n10890), .ZN(n8245) );
  INV_X1 U9964 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n8241) );
  OR2_X1 U9965 ( .A1(n8242), .A2(n8241), .ZN(n8244) );
  OR2_X1 U9966 ( .A1(n8224), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8243) );
  OR2_X1 U9967 ( .A1(n12510), .A2(SI_3_), .ZN(n8253) );
  XNOR2_X1 U9968 ( .A(n8248), .B(n8247), .ZN(n10290) );
  OR2_X1 U9969 ( .A1(n12509), .A2(n10290), .ZN(n8252) );
  NAND2_X1 U9970 ( .A1(n8249), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8250) );
  XNOR2_X1 U9971 ( .A(n8250), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10891) );
  OR2_X1 U9972 ( .A1(n7157), .A2(n10891), .ZN(n8251) );
  INV_X1 U9973 ( .A(n11846), .ZN(n11440) );
  NAND2_X1 U9974 ( .A1(n15847), .A2(n11440), .ZN(n12547) );
  NAND2_X1 U9975 ( .A1(n11662), .A2(n11846), .ZN(n12546) );
  NAND2_X1 U9976 ( .A1(n11332), .A2(n12546), .ZN(n11661) );
  NAND2_X1 U9977 ( .A1(n8665), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8259) );
  INV_X1 U9978 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11670) );
  OR2_X1 U9979 ( .A1(n8495), .A2(n11670), .ZN(n8258) );
  NAND2_X1 U9980 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8254) );
  AND2_X1 U9981 ( .A1(n8268), .A2(n8254), .ZN(n11671) );
  OR2_X1 U9982 ( .A1(n8224), .A2(n11671), .ZN(n8257) );
  INV_X1 U9983 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n8255) );
  OR2_X1 U9984 ( .A1(n12503), .A2(n8255), .ZN(n8256) );
  OR2_X1 U9985 ( .A1(n12510), .A2(SI_4_), .ZN(n8265) );
  XNOR2_X1 U9986 ( .A(n8261), .B(n8260), .ZN(n10293) );
  OR2_X1 U9987 ( .A1(n12509), .A2(n10293), .ZN(n8264) );
  OR2_X1 U9988 ( .A1(n8249), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n8277) );
  NAND2_X1 U9989 ( .A1(n8277), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8262) );
  OR2_X1 U9990 ( .A1(n10850), .A2(n10985), .ZN(n8263) );
  NAND2_X1 U9991 ( .A1(n11856), .A2(n15906), .ZN(n12552) );
  INV_X1 U9992 ( .A(n15906), .ZN(n8266) );
  NAND2_X1 U9993 ( .A1(n13251), .A2(n8266), .ZN(n12553) );
  NAND2_X1 U9994 ( .A1(n12552), .A2(n12553), .ZN(n11664) );
  INV_X1 U9995 ( .A(n11664), .ZN(n12663) );
  NAND2_X1 U9996 ( .A1(n11661), .A2(n12663), .ZN(n11660) );
  NAND2_X1 U9997 ( .A1(n11660), .A2(n12552), .ZN(n11851) );
  NAND2_X1 U9998 ( .A1(n8567), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8274) );
  INV_X1 U9999 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n8267) );
  OR2_X1 U10000 ( .A1(n8240), .A2(n8267), .ZN(n8273) );
  NAND2_X1 U10001 ( .A1(n8268), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8269) );
  AND2_X1 U10002 ( .A1(n8289), .A2(n8269), .ZN(n13130) );
  OR2_X1 U10003 ( .A1(n8224), .A2(n13130), .ZN(n8272) );
  INV_X1 U10004 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n8270) );
  OR2_X1 U10005 ( .A1(n12503), .A2(n8270), .ZN(n8271) );
  OR2_X1 U10006 ( .A1(n12510), .A2(SI_5_), .ZN(n8287) );
  XNOR2_X1 U10007 ( .A(n8276), .B(n8275), .ZN(n10288) );
  OR2_X1 U10008 ( .A1(n12509), .A2(n10288), .ZN(n8286) );
  INV_X1 U10009 ( .A(n8277), .ZN(n8279) );
  NAND2_X1 U10010 ( .A1(n8279), .A2(n8278), .ZN(n8281) );
  NAND2_X1 U10011 ( .A1(n8281), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8280) );
  MUX2_X1 U10012 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8280), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n8284) );
  INV_X1 U10013 ( .A(n8281), .ZN(n8283) );
  NAND2_X1 U10014 ( .A1(n8283), .A2(n8282), .ZN(n8296) );
  OR2_X1 U10015 ( .A1(n7157), .A2(n10978), .ZN(n8285) );
  NAND2_X1 U10016 ( .A1(n11724), .A2(n13129), .ZN(n12556) );
  INV_X1 U10017 ( .A(n13129), .ZN(n12021) );
  NAND2_X1 U10018 ( .A1(n13250), .A2(n12021), .ZN(n12557) );
  NAND2_X1 U10019 ( .A1(n11851), .A2(n12662), .ZN(n11850) );
  NAND2_X1 U10020 ( .A1(n8665), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8295) );
  INV_X1 U10021 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n8288) );
  OR2_X1 U10022 ( .A1(n8495), .A2(n8288), .ZN(n8294) );
  NAND2_X1 U10023 ( .A1(n8289), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8290) );
  AND2_X1 U10024 ( .A1(n8304), .A2(n8290), .ZN(n12043) );
  OR2_X1 U10025 ( .A1(n8224), .A2(n12043), .ZN(n8293) );
  INV_X1 U10026 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n8291) );
  OR2_X1 U10027 ( .A1(n12503), .A2(n8291), .ZN(n8292) );
  NAND2_X1 U10028 ( .A1(n8296), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8298) );
  XNOR2_X1 U10029 ( .A(n8297), .B(n8298), .ZN(n10991) );
  INV_X1 U10030 ( .A(SI_6_), .ZN(n15278) );
  OR2_X1 U10031 ( .A1(n7158), .A2(n15278), .ZN(n8302) );
  XNOR2_X1 U10032 ( .A(n10318), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8299) );
  XNOR2_X1 U10033 ( .A(n8300), .B(n8299), .ZN(n10275) );
  OR2_X1 U10034 ( .A1(n12509), .A2(n10275), .ZN(n8301) );
  OAI211_X1 U10035 ( .C1(n7157), .C2(n10991), .A(n8302), .B(n8301), .ZN(n11908) );
  NAND2_X1 U10036 ( .A1(n11918), .A2(n11908), .ZN(n12560) );
  INV_X1 U10037 ( .A(n11908), .ZN(n12044) );
  NAND2_X1 U10038 ( .A1(n13249), .A2(n12044), .ZN(n12561) );
  NAND2_X1 U10039 ( .A1(n8567), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8310) );
  INV_X1 U10040 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n8303) );
  OR2_X1 U10041 ( .A1(n8240), .A2(n8303), .ZN(n8309) );
  NAND2_X1 U10042 ( .A1(n8304), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8305) );
  AND2_X1 U10043 ( .A1(n8333), .A2(n8305), .ZN(n12207) );
  OR2_X1 U10044 ( .A1(n8224), .A2(n12207), .ZN(n8308) );
  INV_X1 U10045 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n8306) );
  OR2_X1 U10046 ( .A1(n12503), .A2(n8306), .ZN(n8307) );
  INV_X1 U10047 ( .A(n8311), .ZN(n8312) );
  XNOR2_X1 U10048 ( .A(n8313), .B(n8312), .ZN(n10282) );
  OR2_X1 U10049 ( .A1(n12509), .A2(n10282), .ZN(n8318) );
  OR2_X1 U10050 ( .A1(n7158), .A2(SI_7_), .ZN(n8317) );
  NAND2_X1 U10051 ( .A1(n8314), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8315) );
  XNOR2_X1 U10052 ( .A(n8315), .B(P3_IR_REG_7__SCAN_IN), .ZN(n11808) );
  OR2_X1 U10053 ( .A1(n7157), .A2(n11808), .ZN(n8316) );
  NAND2_X1 U10054 ( .A1(n12242), .A2(n11994), .ZN(n12565) );
  INV_X1 U10055 ( .A(n11994), .ZN(n12208) );
  NAND2_X1 U10056 ( .A1(n13248), .A2(n12208), .ZN(n12566) );
  NAND2_X1 U10057 ( .A1(n12565), .A2(n12566), .ZN(n12562) );
  INV_X1 U10058 ( .A(n12562), .ZN(n12659) );
  NAND2_X1 U10059 ( .A1(n11986), .A2(n12565), .ZN(n12244) );
  NAND2_X1 U10060 ( .A1(n8665), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8323) );
  INV_X1 U10061 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n12245) );
  OR2_X1 U10062 ( .A1(n8495), .A2(n12245), .ZN(n8322) );
  XNOR2_X1 U10063 ( .A(n8333), .B(n15269), .ZN(n12246) );
  OR2_X1 U10064 ( .A1(n8224), .A2(n12246), .ZN(n8321) );
  INV_X1 U10065 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n8319) );
  OR2_X1 U10066 ( .A1(n12503), .A2(n8319), .ZN(n8320) );
  NAND4_X1 U10067 ( .A1(n8323), .A2(n8322), .A3(n8321), .A4(n8320), .ZN(n13247) );
  OR2_X1 U10068 ( .A1(n8324), .A2(n8344), .ZN(n8325) );
  XNOR2_X1 U10069 ( .A(n8325), .B(P3_IR_REG_8__SCAN_IN), .ZN(n15755) );
  INV_X1 U10070 ( .A(n15755), .ZN(n11825) );
  XNOR2_X1 U10071 ( .A(n8327), .B(n8326), .ZN(n10279) );
  OR2_X1 U10072 ( .A1(n12509), .A2(n10279), .ZN(n8329) );
  INV_X1 U10073 ( .A(SI_8_), .ZN(n15207) );
  OR2_X1 U10074 ( .A1(n7158), .A2(n15207), .ZN(n8328) );
  OAI211_X1 U10075 ( .C1(n10850), .C2(n11825), .A(n8329), .B(n8328), .ZN(
        n12269) );
  XNOR2_X1 U10076 ( .A(n13247), .B(n12269), .ZN(n12664) );
  NAND2_X1 U10077 ( .A1(n12568), .A2(n12269), .ZN(n8330) );
  NAND2_X1 U10078 ( .A1(n8506), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8338) );
  INV_X1 U10079 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n8331) );
  OR2_X1 U10080 ( .A1(n8240), .A2(n8331), .ZN(n8337) );
  INV_X1 U10081 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n8332) );
  OR2_X1 U10082 ( .A1(n8495), .A2(n8332), .ZN(n8336) );
  OAI21_X1 U10083 ( .B1(n8333), .B2(P3_REG3_REG_8__SCAN_IN), .A(
        P3_REG3_REG_9__SCAN_IN), .ZN(n8334) );
  AND2_X1 U10084 ( .A1(n8334), .A2(n8354), .ZN(n12257) );
  OR2_X1 U10085 ( .A1(n8224), .A2(n12257), .ZN(n8335) );
  NAND4_X1 U10086 ( .A1(n8338), .A2(n8337), .A3(n8336), .A4(n8335), .ZN(n13246) );
  INV_X1 U10087 ( .A(n8339), .ZN(n8340) );
  XNOR2_X1 U10088 ( .A(n8341), .B(n8340), .ZN(n10280) );
  OR2_X1 U10089 ( .A1(n12509), .A2(n10280), .ZN(n8351) );
  OR2_X1 U10090 ( .A1(n7158), .A2(SI_9_), .ZN(n8350) );
  INV_X1 U10091 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8342) );
  AND2_X1 U10092 ( .A1(n8324), .A2(n8342), .ZN(n8346) );
  NOR2_X1 U10093 ( .A1(n8346), .A2(n8344), .ZN(n8343) );
  MUX2_X1 U10094 ( .A(n8344), .B(n8343), .S(P3_IR_REG_9__SCAN_IN), .Z(n8348)
         );
  NAND2_X1 U10095 ( .A1(n8346), .A2(n8345), .ZN(n8364) );
  INV_X1 U10096 ( .A(n8364), .ZN(n8347) );
  OR2_X1 U10097 ( .A1(n7157), .A2(n15780), .ZN(n8349) );
  NOR2_X1 U10098 ( .A1(n13246), .A2(n15929), .ZN(n12575) );
  NAND2_X1 U10099 ( .A1(n13246), .A2(n15929), .ZN(n12251) );
  NAND2_X1 U10100 ( .A1(n8506), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8360) );
  INV_X1 U10101 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n8353) );
  OR2_X1 U10102 ( .A1(n8495), .A2(n8353), .ZN(n8359) );
  NAND2_X1 U10103 ( .A1(n8354), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8355) );
  AND2_X1 U10104 ( .A1(n8369), .A2(n8355), .ZN(n12418) );
  OR2_X1 U10105 ( .A1(n8224), .A2(n12418), .ZN(n8358) );
  INV_X1 U10106 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n8356) );
  OR2_X1 U10107 ( .A1(n8240), .A2(n8356), .ZN(n8357) );
  XNOR2_X1 U10108 ( .A(n8362), .B(n8361), .ZN(n10285) );
  NAND2_X1 U10109 ( .A1(n10285), .A2(n12496), .ZN(n8368) );
  OR2_X1 U10110 ( .A1(n7158), .A2(SI_10_), .ZN(n8367) );
  NAND2_X1 U10111 ( .A1(n8364), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8363) );
  MUX2_X1 U10112 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8363), .S(
        P3_IR_REG_10__SCAN_IN), .Z(n8365) );
  NAND2_X1 U10113 ( .A1(n8365), .A2(n8390), .ZN(n11830) );
  INV_X1 U10114 ( .A(n11830), .ZN(n15789) );
  OR2_X1 U10115 ( .A1(n10850), .A2(n15789), .ZN(n8366) );
  NAND2_X1 U10116 ( .A1(n12423), .A2(n12422), .ZN(n12532) );
  INV_X1 U10117 ( .A(n12422), .ZN(n15957) );
  NAND2_X1 U10118 ( .A1(n13245), .A2(n15957), .ZN(n12579) );
  NAND2_X1 U10119 ( .A1(n12532), .A2(n12579), .ZN(n12576) );
  NAND2_X1 U10120 ( .A1(n8506), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8374) );
  INV_X1 U10121 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11800) );
  OR2_X1 U10122 ( .A1(n8495), .A2(n11800), .ZN(n8373) );
  NAND2_X1 U10123 ( .A1(n8369), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8370) );
  AND2_X1 U10124 ( .A1(n8381), .A2(n8370), .ZN(n13189) );
  OR2_X1 U10125 ( .A1(n8224), .A2(n13189), .ZN(n8372) );
  INV_X1 U10126 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n11799) );
  OR2_X1 U10127 ( .A1(n8240), .A2(n11799), .ZN(n8371) );
  NAND4_X1 U10128 ( .A1(n8374), .A2(n8373), .A3(n8372), .A4(n8371), .ZN(n13244) );
  XNOR2_X1 U10129 ( .A(n8376), .B(n8375), .ZN(n10295) );
  NAND2_X1 U10130 ( .A1(n10295), .A2(n12496), .ZN(n8380) );
  NAND2_X1 U10131 ( .A1(n8390), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8378) );
  XNOR2_X1 U10132 ( .A(n8378), .B(n8377), .ZN(n11814) );
  AOI22_X1 U10133 ( .A1(n8490), .A2(n15275), .B1(n8489), .B2(n11814), .ZN(
        n8379) );
  NAND2_X1 U10134 ( .A1(n13048), .A2(n13191), .ZN(n12581) );
  NAND2_X1 U10135 ( .A1(n13244), .A2(n12471), .ZN(n12583) );
  NAND2_X1 U10136 ( .A1(n12581), .A2(n12583), .ZN(n12968) );
  NAND2_X1 U10137 ( .A1(n8567), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8387) );
  INV_X1 U10138 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n15978) );
  OR2_X1 U10139 ( .A1(n8240), .A2(n15978), .ZN(n8386) );
  NAND2_X1 U10140 ( .A1(n8381), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8382) );
  AND2_X1 U10141 ( .A1(n8405), .A2(n8382), .ZN(n12436) );
  OR2_X1 U10142 ( .A1(n8224), .A2(n12436), .ZN(n8385) );
  INV_X1 U10143 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n8383) );
  OR2_X1 U10144 ( .A1(n12503), .A2(n8383), .ZN(n8384) );
  XNOR2_X1 U10145 ( .A(n8389), .B(n8388), .ZN(n10299) );
  NAND2_X1 U10146 ( .A1(n10299), .A2(n12496), .ZN(n8393) );
  OR2_X1 U10147 ( .A1(n8397), .A2(n8344), .ZN(n8391) );
  XNOR2_X1 U10148 ( .A(n8391), .B(n8396), .ZN(n12114) );
  AOI22_X1 U10149 ( .A1(n8490), .A2(n15172), .B1(n8489), .B2(n12114), .ZN(
        n8392) );
  NAND2_X1 U10150 ( .A1(n8393), .A2(n8392), .ZN(n15971) );
  NAND2_X1 U10151 ( .A1(n15971), .A2(n13243), .ZN(n12972) );
  NAND2_X1 U10152 ( .A1(n13054), .A2(n12972), .ZN(n12580) );
  INV_X1 U10153 ( .A(n12583), .ZN(n8394) );
  XNOR2_X1 U10154 ( .A(n8395), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n10333) );
  NAND2_X1 U10155 ( .A1(n10333), .A2(n12496), .ZN(n8404) );
  INV_X1 U10156 ( .A(SI_13_), .ZN(n15318) );
  NOR2_X1 U10157 ( .A1(n8401), .A2(n8344), .ZN(n8398) );
  MUX2_X1 U10158 ( .A(n8344), .B(n8398), .S(P3_IR_REG_13__SCAN_IN), .Z(n8399)
         );
  INV_X1 U10159 ( .A(n8399), .ZN(n8402) );
  INV_X1 U10160 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8400) );
  NAND2_X1 U10161 ( .A1(n8401), .A2(n8400), .ZN(n8415) );
  NAND2_X1 U10162 ( .A1(n8402), .A2(n8415), .ZN(n12182) );
  AOI22_X1 U10163 ( .A1(n8490), .A2(n15318), .B1(n8489), .B2(n12182), .ZN(
        n8403) );
  NAND2_X1 U10164 ( .A1(n8404), .A2(n8403), .ZN(n12589) );
  NAND2_X1 U10165 ( .A1(n8506), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8410) );
  INV_X1 U10166 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12475) );
  OR2_X1 U10167 ( .A1(n8495), .A2(n12475), .ZN(n8409) );
  NAND2_X1 U10168 ( .A1(n8405), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8406) );
  AND2_X1 U10169 ( .A1(n8419), .A2(n8406), .ZN(n13176) );
  OR2_X1 U10170 ( .A1(n8224), .A2(n13176), .ZN(n8408) );
  INV_X1 U10171 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n12121) );
  OR2_X1 U10172 ( .A1(n8240), .A2(n12121), .ZN(n8407) );
  XNOR2_X1 U10173 ( .A(n12589), .B(n13581), .ZN(n13056) );
  INV_X1 U10174 ( .A(n13581), .ZN(n13242) );
  OR2_X1 U10175 ( .A1(n12589), .A2(n13242), .ZN(n12588) );
  XNOR2_X1 U10176 ( .A(n8413), .B(n8412), .ZN(n10374) );
  NAND2_X1 U10177 ( .A1(n10374), .A2(n12496), .ZN(n8418) );
  NAND2_X1 U10178 ( .A1(n8415), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8414) );
  MUX2_X1 U10179 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8414), .S(
        P3_IR_REG_14__SCAN_IN), .Z(n8416) );
  NAND2_X1 U10180 ( .A1(n8416), .A2(n8439), .ZN(n13263) );
  AOI22_X1 U10181 ( .A1(n8490), .A2(n15315), .B1(n8489), .B2(n13263), .ZN(
        n8417) );
  NAND2_X1 U10182 ( .A1(n8506), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8424) );
  INV_X1 U10183 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n13589) );
  OR2_X1 U10184 ( .A1(n8495), .A2(n13589), .ZN(n8423) );
  NAND2_X1 U10185 ( .A1(n8419), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8420) );
  AND2_X1 U10186 ( .A1(n8431), .A2(n8420), .ZN(n13588) );
  OR2_X1 U10187 ( .A1(n8224), .A2(n13588), .ZN(n8422) );
  INV_X1 U10188 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13654) );
  OR2_X1 U10189 ( .A1(n8240), .A2(n13654), .ZN(n8421) );
  NAND4_X1 U10190 ( .A1(n8424), .A2(n8423), .A3(n8422), .A4(n8421), .ZN(n13564) );
  OR2_X1 U10191 ( .A1(n13706), .A2(n13564), .ZN(n12594) );
  NAND2_X1 U10192 ( .A1(n13706), .A2(n13564), .ZN(n12595) );
  XNOR2_X1 U10193 ( .A(n8426), .B(n8425), .ZN(n10435) );
  NAND2_X1 U10194 ( .A1(n10435), .A2(n12496), .ZN(n8430) );
  NAND2_X1 U10195 ( .A1(n8439), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8428) );
  XNOR2_X1 U10196 ( .A(n8427), .B(n8428), .ZN(n13285) );
  AOI22_X1 U10197 ( .A1(n8490), .A2(n15313), .B1(n8489), .B2(n13285), .ZN(
        n8429) );
  NAND2_X1 U10198 ( .A1(n8430), .A2(n8429), .ZN(n13651) );
  NAND2_X1 U10199 ( .A1(n8506), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8436) );
  INV_X1 U10200 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n13571) );
  OR2_X1 U10201 ( .A1(n8495), .A2(n13571), .ZN(n8435) );
  NAND2_X1 U10202 ( .A1(n8431), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8432) );
  AND2_X1 U10203 ( .A1(n8445), .A2(n8432), .ZN(n13570) );
  OR2_X1 U10204 ( .A1(n8224), .A2(n13570), .ZN(n8434) );
  INV_X1 U10205 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13265) );
  OR2_X1 U10206 ( .A1(n8240), .A2(n13265), .ZN(n8433) );
  NAND4_X1 U10207 ( .A1(n8436), .A2(n8435), .A3(n8434), .A4(n8433), .ZN(n13551) );
  OR2_X1 U10208 ( .A1(n13651), .A2(n13551), .ZN(n12603) );
  NAND2_X1 U10209 ( .A1(n13651), .A2(n13551), .ZN(n12600) );
  NAND2_X1 U10210 ( .A1(n12603), .A2(n12600), .ZN(n13567) );
  NAND2_X1 U10211 ( .A1(n13569), .A2(n8437), .ZN(n13568) );
  NAND2_X1 U10212 ( .A1(n13568), .A2(n12603), .ZN(n13559) );
  XNOR2_X1 U10213 ( .A(n8438), .B(n7288), .ZN(n10608) );
  NAND2_X1 U10214 ( .A1(n10608), .A2(n12496), .ZN(n8444) );
  OAI21_X1 U10215 ( .B1(n8439), .B2(P3_IR_REG_15__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8441) );
  NAND2_X1 U10216 ( .A1(n8441), .A2(n8440), .ZN(n8455) );
  OR2_X1 U10217 ( .A1(n8441), .A2(n8440), .ZN(n8442) );
  AND2_X1 U10218 ( .A1(n8455), .A2(n8442), .ZN(n13289) );
  AOI22_X1 U10219 ( .A1(n13289), .A2(n8489), .B1(n8490), .B2(SI_16_), .ZN(
        n8443) );
  NAND2_X1 U10220 ( .A1(n8444), .A2(n8443), .ZN(n13644) );
  NAND2_X1 U10221 ( .A1(n8506), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8451) );
  INV_X1 U10222 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13555) );
  OR2_X1 U10223 ( .A1(n8495), .A2(n13555), .ZN(n8450) );
  NAND2_X1 U10224 ( .A1(n8445), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8446) );
  AND2_X1 U10225 ( .A1(n8461), .A2(n8446), .ZN(n13554) );
  OR2_X1 U10226 ( .A1(n8224), .A2(n13554), .ZN(n8449) );
  INV_X1 U10227 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n8447) );
  OR2_X1 U10228 ( .A1(n8240), .A2(n8447), .ZN(n8448) );
  OR2_X1 U10229 ( .A1(n13644), .A2(n13535), .ZN(n12601) );
  NAND2_X1 U10230 ( .A1(n13644), .A2(n13535), .ZN(n12598) );
  NAND2_X1 U10231 ( .A1(n12601), .A2(n12598), .ZN(n13549) );
  NAND2_X1 U10232 ( .A1(n13559), .A2(n13558), .ZN(n8452) );
  NAND2_X1 U10233 ( .A1(n8452), .A2(n12598), .ZN(n13539) );
  XNOR2_X1 U10234 ( .A(n8454), .B(n8453), .ZN(n10612) );
  NAND2_X1 U10235 ( .A1(n10612), .A2(n12496), .ZN(n8460) );
  NAND2_X1 U10236 ( .A1(n8455), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8457) );
  INV_X1 U10237 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8456) );
  XNOR2_X1 U10238 ( .A(n8457), .B(n8456), .ZN(n13318) );
  NOR2_X1 U10239 ( .A1(n7158), .A2(SI_17_), .ZN(n8458) );
  AOI21_X1 U10240 ( .B1(n13318), .B2(n8489), .A(n8458), .ZN(n8459) );
  NAND2_X1 U10241 ( .A1(n8461), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8462) );
  NAND2_X1 U10242 ( .A1(n8477), .A2(n8462), .ZN(n13540) );
  NAND2_X1 U10243 ( .A1(n8597), .A2(n13540), .ZN(n8467) );
  INV_X1 U10244 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n8463) );
  OR2_X1 U10245 ( .A1(n8495), .A2(n8463), .ZN(n8466) );
  INV_X1 U10246 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13698) );
  OR2_X1 U10247 ( .A1(n12503), .A2(n13698), .ZN(n8465) );
  INV_X1 U10248 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13642) );
  OR2_X1 U10249 ( .A1(n8240), .A2(n13642), .ZN(n8464) );
  NAND4_X1 U10250 ( .A1(n8467), .A2(n8466), .A3(n8465), .A4(n8464), .ZN(n13552) );
  NAND2_X1 U10251 ( .A1(n13700), .A2(n13552), .ZN(n12612) );
  INV_X1 U10252 ( .A(n8468), .ZN(n8469) );
  XNOR2_X1 U10253 ( .A(n8470), .B(n8469), .ZN(n10700) );
  NAND2_X1 U10254 ( .A1(n10700), .A2(n12496), .ZN(n8476) );
  NAND2_X1 U10255 ( .A1(n8472), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8473) );
  MUX2_X1 U10256 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8473), .S(
        P3_IR_REG_18__SCAN_IN), .Z(n8474) );
  AND2_X1 U10257 ( .A1(n8474), .A2(n7195), .ZN(n13350) );
  AOI22_X1 U10258 ( .A1(n8490), .A2(SI_18_), .B1(n8489), .B2(n13350), .ZN(
        n8475) );
  NAND2_X1 U10259 ( .A1(n8477), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8478) );
  NAND2_X1 U10260 ( .A1(n8493), .A2(n8478), .ZN(n13526) );
  NAND2_X1 U10261 ( .A1(n8597), .A2(n13526), .ZN(n8483) );
  INV_X1 U10262 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13528) );
  OR2_X1 U10263 ( .A1(n8495), .A2(n13528), .ZN(n8482) );
  INV_X1 U10264 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13335) );
  OR2_X1 U10265 ( .A1(n8240), .A2(n13335), .ZN(n8481) );
  INV_X1 U10266 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n8479) );
  OR2_X1 U10267 ( .A1(n12503), .A2(n8479), .ZN(n8480) );
  NAND2_X1 U10268 ( .A1(n13636), .A2(n13536), .ZN(n12608) );
  INV_X1 U10269 ( .A(n8484), .ZN(n8485) );
  XNOR2_X1 U10270 ( .A(n8486), .B(n8485), .ZN(n10793) );
  NAND2_X1 U10271 ( .A1(n10793), .A2(n12496), .ZN(n8492) );
  NAND2_X1 U10272 ( .A1(n7195), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8487) );
  MUX2_X1 U10273 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8487), .S(
        P3_IR_REG_19__SCAN_IN), .Z(n8488) );
  AOI22_X1 U10274 ( .A1(n8490), .A2(SI_19_), .B1(n8489), .B2(n12686), .ZN(
        n8491) );
  NAND2_X1 U10275 ( .A1(n8493), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8494) );
  NAND2_X1 U10276 ( .A1(n8504), .A2(n8494), .ZN(n13506) );
  NAND2_X1 U10277 ( .A1(n13506), .A2(n8597), .ZN(n8499) );
  NAND2_X1 U10278 ( .A1(n8506), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8498) );
  INV_X1 U10279 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13633) );
  OR2_X1 U10280 ( .A1(n8240), .A2(n13633), .ZN(n8497) );
  INV_X1 U10281 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13508) );
  OR2_X1 U10282 ( .A1(n8495), .A2(n13508), .ZN(n8496) );
  NAND4_X1 U10283 ( .A1(n8499), .A2(n8498), .A3(n8497), .A4(n8496), .ZN(n13492) );
  NAND2_X1 U10284 ( .A1(n13514), .A2(n13525), .ZN(n12620) );
  NAND2_X1 U10285 ( .A1(n12621), .A2(n12620), .ZN(n13509) );
  INV_X1 U10286 ( .A(n13509), .ZN(n8500) );
  NAND2_X1 U10287 ( .A1(n13631), .A2(n12621), .ZN(n13486) );
  XNOR2_X1 U10288 ( .A(n8501), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n11235) );
  NAND2_X1 U10289 ( .A1(n11235), .A2(n12496), .ZN(n8503) );
  OR2_X1 U10290 ( .A1(n7158), .A2(n15191), .ZN(n8502) );
  NAND2_X1 U10291 ( .A1(n8504), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8505) );
  NAND2_X1 U10292 ( .A1(n8515), .A2(n8505), .ZN(n13497) );
  NAND2_X1 U10293 ( .A1(n13497), .A2(n8597), .ZN(n8509) );
  AOI22_X1 U10294 ( .A1(n8665), .A2(P3_REG1_REG_20__SCAN_IN), .B1(n8567), .B2(
        P3_REG2_REG_20__SCAN_IN), .ZN(n8508) );
  NAND2_X1 U10295 ( .A1(n8506), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8507) );
  XNOR2_X1 U10296 ( .A(n12999), .B(n13505), .ZN(n12674) );
  NAND2_X1 U10297 ( .A1(n13691), .A2(n13473), .ZN(n12619) );
  INV_X1 U10298 ( .A(n8510), .ZN(n8511) );
  XNOR2_X1 U10299 ( .A(n8512), .B(n8511), .ZN(n11366) );
  NAND2_X1 U10300 ( .A1(n11366), .A2(n12496), .ZN(n8514) );
  INV_X1 U10301 ( .A(SI_21_), .ZN(n11368) );
  OR2_X1 U10302 ( .A1(n7158), .A2(n11368), .ZN(n8513) );
  INV_X1 U10303 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13685) );
  NAND2_X1 U10304 ( .A1(n8515), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8516) );
  NAND2_X1 U10305 ( .A1(n8524), .A2(n8516), .ZN(n13481) );
  NAND2_X1 U10306 ( .A1(n13481), .A2(n8597), .ZN(n8518) );
  AOI22_X1 U10307 ( .A1(n8665), .A2(P3_REG1_REG_21__SCAN_IN), .B1(n8567), .B2(
        P3_REG2_REG_21__SCAN_IN), .ZN(n8517) );
  OAI211_X1 U10308 ( .C1(n12503), .C2(n13685), .A(n8518), .B(n8517), .ZN(
        n13493) );
  INV_X1 U10309 ( .A(n13493), .ZN(n13461) );
  NAND2_X1 U10310 ( .A1(n13480), .A2(n13461), .ZN(n13005) );
  INV_X1 U10311 ( .A(n8519), .ZN(n8520) );
  XNOR2_X1 U10312 ( .A(n8521), .B(n8520), .ZN(n11541) );
  NAND2_X1 U10313 ( .A1(n11541), .A2(n12496), .ZN(n8523) );
  INV_X1 U10314 ( .A(SI_22_), .ZN(n15297) );
  OR2_X1 U10315 ( .A1(n7158), .A2(n15297), .ZN(n8522) );
  NAND2_X1 U10316 ( .A1(n8524), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8525) );
  NAND2_X1 U10317 ( .A1(n8536), .A2(n8525), .ZN(n13467) );
  NAND2_X1 U10318 ( .A1(n13467), .A2(n8597), .ZN(n8530) );
  INV_X1 U10319 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13681) );
  NAND2_X1 U10320 ( .A1(n8665), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8527) );
  NAND2_X1 U10321 ( .A1(n8567), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8526) );
  OAI211_X1 U10322 ( .C1(n13681), .C2(n12503), .A(n8527), .B(n8526), .ZN(n8528) );
  INV_X1 U10323 ( .A(n8528), .ZN(n8529) );
  XNOR2_X1 U10324 ( .A(n13186), .B(n13474), .ZN(n13460) );
  NAND2_X1 U10325 ( .A1(n13458), .A2(n13460), .ZN(n8531) );
  OR2_X1 U10326 ( .A1(n13186), .A2(n13449), .ZN(n12628) );
  NAND2_X1 U10327 ( .A1(n8531), .A2(n12628), .ZN(n13451) );
  XNOR2_X1 U10328 ( .A(n8533), .B(n8532), .ZN(n11715) );
  NAND2_X1 U10329 ( .A1(n11715), .A2(n12496), .ZN(n8535) );
  INV_X1 U10330 ( .A(SI_23_), .ZN(n15294) );
  OR2_X1 U10331 ( .A1(n7158), .A2(n15294), .ZN(n8534) );
  NAND2_X1 U10332 ( .A1(n8536), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8537) );
  NAND2_X1 U10333 ( .A1(n8551), .A2(n8537), .ZN(n13453) );
  NAND2_X1 U10334 ( .A1(n13453), .A2(n8597), .ZN(n8542) );
  INV_X1 U10335 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13677) );
  NAND2_X1 U10336 ( .A1(n8665), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8539) );
  NAND2_X1 U10337 ( .A1(n8567), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8538) );
  OAI211_X1 U10338 ( .C1(n13677), .C2(n12503), .A(n8539), .B(n8538), .ZN(n8540) );
  INV_X1 U10339 ( .A(n8540), .ZN(n8541) );
  XNOR2_X1 U10340 ( .A(n13073), .B(n13462), .ZN(n13452) );
  INV_X1 U10341 ( .A(n13452), .ZN(n12675) );
  NAND2_X1 U10342 ( .A1(n13451), .A2(n12675), .ZN(n8544) );
  NAND2_X1 U10343 ( .A1(n13679), .A2(n13239), .ZN(n8543) );
  NAND2_X1 U10344 ( .A1(n8544), .A2(n8543), .ZN(n13434) );
  NAND2_X1 U10345 ( .A1(n8545), .A2(n10276), .ZN(n8546) );
  OR2_X1 U10346 ( .A1(n8547), .A2(n8546), .ZN(n8550) );
  MUX2_X1 U10347 ( .A(n7394), .B(SI_24_), .S(n10297), .Z(n8548) );
  NAND2_X1 U10348 ( .A1(n8550), .A2(n8548), .ZN(n8549) );
  OAI21_X1 U10349 ( .B1(n8550), .B2(n7394), .A(n8549), .ZN(n13036) );
  INV_X1 U10350 ( .A(n13675), .ZN(n8558) );
  NAND2_X1 U10351 ( .A1(n8551), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8552) );
  NAND2_X1 U10352 ( .A1(n8565), .A2(n8552), .ZN(n13442) );
  NAND2_X1 U10353 ( .A1(n13442), .A2(n8597), .ZN(n8557) );
  INV_X1 U10354 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13673) );
  NAND2_X1 U10355 ( .A1(n8665), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8554) );
  NAND2_X1 U10356 ( .A1(n8567), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8553) );
  OAI211_X1 U10357 ( .C1(n13673), .C2(n12503), .A(n8554), .B(n8553), .ZN(n8555) );
  INV_X1 U10358 ( .A(n8555), .ZN(n8556) );
  NAND2_X1 U10359 ( .A1(n8558), .A2(n13450), .ZN(n12528) );
  NAND2_X1 U10360 ( .A1(n13675), .A2(n13423), .ZN(n12530) );
  INV_X1 U10361 ( .A(n12530), .ZN(n8559) );
  INV_X1 U10362 ( .A(n8560), .ZN(n8561) );
  XNOR2_X1 U10363 ( .A(n8562), .B(n8561), .ZN(n12193) );
  NAND2_X1 U10364 ( .A1(n12193), .A2(n12496), .ZN(n8564) );
  INV_X1 U10365 ( .A(SI_25_), .ZN(n15174) );
  OR2_X1 U10366 ( .A1(n7158), .A2(n15174), .ZN(n8563) );
  NAND2_X1 U10367 ( .A1(n8565), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8566) );
  NAND2_X1 U10368 ( .A1(n8578), .A2(n8566), .ZN(n13429) );
  NAND2_X1 U10369 ( .A1(n13429), .A2(n8597), .ZN(n8572) );
  INV_X1 U10370 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13669) );
  NAND2_X1 U10371 ( .A1(n8665), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8569) );
  NAND2_X1 U10372 ( .A1(n8567), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8568) );
  OAI211_X1 U10373 ( .C1(n13669), .C2(n12503), .A(n8569), .B(n8568), .ZN(n8570) );
  INV_X1 U10374 ( .A(n8570), .ZN(n8571) );
  NAND2_X1 U10375 ( .A1(n13105), .A2(n13437), .ZN(n12519) );
  OR2_X1 U10376 ( .A1(n13105), .A2(n13437), .ZN(n8573) );
  INV_X1 U10377 ( .A(n13427), .ZN(n13422) );
  INV_X1 U10378 ( .A(n8574), .ZN(n8575) );
  INV_X1 U10379 ( .A(SI_26_), .ZN(n12263) );
  OR2_X1 U10380 ( .A1(n7158), .A2(n12263), .ZN(n8577) );
  NAND2_X1 U10381 ( .A1(n8578), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8579) );
  NAND2_X1 U10382 ( .A1(n8580), .A2(n8579), .ZN(n13416) );
  NAND2_X1 U10383 ( .A1(n13416), .A2(n8597), .ZN(n8585) );
  INV_X1 U10384 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13666) );
  NAND2_X1 U10385 ( .A1(n8665), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8582) );
  NAND2_X1 U10386 ( .A1(n8567), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8581) );
  OAI211_X1 U10387 ( .C1(n13666), .C2(n12503), .A(n8582), .B(n8581), .ZN(n8583) );
  INV_X1 U10388 ( .A(n8583), .ZN(n8584) );
  XNOR2_X1 U10389 ( .A(n12518), .B(n13396), .ZN(n13413) );
  INV_X1 U10390 ( .A(n12521), .ZN(n8586) );
  NAND2_X1 U10391 ( .A1(n13398), .A2(n13395), .ZN(n13394) );
  NAND2_X1 U10392 ( .A1(n13394), .A2(n12524), .ZN(n9573) );
  INV_X1 U10393 ( .A(n8587), .ZN(n8588) );
  XNOR2_X1 U10394 ( .A(n8589), .B(n8588), .ZN(n12485) );
  NAND2_X1 U10395 ( .A1(n12485), .A2(n12496), .ZN(n8591) );
  INV_X1 U10396 ( .A(SI_28_), .ZN(n15281) );
  OR2_X1 U10397 ( .A1(n7158), .A2(n15281), .ZN(n8590) );
  NAND2_X1 U10398 ( .A1(n8592), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8593) );
  NAND2_X1 U10399 ( .A1(n13371), .A2(n8593), .ZN(n13388) );
  INV_X1 U10400 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n9577) );
  NAND2_X1 U10401 ( .A1(n8665), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8595) );
  NAND2_X1 U10402 ( .A1(n8567), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8594) );
  OAI211_X1 U10403 ( .C1(n9577), .C2(n12503), .A(n8595), .B(n8594), .ZN(n8596)
         );
  OR2_X1 U10404 ( .A1(n13033), .A2(n13397), .ZN(n12640) );
  NAND2_X1 U10405 ( .A1(n13033), .A2(n13397), .ZN(n12634) );
  XOR2_X1 U10406 ( .A(n12656), .B(n12487), .Z(n13385) );
  INV_X1 U10407 ( .A(n8603), .ZN(n8599) );
  NAND2_X1 U10408 ( .A1(n8599), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8600) );
  MUX2_X1 U10409 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8600), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n8601) );
  NAND2_X1 U10410 ( .A1(n8603), .A2(n8602), .ZN(n8677) );
  INV_X1 U10411 ( .A(n8604), .ZN(n8605) );
  NAND2_X1 U10412 ( .A1(n12697), .A2(n12686), .ZN(n8662) );
  NAND2_X1 U10413 ( .A1(n8598), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8608) );
  NAND2_X1 U10414 ( .A1(n11308), .A2(n13361), .ZN(n8728) );
  NAND2_X1 U10415 ( .A1(n8662), .A2(n8728), .ZN(n8715) );
  INV_X1 U10416 ( .A(n8715), .ZN(n8609) );
  NAND2_X1 U10417 ( .A1(n8609), .A2(n12697), .ZN(n8712) );
  NAND2_X1 U10418 ( .A1(n7895), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8611) );
  NAND2_X1 U10419 ( .A1(n11367), .A2(n11308), .ZN(n8713) );
  INV_X1 U10420 ( .A(n8713), .ZN(n8612) );
  XNOR2_X1 U10421 ( .A(n8714), .B(n8612), .ZN(n8614) );
  NAND2_X1 U10422 ( .A1(n11367), .A2(n13361), .ZN(n8613) );
  NAND2_X1 U10423 ( .A1(n8614), .A2(n8613), .ZN(n11101) );
  NOR2_X1 U10424 ( .A1(n15907), .A2(n8728), .ZN(n8615) );
  NAND2_X1 U10425 ( .A1(n11101), .A2(n8615), .ZN(n8616) );
  NAND2_X1 U10426 ( .A1(n8714), .A2(n15861), .ZN(n15972) );
  NAND2_X1 U10427 ( .A1(n11316), .A2(n11326), .ZN(n8617) );
  NAND2_X1 U10428 ( .A1(n15850), .A2(n15849), .ZN(n8620) );
  NAND2_X1 U10429 ( .A1(n11334), .A2(n15845), .ZN(n8619) );
  NAND2_X1 U10430 ( .A1(n8620), .A2(n8619), .ZN(n11333) );
  NAND2_X1 U10431 ( .A1(n15847), .A2(n11846), .ZN(n8623) );
  NAND2_X1 U10432 ( .A1(n13251), .A2(n15906), .ZN(n8624) );
  NAND2_X1 U10433 ( .A1(n11724), .A2(n12021), .ZN(n8625) );
  NAND2_X1 U10434 ( .A1(n13249), .A2(n11908), .ZN(n8627) );
  NAND2_X1 U10435 ( .A1(n13248), .A2(n11994), .ZN(n8628) );
  INV_X1 U10436 ( .A(n12269), .ZN(n12569) );
  NAND2_X1 U10437 ( .A1(n12568), .A2(n12569), .ZN(n8630) );
  NAND2_X1 U10438 ( .A1(n12238), .A2(n8630), .ZN(n12253) );
  NOR2_X1 U10439 ( .A1(n13246), .A2(n12225), .ZN(n8631) );
  INV_X1 U10440 ( .A(n13246), .ZN(n12285) );
  NAND2_X1 U10441 ( .A1(n12284), .A2(n12576), .ZN(n8633) );
  NAND2_X1 U10442 ( .A1(n13245), .A2(n12422), .ZN(n8632) );
  AND2_X1 U10443 ( .A1(n13244), .A2(n13191), .ZN(n8635) );
  NAND2_X1 U10444 ( .A1(n13048), .A2(n12471), .ZN(n8634) );
  OR2_X1 U10445 ( .A1(n13193), .A2(n15971), .ZN(n13049) );
  NAND2_X1 U10446 ( .A1(n12433), .A2(n13049), .ZN(n8636) );
  NAND2_X1 U10447 ( .A1(n15971), .A2(n13193), .ZN(n13055) );
  OR2_X1 U10448 ( .A1(n12589), .A2(n13581), .ZN(n8637) );
  NAND2_X1 U10449 ( .A1(n12589), .A2(n13581), .ZN(n8638) );
  AND2_X1 U10450 ( .A1(n13567), .A2(n13549), .ZN(n8640) );
  INV_X1 U10451 ( .A(n13564), .ZN(n13228) );
  OR2_X1 U10452 ( .A1(n13706), .A2(n13228), .ZN(n13546) );
  AND2_X1 U10453 ( .A1(n8640), .A2(n13546), .ZN(n8641) );
  INV_X1 U10454 ( .A(n13535), .ZN(n13565) );
  INV_X1 U10455 ( .A(n13551), .ZN(n13579) );
  NAND2_X1 U10456 ( .A1(n13651), .A2(n13579), .ZN(n13548) );
  INV_X1 U10457 ( .A(n13552), .ZN(n13524) );
  INV_X1 U10458 ( .A(n13536), .ZN(n13241) );
  OR2_X1 U10459 ( .A1(n13636), .A2(n13241), .ZN(n8644) );
  NAND2_X1 U10460 ( .A1(n13514), .A2(n13492), .ZN(n8645) );
  NAND2_X1 U10461 ( .A1(n12999), .A2(n13473), .ZN(n8647) );
  OR2_X1 U10462 ( .A1(n13480), .A2(n13493), .ZN(n13006) );
  NAND2_X1 U10463 ( .A1(n13683), .A2(n13449), .ZN(n8648) );
  NAND2_X1 U10464 ( .A1(n13459), .A2(n8648), .ZN(n8650) );
  NAND2_X1 U10465 ( .A1(n13186), .A2(n13474), .ZN(n8649) );
  NAND2_X1 U10466 ( .A1(n8650), .A2(n8649), .ZN(n13447) );
  NAND2_X1 U10467 ( .A1(n13073), .A2(n13239), .ZN(n8651) );
  NOR2_X1 U10468 ( .A1(n13675), .A2(n13450), .ZN(n8653) );
  NAND2_X1 U10469 ( .A1(n13675), .A2(n13450), .ZN(n8654) );
  NAND2_X1 U10470 ( .A1(n13105), .A2(n13238), .ZN(n8655) );
  NAND2_X1 U10471 ( .A1(n7564), .A2(n13396), .ZN(n8656) );
  NAND2_X1 U10472 ( .A1(n13410), .A2(n8656), .ZN(n8658) );
  NAND2_X1 U10473 ( .A1(n12518), .A2(n7563), .ZN(n8657) );
  NAND2_X1 U10474 ( .A1(n13664), .A2(n13412), .ZN(n8661) );
  NAND2_X1 U10475 ( .A1(n9569), .A2(n12678), .ZN(n9568) );
  INV_X1 U10476 ( .A(n8662), .ZN(n8730) );
  INV_X1 U10477 ( .A(n11308), .ZN(n8729) );
  NOR2_X2 U10478 ( .A1(n8730), .A2(n12685), .ZN(n13578) );
  INV_X1 U10479 ( .A(n8663), .ZN(n10853) );
  NAND2_X1 U10480 ( .A1(n10853), .A2(n12695), .ZN(n10868) );
  INV_X1 U10481 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n8668) );
  NAND2_X1 U10482 ( .A1(n8665), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8667) );
  NAND2_X1 U10483 ( .A1(n8567), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8666) );
  OAI211_X1 U10484 ( .C1(n8668), .C2(n12503), .A(n8667), .B(n8666), .ZN(n8669)
         );
  INV_X1 U10485 ( .A(n8669), .ZN(n8670) );
  AND2_X1 U10486 ( .A1(n12506), .A2(n8670), .ZN(n12643) );
  INV_X1 U10487 ( .A(P3_B_REG_SCAN_IN), .ZN(n8672) );
  NAND2_X1 U10488 ( .A1(n10850), .A2(n10868), .ZN(n8671) );
  OAI21_X1 U10489 ( .B1(n8663), .B2(n8672), .A(n15846), .ZN(n13373) );
  NOR2_X1 U10490 ( .A1(n12643), .A2(n13373), .ZN(n8673) );
  NOR2_X2 U10491 ( .A1(n8677), .A2(P3_IR_REG_23__SCAN_IN), .ZN(n8680) );
  INV_X1 U10492 ( .A(n8680), .ZN(n8709) );
  NAND2_X1 U10493 ( .A1(n8683), .A2(n12194), .ZN(n8688) );
  NAND2_X1 U10494 ( .A1(n7235), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8684) );
  INV_X1 U10495 ( .A(n12262), .ZN(n8687) );
  NAND2_X1 U10496 ( .A1(n8688), .A2(n8687), .ZN(n8692) );
  NAND2_X1 U10497 ( .A1(n8690), .A2(n12262), .ZN(n8691) );
  OR2_X1 U10498 ( .A1(n8693), .A2(P3_D_REG_1__SCAN_IN), .ZN(n8695) );
  NAND2_X1 U10499 ( .A1(n12194), .A2(n12262), .ZN(n8694) );
  XNOR2_X1 U10500 ( .A(n11307), .B(n13709), .ZN(n8711) );
  NOR2_X1 U10501 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .ZN(
        n8699) );
  NOR4_X1 U10502 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n8698) );
  NOR4_X1 U10503 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n8697) );
  NOR4_X1 U10504 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8696) );
  NAND4_X1 U10505 ( .A1(n8699), .A2(n8698), .A3(n8697), .A4(n8696), .ZN(n8705)
         );
  NOR4_X1 U10506 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n8703) );
  NOR4_X1 U10507 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n8702) );
  NOR4_X1 U10508 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n8701) );
  NOR4_X1 U10509 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_8__SCAN_IN), .ZN(n8700) );
  NAND4_X1 U10510 ( .A1(n8703), .A2(n8702), .A3(n8701), .A4(n8700), .ZN(n8704)
         );
  NOR2_X1 U10511 ( .A1(n8705), .A2(n8704), .ZN(n8706) );
  NAND2_X1 U10512 ( .A1(n8604), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8707) );
  MUX2_X1 U10513 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8707), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n8708) );
  INV_X1 U10514 ( .A(n13709), .ZN(n8719) );
  NAND2_X1 U10515 ( .A1(n8712), .A2(n12635), .ZN(n11186) );
  NAND2_X1 U10516 ( .A1(n12641), .A2(n8728), .ZN(n11184) );
  AND2_X1 U10517 ( .A1(n11186), .A2(n11184), .ZN(n8718) );
  AOI22_X1 U10518 ( .A1(n8715), .A2(n11367), .B1(n8714), .B2(n8713), .ZN(n8716) );
  NAND2_X1 U10519 ( .A1(n8719), .A2(n8716), .ZN(n8717) );
  OAI21_X1 U10520 ( .B1(n8719), .B2(n8718), .A(n8717), .ZN(n8720) );
  INV_X1 U10521 ( .A(n8720), .ZN(n8721) );
  INV_X1 U10522 ( .A(n8722), .ZN(n13383) );
  INV_X1 U10523 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n8723) );
  NOR2_X1 U10524 ( .A1(n16039), .A2(n8723), .ZN(n8724) );
  INV_X1 U10525 ( .A(n11307), .ZN(n13711) );
  NAND3_X1 U10526 ( .A1(n13711), .A2(n13709), .A3(n8731), .ZN(n11106) );
  INV_X1 U10527 ( .A(n8728), .ZN(n12654) );
  NAND2_X1 U10528 ( .A1(n12641), .A2(n12654), .ZN(n11095) );
  AND2_X1 U10529 ( .A1(n11367), .A2(n8729), .ZN(n12692) );
  NAND2_X1 U10530 ( .A1(n8730), .A2(n12692), .ZN(n11102) );
  AND2_X1 U10531 ( .A1(n11095), .A2(n11102), .ZN(n8734) );
  INV_X1 U10532 ( .A(n8731), .ZN(n8732) );
  INV_X1 U10533 ( .A(n11101), .ZN(n8733) );
  OAI22_X1 U10534 ( .A1(n11106), .A2(n8734), .B1(n11111), .B2(n8733), .ZN(
        n8735) );
  NOR2_X1 U10535 ( .A1(n16042), .A2(n8736), .ZN(n8737) );
  NAND2_X1 U10536 ( .A1(n10297), .A2(SI_0_), .ZN(n8740) );
  XNOR2_X1 U10537 ( .A(n8740), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n14424) );
  NAND4_X1 U10538 ( .A1(n9012), .A2(n8743), .A3(n8742), .A4(n8741), .ZN(n9113)
         );
  INV_X1 U10539 ( .A(n9113), .ZN(n8746) );
  NAND2_X1 U10540 ( .A1(n8800), .A2(n8747), .ZN(n8850) );
  INV_X1 U10541 ( .A(n8850), .ZN(n8749) );
  INV_X1 U10542 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8750) );
  INV_X1 U10543 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8751) );
  NOR2_X1 U10544 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n8753) );
  NOR2_X1 U10545 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), 
        .ZN(n8752) );
  INV_X1 U10546 ( .A(n8758), .ZN(n8759) );
  NAND2_X1 U10547 ( .A1(n8763), .A2(n8765), .ZN(n8766) );
  MUX2_X1 U10548 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8770), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n8769) );
  NAND2_X1 U10549 ( .A1(n8769), .A2(n9525), .ZN(n12356) );
  INV_X2 U10550 ( .A(n12356), .ZN(n10183) );
  INV_X1 U10551 ( .A(n8770), .ZN(n8776) );
  INV_X1 U10552 ( .A(n8763), .ZN(n9135) );
  NAND2_X1 U10553 ( .A1(n9179), .A2(n8771), .ZN(n8772) );
  NAND2_X1 U10554 ( .A1(n8779), .A2(n8773), .ZN(n8774) );
  NAND2_X1 U10555 ( .A1(n8774), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8775) );
  MUX2_X2 U10556 ( .A(n8776), .B(n8775), .S(P2_IR_REG_20__SCAN_IN), .Z(n10264)
         );
  INV_X1 U10557 ( .A(n10264), .ZN(n8777) );
  XNOR2_X2 U10558 ( .A(n8778), .B(P2_IR_REG_22__SCAN_IN), .ZN(n9398) );
  XNOR2_X2 U10559 ( .A(n8779), .B(P2_IR_REG_19__SCAN_IN), .ZN(n12085) );
  INV_X2 U10560 ( .A(n10264), .ZN(n9563) );
  AND2_X2 U10561 ( .A1(n16024), .A2(n10183), .ZN(n8816) );
  INV_X1 U10562 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n8781) );
  NOR2_X1 U10563 ( .A1(n8794), .A2(n8781), .ZN(n8783) );
  NOR2_X1 U10564 ( .A1(n8783), .A2(n8782), .ZN(n8789) );
  INV_X1 U10565 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n8784) );
  NAND2_X1 U10566 ( .A1(n8786), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8787) );
  NAND3_X1 U10567 ( .A1(n8789), .A2(n8788), .A3(n8787), .ZN(n9548) );
  INV_X1 U10568 ( .A(n9548), .ZN(n10108) );
  AOI211_X1 U10569 ( .C1(n11250), .C2(n11242), .A(n8883), .B(n10108), .ZN(
        n8792) );
  NAND2_X1 U10570 ( .A1(n9548), .A2(n10642), .ZN(n9549) );
  BUF_X1 U10571 ( .A(n8816), .Z(n9240) );
  AOI21_X1 U10572 ( .B1(n9549), .B2(n9240), .A(n10235), .ZN(n8790) );
  AOI21_X1 U10573 ( .B1(n11250), .B2(n9484), .A(n8790), .ZN(n8791) );
  INV_X1 U10574 ( .A(n8815), .ZN(n8821) );
  NAND2_X1 U10575 ( .A1(n8793), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8798) );
  INV_X1 U10576 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10456) );
  INV_X1 U10577 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10447) );
  OR2_X1 U10578 ( .A1(n9145), .A2(n10447), .ZN(n8796) );
  INV_X1 U10579 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10545) );
  NAND2_X1 U10580 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8799) );
  MUX2_X1 U10581 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8799), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8801) );
  INV_X1 U10582 ( .A(n8800), .ZN(n8828) );
  NAND2_X1 U10583 ( .A1(n8801), .A2(n8828), .ZN(n15461) );
  INV_X1 U10584 ( .A(n15461), .ZN(n10457) );
  NAND2_X1 U10585 ( .A1(n8849), .A2(n10457), .ZN(n8813) );
  OAI21_X1 U10586 ( .B1(n8806), .B2(n8804), .A(n8803), .ZN(n8805) );
  INV_X1 U10587 ( .A(SI_0_), .ZN(n9657) );
  NAND2_X1 U10588 ( .A1(n8810), .A2(n8047), .ZN(n8811) );
  NAND2_X1 U10589 ( .A1(n8823), .A2(n8811), .ZN(n10305) );
  OAI211_X2 U10590 ( .C1(n9040), .C2(n10304), .A(n8813), .B(n8812), .ZN(n10721) );
  INV_X1 U10591 ( .A(n8820), .ZN(n8814) );
  NAND2_X1 U10592 ( .A1(n8815), .A2(n8814), .ZN(n8819) );
  BUF_X1 U10593 ( .A(n8816), .Z(n9482) );
  AOI22_X1 U10594 ( .A1(n13932), .A2(n9484), .B1(n9482), .B2(n10721), .ZN(
        n8817) );
  INV_X1 U10595 ( .A(n8817), .ZN(n8818) );
  AOI22_X1 U10596 ( .A1(n8821), .A2(n8820), .B1(n8819), .B2(n8818), .ZN(n8838)
         );
  NAND2_X1 U10597 ( .A1(n8824), .A2(SI_2_), .ZN(n8841) );
  INV_X1 U10598 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10278) );
  MUX2_X1 U10599 ( .A(n10278), .B(n10310), .S(n9648), .Z(n8825) );
  NAND2_X1 U10600 ( .A1(n8826), .A2(n8825), .ZN(n8827) );
  AND2_X1 U10601 ( .A1(n8842), .A2(n8827), .ZN(n10277) );
  NAND2_X1 U10602 ( .A1(n10277), .A2(n9467), .ZN(n8831) );
  NAND2_X1 U10603 ( .A1(n8828), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8829) );
  XNOR2_X1 U10604 ( .A(n8829), .B(P2_IR_REG_2__SCAN_IN), .ZN(n10496) );
  AOI22_X1 U10605 ( .A1(n8897), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n8849), .B2(
        n10496), .ZN(n8830) );
  AND2_X2 U10606 ( .A1(n8831), .A2(n8830), .ZN(n11374) );
  INV_X1 U10607 ( .A(n11374), .ZN(n13876) );
  NAND2_X1 U10608 ( .A1(n8793), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8835) );
  INV_X1 U10609 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10465) );
  OR2_X1 U10610 ( .A1(n8856), .A2(n10465), .ZN(n8834) );
  INV_X1 U10611 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10458) );
  OR2_X1 U10612 ( .A1(n8794), .A2(n10458), .ZN(n8832) );
  AOI22_X1 U10613 ( .A1(n9482), .A2(n13876), .B1(n13931), .B2(n9484), .ZN(
        n8837) );
  INV_X1 U10614 ( .A(n9419), .ZN(n9315) );
  OAI22_X1 U10615 ( .A1(n11374), .A2(n9315), .B1(n10241), .B2(n9362), .ZN(
        n8836) );
  NAND2_X1 U10616 ( .A1(n8838), .A2(n8837), .ZN(n8839) );
  MUX2_X1 U10617 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n9648), .Z(n8843) );
  NAND2_X1 U10618 ( .A1(n8843), .A2(SI_3_), .ZN(n8865) );
  OAI21_X1 U10619 ( .B1(n8843), .B2(SI_3_), .A(n8865), .ZN(n8846) );
  INV_X1 U10620 ( .A(n8846), .ZN(n8844) );
  INV_X1 U10621 ( .A(n8845), .ZN(n8847) );
  NAND2_X1 U10622 ( .A1(n8847), .A2(n8846), .ZN(n8848) );
  NAND2_X1 U10623 ( .A1(n10302), .A2(n9467), .ZN(n8855) );
  NAND2_X1 U10624 ( .A1(n8850), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8851) );
  MUX2_X1 U10625 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8851), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n8853) );
  AND2_X1 U10626 ( .A1(n8853), .A2(n8852), .ZN(n15473) );
  AOI22_X1 U10627 ( .A1(n8897), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n9229), .B2(
        n15473), .ZN(n8854) );
  AND2_X2 U10628 ( .A1(n8855), .A2(n8854), .ZN(n11415) );
  CLKBUF_X3 U10629 ( .A(n8793), .Z(n9453) );
  NAND2_X1 U10630 ( .A1(n9453), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8862) );
  INV_X1 U10631 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10476) );
  OR2_X1 U10632 ( .A1(n8794), .A2(n10476), .ZN(n8860) );
  OR2_X1 U10633 ( .A1(n8856), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8858) );
  INV_X1 U10634 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10499) );
  OR2_X1 U10635 ( .A1(n9145), .A2(n10499), .ZN(n8857) );
  OAI22_X1 U10636 ( .A1(n11415), .A2(n9315), .B1(n10758), .B2(n9489), .ZN(
        n8864) );
  AOI22_X1 U10637 ( .A1(n10750), .A2(n8883), .B1(n13929), .B2(n9484), .ZN(
        n8863) );
  NAND2_X1 U10638 ( .A1(n8866), .A2(n8865), .ZN(n8871) );
  INV_X1 U10639 ( .A(n8871), .ZN(n8868) );
  MUX2_X1 U10640 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n9648), .Z(n8867) );
  NAND2_X1 U10641 ( .A1(n8867), .A2(SI_4_), .ZN(n8890) );
  OAI21_X1 U10642 ( .B1(SI_4_), .B2(n8867), .A(n8890), .ZN(n8869) );
  NAND2_X1 U10643 ( .A1(n8868), .A2(n8869), .ZN(n8872) );
  INV_X1 U10644 ( .A(n8869), .ZN(n8870) );
  NAND2_X1 U10645 ( .A1(n8871), .A2(n8870), .ZN(n8891) );
  NAND2_X1 U10646 ( .A1(n10296), .A2(n9467), .ZN(n8878) );
  NAND2_X1 U10647 ( .A1(n8852), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8873) );
  MUX2_X1 U10648 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8873), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n8876) );
  INV_X1 U10649 ( .A(n8852), .ZN(n8875) );
  NAND2_X1 U10650 ( .A1(n8875), .A2(n8874), .ZN(n8899) );
  NAND2_X1 U10651 ( .A1(n8876), .A2(n8899), .ZN(n13940) );
  INV_X1 U10652 ( .A(n13940), .ZN(n13936) );
  AOI22_X1 U10653 ( .A1(n8897), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n9229), .B2(
        n13936), .ZN(n8877) );
  AND2_X2 U10654 ( .A1(n8878), .A2(n8877), .ZN(n11524) );
  NAND2_X1 U10655 ( .A1(n9453), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8882) );
  INV_X1 U10656 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11522) );
  OR2_X1 U10657 ( .A1(n8794), .A2(n11522), .ZN(n8881) );
  NAND2_X1 U10658 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n8906) );
  OAI21_X1 U10659 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n8906), .ZN(n11523) );
  OR2_X1 U10660 ( .A1(n8856), .A2(n11523), .ZN(n8880) );
  INV_X1 U10661 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10500) );
  OR2_X1 U10662 ( .A1(n9145), .A2(n10500), .ZN(n8879) );
  NAND2_X1 U10663 ( .A1(n8884), .A2(n8885), .ZN(n8889) );
  INV_X1 U10664 ( .A(n8884), .ZN(n8887) );
  INV_X1 U10665 ( .A(n8885), .ZN(n8886) );
  AOI22_X1 U10666 ( .A1(n8889), .A2(n8888), .B1(n8887), .B2(n8886), .ZN(n8915)
         );
  INV_X1 U10667 ( .A(n8915), .ZN(n8912) );
  MUX2_X1 U10668 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n9648), .Z(n8892) );
  NAND2_X1 U10669 ( .A1(n8892), .A2(SI_5_), .ZN(n8919) );
  OAI21_X1 U10670 ( .B1(SI_5_), .B2(n8892), .A(n8919), .ZN(n8893) );
  INV_X1 U10671 ( .A(n8893), .ZN(n8894) );
  NAND2_X1 U10672 ( .A1(n10308), .A2(n9467), .ZN(n8902) );
  NAND2_X1 U10673 ( .A1(n8899), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8898) );
  MUX2_X1 U10674 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8898), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n8900) );
  AND2_X1 U10675 ( .A1(n8900), .A2(n9114), .ZN(n13954) );
  AOI22_X1 U10676 ( .A1(n9468), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9229), .B2(
        n13954), .ZN(n8901) );
  NAND2_X1 U10677 ( .A1(n9474), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8911) );
  INV_X1 U10678 ( .A(n8793), .ZN(n9402) );
  INV_X1 U10679 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n8903) );
  OR2_X1 U10680 ( .A1(n9402), .A2(n8903), .ZN(n8910) );
  INV_X1 U10681 ( .A(n8906), .ZN(n8904) );
  NAND2_X1 U10682 ( .A1(n8904), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8927) );
  INV_X1 U10683 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8905) );
  NAND2_X1 U10684 ( .A1(n8906), .A2(n8905), .ZN(n8907) );
  NAND2_X1 U10685 ( .A1(n8927), .A2(n8907), .ZN(n11534) );
  OR2_X1 U10686 ( .A1(n8856), .A2(n11534), .ZN(n8909) );
  INV_X1 U10687 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10503) );
  OR2_X1 U10688 ( .A1(n9145), .A2(n10503), .ZN(n8908) );
  OAI22_X1 U10689 ( .A1(n11535), .A2(n9315), .B1(n11067), .B2(n9489), .ZN(
        n8913) );
  NAND2_X1 U10690 ( .A1(n8912), .A2(n8913), .ZN(n8918) );
  OAI22_X1 U10691 ( .A1(n11535), .A2(n9489), .B1(n11067), .B2(n9315), .ZN(
        n8917) );
  INV_X1 U10692 ( .A(n8913), .ZN(n8914) );
  MUX2_X1 U10693 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n9648), .Z(n8921) );
  NAND2_X1 U10694 ( .A1(n8921), .A2(SI_6_), .ZN(n8939) );
  OAI21_X1 U10695 ( .B1(SI_6_), .B2(n8921), .A(n8939), .ZN(n8936) );
  XNOR2_X1 U10696 ( .A(n8938), .B(n8936), .ZN(n10314) );
  NAND2_X1 U10697 ( .A1(n10314), .A2(n9467), .ZN(n8924) );
  NAND2_X1 U10698 ( .A1(n9114), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8922) );
  XNOR2_X1 U10699 ( .A(n8922), .B(P2_IR_REG_6__SCAN_IN), .ZN(n13969) );
  AOI22_X1 U10700 ( .A1(n9468), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9229), .B2(
        n13969), .ZN(n8923) );
  NAND2_X1 U10701 ( .A1(n9453), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8932) );
  INV_X1 U10702 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10481) );
  OR2_X1 U10703 ( .A1(n8794), .A2(n10481), .ZN(n8931) );
  INV_X1 U10704 ( .A(n8927), .ZN(n8925) );
  NAND2_X1 U10705 ( .A1(n8925), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8951) );
  INV_X1 U10706 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8926) );
  NAND2_X1 U10707 ( .A1(n8927), .A2(n8926), .ZN(n8928) );
  NAND2_X1 U10708 ( .A1(n8951), .A2(n8928), .ZN(n11463) );
  OR2_X1 U10709 ( .A1(n8856), .A2(n11463), .ZN(n8930) );
  INV_X1 U10710 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10506) );
  OR2_X1 U10711 ( .A1(n9145), .A2(n10506), .ZN(n8929) );
  NAND4_X1 U10712 ( .A1(n8932), .A2(n8931), .A3(n8930), .A4(n8929), .ZN(n13926) );
  AOI22_X1 U10713 ( .A1(n11218), .A2(n9240), .B1(n13926), .B2(n9362), .ZN(
        n8934) );
  INV_X1 U10714 ( .A(n11218), .ZN(n11462) );
  INV_X1 U10715 ( .A(n13926), .ZN(n11348) );
  OAI22_X1 U10716 ( .A1(n11462), .A2(n9315), .B1(n11348), .B2(n9489), .ZN(
        n8933) );
  INV_X1 U10717 ( .A(n8936), .ZN(n8937) );
  MUX2_X1 U10718 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9648), .Z(n8940) );
  NAND2_X1 U10719 ( .A1(n8940), .A2(SI_7_), .ZN(n8959) );
  OAI21_X1 U10720 ( .B1(n8940), .B2(SI_7_), .A(n8959), .ZN(n8941) );
  INV_X1 U10721 ( .A(n8941), .ZN(n8942) );
  NAND2_X1 U10722 ( .A1(n8943), .A2(n8942), .ZN(n8960) );
  OR2_X1 U10723 ( .A1(n8943), .A2(n8942), .ZN(n8944) );
  NAND2_X1 U10724 ( .A1(n8960), .A2(n8944), .ZN(n10321) );
  OR2_X1 U10725 ( .A1(n10321), .A2(n9395), .ZN(n8948) );
  INV_X1 U10726 ( .A(n9114), .ZN(n8946) );
  INV_X1 U10727 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8945) );
  NAND2_X1 U10728 ( .A1(n8946), .A2(n8945), .ZN(n9014) );
  NAND2_X1 U10729 ( .A1(n9014), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8967) );
  INV_X1 U10730 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n8966) );
  XNOR2_X1 U10731 ( .A(n8967), .B(P2_IR_REG_7__SCAN_IN), .ZN(n13984) );
  AOI22_X1 U10732 ( .A1(n9468), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n9229), .B2(
        n13984), .ZN(n8947) );
  NAND2_X1 U10733 ( .A1(n9474), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8956) );
  INV_X1 U10734 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n8949) );
  OR2_X1 U10735 ( .A1(n9402), .A2(n8949), .ZN(n8955) );
  NAND2_X1 U10736 ( .A1(n8951), .A2(n8950), .ZN(n8952) );
  NAND2_X1 U10737 ( .A1(n8972), .A2(n8952), .ZN(n11545) );
  OR2_X1 U10738 ( .A1(n8856), .A2(n11545), .ZN(n8954) );
  INV_X1 U10739 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10509) );
  OR2_X1 U10740 ( .A1(n9478), .A2(n10509), .ZN(n8953) );
  OAI22_X1 U10741 ( .A1(n11546), .A2(n9315), .B1(n11391), .B2(n9489), .ZN(
        n8957) );
  OAI22_X1 U10742 ( .A1(n11546), .A2(n9489), .B1(n11391), .B2(n9482), .ZN(
        n8958) );
  INV_X1 U10743 ( .A(n8981), .ZN(n8978) );
  MUX2_X1 U10744 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n10297), .Z(n8961) );
  NAND2_X1 U10745 ( .A1(n8961), .A2(SI_8_), .ZN(n8984) );
  OAI21_X1 U10746 ( .B1(SI_8_), .B2(n8961), .A(n8984), .ZN(n8962) );
  INV_X1 U10747 ( .A(n8962), .ZN(n8963) );
  NAND2_X1 U10748 ( .A1(n8985), .A2(n8965), .ZN(n10372) );
  OR2_X1 U10749 ( .A1(n10372), .A2(n9395), .ZN(n8970) );
  NAND2_X1 U10750 ( .A1(n8967), .A2(n8966), .ZN(n8968) );
  NAND2_X1 U10751 ( .A1(n8968), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8992) );
  XNOR2_X1 U10752 ( .A(n8992), .B(P2_IR_REG_8__SCAN_IN), .ZN(n14000) );
  AOI22_X1 U10753 ( .A1(n9468), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n9229), .B2(
        n14000), .ZN(n8969) );
  NAND2_X1 U10754 ( .A1(n9453), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8977) );
  INV_X1 U10755 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11400) );
  OR2_X1 U10756 ( .A1(n8794), .A2(n11400), .ZN(n8976) );
  NAND2_X1 U10757 ( .A1(n8972), .A2(n8971), .ZN(n8973) );
  NAND2_X1 U10758 ( .A1(n8997), .A2(n8973), .ZN(n11655) );
  OR2_X1 U10759 ( .A1(n8856), .A2(n11655), .ZN(n8975) );
  INV_X1 U10760 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10512) );
  OR2_X1 U10761 ( .A1(n9478), .A2(n10512), .ZN(n8974) );
  OAI22_X1 U10762 ( .A1(n11643), .A2(n9489), .B1(n11644), .B2(n9482), .ZN(
        n8979) );
  NAND2_X1 U10763 ( .A1(n8978), .A2(n8979), .ZN(n8983) );
  OAI22_X1 U10764 ( .A1(n11643), .A2(n9315), .B1(n11644), .B2(n9489), .ZN(
        n8982) );
  INV_X1 U10765 ( .A(n8979), .ZN(n8980) );
  MUX2_X1 U10766 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9648), .Z(n8986) );
  NAND2_X1 U10767 ( .A1(n8986), .A2(SI_9_), .ZN(n9005) );
  OAI21_X1 U10768 ( .B1(SI_9_), .B2(n8986), .A(n9005), .ZN(n8987) );
  INV_X1 U10769 ( .A(n8987), .ZN(n8988) );
  NAND2_X1 U10770 ( .A1(n9006), .A2(n8990), .ZN(n10433) );
  INV_X1 U10771 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n8991) );
  NAND2_X1 U10772 ( .A1(n8992), .A2(n8991), .ZN(n8993) );
  NAND2_X1 U10773 ( .A1(n8993), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8994) );
  XNOR2_X1 U10774 ( .A(n8994), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10530) );
  AOI22_X1 U10775 ( .A1(n10530), .A2(n9229), .B1(n8897), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n8995) );
  NAND2_X1 U10776 ( .A1(n9453), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n9002) );
  NAND2_X1 U10777 ( .A1(n8997), .A2(n8996), .ZN(n8998) );
  NAND2_X1 U10778 ( .A1(n9019), .A2(n8998), .ZN(n11749) );
  OR2_X1 U10779 ( .A1(n8856), .A2(n11749), .ZN(n9001) );
  INV_X1 U10780 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10516) );
  OR2_X1 U10781 ( .A1(n9478), .A2(n10516), .ZN(n9000) );
  INV_X1 U10782 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11595) );
  OR2_X1 U10783 ( .A1(n8794), .A2(n11595), .ZN(n8999) );
  NAND4_X1 U10784 ( .A1(n9002), .A2(n9001), .A3(n9000), .A4(n8999), .ZN(n13923) );
  AOI22_X1 U10785 ( .A1(n11742), .A2(n9362), .B1(n9482), .B2(n13923), .ZN(
        n9003) );
  INV_X1 U10786 ( .A(n11742), .ZN(n15951) );
  INV_X1 U10787 ( .A(n13923), .ZN(n11780) );
  OAI22_X1 U10788 ( .A1(n15951), .A2(n9362), .B1(n11780), .B2(n8883), .ZN(
        n9004) );
  MUX2_X1 U10789 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10297), .Z(n9007) );
  NAND2_X1 U10790 ( .A1(n9007), .A2(SI_10_), .ZN(n9030) );
  OAI21_X1 U10791 ( .B1(SI_10_), .B2(n9007), .A(n9030), .ZN(n9008) );
  INV_X1 U10792 ( .A(n9008), .ZN(n9009) );
  INV_X1 U10793 ( .A(n9012), .ZN(n9013) );
  NAND2_X1 U10794 ( .A1(n9032), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9015) );
  XNOR2_X1 U10795 ( .A(n9015), .B(P2_IR_REG_10__SCAN_IN), .ZN(n11137) );
  AOI22_X1 U10796 ( .A1(n9468), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n9229), 
        .B2(n11137), .ZN(n9016) );
  NAND2_X1 U10797 ( .A1(n9453), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n9024) );
  INV_X1 U10798 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11775) );
  OR2_X1 U10799 ( .A1(n8794), .A2(n11775), .ZN(n9023) );
  INV_X1 U10800 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9018) );
  NAND2_X1 U10801 ( .A1(n9019), .A2(n9018), .ZN(n9020) );
  NAND2_X1 U10802 ( .A1(n9044), .A2(n9020), .ZN(n11881) );
  OR2_X1 U10803 ( .A1(n8856), .A2(n11881), .ZN(n9022) );
  INV_X1 U10804 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10518) );
  OR2_X1 U10805 ( .A1(n9478), .A2(n10518), .ZN(n9021) );
  NAND4_X1 U10806 ( .A1(n9024), .A2(n9023), .A3(n9022), .A4(n9021), .ZN(n13922) );
  AOI22_X1 U10807 ( .A1(n11938), .A2(n8883), .B1(n13922), .B2(n9362), .ZN(
        n9026) );
  INV_X1 U10808 ( .A(n13922), .ZN(n11591) );
  OAI22_X1 U10809 ( .A1(n7597), .A2(n8883), .B1(n11591), .B2(n9489), .ZN(n9025) );
  OAI21_X1 U10810 ( .B1(n9027), .B2(n9026), .A(n9025), .ZN(n9029) );
  NAND2_X1 U10811 ( .A1(n9027), .A2(n9026), .ZN(n9028) );
  NAND2_X1 U10812 ( .A1(n9029), .A2(n9028), .ZN(n9053) );
  MUX2_X1 U10813 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n10297), .Z(n9059) );
  XNOR2_X1 U10814 ( .A(n9059), .B(SI_11_), .ZN(n9061) );
  INV_X1 U10815 ( .A(n9032), .ZN(n9034) );
  INV_X1 U10816 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n9033) );
  NAND2_X1 U10817 ( .A1(n9034), .A2(n9033), .ZN(n9036) );
  NAND2_X1 U10818 ( .A1(n9036), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9035) );
  MUX2_X1 U10819 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9035), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n9039) );
  INV_X1 U10820 ( .A(n9036), .ZN(n9038) );
  INV_X1 U10821 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n9037) );
  NAND2_X1 U10822 ( .A1(n9038), .A2(n9037), .ZN(n9091) );
  NAND2_X1 U10823 ( .A1(n9039), .A2(n9091), .ZN(n14015) );
  INV_X1 U10824 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10631) );
  OAI22_X1 U10825 ( .A1(n14015), .A2(n8802), .B1(n9040), .B2(n10631), .ZN(
        n9041) );
  NAND2_X1 U10826 ( .A1(n9474), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n9049) );
  INV_X1 U10827 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9042) );
  OR2_X1 U10828 ( .A1(n9402), .A2(n9042), .ZN(n9048) );
  NAND2_X1 U10829 ( .A1(n9044), .A2(n9043), .ZN(n9045) );
  NAND2_X1 U10830 ( .A1(n9067), .A2(n9045), .ZN(n11955) );
  OR2_X1 U10831 ( .A1(n8856), .A2(n11955), .ZN(n9047) );
  INV_X1 U10832 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11138) );
  OR2_X1 U10833 ( .A1(n9145), .A2(n11138), .ZN(n9046) );
  NAND2_X1 U10834 ( .A1(n9053), .A2(n9054), .ZN(n9052) );
  INV_X1 U10835 ( .A(n15965), .ZN(n11737) );
  INV_X1 U10836 ( .A(n11948), .ZN(n13921) );
  AOI22_X1 U10837 ( .A1(n11737), .A2(n8883), .B1(n13921), .B2(n9484), .ZN(
        n9050) );
  INV_X1 U10838 ( .A(n9050), .ZN(n9051) );
  NAND2_X1 U10839 ( .A1(n9052), .A2(n9051), .ZN(n9058) );
  NAND2_X1 U10840 ( .A1(n9056), .A2(n9055), .ZN(n9057) );
  NAND2_X1 U10841 ( .A1(n9058), .A2(n9057), .ZN(n9075) );
  INV_X1 U10842 ( .A(n9059), .ZN(n9060) );
  MUX2_X1 U10843 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n10297), .Z(n9083) );
  XNOR2_X1 U10844 ( .A(n9083), .B(n15172), .ZN(n9081) );
  XNOR2_X1 U10845 ( .A(n9082), .B(n9081), .ZN(n10739) );
  NAND2_X1 U10846 ( .A1(n10739), .A2(n9467), .ZN(n9065) );
  NAND2_X1 U10847 ( .A1(n9091), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9063) );
  XNOR2_X1 U10848 ( .A(n9063), .B(P2_IR_REG_12__SCAN_IN), .ZN(n15522) );
  AOI22_X1 U10849 ( .A1(n15522), .A2(n9229), .B1(n8897), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n9064) );
  AND2_X2 U10850 ( .A1(n9065), .A2(n9064), .ZN(n12203) );
  NAND2_X1 U10851 ( .A1(n8793), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9072) );
  INV_X1 U10852 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n12009) );
  OR2_X1 U10853 ( .A1(n8794), .A2(n12009), .ZN(n9071) );
  INV_X1 U10854 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9066) );
  NAND2_X1 U10855 ( .A1(n9067), .A2(n9066), .ZN(n9068) );
  NAND2_X1 U10856 ( .A1(n9096), .A2(n9068), .ZN(n12062) );
  OR2_X1 U10857 ( .A1(n8856), .A2(n12062), .ZN(n9070) );
  INV_X1 U10858 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11142) );
  OR2_X1 U10859 ( .A1(n9145), .A2(n11142), .ZN(n9069) );
  NAND2_X1 U10860 ( .A1(n9075), .A2(n9076), .ZN(n9074) );
  OAI22_X1 U10861 ( .A1(n12203), .A2(n8883), .B1(n12144), .B2(n9489), .ZN(
        n9073) );
  NAND2_X1 U10862 ( .A1(n9074), .A2(n9073), .ZN(n9080) );
  INV_X1 U10863 ( .A(n9075), .ZN(n9078) );
  INV_X1 U10864 ( .A(n9076), .ZN(n9077) );
  NAND2_X1 U10865 ( .A1(n9078), .A2(n9077), .ZN(n9079) );
  NAND2_X1 U10866 ( .A1(n9080), .A2(n9079), .ZN(n9105) );
  INV_X1 U10867 ( .A(n9083), .ZN(n9084) );
  NAND2_X1 U10868 ( .A1(n9084), .A2(n15172), .ZN(n9085) );
  MUX2_X1 U10869 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n9648), .Z(n9087) );
  OAI21_X1 U10870 ( .B1(SI_13_), .B2(n9087), .A(n9111), .ZN(n9088) );
  NAND2_X1 U10871 ( .A1(n9089), .A2(n9088), .ZN(n9090) );
  OAI21_X1 U10872 ( .B1(n9091), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9092) );
  XNOR2_X1 U10873 ( .A(n9092), .B(P2_IR_REG_13__SCAN_IN), .ZN(n15507) );
  AOI22_X1 U10874 ( .A1(n15507), .A2(n9229), .B1(n8897), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n9093) );
  NAND2_X1 U10875 ( .A1(n9453), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n9101) );
  NAND2_X1 U10876 ( .A1(n9096), .A2(n9095), .ZN(n9097) );
  NAND2_X1 U10877 ( .A1(n9119), .A2(n9097), .ZN(n12135) );
  OR2_X1 U10878 ( .A1(n12135), .A2(n8856), .ZN(n9100) );
  INV_X1 U10879 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n12136) );
  OR2_X1 U10880 ( .A1(n8794), .A2(n12136), .ZN(n9099) );
  INV_X1 U10881 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11144) );
  OR2_X1 U10882 ( .A1(n9478), .A2(n11144), .ZN(n9098) );
  OAI22_X1 U10883 ( .A1(n15997), .A2(n9315), .B1(n12216), .B2(n9489), .ZN(
        n9106) );
  NAND2_X1 U10884 ( .A1(n9105), .A2(n9106), .ZN(n9104) );
  INV_X1 U10885 ( .A(n12216), .ZN(n12351) );
  AOI22_X1 U10886 ( .A1(n12141), .A2(n9240), .B1(n12351), .B2(n9362), .ZN(
        n9102) );
  INV_X1 U10887 ( .A(n9102), .ZN(n9103) );
  NAND2_X1 U10888 ( .A1(n9104), .A2(n9103), .ZN(n9110) );
  INV_X1 U10889 ( .A(n9105), .ZN(n9108) );
  INV_X1 U10890 ( .A(n9106), .ZN(n9107) );
  NAND2_X1 U10891 ( .A1(n9108), .A2(n9107), .ZN(n9109) );
  MUX2_X1 U10892 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n10297), .Z(n9131) );
  XNOR2_X1 U10893 ( .A(n9131), .B(SI_14_), .ZN(n9129) );
  XNOR2_X1 U10894 ( .A(n9130), .B(n9129), .ZN(n10817) );
  NAND2_X1 U10895 ( .A1(n10817), .A2(n9467), .ZN(n9117) );
  OAI21_X1 U10896 ( .B1(n9114), .B2(n9113), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n9115) );
  XNOR2_X1 U10897 ( .A(n9115), .B(P2_IR_REG_14__SCAN_IN), .ZN(n14032) );
  AOI22_X1 U10898 ( .A1(n8897), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n9229), 
        .B2(n14032), .ZN(n9116) );
  NAND2_X1 U10899 ( .A1(n9119), .A2(n9118), .ZN(n9120) );
  AND2_X1 U10900 ( .A1(n9140), .A2(n9120), .ZN(n12346) );
  NAND2_X1 U10901 ( .A1(n12346), .A2(n9452), .ZN(n9126) );
  INV_X1 U10902 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n14024) );
  OR2_X1 U10903 ( .A1(n8794), .A2(n14024), .ZN(n9125) );
  INV_X1 U10904 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9121) );
  OR2_X1 U10905 ( .A1(n9402), .A2(n9121), .ZN(n9124) );
  INV_X1 U10906 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9122) );
  OR2_X1 U10907 ( .A1(n9145), .A2(n9122), .ZN(n9123) );
  OAI22_X1 U10908 ( .A1(n12348), .A2(n9489), .B1(n12334), .B2(n9315), .ZN(
        n9128) );
  AOI22_X1 U10909 ( .A1(n12279), .A2(n9362), .B1(n9482), .B2(n13919), .ZN(
        n9127) );
  INV_X1 U10910 ( .A(n9131), .ZN(n9132) );
  NAND2_X1 U10911 ( .A1(n9132), .A2(n15315), .ZN(n9133) );
  MUX2_X1 U10912 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n10297), .Z(n9156) );
  XNOR2_X1 U10913 ( .A(n9156), .B(n15313), .ZN(n9154) );
  XNOR2_X1 U10914 ( .A(n9155), .B(n9154), .ZN(n11290) );
  NAND2_X1 U10915 ( .A1(n11290), .A2(n9467), .ZN(n9137) );
  NAND2_X1 U10916 ( .A1(n9135), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9180) );
  XNOR2_X1 U10917 ( .A(n9180), .B(P2_IR_REG_15__SCAN_IN), .ZN(n11610) );
  AOI22_X1 U10918 ( .A1(n9468), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n9229), 
        .B2(n11610), .ZN(n9136) );
  AND2_X2 U10919 ( .A1(n9137), .A2(n9136), .ZN(n16020) );
  INV_X1 U10920 ( .A(n9140), .ZN(n9138) );
  INV_X1 U10921 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9139) );
  NAND2_X1 U10922 ( .A1(n9140), .A2(n9139), .ZN(n9141) );
  NAND2_X1 U10923 ( .A1(n9168), .A2(n9141), .ZN(n12414) );
  OR2_X1 U10924 ( .A1(n12414), .A2(n8856), .ZN(n9148) );
  NAND2_X1 U10925 ( .A1(n9474), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n9143) );
  NAND2_X1 U10926 ( .A1(n9453), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n9142) );
  AND2_X1 U10927 ( .A1(n9143), .A2(n9142), .ZN(n9147) );
  INV_X1 U10928 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9144) );
  OR2_X1 U10929 ( .A1(n9145), .A2(n9144), .ZN(n9146) );
  OAI22_X1 U10930 ( .A1(n16020), .A2(n8883), .B1(n12401), .B2(n9489), .ZN(
        n9151) );
  AOI22_X1 U10931 ( .A1(n12382), .A2(n9240), .B1(n14273), .B2(n9362), .ZN(
        n9149) );
  INV_X1 U10932 ( .A(n9150), .ZN(n9153) );
  INV_X1 U10933 ( .A(n9156), .ZN(n9157) );
  NAND2_X1 U10934 ( .A1(n9157), .A2(n15313), .ZN(n9158) );
  MUX2_X1 U10935 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(P1_DATAO_REG_16__SCAN_IN), 
        .S(n9648), .Z(n9160) );
  OAI21_X1 U10936 ( .B1(SI_16_), .B2(n9160), .A(n9176), .ZN(n9177) );
  INV_X1 U10937 ( .A(n9177), .ZN(n9161) );
  XNOR2_X1 U10938 ( .A(n9178), .B(n9161), .ZN(n11423) );
  NAND2_X1 U10939 ( .A1(n11423), .A2(n9467), .ZN(n9166) );
  NAND2_X1 U10940 ( .A1(n9180), .A2(n9162), .ZN(n9163) );
  NAND2_X1 U10941 ( .A1(n9163), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9164) );
  XNOR2_X1 U10942 ( .A(n9164), .B(P2_IR_REG_16__SCAN_IN), .ZN(n11674) );
  AOI22_X1 U10943 ( .A1(n9468), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n9229), 
        .B2(n11674), .ZN(n9165) );
  INV_X1 U10944 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9167) );
  NAND2_X1 U10945 ( .A1(n9168), .A2(n9167), .ZN(n9169) );
  AND2_X1 U10946 ( .A1(n9186), .A2(n9169), .ZN(n14286) );
  NAND2_X1 U10947 ( .A1(n14286), .A2(n9452), .ZN(n9172) );
  AOI22_X1 U10948 ( .A1(n9474), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n9453), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n9171) );
  NAND2_X1 U10949 ( .A1(n8786), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n9170) );
  OAI22_X1 U10950 ( .A1(n14403), .A2(n9362), .B1(n12441), .B2(n8883), .ZN(
        n9174) );
  AOI22_X1 U10951 ( .A1(n14284), .A2(n9362), .B1(n9482), .B2(n14249), .ZN(
        n9173) );
  MUX2_X1 U10952 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n9648), .Z(n9201) );
  XNOR2_X1 U10953 ( .A(n9201), .B(SI_17_), .ZN(n9199) );
  XNOR2_X1 U10954 ( .A(n9200), .B(n9199), .ZN(n11569) );
  NAND2_X1 U10955 ( .A1(n11569), .A2(n9467), .ZN(n9183) );
  NAND2_X1 U10956 ( .A1(n9180), .A2(n9179), .ZN(n9181) );
  NAND2_X1 U10957 ( .A1(n9181), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9213) );
  XNOR2_X1 U10958 ( .A(n9213), .B(P2_IR_REG_17__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U10959 ( .A1(n9468), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n9229), 
        .B2(n11693), .ZN(n9182) );
  INV_X1 U10960 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9185) );
  NAND2_X1 U10961 ( .A1(n9186), .A2(n9185), .ZN(n9187) );
  NAND2_X1 U10962 ( .A1(n9218), .A2(n9187), .ZN(n14256) );
  OR2_X1 U10963 ( .A1(n14256), .A2(n8856), .ZN(n9192) );
  INV_X1 U10964 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n11682) );
  NAND2_X1 U10965 ( .A1(n9474), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n9189) );
  NAND2_X1 U10966 ( .A1(n9453), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n9188) );
  OAI211_X1 U10967 ( .C1(n11682), .C2(n9478), .A(n9189), .B(n9188), .ZN(n9190)
         );
  INV_X1 U10968 ( .A(n9190), .ZN(n9191) );
  OAI22_X1 U10969 ( .A1(n16030), .A2(n9315), .B1(n14236), .B2(n9362), .ZN(
        n9196) );
  NAND2_X1 U10970 ( .A1(n9194), .A2(n9193), .ZN(n9198) );
  INV_X1 U10971 ( .A(n9201), .ZN(n9202) );
  NAND2_X1 U10972 ( .A1(n9202), .A2(n15301), .ZN(n9203) );
  NAND2_X1 U10973 ( .A1(n9204), .A2(n15300), .ZN(n9206) );
  MUX2_X1 U10974 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n10297), .Z(n9208) );
  INV_X1 U10975 ( .A(n9207), .ZN(n9210) );
  INV_X1 U10976 ( .A(n9208), .ZN(n9209) );
  NAND2_X1 U10977 ( .A1(n9210), .A2(n9209), .ZN(n9211) );
  NAND2_X1 U10978 ( .A1(n9213), .A2(n9212), .ZN(n9214) );
  NAND2_X1 U10979 ( .A1(n9214), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9215) );
  XNOR2_X1 U10980 ( .A(n9215), .B(P2_IR_REG_18__SCAN_IN), .ZN(n15497) );
  AOI22_X1 U10981 ( .A1(n8897), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n9229), 
        .B2(n15497), .ZN(n9216) );
  INV_X1 U10982 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9217) );
  NAND2_X1 U10983 ( .A1(n9218), .A2(n9217), .ZN(n9219) );
  NAND2_X1 U10984 ( .A1(n9233), .A2(n9219), .ZN(n14229) );
  OR2_X1 U10985 ( .A1(n14229), .A2(n8856), .ZN(n9224) );
  INV_X1 U10986 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n15490) );
  NAND2_X1 U10987 ( .A1(n9474), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9221) );
  NAND2_X1 U10988 ( .A1(n8793), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n9220) );
  OAI211_X1 U10989 ( .C1(n15490), .C2(n9478), .A(n9221), .B(n9220), .ZN(n9222)
         );
  INV_X1 U10990 ( .A(n9222), .ZN(n9223) );
  NAND2_X1 U10991 ( .A1(n9224), .A2(n9223), .ZN(n14250) );
  AOI22_X1 U10992 ( .A1(n14228), .A2(n8883), .B1(n14250), .B2(n9362), .ZN(
        n9226) );
  OAI22_X1 U10993 ( .A1(n14397), .A2(n8883), .B1(n14209), .B2(n9362), .ZN(
        n9225) );
  MUX2_X1 U10994 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n10297), .Z(n9249) );
  XNOR2_X1 U10995 ( .A(n9249), .B(SI_19_), .ZN(n9252) );
  XNOR2_X1 U10996 ( .A(n9253), .B(n9252), .ZN(n12066) );
  NAND2_X1 U10997 ( .A1(n12066), .A2(n9467), .ZN(n9231) );
  AOI22_X1 U10998 ( .A1(n8897), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9229), 
        .B2(n12085), .ZN(n9230) );
  INV_X1 U10999 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9232) );
  NAND2_X1 U11000 ( .A1(n9233), .A2(n9232), .ZN(n9234) );
  NAND2_X1 U11001 ( .A1(n9258), .A2(n9234), .ZN(n14217) );
  INV_X1 U11002 ( .A(n14217), .ZN(n13795) );
  NAND2_X1 U11003 ( .A1(n13795), .A2(n9452), .ZN(n9239) );
  INV_X1 U11004 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n14218) );
  NAND2_X1 U11005 ( .A1(n8786), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n9236) );
  NAND2_X1 U11006 ( .A1(n9453), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n9235) );
  OAI211_X1 U11007 ( .C1(n8794), .C2(n14218), .A(n9236), .B(n9235), .ZN(n9237)
         );
  INV_X1 U11008 ( .A(n9237), .ZN(n9238) );
  OAI22_X1 U11009 ( .A1(n14355), .A2(n9315), .B1(n14238), .B2(n9362), .ZN(
        n9244) );
  AOI22_X1 U11010 ( .A1(n14220), .A2(n9240), .B1(n14188), .B2(n9362), .ZN(
        n9241) );
  AOI21_X1 U11011 ( .B1(n9243), .B2(n9244), .A(n9241), .ZN(n9242) );
  INV_X1 U11012 ( .A(n9242), .ZN(n9248) );
  INV_X1 U11013 ( .A(n9243), .ZN(n9246) );
  INV_X1 U11014 ( .A(n9244), .ZN(n9245) );
  NAND2_X1 U11015 ( .A1(n9248), .A2(n9247), .ZN(n9268) );
  INV_X1 U11016 ( .A(n9249), .ZN(n9250) );
  INV_X1 U11017 ( .A(SI_19_), .ZN(n15303) );
  NAND2_X1 U11018 ( .A1(n9250), .A2(n15303), .ZN(n9251) );
  MUX2_X1 U11019 ( .A(n12273), .B(n7692), .S(n9648), .Z(n9270) );
  XNOR2_X1 U11020 ( .A(n9270), .B(SI_20_), .ZN(n9254) );
  XNOR2_X1 U11021 ( .A(n9271), .B(n9254), .ZN(n12272) );
  NAND2_X1 U11022 ( .A1(n12272), .A2(n9467), .ZN(n9256) );
  NAND2_X1 U11023 ( .A1(n9468), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9255) );
  INV_X1 U11024 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9257) );
  NAND2_X1 U11025 ( .A1(n9258), .A2(n9257), .ZN(n9259) );
  AND2_X1 U11026 ( .A1(n9275), .A2(n9259), .ZN(n14193) );
  NAND2_X1 U11027 ( .A1(n14193), .A2(n9452), .ZN(n9265) );
  INV_X1 U11028 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9262) );
  NAND2_X1 U11029 ( .A1(n9474), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n9261) );
  NAND2_X1 U11030 ( .A1(n9453), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n9260) );
  OAI211_X1 U11031 ( .C1(n9262), .C2(n9478), .A(n9261), .B(n9260), .ZN(n9263)
         );
  INV_X1 U11032 ( .A(n9263), .ZN(n9264) );
  OAI22_X1 U11033 ( .A1(n14195), .A2(n9362), .B1(n14210), .B2(n9482), .ZN(
        n9267) );
  AOI22_X1 U11034 ( .A1(n14346), .A2(n9362), .B1(n9482), .B2(n13918), .ZN(
        n9266) );
  INV_X1 U11035 ( .A(n9270), .ZN(n9269) );
  MUX2_X1 U11036 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n10297), .Z(n9287) );
  XNOR2_X1 U11037 ( .A(n9287), .B(SI_21_), .ZN(n9284) );
  XNOR2_X1 U11038 ( .A(n9286), .B(n9284), .ZN(n12354) );
  NAND2_X1 U11039 ( .A1(n12354), .A2(n9467), .ZN(n9273) );
  NAND2_X1 U11040 ( .A1(n9468), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9272) );
  INV_X1 U11041 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13820) );
  NAND2_X1 U11042 ( .A1(n9275), .A2(n13820), .ZN(n9276) );
  NAND2_X1 U11043 ( .A1(n9290), .A2(n9276), .ZN(n14180) );
  OR2_X1 U11044 ( .A1(n14180), .A2(n8856), .ZN(n9281) );
  INV_X1 U11045 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n14344) );
  NAND2_X1 U11046 ( .A1(n9453), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n9278) );
  NAND2_X1 U11047 ( .A1(n9474), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n9277) );
  OAI211_X1 U11048 ( .C1(n14344), .C2(n9478), .A(n9278), .B(n9277), .ZN(n9279)
         );
  INV_X1 U11049 ( .A(n9279), .ZN(n9280) );
  NAND2_X1 U11050 ( .A1(n9281), .A2(n9280), .ZN(n14189) );
  AOI22_X1 U11051 ( .A1(n14182), .A2(n9362), .B1(n9315), .B2(n14189), .ZN(
        n9283) );
  INV_X1 U11052 ( .A(n14189), .ZN(n13867) );
  OAI22_X1 U11053 ( .A1(n14391), .A2(n9362), .B1(n13867), .B2(n9315), .ZN(
        n9282) );
  INV_X1 U11054 ( .A(n9284), .ZN(n9285) );
  MUX2_X1 U11055 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9648), .Z(n9329) );
  XNOR2_X1 U11056 ( .A(n9581), .B(n9329), .ZN(n12461) );
  NAND2_X1 U11057 ( .A1(n12461), .A2(n9467), .ZN(n9289) );
  NAND2_X1 U11058 ( .A1(n9468), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9288) );
  INV_X1 U11059 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13869) );
  NAND2_X1 U11060 ( .A1(n9290), .A2(n13869), .ZN(n9291) );
  AND2_X1 U11061 ( .A1(n9307), .A2(n9291), .ZN(n14160) );
  INV_X1 U11062 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9294) );
  NAND2_X1 U11063 ( .A1(n9474), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U11064 ( .A1(n9453), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9292) );
  OAI211_X1 U11065 ( .C1(n9294), .C2(n9478), .A(n9293), .B(n9292), .ZN(n9295)
         );
  AOI21_X1 U11066 ( .B1(n14160), .B2(n9452), .A(n9295), .ZN(n13817) );
  OAI22_X1 U11067 ( .A1(n14162), .A2(n9362), .B1(n13817), .B2(n9482), .ZN(
        n9298) );
  INV_X1 U11068 ( .A(n13817), .ZN(n13917) );
  AOI22_X1 U11069 ( .A1(n14336), .A2(n9362), .B1(n8883), .B2(n13917), .ZN(
        n9296) );
  AOI21_X1 U11070 ( .B1(n9299), .B2(n9298), .A(n9296), .ZN(n9297) );
  INV_X1 U11071 ( .A(n9297), .ZN(n9300) );
  NAND2_X1 U11072 ( .A1(n9300), .A2(n7207), .ZN(n9319) );
  INV_X1 U11073 ( .A(n9329), .ZN(n9301) );
  NAND2_X1 U11074 ( .A1(n9328), .A2(SI_22_), .ZN(n9302) );
  MUX2_X1 U11075 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n10297), .Z(n9330) );
  XNOR2_X1 U11076 ( .A(n9330), .B(SI_23_), .ZN(n9304) );
  NAND2_X1 U11077 ( .A1(n9468), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n9306) );
  INV_X1 U11078 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13789) );
  NAND2_X1 U11079 ( .A1(n9307), .A2(n13789), .ZN(n9308) );
  NAND2_X1 U11080 ( .A1(n9339), .A2(n9308), .ZN(n14147) );
  OR2_X1 U11081 ( .A1(n14147), .A2(n8856), .ZN(n9314) );
  INV_X1 U11082 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9311) );
  NAND2_X1 U11083 ( .A1(n9474), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n9310) );
  NAND2_X1 U11084 ( .A1(n9453), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n9309) );
  OAI211_X1 U11085 ( .C1(n9311), .C2(n9478), .A(n9310), .B(n9309), .ZN(n9312)
         );
  INV_X1 U11086 ( .A(n9312), .ZN(n9313) );
  OAI22_X1 U11087 ( .A1(n14149), .A2(n9315), .B1(n13868), .B2(n9362), .ZN(
        n9320) );
  NAND2_X1 U11088 ( .A1(n9319), .A2(n9320), .ZN(n9318) );
  AOI22_X1 U11089 ( .A1(n14331), .A2(n8883), .B1(n13916), .B2(n9362), .ZN(
        n9316) );
  INV_X1 U11090 ( .A(n9316), .ZN(n9317) );
  NAND2_X1 U11091 ( .A1(n9318), .A2(n9317), .ZN(n9324) );
  INV_X1 U11092 ( .A(n9319), .ZN(n9322) );
  INV_X1 U11093 ( .A(n9320), .ZN(n9321) );
  NAND2_X1 U11094 ( .A1(n9322), .A2(n9321), .ZN(n9323) );
  NAND2_X1 U11095 ( .A1(n9324), .A2(n9323), .ZN(n9365) );
  INV_X1 U11096 ( .A(n9330), .ZN(n9325) );
  NAND2_X1 U11097 ( .A1(n9325), .A2(n15294), .ZN(n9331) );
  OAI21_X1 U11098 ( .B1(n9329), .B2(SI_22_), .A(n9331), .ZN(n9326) );
  INV_X1 U11099 ( .A(n9326), .ZN(n9327) );
  NOR2_X1 U11100 ( .A1(n9301), .A2(n15297), .ZN(n9332) );
  AOI22_X1 U11101 ( .A1(n9332), .A2(n9331), .B1(n9330), .B2(SI_23_), .ZN(n9333) );
  MUX2_X1 U11102 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9648), .Z(n9347) );
  INV_X1 U11103 ( .A(SI_24_), .ZN(n15185) );
  XNOR2_X1 U11104 ( .A(n9347), .B(n15185), .ZN(n9345) );
  INV_X1 U11105 ( .A(n9345), .ZN(n9335) );
  XNOR2_X1 U11106 ( .A(n9346), .B(n9335), .ZN(n12457) );
  NAND2_X1 U11107 ( .A1(n12457), .A2(n9467), .ZN(n9337) );
  NAND2_X1 U11108 ( .A1(n8897), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9336) );
  INV_X1 U11109 ( .A(n9339), .ZN(n9338) );
  INV_X1 U11110 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13847) );
  NAND2_X1 U11111 ( .A1(n9339), .A2(n13847), .ZN(n9340) );
  AND2_X1 U11112 ( .A1(n9355), .A2(n9340), .ZN(n14132) );
  INV_X1 U11113 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9343) );
  NAND2_X1 U11114 ( .A1(n9474), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9342) );
  NAND2_X1 U11115 ( .A1(n9453), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9341) );
  OAI211_X1 U11116 ( .C1(n9343), .C2(n9478), .A(n9342), .B(n9341), .ZN(n9344)
         );
  AOI21_X1 U11117 ( .B1(n14132), .B2(n9452), .A(n9344), .ZN(n13828) );
  OAI22_X1 U11118 ( .A1(n14134), .A2(n9362), .B1(n13828), .B2(n8883), .ZN(
        n9364) );
  NAND2_X1 U11119 ( .A1(n9347), .A2(SI_24_), .ZN(n9348) );
  MUX2_X1 U11120 ( .A(n7369), .B(n12481), .S(n10297), .Z(n9350) );
  NAND2_X1 U11121 ( .A1(n9350), .A2(n15174), .ZN(n9368) );
  INV_X1 U11122 ( .A(n9350), .ZN(n9351) );
  NAND2_X1 U11123 ( .A1(n9351), .A2(SI_25_), .ZN(n9352) );
  NAND2_X1 U11124 ( .A1(n9368), .A2(n9352), .ZN(n9366) );
  XNOR2_X1 U11125 ( .A(n9367), .B(n9366), .ZN(n12479) );
  NAND2_X1 U11126 ( .A1(n12479), .A2(n9467), .ZN(n9354) );
  NAND2_X1 U11127 ( .A1(n9468), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9353) );
  INV_X1 U11128 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13830) );
  NAND2_X1 U11129 ( .A1(n9355), .A2(n13830), .ZN(n9356) );
  NAND2_X1 U11130 ( .A1(n14120), .A2(n9452), .ZN(n9361) );
  INV_X1 U11131 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n14323) );
  NAND2_X1 U11132 ( .A1(n9453), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9358) );
  NAND2_X1 U11133 ( .A1(n9474), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9357) );
  OAI211_X1 U11134 ( .C1(n9478), .C2(n14323), .A(n9358), .B(n9357), .ZN(n9359)
         );
  INV_X1 U11135 ( .A(n9359), .ZN(n9360) );
  AOI22_X1 U11136 ( .A1(n14119), .A2(n9362), .B1(n9482), .B2(n13914), .ZN(
        n9488) );
  OAI22_X1 U11137 ( .A1(n14384), .A2(n9362), .B1(n13898), .B2(n9482), .ZN(
        n9487) );
  INV_X1 U11138 ( .A(n13828), .ZN(n13915) );
  AOI22_X1 U11139 ( .A1(n14326), .A2(n9362), .B1(n9240), .B2(n13915), .ZN(
        n9363) );
  MUX2_X1 U11140 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n9648), .Z(n9465) );
  MUX2_X1 U11141 ( .A(n15434), .B(n14413), .S(n10297), .Z(n9371) );
  NAND2_X1 U11142 ( .A1(n9371), .A2(n15289), .ZN(n9372) );
  OAI21_X1 U11143 ( .B1(n9465), .B2(SI_26_), .A(n9372), .ZN(n9369) );
  INV_X1 U11144 ( .A(n9465), .ZN(n9370) );
  NOR2_X1 U11145 ( .A1(n9370), .A2(n12263), .ZN(n9373) );
  INV_X1 U11146 ( .A(n9371), .ZN(n9444) );
  AOI22_X1 U11147 ( .A1(n9373), .A2(n9372), .B1(n9444), .B2(SI_27_), .ZN(n9374) );
  MUX2_X1 U11148 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n9648), .Z(n9376) );
  XNOR2_X1 U11149 ( .A(n9376), .B(SI_28_), .ZN(n9424) );
  MUX2_X1 U11150 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n10297), .Z(n9377) );
  XNOR2_X1 U11151 ( .A(n9377), .B(n13724), .ZN(n9411) );
  NAND2_X1 U11152 ( .A1(n9410), .A2(n9411), .ZN(n9380) );
  INV_X1 U11153 ( .A(n9377), .ZN(n9378) );
  NAND2_X1 U11154 ( .A1(n9378), .A2(n13724), .ZN(n9379) );
  NAND2_X1 U11155 ( .A1(n9380), .A2(n9379), .ZN(n9392) );
  MUX2_X1 U11156 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n10297), .Z(n9381) );
  NAND2_X1 U11157 ( .A1(n9381), .A2(SI_30_), .ZN(n9382) );
  OAI21_X1 U11158 ( .B1(SI_30_), .B2(n9381), .A(n9382), .ZN(n9391) );
  MUX2_X1 U11159 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10297), .Z(n9383) );
  XNOR2_X1 U11160 ( .A(n9383), .B(SI_31_), .ZN(n9384) );
  NAND2_X1 U11161 ( .A1(n12861), .A2(n9467), .ZN(n9387) );
  NAND2_X1 U11162 ( .A1(n9468), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n9386) );
  INV_X1 U11163 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9390) );
  NAND2_X1 U11164 ( .A1(n9474), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9389) );
  NAND2_X1 U11165 ( .A1(n9453), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9388) );
  OAI211_X1 U11166 ( .C1(n9478), .C2(n9390), .A(n9389), .B(n9388), .ZN(n14046)
         );
  XNOR2_X1 U11167 ( .A(n14295), .B(n14046), .ZN(n9499) );
  NAND2_X1 U11168 ( .A1(n9392), .A2(n9391), .ZN(n9393) );
  OR2_X1 U11169 ( .A1(n15427), .A2(n9395), .ZN(n9397) );
  NAND2_X1 U11170 ( .A1(n9468), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n9396) );
  NAND2_X1 U11171 ( .A1(n9398), .A2(n12085), .ZN(n10185) );
  INV_X1 U11172 ( .A(n10185), .ZN(n9399) );
  NAND2_X1 U11173 ( .A1(n9563), .A2(n14076), .ZN(n10210) );
  AOI21_X1 U11174 ( .B1(n9563), .B2(n9399), .A(n7290), .ZN(n9406) );
  NAND2_X1 U11175 ( .A1(n14046), .A2(n9362), .ZN(n9490) );
  INV_X1 U11176 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9400) );
  OR2_X1 U11177 ( .A1(n9478), .A2(n9400), .ZN(n9405) );
  INV_X1 U11178 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n14052) );
  OR2_X1 U11179 ( .A1(n8794), .A2(n14052), .ZN(n9404) );
  INV_X1 U11180 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9401) );
  OR2_X1 U11181 ( .A1(n9402), .A2(n9401), .ZN(n9403) );
  AND3_X1 U11182 ( .A1(n9405), .A2(n9404), .A3(n9403), .ZN(n10189) );
  AOI21_X1 U11183 ( .B1(n9406), .B2(n9490), .A(n10189), .ZN(n9407) );
  AOI21_X1 U11184 ( .B1(n14299), .B2(n9240), .A(n9407), .ZN(n9498) );
  NAND2_X1 U11185 ( .A1(n14299), .A2(n9362), .ZN(n9409) );
  INV_X1 U11186 ( .A(n10189), .ZN(n13909) );
  NAND2_X1 U11187 ( .A1(n13909), .A2(n9482), .ZN(n9408) );
  NAND2_X1 U11188 ( .A1(n9409), .A2(n9408), .ZN(n9497) );
  XNOR2_X1 U11189 ( .A(n9410), .B(n9411), .ZN(n12956) );
  NAND2_X1 U11190 ( .A1(n12956), .A2(n9467), .ZN(n9413) );
  NAND2_X1 U11191 ( .A1(n9468), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n9412) );
  INV_X1 U11192 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n13901) );
  NAND2_X1 U11193 ( .A1(n9428), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n14058) );
  OR2_X1 U11194 ( .A1(n14058), .A2(n8856), .ZN(n9418) );
  INV_X1 U11195 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n10217) );
  NAND2_X1 U11196 ( .A1(n9474), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9415) );
  NAND2_X1 U11197 ( .A1(n9453), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9414) );
  OAI211_X1 U11198 ( .C1(n10217), .C2(n9478), .A(n9415), .B(n9414), .ZN(n9416)
         );
  INV_X1 U11199 ( .A(n9416), .ZN(n9417) );
  NAND2_X1 U11200 ( .A1(n9418), .A2(n9417), .ZN(n13910) );
  AND2_X1 U11201 ( .A1(n13910), .A2(n9419), .ZN(n9420) );
  AOI21_X1 U11202 ( .B1(n14060), .B2(n8883), .A(n9420), .ZN(n9501) );
  NAND2_X1 U11203 ( .A1(n14060), .A2(n9362), .ZN(n9422) );
  NAND2_X1 U11204 ( .A1(n13910), .A2(n8883), .ZN(n9421) );
  NAND2_X1 U11205 ( .A1(n9422), .A2(n9421), .ZN(n9500) );
  OAI22_X1 U11206 ( .A1(n9498), .A2(n9497), .B1(n9501), .B2(n9500), .ZN(n9423)
         );
  NAND2_X1 U11207 ( .A1(n9499), .A2(n9423), .ZN(n9506) );
  NAND2_X1 U11208 ( .A1(n15428), .A2(n9467), .ZN(n9427) );
  NAND2_X1 U11209 ( .A1(n8897), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9426) );
  INV_X1 U11210 ( .A(n9428), .ZN(n9451) );
  INV_X1 U11211 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9429) );
  NAND2_X1 U11212 ( .A1(n9451), .A2(n9429), .ZN(n9430) );
  NAND2_X1 U11213 ( .A1(n14058), .A2(n9430), .ZN(n14069) );
  INV_X1 U11214 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9433) );
  NAND2_X1 U11215 ( .A1(n9474), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9432) );
  NAND2_X1 U11216 ( .A1(n9453), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9431) );
  OAI211_X1 U11217 ( .C1(n9433), .C2(n9478), .A(n9432), .B(n9431), .ZN(n9434)
         );
  INV_X1 U11218 ( .A(n9434), .ZN(n9435) );
  AND2_X1 U11219 ( .A1(n13911), .A2(n9482), .ZN(n9437) );
  AOI21_X1 U11220 ( .B1(n14305), .B2(n9362), .A(n9437), .ZN(n9503) );
  NAND2_X1 U11221 ( .A1(n14305), .A2(n9315), .ZN(n9439) );
  NAND2_X1 U11222 ( .A1(n13911), .A2(n9362), .ZN(n9438) );
  NAND2_X1 U11223 ( .A1(n9439), .A2(n9438), .ZN(n9502) );
  NAND2_X1 U11224 ( .A1(n9503), .A2(n9502), .ZN(n9440) );
  NAND2_X1 U11225 ( .A1(n9506), .A2(n9440), .ZN(n9513) );
  XNOR2_X1 U11226 ( .A(n9441), .B(SI_26_), .ZN(n9464) );
  NAND2_X1 U11227 ( .A1(n9464), .A2(n9465), .ZN(n9443) );
  OR2_X1 U11228 ( .A1(n9441), .A2(n12263), .ZN(n9442) );
  XNOR2_X1 U11229 ( .A(n9444), .B(SI_27_), .ZN(n9445) );
  NAND2_X1 U11230 ( .A1(n14410), .A2(n9467), .ZN(n9448) );
  NAND2_X1 U11231 ( .A1(n9468), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9447) );
  INV_X1 U11232 ( .A(n9449), .ZN(n9473) );
  INV_X1 U11233 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13779) );
  NAND2_X1 U11234 ( .A1(n9473), .A2(n13779), .ZN(n9450) );
  NAND2_X1 U11235 ( .A1(n14090), .A2(n9452), .ZN(n9459) );
  INV_X1 U11236 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9456) );
  NAND2_X1 U11237 ( .A1(n9474), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9455) );
  NAND2_X1 U11238 ( .A1(n9453), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9454) );
  OAI211_X1 U11239 ( .C1(n9456), .C2(n9478), .A(n9455), .B(n9454), .ZN(n9457)
         );
  INV_X1 U11240 ( .A(n9457), .ZN(n9458) );
  AND2_X1 U11241 ( .A1(n13912), .A2(n9482), .ZN(n9460) );
  AOI21_X1 U11242 ( .B1(n14309), .B2(n9362), .A(n9460), .ZN(n9512) );
  NAND2_X1 U11243 ( .A1(n14309), .A2(n8883), .ZN(n9462) );
  NAND2_X1 U11244 ( .A1(n13912), .A2(n9362), .ZN(n9461) );
  NAND2_X1 U11245 ( .A1(n9462), .A2(n9461), .ZN(n9511) );
  AND2_X1 U11246 ( .A1(n9512), .A2(n9511), .ZN(n9463) );
  NOR2_X1 U11247 ( .A1(n9513), .A2(n9463), .ZN(n9516) );
  INV_X1 U11248 ( .A(n9464), .ZN(n9466) );
  NAND2_X1 U11249 ( .A1(n14414), .A2(n9467), .ZN(n9470) );
  NAND2_X1 U11250 ( .A1(n9468), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9469) );
  NAND2_X2 U11251 ( .A1(n9470), .A2(n9469), .ZN(n14314) );
  NAND2_X1 U11252 ( .A1(n9471), .A2(n13901), .ZN(n9472) );
  NAND2_X1 U11253 ( .A1(n9473), .A2(n9472), .ZN(n14103) );
  OR2_X1 U11254 ( .A1(n14103), .A2(n8856), .ZN(n9481) );
  INV_X1 U11255 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9477) );
  NAND2_X1 U11256 ( .A1(n9453), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n9476) );
  NAND2_X1 U11257 ( .A1(n9474), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n9475) );
  OAI211_X1 U11258 ( .C1(n9478), .C2(n9477), .A(n9476), .B(n9475), .ZN(n9479)
         );
  INV_X1 U11259 ( .A(n9479), .ZN(n9480) );
  NAND2_X1 U11260 ( .A1(n9481), .A2(n9480), .ZN(n13913) );
  AND2_X1 U11261 ( .A1(n13913), .A2(n9482), .ZN(n9483) );
  AOI21_X1 U11262 ( .B1(n14314), .B2(n9484), .A(n9483), .ZN(n9496) );
  NAND2_X1 U11263 ( .A1(n14314), .A2(n8883), .ZN(n9486) );
  NAND2_X1 U11264 ( .A1(n13913), .A2(n9362), .ZN(n9485) );
  NAND2_X1 U11265 ( .A1(n9486), .A2(n9485), .ZN(n9495) );
  AOI22_X1 U11266 ( .A1(n9496), .A2(n9495), .B1(n9488), .B2(n9487), .ZN(n9493)
         );
  NAND2_X1 U11267 ( .A1(n14046), .A2(n9315), .ZN(n9492) );
  NAND2_X1 U11268 ( .A1(n9490), .A2(n9489), .ZN(n9491) );
  MUX2_X1 U11269 ( .A(n9492), .B(n9491), .S(n14295), .Z(n9518) );
  AND3_X1 U11270 ( .A1(n9516), .A2(n9493), .A3(n9518), .ZN(n9494) );
  NOR2_X1 U11271 ( .A1(n9496), .A2(n9495), .ZN(n9517) );
  INV_X1 U11272 ( .A(n9497), .ZN(n9510) );
  INV_X1 U11273 ( .A(n9498), .ZN(n9509) );
  INV_X1 U11274 ( .A(n9499), .ZN(n9560) );
  INV_X1 U11275 ( .A(n9500), .ZN(n9505) );
  INV_X1 U11276 ( .A(n9501), .ZN(n9504) );
  OAI22_X1 U11277 ( .A1(n9505), .A2(n9504), .B1(n9503), .B2(n9502), .ZN(n9507)
         );
  OAI21_X1 U11278 ( .B1(n9560), .B2(n9507), .A(n9506), .ZN(n9508) );
  OAI21_X1 U11279 ( .B1(n9510), .B2(n9509), .A(n9508), .ZN(n9515) );
  NOR3_X1 U11280 ( .A1(n9513), .A2(n9512), .A3(n9511), .ZN(n9514) );
  AOI211_X1 U11281 ( .C1(n9517), .C2(n9516), .A(n9515), .B(n9514), .ZN(n9520)
         );
  INV_X1 U11282 ( .A(n9518), .ZN(n9519) );
  NAND2_X1 U11283 ( .A1(n10183), .A2(n14076), .ZN(n9522) );
  OAI211_X1 U11284 ( .C1(n10235), .C2(n9398), .A(n10210), .B(n9522), .ZN(n9523) );
  INV_X1 U11285 ( .A(n9523), .ZN(n9524) );
  NAND2_X1 U11286 ( .A1(n9534), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9527) );
  INV_X1 U11287 ( .A(n10438), .ZN(n9528) );
  AND2_X1 U11288 ( .A1(n9528), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9533) );
  MUX2_X1 U11289 ( .A(n12356), .B(n9530), .S(n9563), .Z(n9531) );
  NOR2_X1 U11290 ( .A1(n9531), .A2(n14076), .ZN(n9532) );
  INV_X1 U11291 ( .A(n9533), .ZN(n14420) );
  INV_X1 U11292 ( .A(n10443), .ZN(n10444) );
  INV_X1 U11293 ( .A(n14411), .ZN(n10445) );
  NAND2_X1 U11294 ( .A1(n9536), .A2(n9535), .ZN(n9537) );
  INV_X1 U11295 ( .A(n10233), .ZN(n10261) );
  AND2_X1 U11296 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10261), .ZN(n9544) );
  INV_X1 U11297 ( .A(n10210), .ZN(n10267) );
  NAND4_X1 U11298 ( .A1(n14274), .A2(n10445), .A3(n15455), .A4(n10267), .ZN(
        n9545) );
  OAI211_X1 U11299 ( .C1(n9398), .C2(n14420), .A(n9545), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9565) );
  XNOR2_X1 U11300 ( .A(n14299), .B(n13909), .ZN(n9559) );
  NAND2_X1 U11301 ( .A1(n14305), .A2(n13778), .ZN(n9546) );
  XNOR2_X1 U11302 ( .A(n14336), .B(n13817), .ZN(n14164) );
  XNOR2_X1 U11303 ( .A(n14119), .B(n13898), .ZN(n14116) );
  XNOR2_X1 U11304 ( .A(n14326), .B(n13915), .ZN(n14127) );
  XNOR2_X1 U11305 ( .A(n14220), .B(n14238), .ZN(n14206) );
  XNOR2_X1 U11306 ( .A(n14228), .B(n14209), .ZN(n14233) );
  INV_X1 U11307 ( .A(n16030), .ZN(n14259) );
  XNOR2_X1 U11308 ( .A(n14259), .B(n14236), .ZN(n14247) );
  XNOR2_X1 U11309 ( .A(n14284), .B(n14249), .ZN(n14270) );
  XNOR2_X1 U11310 ( .A(n12141), .B(n12216), .ZN(n12142) );
  NAND2_X1 U11311 ( .A1(n12200), .A2(n12144), .ZN(n9547) );
  NAND2_X1 U11312 ( .A1(n10159), .A2(n9547), .ZN(n12012) );
  XNOR2_X1 U11313 ( .A(n11737), .B(n11948), .ZN(n11730) );
  XNOR2_X1 U11314 ( .A(n11938), .B(n13922), .ZN(n10157) );
  XNOR2_X1 U11315 ( .A(n11387), .B(n11391), .ZN(n11346) );
  XNOR2_X1 U11316 ( .A(n11218), .B(n11348), .ZN(n11214) );
  INV_X1 U11317 ( .A(n11535), .ZN(n10969) );
  INV_X1 U11318 ( .A(n11067), .ZN(n13927) );
  XNOR2_X1 U11319 ( .A(n10969), .B(n13927), .ZN(n10146) );
  INV_X1 U11320 ( .A(n10721), .ZN(n11503) );
  NAND2_X1 U11321 ( .A1(n10718), .A2(n9549), .ZN(n11243) );
  NOR4_X1 U11322 ( .A1(n10703), .A2(n10717), .A3(n11243), .A4(n9563), .ZN(
        n9550) );
  INV_X1 U11323 ( .A(n11524), .ZN(n10755) );
  NAND4_X1 U11324 ( .A1(n10146), .A2(n9550), .A3(n10756), .A4(n10142), .ZN(
        n9551) );
  NOR3_X1 U11325 ( .A1(n11346), .A2(n11214), .A3(n9551), .ZN(n9552) );
  XNOR2_X1 U11326 ( .A(n11742), .B(n13923), .ZN(n10154) );
  XNOR2_X1 U11327 ( .A(n11657), .B(n13924), .ZN(n11402) );
  NAND4_X1 U11328 ( .A1(n10157), .A2(n9552), .A3(n10154), .A4(n11402), .ZN(
        n9553) );
  NOR4_X1 U11329 ( .A1(n12142), .A2(n12012), .A3(n11730), .A4(n9553), .ZN(
        n9554) );
  XNOR2_X1 U11330 ( .A(n12382), .B(n14273), .ZN(n12372) );
  XNOR2_X1 U11331 ( .A(n12279), .B(n13919), .ZN(n12217) );
  NAND4_X1 U11332 ( .A1(n14270), .A2(n9554), .A3(n12372), .A4(n12217), .ZN(
        n9555) );
  NOR4_X1 U11333 ( .A1(n14206), .A2(n14233), .A3(n14247), .A4(n9555), .ZN(
        n9556) );
  XNOR2_X1 U11334 ( .A(n14182), .B(n14189), .ZN(n14175) );
  XNOR2_X1 U11335 ( .A(n14346), .B(n13918), .ZN(n14197) );
  NAND4_X1 U11336 ( .A1(n14127), .A2(n9556), .A3(n14175), .A4(n14197), .ZN(
        n9557) );
  NOR4_X1 U11337 ( .A1(n14078), .A2(n14164), .A3(n14116), .A4(n9557), .ZN(
        n9558) );
  XNOR2_X1 U11338 ( .A(n14060), .B(n13910), .ZN(n10180) );
  INV_X1 U11339 ( .A(n13912), .ZN(n10178) );
  XNOR2_X1 U11340 ( .A(n14309), .B(n10178), .ZN(n14086) );
  XNOR2_X1 U11341 ( .A(n14314), .B(n13829), .ZN(n14097) );
  XNOR2_X1 U11342 ( .A(n9561), .B(n12085), .ZN(n9562) );
  OAI211_X1 U11343 ( .C1(n9567), .C2(n9566), .A(n9565), .B(n7729), .ZN(
        P2_U3328) );
  OAI22_X1 U11344 ( .A1(n13031), .A2(n13580), .B1(n13412), .B2(n13582), .ZN(
        n9570) );
  INV_X1 U11345 ( .A(n9570), .ZN(n9571) );
  NAND2_X1 U11346 ( .A1(n9575), .A2(n9574), .ZN(n13391) );
  NAND2_X1 U11347 ( .A1(n13391), .A2(n13658), .ZN(n9576) );
  NAND2_X1 U11348 ( .A1(n13393), .A2(n9576), .ZN(n13595) );
  INV_X1 U11349 ( .A(n13595), .ZN(n9580) );
  NOR3_X1 U11350 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), 
        .A3(P1_IR_REG_24__SCAN_IN), .ZN(n9586) );
  NAND2_X1 U11351 ( .A1(n10061), .A2(n9586), .ZN(n9601) );
  NAND2_X1 U11352 ( .A1(n9596), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n9587) );
  NOR2_X1 U11353 ( .A1(n9601), .A2(n9587), .ZN(n9604) );
  XNOR2_X1 U11354 ( .A(n9597), .B(P1_IR_REG_31__SCAN_IN), .ZN(n9603) );
  NOR2_X1 U11355 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n9593) );
  NOR2_X1 U11356 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), 
        .ZN(n9592) );
  NOR2_X1 U11357 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), 
        .ZN(n9591) );
  AND2_X1 U11358 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n9595) );
  NAND3_X1 U11359 ( .A1(n9599), .A2(n9996), .A3(n9598), .ZN(n9600) );
  NOR2_X2 U11360 ( .A1(n9601), .A2(n9600), .ZN(n9602) );
  NAND2_X1 U11361 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9692) );
  NOR2_X1 U11362 ( .A1(n9692), .A2(n9691), .ZN(n9690) );
  NAND2_X1 U11363 ( .A1(n9690), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9718) );
  NAND2_X1 U11364 ( .A1(n9746), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9775) );
  NAND2_X1 U11365 ( .A1(n9787), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9819) );
  INV_X1 U11366 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9885) );
  INV_X1 U11367 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14658) );
  OR2_X1 U11368 ( .A1(n9911), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9606) );
  NAND2_X1 U11369 ( .A1(n9911), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9922) );
  AND2_X1 U11370 ( .A1(n9606), .A2(n9922), .ZN(n14936) );
  INV_X1 U11371 ( .A(n12957), .ZN(n9611) );
  NAND2_X1 U11372 ( .A1(n14936), .A2(n9899), .ZN(n9618) );
  INV_X1 U11373 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9615) );
  NAND2_X1 U11374 ( .A1(n10336), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n9614) );
  NAND2_X1 U11375 ( .A1(n10335), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9613) );
  OAI211_X1 U11376 ( .C1(n10057), .C2(n9615), .A(n9614), .B(n9613), .ZN(n9616)
         );
  INV_X1 U11377 ( .A(n9616), .ZN(n9617) );
  XNOR2_X1 U11378 ( .A(n15108), .B(n14608), .ZN(n14934) );
  NAND2_X1 U11379 ( .A1(n10336), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9625) );
  INV_X1 U11380 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9619) );
  OR2_X1 U11381 ( .A1(n9620), .A2(n9619), .ZN(n9624) );
  INV_X1 U11382 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9621) );
  OR2_X1 U11383 ( .A1(n9679), .A2(n9621), .ZN(n9623) );
  INV_X1 U11384 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10651) );
  OR2_X1 U11385 ( .A1(n9653), .A2(n10651), .ZN(n9622) );
  AND2_X4 U11386 ( .A1(n10323), .A2(n10276), .ZN(n12860) );
  NAND2_X1 U11387 ( .A1(n10277), .A2(n12860), .ZN(n9631) );
  AND2_X4 U11388 ( .A1(n10323), .A2(n10297), .ZN(n9893) );
  INV_X1 U11389 ( .A(n9626), .ZN(n9642) );
  NAND2_X1 U11390 ( .A1(n9642), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9627) );
  MUX2_X1 U11391 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9627), .S(
        P1_IR_REG_2__SCAN_IN), .Z(n9629) );
  INV_X1 U11392 ( .A(n9628), .ZN(n9661) );
  NAND2_X1 U11393 ( .A1(n9629), .A2(n9661), .ZN(n10681) );
  INV_X1 U11394 ( .A(n10681), .ZN(n10358) );
  AOI22_X1 U11395 ( .A1(n9893), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n9882), .B2(
        n10358), .ZN(n9630) );
  AND2_X2 U11396 ( .A1(n9631), .A2(n9630), .ZN(n15880) );
  NAND2_X1 U11397 ( .A1(n15880), .A2(n14742), .ZN(n12716) );
  INV_X1 U11398 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9632) );
  OR2_X1 U11399 ( .A1(n9679), .A2(n11159), .ZN(n9634) );
  INV_X1 U11400 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n11158) );
  OR2_X1 U11401 ( .A1(n9653), .A2(n11158), .ZN(n9633) );
  NAND2_X1 U11402 ( .A1(n9634), .A2(n9633), .ZN(n9635) );
  INV_X1 U11403 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9637) );
  NAND2_X1 U11404 ( .A1(n10305), .A2(n10276), .ZN(n9646) );
  AND2_X1 U11405 ( .A1(n9648), .A2(n8804), .ZN(n9640) );
  NOR2_X1 U11406 ( .A1(n15432), .A2(n9640), .ZN(n9645) );
  NAND2_X1 U11407 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9641) );
  MUX2_X1 U11408 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9641), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n9643) );
  NAND2_X1 U11409 ( .A1(n9643), .A2(n9642), .ZN(n14745) );
  INV_X1 U11410 ( .A(n14745), .ZN(n14753) );
  AND3_X1 U11411 ( .A1(n15432), .A2(n14753), .A3(n15429), .ZN(n9644) );
  NAND2_X1 U11412 ( .A1(n9648), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9647) );
  OAI21_X1 U11413 ( .B1(n10305), .B2(n9648), .A(n9647), .ZN(n9649) );
  INV_X1 U11414 ( .A(n15429), .ZN(n10353) );
  NAND2_X1 U11415 ( .A1(n9649), .A2(n10353), .ZN(n9650) );
  NAND2_X1 U11416 ( .A1(n9985), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9656) );
  INV_X1 U11417 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10574) );
  INV_X1 U11418 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10356) );
  OR2_X1 U11419 ( .A1(n9679), .A2(n10356), .ZN(n9655) );
  INV_X1 U11420 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9652) );
  OR2_X1 U11421 ( .A1(n9653), .A2(n9652), .ZN(n9654) );
  INV_X1 U11422 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10657) );
  NOR2_X1 U11423 ( .A1(n9648), .A2(n9657), .ZN(n9658) );
  XNOR2_X1 U11424 ( .A(n9658), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n15445) );
  MUX2_X1 U11425 ( .A(n10657), .B(n15445), .S(n10323), .Z(n10634) );
  INV_X1 U11426 ( .A(n10634), .ZN(n11155) );
  AND2_X1 U11427 ( .A1(n10632), .A2(n11155), .ZN(n11163) );
  NAND2_X1 U11428 ( .A1(n10302), .A2(n12860), .ZN(n9664) );
  NAND2_X1 U11429 ( .A1(n9661), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9662) );
  XNOR2_X1 U11430 ( .A(n9662), .B(P1_IR_REG_3__SCAN_IN), .ZN(n14760) );
  AOI22_X1 U11431 ( .A1(n9893), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n9882), .B2(
        n14760), .ZN(n9663) );
  NAND2_X1 U11432 ( .A1(n9985), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9669) );
  INV_X1 U11433 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10359) );
  OR2_X1 U11434 ( .A1(n9679), .A2(n10359), .ZN(n9668) );
  OR2_X1 U11435 ( .A1(n9653), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9667) );
  INV_X1 U11436 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10344) );
  OR2_X1 U11437 ( .A1(n9665), .A2(n10344), .ZN(n9666) );
  INV_X1 U11438 ( .A(n12876), .ZN(n9670) );
  INV_X1 U11439 ( .A(n12723), .ZN(n15898) );
  INV_X1 U11440 ( .A(n14741), .ZN(n12721) );
  NAND2_X1 U11441 ( .A1(n10296), .A2(n12860), .ZN(n9678) );
  AND2_X1 U11442 ( .A1(n9628), .A2(n9671), .ZN(n9675) );
  INV_X1 U11443 ( .A(n9675), .ZN(n9672) );
  NAND2_X1 U11444 ( .A1(n9672), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9673) );
  MUX2_X1 U11445 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9673), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n9676) );
  INV_X1 U11446 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9674) );
  NAND2_X1 U11447 ( .A1(n9675), .A2(n9674), .ZN(n9699) );
  NAND2_X1 U11448 ( .A1(n9676), .A2(n9699), .ZN(n10668) );
  INV_X1 U11449 ( .A(n10668), .ZN(n10361) );
  AOI22_X1 U11450 ( .A1(n9893), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n9882), .B2(
        n10361), .ZN(n9677) );
  NAND2_X1 U11451 ( .A1(n9985), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9683) );
  INV_X1 U11452 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10347) );
  OR2_X1 U11453 ( .A1(n9665), .A2(n10347), .ZN(n9682) );
  OAI21_X1 U11454 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n9692), .ZN(n11117) );
  OR2_X1 U11455 ( .A1(n9988), .A2(n11117), .ZN(n9681) );
  INV_X1 U11456 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n11116) );
  OR2_X1 U11457 ( .A1(n9987), .A2(n11116), .ZN(n9680) );
  NAND4_X1 U11458 ( .A1(n9683), .A2(n9682), .A3(n9681), .A4(n9680), .ZN(n14740) );
  NAND2_X1 U11459 ( .A1(n12729), .A2(n14740), .ZN(n9684) );
  AND2_X1 U11460 ( .A1(n9685), .A2(n9684), .ZN(n11075) );
  NAND2_X1 U11461 ( .A1(n9699), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9686) );
  XNOR2_X1 U11462 ( .A(n9686), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10375) );
  AOI22_X1 U11463 ( .A1(n9893), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n9882), .B2(
        n10375), .ZN(n9687) );
  NAND2_X1 U11464 ( .A1(n9985), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9697) );
  INV_X1 U11465 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9689) );
  OR2_X1 U11466 ( .A1(n9665), .A2(n9689), .ZN(n9696) );
  INV_X1 U11467 ( .A(n9690), .ZN(n9705) );
  NAND2_X1 U11468 ( .A1(n9692), .A2(n9691), .ZN(n9693) );
  NAND2_X1 U11469 ( .A1(n9705), .A2(n9693), .ZN(n15912) );
  OR2_X1 U11470 ( .A1(n9653), .A2(n15912), .ZN(n9695) );
  INV_X1 U11471 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10389) );
  OR2_X1 U11472 ( .A1(n9987), .A2(n10389), .ZN(n9694) );
  NAND4_X1 U11473 ( .A1(n9697), .A2(n9696), .A3(n9695), .A4(n9694), .ZN(n14739) );
  INV_X1 U11474 ( .A(n12879), .ZN(n11079) );
  NAND2_X1 U11475 ( .A1(n11075), .A2(n11079), .ZN(n11074) );
  INV_X1 U11476 ( .A(n12738), .ZN(n15916) );
  INV_X1 U11477 ( .A(n14739), .ZN(n10013) );
  NAND2_X1 U11478 ( .A1(n15916), .A2(n10013), .ZN(n9698) );
  NAND2_X1 U11479 ( .A1(n11074), .A2(n9698), .ZN(n10801) );
  NAND2_X1 U11480 ( .A1(n10314), .A2(n12860), .ZN(n9702) );
  NAND2_X1 U11481 ( .A1(n9712), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9700) );
  XNOR2_X1 U11482 ( .A(n9700), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10391) );
  AOI22_X1 U11483 ( .A1(n9893), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9882), .B2(
        n10391), .ZN(n9701) );
  NAND2_X1 U11484 ( .A1(n10336), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9710) );
  INV_X1 U11485 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9703) );
  OR2_X1 U11486 ( .A1(n10057), .A2(n9703), .ZN(n9709) );
  INV_X1 U11487 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9704) );
  NAND2_X1 U11488 ( .A1(n9705), .A2(n9704), .ZN(n9706) );
  NAND2_X1 U11489 ( .A1(n9718), .A2(n9706), .ZN(n11302) );
  OR2_X1 U11490 ( .A1(n9988), .A2(n11302), .ZN(n9708) );
  INV_X1 U11491 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10809) );
  OR2_X1 U11492 ( .A1(n9987), .A2(n10809), .ZN(n9707) );
  NAND4_X1 U11493 ( .A1(n9710), .A2(n9709), .A3(n9708), .A4(n9707), .ZN(n14738) );
  XNOR2_X1 U11494 ( .A(n12741), .B(n14738), .ZN(n12880) );
  INV_X1 U11495 ( .A(n12880), .ZN(n10802) );
  NAND2_X1 U11496 ( .A1(n10801), .A2(n10802), .ZN(n10800) );
  OR2_X1 U11497 ( .A1(n12741), .A2(n14738), .ZN(n9711) );
  NAND2_X1 U11498 ( .A1(n10800), .A2(n9711), .ZN(n11044) );
  OR2_X1 U11499 ( .A1(n10321), .A2(n12853), .ZN(n9715) );
  OAI21_X1 U11500 ( .B1(n9712), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9713) );
  XNOR2_X1 U11501 ( .A(n9713), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10407) );
  AOI22_X1 U11502 ( .A1(n9893), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9882), .B2(
        n10407), .ZN(n9714) );
  NAND2_X1 U11503 ( .A1(n9715), .A2(n9714), .ZN(n12749) );
  NAND2_X1 U11504 ( .A1(n10336), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9723) );
  INV_X1 U11505 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9716) );
  OR2_X1 U11506 ( .A1(n10057), .A2(n9716), .ZN(n9722) );
  NAND2_X1 U11507 ( .A1(n9718), .A2(n9717), .ZN(n9719) );
  NAND2_X1 U11508 ( .A1(n9733), .A2(n9719), .ZN(n11493) );
  OR2_X1 U11509 ( .A1(n9988), .A2(n11493), .ZN(n9721) );
  INV_X1 U11510 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n11357) );
  OR2_X1 U11511 ( .A1(n9987), .A2(n11357), .ZN(n9720) );
  NAND4_X1 U11512 ( .A1(n9723), .A2(n9722), .A3(n9721), .A4(n9720), .ZN(n14737) );
  XNOR2_X1 U11513 ( .A(n12749), .B(n14737), .ZN(n12882) );
  INV_X1 U11514 ( .A(n12882), .ZN(n11043) );
  NAND2_X1 U11515 ( .A1(n11044), .A2(n11043), .ZN(n11042) );
  INV_X1 U11516 ( .A(n14737), .ZN(n11489) );
  NAND2_X1 U11517 ( .A1(n11499), .A2(n11489), .ZN(n9724) );
  NAND2_X1 U11518 ( .A1(n11042), .A2(n9724), .ZN(n11444) );
  OR2_X1 U11519 ( .A1(n10372), .A2(n12853), .ZN(n9731) );
  INV_X1 U11520 ( .A(n9725), .ZN(n9726) );
  NAND2_X1 U11521 ( .A1(n9726), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9727) );
  MUX2_X1 U11522 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9727), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n9729) );
  INV_X1 U11523 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9728) );
  NAND2_X1 U11524 ( .A1(n9725), .A2(n9728), .ZN(n9741) );
  NAND2_X1 U11525 ( .A1(n9729), .A2(n9741), .ZN(n10392) );
  INV_X1 U11526 ( .A(n10392), .ZN(n10428) );
  AOI22_X1 U11527 ( .A1(n9893), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9882), .B2(
        n10428), .ZN(n9730) );
  NAND2_X1 U11528 ( .A1(n9985), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n9738) );
  INV_X1 U11529 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10383) );
  OR2_X1 U11530 ( .A1(n9665), .A2(n10383), .ZN(n9737) );
  NAND2_X1 U11531 ( .A1(n9733), .A2(n9732), .ZN(n9734) );
  NAND2_X1 U11532 ( .A1(n9748), .A2(n9734), .ZN(n11768) );
  OR2_X1 U11533 ( .A1(n9988), .A2(n11768), .ZN(n9736) );
  INV_X1 U11534 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10393) );
  OR2_X1 U11535 ( .A1(n9987), .A2(n10393), .ZN(n9735) );
  NAND4_X1 U11536 ( .A1(n9738), .A2(n9737), .A3(n9736), .A4(n9735), .ZN(n14736) );
  INV_X1 U11537 ( .A(n14736), .ZN(n11756) );
  XNOR2_X1 U11538 ( .A(n12753), .B(n11756), .ZN(n12884) );
  NAND2_X1 U11539 ( .A1(n11444), .A2(n12884), .ZN(n11446) );
  OR2_X1 U11540 ( .A1(n12753), .A2(n14736), .ZN(n9739) );
  NAND2_X1 U11541 ( .A1(n11446), .A2(n9739), .ZN(n11698) );
  OR2_X1 U11542 ( .A1(n10433), .A2(n12853), .ZN(n9744) );
  NAND2_X1 U11543 ( .A1(n9741), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9740) );
  MUX2_X1 U11544 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9740), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n9742) );
  AOI22_X1 U11545 ( .A1(n9893), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9882), .B2(
        n10432), .ZN(n9743) );
  NAND2_X1 U11546 ( .A1(n9985), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9754) );
  INV_X1 U11547 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9745) );
  OR2_X1 U11548 ( .A1(n9665), .A2(n9745), .ZN(n9753) );
  INV_X1 U11549 ( .A(n9746), .ZN(n9761) );
  NAND2_X1 U11550 ( .A1(n9748), .A2(n9747), .ZN(n9749) );
  NAND2_X1 U11551 ( .A1(n9761), .A2(n9749), .ZN(n15937) );
  OR2_X1 U11552 ( .A1(n9988), .A2(n15937), .ZN(n9752) );
  INV_X1 U11553 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9750) );
  OR2_X1 U11554 ( .A1(n9987), .A2(n9750), .ZN(n9751) );
  NAND4_X1 U11555 ( .A1(n9754), .A2(n9753), .A3(n9752), .A4(n9751), .ZN(n14735) );
  XNOR2_X1 U11556 ( .A(n12760), .B(n14735), .ZN(n12885) );
  INV_X1 U11557 ( .A(n12885), .ZN(n11697) );
  NAND2_X1 U11558 ( .A1(n11698), .A2(n11697), .ZN(n11696) );
  OR2_X1 U11559 ( .A1(n12760), .A2(n14735), .ZN(n9755) );
  NAND2_X1 U11560 ( .A1(n11696), .A2(n9755), .ZN(n11509) );
  OR2_X1 U11561 ( .A1(n10471), .A2(n12853), .ZN(n9758) );
  NAND2_X1 U11562 ( .A1(n9768), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9756) );
  XNOR2_X1 U11563 ( .A(n9756), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10599) );
  AOI22_X1 U11564 ( .A1(n9893), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n9882), 
        .B2(n10599), .ZN(n9757) );
  NAND2_X1 U11565 ( .A1(n10336), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9766) );
  INV_X1 U11566 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9759) );
  OR2_X1 U11567 ( .A1(n10057), .A2(n9759), .ZN(n9765) );
  INV_X1 U11568 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9760) );
  NAND2_X1 U11569 ( .A1(n9761), .A2(n9760), .ZN(n9762) );
  NAND2_X1 U11570 ( .A1(n9775), .A2(n9762), .ZN(n12164) );
  OR2_X1 U11571 ( .A1(n9988), .A2(n12164), .ZN(n9764) );
  INV_X1 U11572 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10550) );
  OR2_X1 U11573 ( .A1(n9987), .A2(n10550), .ZN(n9763) );
  NAND4_X1 U11574 ( .A1(n9766), .A2(n9765), .A3(n9764), .A4(n9763), .ZN(n14734) );
  XNOR2_X1 U11575 ( .A(n12764), .B(n14734), .ZN(n12886) );
  INV_X1 U11576 ( .A(n12886), .ZN(n11511) );
  OR2_X1 U11577 ( .A1(n12764), .A2(n14734), .ZN(n9767) );
  NAND2_X1 U11578 ( .A1(n10610), .A2(n12860), .ZN(n9773) );
  INV_X1 U11579 ( .A(n9768), .ZN(n9770) );
  INV_X1 U11580 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9769) );
  NAND2_X1 U11581 ( .A1(n9770), .A2(n9769), .ZN(n9782) );
  NAND2_X1 U11582 ( .A1(n9782), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9771) );
  XNOR2_X1 U11583 ( .A(n9771), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U11584 ( .A1(n9893), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9882), 
        .B2(n10773), .ZN(n9772) );
  NAND2_X1 U11585 ( .A1(n9985), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n9780) );
  INV_X1 U11586 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9774) );
  OR2_X1 U11587 ( .A1(n9665), .A2(n9774), .ZN(n9779) );
  NAND2_X1 U11588 ( .A1(n9775), .A2(n10596), .ZN(n9776) );
  NAND2_X1 U11589 ( .A1(n9789), .A2(n9776), .ZN(n12311) );
  OR2_X1 U11590 ( .A1(n9988), .A2(n12311), .ZN(n9778) );
  INV_X1 U11591 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11579) );
  OR2_X1 U11592 ( .A1(n9987), .A2(n11579), .ZN(n9777) );
  NAND4_X1 U11593 ( .A1(n9780), .A2(n9779), .A3(n9778), .A4(n9777), .ZN(n14733) );
  INV_X1 U11594 ( .A(n9781), .ZN(n11866) );
  NAND2_X1 U11595 ( .A1(n10739), .A2(n12860), .ZN(n9785) );
  NAND2_X1 U11596 ( .A1(n9783), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9798) );
  XNOR2_X1 U11597 ( .A(n9798), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11001) );
  AOI22_X1 U11598 ( .A1(n9893), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n11001), 
        .B2(n9882), .ZN(n9784) );
  NAND2_X1 U11599 ( .A1(n9985), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9795) );
  INV_X1 U11600 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9786) );
  OR2_X1 U11601 ( .A1(n9987), .A2(n9786), .ZN(n9794) );
  INV_X1 U11602 ( .A(n9787), .ZN(n9803) );
  NAND2_X1 U11603 ( .A1(n9789), .A2(n9788), .ZN(n9790) );
  NAND2_X1 U11604 ( .A1(n9803), .A2(n9790), .ZN(n11869) );
  OR2_X1 U11605 ( .A1(n9988), .A2(n11869), .ZN(n9793) );
  INV_X1 U11606 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9791) );
  OR2_X1 U11607 ( .A1(n9665), .A2(n9791), .ZN(n9792) );
  NAND4_X1 U11608 ( .A1(n9795), .A2(n9794), .A3(n9793), .A4(n9792), .ZN(n14732) );
  INV_X1 U11609 ( .A(n14732), .ZN(n12320) );
  XNOR2_X1 U11610 ( .A(n12777), .B(n12320), .ZN(n12890) );
  INV_X1 U11611 ( .A(n12890), .ZN(n11862) );
  OR2_X1 U11612 ( .A1(n12777), .A2(n14732), .ZN(n9796) );
  INV_X1 U11613 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9797) );
  NAND2_X1 U11614 ( .A1(n9798), .A2(n9797), .ZN(n9799) );
  NAND2_X1 U11615 ( .A1(n9799), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9813) );
  XNOR2_X1 U11616 ( .A(n9813), .B(P1_IR_REG_13__SCAN_IN), .ZN(n11630) );
  AOI22_X1 U11617 ( .A1(n11630), .A2(n9882), .B1(P2_DATAO_REG_13__SCAN_IN), 
        .B2(n9893), .ZN(n9800) );
  INV_X1 U11618 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9802) );
  NAND2_X1 U11619 ( .A1(n9803), .A2(n9802), .ZN(n9804) );
  AND2_X1 U11620 ( .A1(n9819), .A2(n9804), .ZN(n12395) );
  NAND2_X1 U11621 ( .A1(n12395), .A2(n9899), .ZN(n9810) );
  NAND2_X1 U11622 ( .A1(n9985), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n9809) );
  INV_X1 U11623 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9805) );
  OR2_X1 U11624 ( .A1(n9665), .A2(n9805), .ZN(n9808) );
  INV_X1 U11625 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9806) );
  OR2_X1 U11626 ( .A1(n9987), .A2(n9806), .ZN(n9807) );
  NAND4_X1 U11627 ( .A1(n9810), .A2(n9809), .A3(n9808), .A4(n9807), .ZN(n14731) );
  INV_X1 U11628 ( .A(n14731), .ZN(n12393) );
  XNOR2_X1 U11629 ( .A(n15983), .B(n12393), .ZN(n12891) );
  OR2_X1 U11630 ( .A1(n15983), .A2(n14731), .ZN(n9811) );
  NAND2_X1 U11631 ( .A1(n10817), .A2(n12860), .ZN(n9817) );
  INV_X1 U11632 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9812) );
  NAND2_X1 U11633 ( .A1(n9813), .A2(n9812), .ZN(n9814) );
  NAND2_X1 U11634 ( .A1(n9814), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9815) );
  XNOR2_X1 U11635 ( .A(n9815), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11888) );
  AOI22_X1 U11636 ( .A1(n11888), .A2(n9882), .B1(n9893), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n9816) );
  NAND2_X1 U11637 ( .A1(n9819), .A2(n9818), .ZN(n9820) );
  NAND2_X1 U11638 ( .A1(n9832), .A2(n9820), .ZN(n14557) );
  NAND2_X1 U11639 ( .A1(n10336), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9822) );
  NAND2_X1 U11640 ( .A1(n9985), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n9821) );
  AND2_X1 U11641 ( .A1(n9822), .A2(n9821), .ZN(n9824) );
  NAND2_X1 U11642 ( .A1(n10335), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9823) );
  OAI211_X1 U11643 ( .C1(n14557), .C2(n9988), .A(n9824), .B(n9823), .ZN(n14730) );
  INV_X1 U11644 ( .A(n14730), .ZN(n14446) );
  NAND2_X1 U11645 ( .A1(n14561), .A2(n14446), .ZN(n10026) );
  OR2_X1 U11646 ( .A1(n14561), .A2(n14446), .ZN(n9825) );
  NAND2_X1 U11647 ( .A1(n10026), .A2(n9825), .ZN(n12892) );
  NAND2_X1 U11648 ( .A1(n11290), .A2(n12860), .ZN(n9830) );
  NAND2_X1 U11649 ( .A1(n9827), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9828) );
  XNOR2_X1 U11650 ( .A(n9828), .B(P1_IR_REG_15__SCAN_IN), .ZN(n14790) );
  AOI22_X1 U11651 ( .A1(n9893), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9882), 
        .B2(n14790), .ZN(n9829) );
  INV_X1 U11652 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n15053) );
  INV_X1 U11653 ( .A(n9831), .ZN(n9845) );
  NAND2_X1 U11654 ( .A1(n9832), .A2(n14705), .ZN(n9833) );
  NAND2_X1 U11655 ( .A1(n9845), .A2(n9833), .ZN(n15052) );
  OR2_X1 U11656 ( .A1(n15052), .A2(n9988), .ZN(n9835) );
  AOI22_X1 U11657 ( .A1(n9985), .A2(P1_REG0_REG_15__SCAN_IN), .B1(n10336), 
        .B2(P1_REG1_REG_15__SCAN_IN), .ZN(n9834) );
  OAI211_X1 U11658 ( .C1(n9987), .C2(n15053), .A(n9835), .B(n9834), .ZN(n14729) );
  INV_X1 U11659 ( .A(n14729), .ZN(n14455) );
  XNOR2_X1 U11660 ( .A(n15413), .B(n14455), .ZN(n15042) );
  INV_X1 U11661 ( .A(n15042), .ZN(n15045) );
  OR2_X1 U11662 ( .A1(n15413), .A2(n14729), .ZN(n9836) );
  NAND2_X1 U11663 ( .A1(n9837), .A2(n9836), .ZN(n15027) );
  NAND2_X1 U11664 ( .A1(n11423), .A2(n12860), .ZN(n9842) );
  NAND2_X1 U11665 ( .A1(n9838), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9839) );
  MUX2_X1 U11666 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9839), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n9840) );
  NAND2_X1 U11667 ( .A1(n9840), .A2(n10068), .ZN(n15563) );
  INV_X1 U11668 ( .A(n15563), .ZN(n14793) );
  AOI22_X1 U11669 ( .A1(n9893), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9882), 
        .B2(n14793), .ZN(n9841) );
  INV_X1 U11670 ( .A(n9843), .ZN(n9858) );
  INV_X1 U11671 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9844) );
  NAND2_X1 U11672 ( .A1(n9845), .A2(n9844), .ZN(n9846) );
  AND2_X1 U11673 ( .A1(n9858), .A2(n9846), .ZN(n15037) );
  NAND2_X1 U11674 ( .A1(n15037), .A2(n9899), .ZN(n9852) );
  INV_X1 U11675 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9849) );
  NAND2_X1 U11676 ( .A1(n10336), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9848) );
  NAND2_X1 U11677 ( .A1(n10335), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9847) );
  OAI211_X1 U11678 ( .C1(n10057), .C2(n9849), .A(n9848), .B(n9847), .ZN(n9850)
         );
  INV_X1 U11679 ( .A(n9850), .ZN(n9851) );
  NAND2_X1 U11680 ( .A1(n9852), .A2(n9851), .ZN(n14728) );
  XNOR2_X1 U11681 ( .A(n15150), .B(n14728), .ZN(n15030) );
  INV_X1 U11682 ( .A(n15030), .ZN(n15026) );
  NAND2_X1 U11683 ( .A1(n15027), .A2(n15026), .ZN(n15025) );
  OR2_X1 U11684 ( .A1(n15150), .A2(n14728), .ZN(n9853) );
  NAND2_X1 U11685 ( .A1(n15025), .A2(n9853), .ZN(n15012) );
  INV_X1 U11686 ( .A(n15012), .ZN(n9866) );
  NAND2_X1 U11687 ( .A1(n11569), .A2(n12860), .ZN(n9856) );
  NAND2_X1 U11688 ( .A1(n10068), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9854) );
  XNOR2_X1 U11689 ( .A(n9854), .B(P1_IR_REG_17__SCAN_IN), .ZN(n15540) );
  AOI22_X1 U11690 ( .A1(n9893), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9882), 
        .B2(n15540), .ZN(n9855) );
  INV_X1 U11691 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9857) );
  NAND2_X1 U11692 ( .A1(n9858), .A2(n9857), .ZN(n9859) );
  NAND2_X1 U11693 ( .A1(n9872), .A2(n9859), .ZN(n15017) );
  OR2_X1 U11694 ( .A1(n15017), .A2(n9988), .ZN(n9864) );
  INV_X1 U11695 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n15016) );
  NAND2_X1 U11696 ( .A1(n9985), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n9861) );
  NAND2_X1 U11697 ( .A1(n10336), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9860) );
  OAI211_X1 U11698 ( .C1(n9987), .C2(n15016), .A(n9861), .B(n9860), .ZN(n9862)
         );
  INV_X1 U11699 ( .A(n9862), .ZN(n9863) );
  NAND2_X1 U11700 ( .A1(n9864), .A2(n9863), .ZN(n14726) );
  XNOR2_X1 U11701 ( .A(n15142), .B(n14726), .ZN(n15013) );
  NAND2_X1 U11702 ( .A1(n15142), .A2(n14726), .ZN(n9867) );
  OR2_X1 U11703 ( .A1(n11975), .A2(n12853), .ZN(n9871) );
  NAND2_X1 U11704 ( .A1(n10060), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9869) );
  XNOR2_X1 U11705 ( .A(n9869), .B(P1_IR_REG_18__SCAN_IN), .ZN(n15547) );
  AOI22_X1 U11706 ( .A1(n9893), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n15547), 
        .B2(n9882), .ZN(n9870) );
  NAND2_X1 U11707 ( .A1(n9872), .A2(n14681), .ZN(n9873) );
  NAND2_X1 U11708 ( .A1(n9886), .A2(n9873), .ZN(n15001) );
  OR2_X1 U11709 ( .A1(n15001), .A2(n9988), .ZN(n9879) );
  INV_X1 U11710 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9876) );
  NAND2_X1 U11711 ( .A1(n10336), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9875) );
  NAND2_X1 U11712 ( .A1(n10335), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9874) );
  OAI211_X1 U11713 ( .C1(n10057), .C2(n9876), .A(n9875), .B(n9874), .ZN(n9877)
         );
  INV_X1 U11714 ( .A(n9877), .ZN(n9878) );
  NAND2_X1 U11715 ( .A1(n9879), .A2(n9878), .ZN(n14725) );
  XNOR2_X1 U11716 ( .A(n15407), .B(n14725), .ZN(n14998) );
  INV_X1 U11717 ( .A(n14998), .ZN(n14994) );
  INV_X1 U11718 ( .A(n14725), .ZN(n14432) );
  NAND2_X1 U11719 ( .A1(n14686), .A2(n14432), .ZN(n9880) );
  NAND2_X1 U11720 ( .A1(n12066), .A2(n12860), .ZN(n9884) );
  XNOR2_X1 U11721 ( .A(n9881), .B(P1_IR_REG_19__SCAN_IN), .ZN(n10000) );
  AOI22_X1 U11722 ( .A1(n10000), .A2(n9882), .B1(n9893), .B2(
        P2_DATAO_REG_19__SCAN_IN), .ZN(n9883) );
  NAND2_X1 U11723 ( .A1(n9886), .A2(n9885), .ZN(n9887) );
  NAND2_X1 U11724 ( .A1(n9896), .A2(n9887), .ZN(n14984) );
  INV_X1 U11725 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14798) );
  NAND2_X1 U11726 ( .A1(n10335), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n9889) );
  NAND2_X1 U11727 ( .A1(n9985), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9888) );
  OAI211_X1 U11728 ( .C1(n9665), .C2(n14798), .A(n9889), .B(n9888), .ZN(n9890)
         );
  INV_X1 U11729 ( .A(n9890), .ZN(n9891) );
  OAI21_X1 U11730 ( .B1(n14984), .B2(n9988), .A(n9891), .ZN(n14724) );
  INV_X1 U11731 ( .A(n14724), .ZN(n10032) );
  XNOR2_X1 U11732 ( .A(n14980), .B(n10032), .ZN(n14978) );
  OR2_X1 U11733 ( .A1(n14980), .A2(n14724), .ZN(n9892) );
  NAND2_X1 U11734 ( .A1(n14977), .A2(n9892), .ZN(n14961) );
  NAND2_X1 U11735 ( .A1(n12272), .A2(n12860), .ZN(n9895) );
  OR2_X1 U11736 ( .A1(n12863), .A2(n12273), .ZN(n9894) );
  INV_X1 U11737 ( .A(n9909), .ZN(n9898) );
  NAND2_X1 U11738 ( .A1(n9896), .A2(n14658), .ZN(n9897) );
  NAND2_X1 U11739 ( .A1(n14968), .A2(n9899), .ZN(n9904) );
  INV_X1 U11740 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n15400) );
  NAND2_X1 U11741 ( .A1(n10336), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n9901) );
  NAND2_X1 U11742 ( .A1(n10335), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9900) );
  OAI211_X1 U11743 ( .C1(n10057), .C2(n15400), .A(n9901), .B(n9900), .ZN(n9902) );
  INV_X1 U11744 ( .A(n9902), .ZN(n9903) );
  NAND2_X1 U11745 ( .A1(n9904), .A2(n9903), .ZN(n14723) );
  INV_X1 U11746 ( .A(n14723), .ZN(n14606) );
  XNOR2_X1 U11747 ( .A(n14967), .B(n14606), .ZN(n12896) );
  NAND2_X1 U11748 ( .A1(n14967), .A2(n14723), .ZN(n9906) );
  NAND2_X1 U11749 ( .A1(n12354), .A2(n12860), .ZN(n9908) );
  OR2_X1 U11750 ( .A1(n12863), .A2(n12355), .ZN(n9907) );
  NOR2_X1 U11751 ( .A1(n9909), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9910) );
  OR2_X1 U11752 ( .A1(n9911), .A2(n9910), .ZN(n14950) );
  INV_X1 U11753 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9914) );
  NAND2_X1 U11754 ( .A1(n10336), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n9913) );
  NAND2_X1 U11755 ( .A1(n10335), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9912) );
  OAI211_X1 U11756 ( .C1(n10057), .C2(n9914), .A(n9913), .B(n9912), .ZN(n9915)
         );
  INV_X1 U11757 ( .A(n9915), .ZN(n9916) );
  INV_X1 U11758 ( .A(n14722), .ZN(n10035) );
  XNOR2_X1 U11759 ( .A(n15115), .B(n10035), .ZN(n14943) );
  NOR2_X1 U11760 ( .A1(n15115), .A2(n14722), .ZN(n9917) );
  NAND2_X1 U11761 ( .A1(n15108), .A2(n14608), .ZN(n9918) );
  NAND2_X1 U11762 ( .A1(n14418), .A2(n12860), .ZN(n9920) );
  OR2_X1 U11763 ( .A1(n12863), .A2(n15442), .ZN(n9919) );
  NAND2_X1 U11764 ( .A1(n10336), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n9927) );
  INV_X1 U11765 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9921) );
  OR2_X1 U11766 ( .A1(n10057), .A2(n9921), .ZN(n9926) );
  OAI21_X1 U11767 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n9923), .A(n9932), .ZN(
        n14919) );
  OR2_X1 U11768 ( .A1(n9988), .A2(n14919), .ZN(n9925) );
  INV_X1 U11769 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n14920) );
  OR2_X1 U11770 ( .A1(n9987), .A2(n14920), .ZN(n9924) );
  NAND4_X1 U11771 ( .A1(n9927), .A2(n9926), .A3(n9925), .A4(n9924), .ZN(n14720) );
  INV_X1 U11772 ( .A(n14720), .ZN(n10038) );
  XNOR2_X1 U11773 ( .A(n15100), .B(n10038), .ZN(n14926) );
  NAND2_X1 U11774 ( .A1(n15100), .A2(n14720), .ZN(n9928) );
  NAND2_X1 U11775 ( .A1(n12457), .A2(n12860), .ZN(n9930) );
  OR2_X1 U11776 ( .A1(n12863), .A2(n7394), .ZN(n9929) );
  NAND2_X1 U11777 ( .A1(n10336), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n9937) );
  INV_X1 U11778 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n15394) );
  OR2_X1 U11779 ( .A1(n10057), .A2(n15394), .ZN(n9936) );
  INV_X1 U11780 ( .A(n9932), .ZN(n9931) );
  NAND2_X1 U11781 ( .A1(n9931), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9942) );
  INV_X1 U11782 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n14650) );
  NAND2_X1 U11783 ( .A1(n9932), .A2(n14650), .ZN(n9933) );
  NAND2_X1 U11784 ( .A1(n9942), .A2(n9933), .ZN(n14906) );
  OR2_X1 U11785 ( .A1(n9988), .A2(n14906), .ZN(n9935) );
  INV_X1 U11786 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n14907) );
  OR2_X1 U11787 ( .A1(n9987), .A2(n14907), .ZN(n9934) );
  NAND4_X1 U11788 ( .A1(n9937), .A2(n9936), .A3(n9935), .A4(n9934), .ZN(n14719) );
  XNOR2_X1 U11789 ( .A(n14905), .B(n14719), .ZN(n12897) );
  OR2_X1 U11790 ( .A1(n14905), .A2(n14719), .ZN(n9938) );
  NAND2_X1 U11791 ( .A1(n12479), .A2(n12860), .ZN(n9940) );
  OR2_X1 U11792 ( .A1(n12863), .A2(n7369), .ZN(n9939) );
  NAND2_X1 U11793 ( .A1(n10336), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n9947) );
  INV_X1 U11794 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n15390) );
  OR2_X1 U11795 ( .A1(n10057), .A2(n15390), .ZN(n9946) );
  INV_X1 U11796 ( .A(n9942), .ZN(n9941) );
  NAND2_X1 U11797 ( .A1(n9941), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9953) );
  INV_X1 U11798 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14621) );
  NAND2_X1 U11799 ( .A1(n9942), .A2(n14621), .ZN(n9943) );
  NAND2_X1 U11800 ( .A1(n9953), .A2(n9943), .ZN(n14894) );
  OR2_X1 U11801 ( .A1(n9988), .A2(n14894), .ZN(n9945) );
  INV_X1 U11802 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n14893) );
  OR2_X1 U11803 ( .A1(n9987), .A2(n14893), .ZN(n9944) );
  NAND4_X1 U11804 ( .A1(n9947), .A2(n9946), .A3(n9945), .A4(n9944), .ZN(n14718) );
  XNOR2_X1 U11805 ( .A(n14897), .B(n14718), .ZN(n12899) );
  NAND2_X1 U11806 ( .A1(n14897), .A2(n14718), .ZN(n9948) );
  NAND2_X1 U11807 ( .A1(n14414), .A2(n12860), .ZN(n9950) );
  OR2_X1 U11808 ( .A1(n12863), .A2(n8134), .ZN(n9949) );
  NAND2_X1 U11809 ( .A1(n10336), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n9959) );
  INV_X1 U11810 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9951) );
  OR2_X1 U11811 ( .A1(n10057), .A2(n9951), .ZN(n9958) );
  INV_X1 U11812 ( .A(n9953), .ZN(n9952) );
  NAND2_X1 U11813 ( .A1(n9952), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n9972) );
  INV_X1 U11814 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14692) );
  NAND2_X1 U11815 ( .A1(n9953), .A2(n14692), .ZN(n9954) );
  NAND2_X1 U11816 ( .A1(n9972), .A2(n9954), .ZN(n14880) );
  OR2_X1 U11817 ( .A1(n9988), .A2(n14880), .ZN(n9957) );
  INV_X1 U11818 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9955) );
  OR2_X1 U11819 ( .A1(n9987), .A2(n9955), .ZN(n9956) );
  NAND4_X1 U11820 ( .A1(n9959), .A2(n9958), .A3(n9957), .A4(n9956), .ZN(n14717) );
  INV_X1 U11821 ( .A(n14717), .ZN(n9960) );
  OR2_X1 U11822 ( .A1(n15079), .A2(n9960), .ZN(n10044) );
  NAND2_X1 U11823 ( .A1(n15079), .A2(n9960), .ZN(n9961) );
  NAND2_X1 U11824 ( .A1(n10044), .A2(n9961), .ZN(n12902) );
  NAND2_X1 U11825 ( .A1(n14886), .A2(n12902), .ZN(n9963) );
  NAND2_X1 U11826 ( .A1(n15079), .A2(n14717), .ZN(n9962) );
  NAND2_X1 U11827 ( .A1(n9963), .A2(n9962), .ZN(n14859) );
  NAND2_X1 U11828 ( .A1(n14410), .A2(n12860), .ZN(n9965) );
  OR2_X1 U11829 ( .A1(n12863), .A2(n15434), .ZN(n9964) );
  NAND2_X1 U11830 ( .A1(n9985), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n9969) );
  INV_X1 U11831 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n14868) );
  OR2_X1 U11832 ( .A1(n9987), .A2(n14868), .ZN(n9968) );
  INV_X1 U11833 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n14549) );
  XNOR2_X1 U11834 ( .A(n9972), .B(n14549), .ZN(n14867) );
  OR2_X1 U11835 ( .A1(n9988), .A2(n14867), .ZN(n9967) );
  INV_X1 U11836 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n15074) );
  OR2_X1 U11837 ( .A1(n9665), .A2(n15074), .ZN(n9966) );
  NAND4_X1 U11838 ( .A1(n9969), .A2(n9968), .A3(n9967), .A4(n9966), .ZN(n14716) );
  XNOR2_X1 U11839 ( .A(n14870), .B(n14716), .ZN(n14861) );
  OAI22_X1 U11840 ( .A1(n14859), .A2(n14861), .B1(n14716), .B2(n14870), .ZN(
        n10218) );
  NAND2_X1 U11841 ( .A1(n15428), .A2(n12860), .ZN(n9971) );
  OR2_X1 U11842 ( .A1(n12863), .A2(n15431), .ZN(n9970) );
  NAND2_X1 U11843 ( .A1(n9985), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n9979) );
  INV_X1 U11844 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n10228) );
  OR2_X1 U11845 ( .A1(n9665), .A2(n10228), .ZN(n9978) );
  INV_X1 U11846 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n14595) );
  OAI21_X1 U11847 ( .B1(n9972), .B2(n14549), .A(n14595), .ZN(n9975) );
  INV_X1 U11848 ( .A(n9972), .ZN(n9974) );
  AND2_X1 U11849 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n9973) );
  NAND2_X1 U11850 ( .A1(n9974), .A2(n9973), .ZN(n14835) );
  NAND2_X1 U11851 ( .A1(n9975), .A2(n14835), .ZN(n14850) );
  OR2_X1 U11852 ( .A1(n9988), .A2(n14850), .ZN(n9977) );
  INV_X1 U11853 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n14851) );
  OR2_X1 U11854 ( .A1(n9987), .A2(n14851), .ZN(n9976) );
  NAND4_X1 U11855 ( .A1(n9979), .A2(n9978), .A3(n9977), .A4(n9976), .ZN(n14715) );
  INV_X1 U11856 ( .A(n14715), .ZN(n14589) );
  NAND2_X1 U11857 ( .A1(n14599), .A2(n14589), .ZN(n10047) );
  OR2_X1 U11858 ( .A1(n14599), .A2(n14589), .ZN(n9980) );
  NAND2_X1 U11859 ( .A1(n10047), .A2(n9980), .ZN(n12901) );
  INV_X1 U11860 ( .A(n12901), .ZN(n9981) );
  NAND2_X1 U11861 ( .A1(n14599), .A2(n14715), .ZN(n9982) );
  NAND2_X1 U11862 ( .A1(n7190), .A2(n9982), .ZN(n9994) );
  NAND2_X1 U11863 ( .A1(n12956), .A2(n12860), .ZN(n9984) );
  OR2_X1 U11864 ( .A1(n12863), .A2(n12958), .ZN(n9983) );
  NAND2_X1 U11865 ( .A1(n9985), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9993) );
  INV_X1 U11866 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9986) );
  OR2_X1 U11867 ( .A1(n9987), .A2(n9986), .ZN(n9992) );
  OR2_X1 U11868 ( .A1(n9653), .A2(n14835), .ZN(n9991) );
  INV_X1 U11869 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9989) );
  OR2_X1 U11870 ( .A1(n9665), .A2(n9989), .ZN(n9990) );
  AND4_X1 U11871 ( .A1(n9993), .A2(n9992), .A3(n9991), .A4(n9990), .ZN(n12872)
         );
  XNOR2_X1 U11872 ( .A(n10099), .B(n14714), .ZN(n12904) );
  XNOR2_X1 U11873 ( .A(n9994), .B(n12904), .ZN(n14833) );
  INV_X2 U11874 ( .A(n10000), .ZN(n14816) );
  NAND2_X1 U11875 ( .A1(n10002), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10003) );
  INV_X1 U11876 ( .A(n10005), .ZN(n10006) );
  NAND2_X1 U11877 ( .A1(n10006), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10008) );
  NAND2_X2 U11878 ( .A1(n10633), .A2(n15827), .ZN(n12706) );
  OAI21_X1 U11879 ( .B1(n12702), .B2(n12706), .A(n14586), .ZN(n10799) );
  NAND2_X1 U11880 ( .A1(n10051), .A2(n10000), .ZN(n12703) );
  NAND2_X1 U11881 ( .A1(n14833), .A2(n15992), .ZN(n10059) );
  INV_X1 U11882 ( .A(n14943), .ZN(n14947) );
  INV_X1 U11883 ( .A(n15835), .ZN(n11160) );
  OR2_X1 U11884 ( .A1(n14743), .A2(n11160), .ZN(n10009) );
  NAND2_X1 U11885 ( .A1(n15871), .A2(n10010), .ZN(n11224) );
  NAND2_X1 U11886 ( .A1(n12723), .A2(n12721), .ZN(n12715) );
  NAND2_X1 U11887 ( .A1(n11223), .A2(n12715), .ZN(n10686) );
  INV_X1 U11888 ( .A(n14740), .ZN(n10928) );
  OR2_X1 U11889 ( .A1(n12729), .A2(n10928), .ZN(n10011) );
  NAND2_X1 U11890 ( .A1(n12729), .A2(n10928), .ZN(n10012) );
  NAND2_X1 U11891 ( .A1(n10803), .A2(n12880), .ZN(n10015) );
  INV_X1 U11892 ( .A(n14738), .ZN(n12743) );
  NAND2_X1 U11893 ( .A1(n12741), .A2(n12743), .ZN(n10014) );
  AND2_X1 U11894 ( .A1(n12749), .A2(n11489), .ZN(n10016) );
  NAND2_X1 U11895 ( .A1(n11499), .A2(n14737), .ZN(n10017) );
  INV_X1 U11896 ( .A(n12884), .ZN(n11447) );
  OR2_X1 U11897 ( .A1(n12753), .A2(n11756), .ZN(n10018) );
  NAND2_X1 U11898 ( .A1(n10019), .A2(n10018), .ZN(n11702) );
  INV_X1 U11899 ( .A(n11702), .ZN(n10021) );
  INV_X1 U11900 ( .A(n14735), .ZN(n10020) );
  INV_X1 U11901 ( .A(n14734), .ZN(n12158) );
  OR2_X1 U11902 ( .A1(n12764), .A2(n12158), .ZN(n10022) );
  INV_X1 U11903 ( .A(n14733), .ZN(n12296) );
  NAND2_X1 U11904 ( .A1(n12773), .A2(n12296), .ZN(n10023) );
  OR2_X1 U11905 ( .A1(n12777), .A2(n12320), .ZN(n10024) );
  NAND2_X1 U11906 ( .A1(n11861), .A2(n10024), .ZN(n11962) );
  INV_X1 U11907 ( .A(n12891), .ZN(n11961) );
  NAND2_X1 U11908 ( .A1(n11962), .A2(n11961), .ZN(n11960) );
  OR2_X1 U11909 ( .A1(n15983), .A2(n12393), .ZN(n10025) );
  OR2_X1 U11910 ( .A1(n15413), .A2(n14455), .ZN(n10027) );
  INV_X1 U11911 ( .A(n14728), .ZN(n10028) );
  INV_X1 U11912 ( .A(n14726), .ZN(n10029) );
  AND2_X1 U11913 ( .A1(n15142), .A2(n10029), .ZN(n10030) );
  NAND2_X1 U11914 ( .A1(n14999), .A2(n14998), .ZN(n15134) );
  NAND2_X1 U11915 ( .A1(n14686), .A2(n14725), .ZN(n10031) );
  NAND2_X1 U11916 ( .A1(n14980), .A2(n10032), .ZN(n10033) );
  OR2_X1 U11917 ( .A1(n14967), .A2(n14606), .ZN(n10034) );
  OR2_X1 U11918 ( .A1(n15115), .A2(n10035), .ZN(n10036) );
  NAND2_X1 U11919 ( .A1(n14932), .A2(n14934), .ZN(n14931) );
  OR2_X1 U11920 ( .A1(n14721), .A2(n15108), .ZN(n10037) );
  INV_X1 U11921 ( .A(n14926), .ZN(n14915) );
  NAND2_X1 U11922 ( .A1(n15100), .A2(n10038), .ZN(n10039) );
  INV_X1 U11923 ( .A(n14719), .ZN(n14568) );
  AND2_X1 U11924 ( .A1(n14905), .A2(n14568), .ZN(n10040) );
  OR2_X1 U11925 ( .A1(n14905), .A2(n14568), .ZN(n10041) );
  INV_X1 U11926 ( .A(n12899), .ZN(n14890) );
  INV_X1 U11927 ( .A(n14718), .ZN(n14524) );
  NAND2_X1 U11928 ( .A1(n14897), .A2(n14524), .ZN(n10042) );
  OAI21_X1 U11929 ( .B1(n14891), .B2(n14890), .A(n10042), .ZN(n10043) );
  INV_X1 U11930 ( .A(n14716), .ZN(n10045) );
  NAND2_X1 U11931 ( .A1(n14870), .A2(n10045), .ZN(n10222) );
  NAND2_X1 U11932 ( .A1(n10046), .A2(n9981), .ZN(n10221) );
  NAND2_X1 U11933 ( .A1(n10221), .A2(n10047), .ZN(n10048) );
  XNOR2_X1 U11934 ( .A(n10048), .B(n12904), .ZN(n14845) );
  OR2_X1 U11935 ( .A1(n14816), .A2(n10051), .ZN(n10050) );
  NAND2_X1 U11936 ( .A1(n10633), .A2(n7429), .ZN(n10049) );
  INV_X1 U11937 ( .A(n15413), .ZN(n15050) );
  INV_X1 U11938 ( .A(n15983), .ZN(n11970) );
  INV_X1 U11939 ( .A(n12773), .ZN(n11930) );
  AND2_X1 U11940 ( .A1(n11160), .A2(n10634), .ZN(n15879) );
  NAND2_X1 U11941 ( .A1(n15898), .A2(n15881), .ZN(n11230) );
  NOR2_X1 U11942 ( .A1(n12729), .A2(n11230), .ZN(n11076) );
  NAND2_X1 U11943 ( .A1(n15916), .A2(n11076), .ZN(n11077) );
  INV_X1 U11944 ( .A(n11701), .ZN(n11455) );
  OR2_X1 U11945 ( .A1(n11868), .A2(n12777), .ZN(n11965) );
  NAND2_X1 U11946 ( .A1(n14686), .A2(n15015), .ZN(n14997) );
  NAND2_X1 U11947 ( .A1(n15403), .A2(n14983), .ZN(n14964) );
  AND2_X1 U11948 ( .A1(n12704), .A2(n15827), .ZN(n10052) );
  AND2_X2 U11949 ( .A1(n10052), .A2(n10051), .ZN(n15878) );
  NAND2_X1 U11950 ( .A1(n10220), .A2(n14842), .ZN(n14826) );
  OAI211_X1 U11951 ( .C1(n10220), .C2(n14842), .A(n15878), .B(n14826), .ZN(
        n14834) );
  NAND2_X1 U11952 ( .A1(n15443), .A2(n10633), .ZN(n12868) );
  INV_X1 U11953 ( .A(n15432), .ZN(n12925) );
  NAND2_X1 U11954 ( .A1(n12925), .A2(P1_B_REG_SCAN_IN), .ZN(n10053) );
  NAND2_X1 U11955 ( .A1(n14704), .A2(n10053), .ZN(n14822) );
  INV_X1 U11956 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10056) );
  NAND2_X1 U11957 ( .A1(n10335), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n10055) );
  NAND2_X1 U11958 ( .A1(n10336), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n10054) );
  OAI211_X1 U11959 ( .C1(n10057), .C2(n10056), .A(n10055), .B(n10054), .ZN(
        n14713) );
  INV_X1 U11960 ( .A(n14713), .ZN(n12857) );
  OR2_X1 U11961 ( .A1(n14822), .A2(n12857), .ZN(n14836) );
  INV_X1 U11962 ( .A(n12868), .ZN(n10088) );
  NAND2_X1 U11963 ( .A1(n14702), .A2(n14715), .ZN(n14838) );
  INV_X1 U11964 ( .A(n10092), .ZN(n12482) );
  NAND2_X1 U11965 ( .A1(n10064), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10065) );
  MUX2_X1 U11966 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10065), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n10067) );
  NAND3_X1 U11967 ( .A1(n12482), .A2(P1_B_REG_SCAN_IN), .A3(n12458), .ZN(
        n10071) );
  INV_X1 U11968 ( .A(P1_B_REG_SCAN_IN), .ZN(n12926) );
  OAI21_X1 U11969 ( .B1(n10068), .B2(n9601), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n10069) );
  AOI21_X1 U11970 ( .B1(n10083), .B2(n12926), .A(n15438), .ZN(n10070) );
  NAND2_X1 U11971 ( .A1(n10071), .A2(n10070), .ZN(n15416) );
  NOR2_X1 U11972 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n10075) );
  NOR4_X1 U11973 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n10074) );
  NOR4_X1 U11974 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n10073) );
  NOR4_X1 U11975 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n10072) );
  NAND4_X1 U11976 ( .A1(n10075), .A2(n10074), .A3(n10073), .A4(n10072), .ZN(
        n10081) );
  NOR4_X1 U11977 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n10079) );
  NOR4_X1 U11978 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n10078) );
  NOR4_X1 U11979 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n10077) );
  NOR4_X1 U11980 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n10076) );
  NAND4_X1 U11981 ( .A1(n10079), .A2(n10078), .A3(n10077), .A4(n10076), .ZN(
        n10080) );
  NOR2_X1 U11982 ( .A1(n10081), .A2(n10080), .ZN(n10082) );
  OR2_X1 U11983 ( .A1(n15416), .A2(n10082), .ZN(n10568) );
  INV_X1 U11984 ( .A(n10324), .ZN(n10086) );
  NAND2_X1 U11985 ( .A1(n14816), .A2(n15827), .ZN(n10087) );
  NAND2_X1 U11986 ( .A1(n10088), .A2(n10087), .ZN(n12924) );
  INV_X1 U11987 ( .A(n12924), .ZN(n10089) );
  NOR2_X1 U11988 ( .A1(n15415), .A2(n10089), .ZN(n10090) );
  AND2_X1 U11989 ( .A1(n10568), .A2(n10090), .ZN(n10797) );
  OR2_X1 U11990 ( .A1(n15416), .A2(P1_D_REG_1__SCAN_IN), .ZN(n10093) );
  OR2_X1 U11991 ( .A1(n10092), .A2(n10091), .ZN(n15418) );
  NAND2_X1 U11992 ( .A1(n10093), .A2(n15418), .ZN(n10795) );
  AND2_X1 U11993 ( .A1(n10797), .A2(n10795), .ZN(n10103) );
  OR2_X1 U11994 ( .A1(n15416), .A2(P1_D_REG_0__SCAN_IN), .ZN(n10094) );
  NAND2_X1 U11995 ( .A1(n12458), .A2(n15438), .ZN(n15419) );
  NAND2_X1 U11996 ( .A1(n10094), .A2(n15419), .ZN(n10796) );
  INV_X1 U11997 ( .A(n10581), .ZN(n10095) );
  NOR2_X1 U11998 ( .A1(n10796), .A2(n10095), .ZN(n10096) );
  OR2_X1 U11999 ( .A1(n10633), .A2(n12703), .ZN(n10098) );
  NAND2_X1 U12000 ( .A1(n12704), .A2(n7429), .ZN(n12912) );
  INV_X1 U12001 ( .A(n12912), .ZN(n10097) );
  NAND2_X1 U12002 ( .A1(n10097), .A2(n10051), .ZN(n10811) );
  NAND2_X1 U12003 ( .A1(n16014), .A2(n15982), .ZN(n15125) );
  NAND2_X1 U12004 ( .A1(n10101), .A2(n10100), .ZN(P1_U3557) );
  AND2_X1 U12005 ( .A1(n10796), .A2(n10581), .ZN(n10102) );
  NAND2_X1 U12006 ( .A1(n10099), .A2(n10105), .ZN(n10106) );
  NAND2_X1 U12007 ( .A1(n10107), .A2(n10106), .ZN(P1_U3525) );
  INV_X1 U12008 ( .A(n14314), .ZN(n14106) );
  OR2_X1 U12009 ( .A1(n10108), .A2(n10642), .ZN(n10713) );
  OR2_X1 U12010 ( .A1(n13932), .A2(n10721), .ZN(n10109) );
  NAND2_X1 U12011 ( .A1(n10241), .A2(n11374), .ZN(n10110) );
  NAND2_X1 U12012 ( .A1(n11415), .A2(n10758), .ZN(n10111) );
  INV_X1 U12013 ( .A(n10756), .ZN(n10112) );
  NAND2_X1 U12014 ( .A1(n11524), .A2(n10785), .ZN(n10113) );
  INV_X1 U12015 ( .A(n10146), .ZN(n10965) );
  NAND2_X1 U12016 ( .A1(n10962), .A2(n10965), .ZN(n10961) );
  NAND2_X1 U12017 ( .A1(n11535), .A2(n11067), .ZN(n10115) );
  NAND2_X1 U12018 ( .A1(n10961), .A2(n10115), .ZN(n11212) );
  OR2_X1 U12019 ( .A1(n11218), .A2(n13926), .ZN(n10116) );
  INV_X1 U12020 ( .A(n11346), .ZN(n11343) );
  INV_X1 U12021 ( .A(n11391), .ZN(n13925) );
  NAND2_X1 U12022 ( .A1(n11387), .A2(n13925), .ZN(n10117) );
  NAND2_X1 U12023 ( .A1(n11657), .A2(n13924), .ZN(n10118) );
  NAND2_X1 U12024 ( .A1(n11742), .A2(n13923), .ZN(n10119) );
  INV_X2 U12025 ( .A(n10157), .ZN(n11779) );
  OR2_X1 U12026 ( .A1(n15965), .A2(n11948), .ZN(n10120) );
  OR2_X1 U12027 ( .A1(n15997), .A2(n12216), .ZN(n10122) );
  INV_X1 U12028 ( .A(n12217), .ZN(n10124) );
  NAND2_X1 U12029 ( .A1(n12218), .A2(n10124), .ZN(n10126) );
  OR2_X1 U12030 ( .A1(n12348), .A2(n12334), .ZN(n10125) );
  NAND2_X1 U12031 ( .A1(n10126), .A2(n10125), .ZN(n12371) );
  NAND2_X1 U12032 ( .A1(n16020), .A2(n12401), .ZN(n10127) );
  OR2_X1 U12033 ( .A1(n14403), .A2(n12441), .ZN(n10128) );
  INV_X1 U12034 ( .A(n14247), .ZN(n14252) );
  NAND2_X1 U12035 ( .A1(n16030), .A2(n14236), .ZN(n10129) );
  NAND2_X1 U12036 ( .A1(n14397), .A2(n14209), .ZN(n10130) );
  NAND2_X1 U12037 ( .A1(n14355), .A2(n14238), .ZN(n10131) );
  NAND2_X1 U12038 ( .A1(n14195), .A2(n14210), .ZN(n10132) );
  NAND2_X1 U12039 ( .A1(n14182), .A2(n14189), .ZN(n10133) );
  NAND2_X1 U12040 ( .A1(n14177), .A2(n10133), .ZN(n14163) );
  OR2_X1 U12041 ( .A1(n14162), .A2(n13817), .ZN(n10134) );
  OR2_X1 U12042 ( .A1(n14149), .A2(n13868), .ZN(n10135) );
  INV_X1 U12043 ( .A(n14116), .ZN(n10177) );
  NAND2_X1 U12044 ( .A1(n14384), .A2(n13898), .ZN(n10136) );
  NAND2_X1 U12045 ( .A1(n14115), .A2(n10136), .ZN(n14108) );
  NAND2_X1 U12046 ( .A1(n10137), .A2(n14076), .ZN(n10236) );
  INV_X1 U12047 ( .A(n16024), .ZN(n10138) );
  NOR2_X1 U12048 ( .A1(n10721), .A2(n11250), .ZN(n10716) );
  AND2_X1 U12049 ( .A1(n11374), .A2(n10716), .ZN(n10744) );
  NAND2_X1 U12050 ( .A1(n11643), .A2(n11397), .ZN(n11398) );
  NOR2_X2 U12051 ( .A1(n9398), .A2(n10183), .ZN(n10834) );
  AOI21_X1 U12052 ( .B1(n14067), .B2(n14060), .A(n14282), .ZN(n10139) );
  NAND2_X1 U12053 ( .A1(n14162), .A2(n13917), .ZN(n10173) );
  OAI22_X1 U12054 ( .A1(n10717), .A2(n10718), .B1(n11503), .B2(n13932), .ZN(
        n10707) );
  INV_X1 U12055 ( .A(n10703), .ZN(n10706) );
  NAND2_X1 U12056 ( .A1(n10707), .A2(n10706), .ZN(n10141) );
  NAND2_X1 U12057 ( .A1(n13876), .A2(n10241), .ZN(n10140) );
  NAND2_X1 U12058 ( .A1(n10141), .A2(n10140), .ZN(n10747) );
  NAND2_X1 U12059 ( .A1(n10747), .A2(n10142), .ZN(n10144) );
  NAND2_X1 U12060 ( .A1(n10750), .A2(n10758), .ZN(n10143) );
  OR2_X1 U12061 ( .A1(n11524), .A2(n13928), .ZN(n10145) );
  NAND2_X1 U12062 ( .A1(n10969), .A2(n11067), .ZN(n10147) );
  NAND2_X1 U12063 ( .A1(n10148), .A2(n10147), .ZN(n11215) );
  INV_X1 U12064 ( .A(n11214), .ZN(n10149) );
  NAND2_X1 U12065 ( .A1(n11215), .A2(n10149), .ZN(n10151) );
  NAND2_X1 U12066 ( .A1(n11218), .A2(n11348), .ZN(n10150) );
  NAND2_X1 U12067 ( .A1(n11387), .A2(n11391), .ZN(n10152) );
  NAND2_X1 U12068 ( .A1(n11643), .A2(n13924), .ZN(n10153) );
  OR2_X1 U12069 ( .A1(n11742), .A2(n11780), .ZN(n10155) );
  OR2_X1 U12070 ( .A1(n11938), .A2(n11591), .ZN(n10158) );
  NOR2_X1 U12071 ( .A1(n15965), .A2(n13921), .ZN(n12013) );
  INV_X1 U12072 ( .A(n12142), .ZN(n10160) );
  NAND2_X1 U12073 ( .A1(n12143), .A2(n10160), .ZN(n10162) );
  NAND2_X1 U12074 ( .A1(n15997), .A2(n12351), .ZN(n10161) );
  AND2_X1 U12075 ( .A1(n12348), .A2(n13919), .ZN(n10163) );
  OR2_X1 U12076 ( .A1(n12348), .A2(n13919), .ZN(n10164) );
  NOR2_X1 U12077 ( .A1(n16020), .A2(n14273), .ZN(n10165) );
  NAND2_X1 U12078 ( .A1(n14403), .A2(n14249), .ZN(n10166) );
  INV_X1 U12079 ( .A(n14236), .ZN(n14276) );
  NAND2_X1 U12080 ( .A1(n16030), .A2(n14276), .ZN(n10168) );
  NAND2_X1 U12081 ( .A1(n14355), .A2(n14188), .ZN(n10170) );
  OR2_X1 U12082 ( .A1(n14182), .A2(n13867), .ZN(n10172) );
  NAND2_X1 U12083 ( .A1(n10173), .A2(n14157), .ZN(n10175) );
  OR2_X1 U12084 ( .A1(n14162), .A2(n13917), .ZN(n10174) );
  NAND2_X1 U12085 ( .A1(n10175), .A2(n10174), .ZN(n14141) );
  INV_X1 U12086 ( .A(n14078), .ZN(n14071) );
  NAND2_X1 U12087 ( .A1(n14070), .A2(n10179), .ZN(n10182) );
  XNOR2_X1 U12088 ( .A(n10182), .B(n10181), .ZN(n10186) );
  NAND2_X1 U12089 ( .A1(n10264), .A2(n10183), .ZN(n10184) );
  INV_X1 U12090 ( .A(P2_B_REG_SCAN_IN), .ZN(n10187) );
  OR2_X1 U12091 ( .A1(n14411), .A2(n10187), .ZN(n10188) );
  NAND2_X1 U12092 ( .A1(n14275), .A2(n10188), .ZN(n14044) );
  OAI22_X1 U12093 ( .A1(n13778), .A2(n14235), .B1(n14044), .B2(n10189), .ZN(
        n10190) );
  NOR4_X1 U12094 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n10196) );
  NOR4_X1 U12095 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n10195) );
  NOR4_X1 U12096 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n10194) );
  NOR4_X1 U12097 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n10193) );
  NAND4_X1 U12098 ( .A1(n10196), .A2(n10195), .A3(n10194), .A4(n10193), .ZN(
        n10204) );
  NOR2_X1 U12099 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n10200) );
  NOR4_X1 U12100 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n10199) );
  NOR4_X1 U12101 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n10198) );
  NOR4_X1 U12102 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n10197) );
  NAND4_X1 U12103 ( .A1(n10200), .A2(n10199), .A3(n10198), .A4(n10197), .ZN(
        n10203) );
  XNOR2_X1 U12104 ( .A(n12459), .B(P2_B_REG_SCAN_IN), .ZN(n10201) );
  AND2_X1 U12105 ( .A1(n12480), .A2(n10201), .ZN(n10202) );
  INV_X1 U12106 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15449) );
  NAND2_X1 U12107 ( .A1(n15450), .A2(n15449), .ZN(n10206) );
  NAND2_X1 U12108 ( .A1(n14417), .A2(n12480), .ZN(n10205) );
  AND2_X1 U12109 ( .A1(n10206), .A2(n10205), .ZN(n10260) );
  NAND2_X1 U12110 ( .A1(n14151), .A2(n12085), .ZN(n10265) );
  NAND2_X1 U12111 ( .A1(n10439), .A2(n10210), .ZN(n11239) );
  AND2_X1 U12112 ( .A1(n10265), .A2(n11239), .ZN(n10207) );
  NAND2_X1 U12113 ( .A1(n14417), .A2(n12459), .ZN(n10208) );
  NAND2_X1 U12114 ( .A1(n10834), .A2(n10210), .ZN(n16029) );
  INV_X1 U12115 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n10211) );
  OAI21_X1 U12116 ( .B1(n7594), .B2(n14402), .A(n10212), .ZN(n10213) );
  INV_X1 U12117 ( .A(n10213), .ZN(n10214) );
  INV_X1 U12118 ( .A(n15454), .ZN(n10251) );
  NAND2_X1 U12119 ( .A1(n16035), .A2(n14347), .ZN(n14369) );
  NAND2_X1 U12120 ( .A1(n10218), .A2(n9981), .ZN(n10219) );
  NAND2_X1 U12121 ( .A1(n7190), .A2(n10219), .ZN(n14858) );
  AOI211_X1 U12122 ( .C1(n14599), .C2(n14865), .A(n15985), .B(n10220), .ZN(
        n14854) );
  INV_X1 U12123 ( .A(n14854), .ZN(n10227) );
  INV_X1 U12124 ( .A(n10221), .ZN(n10224) );
  AND3_X1 U12125 ( .A1(n14860), .A2(n12901), .A3(n10222), .ZN(n10223) );
  OAI21_X1 U12126 ( .B1(n10224), .B2(n10223), .A(n16013), .ZN(n10225) );
  AOI22_X1 U12127 ( .A1(n14714), .A2(n14704), .B1(n14702), .B2(n14716), .ZN(
        n14596) );
  NAND2_X1 U12128 ( .A1(n14599), .A2(n10105), .ZN(n10232) );
  AND2_X1 U12129 ( .A1(n10438), .A2(n10233), .ZN(n10437) );
  INV_X1 U12130 ( .A(n10583), .ZN(n10570) );
  INV_X1 U12131 ( .A(n13710), .ZN(n10234) );
  INV_X2 U12132 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NAND2_X1 U12133 ( .A1(n13932), .A2(n14282), .ZN(n10237) );
  OAI22_X1 U12134 ( .A1(n10713), .A2(n14151), .B1(n11250), .B2(n13805), .ZN(
        n10542) );
  NAND2_X1 U12135 ( .A1(n10238), .A2(n10237), .ZN(n10239) );
  NAND2_X1 U12136 ( .A1(n10540), .A2(n10239), .ZN(n13878) );
  XNOR2_X1 U12137 ( .A(n11374), .B(n13773), .ZN(n10242) );
  OR2_X1 U12138 ( .A1(n10241), .A2(n14151), .ZN(n10243) );
  XNOR2_X1 U12139 ( .A(n10242), .B(n10243), .ZN(n13879) );
  INV_X1 U12140 ( .A(n10242), .ZN(n10244) );
  NAND2_X1 U12141 ( .A1(n10244), .A2(n10243), .ZN(n10245) );
  XNOR2_X1 U12142 ( .A(n11415), .B(n13773), .ZN(n10246) );
  NAND2_X1 U12143 ( .A1(n10246), .A2(n10247), .ZN(n10782) );
  INV_X1 U12144 ( .A(n10246), .ZN(n10249) );
  INV_X1 U12145 ( .A(n10247), .ZN(n10248) );
  NAND2_X1 U12146 ( .A1(n10249), .A2(n10248), .ZN(n10250) );
  NAND2_X1 U12147 ( .A1(n10782), .A2(n10250), .ZN(n10257) );
  AND3_X1 U12148 ( .A1(n10251), .A2(n15455), .A3(n10260), .ZN(n10252) );
  AND2_X1 U12149 ( .A1(n10259), .A2(n10252), .ZN(n10268) );
  INV_X1 U12150 ( .A(n10439), .ZN(n10253) );
  AND2_X1 U12151 ( .A1(n16029), .A2(n10253), .ZN(n10254) );
  AOI211_X1 U12152 ( .C1(n10258), .C2(n10257), .A(n13907), .B(n10256), .ZN(
        n10271) );
  NAND2_X1 U12153 ( .A1(n10260), .A2(n10259), .ZN(n11238) );
  OAI21_X1 U12154 ( .B1(n15454), .B2(n11238), .A(n10265), .ZN(n10263) );
  AND3_X1 U12155 ( .A1(n11239), .A2(n10438), .A3(n10261), .ZN(n10262) );
  NAND2_X1 U12156 ( .A1(n10263), .A2(n10262), .ZN(n10544) );
  MUX2_X1 U12157 ( .A(n13856), .B(P2_U3088), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n10270) );
  AND2_X1 U12158 ( .A1(n10834), .A2(n10264), .ZN(n11249) );
  NAND2_X1 U12159 ( .A1(n10268), .A2(n11249), .ZN(n10266) );
  AOI22_X1 U12160 ( .A1(n14274), .A2(n13931), .B1(n13928), .B2(n14275), .ZN(
        n10748) );
  NAND2_X1 U12161 ( .A1(n10268), .A2(n10267), .ZN(n13900) );
  OAI22_X1 U12162 ( .A1(n13889), .A2(n11415), .B1(n10748), .B2(n13900), .ZN(
        n10269) );
  OR3_X1 U12163 ( .A1(n10271), .A2(n10270), .A3(n10269), .ZN(P2_U3190) );
  INV_X1 U12164 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10862) );
  NAND2_X1 U12165 ( .A1(n10272), .A2(P3_U3151), .ZN(n10273) );
  OAI21_X1 U12166 ( .B1(n10862), .B2(P3_U3151), .A(n10273), .ZN(P3_U3295) );
  NOR2_X1 U12167 ( .A1(n10297), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13717) );
  INV_X2 U12168 ( .A(n13717), .ZN(n13730) );
  OAI222_X1 U12169 ( .A1(P3_U3151), .A2(n11274), .B1(n13730), .B2(n10274), 
        .C1(n8049), .C2(n13723), .ZN(P3_U3294) );
  OAI222_X1 U12170 ( .A1(P3_U3151), .A2(n10991), .B1(n13730), .B2(n10275), 
        .C1(n15278), .C2(n13723), .ZN(P3_U3289) );
  AND2_X1 U12171 ( .A1(n10276), .A2(P1_U3086), .ZN(n15439) );
  INV_X2 U12172 ( .A(n15439), .ZN(n15437) );
  INV_X1 U12173 ( .A(n10277), .ZN(n10311) );
  OAI222_X1 U12174 ( .A1(n15435), .A2(n10278), .B1(n15437), .B2(n10311), .C1(
        n10681), .C2(P1_U3086), .ZN(P1_U3353) );
  OAI222_X1 U12175 ( .A1(P3_U3151), .A2(n11825), .B1(n13723), .B2(n15207), 
        .C1(n13730), .C2(n10279), .ZN(P3_U3287) );
  INV_X1 U12176 ( .A(n15780), .ZN(n11828) );
  INV_X1 U12177 ( .A(SI_9_), .ZN(n15320) );
  INV_X1 U12178 ( .A(n10280), .ZN(n10281) );
  OAI222_X1 U12179 ( .A1(P3_U3151), .A2(n11828), .B1(n13723), .B2(n15320), 
        .C1(n13730), .C2(n10281), .ZN(P3_U3286) );
  INV_X1 U12180 ( .A(n11808), .ZN(n11820) );
  INV_X1 U12181 ( .A(SI_7_), .ZN(n10284) );
  INV_X1 U12182 ( .A(n10282), .ZN(n10283) );
  OAI222_X1 U12183 ( .A1(P3_U3151), .A2(n11820), .B1(n13723), .B2(n10284), 
        .C1(n13730), .C2(n10283), .ZN(P3_U3288) );
  INV_X1 U12184 ( .A(SI_10_), .ZN(n15321) );
  OAI222_X1 U12185 ( .A1(P3_U3151), .A2(n11830), .B1(n13723), .B2(n15321), 
        .C1(n13730), .C2(n10285), .ZN(P3_U3285) );
  INV_X1 U12186 ( .A(n10885), .ZN(n11038) );
  INV_X1 U12187 ( .A(n10286), .ZN(n10287) );
  OAI222_X1 U12188 ( .A1(n11038), .A2(P3_U3151), .B1(n13730), .B2(n10287), 
        .C1(n7319), .C2(n13723), .ZN(P3_U3293) );
  INV_X1 U12189 ( .A(n10288), .ZN(n10289) );
  INV_X1 U12190 ( .A(SI_5_), .ZN(n15206) );
  OAI222_X1 U12191 ( .A1(n11206), .A2(P3_U3151), .B1(n13730), .B2(n10289), 
        .C1(n15206), .C2(n13723), .ZN(P3_U3290) );
  INV_X1 U12192 ( .A(n10891), .ZN(n10949) );
  INV_X1 U12193 ( .A(n10290), .ZN(n10292) );
  INV_X1 U12194 ( .A(SI_3_), .ZN(n10291) );
  OAI222_X1 U12195 ( .A1(n10949), .A2(P3_U3151), .B1(n13730), .B2(n10292), 
        .C1(n10291), .C2(n13723), .ZN(P3_U3292) );
  INV_X1 U12196 ( .A(n10985), .ZN(n10902) );
  INV_X1 U12197 ( .A(n10293), .ZN(n10294) );
  INV_X1 U12198 ( .A(SI_4_), .ZN(n15323) );
  OAI222_X1 U12199 ( .A1(n10902), .A2(P3_U3151), .B1(n13730), .B2(n10294), 
        .C1(n15323), .C2(n13723), .ZN(P3_U3291) );
  OAI222_X1 U12200 ( .A1(n11814), .A2(P3_U3151), .B1(n13730), .B2(n10295), 
        .C1(n13723), .C2(n15275), .ZN(P3_U3284) );
  NAND2_X1 U12201 ( .A1(n10297), .A2(P2_U3088), .ZN(n12358) );
  INV_X1 U12202 ( .A(n10296), .ZN(n10301) );
  NOR2_X1 U12203 ( .A1(n10297), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12961) );
  INV_X2 U12204 ( .A(n12961), .ZN(n14422) );
  OAI222_X1 U12205 ( .A1(P2_U3088), .A2(n13940), .B1(n12358), .B2(n10301), 
        .C1(n10298), .C2(n14422), .ZN(P2_U3323) );
  OAI222_X1 U12206 ( .A1(n12114), .A2(P3_U3151), .B1(n13730), .B2(n10299), 
        .C1(n13723), .C2(n15172), .ZN(P3_U3283) );
  OAI222_X1 U12207 ( .A1(P1_U3086), .A2(n14745), .B1(n15437), .B2(n10305), 
        .C1(n8804), .C2(n15435), .ZN(P1_U3354) );
  INV_X1 U12208 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10300) );
  OAI222_X1 U12209 ( .A1(P1_U3086), .A2(n10668), .B1(n15437), .B2(n10301), 
        .C1(n10300), .C2(n15435), .ZN(P1_U3351) );
  INV_X1 U12210 ( .A(n14760), .ZN(n10360) );
  INV_X1 U12211 ( .A(n10302), .ZN(n10307) );
  INV_X1 U12212 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10303) );
  OAI222_X1 U12213 ( .A1(P1_U3086), .A2(n10360), .B1(n15437), .B2(n10307), 
        .C1(n10303), .C2(n15435), .ZN(P1_U3352) );
  INV_X1 U12214 ( .A(n14419), .ZN(n14416) );
  OAI222_X1 U12215 ( .A1(n14416), .A2(n10305), .B1(n14422), .B2(n10304), .C1(
        P2_U3088), .C2(n15461), .ZN(P2_U3326) );
  AOI22_X1 U12216 ( .A1(n15473), .A2(P2_STATE_REG_SCAN_IN), .B1(n12961), .B2(
        P1_DATAO_REG_3__SCAN_IN), .ZN(n10306) );
  OAI21_X1 U12217 ( .B1(n10307), .B2(n14416), .A(n10306), .ZN(P2_U3324) );
  INV_X1 U12218 ( .A(n10308), .ZN(n10313) );
  AOI22_X1 U12219 ( .A1(n13954), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n12961), .ZN(n10309) );
  OAI21_X1 U12220 ( .B1(n10313), .B2(n12358), .A(n10309), .ZN(P2_U3322) );
  INV_X1 U12221 ( .A(n10496), .ZN(n10469) );
  OAI222_X1 U12222 ( .A1(P2_U3088), .A2(n10469), .B1(n14416), .B2(n10311), 
        .C1(n10310), .C2(n14422), .ZN(P2_U3325) );
  INV_X1 U12223 ( .A(n10375), .ZN(n10390) );
  INV_X1 U12224 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10312) );
  OAI222_X1 U12225 ( .A1(P1_U3086), .A2(n10390), .B1(n15437), .B2(n10313), 
        .C1(n10312), .C2(n15435), .ZN(P1_U3350) );
  INV_X1 U12226 ( .A(n10314), .ZN(n10317) );
  INV_X1 U12227 ( .A(n10391), .ZN(n14775) );
  OAI222_X1 U12228 ( .A1(n15435), .A2(n10315), .B1(n15437), .B2(n10317), .C1(
        P1_U3086), .C2(n14775), .ZN(P1_U3349) );
  INV_X1 U12229 ( .A(n13969), .ZN(n10316) );
  OAI222_X1 U12230 ( .A1(n14422), .A2(n10318), .B1(n14416), .B2(n10317), .C1(
        P2_U3088), .C2(n10316), .ZN(P2_U3321) );
  INV_X1 U12231 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10320) );
  INV_X1 U12232 ( .A(n13984), .ZN(n10319) );
  OAI222_X1 U12233 ( .A1(n14422), .A2(n10320), .B1(n12358), .B2(n10321), .C1(
        n10319), .C2(P2_U3088), .ZN(P2_U3320) );
  INV_X1 U12234 ( .A(n10407), .ZN(n10405) );
  OAI222_X1 U12235 ( .A1(n15435), .A2(n10322), .B1(n15437), .B2(n10321), .C1(
        n10405), .C2(P1_U3086), .ZN(P1_U3348) );
  NAND2_X1 U12236 ( .A1(n10324), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15440) );
  NAND2_X1 U12237 ( .A1(n15415), .A2(n15440), .ZN(n10327) );
  OAI21_X1 U12238 ( .B1(n12868), .B2(n10324), .A(n10323), .ZN(n10325) );
  AND2_X1 U12239 ( .A1(n10327), .A2(n10325), .ZN(n15544) );
  NOR2_X1 U12240 ( .A1(n15544), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12241 ( .A(n10325), .ZN(n10326) );
  NAND2_X1 U12242 ( .A1(n10327), .A2(n10326), .ZN(n10355) );
  INV_X1 U12243 ( .A(n10355), .ZN(n10330) );
  NAND3_X1 U12244 ( .A1(n15566), .A2(P1_IR_REG_0__SCAN_IN), .A3(n10574), .ZN(
        n10332) );
  OAI21_X1 U12245 ( .B1(n15432), .B2(P1_REG2_REG_0__SCAN_IN), .A(n10353), .ZN(
        n10656) );
  AOI21_X1 U12246 ( .B1(n15432), .B2(n10574), .A(n10656), .ZN(n10328) );
  MUX2_X1 U12247 ( .A(n10656), .B(n10328), .S(n10657), .Z(n10329) );
  AOI22_X1 U12248 ( .A1(n10330), .A2(n10329), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10331) );
  OAI211_X1 U12249 ( .C1(n15570), .C2(n7607), .A(n10332), .B(n10331), .ZN(
        P1_U3243) );
  OAI222_X1 U12250 ( .A1(n12182), .A2(P3_U3151), .B1(n13730), .B2(n10333), 
        .C1(n15318), .C2(n13723), .ZN(P3_U3282) );
  NAND2_X1 U12251 ( .A1(n12351), .A2(P2_U3947), .ZN(n10334) );
  OAI21_X1 U12252 ( .B1(n10765), .B2(P2_U3947), .A(n10334), .ZN(P2_U3544) );
  INV_X1 U12253 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n12493) );
  INV_X1 U12254 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n15161) );
  NAND2_X1 U12255 ( .A1(n10335), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n10338) );
  NAND2_X1 U12256 ( .A1(n10336), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n10337) );
  OAI211_X1 U12257 ( .C1(n10057), .C2(n15161), .A(n10338), .B(n10337), .ZN(
        n12866) );
  NAND2_X1 U12258 ( .A1(P1_U4016), .A2(n12866), .ZN(n10339) );
  OAI21_X1 U12259 ( .B1(P1_U4016), .B2(n12493), .A(n10339), .ZN(P1_U3591) );
  NAND2_X1 U12260 ( .A1(P1_U4016), .A2(n10632), .ZN(n10340) );
  OAI21_X1 U12261 ( .B1(P1_U4016), .B2(n8807), .A(n10340), .ZN(P1_U3560) );
  MUX2_X1 U12262 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9689), .S(n10375), .Z(
        n10352) );
  MUX2_X1 U12263 ( .A(n9632), .B(P1_REG1_REG_1__SCAN_IN), .S(n14745), .Z(
        n14751) );
  AND2_X1 U12264 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14752) );
  NAND2_X1 U12265 ( .A1(n14751), .A2(n14752), .ZN(n14750) );
  NAND2_X1 U12266 ( .A1(n14753), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10341) );
  NAND2_X1 U12267 ( .A1(n14750), .A2(n10341), .ZN(n10675) );
  INV_X1 U12268 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10342) );
  MUX2_X1 U12269 ( .A(n10342), .B(P1_REG1_REG_2__SCAN_IN), .S(n10681), .Z(
        n10343) );
  NAND2_X1 U12270 ( .A1(n10675), .A2(n10343), .ZN(n14763) );
  NAND2_X1 U12271 ( .A1(n10358), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n14762) );
  NAND2_X1 U12272 ( .A1(n14763), .A2(n14762), .ZN(n10346) );
  MUX2_X1 U12273 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10344), .S(n14760), .Z(
        n10345) );
  NAND2_X1 U12274 ( .A1(n10346), .A2(n10345), .ZN(n14765) );
  NAND2_X1 U12275 ( .A1(n14760), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n10658) );
  NAND2_X1 U12276 ( .A1(n14765), .A2(n10658), .ZN(n10349) );
  MUX2_X1 U12277 ( .A(n10347), .B(P1_REG1_REG_4__SCAN_IN), .S(n10668), .Z(
        n10348) );
  NAND2_X1 U12278 ( .A1(n10349), .A2(n10348), .ZN(n10661) );
  NAND2_X1 U12279 ( .A1(n10361), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10350) );
  AND2_X1 U12280 ( .A1(n10661), .A2(n10350), .ZN(n10351) );
  NAND2_X1 U12281 ( .A1(n10351), .A2(n10352), .ZN(n10377) );
  OAI21_X1 U12282 ( .B1(n10352), .B2(n10351), .A(n10377), .ZN(n10366) );
  NAND2_X1 U12283 ( .A1(n12925), .A2(n10353), .ZN(n10354) );
  OR2_X1 U12284 ( .A1(n10355), .A2(n10354), .ZN(n14811) );
  INV_X1 U12285 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n11159) );
  MUX2_X1 U12286 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n11159), .S(n14745), .Z(
        n10357) );
  NOR3_X1 U12287 ( .A1(n10357), .A2(n10356), .A3(n10657), .ZN(n14746) );
  AOI21_X1 U12288 ( .B1(n14753), .B2(P1_REG2_REG_1__SCAN_IN), .A(n14746), .ZN(
        n10674) );
  MUX2_X1 U12289 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9621), .S(n10681), .Z(
        n10673) );
  OR2_X1 U12290 ( .A1(n10674), .A2(n10673), .ZN(n14769) );
  NAND2_X1 U12291 ( .A1(n10358), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14768) );
  MUX2_X1 U12292 ( .A(n10359), .B(P1_REG2_REG_3__SCAN_IN), .S(n14760), .Z(
        n14767) );
  AOI21_X1 U12293 ( .B1(n14769), .B2(n14768), .A(n14767), .ZN(n14766) );
  NOR2_X1 U12294 ( .A1(n10360), .A2(n10359), .ZN(n10664) );
  MUX2_X1 U12295 ( .A(n11116), .B(P1_REG2_REG_4__SCAN_IN), .S(n10668), .Z(
        n10663) );
  OAI21_X1 U12296 ( .B1(n14766), .B2(n10664), .A(n10663), .ZN(n10662) );
  NAND2_X1 U12297 ( .A1(n10361), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10363) );
  MUX2_X1 U12298 ( .A(n10389), .B(P1_REG2_REG_5__SCAN_IN), .S(n10375), .Z(
        n10362) );
  AOI21_X1 U12299 ( .B1(n10662), .B2(n10363), .A(n10362), .ZN(n14783) );
  AND3_X1 U12300 ( .A1(n10662), .A2(n10363), .A3(n10362), .ZN(n10364) );
  NOR3_X1 U12301 ( .A1(n14811), .A2(n14783), .A3(n10364), .ZN(n10365) );
  AOI21_X1 U12302 ( .B1(n15566), .B2(n10366), .A(n10365), .ZN(n10369) );
  NAND2_X1 U12303 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10930) );
  INV_X1 U12304 ( .A(n10930), .ZN(n10367) );
  AOI21_X1 U12305 ( .B1(n15544), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10367), .ZN(
        n10368) );
  OAI211_X1 U12306 ( .C1(n10390), .C2(n15564), .A(n10369), .B(n10368), .ZN(
        P1_U3248) );
  OAI222_X1 U12307 ( .A1(P1_U3086), .A2(n10392), .B1(n15437), .B2(n10372), 
        .C1(n10370), .C2(n15435), .ZN(P1_U3347) );
  INV_X1 U12308 ( .A(n14000), .ZN(n10373) );
  INV_X1 U12309 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10371) );
  OAI222_X1 U12310 ( .A1(P2_U3088), .A2(n10373), .B1(n14416), .B2(n10372), 
        .C1(n10371), .C2(n14422), .ZN(P2_U3319) );
  OAI222_X1 U12311 ( .A1(n13263), .A2(P3_U3151), .B1(n13730), .B2(n10374), 
        .C1(n13723), .C2(n15315), .ZN(P3_U3281) );
  OR2_X1 U12312 ( .A1(n10375), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n10376) );
  AND2_X1 U12313 ( .A1(n10377), .A2(n10376), .ZN(n14780) );
  INV_X1 U12314 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10378) );
  MUX2_X1 U12315 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10378), .S(n10391), .Z(
        n14779) );
  NAND2_X1 U12316 ( .A1(n14780), .A2(n14779), .ZN(n14778) );
  NAND2_X1 U12317 ( .A1(n10391), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10409) );
  NAND2_X1 U12318 ( .A1(n14778), .A2(n10409), .ZN(n10381) );
  INV_X1 U12319 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10379) );
  MUX2_X1 U12320 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n10379), .S(n10407), .Z(
        n10380) );
  NAND2_X1 U12321 ( .A1(n10381), .A2(n10380), .ZN(n10411) );
  NAND2_X1 U12322 ( .A1(n10407), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10382) );
  NAND2_X1 U12323 ( .A1(n10411), .A2(n10382), .ZN(n10417) );
  MUX2_X1 U12324 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10383), .S(n10392), .Z(
        n10418) );
  NAND2_X1 U12325 ( .A1(n10392), .A2(n10383), .ZN(n10386) );
  NAND2_X1 U12326 ( .A1(n10415), .A2(n10386), .ZN(n10384) );
  MUX2_X1 U12327 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9745), .S(n10432), .Z(
        n10385) );
  NAND2_X1 U12328 ( .A1(n10384), .A2(n10385), .ZN(n10558) );
  INV_X1 U12329 ( .A(n10385), .ZN(n10387) );
  NAND3_X1 U12330 ( .A1(n10415), .A2(n10387), .A3(n10386), .ZN(n10388) );
  AND2_X1 U12331 ( .A1(n10558), .A2(n10388), .ZN(n10401) );
  NOR2_X1 U12332 ( .A1(n10390), .A2(n10389), .ZN(n14782) );
  MUX2_X1 U12333 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10809), .S(n10391), .Z(
        n14781) );
  OAI21_X1 U12334 ( .B1(n14783), .B2(n14782), .A(n14781), .ZN(n14785) );
  NAND2_X1 U12335 ( .A1(n10391), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10403) );
  MUX2_X1 U12336 ( .A(n11357), .B(P1_REG2_REG_7__SCAN_IN), .S(n10407), .Z(
        n10402) );
  AOI21_X1 U12337 ( .B1(n14785), .B2(n10403), .A(n10402), .ZN(n10423) );
  NOR2_X1 U12338 ( .A1(n10405), .A2(n11357), .ZN(n10422) );
  MUX2_X1 U12339 ( .A(n10393), .B(P1_REG2_REG_8__SCAN_IN), .S(n10392), .Z(
        n10421) );
  OAI21_X1 U12340 ( .B1(n10423), .B2(n10422), .A(n10421), .ZN(n10420) );
  NAND2_X1 U12341 ( .A1(n10428), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10395) );
  MUX2_X1 U12342 ( .A(n9750), .B(P1_REG2_REG_9__SCAN_IN), .S(n10432), .Z(
        n10394) );
  AOI21_X1 U12343 ( .B1(n10420), .B2(n10395), .A(n10394), .ZN(n10553) );
  INV_X1 U12344 ( .A(n10553), .ZN(n10397) );
  INV_X1 U12345 ( .A(n14811), .ZN(n15558) );
  NAND3_X1 U12346 ( .A1(n10420), .A2(n10395), .A3(n10394), .ZN(n10396) );
  NAND3_X1 U12347 ( .A1(n10397), .A2(n15558), .A3(n10396), .ZN(n10400) );
  INV_X1 U12348 ( .A(n15564), .ZN(n15548) );
  AND2_X1 U12349 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n12039) );
  NOR2_X1 U12350 ( .A1(n15570), .A2(n15642), .ZN(n10398) );
  AOI211_X1 U12351 ( .C1(n15548), .C2(n10432), .A(n12039), .B(n10398), .ZN(
        n10399) );
  OAI211_X1 U12352 ( .C1(n10401), .C2(n11897), .A(n10400), .B(n10399), .ZN(
        P1_U3252) );
  NAND3_X1 U12353 ( .A1(n14785), .A2(n10403), .A3(n10402), .ZN(n10404) );
  NAND2_X1 U12354 ( .A1(n10404), .A2(n15558), .ZN(n10414) );
  AND2_X1 U12355 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n11495) );
  NOR2_X1 U12356 ( .A1(n15564), .A2(n10405), .ZN(n10406) );
  AOI211_X1 U12357 ( .C1(n15544), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n11495), .B(
        n10406), .ZN(n10413) );
  MUX2_X1 U12358 ( .A(n10379), .B(P1_REG1_REG_7__SCAN_IN), .S(n10407), .Z(
        n10408) );
  NAND3_X1 U12359 ( .A1(n14778), .A2(n10409), .A3(n10408), .ZN(n10410) );
  NAND3_X1 U12360 ( .A1(n15566), .A2(n10411), .A3(n10410), .ZN(n10412) );
  OAI211_X1 U12361 ( .C1(n10423), .C2(n10414), .A(n10413), .B(n10412), .ZN(
        P1_U3250) );
  INV_X1 U12362 ( .A(n10415), .ZN(n10416) );
  AOI21_X1 U12363 ( .B1(n10418), .B2(n10417), .A(n10416), .ZN(n10430) );
  NAND2_X1 U12364 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n10419) );
  OAI21_X1 U12365 ( .B1(n15570), .B2(n15637), .A(n10419), .ZN(n10427) );
  INV_X1 U12366 ( .A(n10420), .ZN(n10425) );
  NOR3_X1 U12367 ( .A1(n10423), .A2(n10422), .A3(n10421), .ZN(n10424) );
  NOR3_X1 U12368 ( .A1(n10425), .A2(n10424), .A3(n14811), .ZN(n10426) );
  AOI211_X1 U12369 ( .C1(n15548), .C2(n10428), .A(n10427), .B(n10426), .ZN(
        n10429) );
  OAI21_X1 U12370 ( .B1(n10430), .B2(n11897), .A(n10429), .ZN(P1_U3251) );
  INV_X1 U12371 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10431) );
  INV_X1 U12372 ( .A(n10530), .ZN(n10535) );
  OAI222_X1 U12373 ( .A1(n14422), .A2(n10431), .B1(n14416), .B2(n10433), .C1(
        n10535), .C2(P2_U3088), .ZN(P2_U3318) );
  INV_X1 U12374 ( .A(n10432), .ZN(n10556) );
  OAI222_X1 U12375 ( .A1(n15435), .A2(n10434), .B1(n15437), .B2(n10433), .C1(
        n10556), .C2(P1_U3086), .ZN(P1_U3346) );
  OAI222_X1 U12376 ( .A1(n13285), .A2(P3_U3151), .B1(n13730), .B2(n10435), 
        .C1(n13723), .C2(n15313), .ZN(P3_U3280) );
  AND2_X1 U12377 ( .A1(n10638), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U12378 ( .A1(n10638), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U12379 ( .A1(n10638), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U12380 ( .A1(n10638), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U12381 ( .A1(n10638), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U12382 ( .A1(n10638), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U12383 ( .A1(n10638), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U12384 ( .A1(n10638), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U12385 ( .A1(n10638), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U12386 ( .A1(n10638), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U12387 ( .A1(n10638), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U12388 ( .A1(n10638), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U12389 ( .A1(n10638), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U12390 ( .A1(n10638), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U12391 ( .A1(n10638), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U12392 ( .A1(n10638), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U12393 ( .A1(n10638), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  INV_X1 U12394 ( .A(n15435), .ZN(n15423) );
  AOI22_X1 U12395 ( .A1(n10599), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n15423), .ZN(n10436) );
  OAI21_X1 U12396 ( .B1(n10471), .B2(n15437), .A(n10436), .ZN(P1_U3345) );
  INV_X1 U12397 ( .A(n10437), .ZN(n10442) );
  NAND2_X1 U12398 ( .A1(n10439), .A2(n10438), .ZN(n10440) );
  NAND2_X1 U12399 ( .A1(n10440), .A2(n8802), .ZN(n10441) );
  NAND2_X1 U12400 ( .A1(n10442), .A2(n10441), .ZN(n10455) );
  AND2_X1 U12401 ( .A1(n10443), .A2(n10455), .ZN(n15460) );
  INV_X1 U12402 ( .A(n15521), .ZN(n12095) );
  INV_X1 U12403 ( .A(n15534), .ZN(n15501) );
  NAND2_X1 U12404 ( .A1(n10444), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14407) );
  NOR2_X1 U12405 ( .A1(n14407), .A2(n10445), .ZN(n10446) );
  NAND2_X1 U12406 ( .A1(n10455), .A2(n10446), .ZN(n15488) );
  INV_X1 U12407 ( .A(n15488), .ZN(n15527) );
  MUX2_X1 U12408 ( .A(n10447), .B(P2_REG1_REG_1__SCAN_IN), .S(n15461), .Z(
        n15467) );
  AND2_X1 U12409 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n15468) );
  NAND2_X1 U12410 ( .A1(n15467), .A2(n15468), .ZN(n15466) );
  NAND2_X1 U12411 ( .A1(n10457), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10452) );
  NAND2_X1 U12412 ( .A1(n15466), .A2(n10452), .ZN(n10450) );
  INV_X1 U12413 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10448) );
  MUX2_X1 U12414 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n10448), .S(n10496), .Z(
        n10449) );
  NAND2_X1 U12415 ( .A1(n10450), .A2(n10449), .ZN(n10498) );
  MUX2_X1 U12416 ( .A(n10448), .B(P2_REG1_REG_2__SCAN_IN), .S(n10496), .Z(
        n10451) );
  NAND3_X1 U12417 ( .A1(n15466), .A2(n10452), .A3(n10451), .ZN(n10453) );
  AND3_X1 U12418 ( .A1(n15527), .A2(n10498), .A3(n10453), .ZN(n10467) );
  NOR2_X1 U12419 ( .A1(n14407), .A2(n14411), .ZN(n10454) );
  NAND2_X1 U12420 ( .A1(n10455), .A2(n10454), .ZN(n15502) );
  MUX2_X1 U12421 ( .A(n10456), .B(P2_REG2_REG_1__SCAN_IN), .S(n15461), .Z(
        n15464) );
  AND2_X1 U12422 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n15465) );
  NAND2_X1 U12423 ( .A1(n15464), .A2(n15465), .ZN(n15463) );
  NAND2_X1 U12424 ( .A1(n10457), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10462) );
  NAND2_X1 U12425 ( .A1(n15463), .A2(n10462), .ZN(n10460) );
  MUX2_X1 U12426 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10458), .S(n10496), .Z(
        n10459) );
  NAND2_X1 U12427 ( .A1(n10460), .A2(n10459), .ZN(n10475) );
  MUX2_X1 U12428 ( .A(n10458), .B(P2_REG2_REG_2__SCAN_IN), .S(n10496), .Z(
        n10461) );
  NAND3_X1 U12429 ( .A1(n15463), .A2(n10462), .A3(n10461), .ZN(n10463) );
  NAND3_X1 U12430 ( .A1(n15523), .A2(n10475), .A3(n10463), .ZN(n10464) );
  OAI21_X1 U12431 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n10465), .A(n10464), .ZN(
        n10466) );
  AOI211_X1 U12432 ( .C1(n15501), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n10467), .B(
        n10466), .ZN(n10468) );
  OAI21_X1 U12433 ( .B1(n10469), .B2(n12095), .A(n10468), .ZN(P2_U3216) );
  INV_X1 U12434 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10472) );
  INV_X1 U12435 ( .A(n11137), .ZN(n10470) );
  OAI222_X1 U12436 ( .A1(n14422), .A2(n10472), .B1(n14416), .B2(n10471), .C1(
        n10470), .C2(P2_U3088), .ZN(P2_U3317) );
  INV_X1 U12437 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10473) );
  NAND2_X1 U12438 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n11880)
         );
  OAI21_X1 U12439 ( .B1(n15534), .B2(n10473), .A(n11880), .ZN(n10495) );
  NAND2_X1 U12440 ( .A1(n10496), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10474) );
  NAND2_X1 U12441 ( .A1(n10475), .A2(n10474), .ZN(n15482) );
  MUX2_X1 U12442 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10476), .S(n15473), .Z(
        n15481) );
  NAND2_X1 U12443 ( .A1(n15482), .A2(n15481), .ZN(n15480) );
  NAND2_X1 U12444 ( .A1(n15473), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n13937) );
  NAND2_X1 U12445 ( .A1(n15480), .A2(n13937), .ZN(n10478) );
  MUX2_X1 U12446 ( .A(n11522), .B(P2_REG2_REG_4__SCAN_IN), .S(n13940), .Z(
        n10477) );
  NAND2_X1 U12447 ( .A1(n10478), .A2(n10477), .ZN(n13952) );
  NAND2_X1 U12448 ( .A1(n13936), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n13951) );
  NAND2_X1 U12449 ( .A1(n13952), .A2(n13951), .ZN(n10480) );
  INV_X1 U12450 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11533) );
  MUX2_X1 U12451 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11533), .S(n13954), .Z(
        n10479) );
  NAND2_X1 U12452 ( .A1(n10480), .A2(n10479), .ZN(n13972) );
  NAND2_X1 U12453 ( .A1(n13954), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n13971) );
  NAND2_X1 U12454 ( .A1(n13972), .A2(n13971), .ZN(n10483) );
  MUX2_X1 U12455 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10481), .S(n13969), .Z(
        n10482) );
  NAND2_X1 U12456 ( .A1(n10483), .A2(n10482), .ZN(n13987) );
  NAND2_X1 U12457 ( .A1(n13969), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n13986) );
  NAND2_X1 U12458 ( .A1(n13987), .A2(n13986), .ZN(n10485) );
  INV_X1 U12459 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11551) );
  MUX2_X1 U12460 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11551), .S(n13984), .Z(
        n10484) );
  NAND2_X1 U12461 ( .A1(n10485), .A2(n10484), .ZN(n14003) );
  NAND2_X1 U12462 ( .A1(n13984), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n14002) );
  NAND2_X1 U12463 ( .A1(n14003), .A2(n14002), .ZN(n10487) );
  MUX2_X1 U12464 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n11400), .S(n14000), .Z(
        n10486) );
  NAND2_X1 U12465 ( .A1(n10487), .A2(n10486), .ZN(n14005) );
  NAND2_X1 U12466 ( .A1(n14000), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10488) );
  NAND2_X1 U12467 ( .A1(n14005), .A2(n10488), .ZN(n10529) );
  MUX2_X1 U12468 ( .A(n11595), .B(P2_REG2_REG_9__SCAN_IN), .S(n10530), .Z(
        n10489) );
  OR2_X1 U12469 ( .A1(n10529), .A2(n10489), .ZN(n10531) );
  OR2_X1 U12470 ( .A1(n10530), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n10490) );
  NAND2_X1 U12471 ( .A1(n10531), .A2(n10490), .ZN(n10493) );
  MUX2_X1 U12472 ( .A(n11775), .B(P2_REG2_REG_10__SCAN_IN), .S(n11137), .Z(
        n10492) );
  OR2_X1 U12473 ( .A1(n10493), .A2(n10492), .ZN(n11129) );
  INV_X1 U12474 ( .A(n11129), .ZN(n10491) );
  AOI211_X1 U12475 ( .C1(n10493), .C2(n10492), .A(n15502), .B(n10491), .ZN(
        n10494) );
  AOI211_X1 U12476 ( .C1(n15521), .C2(n11137), .A(n10495), .B(n10494), .ZN(
        n10524) );
  NAND2_X1 U12477 ( .A1(n10496), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10497) );
  NAND2_X1 U12478 ( .A1(n10498), .A2(n10497), .ZN(n15479) );
  MUX2_X1 U12479 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10499), .S(n15473), .Z(
        n15478) );
  NAND2_X1 U12480 ( .A1(n15479), .A2(n15478), .ZN(n15477) );
  NAND2_X1 U12481 ( .A1(n15473), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n13941) );
  NAND2_X1 U12482 ( .A1(n15477), .A2(n13941), .ZN(n10502) );
  MUX2_X1 U12483 ( .A(n10500), .B(P2_REG1_REG_4__SCAN_IN), .S(n13940), .Z(
        n10501) );
  NAND2_X1 U12484 ( .A1(n10502), .A2(n10501), .ZN(n13957) );
  NAND2_X1 U12485 ( .A1(n13936), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n13956) );
  NAND2_X1 U12486 ( .A1(n13957), .A2(n13956), .ZN(n10505) );
  MUX2_X1 U12487 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n10503), .S(n13954), .Z(
        n10504) );
  NAND2_X1 U12488 ( .A1(n10505), .A2(n10504), .ZN(n13967) );
  NAND2_X1 U12489 ( .A1(n13954), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n13966) );
  NAND2_X1 U12490 ( .A1(n13967), .A2(n13966), .ZN(n10508) );
  MUX2_X1 U12491 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10506), .S(n13969), .Z(
        n10507) );
  NAND2_X1 U12492 ( .A1(n10508), .A2(n10507), .ZN(n13982) );
  NAND2_X1 U12493 ( .A1(n13969), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n13981) );
  NAND2_X1 U12494 ( .A1(n13982), .A2(n13981), .ZN(n10511) );
  MUX2_X1 U12495 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10509), .S(n13984), .Z(
        n10510) );
  NAND2_X1 U12496 ( .A1(n10511), .A2(n10510), .ZN(n13997) );
  NAND2_X1 U12497 ( .A1(n13984), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n13996) );
  NAND2_X1 U12498 ( .A1(n13997), .A2(n13996), .ZN(n10514) );
  MUX2_X1 U12499 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10512), .S(n14000), .Z(
        n10513) );
  NAND2_X1 U12500 ( .A1(n10514), .A2(n10513), .ZN(n13999) );
  NAND2_X1 U12501 ( .A1(n14000), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10515) );
  NAND2_X1 U12502 ( .A1(n13999), .A2(n10515), .ZN(n10528) );
  MUX2_X1 U12503 ( .A(n10516), .B(P2_REG1_REG_9__SCAN_IN), .S(n10530), .Z(
        n10527) );
  OR2_X1 U12504 ( .A1(n10528), .A2(n10527), .ZN(n10525) );
  OR2_X1 U12505 ( .A1(n10530), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n10517) );
  NAND2_X1 U12506 ( .A1(n10525), .A2(n10517), .ZN(n10520) );
  INV_X1 U12507 ( .A(n10520), .ZN(n10522) );
  MUX2_X1 U12508 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n10518), .S(n11137), .Z(
        n10521) );
  MUX2_X1 U12509 ( .A(n10518), .B(P2_REG1_REG_10__SCAN_IN), .S(n11137), .Z(
        n10519) );
  OR2_X1 U12510 ( .A1(n10520), .A2(n10519), .ZN(n14018) );
  OAI211_X1 U12511 ( .C1(n10522), .C2(n10521), .A(n15527), .B(n14018), .ZN(
        n10523) );
  NAND2_X1 U12512 ( .A1(n10524), .A2(n10523), .ZN(P2_U3224) );
  INV_X1 U12513 ( .A(n10525), .ZN(n10526) );
  AOI21_X1 U12514 ( .B1(n10528), .B2(n10527), .A(n10526), .ZN(n10539) );
  INV_X1 U12515 ( .A(n10529), .ZN(n10533) );
  MUX2_X1 U12516 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n11595), .S(n10530), .Z(
        n10532) );
  OAI21_X1 U12517 ( .B1(n10533), .B2(n10532), .A(n10531), .ZN(n10537) );
  NAND2_X1 U12518 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n11747) );
  NAND2_X1 U12519 ( .A1(n15501), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n10534) );
  OAI211_X1 U12520 ( .C1(n12095), .C2(n10535), .A(n11747), .B(n10534), .ZN(
        n10536) );
  AOI21_X1 U12521 ( .B1(n10537), .B2(n15523), .A(n10536), .ZN(n10538) );
  OAI21_X1 U12522 ( .B1(n10539), .B2(n15488), .A(n10538), .ZN(P2_U3223) );
  INV_X1 U12523 ( .A(n10540), .ZN(n10541) );
  AOI21_X1 U12524 ( .B1(n10543), .B2(n10542), .A(n10541), .ZN(n10549) );
  OR2_X1 U12525 ( .A1(n10544), .A2(P2_U3088), .ZN(n13875) );
  INV_X1 U12526 ( .A(n13875), .ZN(n10546) );
  OAI22_X1 U12527 ( .A1(n13900), .A2(n10719), .B1(n10546), .B2(n10545), .ZN(
        n10547) );
  AOI21_X1 U12528 ( .B1(n10721), .B2(n13905), .A(n10547), .ZN(n10548) );
  OAI21_X1 U12529 ( .B1(n10549), .B2(n13907), .A(n10548), .ZN(P2_U3194) );
  NOR2_X1 U12530 ( .A1(n10556), .A2(n9750), .ZN(n10552) );
  MUX2_X1 U12531 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10550), .S(n10599), .Z(
        n10551) );
  OAI21_X1 U12532 ( .B1(n10553), .B2(n10552), .A(n10551), .ZN(n10594) );
  INV_X1 U12533 ( .A(n10594), .ZN(n10555) );
  NOR3_X1 U12534 ( .A1(n10553), .A2(n10552), .A3(n10551), .ZN(n10554) );
  NOR3_X1 U12535 ( .A1(n10555), .A2(n10554), .A3(n14811), .ZN(n10567) );
  NAND2_X1 U12536 ( .A1(n10556), .A2(n9745), .ZN(n10557) );
  NAND2_X1 U12537 ( .A1(n10558), .A2(n10557), .ZN(n10562) );
  INV_X1 U12538 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10559) );
  MUX2_X1 U12539 ( .A(n10559), .B(P1_REG1_REG_10__SCAN_IN), .S(n10599), .Z(
        n10561) );
  INV_X1 U12540 ( .A(n10601), .ZN(n10560) );
  AOI211_X1 U12541 ( .C1(n10562), .C2(n10561), .A(n11897), .B(n10560), .ZN(
        n10566) );
  INV_X1 U12542 ( .A(n10599), .ZN(n10564) );
  NAND2_X1 U12543 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n12163)
         );
  NAND2_X1 U12544 ( .A1(n15544), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n10563) );
  OAI211_X1 U12545 ( .C1(n15564), .C2(n10564), .A(n12163), .B(n10563), .ZN(
        n10565) );
  OR3_X1 U12546 ( .A1(n10567), .A2(n10566), .A3(n10565), .ZN(P1_U3253) );
  NOR2_X1 U12547 ( .A1(n10796), .A2(n10795), .ZN(n10580) );
  NAND2_X1 U12548 ( .A1(n10580), .A2(n10568), .ZN(n10582) );
  OR2_X1 U12549 ( .A1(n10582), .A2(n15415), .ZN(n10578) );
  INV_X1 U12550 ( .A(n15982), .ZN(n16006) );
  NAND2_X1 U12551 ( .A1(n16006), .A2(n12868), .ZN(n10569) );
  INV_X1 U12552 ( .A(n12706), .ZN(n11221) );
  AOI22_X1 U12553 ( .A1(n14533), .A2(n11155), .B1(n10570), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n10573) );
  NAND2_X1 U12554 ( .A1(n15878), .A2(n14816), .ZN(n15036) );
  INV_X1 U12555 ( .A(n10632), .ZN(n10571) );
  OR2_X1 U12556 ( .A1(n14588), .A2(n10571), .ZN(n10572) );
  NAND2_X1 U12557 ( .A1(n14533), .A2(n10632), .ZN(n10576) );
  OR2_X1 U12558 ( .A1(n10583), .A2(n10574), .ZN(n10575) );
  OAI211_X1 U12559 ( .C1(n14585), .C2(n10634), .A(n10576), .B(n10575), .ZN(
        n10617) );
  INV_X1 U12560 ( .A(n10617), .ZN(n10577) );
  XNOR2_X1 U12561 ( .A(n10618), .B(n10577), .ZN(n10653) );
  INV_X1 U12562 ( .A(n10653), .ZN(n10591) );
  OR2_X1 U12563 ( .A1(n10578), .A2(n10811), .ZN(n10579) );
  NAND2_X1 U12564 ( .A1(n10580), .A2(n10797), .ZN(n14706) );
  NAND2_X1 U12565 ( .A1(n14704), .A2(n14743), .ZN(n10635) );
  NAND2_X1 U12566 ( .A1(n10582), .A2(n10581), .ZN(n10585) );
  AND2_X1 U12567 ( .A1(n10583), .A2(n12924), .ZN(n10584) );
  NAND2_X1 U12568 ( .A1(n10585), .A2(n10584), .ZN(n10731) );
  INV_X1 U12569 ( .A(n10586), .ZN(n10587) );
  OR2_X1 U12570 ( .A1(n10731), .A2(n10587), .ZN(n10613) );
  NAND2_X1 U12571 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n10613), .ZN(n10588) );
  OAI21_X1 U12572 ( .B1(n14706), .B2(n10635), .A(n10588), .ZN(n10589) );
  AOI21_X1 U12573 ( .B1(n14709), .B2(n11155), .A(n10589), .ZN(n10590) );
  OAI21_X1 U12574 ( .B1(n14711), .B2(n10591), .A(n10590), .ZN(P1_U3232) );
  NAND2_X1 U12575 ( .A1(n10599), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10593) );
  MUX2_X1 U12576 ( .A(n11579), .B(P1_REG2_REG_11__SCAN_IN), .S(n10773), .Z(
        n10592) );
  AOI21_X1 U12577 ( .B1(n10594), .B2(n10593), .A(n10592), .ZN(n10772) );
  NAND3_X1 U12578 ( .A1(n10594), .A2(n10593), .A3(n10592), .ZN(n10595) );
  NAND2_X1 U12579 ( .A1(n10595), .A2(n15558), .ZN(n10607) );
  NOR2_X1 U12580 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10596), .ZN(n12308) );
  INV_X1 U12581 ( .A(n10773), .ZN(n10597) );
  NOR2_X1 U12582 ( .A1(n15564), .A2(n10597), .ZN(n10598) );
  AOI211_X1 U12583 ( .C1(n15544), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n12308), 
        .B(n10598), .ZN(n10606) );
  MUX2_X1 U12584 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9774), .S(n10773), .Z(
        n10603) );
  NAND2_X1 U12585 ( .A1(n10599), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10600) );
  NAND2_X1 U12586 ( .A1(n10602), .A2(n10603), .ZN(n10767) );
  OAI21_X1 U12587 ( .B1(n10603), .B2(n10602), .A(n10767), .ZN(n10604) );
  NAND2_X1 U12588 ( .A1(n10604), .A2(n15566), .ZN(n10605) );
  OAI211_X1 U12589 ( .C1(n10772), .C2(n10607), .A(n10606), .B(n10605), .ZN(
        P1_U3254) );
  INV_X1 U12590 ( .A(n13289), .ZN(n13309) );
  INV_X1 U12591 ( .A(SI_16_), .ZN(n15310) );
  INV_X1 U12592 ( .A(n10608), .ZN(n10609) );
  OAI222_X1 U12593 ( .A1(P3_U3151), .A2(n13309), .B1(n13723), .B2(n15310), 
        .C1(n13730), .C2(n10609), .ZN(P3_U3279) );
  INV_X1 U12594 ( .A(n10610), .ZN(n10630) );
  AOI22_X1 U12595 ( .A1(n10773), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n15423), .ZN(n10611) );
  OAI21_X1 U12596 ( .B1(n10630), .B2(n15437), .A(n10611), .ZN(P1_U3344) );
  OAI222_X1 U12597 ( .A1(n13318), .A2(P3_U3151), .B1(n13730), .B2(n10612), 
        .C1(n13723), .C2(n15301), .ZN(P3_U3278) );
  INV_X1 U12598 ( .A(n10613), .ZN(n10652) );
  NAND2_X1 U12599 ( .A1(n14704), .A2(n14742), .ZN(n10615) );
  NAND2_X1 U12600 ( .A1(n14702), .A2(n10632), .ZN(n10614) );
  NAND2_X1 U12601 ( .A1(n10615), .A2(n10614), .ZN(n11153) );
  AOI22_X1 U12602 ( .A1(n14709), .A2(n15835), .B1(n14671), .B2(n11153), .ZN(
        n10629) );
  NAND2_X1 U12603 ( .A1(n14492), .A2(n15835), .ZN(n10620) );
  NAND2_X1 U12604 ( .A1(n14533), .A2(n14743), .ZN(n10619) );
  NAND2_X1 U12605 ( .A1(n10620), .A2(n10619), .ZN(n10621) );
  XNOR2_X1 U12606 ( .A(n10621), .B(n14522), .ZN(n10623) );
  INV_X1 U12607 ( .A(n14743), .ZN(n12710) );
  NAND2_X1 U12608 ( .A1(n14533), .A2(n15835), .ZN(n10622) );
  NAND2_X1 U12609 ( .A1(n10623), .A2(n10624), .ZN(n10644) );
  NAND2_X1 U12610 ( .A1(n10627), .A2(n14690), .ZN(n10628) );
  OAI211_X1 U12611 ( .C1(n10652), .C2(n11158), .A(n10629), .B(n10628), .ZN(
        P1_U3222) );
  OAI222_X1 U12612 ( .A1(n14422), .A2(n10631), .B1(n14416), .B2(n10630), .C1(
        P2_U3088), .C2(n14015), .ZN(P2_U3316) );
  NAND2_X1 U12613 ( .A1(n10632), .A2(n10634), .ZN(n12708) );
  AND2_X1 U12614 ( .A1(n12707), .A2(n12708), .ZN(n12875) );
  INV_X1 U12615 ( .A(n12875), .ZN(n15831) );
  NOR3_X1 U12616 ( .A1(n15443), .A2(n10634), .A3(n10633), .ZN(n15830) );
  INV_X1 U12617 ( .A(n15874), .ZN(n15837) );
  OAI21_X1 U12618 ( .B1(n15837), .B2(n16013), .A(n15831), .ZN(n10636) );
  NAND2_X1 U12619 ( .A1(n10636), .A2(n10635), .ZN(n15828) );
  AOI211_X1 U12620 ( .C1(n15926), .C2(n15831), .A(n15830), .B(n15828), .ZN(
        n15826) );
  NAND2_X1 U12621 ( .A1(n7362), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10637) );
  OAI21_X1 U12622 ( .B1(n15826), .B2(n7362), .A(n10637), .ZN(P1_U3528) );
  AND2_X1 U12623 ( .A1(n10638), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U12624 ( .A1(n10638), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U12625 ( .A1(n10638), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U12626 ( .A1(n10638), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U12627 ( .A1(n10638), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U12628 ( .A1(n10638), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U12629 ( .A1(n10638), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U12630 ( .A1(n10638), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U12631 ( .A1(n10638), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U12632 ( .A1(n10638), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U12633 ( .A1(n10638), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U12634 ( .A1(n10638), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U12635 ( .A1(n10638), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  NAND2_X1 U12636 ( .A1(n13872), .A2(n14275), .ZN(n13859) );
  INV_X1 U12637 ( .A(n13859), .ZN(n13887) );
  NAND2_X1 U12638 ( .A1(n13887), .A2(n13932), .ZN(n10641) );
  MUX2_X1 U12639 ( .A(n11243), .B(n11250), .S(n14151), .Z(n10639) );
  AOI22_X1 U12640 ( .A1(n13881), .A2(n10639), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n13875), .ZN(n10640) );
  OAI211_X1 U12641 ( .C1(n13889), .C2(n10642), .A(n10641), .B(n10640), .ZN(
        P2_U3204) );
  OAI22_X1 U12642 ( .A1(n15880), .A2(n14585), .B1(n14590), .B2(n7903), .ZN(
        n10643) );
  XNOR2_X1 U12643 ( .A(n10643), .B(n14522), .ZN(n10724) );
  OAI22_X1 U12644 ( .A1(n14588), .A2(n7903), .B1(n15880), .B2(n14590), .ZN(
        n10725) );
  XNOR2_X1 U12645 ( .A(n10724), .B(n10725), .ZN(n10647) );
  NAND2_X1 U12646 ( .A1(n10645), .A2(n10644), .ZN(n10646) );
  OAI21_X1 U12647 ( .B1(n10647), .B2(n10646), .A(n10728), .ZN(n10648) );
  NAND2_X1 U12648 ( .A1(n10648), .A2(n14690), .ZN(n10650) );
  INV_X1 U12649 ( .A(n14702), .ZN(n14605) );
  OAI22_X1 U12650 ( .A1(n12721), .A2(n14607), .B1(n14605), .B2(n12710), .ZN(
        n15876) );
  AOI22_X1 U12651 ( .A1(n14709), .A2(n15888), .B1(n14671), .B2(n15876), .ZN(
        n10649) );
  OAI211_X1 U12652 ( .C1(n10652), .C2(n10651), .A(n10650), .B(n10649), .ZN(
        P1_U3237) );
  INV_X1 U12653 ( .A(P1_U4016), .ZN(n14727) );
  NAND2_X1 U12654 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14744) );
  MUX2_X1 U12655 ( .A(n10653), .B(n14744), .S(n12925), .Z(n10654) );
  NOR2_X1 U12656 ( .A1(n10654), .A2(n15429), .ZN(n10655) );
  AOI211_X1 U12657 ( .C1(n10657), .C2(n10656), .A(n14727), .B(n10655), .ZN(
        n10685) );
  MUX2_X1 U12658 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10347), .S(n10668), .Z(
        n10659) );
  NAND3_X1 U12659 ( .A1(n10659), .A2(n14765), .A3(n10658), .ZN(n10660) );
  AND3_X1 U12660 ( .A1(n15566), .A2(n10661), .A3(n10660), .ZN(n10671) );
  INV_X1 U12661 ( .A(n10662), .ZN(n10666) );
  NOR3_X1 U12662 ( .A1(n14766), .A2(n10664), .A3(n10663), .ZN(n10665) );
  NOR3_X1 U12663 ( .A1(n14811), .A2(n10666), .A3(n10665), .ZN(n10670) );
  NAND2_X1 U12664 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10956) );
  NAND2_X1 U12665 ( .A1(n15544), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n10667) );
  OAI211_X1 U12666 ( .C1(n15564), .C2(n10668), .A(n10956), .B(n10667), .ZN(
        n10669) );
  OR4_X1 U12667 ( .A1(n10685), .A2(n10671), .A3(n10670), .A4(n10669), .ZN(
        P1_U3247) );
  INV_X1 U12668 ( .A(n14769), .ZN(n10672) );
  AOI211_X1 U12669 ( .C1(n10674), .C2(n10673), .A(n10672), .B(n14811), .ZN(
        n10684) );
  INV_X1 U12670 ( .A(n10675), .ZN(n10678) );
  MUX2_X1 U12671 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10342), .S(n10681), .Z(
        n10677) );
  INV_X1 U12672 ( .A(n14763), .ZN(n10676) );
  AOI211_X1 U12673 ( .C1(n10678), .C2(n10677), .A(n10676), .B(n11897), .ZN(
        n10683) );
  NAND2_X1 U12674 ( .A1(P1_U3086), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n10680) );
  NAND2_X1 U12675 ( .A1(n15544), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n10679) );
  OAI211_X1 U12676 ( .C1(n15564), .C2(n10681), .A(n10680), .B(n10679), .ZN(
        n10682) );
  OR4_X1 U12677 ( .A1(n10685), .A2(n10684), .A3(n10683), .A4(n10682), .ZN(
        P1_U3245) );
  INV_X1 U12678 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10696) );
  XNOR2_X1 U12679 ( .A(n12729), .B(n10928), .ZN(n12878) );
  XNOR2_X1 U12680 ( .A(n10686), .B(n12878), .ZN(n11127) );
  XNOR2_X1 U12681 ( .A(n10687), .B(n12878), .ZN(n11125) );
  NAND2_X1 U12682 ( .A1(n14704), .A2(n14739), .ZN(n10689) );
  NAND2_X1 U12683 ( .A1(n14702), .A2(n14741), .ZN(n10688) );
  AND2_X1 U12684 ( .A1(n10689), .A2(n10688), .ZN(n11115) );
  INV_X1 U12685 ( .A(n11115), .ZN(n10692) );
  NAND2_X1 U12686 ( .A1(n12729), .A2(n11230), .ZN(n10690) );
  NAND2_X1 U12687 ( .A1(n10690), .A2(n15878), .ZN(n10691) );
  NOR2_X1 U12688 ( .A1(n11076), .A2(n10691), .ZN(n11122) );
  AOI211_X1 U12689 ( .C1(n11125), .C2(n15992), .A(n10692), .B(n11122), .ZN(
        n10693) );
  OAI21_X1 U12690 ( .B1(n15987), .B2(n11127), .A(n10693), .ZN(n10697) );
  NAND2_X1 U12691 ( .A1(n10697), .A2(n16017), .ZN(n10695) );
  NAND2_X1 U12692 ( .A1(n10105), .A2(n12729), .ZN(n10694) );
  OAI211_X1 U12693 ( .C1(n16017), .C2(n10696), .A(n10695), .B(n10694), .ZN(
        P1_U3471) );
  NAND2_X1 U12694 ( .A1(n10697), .A2(n16014), .ZN(n10699) );
  NAND2_X1 U12695 ( .A1(n10229), .A2(n12729), .ZN(n10698) );
  OAI211_X1 U12696 ( .C1(n16014), .C2(n10347), .A(n10699), .B(n10698), .ZN(
        P1_U3532) );
  INV_X1 U12697 ( .A(n13350), .ZN(n13334) );
  INV_X1 U12698 ( .A(n10700), .ZN(n10701) );
  OAI222_X1 U12699 ( .A1(P3_U3151), .A2(n13334), .B1(n13723), .B2(n15300), 
        .C1(n13730), .C2(n10701), .ZN(P3_U3277) );
  OAI21_X1 U12700 ( .B1(n10704), .B2(n10703), .A(n10702), .ZN(n11377) );
  INV_X1 U12701 ( .A(n10716), .ZN(n10705) );
  AOI211_X1 U12702 ( .C1(n13876), .C2(n10705), .A(n14282), .B(n10744), .ZN(
        n11372) );
  XNOR2_X1 U12703 ( .A(n10707), .B(n10706), .ZN(n10708) );
  NAND2_X1 U12704 ( .A1(n10708), .A2(n14271), .ZN(n10710) );
  AOI22_X1 U12705 ( .A1(n13929), .A2(n14275), .B1(n14274), .B2(n13932), .ZN(
        n10709) );
  NAND2_X1 U12706 ( .A1(n10710), .A2(n10709), .ZN(n11371) );
  AOI211_X1 U12707 ( .C1(n16033), .C2(n11377), .A(n11372), .B(n11371), .ZN(
        n11285) );
  AOI22_X1 U12708 ( .A1(n14300), .A2(n13876), .B1(n16034), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n10711) );
  OAI21_X1 U12709 ( .B1(n11285), .B2(n16034), .A(n10711), .ZN(P2_U3501) );
  OAI21_X1 U12710 ( .B1(n10717), .B2(n10713), .A(n10712), .ZN(n11506) );
  NAND2_X1 U12711 ( .A1(n10721), .A2(n11250), .ZN(n10714) );
  NAND2_X1 U12712 ( .A1(n10714), .A2(n14151), .ZN(n10715) );
  NOR2_X1 U12713 ( .A1(n10716), .A2(n10715), .ZN(n11501) );
  XOR2_X1 U12714 ( .A(n10718), .B(n10717), .Z(n10720) );
  OAI21_X1 U12715 ( .B1(n10720), .B2(n14243), .A(n10719), .ZN(n11500) );
  AOI211_X1 U12716 ( .C1(n16033), .C2(n11506), .A(n11501), .B(n11500), .ZN(
        n11289) );
  AOI22_X1 U12717 ( .A1(n14300), .A2(n10721), .B1(n16034), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n10722) );
  OAI21_X1 U12718 ( .B1(n11289), .B2(n16034), .A(n10722), .ZN(P2_U3500) );
  INV_X2 U12719 ( .A(n14533), .ZN(n14590) );
  OAI22_X1 U12720 ( .A1(n15898), .A2(n14585), .B1(n12721), .B2(n14590), .ZN(
        n10723) );
  XNOR2_X1 U12721 ( .A(n10723), .B(n14522), .ZN(n10903) );
  OAI22_X1 U12722 ( .A1(n15898), .A2(n14590), .B1(n12721), .B2(n14588), .ZN(
        n10904) );
  XNOR2_X1 U12723 ( .A(n10903), .B(n10904), .ZN(n10730) );
  INV_X1 U12724 ( .A(n10724), .ZN(n10726) );
  OR2_X1 U12725 ( .A1(n10726), .A2(n10725), .ZN(n10727) );
  OAI211_X1 U12726 ( .C1(n10730), .C2(n10729), .A(n10912), .B(n14690), .ZN(
        n10738) );
  INV_X1 U12727 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n14758) );
  NAND2_X1 U12728 ( .A1(n10731), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10732) );
  INV_X1 U12729 ( .A(n14701), .ZN(n14695) );
  INV_X1 U12730 ( .A(n14709), .ZN(n14698) );
  NAND2_X1 U12731 ( .A1(n14704), .A2(n14740), .ZN(n10734) );
  NAND2_X1 U12732 ( .A1(n14702), .A2(n14742), .ZN(n10733) );
  NAND2_X1 U12733 ( .A1(n10734), .A2(n10733), .ZN(n11225) );
  AOI22_X1 U12734 ( .A1(n14671), .A2(n11225), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10735) );
  OAI21_X1 U12735 ( .B1(n14698), .B2(n15898), .A(n10735), .ZN(n10736) );
  AOI21_X1 U12736 ( .B1(n14758), .B2(n14695), .A(n10736), .ZN(n10737) );
  NAND2_X1 U12737 ( .A1(n10738), .A2(n10737), .ZN(P1_U3218) );
  INV_X1 U12738 ( .A(n10739), .ZN(n10740) );
  INV_X1 U12739 ( .A(n11001), .ZN(n10768) );
  OAI222_X1 U12740 ( .A1(n15435), .A2(n7678), .B1(n15437), .B2(n10740), .C1(
        n10768), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U12741 ( .A(n15522), .ZN(n11143) );
  OAI222_X1 U12742 ( .A1(n14422), .A2(n10741), .B1(n12358), .B2(n10740), .C1(
        n11143), .C2(P2_U3088), .ZN(P2_U3315) );
  OAI21_X1 U12743 ( .B1(n10743), .B2(n10746), .A(n10742), .ZN(n11419) );
  INV_X1 U12744 ( .A(n10744), .ZN(n10745) );
  AOI211_X1 U12745 ( .C1(n10750), .C2(n10745), .A(n14282), .B(n10753), .ZN(
        n11418) );
  XNOR2_X1 U12746 ( .A(n10747), .B(n10746), .ZN(n10749) );
  OAI21_X1 U12747 ( .B1(n10749), .B2(n14243), .A(n10748), .ZN(n11414) );
  AOI211_X1 U12748 ( .C1(n16033), .C2(n11419), .A(n11418), .B(n11414), .ZN(
        n11281) );
  AOI22_X1 U12749 ( .A1(n14300), .A2(n10750), .B1(n16034), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n10751) );
  OAI21_X1 U12750 ( .B1(n11281), .B2(n16034), .A(n10751), .ZN(P2_U3502) );
  XNOR2_X1 U12751 ( .A(n10752), .B(n10756), .ZN(n11529) );
  INV_X1 U12752 ( .A(n10753), .ZN(n10754) );
  AOI211_X1 U12753 ( .C1(n10755), .C2(n10754), .A(n8098), .B(n10963), .ZN(
        n11526) );
  AOI21_X1 U12754 ( .B1(n14347), .B2(n10755), .A(n11526), .ZN(n10760) );
  XNOR2_X1 U12755 ( .A(n10757), .B(n10756), .ZN(n10759) );
  OAI22_X1 U12756 ( .A1(n10758), .A2(n14235), .B1(n11067), .B2(n14237), .ZN(
        n10790) );
  AOI21_X1 U12757 ( .B1(n10759), .B2(n14271), .A(n10790), .ZN(n11521) );
  OAI211_X1 U12758 ( .C1(n14353), .C2(n11529), .A(n10760), .B(n11521), .ZN(
        n10845) );
  NAND2_X1 U12759 ( .A1(n10845), .A2(n16035), .ZN(n10761) );
  OAI21_X1 U12760 ( .B1(n16035), .B2(n10500), .A(n10761), .ZN(P2_U3503) );
  INV_X1 U12761 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10763) );
  INV_X1 U12762 ( .A(n15507), .ZN(n10762) );
  OAI222_X1 U12763 ( .A1(n14422), .A2(n10763), .B1(n12358), .B2(n10764), .C1(
        n10762), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U12764 ( .A(n11630), .ZN(n11010) );
  OAI222_X1 U12765 ( .A1(P1_U3086), .A2(n11010), .B1(n15435), .B2(n10765), 
        .C1(n10764), .C2(n15437), .ZN(P1_U3342) );
  OR2_X1 U12766 ( .A1(n10773), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10766) );
  NAND2_X1 U12767 ( .A1(n10767), .A2(n10766), .ZN(n10769) );
  NAND2_X1 U12768 ( .A1(n10769), .A2(n10768), .ZN(n11005) );
  OAI21_X1 U12769 ( .B1(n10769), .B2(n10768), .A(n11005), .ZN(n10771) );
  OR2_X1 U12770 ( .A1(n10771), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11006) );
  INV_X1 U12771 ( .A(n11006), .ZN(n10770) );
  AOI21_X1 U12772 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n10771), .A(n10770), 
        .ZN(n10781) );
  MUX2_X1 U12773 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n9786), .S(n11001), .Z(
        n10775) );
  AOI21_X1 U12774 ( .B1(n10773), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10772), 
        .ZN(n10774) );
  NAND2_X1 U12775 ( .A1(n10774), .A2(n10775), .ZN(n11000) );
  OAI21_X1 U12776 ( .B1(n10775), .B2(n10774), .A(n11000), .ZN(n10779) );
  INV_X1 U12777 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10777) );
  NAND2_X1 U12778 ( .A1(n15548), .A2(n11001), .ZN(n10776) );
  NAND2_X1 U12779 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n12327)
         );
  OAI211_X1 U12780 ( .C1(n10777), .C2(n15570), .A(n10776), .B(n12327), .ZN(
        n10778) );
  AOI21_X1 U12781 ( .B1(n10779), .B2(n15558), .A(n10778), .ZN(n10780) );
  OAI21_X1 U12782 ( .B1(n10781), .B2(n11897), .A(n10780), .ZN(P1_U3255) );
  XNOR2_X1 U12783 ( .A(n11524), .B(n13764), .ZN(n10821) );
  NOR2_X1 U12784 ( .A1(n10785), .A2(n14348), .ZN(n10819) );
  XNOR2_X1 U12785 ( .A(n10821), .B(n10819), .ZN(n10786) );
  OAI21_X1 U12786 ( .B1(n10787), .B2(n10786), .A(n7335), .ZN(n10788) );
  NAND2_X1 U12787 ( .A1(n10788), .A2(n13881), .ZN(n10792) );
  NAND2_X1 U12788 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n13933) );
  OAI21_X1 U12789 ( .B1(n13902), .B2(n11523), .A(n13933), .ZN(n10789) );
  AOI21_X1 U12790 ( .B1(n13872), .B2(n10790), .A(n10789), .ZN(n10791) );
  OAI211_X1 U12791 ( .C1(n11524), .C2(n13889), .A(n10792), .B(n10791), .ZN(
        P2_U3202) );
  INV_X1 U12792 ( .A(n10793), .ZN(n10794) );
  OAI222_X1 U12793 ( .A1(n13723), .A2(n15303), .B1(P3_U3151), .B2(n13361), 
        .C1(n13730), .C2(n10794), .ZN(P3_U3276) );
  INV_X1 U12794 ( .A(n10795), .ZN(n10798) );
  NAND3_X1 U12795 ( .A1(n10798), .A2(n10797), .A3(n10796), .ZN(n14837) );
  INV_X1 U12796 ( .A(n10799), .ZN(n11558) );
  OAI21_X1 U12797 ( .B1(n10801), .B2(n10802), .A(n10800), .ZN(n10840) );
  INV_X1 U12798 ( .A(n10840), .ZN(n10816) );
  XNOR2_X1 U12799 ( .A(n10803), .B(n10802), .ZN(n10807) );
  NAND2_X1 U12800 ( .A1(n14704), .A2(n14737), .ZN(n10805) );
  NAND2_X1 U12801 ( .A1(n14702), .A2(n14739), .ZN(n10804) );
  NAND2_X1 U12802 ( .A1(n10805), .A2(n10804), .ZN(n11304) );
  INV_X1 U12803 ( .A(n11304), .ZN(n10806) );
  OAI21_X1 U12804 ( .B1(n10807), .B2(n15987), .A(n10806), .ZN(n10838) );
  INV_X1 U12805 ( .A(n10838), .ZN(n10808) );
  MUX2_X1 U12806 ( .A(n10809), .B(n10808), .S(n15054), .Z(n10815) );
  AOI211_X1 U12807 ( .C1(n12741), .C2(n11077), .A(n15985), .B(n10810), .ZN(
        n10839) );
  INV_X1 U12808 ( .A(n12741), .ZN(n12742) );
  INV_X1 U12809 ( .A(n10811), .ZN(n10812) );
  OAI22_X1 U12810 ( .A1(n12742), .A2(n15942), .B1(n11302), .B2(n15051), .ZN(
        n10813) );
  AOI21_X1 U12811 ( .B1(n10839), .B2(n15935), .A(n10813), .ZN(n10814) );
  OAI211_X1 U12812 ( .C1(n15061), .C2(n10816), .A(n10815), .B(n10814), .ZN(
        P1_U3287) );
  INV_X1 U12813 ( .A(n10817), .ZN(n10950) );
  AOI22_X1 U12814 ( .A1(n11888), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n15423), .ZN(n10818) );
  OAI21_X1 U12815 ( .B1(n10950), .B2(n15437), .A(n10818), .ZN(P1_U3341) );
  XNOR2_X1 U12816 ( .A(n11535), .B(n13805), .ZN(n11057) );
  NOR2_X1 U12817 ( .A1(n11067), .A2(n14348), .ZN(n11055) );
  XNOR2_X1 U12818 ( .A(n11057), .B(n11055), .ZN(n10825) );
  INV_X1 U12819 ( .A(n10819), .ZN(n10820) );
  NAND2_X1 U12820 ( .A1(n10821), .A2(n10820), .ZN(n10822) );
  OAI21_X1 U12821 ( .B1(n10825), .B2(n10824), .A(n11059), .ZN(n10826) );
  NAND2_X1 U12822 ( .A1(n10826), .A2(n13881), .ZN(n10830) );
  AOI22_X1 U12823 ( .A1(n13928), .A2(n14274), .B1(n14275), .B2(n13926), .ZN(
        n10967) );
  INV_X1 U12824 ( .A(n10967), .ZN(n10828) );
  NAND2_X1 U12825 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n13947) );
  OAI21_X1 U12826 ( .B1(n13902), .B2(n11534), .A(n13947), .ZN(n10827) );
  AOI21_X1 U12827 ( .B1(n13872), .B2(n10828), .A(n10827), .ZN(n10829) );
  OAI211_X1 U12828 ( .C1(n11535), .C2(n13889), .A(n10830), .B(n10829), .ZN(
        P2_U3199) );
  INV_X1 U12829 ( .A(n11314), .ZN(n11413) );
  NOR2_X1 U12830 ( .A1(n11016), .A2(n11314), .ZN(n12535) );
  INV_X1 U12831 ( .A(n11313), .ZN(n11014) );
  NOR2_X1 U12832 ( .A1(n12535), .A2(n11014), .ZN(n12660) );
  NAND2_X1 U12833 ( .A1(n11095), .A2(n15970), .ZN(n10831) );
  OAI22_X1 U12834 ( .A1(n12660), .A2(n10831), .B1(n11316), .B2(n13580), .ZN(
        n11409) );
  NOR2_X1 U12835 ( .A1(n16039), .A2(n10883), .ZN(n10832) );
  AOI21_X1 U12836 ( .B1(n11409), .B2(n16039), .A(n10832), .ZN(n10833) );
  OAI21_X1 U12837 ( .B1(n11413), .B2(n13656), .A(n10833), .ZN(P3_U3459) );
  INV_X1 U12838 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10837) );
  AOI22_X1 U12839 ( .A1(n11243), .A2(n14271), .B1(n14275), .B2(n13932), .ZN(
        n11245) );
  AOI22_X1 U12840 ( .A1(n11243), .A2(n16033), .B1(n10834), .B2(n11250), .ZN(
        n10835) );
  NAND2_X1 U12841 ( .A1(n11245), .A2(n10835), .ZN(n14370) );
  NAND2_X1 U12842 ( .A1(n14371), .A2(n14370), .ZN(n10836) );
  OAI21_X1 U12843 ( .B1(n14398), .B2(n10837), .A(n10836), .ZN(P2_U3430) );
  AOI211_X1 U12844 ( .C1(n15992), .C2(n10840), .A(n10839), .B(n10838), .ZN(
        n10844) );
  OAI22_X1 U12845 ( .A1(n12742), .A2(n15402), .B1(n16017), .B2(n9703), .ZN(
        n10841) );
  INV_X1 U12846 ( .A(n10841), .ZN(n10842) );
  OAI21_X1 U12847 ( .B1(n10844), .B2(n7917), .A(n10842), .ZN(P1_U3477) );
  AOI22_X1 U12848 ( .A1(n10229), .A2(n12741), .B1(n7362), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n10843) );
  OAI21_X1 U12849 ( .B1(n10844), .B2(n7362), .A(n10843), .ZN(P1_U3534) );
  INV_X1 U12850 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10847) );
  NAND2_X1 U12851 ( .A1(n10845), .A2(n14371), .ZN(n10846) );
  OAI21_X1 U12852 ( .B1(n14398), .B2(n10847), .A(n10846), .ZN(P2_U3442) );
  INV_X1 U12853 ( .A(n11109), .ZN(n10848) );
  OR2_X1 U12854 ( .A1(n10849), .A2(P3_U3151), .ZN(n12700) );
  NAND2_X1 U12855 ( .A1(n10848), .A2(n12700), .ZN(n10872) );
  INV_X1 U12856 ( .A(n10849), .ZN(n10851) );
  OAI21_X1 U12857 ( .B1(n12635), .B2(n10851), .A(n10850), .ZN(n10871) );
  INV_X1 U12858 ( .A(n10871), .ZN(n10852) );
  NAND2_X1 U12859 ( .A1(n10872), .A2(n10852), .ZN(n10869) );
  MUX2_X1 U12860 ( .A(n10869), .B(n13240), .S(n10853), .Z(n13362) );
  MUX2_X1 U12861 ( .A(n8201), .B(P3_REG1_REG_2__SCAN_IN), .S(n10885), .Z(
        n11024) );
  AND2_X1 U12862 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n10862), .ZN(n10854) );
  OAI21_X1 U12863 ( .B1(n11274), .B2(n10854), .A(n10855), .ZN(n11265) );
  OR2_X1 U12864 ( .A1(n11265), .A2(n10877), .ZN(n11267) );
  NAND2_X1 U12865 ( .A1(n11267), .A2(n10855), .ZN(n11023) );
  NAND2_X1 U12866 ( .A1(n11038), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10856) );
  NAND2_X1 U12867 ( .A1(n10934), .A2(n10859), .ZN(n10857) );
  INV_X1 U12868 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15910) );
  MUX2_X1 U12869 ( .A(n15910), .B(P3_REG1_REG_4__SCAN_IN), .S(n10985), .Z(
        n10858) );
  NAND2_X1 U12870 ( .A1(n10857), .A2(n10858), .ZN(n10987) );
  INV_X1 U12871 ( .A(n10858), .ZN(n10860) );
  NAND3_X1 U12872 ( .A1(n10934), .A2(n10860), .A3(n10859), .ZN(n10861) );
  AOI21_X1 U12873 ( .B1(n10987), .B2(n10861), .A(n15800), .ZN(n10876) );
  INV_X1 U12874 ( .A(n11274), .ZN(n10879) );
  NAND2_X1 U12875 ( .A1(n10862), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10863) );
  MUX2_X1 U12876 ( .A(n10884), .B(P3_REG2_REG_2__SCAN_IN), .S(n10885), .Z(
        n11027) );
  OAI21_X1 U12877 ( .B1(n10885), .B2(n10884), .A(n11025), .ZN(n10865) );
  XNOR2_X1 U12878 ( .A(n10865), .B(n10891), .ZN(n10935) );
  MUX2_X1 U12879 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n11670), .S(n10985), .Z(
        n10866) );
  NAND2_X1 U12880 ( .A1(n10867), .A2(n10866), .ZN(n10870) );
  AOI21_X1 U12881 ( .B1(n10971), .B2(n10870), .A(n15742), .ZN(n10875) );
  INV_X1 U12882 ( .A(n15806), .ZN(n15787) );
  INV_X1 U12883 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n10873) );
  NOR2_X1 U12884 ( .A1(n15787), .A2(n10873), .ZN(n10874) );
  NOR2_X1 U12885 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15356), .ZN(n13157) );
  NOR4_X1 U12886 ( .A1(n10876), .A2(n10875), .A3(n10874), .A4(n13157), .ZN(
        n10901) );
  INV_X1 U12887 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10878) );
  INV_X1 U12888 ( .A(n12695), .ZN(n11797) );
  MUX2_X1 U12889 ( .A(n10878), .B(n10877), .S(n8664), .Z(n10880) );
  NAND2_X1 U12890 ( .A1(n10880), .A2(n10879), .ZN(n11031) );
  INV_X1 U12891 ( .A(n10880), .ZN(n10881) );
  NAND2_X1 U12892 ( .A1(n10881), .A2(n11274), .ZN(n10882) );
  NAND2_X1 U12893 ( .A1(n11031), .A2(n10882), .ZN(n11263) );
  MUX2_X1 U12894 ( .A(n11411), .B(n10883), .S(n11797), .Z(n15744) );
  NAND2_X1 U12895 ( .A1(n15744), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15743) );
  NAND2_X1 U12896 ( .A1(n11030), .A2(n11031), .ZN(n10889) );
  MUX2_X1 U12897 ( .A(n10884), .B(n8201), .S(n11797), .Z(n10886) );
  NAND2_X1 U12898 ( .A1(n10886), .A2(n10885), .ZN(n10941) );
  INV_X1 U12899 ( .A(n10886), .ZN(n10887) );
  NAND2_X1 U12900 ( .A1(n10887), .A2(n11038), .ZN(n10888) );
  AND2_X1 U12901 ( .A1(n10941), .A2(n10888), .ZN(n11032) );
  NAND2_X1 U12902 ( .A1(n10889), .A2(n11032), .ZN(n10940) );
  NAND2_X1 U12903 ( .A1(n10940), .A2(n10941), .ZN(n10895) );
  INV_X1 U12904 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11845) );
  MUX2_X1 U12905 ( .A(n11845), .B(n10890), .S(n13728), .Z(n10892) );
  NAND2_X1 U12906 ( .A1(n10892), .A2(n10891), .ZN(n10896) );
  INV_X1 U12907 ( .A(n10892), .ZN(n10893) );
  NAND2_X1 U12908 ( .A1(n10893), .A2(n10949), .ZN(n10894) );
  AND2_X1 U12909 ( .A1(n10896), .A2(n10894), .ZN(n10942) );
  MUX2_X1 U12910 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n13728), .Z(n10973) );
  XNOR2_X1 U12911 ( .A(n10973), .B(n10985), .ZN(n10897) );
  NAND2_X1 U12912 ( .A1(n10898), .A2(n10897), .ZN(n10976) );
  OAI21_X1 U12913 ( .B1(n10898), .B2(n10897), .A(n10976), .ZN(n10899) );
  AND2_X1 U12914 ( .A1(P3_U3897), .A2(n8663), .ZN(n15814) );
  NAND2_X1 U12915 ( .A1(n10899), .A2(n15814), .ZN(n10900) );
  OAI211_X1 U12916 ( .C1(n13362), .C2(n10902), .A(n10901), .B(n10900), .ZN(
        P3_U3186) );
  INV_X1 U12917 ( .A(n10903), .ZN(n10905) );
  NAND2_X1 U12918 ( .A1(n10905), .A2(n10904), .ZN(n10911) );
  NOR2_X1 U12919 ( .A1(n14588), .A2(n10928), .ZN(n10906) );
  AOI21_X1 U12920 ( .B1(n12729), .B2(n14442), .A(n10906), .ZN(n10913) );
  AND2_X1 U12921 ( .A1(n10911), .A2(n10913), .ZN(n10907) );
  NAND2_X1 U12922 ( .A1(n10912), .A2(n10907), .ZN(n10952) );
  NAND2_X1 U12923 ( .A1(n12729), .A2(n14532), .ZN(n10909) );
  NAND2_X1 U12924 ( .A1(n14442), .A2(n14740), .ZN(n10908) );
  NAND2_X1 U12925 ( .A1(n10909), .A2(n10908), .ZN(n10910) );
  XNOR2_X1 U12926 ( .A(n10910), .B(n14586), .ZN(n10955) );
  NAND2_X1 U12927 ( .A1(n10952), .A2(n10955), .ZN(n10916) );
  INV_X1 U12928 ( .A(n10913), .ZN(n10914) );
  NAND2_X1 U12929 ( .A1(n10915), .A2(n10914), .ZN(n10953) );
  NAND2_X1 U12930 ( .A1(n12738), .A2(n14532), .ZN(n10918) );
  NAND2_X1 U12931 ( .A1(n14509), .A2(n14739), .ZN(n10917) );
  NAND2_X1 U12932 ( .A1(n10918), .A2(n10917), .ZN(n10919) );
  XNOR2_X1 U12933 ( .A(n10919), .B(n14586), .ZN(n10925) );
  INV_X1 U12934 ( .A(n10925), .ZN(n10923) );
  NAND2_X1 U12935 ( .A1(n12738), .A2(n14509), .ZN(n10921) );
  NAND2_X1 U12936 ( .A1(n14537), .A2(n14739), .ZN(n10920) );
  NAND2_X1 U12937 ( .A1(n10921), .A2(n10920), .ZN(n10924) );
  INV_X1 U12938 ( .A(n10924), .ZN(n10922) );
  NAND2_X1 U12939 ( .A1(n10923), .A2(n10922), .ZN(n11296) );
  INV_X1 U12940 ( .A(n11296), .ZN(n10926) );
  AND2_X1 U12941 ( .A1(n10925), .A2(n10924), .ZN(n11294) );
  NOR2_X1 U12942 ( .A1(n10926), .A2(n11294), .ZN(n10927) );
  XNOR2_X1 U12943 ( .A(n11295), .B(n10927), .ZN(n10933) );
  OAI22_X1 U12944 ( .A1(n12743), .A2(n14607), .B1(n14605), .B2(n10928), .ZN(
        n11083) );
  NAND2_X1 U12945 ( .A1(n14671), .A2(n11083), .ZN(n10929) );
  OAI211_X1 U12946 ( .C1(n14701), .C2(n15912), .A(n10930), .B(n10929), .ZN(
        n10931) );
  AOI21_X1 U12947 ( .B1(n12738), .B2(n14709), .A(n10931), .ZN(n10932) );
  OAI21_X1 U12948 ( .B1(n10933), .B2(n14711), .A(n10932), .ZN(P1_U3227) );
  OAI21_X1 U12949 ( .B1(n7295), .B2(P3_REG1_REG_3__SCAN_IN), .A(n10934), .ZN(
        n10939) );
  XNOR2_X1 U12950 ( .A(n10935), .B(n11845), .ZN(n10937) );
  NOR2_X1 U12951 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15169), .ZN(n11427) );
  AOI21_X1 U12952 ( .B1(n15806), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n11427), .ZN(
        n10936) );
  OAI21_X1 U12953 ( .B1(n10937), .B2(n15742), .A(n10936), .ZN(n10938) );
  AOI21_X1 U12954 ( .B1(n15819), .B2(n10939), .A(n10938), .ZN(n10948) );
  INV_X1 U12955 ( .A(n10940), .ZN(n11034) );
  INV_X1 U12956 ( .A(n10941), .ZN(n10943) );
  NOR3_X1 U12957 ( .A1(n11034), .A2(n10943), .A3(n10942), .ZN(n10946) );
  INV_X1 U12958 ( .A(n10944), .ZN(n10945) );
  OAI21_X1 U12959 ( .B1(n10946), .B2(n10945), .A(n15814), .ZN(n10947) );
  OAI211_X1 U12960 ( .C1(n13362), .C2(n10949), .A(n10948), .B(n10947), .ZN(
        P3_U3185) );
  INV_X1 U12961 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10951) );
  INV_X1 U12962 ( .A(n14032), .ZN(n14035) );
  OAI222_X1 U12963 ( .A1(n14422), .A2(n10951), .B1(n12358), .B2(n10950), .C1(
        P2_U3088), .C2(n14035), .ZN(P2_U3313) );
  NAND2_X1 U12964 ( .A1(n10953), .A2(n10952), .ZN(n10954) );
  XOR2_X1 U12965 ( .A(n10955), .B(n10954), .Z(n10960) );
  OAI21_X1 U12966 ( .B1(n14706), .B2(n11115), .A(n10956), .ZN(n10958) );
  NOR2_X1 U12967 ( .A1(n14701), .A2(n11117), .ZN(n10957) );
  AOI211_X1 U12968 ( .C1(n12729), .C2(n14709), .A(n10958), .B(n10957), .ZN(
        n10959) );
  OAI21_X1 U12969 ( .B1(n10960), .B2(n14711), .A(n10959), .ZN(P1_U3230) );
  OAI21_X1 U12970 ( .B1(n10962), .B2(n10965), .A(n10961), .ZN(n11530) );
  OAI211_X1 U12971 ( .C1(n11535), .C2(n10963), .A(n14348), .B(n11213), .ZN(
        n10964) );
  INV_X1 U12972 ( .A(n10964), .ZN(n11537) );
  XNOR2_X1 U12973 ( .A(n10966), .B(n10965), .ZN(n10968) );
  OAI21_X1 U12974 ( .B1(n10968), .B2(n14243), .A(n10967), .ZN(n11531) );
  AOI211_X1 U12975 ( .C1(n16033), .C2(n11530), .A(n11537), .B(n11531), .ZN(
        n11259) );
  AOI22_X1 U12976 ( .A1(n14300), .A2(n10969), .B1(n16034), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n10970) );
  OAI21_X1 U12977 ( .B1(n11259), .B2(n16034), .A(n10970), .ZN(P2_U3504) );
  INV_X1 U12978 ( .A(n10991), .ZN(n11181) );
  XNOR2_X1 U12979 ( .A(n10972), .B(n10978), .ZN(n11200) );
  AOI22_X1 U12980 ( .A1(n11200), .A2(P3_REG2_REG_5__SCAN_IN), .B1(n11206), 
        .B2(n10972), .ZN(n11169) );
  MUX2_X1 U12981 ( .A(n8288), .B(P3_REG2_REG_6__SCAN_IN), .S(n10991), .Z(
        n11168) );
  XNOR2_X1 U12982 ( .A(n11806), .B(n11820), .ZN(n11810) );
  XNOR2_X1 U12983 ( .A(n11810), .B(P3_REG2_REG_7__SCAN_IN), .ZN(n10999) );
  INV_X1 U12984 ( .A(n10973), .ZN(n10974) );
  NAND2_X1 U12985 ( .A1(n10974), .A2(n10985), .ZN(n10975) );
  MUX2_X1 U12986 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n13728), .Z(n10977) );
  NAND2_X1 U12987 ( .A1(n10977), .A2(n11206), .ZN(n11197) );
  NAND2_X1 U12988 ( .A1(n11199), .A2(n11197), .ZN(n10980) );
  INV_X1 U12989 ( .A(n10977), .ZN(n10979) );
  NAND2_X1 U12990 ( .A1(n10979), .A2(n10978), .ZN(n11196) );
  NAND2_X1 U12991 ( .A1(n10980), .A2(n11196), .ZN(n11166) );
  MUX2_X1 U12992 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n13728), .Z(n10981) );
  XNOR2_X1 U12993 ( .A(n10981), .B(n11181), .ZN(n11167) );
  NAND2_X1 U12994 ( .A1(n11166), .A2(n11167), .ZN(n10984) );
  INV_X1 U12995 ( .A(n10981), .ZN(n10982) );
  NAND2_X1 U12996 ( .A1(n10982), .A2(n11181), .ZN(n10983) );
  MUX2_X1 U12997 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n13728), .Z(n11788) );
  XNOR2_X1 U12998 ( .A(n11788), .B(n11808), .ZN(n11786) );
  XNOR2_X1 U12999 ( .A(n11787), .B(n11786), .ZN(n10997) );
  AND2_X1 U13000 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n11920) );
  AOI21_X1 U13001 ( .B1(n15806), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11920), .ZN(
        n10995) );
  OR2_X1 U13002 ( .A1(n10985), .A2(n15910), .ZN(n10986) );
  NAND2_X1 U13003 ( .A1(n10987), .A2(n10986), .ZN(n10988) );
  NAND2_X1 U13004 ( .A1(n10988), .A2(n11206), .ZN(n10989) );
  OAI21_X1 U13005 ( .B1(n10988), .B2(n11206), .A(n10989), .ZN(n11201) );
  NAND2_X1 U13006 ( .A1(n11203), .A2(n10989), .ZN(n11173) );
  INV_X1 U13007 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10990) );
  MUX2_X1 U13008 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n10990), .S(n10991), .Z(
        n11174) );
  NAND2_X1 U13009 ( .A1(n11173), .A2(n11174), .ZN(n11172) );
  NAND2_X1 U13010 ( .A1(n10991), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n10992) );
  NAND2_X1 U13011 ( .A1(n11172), .A2(n10992), .ZN(n11821) );
  XNOR2_X1 U13012 ( .A(n11821), .B(n11808), .ZN(n11819) );
  XNOR2_X1 U13013 ( .A(n11819), .B(P3_REG1_REG_7__SCAN_IN), .ZN(n10993) );
  NAND2_X1 U13014 ( .A1(n15819), .A2(n10993), .ZN(n10994) );
  OAI211_X1 U13015 ( .C1(n13362), .C2(n11820), .A(n10995), .B(n10994), .ZN(
        n10996) );
  AOI21_X1 U13016 ( .B1(n10997), .B2(n15814), .A(n10996), .ZN(n10998) );
  OAI21_X1 U13017 ( .B1(n10999), .B2(n15742), .A(n10998), .ZN(P3_U3189) );
  OAI21_X1 U13018 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n11001), .A(n11000), 
        .ZN(n11004) );
  MUX2_X1 U13019 ( .A(n9806), .B(P1_REG2_REG_13__SCAN_IN), .S(n11630), .Z(
        n11003) );
  INV_X1 U13020 ( .A(n11626), .ZN(n11002) );
  AOI211_X1 U13021 ( .C1(n11004), .C2(n11003), .A(n14811), .B(n11002), .ZN(
        n11013) );
  NAND2_X1 U13022 ( .A1(n11006), .A2(n11005), .ZN(n11008) );
  MUX2_X1 U13023 ( .A(n9805), .B(P1_REG1_REG_13__SCAN_IN), .S(n11630), .Z(
        n11007) );
  NOR2_X1 U13024 ( .A1(n11008), .A2(n11007), .ZN(n11629) );
  AOI211_X1 U13025 ( .C1(n11008), .C2(n11007), .A(n11897), .B(n11629), .ZN(
        n11012) );
  NAND2_X1 U13026 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n12396)
         );
  NAND2_X1 U13027 ( .A1(n15544), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n11009) );
  OAI211_X1 U13028 ( .C1(n15564), .C2(n11010), .A(n12396), .B(n11009), .ZN(
        n11011) );
  OR3_X1 U13029 ( .A1(n11013), .A2(n11012), .A3(n11011), .ZN(P1_U3256) );
  INV_X1 U13030 ( .A(n15972), .ZN(n15857) );
  INV_X1 U13031 ( .A(n11020), .ZN(n11193) );
  OAI22_X1 U13032 ( .A1(n11016), .A2(n13582), .B1(n11334), .B2(n13580), .ZN(
        n11017) );
  AOI21_X1 U13033 ( .B1(n11018), .B2(n15851), .A(n11017), .ZN(n11019) );
  OAI21_X1 U13034 ( .B1(n11020), .B2(n15855), .A(n11019), .ZN(n11192) );
  AOI21_X1 U13035 ( .B1(n15857), .B2(n11193), .A(n11192), .ZN(n11473) );
  INV_X1 U13036 ( .A(n13656), .ZN(n16045) );
  AOI22_X1 U13037 ( .A1(n16045), .A2(n11471), .B1(n8727), .B2(
        P3_REG1_REG_1__SCAN_IN), .ZN(n11021) );
  OAI21_X1 U13038 ( .B1(n11473), .B2(n8727), .A(n11021), .ZN(P3_U3460) );
  OAI21_X1 U13039 ( .B1(n11024), .B2(n11023), .A(n11022), .ZN(n11029) );
  OAI21_X1 U13040 ( .B1(n11027), .B2(n11026), .A(n11025), .ZN(n11028) );
  AOI22_X1 U13041 ( .A1(n15819), .A2(n11029), .B1(n15815), .B2(n11028), .ZN(
        n11037) );
  INV_X1 U13042 ( .A(n11030), .ZN(n11262) );
  INV_X1 U13043 ( .A(n11031), .ZN(n11033) );
  NOR3_X1 U13044 ( .A1(n11262), .A2(n11033), .A3(n11032), .ZN(n11035) );
  OAI21_X1 U13045 ( .B1(n11035), .B2(n11034), .A(n15814), .ZN(n11036) );
  OAI211_X1 U13046 ( .C1(n13362), .C2(n11038), .A(n11037), .B(n11036), .ZN(
        n11040) );
  OAI22_X1 U13047 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8203), .B1(n15585), .B2(
        n15787), .ZN(n11039) );
  OR2_X1 U13048 ( .A1(n11040), .A2(n11039), .ZN(P3_U3184) );
  XNOR2_X1 U13049 ( .A(n11041), .B(n12882), .ZN(n11355) );
  OAI21_X1 U13050 ( .B1(n11044), .B2(n11043), .A(n11042), .ZN(n11363) );
  INV_X1 U13051 ( .A(n11363), .ZN(n11049) );
  INV_X1 U13052 ( .A(n15992), .ZN(n16008) );
  NAND2_X1 U13053 ( .A1(n14704), .A2(n14736), .ZN(n11046) );
  NAND2_X1 U13054 ( .A1(n14702), .A2(n14738), .ZN(n11045) );
  NAND2_X1 U13055 ( .A1(n11046), .A2(n11045), .ZN(n11496) );
  INV_X1 U13056 ( .A(n11496), .ZN(n11356) );
  AOI21_X1 U13057 ( .B1(n12749), .B2(n11047), .A(n15985), .ZN(n11048) );
  NAND2_X1 U13058 ( .A1(n11456), .A2(n11048), .ZN(n11361) );
  OAI211_X1 U13059 ( .C1(n11049), .C2(n16008), .A(n11356), .B(n11361), .ZN(
        n11050) );
  AOI21_X1 U13060 ( .B1(n16013), .B2(n11355), .A(n11050), .ZN(n11054) );
  OAI22_X1 U13061 ( .A1(n11499), .A2(n15402), .B1(n16017), .B2(n9716), .ZN(
        n11051) );
  INV_X1 U13062 ( .A(n11051), .ZN(n11052) );
  OAI21_X1 U13063 ( .B1(n11054), .B2(n7917), .A(n11052), .ZN(P1_U3480) );
  AOI22_X1 U13064 ( .A1(n12749), .A2(n10229), .B1(n7362), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n11053) );
  OAI21_X1 U13065 ( .B1(n11054), .B2(n7362), .A(n11053), .ZN(P1_U3535) );
  INV_X1 U13066 ( .A(n11055), .ZN(n11056) );
  NAND2_X1 U13067 ( .A1(n11057), .A2(n11056), .ZN(n11058) );
  XNOR2_X1 U13068 ( .A(n11218), .B(n13764), .ZN(n11060) );
  AND2_X1 U13069 ( .A1(n13926), .A2(n8098), .ZN(n11061) );
  NAND2_X1 U13070 ( .A1(n11060), .A2(n11061), .ZN(n11379) );
  INV_X1 U13071 ( .A(n11060), .ZN(n11063) );
  INV_X1 U13072 ( .A(n11061), .ZN(n11062) );
  NAND2_X1 U13073 ( .A1(n11063), .A2(n11062), .ZN(n11064) );
  AND2_X1 U13074 ( .A1(n11379), .A2(n11064), .ZN(n11065) );
  OAI211_X1 U13075 ( .C1(n11066), .C2(n11065), .A(n11380), .B(n13881), .ZN(
        n11073) );
  OR2_X1 U13076 ( .A1(n11391), .A2(n14237), .ZN(n11069) );
  OR2_X1 U13077 ( .A1(n11067), .A2(n14235), .ZN(n11068) );
  AND2_X1 U13078 ( .A1(n11069), .A2(n11068), .ZN(n11216) );
  INV_X1 U13079 ( .A(n11216), .ZN(n11071) );
  NAND2_X1 U13080 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n13962) );
  OAI21_X1 U13081 ( .B1(n13902), .B2(n11463), .A(n13962), .ZN(n11070) );
  AOI21_X1 U13082 ( .B1(n13872), .B2(n11071), .A(n11070), .ZN(n11072) );
  OAI211_X1 U13083 ( .C1(n11462), .C2(n13889), .A(n11073), .B(n11072), .ZN(
        P2_U3211) );
  OAI21_X1 U13084 ( .B1(n11075), .B2(n11079), .A(n11074), .ZN(n15918) );
  INV_X1 U13085 ( .A(n11076), .ZN(n11078) );
  AOI211_X1 U13086 ( .C1(n12738), .C2(n11078), .A(n15985), .B(n7661), .ZN(
        n15911) );
  XNOR2_X1 U13087 ( .A(n11080), .B(n11079), .ZN(n11081) );
  NOR2_X1 U13088 ( .A1(n11081), .A2(n15987), .ZN(n11082) );
  AOI211_X1 U13089 ( .C1(n15837), .C2(n15918), .A(n11083), .B(n11082), .ZN(
        n15920) );
  INV_X1 U13090 ( .A(n15920), .ZN(n11084) );
  AOI211_X1 U13091 ( .C1(n15926), .C2(n15918), .A(n15911), .B(n11084), .ZN(
        n11089) );
  INV_X1 U13092 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n11085) );
  OAI22_X1 U13093 ( .A1(n15402), .A2(n15916), .B1(n16017), .B2(n11085), .ZN(
        n11086) );
  INV_X1 U13094 ( .A(n11086), .ZN(n11087) );
  OAI21_X1 U13095 ( .B1(n11089), .B2(n7917), .A(n11087), .ZN(P1_U3474) );
  AOI22_X1 U13096 ( .A1(n10229), .A2(n12738), .B1(n7362), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n11088) );
  OAI21_X1 U13097 ( .B1(n11089), .B2(n7362), .A(n11088), .ZN(P1_U3533) );
  INV_X1 U13098 ( .A(n11102), .ZN(n11090) );
  NAND2_X1 U13099 ( .A1(n11111), .A2(n11090), .ZN(n11093) );
  NAND2_X1 U13100 ( .A1(n11106), .A2(n11101), .ZN(n11091) );
  NAND4_X1 U13101 ( .A1(n11093), .A2(n11092), .A3(n11091), .A4(n11184), .ZN(
        n11094) );
  NAND2_X1 U13102 ( .A1(n11094), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11100) );
  INV_X1 U13103 ( .A(n11095), .ZN(n11096) );
  NAND2_X1 U13104 ( .A1(n11109), .A2(n11096), .ZN(n12696) );
  INV_X1 U13105 ( .A(n12696), .ZN(n11098) );
  INV_X1 U13106 ( .A(n12700), .ZN(n11097) );
  AOI21_X1 U13107 ( .B1(n11111), .B2(n11098), .A(n11097), .ZN(n11099) );
  NOR2_X1 U13108 ( .A1(n13230), .A2(P3_U3151), .ZN(n11327) );
  NAND2_X1 U13109 ( .A1(n11101), .A2(n15970), .ZN(n11103) );
  OAI22_X1 U13110 ( .A1(n11106), .A2(n11103), .B1(n11111), .B2(n11102), .ZN(
        n11104) );
  INV_X1 U13111 ( .A(n12660), .ZN(n11113) );
  NAND2_X1 U13112 ( .A1(n11109), .A2(n15907), .ZN(n11105) );
  OR2_X1 U13113 ( .A1(n11106), .A2(n11105), .ZN(n11108) );
  INV_X1 U13114 ( .A(n15861), .ZN(n11190) );
  NOR2_X1 U13115 ( .A1(n15970), .A2(n11190), .ZN(n11107) );
  INV_X1 U13116 ( .A(n13190), .ZN(n13234) );
  NAND2_X1 U13117 ( .A1(n11109), .A2(n12654), .ZN(n11110) );
  NOR2_X1 U13118 ( .A1(n11111), .A2(n11110), .ZN(n11318) );
  OAI22_X1 U13119 ( .A1(n11413), .A2(n13234), .B1(n13217), .B2(n11316), .ZN(
        n11112) );
  AOI21_X1 U13120 ( .B1(n13223), .B2(n11113), .A(n11112), .ZN(n11114) );
  OAI21_X1 U13121 ( .B1(n11327), .B2(n8216), .A(n11114), .ZN(P3_U3172) );
  INV_X1 U13122 ( .A(n15000), .ZN(n15024) );
  INV_X1 U13123 ( .A(n12729), .ZN(n11121) );
  MUX2_X1 U13124 ( .A(n11116), .B(n11115), .S(n15054), .Z(n11120) );
  INV_X1 U13125 ( .A(n15051), .ZN(n15938) );
  INV_X1 U13126 ( .A(n11117), .ZN(n11118) );
  NAND2_X1 U13127 ( .A1(n15938), .A2(n11118), .ZN(n11119) );
  OAI211_X1 U13128 ( .C1(n11121), .C2(n15942), .A(n11120), .B(n11119), .ZN(
        n11124) );
  AND2_X1 U13129 ( .A1(n11122), .A2(n15935), .ZN(n11123) );
  AOI211_X1 U13130 ( .C1(n11125), .C2(n15022), .A(n11124), .B(n11123), .ZN(
        n11126) );
  OAI21_X1 U13131 ( .B1(n11127), .B2(n15024), .A(n11126), .ZN(P1_U3289) );
  NAND2_X1 U13132 ( .A1(n11137), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n11128) );
  AND2_X1 U13133 ( .A1(n11129), .A2(n11128), .ZN(n14010) );
  INV_X1 U13134 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11130) );
  MUX2_X1 U13135 ( .A(n11130), .B(P2_REG2_REG_11__SCAN_IN), .S(n14015), .Z(
        n14009) );
  NAND2_X1 U13136 ( .A1(n14010), .A2(n14009), .ZN(n15518) );
  NAND2_X1 U13137 ( .A1(n14015), .A2(n11130), .ZN(n15516) );
  NAND2_X1 U13138 ( .A1(n15518), .A2(n15516), .ZN(n11131) );
  MUX2_X1 U13139 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n12009), .S(n15522), .Z(
        n15515) );
  NAND2_X1 U13140 ( .A1(n11131), .A2(n15515), .ZN(n15520) );
  OR2_X1 U13141 ( .A1(n15522), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n11132) );
  NAND2_X1 U13142 ( .A1(n15520), .A2(n11132), .ZN(n15504) );
  MUX2_X1 U13143 ( .A(n12136), .B(P2_REG2_REG_13__SCAN_IN), .S(n15507), .Z(
        n15503) );
  NAND2_X1 U13144 ( .A1(n15507), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11133) );
  MUX2_X1 U13145 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n14024), .S(n14032), .Z(
        n11134) );
  NAND2_X1 U13146 ( .A1(n14025), .A2(n11134), .ZN(n14027) );
  OR2_X1 U13147 ( .A1(n14032), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n11135) );
  NAND2_X1 U13148 ( .A1(n14027), .A2(n11135), .ZN(n11601) );
  XOR2_X1 U13149 ( .A(n11610), .B(n11601), .Z(n11603) );
  INV_X1 U13150 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n12377) );
  XNOR2_X1 U13151 ( .A(n11603), .B(n12377), .ZN(n11150) );
  INV_X1 U13152 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15697) );
  NAND2_X1 U13153 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n12412)
         );
  OAI21_X1 U13154 ( .B1(n15534), .B2(n15697), .A(n12412), .ZN(n11136) );
  AOI21_X1 U13155 ( .B1(n11610), .B2(n15521), .A(n11136), .ZN(n11149) );
  NAND2_X1 U13156 ( .A1(n11137), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n14017) );
  NAND2_X1 U13157 ( .A1(n14018), .A2(n14017), .ZN(n11140) );
  MUX2_X1 U13158 ( .A(n11138), .B(P2_REG1_REG_11__SCAN_IN), .S(n14015), .Z(
        n11139) );
  NAND2_X1 U13159 ( .A1(n11140), .A2(n11139), .ZN(n14020) );
  INV_X1 U13160 ( .A(n14015), .ZN(n14014) );
  NAND2_X1 U13161 ( .A1(n14014), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n11141) );
  NAND2_X1 U13162 ( .A1(n14020), .A2(n11141), .ZN(n15526) );
  MUX2_X1 U13163 ( .A(n11142), .B(P2_REG1_REG_12__SCAN_IN), .S(n15522), .Z(
        n15525) );
  NOR2_X1 U13164 ( .A1(n15526), .A2(n15525), .ZN(n15529) );
  AOI21_X1 U13165 ( .B1(n11142), .B2(n11143), .A(n15529), .ZN(n15510) );
  MUX2_X1 U13166 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n11144), .S(n15507), .Z(
        n15509) );
  NAND2_X1 U13167 ( .A1(n15510), .A2(n15509), .ZN(n15508) );
  NAND2_X1 U13168 ( .A1(n15507), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n14034) );
  NAND2_X1 U13169 ( .A1(n15508), .A2(n14034), .ZN(n11146) );
  NAND2_X1 U13170 ( .A1(n14032), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n11145) );
  OAI211_X1 U13171 ( .C1(n14032), .C2(P2_REG1_REG_14__SCAN_IN), .A(n11146), 
        .B(n11145), .ZN(n14036) );
  OAI21_X1 U13172 ( .B1(n9122), .B2(n14035), .A(n14036), .ZN(n11609) );
  INV_X1 U13173 ( .A(n11610), .ZN(n11602) );
  XNOR2_X1 U13174 ( .A(n11609), .B(n11602), .ZN(n11147) );
  NAND2_X1 U13175 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n11147), .ZN(n11611) );
  OAI211_X1 U13176 ( .C1(n11147), .C2(P2_REG1_REG_15__SCAN_IN), .A(n15527), 
        .B(n11611), .ZN(n11148) );
  OAI211_X1 U13177 ( .C1(n11150), .C2(n15502), .A(n11149), .B(n11148), .ZN(
        P2_U3229) );
  XNOR2_X1 U13178 ( .A(n11152), .B(n12874), .ZN(n11154) );
  AOI21_X1 U13179 ( .B1(n11154), .B2(n16013), .A(n11153), .ZN(n15840) );
  NAND2_X1 U13180 ( .A1(n11155), .A2(n15835), .ZN(n11156) );
  NAND2_X1 U13181 ( .A1(n11156), .A2(n15878), .ZN(n11157) );
  NOR2_X1 U13182 ( .A1(n15879), .A2(n11157), .ZN(n15834) );
  OAI22_X1 U13183 ( .A1(n15054), .A2(n11159), .B1(n11158), .B2(n15051), .ZN(
        n11162) );
  NOR2_X1 U13184 ( .A1(n15942), .A2(n11160), .ZN(n11161) );
  AOI211_X1 U13185 ( .C1(n15834), .C2(n15935), .A(n11162), .B(n11161), .ZN(
        n11165) );
  XNOR2_X1 U13186 ( .A(n12874), .B(n11163), .ZN(n15836) );
  NAND2_X1 U13187 ( .A1(n15022), .A2(n15836), .ZN(n11164) );
  OAI211_X1 U13188 ( .C1(n15895), .C2(n15840), .A(n11165), .B(n11164), .ZN(
        P1_U3292) );
  XOR2_X1 U13189 ( .A(n11167), .B(n11166), .Z(n11183) );
  NAND2_X1 U13190 ( .A1(n11169), .A2(n11168), .ZN(n11170) );
  AOI21_X1 U13191 ( .B1(n11171), .B2(n11170), .A(n15742), .ZN(n11180) );
  INV_X1 U13192 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n11178) );
  OAI21_X1 U13193 ( .B1(n11174), .B2(n11173), .A(n11172), .ZN(n11175) );
  NAND2_X1 U13194 ( .A1(n15819), .A2(n11175), .ZN(n11177) );
  INV_X1 U13195 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n15252) );
  NOR2_X1 U13196 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15252), .ZN(n11726) );
  INV_X1 U13197 ( .A(n11726), .ZN(n11176) );
  OAI211_X1 U13198 ( .C1(n15787), .C2(n11178), .A(n11177), .B(n11176), .ZN(
        n11179) );
  AOI211_X1 U13199 ( .C1(n15808), .C2(n11181), .A(n11180), .B(n11179), .ZN(
        n11182) );
  OAI21_X1 U13200 ( .B1(n11183), .B2(n15763), .A(n11182), .ZN(P3_U3188) );
  INV_X1 U13201 ( .A(n11184), .ZN(n11185) );
  NOR2_X1 U13202 ( .A1(n13709), .A2(n11185), .ZN(n11187) );
  MUX2_X1 U13203 ( .A(n13709), .B(n11187), .S(n11186), .Z(n11188) );
  NAND2_X1 U13204 ( .A1(n15907), .A2(n11190), .ZN(n11407) );
  OAI22_X1 U13205 ( .A1(n15860), .A2(n8223), .B1(n11326), .B2(n11407), .ZN(
        n11191) );
  OAI21_X1 U13206 ( .B1(n11192), .B2(n11191), .A(n15867), .ZN(n11195) );
  NAND2_X1 U13207 ( .A1(n12536), .A2(n15861), .ZN(n11841) );
  INV_X1 U13208 ( .A(n11841), .ZN(n15866) );
  NAND2_X1 U13209 ( .A1(n13500), .A2(n11193), .ZN(n11194) );
  OAI211_X1 U13210 ( .C1(n10878), .C2(n15867), .A(n11195), .B(n11194), .ZN(
        P3_U3232) );
  NAND2_X1 U13211 ( .A1(n11197), .A2(n11196), .ZN(n11198) );
  XNOR2_X1 U13212 ( .A(n11199), .B(n11198), .ZN(n11210) );
  XNOR2_X1 U13213 ( .A(n11200), .B(P3_REG2_REG_5__SCAN_IN), .ZN(n11208) );
  AND2_X1 U13214 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n13128) );
  NAND2_X1 U13215 ( .A1(n11201), .A2(n8267), .ZN(n11202) );
  AOI21_X1 U13216 ( .B1(n11203), .B2(n11202), .A(n15800), .ZN(n11204) );
  AOI211_X1 U13217 ( .C1(n15806), .C2(P3_ADDR_REG_5__SCAN_IN), .A(n13128), .B(
        n11204), .ZN(n11205) );
  OAI21_X1 U13218 ( .B1(n11206), .B2(n13362), .A(n11205), .ZN(n11207) );
  AOI21_X1 U13219 ( .B1(n15815), .B2(n11208), .A(n11207), .ZN(n11209) );
  OAI21_X1 U13220 ( .B1(n15763), .B2(n11210), .A(n11209), .ZN(P3_U3187) );
  OAI21_X1 U13221 ( .B1(n11212), .B2(n11214), .A(n11211), .ZN(n11467) );
  AOI211_X1 U13222 ( .C1(n11218), .C2(n11213), .A(n14282), .B(n11344), .ZN(
        n11466) );
  XNOR2_X1 U13223 ( .A(n11215), .B(n11214), .ZN(n11217) );
  OAI21_X1 U13224 ( .B1(n11217), .B2(n14243), .A(n11216), .ZN(n11461) );
  AOI211_X1 U13225 ( .C1(n16033), .C2(n11467), .A(n11466), .B(n11461), .ZN(
        n11256) );
  AOI22_X1 U13226 ( .A1(n14300), .A2(n11218), .B1(n16034), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n11219) );
  OAI21_X1 U13227 ( .B1(n11256), .B2(n16034), .A(n11219), .ZN(P2_U3505) );
  XNOR2_X1 U13228 ( .A(n11220), .B(n12876), .ZN(n15896) );
  NAND2_X1 U13229 ( .A1(n11221), .A2(n10000), .ZN(n12869) );
  INV_X1 U13230 ( .A(n12869), .ZN(n11222) );
  NAND2_X1 U13231 ( .A1(n15054), .A2(n11222), .ZN(n14857) );
  OR2_X1 U13232 ( .A1(n15896), .A2(n15874), .ZN(n11228) );
  OAI21_X1 U13233 ( .B1(n11224), .B2(n12876), .A(n11223), .ZN(n11226) );
  AOI21_X1 U13234 ( .B1(n11226), .B2(n16013), .A(n11225), .ZN(n11227) );
  NAND2_X1 U13235 ( .A1(n11228), .A2(n11227), .ZN(n15899) );
  INV_X2 U13236 ( .A(n15054), .ZN(n15895) );
  MUX2_X1 U13237 ( .A(n15899), .B(P1_REG2_REG_3__SCAN_IN), .S(n15895), .Z(
        n11229) );
  INV_X1 U13238 ( .A(n11229), .ZN(n11234) );
  OAI22_X1 U13239 ( .A1(n15942), .A2(n15898), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n15051), .ZN(n11232) );
  OAI211_X1 U13240 ( .C1(n15898), .C2(n15881), .A(n15878), .B(n11230), .ZN(
        n15897) );
  NOR2_X1 U13241 ( .A1(n15057), .A2(n15897), .ZN(n11231) );
  NOR2_X1 U13242 ( .A1(n11232), .A2(n11231), .ZN(n11233) );
  OAI211_X1 U13243 ( .C1(n15896), .C2(n14857), .A(n11234), .B(n11233), .ZN(
        P1_U3290) );
  INV_X1 U13244 ( .A(n11235), .ZN(n11236) );
  OAI222_X1 U13245 ( .A1(P3_U3151), .A2(n11308), .B1(n13730), .B2(n11236), 
        .C1(n15191), .C2(n13723), .ZN(P3_U3275) );
  INV_X1 U13246 ( .A(n11238), .ZN(n11240) );
  AND3_X1 U13247 ( .A1(n15455), .A2(n11240), .A3(n11239), .ZN(n11241) );
  NAND2_X1 U13248 ( .A1(n15454), .A2(n11241), .ZN(n11247) );
  NAND2_X1 U13249 ( .A1(n11242), .A2(n12085), .ZN(n11588) );
  NAND2_X1 U13250 ( .A1(n14279), .A2(n11588), .ZN(n11370) );
  INV_X1 U13251 ( .A(n14255), .ZN(n14285) );
  AOI22_X1 U13252 ( .A1(n11243), .A2(n11370), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n14285), .ZN(n11244) );
  INV_X2 U13253 ( .A(n14280), .ZN(n14265) );
  AOI21_X1 U13254 ( .B1(n11245), .B2(n11244), .A(n14265), .ZN(n11246) );
  AOI21_X1 U13255 ( .B1(n14265), .B2(P2_REG2_REG_0__SCAN_IN), .A(n11246), .ZN(
        n11252) );
  INV_X1 U13256 ( .A(n11247), .ZN(n11248) );
  AND2_X1 U13257 ( .A1(n14290), .A2(n14151), .ZN(n14201) );
  OAI21_X1 U13258 ( .B1(n14201), .B2(n14258), .A(n11250), .ZN(n11251) );
  NAND2_X1 U13259 ( .A1(n11252), .A2(n11251), .ZN(P2_U3265) );
  INV_X1 U13260 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n11253) );
  OAI22_X1 U13261 ( .A1(n14402), .A2(n11462), .B1(n14371), .B2(n11253), .ZN(
        n11254) );
  INV_X1 U13262 ( .A(n11254), .ZN(n11255) );
  OAI21_X1 U13263 ( .B1(n11256), .B2(n16001), .A(n11255), .ZN(P2_U3448) );
  OAI22_X1 U13264 ( .A1(n14402), .A2(n11535), .B1(n14371), .B2(n8903), .ZN(
        n11257) );
  INV_X1 U13265 ( .A(n11257), .ZN(n11258) );
  OAI21_X1 U13266 ( .B1(n11259), .B2(n16001), .A(n11258), .ZN(P2_U3445) );
  OAI21_X1 U13267 ( .B1(P3_REG2_REG_1__SCAN_IN), .B2(n11261), .A(n11260), .ZN(
        n11270) );
  AOI21_X1 U13268 ( .B1(n11263), .B2(n15743), .A(n11262), .ZN(n11264) );
  NOR2_X1 U13269 ( .A1(n11264), .A2(n15763), .ZN(n11269) );
  NAND2_X1 U13270 ( .A1(n11265), .A2(n10877), .ZN(n11266) );
  AOI21_X1 U13271 ( .B1(n11267), .B2(n11266), .A(n15800), .ZN(n11268) );
  AOI211_X1 U13272 ( .C1(n15815), .C2(n11270), .A(n11269), .B(n11268), .ZN(
        n11273) );
  OAI22_X1 U13273 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8223), .B1(n15576), .B2(
        n15787), .ZN(n11271) );
  INV_X1 U13274 ( .A(n11271), .ZN(n11272) );
  OAI211_X1 U13275 ( .C1(n13362), .C2(n11274), .A(n11273), .B(n11272), .ZN(
        P3_U3183) );
  INV_X1 U13276 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11275) );
  NOR2_X1 U13277 ( .A1(n16042), .A2(n11275), .ZN(n11276) );
  AOI21_X1 U13278 ( .B1(n16042), .B2(n11409), .A(n11276), .ZN(n11277) );
  OAI21_X1 U13279 ( .B1(n11413), .B2(n13707), .A(n11277), .ZN(P3_U3390) );
  INV_X1 U13280 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n11278) );
  OAI22_X1 U13281 ( .A1(n14402), .A2(n11415), .B1(n14371), .B2(n11278), .ZN(
        n11279) );
  INV_X1 U13282 ( .A(n11279), .ZN(n11280) );
  OAI21_X1 U13283 ( .B1(n11281), .B2(n16001), .A(n11280), .ZN(P2_U3439) );
  INV_X1 U13284 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n11282) );
  OAI22_X1 U13285 ( .A1(n14402), .A2(n11374), .B1(n14371), .B2(n11282), .ZN(
        n11283) );
  INV_X1 U13286 ( .A(n11283), .ZN(n11284) );
  OAI21_X1 U13287 ( .B1(n11285), .B2(n16001), .A(n11284), .ZN(P2_U3436) );
  INV_X1 U13288 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n11286) );
  OAI22_X1 U13289 ( .A1(n14402), .A2(n11503), .B1(n14371), .B2(n11286), .ZN(
        n11287) );
  INV_X1 U13290 ( .A(n11287), .ZN(n11288) );
  OAI21_X1 U13291 ( .B1(n11289), .B2(n16001), .A(n11288), .ZN(P2_U3433) );
  INV_X1 U13292 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11291) );
  INV_X1 U13293 ( .A(n11290), .ZN(n11292) );
  OAI222_X1 U13294 ( .A1(n14422), .A2(n11291), .B1(n12358), .B2(n11292), .C1(
        n11602), .C2(P2_U3088), .ZN(P2_U3312) );
  INV_X1 U13295 ( .A(n14790), .ZN(n14801) );
  OAI222_X1 U13296 ( .A1(n15435), .A2(n11293), .B1(n15437), .B2(n11292), .C1(
        n14801), .C2(P1_U3086), .ZN(P1_U3340) );
  NAND2_X1 U13297 ( .A1(n12741), .A2(n14532), .ZN(n11298) );
  NAND2_X1 U13298 ( .A1(n14442), .A2(n14738), .ZN(n11297) );
  NAND2_X1 U13299 ( .A1(n11298), .A2(n11297), .ZN(n11299) );
  XNOR2_X1 U13300 ( .A(n11299), .B(n14586), .ZN(n11484) );
  NOR2_X1 U13301 ( .A1(n14588), .A2(n12743), .ZN(n11300) );
  AOI21_X1 U13302 ( .B1(n12741), .B2(n14442), .A(n11300), .ZN(n11482) );
  XNOR2_X1 U13303 ( .A(n11484), .B(n11482), .ZN(n11301) );
  OAI211_X1 U13304 ( .C1(n7294), .C2(n11301), .A(n11485), .B(n14690), .ZN(
        n11306) );
  AND2_X1 U13305 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n14777) );
  NOR2_X1 U13306 ( .A1(n14701), .A2(n11302), .ZN(n11303) );
  AOI211_X1 U13307 ( .C1(n14671), .C2(n11304), .A(n14777), .B(n11303), .ZN(
        n11305) );
  OAI211_X1 U13308 ( .C1(n12742), .C2(n14698), .A(n11306), .B(n11305), .ZN(
        P1_U3239) );
  NAND2_X1 U13309 ( .A1(n11309), .A2(n11308), .ZN(n11310) );
  XNOR2_X1 U13310 ( .A(n11431), .B(n11334), .ZN(n11434) );
  OAI21_X1 U13311 ( .B1(n12986), .B2(n11314), .A(n11313), .ZN(n11325) );
  XOR2_X1 U13312 ( .A(n11434), .B(n11317), .Z(n11322) );
  OAI22_X1 U13313 ( .A1(n13234), .A2(n15845), .B1(n13217), .B2(n11662), .ZN(
        n11320) );
  NOR2_X1 U13314 ( .A1(n11327), .A2(n8203), .ZN(n11319) );
  AOI211_X1 U13315 ( .C1(n13215), .C2(n7349), .A(n11320), .B(n11319), .ZN(
        n11321) );
  OAI21_X1 U13316 ( .B1(n13196), .B2(n11322), .A(n11321), .ZN(P3_U3177) );
  XOR2_X1 U13317 ( .A(n11325), .B(n11324), .Z(n11331) );
  OAI22_X1 U13318 ( .A1(n11326), .A2(n13234), .B1(n13217), .B2(n11334), .ZN(
        n11329) );
  NOR2_X1 U13319 ( .A1(n11327), .A2(n8223), .ZN(n11328) );
  OAI21_X1 U13320 ( .B1(n11331), .B2(n13196), .A(n11330), .ZN(P3_U3162) );
  AOI21_X1 U13321 ( .B1(n11333), .B2(n12658), .A(n13578), .ZN(n11337) );
  OAI22_X1 U13322 ( .A1(n11334), .A2(n13582), .B1(n11856), .B2(n13580), .ZN(
        n11335) );
  AOI21_X1 U13323 ( .B1(n11337), .B2(n11336), .A(n11335), .ZN(n11844) );
  INV_X1 U13324 ( .A(n11844), .ZN(n11338) );
  AOI21_X1 U13325 ( .B1(n13658), .B2(n11843), .A(n11338), .ZN(n11443) );
  AOI22_X1 U13326 ( .A1(n16045), .A2(n11846), .B1(n8727), .B2(
        P3_REG1_REG_3__SCAN_IN), .ZN(n11339) );
  OAI21_X1 U13327 ( .B1(n11443), .B2(n8727), .A(n11339), .ZN(P3_U3462) );
  INV_X1 U13328 ( .A(n11340), .ZN(n11341) );
  AOI21_X1 U13329 ( .B1(n11343), .B2(n11342), .A(n11341), .ZN(n11544) );
  OAI21_X1 U13330 ( .B1(n11344), .B2(n11546), .A(n14348), .ZN(n11345) );
  NOR2_X1 U13331 ( .A1(n11345), .A2(n11397), .ZN(n11548) );
  XNOR2_X1 U13332 ( .A(n11347), .B(n11346), .ZN(n11350) );
  OAI22_X1 U13333 ( .A1(n11348), .A2(n14235), .B1(n11644), .B2(n14237), .ZN(
        n11384) );
  INV_X1 U13334 ( .A(n11384), .ZN(n11349) );
  OAI21_X1 U13335 ( .B1(n11350), .B2(n14243), .A(n11349), .ZN(n11549) );
  AOI211_X1 U13336 ( .C1(n11544), .C2(n16033), .A(n11548), .B(n11549), .ZN(
        n11354) );
  AOI22_X1 U13337 ( .A1(n14300), .A2(n11387), .B1(n16034), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n11351) );
  OAI21_X1 U13338 ( .B1(n11354), .B2(n16034), .A(n11351), .ZN(P2_U3506) );
  OAI22_X1 U13339 ( .A1(n14402), .A2(n11546), .B1(n14371), .B2(n8949), .ZN(
        n11352) );
  INV_X1 U13340 ( .A(n11352), .ZN(n11353) );
  OAI21_X1 U13341 ( .B1(n11354), .B2(n16001), .A(n11353), .ZN(P2_U3451) );
  INV_X1 U13342 ( .A(n11355), .ZN(n11365) );
  MUX2_X1 U13343 ( .A(n11357), .B(n11356), .S(n15054), .Z(n11358) );
  OAI21_X1 U13344 ( .B1(n15051), .B2(n11493), .A(n11358), .ZN(n11359) );
  AOI21_X1 U13345 ( .B1(n15887), .B2(n12749), .A(n11359), .ZN(n11360) );
  OAI21_X1 U13346 ( .B1(n11361), .B2(n15057), .A(n11360), .ZN(n11362) );
  AOI21_X1 U13347 ( .B1(n11363), .B2(n15022), .A(n11362), .ZN(n11364) );
  OAI21_X1 U13348 ( .B1(n11365), .B2(n15024), .A(n11364), .ZN(P1_U3286) );
  INV_X1 U13349 ( .A(n11366), .ZN(n11369) );
  OAI222_X1 U13350 ( .A1(n13730), .A2(n11369), .B1(n13723), .B2(n11368), .C1(
        P3_U3151), .C2(n11367), .ZN(P3_U3274) );
  MUX2_X1 U13351 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n11371), .S(n14280), .Z(
        n11376) );
  AOI22_X1 U13352 ( .A1(n11372), .A2(n14290), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n14285), .ZN(n11373) );
  OAI21_X1 U13353 ( .B1(n11374), .B2(n14288), .A(n11373), .ZN(n11375) );
  AOI211_X1 U13354 ( .C1(n14263), .C2(n11377), .A(n11376), .B(n11375), .ZN(
        n11378) );
  INV_X1 U13355 ( .A(n11378), .ZN(P2_U3263) );
  XNOR2_X1 U13356 ( .A(n11546), .B(n13773), .ZN(n11637) );
  NOR2_X1 U13357 ( .A1(n11391), .A2(n14348), .ZN(n11638) );
  XNOR2_X1 U13358 ( .A(n11637), .B(n11638), .ZN(n11383) );
  INV_X1 U13359 ( .A(n11642), .ZN(n11381) );
  AOI21_X1 U13360 ( .B1(n11383), .B2(n11382), .A(n11381), .ZN(n11389) );
  NAND2_X1 U13361 ( .A1(n13872), .A2(n11384), .ZN(n11385) );
  NAND2_X1 U13362 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n13977) );
  OAI211_X1 U13363 ( .C1(n13902), .C2(n11545), .A(n11385), .B(n13977), .ZN(
        n11386) );
  AOI21_X1 U13364 ( .B1(n11387), .B2(n13905), .A(n11386), .ZN(n11388) );
  OAI21_X1 U13365 ( .B1(n11389), .B2(n13907), .A(n11388), .ZN(P2_U3185) );
  INV_X1 U13366 ( .A(n11655), .ZN(n11396) );
  XNOR2_X1 U13367 ( .A(n11390), .B(n8025), .ZN(n11395) );
  OR2_X1 U13368 ( .A1(n11391), .A2(n14235), .ZN(n11393) );
  NAND2_X1 U13369 ( .A1(n13923), .A2(n14275), .ZN(n11392) );
  NAND2_X1 U13370 ( .A1(n11393), .A2(n11392), .ZN(n11653) );
  INV_X1 U13371 ( .A(n11653), .ZN(n11394) );
  OAI21_X1 U13372 ( .B1(n11395), .B2(n14243), .A(n11394), .ZN(n11474) );
  AOI21_X1 U13373 ( .B1(n11396), .B2(n14285), .A(n11474), .ZN(n11406) );
  INV_X1 U13374 ( .A(n11397), .ZN(n11399) );
  INV_X1 U13375 ( .A(n11398), .ZN(n11596) );
  AOI211_X1 U13376 ( .C1(n11657), .C2(n11399), .A(n8098), .B(n11596), .ZN(
        n11475) );
  OAI22_X1 U13377 ( .A1(n11643), .A2(n14288), .B1(n14280), .B2(n11400), .ZN(
        n11401) );
  AOI21_X1 U13378 ( .B1(n11475), .B2(n14290), .A(n11401), .ZN(n11405) );
  XNOR2_X1 U13379 ( .A(n11403), .B(n11402), .ZN(n11476) );
  NAND2_X1 U13380 ( .A1(n11476), .A2(n14263), .ZN(n11404) );
  OAI211_X1 U13381 ( .C1(n11406), .C2(n14265), .A(n11405), .B(n11404), .ZN(
        P2_U3257) );
  OR2_X2 U13382 ( .A1(n11408), .A2(n11407), .ZN(n13587) );
  AOI21_X1 U13383 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n13541), .A(n11409), .ZN(
        n11410) );
  MUX2_X1 U13384 ( .A(n11411), .B(n11410), .S(n15867), .Z(n11412) );
  OAI21_X1 U13385 ( .B1(n11413), .B2(n13587), .A(n11412), .ZN(P3_U3233) );
  INV_X1 U13386 ( .A(n11414), .ZN(n11422) );
  OAI22_X1 U13387 ( .A1(n14280), .A2(n10476), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n14255), .ZN(n11417) );
  NOR2_X1 U13388 ( .A1(n14288), .A2(n11415), .ZN(n11416) );
  AOI211_X1 U13389 ( .C1(n11418), .C2(n14290), .A(n11417), .B(n11416), .ZN(
        n11421) );
  NAND2_X1 U13390 ( .A1(n11419), .A2(n14263), .ZN(n11420) );
  OAI211_X1 U13391 ( .C1(n14265), .C2(n11422), .A(n11421), .B(n11420), .ZN(
        P2_U3262) );
  INV_X1 U13392 ( .A(n11423), .ZN(n11426) );
  OAI222_X1 U13393 ( .A1(n15435), .A2(n11424), .B1(n15437), .B2(n11426), .C1(
        n15563), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U13394 ( .A(n11674), .ZN(n11622) );
  INV_X1 U13395 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11425) );
  OAI222_X1 U13396 ( .A1(P2_U3088), .A2(n11622), .B1(n12358), .B2(n11426), 
        .C1(n11425), .C2(n14422), .ZN(P2_U3311) );
  NAND2_X1 U13397 ( .A1(n13215), .A2(n13252), .ZN(n11429) );
  AOI21_X1 U13398 ( .B1(n13190), .B2(n11846), .A(n11427), .ZN(n11428) );
  OAI211_X1 U13399 ( .C1(n11856), .C2(n13217), .A(n11429), .B(n11428), .ZN(
        n11438) );
  XNOR2_X1 U13400 ( .A(n12986), .B(n11846), .ZN(n11717) );
  XNOR2_X1 U13401 ( .A(n11717), .B(n11662), .ZN(n11436) );
  INV_X1 U13402 ( .A(n11431), .ZN(n11432) );
  AOI211_X1 U13403 ( .C1(n11436), .C2(n11435), .A(n13196), .B(n11718), .ZN(
        n11437) );
  AOI211_X1 U13404 ( .C1(n15169), .C2(n13230), .A(n11438), .B(n11437), .ZN(
        n11439) );
  INV_X1 U13405 ( .A(n11439), .ZN(P3_U3158) );
  OAI22_X1 U13406 ( .A1(n13707), .A2(n11440), .B1(n16042), .B2(n8241), .ZN(
        n11441) );
  INV_X1 U13407 ( .A(n11441), .ZN(n11442) );
  OAI21_X1 U13408 ( .B1(n11443), .B2(n16048), .A(n11442), .ZN(P3_U3399) );
  OR2_X1 U13409 ( .A1(n11444), .A2(n12884), .ZN(n11445) );
  NAND2_X1 U13410 ( .A1(n11446), .A2(n11445), .ZN(n15925) );
  INV_X1 U13411 ( .A(n15925), .ZN(n11460) );
  XNOR2_X1 U13412 ( .A(n11448), .B(n11447), .ZN(n11453) );
  NAND2_X1 U13413 ( .A1(n15925), .A2(n15837), .ZN(n11452) );
  NAND2_X1 U13414 ( .A1(n14704), .A2(n14735), .ZN(n11450) );
  NAND2_X1 U13415 ( .A1(n14702), .A2(n14737), .ZN(n11449) );
  NAND2_X1 U13416 ( .A1(n11450), .A2(n11449), .ZN(n11766) );
  INV_X1 U13417 ( .A(n11766), .ZN(n11451) );
  OAI211_X1 U13418 ( .C1(n15987), .C2(n11453), .A(n11452), .B(n11451), .ZN(
        n15924) );
  MUX2_X1 U13419 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n15924), .S(n15054), .Z(
        n11454) );
  INV_X1 U13420 ( .A(n11454), .ZN(n11459) );
  AOI211_X1 U13421 ( .C1(n12753), .C2(n11456), .A(n15985), .B(n11455), .ZN(
        n15921) );
  OAI22_X1 U13422 ( .A1(n7659), .A2(n15942), .B1(n11768), .B2(n15051), .ZN(
        n11457) );
  AOI21_X1 U13423 ( .B1(n15921), .B2(n15935), .A(n11457), .ZN(n11458) );
  OAI211_X1 U13424 ( .C1(n11460), .C2(n14857), .A(n11459), .B(n11458), .ZN(
        P1_U3285) );
  INV_X1 U13425 ( .A(n11461), .ZN(n11470) );
  NOR2_X1 U13426 ( .A1(n11462), .A2(n14288), .ZN(n11465) );
  OAI22_X1 U13427 ( .A1(n14280), .A2(n10481), .B1(n11463), .B2(n14255), .ZN(
        n11464) );
  AOI211_X1 U13428 ( .C1(n11466), .C2(n14290), .A(n11465), .B(n11464), .ZN(
        n11469) );
  NAND2_X1 U13429 ( .A1(n11467), .A2(n14263), .ZN(n11468) );
  OAI211_X1 U13430 ( .C1(n14265), .C2(n11470), .A(n11469), .B(n11468), .ZN(
        P2_U3259) );
  INV_X1 U13431 ( .A(n13707), .ZN(n16049) );
  AOI22_X1 U13432 ( .A1(n16049), .A2(n11471), .B1(P3_REG0_REG_1__SCAN_IN), 
        .B2(n16048), .ZN(n11472) );
  OAI21_X1 U13433 ( .B1(n11473), .B2(n16048), .A(n11472), .ZN(P3_U3393) );
  AOI211_X1 U13434 ( .C1(n16033), .C2(n11476), .A(n11475), .B(n11474), .ZN(
        n11481) );
  INV_X1 U13435 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n11477) );
  OAI22_X1 U13436 ( .A1(n11643), .A2(n14402), .B1(n14398), .B2(n11477), .ZN(
        n11478) );
  INV_X1 U13437 ( .A(n11478), .ZN(n11479) );
  OAI21_X1 U13438 ( .B1(n11481), .B2(n16001), .A(n11479), .ZN(P2_U3454) );
  AOI22_X1 U13439 ( .A1(n11657), .A2(n14300), .B1(n16034), .B2(
        P2_REG1_REG_8__SCAN_IN), .ZN(n11480) );
  OAI21_X1 U13440 ( .B1(n11481), .B2(n16034), .A(n11480), .ZN(P2_U3507) );
  INV_X1 U13441 ( .A(n11482), .ZN(n11483) );
  NAND2_X1 U13442 ( .A1(n12749), .A2(n14532), .ZN(n11487) );
  NAND2_X1 U13443 ( .A1(n14442), .A2(n14737), .ZN(n11486) );
  NAND2_X1 U13444 ( .A1(n11487), .A2(n11486), .ZN(n11488) );
  XNOR2_X1 U13445 ( .A(n11488), .B(n14586), .ZN(n11760) );
  NOR2_X1 U13446 ( .A1(n14588), .A2(n11489), .ZN(n11490) );
  AOI21_X1 U13447 ( .B1(n12749), .B2(n14442), .A(n11490), .ZN(n11758) );
  XNOR2_X1 U13448 ( .A(n11760), .B(n11758), .ZN(n11491) );
  NAND2_X1 U13449 ( .A1(n11492), .A2(n11491), .ZN(n11762) );
  OAI211_X1 U13450 ( .C1(n11492), .C2(n11491), .A(n11762), .B(n14690), .ZN(
        n11498) );
  NOR2_X1 U13451 ( .A1(n14701), .A2(n11493), .ZN(n11494) );
  AOI211_X1 U13452 ( .C1(n14671), .C2(n11496), .A(n11495), .B(n11494), .ZN(
        n11497) );
  OAI211_X1 U13453 ( .C1(n11499), .C2(n14698), .A(n11498), .B(n11497), .ZN(
        P1_U3213) );
  MUX2_X1 U13454 ( .A(n11500), .B(P2_REG2_REG_1__SCAN_IN), .S(n14265), .Z(
        n11505) );
  AOI22_X1 U13455 ( .A1(n14290), .A2(n11501), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n14285), .ZN(n11502) );
  OAI21_X1 U13456 ( .B1(n14288), .B2(n11503), .A(n11502), .ZN(n11504) );
  AOI211_X1 U13457 ( .C1(n14263), .C2(n11506), .A(n11505), .B(n11504), .ZN(
        n11507) );
  INV_X1 U13458 ( .A(n11507), .ZN(P2_U3264) );
  OAI21_X1 U13459 ( .B1(n11509), .B2(n11511), .A(n11508), .ZN(n11566) );
  INV_X1 U13460 ( .A(n11510), .ZN(n11512) );
  NAND2_X1 U13461 ( .A1(n11512), .A2(n11511), .ZN(n11560) );
  NAND3_X1 U13462 ( .A1(n11560), .A2(n16013), .A3(n11559), .ZN(n11515) );
  NAND2_X1 U13463 ( .A1(n11699), .A2(n12764), .ZN(n11513) );
  AND3_X1 U13464 ( .A1(n11578), .A2(n15878), .A3(n11513), .ZN(n11556) );
  NAND2_X1 U13465 ( .A1(n14704), .A2(n14733), .ZN(n11555) );
  NAND2_X1 U13466 ( .A1(n14702), .A2(n14735), .ZN(n11561) );
  NAND2_X1 U13467 ( .A1(n11555), .A2(n11561), .ZN(n12161) );
  NOR2_X1 U13468 ( .A1(n11556), .A2(n12161), .ZN(n11514) );
  NAND2_X1 U13469 ( .A1(n11515), .A2(n11514), .ZN(n11516) );
  AOI21_X1 U13470 ( .B1(n15992), .B2(n11566), .A(n11516), .ZN(n11520) );
  OAI22_X1 U13471 ( .A1(n7671), .A2(n15402), .B1(n16017), .B2(n9759), .ZN(
        n11517) );
  INV_X1 U13472 ( .A(n11517), .ZN(n11518) );
  OAI21_X1 U13473 ( .B1(n11520), .B2(n7917), .A(n11518), .ZN(P1_U3489) );
  AOI22_X1 U13474 ( .A1(n12764), .A2(n10229), .B1(n7362), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n11519) );
  OAI21_X1 U13475 ( .B1(n11520), .B2(n7362), .A(n11519), .ZN(P1_U3538) );
  MUX2_X1 U13476 ( .A(n11522), .B(n11521), .S(n14280), .Z(n11528) );
  OAI22_X1 U13477 ( .A1(n14288), .A2(n11524), .B1(n11523), .B2(n14255), .ZN(
        n11525) );
  AOI21_X1 U13478 ( .B1(n11526), .B2(n14290), .A(n11525), .ZN(n11527) );
  OAI211_X1 U13479 ( .C1(n14198), .C2(n11529), .A(n11528), .B(n11527), .ZN(
        P2_U3261) );
  INV_X1 U13480 ( .A(n11530), .ZN(n11540) );
  INV_X1 U13481 ( .A(n11531), .ZN(n11532) );
  MUX2_X1 U13482 ( .A(n11533), .B(n11532), .S(n14280), .Z(n11539) );
  OAI22_X1 U13483 ( .A1(n14288), .A2(n11535), .B1(n14255), .B2(n11534), .ZN(
        n11536) );
  AOI21_X1 U13484 ( .B1(n14290), .B2(n11537), .A(n11536), .ZN(n11538) );
  OAI211_X1 U13485 ( .C1(n14198), .C2(n11540), .A(n11539), .B(n11538), .ZN(
        P2_U3260) );
  INV_X1 U13486 ( .A(n11541), .ZN(n11543) );
  OAI22_X1 U13487 ( .A1(n12697), .A2(P3_U3151), .B1(SI_22_), .B2(n13723), .ZN(
        n11542) );
  AOI21_X1 U13488 ( .B1(n11543), .B2(n13717), .A(n11542), .ZN(P3_U3273) );
  INV_X1 U13489 ( .A(n11544), .ZN(n11554) );
  OAI22_X1 U13490 ( .A1(n11546), .A2(n14288), .B1(n11545), .B2(n14255), .ZN(
        n11547) );
  AOI21_X1 U13491 ( .B1(n11548), .B2(n14290), .A(n11547), .ZN(n11553) );
  INV_X1 U13492 ( .A(n11549), .ZN(n11550) );
  MUX2_X1 U13493 ( .A(n11551), .B(n11550), .S(n14280), .Z(n11552) );
  OAI211_X1 U13494 ( .C1(n11554), .C2(n14198), .A(n11553), .B(n11552), .ZN(
        P2_U3258) );
  INV_X1 U13495 ( .A(n11555), .ZN(n11557) );
  AOI211_X1 U13496 ( .C1(n11566), .C2(n11558), .A(n11557), .B(n11556), .ZN(
        n11568) );
  INV_X1 U13497 ( .A(n14857), .ZN(n15946) );
  NAND3_X1 U13498 ( .A1(n11560), .A2(n15000), .A3(n11559), .ZN(n11564) );
  OAI22_X1 U13499 ( .A1(n15895), .A2(n11561), .B1(n12164), .B2(n15051), .ZN(
        n11562) );
  AOI21_X1 U13500 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n15895), .A(n11562), 
        .ZN(n11563) );
  OAI211_X1 U13501 ( .C1(n7671), .C2(n15942), .A(n11564), .B(n11563), .ZN(
        n11565) );
  AOI21_X1 U13502 ( .B1(n15946), .B2(n11566), .A(n11565), .ZN(n11567) );
  OAI21_X1 U13503 ( .B1(n11568), .B2(n15057), .A(n11567), .ZN(P1_U3283) );
  INV_X1 U13504 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11570) );
  INV_X1 U13505 ( .A(n11569), .ZN(n11571) );
  INV_X1 U13506 ( .A(n11693), .ZN(n12089) );
  OAI222_X1 U13507 ( .A1(n14422), .A2(n11570), .B1(n12358), .B2(n11571), .C1(
        P2_U3088), .C2(n12089), .ZN(P2_U3310) );
  INV_X1 U13508 ( .A(n15540), .ZN(n14794) );
  OAI222_X1 U13509 ( .A1(n15435), .A2(n11572), .B1(n15437), .B2(n11571), .C1(
        P1_U3086), .C2(n14794), .ZN(P1_U3338) );
  NAND2_X1 U13510 ( .A1(n13240), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n11573) );
  OAI21_X1 U13511 ( .B1(n13397), .B2(n13240), .A(n11573), .ZN(P3_U3519) );
  OAI21_X1 U13512 ( .B1(n11575), .B2(n12888), .A(n11574), .ZN(n11576) );
  OAI22_X1 U13513 ( .A1(n12320), .A2(n14607), .B1(n14605), .B2(n12158), .ZN(
        n12309) );
  AOI21_X1 U13514 ( .B1(n11576), .B2(n16013), .A(n12309), .ZN(n11924) );
  INV_X1 U13515 ( .A(n11868), .ZN(n11577) );
  AOI211_X1 U13516 ( .C1(n12773), .C2(n11578), .A(n15985), .B(n11577), .ZN(
        n11926) );
  NOR2_X1 U13517 ( .A1(n11930), .A2(n15942), .ZN(n11581) );
  OAI22_X1 U13518 ( .A1(n15054), .A2(n11579), .B1(n12311), .B2(n15051), .ZN(
        n11580) );
  AOI211_X1 U13519 ( .C1(n11926), .C2(n15935), .A(n11581), .B(n11580), .ZN(
        n11586) );
  NAND2_X1 U13520 ( .A1(n11582), .A2(n12888), .ZN(n11583) );
  AND2_X1 U13521 ( .A1(n11584), .A2(n11583), .ZN(n11927) );
  NAND2_X1 U13522 ( .A1(n11927), .A2(n15022), .ZN(n11585) );
  OAI211_X1 U13523 ( .C1(n15895), .C2(n11924), .A(n11586), .B(n11585), .ZN(
        P1_U3282) );
  XNOR2_X1 U13524 ( .A(n11587), .B(n8022), .ZN(n15949) );
  INV_X1 U13525 ( .A(n11588), .ZN(n11589) );
  NAND2_X1 U13526 ( .A1(n14280), .A2(n11589), .ZN(n14293) );
  XNOR2_X1 U13527 ( .A(n11590), .B(n8022), .ZN(n11593) );
  OAI22_X1 U13528 ( .A1(n11591), .A2(n14237), .B1(n11644), .B2(n14235), .ZN(
        n11592) );
  AOI21_X1 U13529 ( .B1(n11593), .B2(n14271), .A(n11592), .ZN(n11594) );
  OAI21_X1 U13530 ( .B1(n15949), .B2(n14279), .A(n11594), .ZN(n15952) );
  NAND2_X1 U13531 ( .A1(n15952), .A2(n14280), .ZN(n11600) );
  OAI22_X1 U13532 ( .A1(n14280), .A2(n11595), .B1(n11749), .B2(n14255), .ZN(
        n11598) );
  OAI211_X1 U13533 ( .C1(n15951), .C2(n11596), .A(n14348), .B(n11774), .ZN(
        n15950) );
  NOR2_X1 U13534 ( .A1(n15950), .A2(n14261), .ZN(n11597) );
  AOI211_X1 U13535 ( .C1(n14258), .C2(n11742), .A(n11598), .B(n11597), .ZN(
        n11599) );
  OAI211_X1 U13536 ( .C1(n15949), .C2(n14293), .A(n11600), .B(n11599), .ZN(
        P2_U3256) );
  OAI22_X1 U13537 ( .A1(n11603), .A2(n12377), .B1(n11602), .B2(n11601), .ZN(
        n11608) );
  INV_X1 U13538 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11605) );
  NAND2_X1 U13539 ( .A1(n11674), .A2(n11605), .ZN(n11604) );
  OAI21_X1 U13540 ( .B1(n11674), .B2(n11605), .A(n11604), .ZN(n11607) );
  NAND2_X1 U13541 ( .A1(n11622), .A2(n11605), .ZN(n11606) );
  OAI211_X1 U13542 ( .C1(n11605), .C2(n11622), .A(n11608), .B(n11606), .ZN(
        n11677) );
  OAI211_X1 U13543 ( .C1(n11608), .C2(n11607), .A(n11677), .B(n15523), .ZN(
        n11621) );
  NAND2_X1 U13544 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n12453)
         );
  INV_X1 U13545 ( .A(n12453), .ZN(n11619) );
  OR2_X1 U13546 ( .A1(n11674), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n11613) );
  NAND2_X1 U13547 ( .A1(n11674), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n11684) );
  NAND2_X1 U13548 ( .A1(n11610), .A2(n11609), .ZN(n11612) );
  NAND2_X1 U13549 ( .A1(n11612), .A2(n11611), .ZN(n11615) );
  NAND3_X1 U13550 ( .A1(n11613), .A2(n11684), .A3(n11615), .ZN(n11685) );
  INV_X1 U13551 ( .A(n11685), .ZN(n11689) );
  INV_X1 U13552 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n11616) );
  NOR2_X1 U13553 ( .A1(n11674), .A2(n11616), .ZN(n11614) );
  AOI211_X1 U13554 ( .C1(n11674), .C2(n11616), .A(n11615), .B(n11614), .ZN(
        n11617) );
  NOR3_X1 U13555 ( .A1(n15488), .A2(n11689), .A3(n11617), .ZN(n11618) );
  AOI211_X1 U13556 ( .C1(n15501), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n11619), 
        .B(n11618), .ZN(n11620) );
  OAI211_X1 U13557 ( .C1(n12095), .C2(n11622), .A(n11621), .B(n11620), .ZN(
        P2_U3230) );
  INV_X1 U13558 ( .A(n11888), .ZN(n11892) );
  NAND2_X1 U13559 ( .A1(n11630), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11625) );
  INV_X1 U13560 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11623) );
  MUX2_X1 U13561 ( .A(n11623), .B(P1_REG2_REG_14__SCAN_IN), .S(n11888), .Z(
        n11624) );
  AOI21_X1 U13562 ( .B1(n11626), .B2(n11625), .A(n11624), .ZN(n11887) );
  INV_X1 U13563 ( .A(n11887), .ZN(n11628) );
  NAND3_X1 U13564 ( .A1(n11626), .A2(n11625), .A3(n11624), .ZN(n11627) );
  NAND3_X1 U13565 ( .A1(n11628), .A2(n15558), .A3(n11627), .ZN(n11635) );
  NAND2_X1 U13566 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14558)
         );
  AOI21_X1 U13567 ( .B1(n11630), .B2(P1_REG1_REG_13__SCAN_IN), .A(n11629), 
        .ZN(n11893) );
  XOR2_X1 U13568 ( .A(n11888), .B(n11893), .Z(n11895) );
  XNOR2_X1 U13569 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n11895), .ZN(n11631) );
  NAND2_X1 U13570 ( .A1(n15566), .A2(n11631), .ZN(n11632) );
  NAND2_X1 U13571 ( .A1(n14558), .A2(n11632), .ZN(n11633) );
  AOI21_X1 U13572 ( .B1(n15544), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n11633), 
        .ZN(n11634) );
  OAI211_X1 U13573 ( .C1(n15564), .C2(n11892), .A(n11635), .B(n11634), .ZN(
        P1_U3257) );
  NAND2_X1 U13574 ( .A1(n13240), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n11636) );
  OAI21_X1 U13575 ( .B1(n13031), .B2(n13240), .A(n11636), .ZN(P3_U3520) );
  INV_X1 U13576 ( .A(n11637), .ZN(n11640) );
  INV_X1 U13577 ( .A(n11638), .ZN(n11639) );
  NAND2_X1 U13578 ( .A1(n11640), .A2(n11639), .ZN(n11641) );
  XNOR2_X1 U13579 ( .A(n11643), .B(n13805), .ZN(n11645) );
  OR2_X1 U13580 ( .A1(n11644), .A2(n14151), .ZN(n11646) );
  NAND2_X1 U13581 ( .A1(n11645), .A2(n11646), .ZN(n11650) );
  INV_X1 U13582 ( .A(n11645), .ZN(n11648) );
  INV_X1 U13583 ( .A(n11646), .ZN(n11647) );
  NAND2_X1 U13584 ( .A1(n11648), .A2(n11647), .ZN(n11649) );
  NAND2_X1 U13585 ( .A1(n7291), .A2(n11649), .ZN(n11651) );
  AOI22_X1 U13586 ( .A1(n11652), .A2(n11651), .B1(n11745), .B2(n11650), .ZN(
        n11659) );
  NAND2_X1 U13587 ( .A1(n13872), .A2(n11653), .ZN(n11654) );
  NAND2_X1 U13588 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n13992) );
  OAI211_X1 U13589 ( .C1(n13902), .C2(n11655), .A(n11654), .B(n13992), .ZN(
        n11656) );
  AOI21_X1 U13590 ( .B1(n11657), .B2(n13905), .A(n11656), .ZN(n11658) );
  OAI21_X1 U13591 ( .B1(n11659), .B2(n13907), .A(n11658), .ZN(P2_U3193) );
  OAI21_X1 U13592 ( .B1(n11661), .B2(n12663), .A(n11660), .ZN(n11669) );
  INV_X1 U13593 ( .A(n11669), .ZN(n11712) );
  INV_X1 U13594 ( .A(n15855), .ZN(n15977) );
  OAI22_X1 U13595 ( .A1(n11724), .A2(n13580), .B1(n11662), .B2(n13582), .ZN(
        n11668) );
  OAI211_X1 U13596 ( .C1(n11665), .C2(n11664), .A(n11663), .B(n15851), .ZN(
        n11666) );
  INV_X1 U13597 ( .A(n11666), .ZN(n11667) );
  AOI211_X1 U13598 ( .C1(n15977), .C2(n11669), .A(n11668), .B(n11667), .ZN(
        n11711) );
  MUX2_X1 U13599 ( .A(n11670), .B(n11711), .S(n15867), .Z(n11673) );
  INV_X1 U13600 ( .A(n13587), .ZN(n13557) );
  INV_X1 U13601 ( .A(n11671), .ZN(n13158) );
  AOI22_X1 U13602 ( .A1(n13557), .A2(n15906), .B1(n13541), .B2(n13158), .ZN(
        n11672) );
  OAI211_X1 U13603 ( .C1(n11712), .C2(n12292), .A(n11673), .B(n11672), .ZN(
        P3_U3229) );
  INV_X1 U13604 ( .A(n11677), .ZN(n11681) );
  NAND2_X1 U13605 ( .A1(n11674), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n11676) );
  INV_X1 U13606 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n12082) );
  OR2_X1 U13607 ( .A1(n11693), .A2(n12082), .ZN(n11675) );
  OAI211_X1 U13608 ( .C1(n12089), .C2(P2_REG2_REG_17__SCAN_IN), .A(n11676), 
        .B(n11675), .ZN(n11680) );
  NAND2_X1 U13609 ( .A1(n11677), .A2(n11676), .ZN(n11679) );
  NAND2_X1 U13610 ( .A1(n12089), .A2(n12082), .ZN(n11678) );
  OAI211_X1 U13611 ( .C1(n12082), .C2(n12089), .A(n11679), .B(n11678), .ZN(
        n12081) );
  OAI211_X1 U13612 ( .C1(n11681), .C2(n11680), .A(n12081), .B(n15523), .ZN(
        n11695) );
  INV_X1 U13613 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n11691) );
  NAND2_X1 U13614 ( .A1(n11693), .A2(n11682), .ZN(n11683) );
  OAI211_X1 U13615 ( .C1(n11693), .C2(n11682), .A(n11683), .B(n11684), .ZN(
        n11688) );
  NAND2_X1 U13616 ( .A1(n11685), .A2(n11684), .ZN(n11687) );
  NAND2_X1 U13617 ( .A1(n11693), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n11686) );
  OAI211_X1 U13618 ( .C1(n11693), .C2(P2_REG1_REG_17__SCAN_IN), .A(n11687), 
        .B(n11686), .ZN(n12088) );
  OAI211_X1 U13619 ( .C1(n11689), .C2(n11688), .A(n15527), .B(n12088), .ZN(
        n11690) );
  NAND2_X1 U13620 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3088), .ZN(n13839)
         );
  OAI211_X1 U13621 ( .C1(n11691), .C2(n15534), .A(n11690), .B(n13839), .ZN(
        n11692) );
  AOI21_X1 U13622 ( .B1(n11693), .B2(n15521), .A(n11692), .ZN(n11694) );
  NAND2_X1 U13623 ( .A1(n11695), .A2(n11694), .ZN(P2_U3231) );
  OAI21_X1 U13624 ( .B1(n11698), .B2(n11697), .A(n11696), .ZN(n15945) );
  INV_X1 U13625 ( .A(n11699), .ZN(n11700) );
  AOI211_X1 U13626 ( .C1(n12760), .C2(n11701), .A(n15985), .B(n11700), .ZN(
        n15936) );
  OAI22_X1 U13627 ( .A1(n12158), .A2(n14607), .B1(n14605), .B2(n11756), .ZN(
        n12040) );
  XNOR2_X1 U13628 ( .A(n11702), .B(n12885), .ZN(n11703) );
  NOR2_X1 U13629 ( .A1(n11703), .A2(n15987), .ZN(n11704) );
  AOI211_X1 U13630 ( .C1(n15837), .C2(n15945), .A(n12040), .B(n11704), .ZN(
        n15948) );
  INV_X1 U13631 ( .A(n15948), .ZN(n11705) );
  AOI211_X1 U13632 ( .C1(n15926), .C2(n15945), .A(n15936), .B(n11705), .ZN(
        n11710) );
  INV_X1 U13633 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n11706) );
  OAI22_X1 U13634 ( .A1(n15943), .A2(n15402), .B1(n16017), .B2(n11706), .ZN(
        n11707) );
  INV_X1 U13635 ( .A(n11707), .ZN(n11708) );
  OAI21_X1 U13636 ( .B1(n11710), .B2(n7917), .A(n11708), .ZN(P1_U3486) );
  AOI22_X1 U13637 ( .A1(n12760), .A2(n10229), .B1(n7362), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n11709) );
  OAI21_X1 U13638 ( .B1(n11710), .B2(n7362), .A(n11709), .ZN(P1_U3537) );
  INV_X1 U13639 ( .A(n11711), .ZN(n15904) );
  NOR2_X1 U13640 ( .A1(n11712), .A2(n15972), .ZN(n15905) );
  OAI21_X1 U13641 ( .B1(n15904), .B2(n15905), .A(n16042), .ZN(n11714) );
  NAND2_X1 U13642 ( .A1(n16049), .A2(n15906), .ZN(n11713) );
  OAI211_X1 U13643 ( .C1(n16042), .C2(n8255), .A(n11714), .B(n11713), .ZN(
        P3_U3402) );
  NAND2_X1 U13644 ( .A1(n11715), .A2(n13717), .ZN(n11716) );
  OAI211_X1 U13645 ( .C1(n15294), .C2(n13723), .A(n11716), .B(n12700), .ZN(
        P3_U3272) );
  XNOR2_X1 U13646 ( .A(n12986), .B(n15906), .ZN(n11720) );
  INV_X1 U13647 ( .A(n11717), .ZN(n11719) );
  XNOR2_X1 U13648 ( .A(n11720), .B(n13251), .ZN(n13155) );
  XNOR2_X1 U13649 ( .A(n13053), .B(n13129), .ZN(n11721) );
  XNOR2_X1 U13650 ( .A(n11721), .B(n13250), .ZN(n13125) );
  XNOR2_X1 U13651 ( .A(n12986), .B(n12044), .ZN(n11913) );
  XNOR2_X1 U13652 ( .A(n11913), .B(n11918), .ZN(n11722) );
  OAI211_X1 U13653 ( .C1(n11723), .C2(n11722), .A(n11915), .B(n13223), .ZN(
        n11728) );
  INV_X1 U13654 ( .A(n13215), .ZN(n13227) );
  OAI22_X1 U13655 ( .A1(n13227), .A2(n11724), .B1(n12242), .B2(n13217), .ZN(
        n11725) );
  AOI211_X1 U13656 ( .C1(n11908), .C2(n13190), .A(n11726), .B(n11725), .ZN(
        n11727) );
  OAI211_X1 U13657 ( .C1(n12043), .C2(n13175), .A(n11728), .B(n11727), .ZN(
        P3_U3179) );
  XNOR2_X1 U13658 ( .A(n11729), .B(n7490), .ZN(n15963) );
  INV_X1 U13659 ( .A(n15963), .ZN(n11741) );
  AND2_X1 U13660 ( .A1(n11731), .A2(n11730), .ZN(n11732) );
  OAI21_X1 U13661 ( .B1(n12014), .B2(n11732), .A(n14271), .ZN(n11734) );
  INV_X1 U13662 ( .A(n12144), .ZN(n13920) );
  AOI22_X1 U13663 ( .A1(n13920), .A2(n14275), .B1(n14274), .B2(n13922), .ZN(
        n11733) );
  NAND2_X1 U13664 ( .A1(n11734), .A2(n11733), .ZN(n15968) );
  OAI21_X1 U13665 ( .B1(n15965), .B2(n11773), .A(n14348), .ZN(n11735) );
  OR2_X1 U13666 ( .A1(n11735), .A2(n12007), .ZN(n15964) );
  OAI22_X1 U13667 ( .A1(n14280), .A2(n11130), .B1(n11955), .B2(n14255), .ZN(
        n11736) );
  AOI21_X1 U13668 ( .B1(n11737), .B2(n14258), .A(n11736), .ZN(n11738) );
  OAI21_X1 U13669 ( .B1(n15964), .B2(n14261), .A(n11738), .ZN(n11739) );
  AOI21_X1 U13670 ( .B1(n15968), .B2(n14280), .A(n11739), .ZN(n11740) );
  OAI21_X1 U13671 ( .B1(n14198), .B2(n11741), .A(n11740), .ZN(P2_U3254) );
  XNOR2_X1 U13672 ( .A(n11742), .B(n13764), .ZN(n11875) );
  NAND2_X1 U13673 ( .A1(n13923), .A2(n8098), .ZN(n11876) );
  XNOR2_X1 U13674 ( .A(n11875), .B(n11876), .ZN(n11744) );
  OAI21_X1 U13675 ( .B1(n11745), .B2(n11744), .A(n11879), .ZN(n11746) );
  NAND2_X1 U13676 ( .A1(n11746), .A2(n13881), .ZN(n11752) );
  NOR2_X2 U13677 ( .A1(n13900), .A2(n14235), .ZN(n13892) );
  NAND2_X1 U13678 ( .A1(n13887), .A2(n13922), .ZN(n11748) );
  OAI211_X1 U13679 ( .C1(n13902), .C2(n11749), .A(n11748), .B(n11747), .ZN(
        n11750) );
  AOI21_X1 U13680 ( .B1(n13892), .B2(n13924), .A(n11750), .ZN(n11751) );
  OAI211_X1 U13681 ( .C1(n15951), .C2(n13889), .A(n11752), .B(n11751), .ZN(
        P2_U3203) );
  NAND2_X1 U13682 ( .A1(n12753), .A2(n14532), .ZN(n11754) );
  NAND2_X1 U13683 ( .A1(n14442), .A2(n14736), .ZN(n11753) );
  NAND2_X1 U13684 ( .A1(n11754), .A2(n11753), .ZN(n11755) );
  XNOR2_X1 U13685 ( .A(n11755), .B(n14522), .ZN(n12028) );
  NOR2_X1 U13686 ( .A1(n14588), .A2(n11756), .ZN(n11757) );
  AOI21_X1 U13687 ( .B1(n12753), .B2(n14442), .A(n11757), .ZN(n12027) );
  XNOR2_X1 U13688 ( .A(n12028), .B(n12027), .ZN(n11765) );
  INV_X1 U13689 ( .A(n11758), .ZN(n11759) );
  NAND2_X1 U13690 ( .A1(n11760), .A2(n11759), .ZN(n11761) );
  INV_X1 U13691 ( .A(n12030), .ZN(n11763) );
  AOI21_X1 U13692 ( .B1(n11765), .B2(n11764), .A(n11763), .ZN(n11771) );
  AOI22_X1 U13693 ( .A1(n14671), .A2(n11766), .B1(P1_REG3_REG_8__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11767) );
  OAI21_X1 U13694 ( .B1(n14701), .B2(n11768), .A(n11767), .ZN(n11769) );
  AOI21_X1 U13695 ( .B1(n12753), .B2(n14709), .A(n11769), .ZN(n11770) );
  OAI21_X1 U13696 ( .B1(n11771), .B2(n14711), .A(n11770), .ZN(P1_U3221) );
  XNOR2_X1 U13697 ( .A(n11772), .B(n11779), .ZN(n11934) );
  AOI211_X1 U13698 ( .C1(n11938), .C2(n11774), .A(n8098), .B(n11773), .ZN(
        n11936) );
  NOR2_X1 U13699 ( .A1(n7597), .A2(n14288), .ZN(n11777) );
  OAI22_X1 U13700 ( .A1(n14280), .A2(n11775), .B1(n11881), .B2(n14255), .ZN(
        n11776) );
  AOI211_X1 U13701 ( .C1(n11936), .C2(n14290), .A(n11777), .B(n11776), .ZN(
        n11785) );
  XNOR2_X1 U13702 ( .A(n11779), .B(n11778), .ZN(n11782) );
  OAI22_X1 U13703 ( .A1(n11780), .A2(n14235), .B1(n11948), .B2(n14237), .ZN(
        n11781) );
  AOI21_X1 U13704 ( .B1(n11782), .B2(n14271), .A(n11781), .ZN(n11783) );
  OAI21_X1 U13705 ( .B1(n11934), .B2(n14279), .A(n11783), .ZN(n11935) );
  NAND2_X1 U13706 ( .A1(n11935), .A2(n14280), .ZN(n11784) );
  OAI211_X1 U13707 ( .C1(n11934), .C2(n14293), .A(n11785), .B(n11784), .ZN(
        P2_U3255) );
  NAND2_X1 U13708 ( .A1(n11787), .A2(n11786), .ZN(n11791) );
  INV_X1 U13709 ( .A(n11788), .ZN(n11789) );
  NAND2_X1 U13710 ( .A1(n11789), .A2(n11808), .ZN(n11790) );
  NAND2_X1 U13711 ( .A1(n11791), .A2(n11790), .ZN(n15750) );
  MUX2_X1 U13712 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n13728), .Z(n11792) );
  XNOR2_X1 U13713 ( .A(n11792), .B(n15755), .ZN(n15751) );
  INV_X1 U13714 ( .A(n11792), .ZN(n11793) );
  NAND2_X1 U13715 ( .A1(n11793), .A2(n15755), .ZN(n11794) );
  MUX2_X1 U13716 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n13728), .Z(n11795) );
  XNOR2_X1 U13717 ( .A(n11795), .B(n15780), .ZN(n15769) );
  INV_X1 U13718 ( .A(n11795), .ZN(n11796) );
  MUX2_X1 U13719 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n13728), .Z(n11798) );
  XNOR2_X1 U13720 ( .A(n11798), .B(n11830), .ZN(n15790) );
  MUX2_X1 U13721 ( .A(n11800), .B(n11799), .S(n13728), .Z(n11801) );
  XNOR2_X1 U13722 ( .A(n11801), .B(n11814), .ZN(n15811) );
  INV_X1 U13723 ( .A(n11814), .ZN(n15807) );
  AOI22_X1 U13724 ( .A1(n15812), .A2(n15811), .B1(n15807), .B2(n11801), .ZN(
        n11805) );
  NOR2_X1 U13725 ( .A1(n12114), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n11802) );
  AOI21_X1 U13726 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n12114), .A(n11802), 
        .ZN(n11817) );
  NAND2_X1 U13727 ( .A1(n12114), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n12117) );
  OAI21_X1 U13728 ( .B1(n12114), .B2(P3_REG1_REG_12__SCAN_IN), .A(n12117), 
        .ZN(n11834) );
  INV_X1 U13729 ( .A(n11834), .ZN(n11803) );
  MUX2_X1 U13730 ( .A(n11817), .B(n11803), .S(n13728), .Z(n11804) );
  NAND2_X1 U13731 ( .A1(n11805), .A2(n11804), .ZN(n12116) );
  OAI211_X1 U13732 ( .C1(n11805), .C2(n11804), .A(n12116), .B(n15814), .ZN(
        n11840) );
  NAND2_X1 U13733 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n11830), .ZN(n11813) );
  AOI22_X1 U13734 ( .A1(n15789), .A2(n8353), .B1(P3_REG2_REG_10__SCAN_IN), 
        .B2(n11830), .ZN(n15794) );
  AOI22_X1 U13735 ( .A1(n15755), .A2(n12245), .B1(P3_REG2_REG_8__SCAN_IN), 
        .B2(n11825), .ZN(n15753) );
  INV_X1 U13736 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11809) );
  INV_X1 U13737 ( .A(n11806), .ZN(n11807) );
  OAI22_X1 U13738 ( .A1(n11810), .A2(n11809), .B1(n11808), .B2(n11807), .ZN(
        n15754) );
  NAND2_X1 U13739 ( .A1(n15753), .A2(n15754), .ZN(n15752) );
  OAI21_X1 U13740 ( .B1(n15755), .B2(n12245), .A(n15752), .ZN(n11811) );
  NAND2_X1 U13741 ( .A1(n11811), .A2(n11828), .ZN(n11812) );
  XNOR2_X1 U13742 ( .A(n11811), .B(n15780), .ZN(n15773) );
  NAND2_X1 U13743 ( .A1(P3_REG2_REG_9__SCAN_IN), .A2(n15773), .ZN(n15772) );
  NAND2_X1 U13744 ( .A1(n11815), .A2(n11814), .ZN(n11816) );
  XNOR2_X1 U13745 ( .A(n11815), .B(n15807), .ZN(n15810) );
  NAND2_X1 U13746 ( .A1(P3_REG2_REG_11__SCAN_IN), .A2(n15810), .ZN(n15809) );
  OAI21_X1 U13747 ( .B1(n11818), .B2(n11817), .A(n12123), .ZN(n11838) );
  NAND2_X1 U13748 ( .A1(n11819), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n11823) );
  NAND2_X1 U13749 ( .A1(n11821), .A2(n11820), .ZN(n11822) );
  NAND2_X1 U13750 ( .A1(n11823), .A2(n11822), .ZN(n15758) );
  INV_X1 U13751 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n11824) );
  MUX2_X1 U13752 ( .A(n11824), .B(P3_REG1_REG_8__SCAN_IN), .S(n15755), .Z(
        n15759) );
  NAND2_X1 U13753 ( .A1(n15758), .A2(n15759), .ZN(n15757) );
  NAND2_X1 U13754 ( .A1(n11825), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n11826) );
  NAND2_X1 U13755 ( .A1(n15757), .A2(n11826), .ZN(n11827) );
  XNOR2_X1 U13756 ( .A(n11827), .B(n15780), .ZN(n15775) );
  NAND2_X1 U13757 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n11830), .ZN(n11829) );
  OAI21_X1 U13758 ( .B1(n11830), .B2(P3_REG1_REG_10__SCAN_IN), .A(n11829), 
        .ZN(n15798) );
  NOR2_X1 U13759 ( .A1(n11831), .A2(n15807), .ZN(n11832) );
  NOR2_X1 U13760 ( .A1(n11833), .A2(n11834), .ZN(n12118) );
  AOI21_X1 U13761 ( .B1(n11834), .B2(n11833), .A(n12118), .ZN(n11835) );
  NOR2_X1 U13762 ( .A1(n15800), .A2(n11835), .ZN(n11837) );
  INV_X1 U13763 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n15669) );
  INV_X1 U13764 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n15165) );
  OR2_X1 U13765 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15165), .ZN(n13098) );
  OAI21_X1 U13766 ( .B1(n15787), .B2(n15669), .A(n13098), .ZN(n11836) );
  AOI211_X1 U13767 ( .C1(n15815), .C2(n11838), .A(n11837), .B(n11836), .ZN(
        n11839) );
  OAI211_X1 U13768 ( .C1(n13362), .C2(n12114), .A(n11840), .B(n11839), .ZN(
        P3_U3194) );
  NAND2_X1 U13769 ( .A1(n15855), .A2(n11841), .ZN(n11842) );
  INV_X1 U13770 ( .A(n13592), .ZN(n13532) );
  INV_X1 U13771 ( .A(n11843), .ZN(n11849) );
  MUX2_X1 U13772 ( .A(n11845), .B(n11844), .S(n15867), .Z(n11848) );
  AOI22_X1 U13773 ( .A1(n13557), .A2(n11846), .B1(n13541), .B2(n15169), .ZN(
        n11847) );
  OAI211_X1 U13774 ( .C1(n13532), .C2(n11849), .A(n11848), .B(n11847), .ZN(
        P3_U3230) );
  OAI21_X1 U13775 ( .B1(n11851), .B2(n12662), .A(n11850), .ZN(n12025) );
  INV_X1 U13776 ( .A(n11852), .ZN(n11853) );
  AOI21_X1 U13777 ( .B1(n12662), .B2(n11854), .A(n11853), .ZN(n11855) );
  OAI222_X1 U13778 ( .A1(n13580), .A2(n11918), .B1(n13582), .B2(n11856), .C1(
        n13578), .C2(n11855), .ZN(n12022) );
  AOI21_X1 U13779 ( .B1(n13658), .B2(n12025), .A(n12022), .ZN(n11860) );
  OAI22_X1 U13780 ( .A1(n13707), .A2(n12021), .B1(n16042), .B2(n8270), .ZN(
        n11857) );
  INV_X1 U13781 ( .A(n11857), .ZN(n11858) );
  OAI21_X1 U13782 ( .B1(n11860), .B2(n16048), .A(n11858), .ZN(P3_U3405) );
  AOI22_X1 U13783 ( .A1(n16045), .A2(n13129), .B1(n8727), .B2(
        P3_REG1_REG_5__SCAN_IN), .ZN(n11859) );
  OAI21_X1 U13784 ( .B1(n11860), .B2(n8727), .A(n11859), .ZN(P3_U3464) );
  OAI211_X1 U13785 ( .C1(n11863), .C2(n11862), .A(n11861), .B(n16013), .ZN(
        n11864) );
  AOI22_X1 U13786 ( .A1(n14704), .A2(n14731), .B1(n14702), .B2(n14733), .ZN(
        n12328) );
  NAND2_X1 U13787 ( .A1(n11864), .A2(n12328), .ZN(n11977) );
  INV_X1 U13788 ( .A(n11977), .ZN(n11874) );
  OAI21_X1 U13789 ( .B1(n11866), .B2(n12890), .A(n11865), .ZN(n11979) );
  INV_X1 U13790 ( .A(n12777), .ZN(n12333) );
  AOI211_X1 U13791 ( .C1(n12777), .C2(n11868), .A(n15985), .B(n11867), .ZN(
        n11978) );
  NAND2_X1 U13792 ( .A1(n11978), .A2(n15935), .ZN(n11871) );
  INV_X1 U13793 ( .A(n11869), .ZN(n12330) );
  AOI22_X1 U13794 ( .A1(n15895), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n12330), 
        .B2(n15938), .ZN(n11870) );
  OAI211_X1 U13795 ( .C1(n12333), .C2(n15942), .A(n11871), .B(n11870), .ZN(
        n11872) );
  AOI21_X1 U13796 ( .B1(n15022), .B2(n11979), .A(n11872), .ZN(n11873) );
  OAI21_X1 U13797 ( .B1(n15895), .B2(n11874), .A(n11873), .ZN(P1_U3281) );
  INV_X1 U13798 ( .A(n11875), .ZN(n11877) );
  NAND2_X1 U13799 ( .A1(n13922), .A2(n14282), .ZN(n11947) );
  XOR2_X1 U13800 ( .A(n11945), .B(n11944), .Z(n11886) );
  OAI21_X1 U13801 ( .B1(n13902), .B2(n11881), .A(n11880), .ZN(n11882) );
  AOI21_X1 U13802 ( .B1(n13892), .B2(n13923), .A(n11882), .ZN(n11883) );
  OAI21_X1 U13803 ( .B1(n11948), .B2(n13859), .A(n11883), .ZN(n11884) );
  AOI21_X1 U13804 ( .B1(n11938), .B2(n13905), .A(n11884), .ZN(n11885) );
  OAI21_X1 U13805 ( .B1(n11886), .B2(n13907), .A(n11885), .ZN(P2_U3189) );
  AOI21_X1 U13806 ( .B1(n11888), .B2(P1_REG2_REG_14__SCAN_IN), .A(n11887), 
        .ZN(n14802) );
  XNOR2_X1 U13807 ( .A(n14802), .B(n14801), .ZN(n11889) );
  NOR2_X1 U13808 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n11889), .ZN(n14800) );
  AOI21_X1 U13809 ( .B1(n11889), .B2(P1_REG2_REG_15__SCAN_IN), .A(n14800), 
        .ZN(n11901) );
  NOR2_X1 U13810 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14705), .ZN(n11891) );
  NOR2_X1 U13811 ( .A1(n15564), .A2(n14801), .ZN(n11890) );
  AOI211_X1 U13812 ( .C1(n15544), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n11891), 
        .B(n11890), .ZN(n11900) );
  INV_X1 U13813 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11894) );
  OAI22_X1 U13814 ( .A1(n11895), .A2(n11894), .B1(n11893), .B2(n11892), .ZN(
        n14789) );
  XNOR2_X1 U13815 ( .A(n14789), .B(n14790), .ZN(n11896) );
  NOR2_X1 U13816 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n11896), .ZN(n14791) );
  AOI21_X1 U13817 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n11896), .A(n14791), 
        .ZN(n11898) );
  OR2_X1 U13818 ( .A1(n11898), .A2(n11897), .ZN(n11899) );
  OAI211_X1 U13819 ( .C1(n11901), .C2(n14811), .A(n11900), .B(n11899), .ZN(
        P1_U3258) );
  OAI21_X1 U13820 ( .B1(n11903), .B2(n12661), .A(n11902), .ZN(n12048) );
  OAI211_X1 U13821 ( .C1(n11905), .C2(n8626), .A(n15851), .B(n11904), .ZN(
        n11907) );
  AOI22_X1 U13822 ( .A1(n15846), .A2(n13248), .B1(n13250), .B2(n15848), .ZN(
        n11906) );
  NAND2_X1 U13823 ( .A1(n11907), .A2(n11906), .ZN(n12045) );
  AOI21_X1 U13824 ( .B1(n13658), .B2(n12048), .A(n12045), .ZN(n11912) );
  AOI22_X1 U13825 ( .A1(n16045), .A2(n11908), .B1(n8727), .B2(
        P3_REG1_REG_6__SCAN_IN), .ZN(n11909) );
  OAI21_X1 U13826 ( .B1(n11912), .B2(n8727), .A(n11909), .ZN(P3_U3465) );
  OAI22_X1 U13827 ( .A1(n13707), .A2(n12044), .B1(n16042), .B2(n8291), .ZN(
        n11910) );
  INV_X1 U13828 ( .A(n11910), .ZN(n11911) );
  OAI21_X1 U13829 ( .B1(n11912), .B2(n16048), .A(n11911), .ZN(P3_U3408) );
  NAND2_X1 U13830 ( .A1(n11913), .A2(n13249), .ZN(n11914) );
  NAND2_X1 U13831 ( .A1(n11915), .A2(n11914), .ZN(n11917) );
  XNOR2_X1 U13832 ( .A(n13053), .B(n11994), .ZN(n11997) );
  XNOR2_X1 U13833 ( .A(n11997), .B(n13248), .ZN(n11916) );
  OAI211_X1 U13834 ( .C1(n11917), .C2(n11916), .A(n11999), .B(n13223), .ZN(
        n11922) );
  OAI22_X1 U13835 ( .A1(n13227), .A2(n11918), .B1(n12568), .B2(n13217), .ZN(
        n11919) );
  AOI211_X1 U13836 ( .C1(n11994), .C2(n13190), .A(n11920), .B(n11919), .ZN(
        n11921) );
  OAI211_X1 U13837 ( .C1(n12207), .C2(n13175), .A(n11922), .B(n11921), .ZN(
        P3_U3153) );
  AOI22_X1 U13838 ( .A1(n15547), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n15423), .ZN(n11923) );
  OAI21_X1 U13839 ( .B1(n11975), .B2(n15437), .A(n11923), .ZN(P1_U3337) );
  INV_X1 U13840 ( .A(n11924), .ZN(n11925) );
  AOI211_X1 U13841 ( .C1(n11927), .C2(n15992), .A(n11926), .B(n11925), .ZN(
        n11933) );
  AOI22_X1 U13842 ( .A1(n12773), .A2(n10229), .B1(n7362), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n11928) );
  OAI21_X1 U13843 ( .B1(n11933), .B2(n7362), .A(n11928), .ZN(P1_U3539) );
  INV_X1 U13844 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n11929) );
  OAI22_X1 U13845 ( .A1(n11930), .A2(n15402), .B1(n16017), .B2(n11929), .ZN(
        n11931) );
  INV_X1 U13846 ( .A(n11931), .ZN(n11932) );
  OAI21_X1 U13847 ( .B1(n11933), .B2(n7917), .A(n11932), .ZN(P1_U3492) );
  INV_X1 U13848 ( .A(n11934), .ZN(n11937) );
  AOI211_X1 U13849 ( .C1(n16024), .C2(n11937), .A(n11936), .B(n11935), .ZN(
        n11943) );
  AOI22_X1 U13850 ( .A1(n11938), .A2(n14300), .B1(n16034), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n11939) );
  OAI21_X1 U13851 ( .B1(n11943), .B2(n16034), .A(n11939), .ZN(P2_U3509) );
  INV_X1 U13852 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n11940) );
  OAI22_X1 U13853 ( .A1(n7597), .A2(n14402), .B1(n14371), .B2(n11940), .ZN(
        n11941) );
  INV_X1 U13854 ( .A(n11941), .ZN(n11942) );
  OAI21_X1 U13855 ( .B1(n11943), .B2(n16001), .A(n11942), .ZN(P2_U3460) );
  XNOR2_X1 U13856 ( .A(n15965), .B(n13773), .ZN(n11952) );
  INV_X1 U13857 ( .A(n11952), .ZN(n11950) );
  NOR2_X1 U13858 ( .A1(n11948), .A2(n14348), .ZN(n11951) );
  INV_X1 U13859 ( .A(n11951), .ZN(n11949) );
  NAND2_X1 U13860 ( .A1(n11950), .A2(n11949), .ZN(n12057) );
  NAND2_X1 U13861 ( .A1(n11952), .A2(n11951), .ZN(n12055) );
  NAND2_X1 U13862 ( .A1(n12057), .A2(n12055), .ZN(n11953) );
  XNOR2_X1 U13863 ( .A(n12056), .B(n11953), .ZN(n11959) );
  NAND2_X1 U13864 ( .A1(n13887), .A2(n13920), .ZN(n11954) );
  NAND2_X1 U13865 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n14012)
         );
  OAI211_X1 U13866 ( .C1(n13902), .C2(n11955), .A(n11954), .B(n14012), .ZN(
        n11957) );
  NOR2_X1 U13867 ( .A1(n15965), .A2(n13889), .ZN(n11956) );
  AOI211_X1 U13868 ( .C1(n13892), .C2(n13922), .A(n11957), .B(n11956), .ZN(
        n11958) );
  OAI21_X1 U13869 ( .B1(n11959), .B2(n13907), .A(n11958), .ZN(P2_U3208) );
  OAI21_X1 U13870 ( .B1(n11962), .B2(n11961), .A(n11960), .ZN(n15988) );
  OAI21_X1 U13871 ( .B1(n11964), .B2(n12891), .A(n11963), .ZN(n15991) );
  NAND2_X1 U13872 ( .A1(n15991), .A2(n15022), .ZN(n11974) );
  NAND2_X1 U13873 ( .A1(n15983), .A2(n11965), .ZN(n11966) );
  NAND2_X1 U13874 ( .A1(n12072), .A2(n11966), .ZN(n15986) );
  NAND2_X1 U13875 ( .A1(n14730), .A2(n14704), .ZN(n11968) );
  NAND2_X1 U13876 ( .A1(n14702), .A2(n14732), .ZN(n11967) );
  AND2_X1 U13877 ( .A1(n11968), .A2(n11967), .ZN(n15980) );
  NAND2_X1 U13878 ( .A1(n15938), .A2(n12395), .ZN(n11969) );
  OAI211_X1 U13879 ( .C1(n15986), .C2(n15036), .A(n15980), .B(n11969), .ZN(
        n11972) );
  OAI22_X1 U13880 ( .A1(n11970), .A2(n15942), .B1(n9806), .B2(n15054), .ZN(
        n11971) );
  AOI21_X1 U13881 ( .B1(n11972), .B2(n15054), .A(n11971), .ZN(n11973) );
  OAI211_X1 U13882 ( .C1(n15988), .C2(n15024), .A(n11974), .B(n11973), .ZN(
        P1_U3280) );
  INV_X1 U13883 ( .A(n15497), .ZN(n12090) );
  OAI222_X1 U13884 ( .A1(n14422), .A2(n11976), .B1(n12358), .B2(n11975), .C1(
        n12090), .C2(P2_U3088), .ZN(P2_U3309) );
  AOI211_X1 U13885 ( .C1(n15992), .C2(n11979), .A(n11978), .B(n11977), .ZN(
        n11985) );
  INV_X1 U13886 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11980) );
  OAI22_X1 U13887 ( .A1(n12333), .A2(n15402), .B1(n16017), .B2(n11980), .ZN(
        n11981) );
  INV_X1 U13888 ( .A(n11981), .ZN(n11982) );
  OAI21_X1 U13889 ( .B1(n11985), .B2(n7917), .A(n11982), .ZN(P1_U3495) );
  OAI22_X1 U13890 ( .A1(n12333), .A2(n15125), .B1(n16014), .B2(n9791), .ZN(
        n11983) );
  INV_X1 U13891 ( .A(n11983), .ZN(n11984) );
  OAI21_X1 U13892 ( .B1(n11985), .B2(n7362), .A(n11984), .ZN(P1_U3540) );
  OAI21_X1 U13893 ( .B1(n11987), .B2(n12659), .A(n11986), .ZN(n12212) );
  OAI211_X1 U13894 ( .C1(n11989), .C2(n12562), .A(n11988), .B(n15851), .ZN(
        n11991) );
  AOI22_X1 U13895 ( .A1(n13249), .A2(n15848), .B1(n15846), .B2(n13247), .ZN(
        n11990) );
  NAND2_X1 U13896 ( .A1(n11991), .A2(n11990), .ZN(n12209) );
  AOI21_X1 U13897 ( .B1(n13658), .B2(n12212), .A(n12209), .ZN(n11996) );
  OAI22_X1 U13898 ( .A1(n13707), .A2(n12208), .B1(n16042), .B2(n8306), .ZN(
        n11992) );
  INV_X1 U13899 ( .A(n11992), .ZN(n11993) );
  OAI21_X1 U13900 ( .B1(n11996), .B2(n16048), .A(n11993), .ZN(P3_U3411) );
  AOI22_X1 U13901 ( .A1(n16045), .A2(n11994), .B1(n8727), .B2(
        P3_REG1_REG_7__SCAN_IN), .ZN(n11995) );
  OAI21_X1 U13902 ( .B1(n11996), .B2(n8727), .A(n11995), .ZN(P3_U3466) );
  XNOR2_X1 U13903 ( .A(n13053), .B(n12569), .ZN(n12226) );
  XNOR2_X1 U13904 ( .A(n12226), .B(n12568), .ZN(n12000) );
  OAI211_X1 U13905 ( .C1(n12001), .C2(n12000), .A(n12228), .B(n13223), .ZN(
        n12005) );
  NAND2_X1 U13906 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n15766) );
  INV_X1 U13907 ( .A(n15766), .ZN(n12003) );
  OAI22_X1 U13908 ( .A1(n13227), .A2(n12242), .B1(n12285), .B2(n13217), .ZN(
        n12002) );
  AOI211_X1 U13909 ( .C1(n12269), .C2(n13190), .A(n12003), .B(n12002), .ZN(
        n12004) );
  OAI211_X1 U13910 ( .C1(n13175), .C2(n12246), .A(n12005), .B(n12004), .ZN(
        P3_U3161) );
  XNOR2_X1 U13911 ( .A(n12006), .B(n12012), .ZN(n12196) );
  INV_X1 U13912 ( .A(n12007), .ZN(n12008) );
  AOI211_X1 U13913 ( .C1(n12200), .C2(n12008), .A(n8098), .B(n12138), .ZN(
        n12198) );
  NOR2_X1 U13914 ( .A1(n12203), .A2(n14288), .ZN(n12011) );
  OAI22_X1 U13915 ( .A1(n14280), .A2(n12009), .B1(n12062), .B2(n14255), .ZN(
        n12010) );
  AOI211_X1 U13916 ( .C1(n12198), .C2(n14290), .A(n12011), .B(n12010), .ZN(
        n12020) );
  AOI22_X1 U13917 ( .A1(n14274), .A2(n13921), .B1(n12351), .B2(n14275), .ZN(
        n12018) );
  OAI21_X1 U13918 ( .B1(n12014), .B2(n12013), .A(n12012), .ZN(n12016) );
  NAND3_X1 U13919 ( .A1(n12016), .A2(n14271), .A3(n12015), .ZN(n12017) );
  OAI211_X1 U13920 ( .C1(n12196), .C2(n14279), .A(n12018), .B(n12017), .ZN(
        n12197) );
  NAND2_X1 U13921 ( .A1(n12197), .A2(n14280), .ZN(n12019) );
  OAI211_X1 U13922 ( .C1(n12196), .C2(n14293), .A(n12020), .B(n12019), .ZN(
        P2_U3253) );
  OAI22_X1 U13923 ( .A1(n13587), .A2(n12021), .B1(n13130), .B2(n15860), .ZN(
        n12024) );
  MUX2_X1 U13924 ( .A(P3_REG2_REG_5__SCAN_IN), .B(n12022), .S(n15867), .Z(
        n12023) );
  AOI211_X1 U13925 ( .C1(n13592), .C2(n12025), .A(n12024), .B(n12023), .ZN(
        n12026) );
  INV_X1 U13926 ( .A(n12026), .ZN(P3_U3228) );
  NAND2_X1 U13927 ( .A1(n12028), .A2(n12027), .ZN(n12029) );
  NAND2_X1 U13928 ( .A1(n12760), .A2(n14509), .ZN(n12032) );
  NAND2_X1 U13929 ( .A1(n14537), .A2(n14735), .ZN(n12031) );
  NAND2_X1 U13930 ( .A1(n12032), .A2(n12031), .ZN(n12151) );
  NAND2_X1 U13931 ( .A1(n12760), .A2(n14492), .ZN(n12034) );
  NAND2_X1 U13932 ( .A1(n14442), .A2(n14735), .ZN(n12033) );
  NAND2_X1 U13933 ( .A1(n12034), .A2(n12033), .ZN(n12035) );
  XNOR2_X1 U13934 ( .A(n12035), .B(n14586), .ZN(n12036) );
  NAND2_X1 U13935 ( .A1(n12037), .A2(n12036), .ZN(n12154) );
  OAI211_X1 U13936 ( .C1(n12037), .C2(n12036), .A(n12154), .B(n14690), .ZN(
        n12042) );
  NOR2_X1 U13937 ( .A1(n14701), .A2(n15937), .ZN(n12038) );
  AOI211_X1 U13938 ( .C1(n14671), .C2(n12040), .A(n12039), .B(n12038), .ZN(
        n12041) );
  OAI211_X1 U13939 ( .C1(n15943), .C2(n14698), .A(n12042), .B(n12041), .ZN(
        P1_U3231) );
  OAI22_X1 U13940 ( .A1(n13587), .A2(n12044), .B1(n12043), .B2(n15860), .ZN(
        n12047) );
  MUX2_X1 U13941 ( .A(n12045), .B(P3_REG2_REG_6__SCAN_IN), .S(n15869), .Z(
        n12046) );
  AOI211_X1 U13942 ( .C1(n13592), .C2(n12048), .A(n12047), .B(n12046), .ZN(
        n12049) );
  INV_X1 U13943 ( .A(n12049), .ZN(P3_U3227) );
  XNOR2_X1 U13944 ( .A(n12203), .B(n13764), .ZN(n12050) );
  OR2_X1 U13945 ( .A1(n12144), .A2(n14151), .ZN(n12051) );
  NAND2_X1 U13946 ( .A1(n12050), .A2(n12051), .ZN(n12100) );
  INV_X1 U13947 ( .A(n12050), .ZN(n12053) );
  INV_X1 U13948 ( .A(n12051), .ZN(n12052) );
  NAND2_X1 U13949 ( .A1(n12053), .A2(n12052), .ZN(n12054) );
  AND2_X1 U13950 ( .A1(n12100), .A2(n12054), .ZN(n12059) );
  OAI21_X1 U13951 ( .B1(n12059), .B2(n12058), .A(n12101), .ZN(n12060) );
  NAND2_X1 U13952 ( .A1(n12060), .A2(n13881), .ZN(n12065) );
  NAND2_X1 U13953 ( .A1(n13887), .A2(n12351), .ZN(n12061) );
  NAND2_X1 U13954 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n15532)
         );
  OAI211_X1 U13955 ( .C1(n13902), .C2(n12062), .A(n12061), .B(n15532), .ZN(
        n12063) );
  AOI21_X1 U13956 ( .B1(n13892), .B2(n13921), .A(n12063), .ZN(n12064) );
  OAI211_X1 U13957 ( .C1(n12203), .C2(n13889), .A(n12065), .B(n12064), .ZN(
        P2_U3196) );
  INV_X1 U13958 ( .A(n12066), .ZN(n12068) );
  OAI222_X1 U13959 ( .A1(n14422), .A2(n12067), .B1(n12358), .B2(n12068), .C1(
        n14076), .C2(P2_U3088), .ZN(P2_U3308) );
  OAI222_X1 U13960 ( .A1(n15435), .A2(n7694), .B1(n15437), .B2(n12068), .C1(
        P1_U3086), .C2(n14816), .ZN(P1_U3336) );
  XNOR2_X1 U13961 ( .A(n12069), .B(n12071), .ZN(n16009) );
  OAI21_X1 U13962 ( .B1(n7163), .B2(n12071), .A(n12070), .ZN(n16012) );
  NAND2_X1 U13963 ( .A1(n14561), .A2(n12072), .ZN(n12073) );
  NAND2_X1 U13964 ( .A1(n12073), .A2(n15878), .ZN(n12074) );
  OR2_X1 U13965 ( .A1(n7270), .A2(n12074), .ZN(n16005) );
  AND2_X1 U13966 ( .A1(n14702), .A2(n14731), .ZN(n12075) );
  AOI21_X1 U13967 ( .B1(n14729), .B2(n14704), .A(n12075), .ZN(n16004) );
  OAI22_X1 U13968 ( .A1(n15895), .A2(n16004), .B1(n14557), .B2(n15051), .ZN(
        n12077) );
  INV_X1 U13969 ( .A(n14561), .ZN(n16007) );
  NOR2_X1 U13970 ( .A1(n16007), .A2(n15942), .ZN(n12076) );
  AOI211_X1 U13971 ( .C1(n15895), .C2(P1_REG2_REG_14__SCAN_IN), .A(n12077), 
        .B(n12076), .ZN(n12078) );
  OAI21_X1 U13972 ( .B1(n15057), .B2(n16005), .A(n12078), .ZN(n12079) );
  AOI21_X1 U13973 ( .B1(n15000), .B2(n16012), .A(n12079), .ZN(n12080) );
  OAI21_X1 U13974 ( .B1(n16009), .B2(n15061), .A(n12080), .ZN(P1_U3279) );
  OAI21_X1 U13975 ( .B1(n12082), .B2(n12089), .A(n12081), .ZN(n12084) );
  XNOR2_X1 U13976 ( .A(n12084), .B(n15497), .ZN(n15493) );
  NOR2_X1 U13977 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n15493), .ZN(n15492) );
  INV_X1 U13978 ( .A(n15492), .ZN(n12083) );
  OAI21_X1 U13979 ( .B1(n12084), .B2(n15497), .A(n12083), .ZN(n12087) );
  MUX2_X1 U13980 ( .A(n14218), .B(P2_REG2_REG_19__SCAN_IN), .S(n12085), .Z(
        n12086) );
  XNOR2_X1 U13981 ( .A(n12087), .B(n12086), .ZN(n12099) );
  OAI21_X1 U13982 ( .B1(n11682), .B2(n12089), .A(n12088), .ZN(n12091) );
  XNOR2_X1 U13983 ( .A(n12091), .B(n12090), .ZN(n15487) );
  AND2_X1 U13984 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n15487), .ZN(n15489) );
  AOI21_X1 U13985 ( .B1(n12091), .B2(n15497), .A(n15489), .ZN(n12093) );
  XNOR2_X1 U13986 ( .A(n14076), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n12092) );
  XNOR2_X1 U13987 ( .A(n12093), .B(n12092), .ZN(n12097) );
  NAND2_X1 U13988 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13796)
         );
  NAND2_X1 U13989 ( .A1(n15501), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n12094) );
  OAI211_X1 U13990 ( .C1(n12095), .C2(n14076), .A(n13796), .B(n12094), .ZN(
        n12096) );
  AOI21_X1 U13991 ( .B1(n15527), .B2(n12097), .A(n12096), .ZN(n12098) );
  OAI21_X1 U13992 ( .B1(n12099), .B2(n15502), .A(n12098), .ZN(P2_U3233) );
  XNOR2_X1 U13993 ( .A(n15997), .B(n13805), .ZN(n12102) );
  OR2_X1 U13994 ( .A1(n12216), .A2(n14151), .ZN(n12103) );
  AND2_X1 U13995 ( .A1(n12102), .A2(n12103), .ZN(n12341) );
  INV_X1 U13996 ( .A(n12341), .ZN(n12106) );
  INV_X1 U13997 ( .A(n12102), .ZN(n12105) );
  INV_X1 U13998 ( .A(n12103), .ZN(n12104) );
  NAND2_X1 U13999 ( .A1(n12105), .A2(n12104), .ZN(n12342) );
  NAND2_X1 U14000 ( .A1(n12106), .A2(n12342), .ZN(n12107) );
  XNOR2_X1 U14001 ( .A(n12340), .B(n12107), .ZN(n12113) );
  NOR2_X1 U14002 ( .A1(n13859), .A2(n12334), .ZN(n12111) );
  NAND2_X1 U14003 ( .A1(n13892), .A2(n13920), .ZN(n12109) );
  NAND2_X1 U14004 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n12108)
         );
  OAI211_X1 U14005 ( .C1(n13902), .C2(n12135), .A(n12109), .B(n12108), .ZN(
        n12110) );
  AOI211_X1 U14006 ( .C1(n12141), .C2(n13905), .A(n12111), .B(n12110), .ZN(
        n12112) );
  OAI21_X1 U14007 ( .B1(n12113), .B2(n13907), .A(n12112), .ZN(P2_U3206) );
  MUX2_X1 U14008 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13728), .Z(n12183) );
  XNOR2_X1 U14009 ( .A(n12183), .B(n12182), .ZN(n12184) );
  NAND2_X1 U14010 ( .A1(n12114), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12124) );
  MUX2_X1 U14011 ( .A(n12124), .B(n12117), .S(n13728), .Z(n12115) );
  NAND2_X1 U14012 ( .A1(n12116), .A2(n12115), .ZN(n12185) );
  XOR2_X1 U14013 ( .A(n12184), .B(n12185), .Z(n12133) );
  INV_X1 U14014 ( .A(n12182), .ZN(n12131) );
  INV_X1 U14015 ( .A(n12117), .ZN(n12119) );
  AOI21_X1 U14016 ( .B1(n12122), .B2(n12121), .A(n12168), .ZN(n12129) );
  XNOR2_X1 U14017 ( .A(n12131), .B(n12173), .ZN(n12125) );
  NAND2_X1 U14018 ( .A1(P3_REG2_REG_13__SCAN_IN), .A2(n12125), .ZN(n12174) );
  OAI21_X1 U14019 ( .B1(n12125), .B2(P3_REG2_REG_13__SCAN_IN), .A(n12174), 
        .ZN(n12127) );
  AND2_X1 U14020 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n13173) );
  INV_X1 U14021 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15682) );
  NOR2_X1 U14022 ( .A1(n15787), .A2(n15682), .ZN(n12126) );
  AOI211_X1 U14023 ( .C1(n15815), .C2(n12127), .A(n13173), .B(n12126), .ZN(
        n12128) );
  OAI21_X1 U14024 ( .B1(n12129), .B2(n15800), .A(n12128), .ZN(n12130) );
  AOI21_X1 U14025 ( .B1(n12131), .B2(n15808), .A(n12130), .ZN(n12132) );
  OAI21_X1 U14026 ( .B1(n12133), .B2(n15763), .A(n12132), .ZN(P3_U3195) );
  XNOR2_X1 U14027 ( .A(n12134), .B(n12142), .ZN(n15995) );
  OAI22_X1 U14028 ( .A1(n14280), .A2(n12136), .B1(n12135), .B2(n14255), .ZN(
        n12140) );
  INV_X1 U14029 ( .A(n12137), .ZN(n12219) );
  OAI211_X1 U14030 ( .C1(n15997), .C2(n12138), .A(n12219), .B(n14151), .ZN(
        n15996) );
  NOR2_X1 U14031 ( .A1(n15996), .A2(n14261), .ZN(n12139) );
  AOI211_X1 U14032 ( .C1(n14258), .C2(n12141), .A(n12140), .B(n12139), .ZN(
        n12149) );
  XNOR2_X1 U14033 ( .A(n12143), .B(n12142), .ZN(n12146) );
  OAI22_X1 U14034 ( .A1(n12334), .A2(n14237), .B1(n12144), .B2(n14235), .ZN(
        n12145) );
  AOI21_X1 U14035 ( .B1(n12146), .B2(n14271), .A(n12145), .ZN(n12147) );
  OAI21_X1 U14036 ( .B1(n15995), .B2(n14279), .A(n12147), .ZN(n15998) );
  NAND2_X1 U14037 ( .A1(n15998), .A2(n14280), .ZN(n12148) );
  OAI211_X1 U14038 ( .C1(n15995), .C2(n14293), .A(n12149), .B(n12148), .ZN(
        P2_U3252) );
  INV_X1 U14039 ( .A(n12150), .ZN(n12152) );
  NAND2_X1 U14040 ( .A1(n12152), .A2(n12151), .ZN(n12153) );
  NAND2_X1 U14041 ( .A1(n12764), .A2(n14532), .ZN(n12156) );
  NAND2_X1 U14042 ( .A1(n14509), .A2(n14734), .ZN(n12155) );
  NAND2_X1 U14043 ( .A1(n12156), .A2(n12155), .ZN(n12157) );
  XNOR2_X1 U14044 ( .A(n12157), .B(n14522), .ZN(n12301) );
  NOR2_X1 U14045 ( .A1(n14588), .A2(n12158), .ZN(n12159) );
  AOI21_X1 U14046 ( .B1(n12764), .B2(n14442), .A(n12159), .ZN(n12298) );
  INV_X1 U14047 ( .A(n12298), .ZN(n12302) );
  XNOR2_X1 U14048 ( .A(n12301), .B(n12302), .ZN(n12160) );
  XNOR2_X1 U14049 ( .A(n12300), .B(n12160), .ZN(n12167) );
  NAND2_X1 U14050 ( .A1(n14671), .A2(n12161), .ZN(n12162) );
  OAI211_X1 U14051 ( .C1(n14701), .C2(n12164), .A(n12163), .B(n12162), .ZN(
        n12165) );
  AOI21_X1 U14052 ( .B1(n12764), .B2(n14709), .A(n12165), .ZN(n12166) );
  OAI21_X1 U14053 ( .B1(n12167), .B2(n14711), .A(n12166), .ZN(P1_U3217) );
  NAND2_X1 U14054 ( .A1(P3_REG1_REG_14__SCAN_IN), .A2(n13263), .ZN(n12170) );
  OAI21_X1 U14055 ( .B1(P3_REG1_REG_14__SCAN_IN), .B2(n13263), .A(n12170), 
        .ZN(n12171) );
  NOR2_X1 U14056 ( .A1(n12172), .A2(n12171), .ZN(n13254) );
  AOI21_X1 U14057 ( .B1(n12172), .B2(n12171), .A(n13254), .ZN(n12192) );
  INV_X1 U14058 ( .A(n13263), .ZN(n12190) );
  AOI22_X1 U14059 ( .A1(P3_REG2_REG_14__SCAN_IN), .A2(n13263), .B1(n12190), 
        .B2(n13589), .ZN(n12177) );
  NAND2_X1 U14060 ( .A1(n12182), .A2(n12173), .ZN(n12175) );
  OAI21_X1 U14061 ( .B1(n12177), .B2(n12176), .A(n13257), .ZN(n12178) );
  NAND2_X1 U14062 ( .A1(n15815), .A2(n12178), .ZN(n12181) );
  NOR2_X1 U14063 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12179), .ZN(n13062) );
  INV_X1 U14064 ( .A(n13062), .ZN(n12180) );
  OAI211_X1 U14065 ( .C1(n15691), .C2(n15787), .A(n12181), .B(n12180), .ZN(
        n12189) );
  MUX2_X1 U14066 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n13728), .Z(n13264) );
  XNOR2_X1 U14067 ( .A(n13264), .B(n13263), .ZN(n12187) );
  NOR2_X1 U14068 ( .A1(n12186), .A2(n12187), .ZN(n13262) );
  AOI211_X1 U14069 ( .C1(n12187), .C2(n12186), .A(n15763), .B(n13262), .ZN(
        n12188) );
  AOI211_X1 U14070 ( .C1(n15808), .C2(n12190), .A(n12189), .B(n12188), .ZN(
        n12191) );
  OAI21_X1 U14071 ( .B1(n12192), .B2(n15800), .A(n12191), .ZN(P3_U3196) );
  INV_X1 U14072 ( .A(n12193), .ZN(n12195) );
  OAI222_X1 U14073 ( .A1(n13730), .A2(n12195), .B1(n13723), .B2(n15174), .C1(
        P3_U3151), .C2(n12194), .ZN(P3_U3270) );
  INV_X1 U14074 ( .A(n12196), .ZN(n12199) );
  AOI211_X1 U14075 ( .C1(n12199), .C2(n16024), .A(n12198), .B(n12197), .ZN(
        n12206) );
  AOI22_X1 U14076 ( .A1(n12200), .A2(n14300), .B1(n16034), .B2(
        P2_REG1_REG_12__SCAN_IN), .ZN(n12201) );
  OAI21_X1 U14077 ( .B1(n12206), .B2(n16034), .A(n12201), .ZN(P2_U3511) );
  INV_X1 U14078 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n12202) );
  OAI22_X1 U14079 ( .A1(n12203), .A2(n14402), .B1(n14398), .B2(n12202), .ZN(
        n12204) );
  INV_X1 U14080 ( .A(n12204), .ZN(n12205) );
  OAI21_X1 U14081 ( .B1(n12206), .B2(n16001), .A(n12205), .ZN(P2_U3466) );
  OAI22_X1 U14082 ( .A1(n13587), .A2(n12208), .B1(n12207), .B2(n15860), .ZN(
        n12211) );
  MUX2_X1 U14083 ( .A(n12209), .B(P3_REG2_REG_7__SCAN_IN), .S(n15869), .Z(
        n12210) );
  AOI211_X1 U14084 ( .C1(n13592), .C2(n12212), .A(n12211), .B(n12210), .ZN(
        n12213) );
  INV_X1 U14085 ( .A(n12213), .ZN(P3_U3226) );
  XNOR2_X1 U14086 ( .A(n12214), .B(n12217), .ZN(n12215) );
  OAI222_X1 U14087 ( .A1(n14237), .A2(n12401), .B1(n14235), .B2(n12216), .C1(
        n12215), .C2(n14243), .ZN(n12274) );
  INV_X1 U14088 ( .A(n12274), .ZN(n12224) );
  XNOR2_X1 U14089 ( .A(n12218), .B(n12217), .ZN(n12276) );
  AOI211_X1 U14090 ( .C1(n12279), .C2(n12219), .A(n14282), .B(n12379), .ZN(
        n12275) );
  NAND2_X1 U14091 ( .A1(n12275), .A2(n14290), .ZN(n12221) );
  AOI22_X1 U14092 ( .A1(n14265), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n12346), 
        .B2(n14285), .ZN(n12220) );
  OAI211_X1 U14093 ( .C1(n12348), .C2(n14288), .A(n12221), .B(n12220), .ZN(
        n12222) );
  AOI21_X1 U14094 ( .B1(n14263), .B2(n12276), .A(n12222), .ZN(n12223) );
  OAI21_X1 U14095 ( .B1(n14265), .B2(n12224), .A(n12223), .ZN(P2_U3251) );
  XNOR2_X1 U14096 ( .A(n13053), .B(n12225), .ZN(n12424) );
  XNOR2_X1 U14097 ( .A(n12424), .B(n12285), .ZN(n12232) );
  INV_X1 U14098 ( .A(n12226), .ZN(n12227) );
  INV_X1 U14099 ( .A(n12426), .ZN(n12230) );
  AOI21_X1 U14100 ( .B1(n12232), .B2(n12231), .A(n12230), .ZN(n12237) );
  INV_X1 U14101 ( .A(n12257), .ZN(n12235) );
  INV_X1 U14102 ( .A(n13217), .ZN(n13225) );
  AOI22_X1 U14103 ( .A1(n13225), .A2(n13245), .B1(n13215), .B2(n13247), .ZN(
        n12233) );
  NAND2_X1 U14104 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(P3_U3151), .ZN(n15785) );
  OAI211_X1 U14105 ( .C1(n13234), .C2(n15929), .A(n12233), .B(n15785), .ZN(
        n12234) );
  AOI21_X1 U14106 ( .B1(n12235), .B2(n13230), .A(n12234), .ZN(n12236) );
  OAI21_X1 U14107 ( .B1(n12237), .B2(n13196), .A(n12236), .ZN(P3_U3171) );
  INV_X1 U14108 ( .A(n12238), .ZN(n12239) );
  AOI21_X1 U14109 ( .B1(n12664), .B2(n12240), .A(n12239), .ZN(n12241) );
  OAI222_X1 U14110 ( .A1(n13580), .A2(n12285), .B1(n13582), .B2(n12242), .C1(
        n13578), .C2(n12241), .ZN(n12265) );
  INV_X1 U14111 ( .A(n12265), .ZN(n12250) );
  OAI21_X1 U14112 ( .B1(n12244), .B2(n12664), .A(n12243), .ZN(n12266) );
  NOR2_X1 U14113 ( .A1(n15867), .A2(n12245), .ZN(n12248) );
  OAI22_X1 U14114 ( .A1(n13587), .A2(n12569), .B1(n12246), .B2(n15860), .ZN(
        n12247) );
  AOI211_X1 U14115 ( .C1(n12266), .C2(n13592), .A(n12248), .B(n12247), .ZN(
        n12249) );
  OAI21_X1 U14116 ( .B1(n12250), .B2(n15869), .A(n12249), .ZN(P3_U3225) );
  INV_X1 U14117 ( .A(n12251), .ZN(n12574) );
  OR2_X1 U14118 ( .A1(n12574), .A2(n12575), .ZN(n12665) );
  XNOR2_X1 U14119 ( .A(n12252), .B(n12665), .ZN(n15930) );
  XNOR2_X1 U14120 ( .A(n12253), .B(n12665), .ZN(n12255) );
  OAI22_X1 U14121 ( .A1(n12568), .A2(n13582), .B1(n12423), .B2(n13580), .ZN(
        n12254) );
  AOI21_X1 U14122 ( .B1(n12255), .B2(n15851), .A(n12254), .ZN(n12256) );
  OAI21_X1 U14123 ( .B1(n15855), .B2(n15930), .A(n12256), .ZN(n15932) );
  NAND2_X1 U14124 ( .A1(n15932), .A2(n15867), .ZN(n12260) );
  OAI22_X1 U14125 ( .A1(n13587), .A2(n15929), .B1(n12257), .B2(n15860), .ZN(
        n12258) );
  AOI21_X1 U14126 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n15869), .A(n12258), .ZN(
        n12259) );
  OAI211_X1 U14127 ( .C1(n15930), .C2(n12292), .A(n12260), .B(n12259), .ZN(
        P3_U3224) );
  INV_X1 U14128 ( .A(n12261), .ZN(n12264) );
  OAI222_X1 U14129 ( .A1(n13730), .A2(n12264), .B1(n13723), .B2(n12263), .C1(
        P3_U3151), .C2(n12262), .ZN(P3_U3269) );
  AOI21_X1 U14130 ( .B1(n13658), .B2(n12266), .A(n12265), .ZN(n12271) );
  OAI22_X1 U14131 ( .A1(n13707), .A2(n12569), .B1(n16042), .B2(n8319), .ZN(
        n12267) );
  INV_X1 U14132 ( .A(n12267), .ZN(n12268) );
  OAI21_X1 U14133 ( .B1(n12271), .B2(n16048), .A(n12268), .ZN(P3_U3414) );
  AOI22_X1 U14134 ( .A1(n16045), .A2(n12269), .B1(n8727), .B2(
        P3_REG1_REG_8__SCAN_IN), .ZN(n12270) );
  OAI21_X1 U14135 ( .B1(n12271), .B2(n8727), .A(n12270), .ZN(P3_U3467) );
  INV_X1 U14136 ( .A(n12272), .ZN(n12282) );
  OAI222_X1 U14137 ( .A1(n15435), .A2(n12273), .B1(n15437), .B2(n12282), .C1(
        n15827), .C2(P1_U3086), .ZN(P1_U3335) );
  AOI211_X1 U14138 ( .C1(n16033), .C2(n12276), .A(n12275), .B(n12274), .ZN(
        n12281) );
  OAI22_X1 U14139 ( .A1(n12348), .A2(n14402), .B1(n14371), .B2(n9121), .ZN(
        n12277) );
  INV_X1 U14140 ( .A(n12277), .ZN(n12278) );
  OAI21_X1 U14141 ( .B1(n12281), .B2(n16001), .A(n12278), .ZN(P2_U3472) );
  AOI22_X1 U14142 ( .A1(n12279), .A2(n14300), .B1(n16034), .B2(
        P2_REG1_REG_14__SCAN_IN), .ZN(n12280) );
  OAI21_X1 U14143 ( .B1(n12281), .B2(n16034), .A(n12280), .ZN(P2_U3513) );
  OAI222_X1 U14144 ( .A1(n14422), .A2(n7692), .B1(P2_U3088), .B2(n9563), .C1(
        n14416), .C2(n12282), .ZN(P2_U3307) );
  XNOR2_X1 U14145 ( .A(n12283), .B(n7634), .ZN(n15958) );
  XNOR2_X1 U14146 ( .A(n12284), .B(n7634), .ZN(n12287) );
  OAI22_X1 U14147 ( .A1(n13048), .A2(n13580), .B1(n12285), .B2(n13582), .ZN(
        n12286) );
  AOI21_X1 U14148 ( .B1(n12287), .B2(n15851), .A(n12286), .ZN(n12288) );
  OAI21_X1 U14149 ( .B1(n15855), .B2(n15958), .A(n12288), .ZN(n15960) );
  NAND2_X1 U14150 ( .A1(n15960), .A2(n15867), .ZN(n12291) );
  OAI22_X1 U14151 ( .A1(n13587), .A2(n15957), .B1(n12418), .B2(n15860), .ZN(
        n12289) );
  AOI21_X1 U14152 ( .B1(n15869), .B2(P3_REG2_REG_10__SCAN_IN), .A(n12289), 
        .ZN(n12290) );
  OAI211_X1 U14153 ( .C1(n15958), .C2(n12292), .A(n12291), .B(n12290), .ZN(
        P3_U3223) );
  NAND2_X1 U14154 ( .A1(n12773), .A2(n14532), .ZN(n12294) );
  NAND2_X1 U14155 ( .A1(n14442), .A2(n14733), .ZN(n12293) );
  NAND2_X1 U14156 ( .A1(n12294), .A2(n12293), .ZN(n12295) );
  XNOR2_X1 U14157 ( .A(n12295), .B(n14522), .ZN(n12316) );
  NOR2_X1 U14158 ( .A1(n14588), .A2(n12296), .ZN(n12297) );
  AOI21_X1 U14159 ( .B1(n12773), .B2(n14509), .A(n12297), .ZN(n12315) );
  XNOR2_X1 U14160 ( .A(n12316), .B(n12315), .ZN(n12307) );
  NAND2_X1 U14161 ( .A1(n12301), .A2(n12298), .ZN(n12299) );
  INV_X1 U14162 ( .A(n12301), .ZN(n12303) );
  NAND2_X1 U14163 ( .A1(n12303), .A2(n12302), .ZN(n12304) );
  INV_X1 U14164 ( .A(n12324), .ZN(n12305) );
  AOI21_X1 U14165 ( .B1(n12307), .B2(n12306), .A(n12305), .ZN(n12314) );
  AOI21_X1 U14166 ( .B1(n14671), .B2(n12309), .A(n12308), .ZN(n12310) );
  OAI21_X1 U14167 ( .B1(n14701), .B2(n12311), .A(n12310), .ZN(n12312) );
  AOI21_X1 U14168 ( .B1(n12773), .B2(n14709), .A(n12312), .ZN(n12313) );
  OAI21_X1 U14169 ( .B1(n12314), .B2(n14711), .A(n12313), .ZN(P1_U3236) );
  NAND2_X1 U14170 ( .A1(n12316), .A2(n12315), .ZN(n12322) );
  AND2_X1 U14171 ( .A1(n12324), .A2(n12322), .ZN(n12326) );
  NAND2_X1 U14172 ( .A1(n12777), .A2(n14532), .ZN(n12318) );
  NAND2_X1 U14173 ( .A1(n14442), .A2(n14732), .ZN(n12317) );
  NAND2_X1 U14174 ( .A1(n12318), .A2(n12317), .ZN(n12319) );
  XNOR2_X1 U14175 ( .A(n12319), .B(n14586), .ZN(n12387) );
  NOR2_X1 U14176 ( .A1(n14588), .A2(n12320), .ZN(n12321) );
  AOI21_X1 U14177 ( .B1(n12777), .B2(n14509), .A(n12321), .ZN(n12385) );
  XNOR2_X1 U14178 ( .A(n12387), .B(n12385), .ZN(n12325) );
  AND2_X1 U14179 ( .A1(n12325), .A2(n12322), .ZN(n12323) );
  OAI211_X1 U14180 ( .C1(n12326), .C2(n12325), .A(n14690), .B(n12389), .ZN(
        n12332) );
  OAI21_X1 U14181 ( .B1(n14706), .B2(n12328), .A(n12327), .ZN(n12329) );
  AOI21_X1 U14182 ( .B1(n14695), .B2(n12330), .A(n12329), .ZN(n12331) );
  OAI211_X1 U14183 ( .C1(n12333), .C2(n14698), .A(n12332), .B(n12331), .ZN(
        P1_U3224) );
  XNOR2_X1 U14184 ( .A(n12348), .B(n13764), .ZN(n12335) );
  OR2_X1 U14185 ( .A1(n12334), .A2(n14151), .ZN(n12336) );
  NAND2_X1 U14186 ( .A1(n12335), .A2(n12336), .ZN(n12407) );
  INV_X1 U14187 ( .A(n12335), .ZN(n12338) );
  INV_X1 U14188 ( .A(n12336), .ZN(n12337) );
  NAND2_X1 U14189 ( .A1(n12338), .A2(n12337), .ZN(n12339) );
  NAND2_X1 U14190 ( .A1(n12407), .A2(n12339), .ZN(n12345) );
  AOI21_X1 U14191 ( .B1(n12345), .B2(n12344), .A(n7990), .ZN(n12353) );
  NAND2_X1 U14192 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14030)
         );
  NAND2_X1 U14193 ( .A1(n13856), .A2(n12346), .ZN(n12347) );
  OAI211_X1 U14194 ( .C1(n13859), .C2(n12401), .A(n14030), .B(n12347), .ZN(
        n12350) );
  NOR2_X1 U14195 ( .A1(n12348), .A2(n13889), .ZN(n12349) );
  AOI211_X1 U14196 ( .C1(n13892), .C2(n12351), .A(n12350), .B(n12349), .ZN(
        n12352) );
  OAI21_X1 U14197 ( .B1(n12353), .B2(n13907), .A(n12352), .ZN(P2_U3187) );
  INV_X1 U14198 ( .A(n12354), .ZN(n12357) );
  OAI222_X1 U14199 ( .A1(n15435), .A2(n12355), .B1(n15437), .B2(n12357), .C1(
        P1_U3086), .C2(n12704), .ZN(P1_U3334) );
  OAI222_X1 U14200 ( .A1(n14422), .A2(n12359), .B1(n12358), .B2(n12357), .C1(
        n12356), .C2(P2_U3088), .ZN(P2_U3306) );
  XNOR2_X1 U14201 ( .A(n12360), .B(n12968), .ZN(n12361) );
  OAI222_X1 U14202 ( .A1(n13582), .A2(n12423), .B1(n13580), .B2(n13193), .C1(
        n12361), .C2(n13578), .ZN(n12465) );
  INV_X1 U14203 ( .A(n12465), .ZN(n12368) );
  OAI22_X1 U14204 ( .A1(n13587), .A2(n12471), .B1(n13189), .B2(n15860), .ZN(
        n12366) );
  INV_X1 U14205 ( .A(n12362), .ZN(n12364) );
  AND2_X1 U14206 ( .A1(n12363), .A2(n12968), .ZN(n12464) );
  NOR3_X1 U14207 ( .A1(n12364), .A2(n12464), .A3(n13532), .ZN(n12365) );
  AOI211_X1 U14208 ( .C1(n15869), .C2(P3_REG2_REG_11__SCAN_IN), .A(n12366), 
        .B(n12365), .ZN(n12367) );
  OAI21_X1 U14209 ( .B1(n12368), .B2(n15869), .A(n12367), .ZN(P3_U3222) );
  INV_X1 U14210 ( .A(n12369), .ZN(n12370) );
  AOI21_X1 U14211 ( .B1(n12372), .B2(n12371), .A(n12370), .ZN(n16018) );
  AOI22_X1 U14212 ( .A1(n14249), .A2(n14275), .B1(n14274), .B2(n13919), .ZN(
        n12376) );
  XNOR2_X1 U14213 ( .A(n12373), .B(n12372), .ZN(n12374) );
  NAND2_X1 U14214 ( .A1(n12374), .A2(n14271), .ZN(n12375) );
  OAI211_X1 U14215 ( .C1(n16018), .C2(n14279), .A(n12376), .B(n12375), .ZN(
        n16021) );
  NAND2_X1 U14216 ( .A1(n16021), .A2(n14280), .ZN(n12384) );
  OAI22_X1 U14217 ( .A1(n14280), .A2(n12377), .B1(n12414), .B2(n14255), .ZN(
        n12381) );
  INV_X1 U14218 ( .A(n12378), .ZN(n14283) );
  OAI211_X1 U14219 ( .C1(n16020), .C2(n12379), .A(n14283), .B(n14151), .ZN(
        n16019) );
  NOR2_X1 U14220 ( .A1(n16019), .A2(n14261), .ZN(n12380) );
  AOI211_X1 U14221 ( .C1(n14258), .C2(n12382), .A(n12381), .B(n12380), .ZN(
        n12383) );
  OAI211_X1 U14222 ( .C1(n16018), .C2(n14293), .A(n12384), .B(n12383), .ZN(
        P2_U3250) );
  INV_X1 U14223 ( .A(n12385), .ZN(n12386) );
  NAND2_X1 U14224 ( .A1(n12387), .A2(n12386), .ZN(n12388) );
  NAND2_X1 U14225 ( .A1(n15983), .A2(n14532), .ZN(n12391) );
  NAND2_X1 U14226 ( .A1(n14442), .A2(n14731), .ZN(n12390) );
  NAND2_X1 U14227 ( .A1(n12391), .A2(n12390), .ZN(n12392) );
  XNOR2_X1 U14228 ( .A(n12392), .B(n14586), .ZN(n14440) );
  NOR2_X1 U14229 ( .A1(n14588), .A2(n12393), .ZN(n12394) );
  AOI21_X1 U14230 ( .B1(n15983), .B2(n14442), .A(n12394), .ZN(n14438) );
  XNOR2_X1 U14231 ( .A(n14440), .B(n14438), .ZN(n14436) );
  XNOR2_X1 U14232 ( .A(n14437), .B(n14436), .ZN(n12400) );
  NAND2_X1 U14233 ( .A1(n14695), .A2(n12395), .ZN(n12397) );
  OAI211_X1 U14234 ( .C1(n15980), .C2(n14706), .A(n12397), .B(n12396), .ZN(
        n12398) );
  AOI21_X1 U14235 ( .B1(n15983), .B2(n14709), .A(n12398), .ZN(n12399) );
  OAI21_X1 U14236 ( .B1(n12400), .B2(n14711), .A(n12399), .ZN(P1_U3234) );
  XNOR2_X1 U14237 ( .A(n16020), .B(n13805), .ZN(n12402) );
  OR2_X1 U14238 ( .A1(n12401), .A2(n14151), .ZN(n12403) );
  NAND2_X1 U14239 ( .A1(n12402), .A2(n12403), .ZN(n12447) );
  INV_X1 U14240 ( .A(n12402), .ZN(n12405) );
  INV_X1 U14241 ( .A(n12403), .ZN(n12404) );
  NAND2_X1 U14242 ( .A1(n12405), .A2(n12404), .ZN(n12406) );
  AND2_X1 U14243 ( .A1(n12447), .A2(n12406), .ZN(n12410) );
  OAI21_X1 U14244 ( .B1(n12410), .B2(n12409), .A(n12448), .ZN(n12411) );
  NAND2_X1 U14245 ( .A1(n12411), .A2(n13881), .ZN(n12417) );
  NAND2_X1 U14246 ( .A1(n13887), .A2(n14249), .ZN(n12413) );
  OAI211_X1 U14247 ( .C1(n13902), .C2(n12414), .A(n12413), .B(n12412), .ZN(
        n12415) );
  AOI21_X1 U14248 ( .B1(n13892), .B2(n13919), .A(n12415), .ZN(n12416) );
  OAI211_X1 U14249 ( .C1(n16020), .C2(n13889), .A(n12417), .B(n12416), .ZN(
        P2_U3213) );
  INV_X1 U14250 ( .A(n12418), .ZN(n12431) );
  NAND2_X1 U14251 ( .A1(n13215), .A2(n13246), .ZN(n12421) );
  NAND2_X1 U14252 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n15803)
         );
  INV_X1 U14253 ( .A(n15803), .ZN(n12419) );
  AOI21_X1 U14254 ( .B1(n13190), .B2(n12422), .A(n12419), .ZN(n12420) );
  OAI211_X1 U14255 ( .C1(n13048), .C2(n13217), .A(n12421), .B(n12420), .ZN(
        n12430) );
  XNOR2_X1 U14256 ( .A(n13053), .B(n12422), .ZN(n12965) );
  XNOR2_X1 U14257 ( .A(n12965), .B(n12423), .ZN(n12428) );
  NAND2_X1 U14258 ( .A1(n12424), .A2(n12285), .ZN(n12425) );
  AOI211_X1 U14259 ( .C1(n12428), .C2(n12427), .A(n13196), .B(n12966), .ZN(
        n12429) );
  AOI211_X1 U14260 ( .C1(n12431), .C2(n13230), .A(n12430), .B(n12429), .ZN(
        n12432) );
  INV_X1 U14261 ( .A(n12432), .ZN(P3_U3157) );
  INV_X1 U14262 ( .A(n12580), .ZN(n12668) );
  XNOR2_X1 U14263 ( .A(n12433), .B(n12668), .ZN(n12434) );
  OAI222_X1 U14264 ( .A1(n13582), .A2(n13048), .B1(n13580), .B2(n13581), .C1(
        n13578), .C2(n12434), .ZN(n15974) );
  INV_X1 U14265 ( .A(n15974), .ZN(n12440) );
  AOI21_X1 U14266 ( .B1(n12362), .B2(n12583), .A(n12668), .ZN(n12435) );
  NOR2_X1 U14267 ( .A1(n7273), .A2(n12435), .ZN(n15973) );
  INV_X1 U14268 ( .A(n15973), .ZN(n15976) );
  INV_X1 U14269 ( .A(n12436), .ZN(n13102) );
  AOI22_X1 U14270 ( .A1(n15869), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n13541), 
        .B2(n13102), .ZN(n12437) );
  OAI21_X1 U14271 ( .B1(n15971), .B2(n13587), .A(n12437), .ZN(n12438) );
  AOI21_X1 U14272 ( .B1(n15976), .B2(n13592), .A(n12438), .ZN(n12439) );
  OAI21_X1 U14273 ( .B1(n12440), .B2(n15869), .A(n12439), .ZN(P3_U3221) );
  XNOR2_X1 U14274 ( .A(n14403), .B(n13764), .ZN(n12442) );
  OR2_X1 U14275 ( .A1(n12441), .A2(n14151), .ZN(n12443) );
  NAND2_X1 U14276 ( .A1(n12442), .A2(n12443), .ZN(n13731) );
  INV_X1 U14277 ( .A(n12442), .ZN(n12445) );
  INV_X1 U14278 ( .A(n12443), .ZN(n12444) );
  NAND2_X1 U14279 ( .A1(n12445), .A2(n12444), .ZN(n12446) );
  AND2_X1 U14280 ( .A1(n13731), .A2(n12446), .ZN(n12450) );
  OAI21_X1 U14281 ( .B1(n12450), .B2(n12449), .A(n13732), .ZN(n12451) );
  NAND2_X1 U14282 ( .A1(n12451), .A2(n13881), .ZN(n12456) );
  NAND2_X1 U14283 ( .A1(n13856), .A2(n14286), .ZN(n12452) );
  OAI211_X1 U14284 ( .C1(n13859), .C2(n14236), .A(n12453), .B(n12452), .ZN(
        n12454) );
  AOI21_X1 U14285 ( .B1(n13892), .B2(n14273), .A(n12454), .ZN(n12455) );
  OAI211_X1 U14286 ( .C1(n14403), .C2(n13889), .A(n12456), .B(n12455), .ZN(
        P2_U3198) );
  INV_X1 U14287 ( .A(n12457), .ZN(n12460) );
  OAI222_X1 U14288 ( .A1(n15435), .A2(n7394), .B1(n15437), .B2(n12460), .C1(
        P1_U3086), .C2(n12458), .ZN(P1_U3331) );
  OAI222_X1 U14289 ( .A1(n14422), .A2(n7395), .B1(n14416), .B2(n12460), .C1(
        P2_U3088), .C2(n12459), .ZN(P2_U3303) );
  INV_X1 U14290 ( .A(n12461), .ZN(n12462) );
  OAI222_X1 U14291 ( .A1(n14422), .A2(n12463), .B1(n14416), .B2(n12462), .C1(
        n9530), .C2(P2_U3088), .ZN(P2_U3305) );
  INV_X1 U14292 ( .A(n13658), .ZN(n13639) );
  NOR2_X1 U14293 ( .A1(n12464), .A2(n13639), .ZN(n12466) );
  AOI21_X1 U14294 ( .B1(n12466), .B2(n12362), .A(n12465), .ZN(n12468) );
  MUX2_X1 U14295 ( .A(n11799), .B(n12468), .S(n16039), .Z(n12467) );
  OAI21_X1 U14296 ( .B1(n13656), .B2(n12471), .A(n12467), .ZN(P3_U3470) );
  INV_X1 U14297 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n12469) );
  MUX2_X1 U14298 ( .A(n12469), .B(n12468), .S(n16042), .Z(n12470) );
  OAI21_X1 U14299 ( .B1(n13707), .B2(n12471), .A(n12470), .ZN(P3_U3423) );
  INV_X1 U14300 ( .A(n13056), .ZN(n12975) );
  XNOR2_X1 U14301 ( .A(n12472), .B(n12975), .ZN(n12473) );
  AOI222_X1 U14302 ( .A1(n15851), .A2(n12473), .B1(n13564), .B2(n15846), .C1(
        n13243), .C2(n15848), .ZN(n13661) );
  XNOR2_X1 U14303 ( .A(n12474), .B(n13056), .ZN(n13659) );
  NOR2_X1 U14304 ( .A1(n12589), .A2(n13587), .ZN(n12477) );
  OAI22_X1 U14305 ( .A1(n15867), .A2(n12475), .B1(n13176), .B2(n15860), .ZN(
        n12476) );
  AOI211_X1 U14306 ( .C1(n13659), .C2(n13592), .A(n12477), .B(n12476), .ZN(
        n12478) );
  OAI21_X1 U14307 ( .B1(n13661), .B2(n15869), .A(n12478), .ZN(P3_U3220) );
  INV_X1 U14308 ( .A(n12479), .ZN(n12483) );
  OAI222_X1 U14309 ( .A1(n14422), .A2(n12481), .B1(n14416), .B2(n12483), .C1(
        P2_U3088), .C2(n12480), .ZN(P2_U3302) );
  OAI222_X1 U14310 ( .A1(n15435), .A2(n7369), .B1(n15437), .B2(n12483), .C1(
        P1_U3086), .C2(n12482), .ZN(P1_U3330) );
  INV_X1 U14311 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12492) );
  OAI222_X1 U14312 ( .A1(n14416), .A2(n15427), .B1(P2_U3088), .B2(n12484), 
        .C1(n12492), .C2(n14422), .ZN(P2_U3297) );
  INV_X1 U14313 ( .A(n12485), .ZN(n12486) );
  OAI222_X1 U14314 ( .A1(n13723), .A2(n15281), .B1(P3_U3151), .B2(n8663), .C1(
        n13730), .C2(n12486), .ZN(P3_U3267) );
  INV_X1 U14315 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n15426) );
  AOI22_X1 U14316 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n12492), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n15426), .ZN(n12507) );
  AOI22_X1 U14317 ( .A1(n12958), .A2(P1_DATAO_REG_29__SCAN_IN), .B1(n12489), 
        .B2(n12488), .ZN(n12490) );
  INV_X1 U14318 ( .A(n12490), .ZN(n12508) );
  NAND2_X1 U14319 ( .A1(n12507), .A2(n12508), .ZN(n12491) );
  OAI21_X1 U14320 ( .B1(n12492), .B2(P2_DATAO_REG_30__SCAN_IN), .A(n12491), 
        .ZN(n12495) );
  INV_X1 U14321 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n12862) );
  AOI22_X1 U14322 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(
        P1_DATAO_REG_31__SCAN_IN), .B1(n12493), .B2(n12862), .ZN(n12494) );
  XNOR2_X1 U14323 ( .A(n12495), .B(n12494), .ZN(n13718) );
  NAND2_X1 U14324 ( .A1(n13718), .A2(n12496), .ZN(n12498) );
  INV_X1 U14325 ( .A(SI_31_), .ZN(n13713) );
  OR2_X1 U14326 ( .A1(n7158), .A2(n13713), .ZN(n12497) );
  INV_X1 U14327 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12502) );
  NAND2_X1 U14328 ( .A1(n8567), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12501) );
  INV_X1 U14329 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n12499) );
  OR2_X1 U14330 ( .A1(n8240), .A2(n12499), .ZN(n12500) );
  OAI211_X1 U14331 ( .C1(n12503), .C2(n12502), .A(n12501), .B(n12500), .ZN(
        n12504) );
  INV_X1 U14332 ( .A(n12504), .ZN(n12505) );
  NAND2_X1 U14333 ( .A1(n12506), .A2(n12505), .ZN(n13235) );
  INV_X1 U14334 ( .A(n13235), .ZN(n13374) );
  NAND2_X1 U14335 ( .A1(n16050), .A2(n13374), .ZN(n12514) );
  INV_X1 U14336 ( .A(n12643), .ZN(n13236) );
  XNOR2_X1 U14337 ( .A(n12508), .B(n12507), .ZN(n13720) );
  OR2_X1 U14338 ( .A1(n12509), .A2(n13720), .ZN(n12512) );
  INV_X1 U14339 ( .A(SI_30_), .ZN(n15284) );
  OR2_X1 U14340 ( .A1(n7158), .A2(n15284), .ZN(n12511) );
  INV_X1 U14341 ( .A(n16041), .ZN(n13379) );
  NAND2_X1 U14342 ( .A1(n13236), .A2(n13379), .ZN(n12513) );
  NAND2_X1 U14343 ( .A1(n12514), .A2(n12513), .ZN(n12516) );
  NAND2_X1 U14344 ( .A1(n12516), .A2(n16050), .ZN(n12648) );
  NAND4_X1 U14345 ( .A1(n12515), .A2(n12685), .A3(n13361), .A4(n12648), .ZN(
        n12655) );
  INV_X1 U14346 ( .A(n12516), .ZN(n12681) );
  INV_X1 U14347 ( .A(n13413), .ZN(n12517) );
  AND3_X1 U14348 ( .A1(n13398), .A2(n13427), .A3(n12517), .ZN(n12633) );
  INV_X1 U14349 ( .A(n12633), .ZN(n12679) );
  NAND2_X1 U14350 ( .A1(n12518), .A2(n13396), .ZN(n12523) );
  INV_X1 U14351 ( .A(n12519), .ZN(n12520) );
  NAND2_X1 U14352 ( .A1(n12521), .A2(n12520), .ZN(n12522) );
  NAND3_X1 U14353 ( .A1(n12524), .A2(n12523), .A3(n12522), .ZN(n12526) );
  AND2_X1 U14354 ( .A1(n12526), .A2(n12525), .ZN(n12529) );
  INV_X1 U14355 ( .A(n12529), .ZN(n12527) );
  OAI21_X1 U14356 ( .B1(n12679), .B2(n12528), .A(n12527), .ZN(n12531) );
  INV_X1 U14357 ( .A(n12533), .ZN(n12534) );
  NOR2_X1 U14358 ( .A1(n12535), .A2(n12534), .ZN(n12537) );
  OAI211_X1 U14359 ( .C1(n12537), .C2(n12697), .A(n12536), .B(n8239), .ZN(
        n12541) );
  INV_X1 U14360 ( .A(n12537), .ZN(n12539) );
  AOI21_X1 U14361 ( .B1(n12539), .B2(n12538), .A(n12635), .ZN(n12540) );
  AOI21_X1 U14362 ( .B1(n12541), .B2(n15842), .A(n12540), .ZN(n12550) );
  NAND2_X1 U14363 ( .A1(n12547), .A2(n12542), .ZN(n12545) );
  NAND2_X1 U14364 ( .A1(n12546), .A2(n12543), .ZN(n12544) );
  MUX2_X1 U14365 ( .A(n12545), .B(n12544), .S(n12635), .Z(n12549) );
  MUX2_X1 U14366 ( .A(n12547), .B(n12546), .S(n12641), .Z(n12548) );
  OAI21_X1 U14367 ( .B1(n12550), .B2(n12549), .A(n12548), .ZN(n12551) );
  NAND2_X1 U14368 ( .A1(n12551), .A2(n12663), .ZN(n12555) );
  MUX2_X1 U14369 ( .A(n12553), .B(n12552), .S(n12641), .Z(n12554) );
  NAND3_X1 U14370 ( .A1(n12555), .A2(n12662), .A3(n12554), .ZN(n12559) );
  MUX2_X1 U14371 ( .A(n12557), .B(n12556), .S(n12635), .Z(n12558) );
  NAND3_X1 U14372 ( .A1(n12559), .A2(n12661), .A3(n12558), .ZN(n12564) );
  MUX2_X1 U14373 ( .A(n12561), .B(n12560), .S(n12641), .Z(n12563) );
  MUX2_X1 U14374 ( .A(n12566), .B(n12565), .S(n12641), .Z(n12567) );
  NAND2_X1 U14375 ( .A1(n12567), .A2(n12664), .ZN(n12573) );
  NAND2_X1 U14376 ( .A1(n12568), .A2(n12635), .ZN(n12571) );
  NAND2_X1 U14377 ( .A1(n13247), .A2(n12641), .ZN(n12570) );
  MUX2_X1 U14378 ( .A(n12571), .B(n12570), .S(n12569), .Z(n12572) );
  INV_X1 U14379 ( .A(n12665), .ZN(n12578) );
  MUX2_X1 U14380 ( .A(n12575), .B(n12574), .S(n12641), .Z(n12577) );
  NAND2_X1 U14381 ( .A1(n12585), .A2(n12579), .ZN(n12582) );
  AOI21_X1 U14382 ( .B1(n12582), .B2(n12581), .A(n12580), .ZN(n12587) );
  XNOR2_X1 U14383 ( .A(n13054), .B(n12641), .ZN(n12586) );
  NAND3_X1 U14384 ( .A1(n12972), .A2(n12641), .A3(n12583), .ZN(n12584) );
  OAI22_X1 U14385 ( .A1(n12587), .A2(n12586), .B1(n12585), .B2(n12584), .ZN(
        n12592) );
  INV_X1 U14386 ( .A(n12589), .ZN(n13657) );
  NOR2_X1 U14387 ( .A1(n13657), .A2(n13581), .ZN(n12590) );
  MUX2_X1 U14388 ( .A(n7639), .B(n12590), .S(n12635), .Z(n12591) );
  AOI211_X1 U14389 ( .C1(n12592), .C2(n13056), .A(n12591), .B(n13586), .ZN(
        n12593) );
  NOR2_X1 U14390 ( .A1(n12593), .A2(n13567), .ZN(n12597) );
  MUX2_X1 U14391 ( .A(n12595), .B(n12594), .S(n12635), .Z(n12596) );
  INV_X1 U14392 ( .A(n12598), .ZN(n12599) );
  INV_X1 U14393 ( .A(n12601), .ZN(n12602) );
  NAND2_X1 U14394 ( .A1(n13536), .A2(n12641), .ZN(n12604) );
  NAND2_X1 U14395 ( .A1(n12611), .A2(n12604), .ZN(n12606) );
  OR2_X1 U14396 ( .A1(n13636), .A2(n12635), .ZN(n12605) );
  AND2_X1 U14397 ( .A1(n12606), .A2(n12605), .ZN(n12613) );
  INV_X1 U14398 ( .A(n13538), .ZN(n12607) );
  INV_X1 U14399 ( .A(n12611), .ZN(n12610) );
  OAI211_X1 U14400 ( .C1(n12610), .C2(n12609), .A(n12620), .B(n12608), .ZN(
        n12615) );
  OAI211_X1 U14401 ( .C1(n12613), .C2(n12612), .A(n12621), .B(n12611), .ZN(
        n12614) );
  MUX2_X1 U14402 ( .A(n12615), .B(n12614), .S(n12641), .Z(n12616) );
  OAI21_X1 U14403 ( .B1(n12617), .B2(n12616), .A(n13489), .ZN(n12618) );
  INV_X1 U14404 ( .A(n12618), .ZN(n12622) );
  AOI21_X1 U14405 ( .B1(n12622), .B2(n12620), .A(n7465), .ZN(n12624) );
  AOI22_X1 U14406 ( .A1(n12622), .A2(n12621), .B1(n13505), .B2(n12999), .ZN(
        n12623) );
  MUX2_X1 U14407 ( .A(n12624), .B(n12623), .S(n12635), .Z(n12626) );
  NAND2_X1 U14408 ( .A1(n13003), .A2(n13005), .ZN(n13475) );
  MUX2_X1 U14409 ( .A(n13003), .B(n13005), .S(n12635), .Z(n12625) );
  OAI211_X1 U14410 ( .C1(n12626), .C2(n13475), .A(n13460), .B(n12625), .ZN(
        n12630) );
  NAND2_X1 U14411 ( .A1(n13186), .A2(n13449), .ZN(n12627) );
  MUX2_X1 U14412 ( .A(n12628), .B(n12627), .S(n12641), .Z(n12629) );
  NAND3_X1 U14413 ( .A1(n13073), .A2(n13462), .A3(n12635), .ZN(n12632) );
  NAND3_X1 U14414 ( .A1(n13679), .A2(n12641), .A3(n13239), .ZN(n12631) );
  NAND2_X1 U14415 ( .A1(n12638), .A2(n12637), .ZN(n12642) );
  INV_X1 U14416 ( .A(n12687), .ZN(n12639) );
  NAND2_X1 U14417 ( .A1(n13376), .A2(n13235), .ZN(n12645) );
  NAND2_X1 U14418 ( .A1(n12643), .A2(n16041), .ZN(n12644) );
  NAND2_X1 U14419 ( .A1(n12646), .A2(n12682), .ZN(n12647) );
  OAI211_X1 U14420 ( .C1(n12681), .C2(n13235), .A(n12647), .B(n12648), .ZN(
        n12653) );
  INV_X1 U14421 ( .A(n12682), .ZN(n12689) );
  NAND2_X1 U14422 ( .A1(n13374), .A2(n16041), .ZN(n12684) );
  NAND3_X1 U14423 ( .A1(n12687), .A2(n13361), .A3(n12684), .ZN(n12651) );
  INV_X1 U14424 ( .A(n12648), .ZN(n12649) );
  XNOR2_X1 U14425 ( .A(n12649), .B(n12686), .ZN(n12650) );
  OAI211_X1 U14426 ( .C1(n12689), .C2(n12651), .A(n12650), .B(n12685), .ZN(
        n12652) );
  NAND4_X1 U14427 ( .A1(n12660), .A2(n12659), .A3(n12658), .A4(n12657), .ZN(
        n12667) );
  NAND4_X1 U14428 ( .A1(n12663), .A2(n8239), .A3(n12662), .A4(n12661), .ZN(
        n12666) );
  NOR4_X1 U14429 ( .A1(n12667), .A2(n12666), .A3(n8629), .A4(n12665), .ZN(
        n12670) );
  INV_X1 U14430 ( .A(n12968), .ZN(n12669) );
  NAND4_X1 U14431 ( .A1(n12670), .A2(n12669), .A3(n7634), .A4(n12668), .ZN(
        n12671) );
  NOR4_X1 U14432 ( .A1(n13567), .A2(n13586), .A3(n12975), .A4(n12671), .ZN(
        n12672) );
  NAND4_X1 U14433 ( .A1(n13522), .A2(n13558), .A3(n13538), .A4(n12672), .ZN(
        n12673) );
  NOR4_X1 U14434 ( .A1(n13475), .A2(n12674), .A3(n13509), .A4(n12673), .ZN(
        n12676) );
  NAND4_X1 U14435 ( .A1(n13435), .A2(n12676), .A3(n13460), .A4(n12675), .ZN(
        n12677) );
  NOR3_X1 U14436 ( .A1(n12679), .A2(n12678), .A3(n12677), .ZN(n12680) );
  NAND4_X1 U14437 ( .A1(n12682), .A2(n12636), .A3(n12681), .A4(n12680), .ZN(
        n12683) );
  XNOR2_X1 U14438 ( .A(n12683), .B(n12686), .ZN(n12693) );
  NAND4_X1 U14439 ( .A1(n12687), .A2(n12686), .A3(n12685), .A4(n12684), .ZN(
        n12688) );
  NOR2_X1 U14440 ( .A1(n12689), .A2(n12688), .ZN(n12691) );
  AOI22_X1 U14441 ( .A1(n12693), .A2(n12692), .B1(n12691), .B2(n12690), .ZN(
        n12694) );
  NOR3_X1 U14442 ( .A1(n12696), .A2(n12695), .A3(n8663), .ZN(n12699) );
  OAI21_X1 U14443 ( .B1(n12700), .B2(n12697), .A(P3_B_REG_SCAN_IN), .ZN(n12698) );
  OAI22_X1 U14444 ( .A1(n12701), .A2(n12700), .B1(n12699), .B2(n12698), .ZN(
        P3_U3296) );
  NAND2_X1 U14445 ( .A1(n12705), .A2(n12704), .ZN(n12858) );
  NAND2_X1 U14446 ( .A1(n12707), .A2(n12706), .ZN(n12709) );
  NAND2_X1 U14447 ( .A1(n12709), .A2(n12708), .ZN(n12712) );
  NAND4_X1 U14448 ( .A1(n12715), .A2(n12873), .A3(n12714), .A4(n10010), .ZN(
        n12727) );
  AND2_X1 U14449 ( .A1(n12716), .A2(n12728), .ZN(n12720) );
  NAND2_X1 U14450 ( .A1(n15898), .A2(n14741), .ZN(n12717) );
  NAND2_X1 U14451 ( .A1(n12720), .A2(n12719), .ZN(n12726) );
  NOR2_X1 U14452 ( .A1(n12728), .A2(n12721), .ZN(n12724) );
  OAI21_X1 U14453 ( .B1(n12873), .B2(n14741), .A(n12723), .ZN(n12722) );
  OAI21_X1 U14454 ( .B1(n12724), .B2(n12723), .A(n12722), .ZN(n12725) );
  NAND3_X1 U14455 ( .A1(n12727), .A2(n12726), .A3(n12725), .ZN(n12732) );
  MUX2_X1 U14456 ( .A(n12729), .B(n14740), .S(n12873), .Z(n12733) );
  NAND2_X1 U14457 ( .A1(n12732), .A2(n12733), .ZN(n12731) );
  MUX2_X1 U14458 ( .A(n12729), .B(n14740), .S(n12728), .Z(n12730) );
  NAND2_X1 U14459 ( .A1(n12731), .A2(n12730), .ZN(n12737) );
  INV_X1 U14460 ( .A(n12732), .ZN(n12735) );
  INV_X1 U14461 ( .A(n12733), .ZN(n12734) );
  NAND2_X1 U14462 ( .A1(n12735), .A2(n12734), .ZN(n12736) );
  MUX2_X1 U14463 ( .A(n12738), .B(n14739), .S(n12728), .Z(n12740) );
  MUX2_X1 U14464 ( .A(n14739), .B(n12738), .S(n12728), .Z(n12739) );
  MUX2_X1 U14465 ( .A(n14738), .B(n12741), .S(n12728), .Z(n12745) );
  MUX2_X1 U14466 ( .A(n12743), .B(n12742), .S(n12873), .Z(n12744) );
  AOI21_X1 U14467 ( .B1(n12746), .B2(n12745), .A(n12744), .ZN(n12748) );
  NOR2_X1 U14468 ( .A1(n12746), .A2(n12745), .ZN(n12747) );
  MUX2_X1 U14469 ( .A(n12749), .B(n14737), .S(n12728), .Z(n12751) );
  MUX2_X1 U14470 ( .A(n12749), .B(n14737), .S(n12873), .Z(n12750) );
  MUX2_X1 U14471 ( .A(n14736), .B(n12753), .S(n12871), .Z(n12756) );
  NAND2_X1 U14472 ( .A1(n12757), .A2(n12756), .ZN(n12755) );
  MUX2_X1 U14473 ( .A(n12753), .B(n14736), .S(n12871), .Z(n12754) );
  NAND2_X1 U14474 ( .A1(n12755), .A2(n12754), .ZN(n12759) );
  MUX2_X1 U14475 ( .A(n14735), .B(n12760), .S(n12873), .Z(n12762) );
  MUX2_X1 U14476 ( .A(n14735), .B(n12760), .S(n12871), .Z(n12761) );
  INV_X1 U14477 ( .A(n12762), .ZN(n12763) );
  MUX2_X1 U14478 ( .A(n14734), .B(n12764), .S(n12871), .Z(n12768) );
  NAND2_X1 U14479 ( .A1(n12767), .A2(n12768), .ZN(n12766) );
  MUX2_X1 U14480 ( .A(n14734), .B(n12764), .S(n12873), .Z(n12765) );
  NAND2_X1 U14481 ( .A1(n12766), .A2(n12765), .ZN(n12772) );
  INV_X1 U14482 ( .A(n12767), .ZN(n12770) );
  INV_X1 U14483 ( .A(n12768), .ZN(n12769) );
  NAND2_X1 U14484 ( .A1(n12770), .A2(n12769), .ZN(n12771) );
  MUX2_X1 U14485 ( .A(n14733), .B(n12773), .S(n12873), .Z(n12775) );
  MUX2_X1 U14486 ( .A(n14733), .B(n12773), .S(n12871), .Z(n12774) );
  INV_X1 U14487 ( .A(n12775), .ZN(n12776) );
  MUX2_X1 U14488 ( .A(n14732), .B(n12777), .S(n12871), .Z(n12781) );
  NAND2_X1 U14489 ( .A1(n12780), .A2(n12781), .ZN(n12779) );
  MUX2_X1 U14490 ( .A(n14732), .B(n12777), .S(n12873), .Z(n12778) );
  NAND2_X1 U14491 ( .A1(n12779), .A2(n12778), .ZN(n12785) );
  INV_X1 U14492 ( .A(n12780), .ZN(n12783) );
  INV_X1 U14493 ( .A(n12781), .ZN(n12782) );
  NAND2_X1 U14494 ( .A1(n12783), .A2(n12782), .ZN(n12784) );
  MUX2_X1 U14495 ( .A(n14731), .B(n15983), .S(n12873), .Z(n12787) );
  MUX2_X1 U14496 ( .A(n14731), .B(n15983), .S(n12871), .Z(n12786) );
  MUX2_X1 U14497 ( .A(n14730), .B(n14561), .S(n12871), .Z(n12791) );
  NAND2_X1 U14498 ( .A1(n12790), .A2(n12791), .ZN(n12789) );
  MUX2_X1 U14499 ( .A(n14730), .B(n14561), .S(n12873), .Z(n12788) );
  NAND2_X1 U14500 ( .A1(n12789), .A2(n12788), .ZN(n12795) );
  INV_X1 U14501 ( .A(n12790), .ZN(n12793) );
  INV_X1 U14502 ( .A(n12791), .ZN(n12792) );
  NAND2_X1 U14503 ( .A1(n12793), .A2(n12792), .ZN(n12794) );
  MUX2_X1 U14504 ( .A(n14729), .B(n15413), .S(n12873), .Z(n12797) );
  MUX2_X1 U14505 ( .A(n14729), .B(n15413), .S(n12871), .Z(n12796) );
  MUX2_X1 U14506 ( .A(n14728), .B(n15150), .S(n12871), .Z(n12799) );
  MUX2_X1 U14507 ( .A(n14728), .B(n15150), .S(n12873), .Z(n12798) );
  INV_X1 U14508 ( .A(n12799), .ZN(n12800) );
  MUX2_X1 U14509 ( .A(n14726), .B(n15142), .S(n12873), .Z(n12802) );
  MUX2_X1 U14510 ( .A(n14726), .B(n15142), .S(n12871), .Z(n12801) );
  INV_X1 U14511 ( .A(n12802), .ZN(n12803) );
  MUX2_X1 U14512 ( .A(n14725), .B(n15407), .S(n12871), .Z(n12807) );
  NAND2_X1 U14513 ( .A1(n12806), .A2(n12807), .ZN(n12805) );
  MUX2_X1 U14514 ( .A(n15407), .B(n14725), .S(n12871), .Z(n12804) );
  NAND2_X1 U14515 ( .A1(n12805), .A2(n12804), .ZN(n12811) );
  INV_X1 U14516 ( .A(n12806), .ZN(n12809) );
  INV_X1 U14517 ( .A(n12807), .ZN(n12808) );
  NAND2_X1 U14518 ( .A1(n12809), .A2(n12808), .ZN(n12810) );
  MUX2_X1 U14519 ( .A(n14724), .B(n14980), .S(n12873), .Z(n12813) );
  MUX2_X1 U14520 ( .A(n14724), .B(n14980), .S(n12871), .Z(n12812) );
  MUX2_X1 U14521 ( .A(n14723), .B(n14967), .S(n12728), .Z(n12815) );
  MUX2_X1 U14522 ( .A(n14967), .B(n14723), .S(n12728), .Z(n12814) );
  MUX2_X1 U14523 ( .A(n14722), .B(n15115), .S(n12873), .Z(n12816) );
  MUX2_X1 U14524 ( .A(n14722), .B(n15115), .S(n12728), .Z(n12818) );
  NOR2_X1 U14525 ( .A1(n14721), .A2(n12871), .ZN(n12821) );
  NAND2_X1 U14526 ( .A1(n14721), .A2(n12728), .ZN(n12819) );
  NAND2_X1 U14527 ( .A1(n15108), .A2(n12819), .ZN(n12820) );
  OAI21_X1 U14528 ( .B1(n15108), .B2(n12821), .A(n12820), .ZN(n12822) );
  MUX2_X1 U14529 ( .A(n14720), .B(n15100), .S(n12873), .Z(n12826) );
  NAND2_X1 U14530 ( .A1(n12825), .A2(n12826), .ZN(n12824) );
  MUX2_X1 U14531 ( .A(n14720), .B(n15100), .S(n12728), .Z(n12823) );
  INV_X1 U14532 ( .A(n12825), .ZN(n12828) );
  INV_X1 U14533 ( .A(n12826), .ZN(n12827) );
  NAND2_X1 U14534 ( .A1(n12828), .A2(n12827), .ZN(n12829) );
  MUX2_X1 U14535 ( .A(n14719), .B(n14905), .S(n12728), .Z(n12831) );
  MUX2_X1 U14536 ( .A(n14719), .B(n14905), .S(n12873), .Z(n12830) );
  MUX2_X1 U14537 ( .A(n14718), .B(n14897), .S(n12873), .Z(n12835) );
  NAND2_X1 U14538 ( .A1(n12834), .A2(n12835), .ZN(n12833) );
  MUX2_X1 U14539 ( .A(n14718), .B(n14897), .S(n12728), .Z(n12832) );
  NAND2_X1 U14540 ( .A1(n12833), .A2(n12832), .ZN(n12839) );
  INV_X1 U14541 ( .A(n12834), .ZN(n12837) );
  INV_X1 U14542 ( .A(n12835), .ZN(n12836) );
  NAND2_X1 U14543 ( .A1(n12837), .A2(n12836), .ZN(n12838) );
  MUX2_X1 U14544 ( .A(n14717), .B(n15079), .S(n12728), .Z(n12841) );
  MUX2_X1 U14545 ( .A(n14717), .B(n15079), .S(n12873), .Z(n12840) );
  MUX2_X1 U14546 ( .A(n14716), .B(n14870), .S(n12873), .Z(n12845) );
  NAND2_X1 U14547 ( .A1(n12844), .A2(n12845), .ZN(n12843) );
  MUX2_X1 U14548 ( .A(n14716), .B(n14870), .S(n12871), .Z(n12842) );
  NAND2_X1 U14549 ( .A1(n12843), .A2(n12842), .ZN(n12849) );
  INV_X1 U14550 ( .A(n12844), .ZN(n12847) );
  INV_X1 U14551 ( .A(n12845), .ZN(n12846) );
  NAND2_X1 U14552 ( .A1(n12847), .A2(n12846), .ZN(n12848) );
  MUX2_X1 U14553 ( .A(n14715), .B(n14599), .S(n12728), .Z(n12850) );
  MUX2_X1 U14554 ( .A(n14599), .B(n14715), .S(n12871), .Z(n12851) );
  OAI21_X1 U14555 ( .B1(n12866), .B2(n15827), .A(n14713), .ZN(n12852) );
  INV_X1 U14556 ( .A(n12852), .ZN(n12856) );
  OR2_X1 U14557 ( .A1(n12863), .A2(n15426), .ZN(n12854) );
  MUX2_X1 U14558 ( .A(n12856), .B(n15382), .S(n12871), .Z(n12919) );
  INV_X1 U14559 ( .A(n12919), .ZN(n12922) );
  INV_X1 U14560 ( .A(n12866), .ZN(n14821) );
  AOI21_X1 U14561 ( .B1(n14821), .B2(n12858), .A(n12857), .ZN(n12859) );
  MUX2_X1 U14562 ( .A(n15382), .B(n12859), .S(n12728), .Z(n12939) );
  NAND2_X1 U14563 ( .A1(n12861), .A2(n12860), .ZN(n12865) );
  OR2_X1 U14564 ( .A1(n12863), .A2(n12862), .ZN(n12864) );
  XNOR2_X1 U14565 ( .A(n15064), .B(n12866), .ZN(n12923) );
  NAND2_X1 U14566 ( .A1(n10051), .A2(n15827), .ZN(n12867) );
  NAND2_X1 U14567 ( .A1(n12868), .A2(n12867), .ZN(n12870) );
  NAND2_X1 U14568 ( .A1(n12870), .A2(n12869), .ZN(n12913) );
  NOR2_X1 U14569 ( .A1(n12913), .A2(n15440), .ZN(n12921) );
  OAI211_X1 U14570 ( .C1(n12922), .C2(n12939), .A(n12923), .B(n12921), .ZN(
        n12934) );
  MUX2_X1 U14571 ( .A(n12872), .B(n14842), .S(n12871), .Z(n12933) );
  MUX2_X1 U14572 ( .A(n14714), .B(n10099), .S(n12873), .Z(n12932) );
  NOR2_X1 U14573 ( .A1(n12933), .A2(n12932), .ZN(n12946) );
  NOR2_X1 U14574 ( .A1(n12934), .A2(n12946), .ZN(n12949) );
  INV_X1 U14575 ( .A(n12923), .ZN(n12914) );
  NAND4_X1 U14576 ( .A1(n12876), .A2(n15873), .A3(n12875), .A4(n12874), .ZN(
        n12877) );
  NOR2_X1 U14577 ( .A1(n12878), .A2(n12877), .ZN(n12881) );
  NAND4_X1 U14578 ( .A1(n12882), .A2(n12881), .A3(n12880), .A4(n12879), .ZN(
        n12883) );
  NOR2_X1 U14579 ( .A1(n12884), .A2(n12883), .ZN(n12887) );
  NAND4_X1 U14580 ( .A1(n12888), .A2(n12887), .A3(n12886), .A4(n12885), .ZN(
        n12889) );
  OR4_X1 U14581 ( .A1(n12892), .A2(n12891), .A3(n12890), .A4(n12889), .ZN(
        n12893) );
  NOR2_X1 U14582 ( .A1(n15042), .A2(n12893), .ZN(n12894) );
  NAND4_X1 U14583 ( .A1(n14998), .A2(n12894), .A3(n15013), .A4(n15030), .ZN(
        n12895) );
  NOR4_X1 U14584 ( .A1(n14943), .A2(n12896), .A3(n14978), .A4(n12895), .ZN(
        n12898) );
  NAND4_X1 U14585 ( .A1(n12899), .A2(n14934), .A3(n12898), .A4(n12897), .ZN(
        n12900) );
  NOR4_X1 U14586 ( .A1(n12902), .A2(n12901), .A3(n14926), .A4(n12900), .ZN(
        n12905) );
  XNOR2_X1 U14587 ( .A(n15382), .B(n14713), .ZN(n12903) );
  NAND4_X1 U14588 ( .A1(n12905), .A2(n12904), .A3(n14861), .A4(n12903), .ZN(
        n12906) );
  NOR2_X1 U14589 ( .A1(n12914), .A2(n12906), .ZN(n12907) );
  XOR2_X1 U14590 ( .A(n10000), .B(n12907), .Z(n12911) );
  OR2_X1 U14591 ( .A1(n15064), .A2(n14821), .ZN(n12909) );
  NAND2_X1 U14592 ( .A1(n15064), .A2(n14821), .ZN(n12908) );
  XNOR2_X1 U14593 ( .A(n12938), .B(n12913), .ZN(n12910) );
  MUX2_X1 U14594 ( .A(n12911), .B(n12910), .S(n12912), .Z(n12942) );
  NAND2_X1 U14595 ( .A1(n12913), .A2(n12912), .ZN(n12917) );
  INV_X1 U14596 ( .A(n15440), .ZN(n12941) );
  NOR2_X1 U14597 ( .A1(n12917), .A2(n15440), .ZN(n12918) );
  NAND2_X1 U14598 ( .A1(n12919), .A2(n12918), .ZN(n12944) );
  NOR2_X1 U14599 ( .A1(n12944), .A2(n12939), .ZN(n12920) );
  NAND2_X1 U14600 ( .A1(n12938), .A2(n12920), .ZN(n12931) );
  NAND4_X1 U14601 ( .A1(n12923), .A2(n12922), .A3(n12939), .A4(n12921), .ZN(
        n12930) );
  NAND3_X1 U14602 ( .A1(n14702), .A2(n12925), .A3(n12924), .ZN(n12928) );
  AOI21_X1 U14603 ( .B1(n12941), .B2(n10051), .A(n12926), .ZN(n12927) );
  OAI21_X1 U14604 ( .B1(n12928), .B2(n15415), .A(n12927), .ZN(n12929) );
  AND3_X1 U14605 ( .A1(n12931), .A2(n12930), .A3(n12929), .ZN(n12935) );
  NAND2_X1 U14606 ( .A1(n12933), .A2(n12932), .ZN(n12951) );
  INV_X1 U14607 ( .A(n12938), .ZN(n12945) );
  INV_X1 U14608 ( .A(n12939), .ZN(n12940) );
  NAND3_X1 U14609 ( .A1(n12942), .A2(n12941), .A3(n12940), .ZN(n12943) );
  OAI21_X1 U14610 ( .B1(n12945), .B2(n12944), .A(n12943), .ZN(n12952) );
  NAND2_X1 U14611 ( .A1(n8099), .A2(n12947), .ZN(n12948) );
  AOI21_X1 U14612 ( .B1(n12950), .B2(n12949), .A(n12948), .ZN(n12955) );
  NAND3_X1 U14613 ( .A1(n12953), .A2(n12952), .A3(n12951), .ZN(n12954) );
  NAND2_X1 U14614 ( .A1(n12955), .A2(n12954), .ZN(P1_U3242) );
  INV_X1 U14615 ( .A(n12956), .ZN(n14406) );
  OAI222_X1 U14616 ( .A1(n15435), .A2(n12958), .B1(n15437), .B2(n14406), .C1(
        n12957), .C2(P1_U3086), .ZN(P1_U3326) );
  NAND3_X1 U14617 ( .A1(n12960), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n12964) );
  NAND2_X1 U14618 ( .A1(n12861), .A2(n14419), .ZN(n12963) );
  NAND2_X1 U14619 ( .A1(n12961), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n12962) );
  OAI211_X1 U14620 ( .C1(n12959), .C2(n12964), .A(n12963), .B(n12962), .ZN(
        P2_U3296) );
  INV_X1 U14621 ( .A(n12965), .ZN(n12967) );
  XNOR2_X1 U14622 ( .A(n12968), .B(n13050), .ZN(n13047) );
  NAND2_X1 U14623 ( .A1(n12975), .A2(n13049), .ZN(n12971) );
  NAND3_X1 U14624 ( .A1(n13056), .A2(n13053), .A3(n12972), .ZN(n12969) );
  OAI21_X1 U14625 ( .B1(n12971), .B2(n13053), .A(n12969), .ZN(n12970) );
  NOR3_X1 U14626 ( .A1(n12971), .A2(n13053), .A3(n13244), .ZN(n12974) );
  INV_X1 U14627 ( .A(n12972), .ZN(n13052) );
  NOR4_X1 U14628 ( .A1(n12975), .A2(n13050), .A3(n13052), .A4(n13244), .ZN(
        n12973) );
  INV_X1 U14629 ( .A(n13047), .ZN(n13197) );
  OAI21_X1 U14630 ( .B1(n12974), .B2(n12973), .A(n13197), .ZN(n12981) );
  NOR2_X1 U14631 ( .A1(n13050), .A2(n13054), .ZN(n12976) );
  AOI211_X1 U14632 ( .C1(n13581), .C2(n13050), .A(n12976), .B(n12975), .ZN(
        n12979) );
  NOR2_X1 U14633 ( .A1(n13055), .A2(n13053), .ZN(n12977) );
  AOI211_X1 U14634 ( .C1(n13581), .C2(n13053), .A(n12977), .B(n13056), .ZN(
        n12978) );
  XNOR2_X1 U14635 ( .A(n13706), .B(n13050), .ZN(n12982) );
  NAND2_X1 U14636 ( .A1(n12982), .A2(n13228), .ZN(n12985) );
  INV_X1 U14637 ( .A(n12982), .ZN(n12983) );
  NAND2_X1 U14638 ( .A1(n12983), .A2(n13564), .ZN(n12984) );
  AND2_X1 U14639 ( .A1(n12985), .A2(n12984), .ZN(n13058) );
  NAND2_X1 U14640 ( .A1(n13059), .A2(n12985), .ZN(n13221) );
  XNOR2_X1 U14641 ( .A(n13651), .B(n13053), .ZN(n12987) );
  XNOR2_X1 U14642 ( .A(n12987), .B(n13579), .ZN(n13222) );
  XNOR2_X1 U14643 ( .A(n13644), .B(n13053), .ZN(n12989) );
  XNOR2_X1 U14644 ( .A(n12989), .B(n13535), .ZN(n13121) );
  NOR2_X1 U14645 ( .A1(n12989), .A2(n13535), .ZN(n12990) );
  XNOR2_X1 U14646 ( .A(n13700), .B(n13053), .ZN(n13136) );
  NAND2_X1 U14647 ( .A1(n13136), .A2(n13552), .ZN(n12992) );
  INV_X1 U14648 ( .A(n13136), .ZN(n12991) );
  XNOR2_X1 U14649 ( .A(n13636), .B(n13053), .ZN(n12993) );
  XNOR2_X1 U14650 ( .A(n12993), .B(n13241), .ZN(n13204) );
  INV_X1 U14651 ( .A(n12993), .ZN(n12994) );
  NAND2_X1 U14652 ( .A1(n12994), .A2(n13241), .ZN(n12995) );
  XNOR2_X1 U14653 ( .A(n13514), .B(n13053), .ZN(n12996) );
  XNOR2_X1 U14654 ( .A(n12996), .B(n13492), .ZN(n13077) );
  NAND2_X1 U14655 ( .A1(n13078), .A2(n13077), .ZN(n13076) );
  INV_X1 U14656 ( .A(n12996), .ZN(n12997) );
  NAND2_X1 U14657 ( .A1(n12997), .A2(n13492), .ZN(n12998) );
  XNOR2_X1 U14658 ( .A(n12999), .B(n13053), .ZN(n13000) );
  XNOR2_X1 U14659 ( .A(n13000), .B(n13473), .ZN(n13164) );
  INV_X1 U14660 ( .A(n13000), .ZN(n13001) );
  NAND2_X1 U14661 ( .A1(n13001), .A2(n13473), .ZN(n13002) );
  MUX2_X1 U14662 ( .A(n7271), .B(n7462), .S(n13053), .Z(n13085) );
  INV_X1 U14663 ( .A(n13085), .ZN(n13004) );
  MUX2_X1 U14664 ( .A(n13006), .B(n13005), .S(n13053), .Z(n13083) );
  NAND2_X1 U14665 ( .A1(n13007), .A2(n13083), .ZN(n13009) );
  XNOR2_X1 U14666 ( .A(n13186), .B(n13053), .ZN(n13008) );
  XNOR2_X1 U14667 ( .A(n13073), .B(n13053), .ZN(n13010) );
  NAND2_X1 U14668 ( .A1(n13012), .A2(n13144), .ZN(n13068) );
  XNOR2_X1 U14669 ( .A(n13675), .B(n13050), .ZN(n13013) );
  NAND2_X1 U14670 ( .A1(n13013), .A2(n13450), .ZN(n13108) );
  INV_X1 U14671 ( .A(n13013), .ZN(n13014) );
  NAND2_X1 U14672 ( .A1(n13014), .A2(n13423), .ZN(n13015) );
  NAND2_X1 U14673 ( .A1(n13106), .A2(n13108), .ZN(n13019) );
  XNOR2_X1 U14674 ( .A(n13105), .B(n13053), .ZN(n13016) );
  NAND2_X1 U14675 ( .A1(n13016), .A2(n13437), .ZN(n13020) );
  INV_X1 U14676 ( .A(n13016), .ZN(n13017) );
  NAND2_X1 U14677 ( .A1(n13017), .A2(n13238), .ZN(n13018) );
  XNOR2_X1 U14678 ( .A(n7564), .B(n13053), .ZN(n13021) );
  NOR2_X1 U14679 ( .A1(n13021), .A2(n7563), .ZN(n13022) );
  AOI21_X1 U14680 ( .B1(n13021), .B2(n7563), .A(n13022), .ZN(n13213) );
  XNOR2_X1 U14681 ( .A(n8660), .B(n13050), .ZN(n13023) );
  INV_X1 U14682 ( .A(n13412), .ZN(n13237) );
  NOR2_X1 U14683 ( .A1(n13023), .A2(n13237), .ZN(n13024) );
  AOI21_X1 U14684 ( .B1(n13023), .B2(n13237), .A(n13024), .ZN(n13040) );
  INV_X1 U14685 ( .A(n13024), .ZN(n13025) );
  NAND2_X1 U14686 ( .A1(n13039), .A2(n13025), .ZN(n13027) );
  XNOR2_X1 U14687 ( .A(n7543), .B(n13053), .ZN(n13026) );
  XNOR2_X1 U14688 ( .A(n13027), .B(n13026), .ZN(n13028) );
  NAND2_X1 U14689 ( .A1(n13028), .A2(n13223), .ZN(n13035) );
  AOI22_X1 U14690 ( .A1(n13237), .A2(n13215), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13030) );
  NAND2_X1 U14691 ( .A1(n13388), .A2(n13230), .ZN(n13029) );
  OAI211_X1 U14692 ( .C1(n13031), .C2(n13217), .A(n13030), .B(n13029), .ZN(
        n13032) );
  AOI21_X1 U14693 ( .B1(n13033), .B2(n13190), .A(n13032), .ZN(n13034) );
  NAND2_X1 U14694 ( .A1(n13035), .A2(n13034), .ZN(P3_U3160) );
  NAND2_X1 U14695 ( .A1(n13036), .A2(P3_U3151), .ZN(n13037) );
  OAI21_X1 U14696 ( .B1(P3_U3151), .B2(n8690), .A(n13037), .ZN(P3_U3271) );
  OAI21_X1 U14697 ( .B1(n13040), .B2(n13038), .A(n13039), .ZN(n13041) );
  NAND2_X1 U14698 ( .A1(n13041), .A2(n13223), .ZN(n13045) );
  INV_X1 U14699 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n15272) );
  OAI22_X1 U14700 ( .A1(n13396), .A2(n13227), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15272), .ZN(n13043) );
  NOR2_X1 U14701 ( .A1(n13397), .A2(n13217), .ZN(n13042) );
  AOI211_X1 U14702 ( .C1(n13405), .C2(n13230), .A(n13043), .B(n13042), .ZN(
        n13044) );
  OAI211_X1 U14703 ( .C1(n13664), .C2(n13234), .A(n13045), .B(n13044), .ZN(
        P3_U3154) );
  INV_X1 U14704 ( .A(n13198), .ZN(n13046) );
  NAND2_X1 U14705 ( .A1(n13046), .A2(n13047), .ZN(n13194) );
  OAI21_X1 U14706 ( .B1(n13048), .B2(n13047), .A(n13194), .ZN(n13097) );
  INV_X1 U14707 ( .A(n13049), .ZN(n13051) );
  MUX2_X1 U14708 ( .A(n13052), .B(n13051), .S(n13050), .Z(n13095) );
  MUX2_X1 U14709 ( .A(n13055), .B(n13054), .S(n13053), .Z(n13093) );
  OAI21_X1 U14710 ( .B1(n13097), .B2(n13095), .A(n13093), .ZN(n13170) );
  XNOR2_X1 U14711 ( .A(n13056), .B(n13053), .ZN(n13171) );
  NOR2_X1 U14712 ( .A1(n13171), .A2(n13242), .ZN(n13057) );
  AOI211_X1 U14713 ( .C1(n13170), .C2(n13171), .A(n13058), .B(n13057), .ZN(
        n13061) );
  INV_X1 U14714 ( .A(n13059), .ZN(n13060) );
  OAI21_X1 U14715 ( .B1(n13061), .B2(n13060), .A(n13223), .ZN(n13067) );
  INV_X1 U14716 ( .A(n13588), .ZN(n13065) );
  AOI21_X1 U14717 ( .B1(n13215), .B2(n13242), .A(n13062), .ZN(n13063) );
  OAI21_X1 U14718 ( .B1(n13579), .B2(n13217), .A(n13063), .ZN(n13064) );
  AOI21_X1 U14719 ( .B1(n13065), .B2(n13230), .A(n13064), .ZN(n13066) );
  OAI211_X1 U14720 ( .C1(n13234), .C2(n13706), .A(n13067), .B(n13066), .ZN(
        P3_U3155) );
  AOI21_X1 U14721 ( .B1(n13239), .B2(n13069), .A(n7187), .ZN(n13075) );
  AOI22_X1 U14722 ( .A1(n13215), .A2(n13474), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13071) );
  NAND2_X1 U14723 ( .A1(n13230), .A2(n13453), .ZN(n13070) );
  OAI211_X1 U14724 ( .C1(n13450), .C2(n13217), .A(n13071), .B(n13070), .ZN(
        n13072) );
  AOI21_X1 U14725 ( .B1(n13073), .B2(n13190), .A(n13072), .ZN(n13074) );
  OAI21_X1 U14726 ( .B1(n13075), .B2(n13196), .A(n13074), .ZN(P3_U3156) );
  INV_X1 U14727 ( .A(n13514), .ZN(n13695) );
  OAI211_X1 U14728 ( .C1(n13078), .C2(n13077), .A(n13076), .B(n13223), .ZN(
        n13082) );
  INV_X1 U14729 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n15232) );
  NOR2_X1 U14730 ( .A1(n15232), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13364) );
  AOI21_X1 U14731 ( .B1(n13225), .B2(n13473), .A(n13364), .ZN(n13079) );
  OAI21_X1 U14732 ( .B1(n13536), .B2(n13227), .A(n13079), .ZN(n13080) );
  AOI21_X1 U14733 ( .B1(n13506), .B2(n13230), .A(n13080), .ZN(n13081) );
  OAI211_X1 U14734 ( .C1(n13695), .C2(n13234), .A(n13082), .B(n13081), .ZN(
        P3_U3159) );
  INV_X1 U14735 ( .A(n13083), .ZN(n13084) );
  NOR2_X1 U14736 ( .A1(n13085), .A2(n13084), .ZN(n13086) );
  XNOR2_X1 U14737 ( .A(n13087), .B(n13086), .ZN(n13092) );
  AOI22_X1 U14738 ( .A1(n13215), .A2(n13473), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13089) );
  NAND2_X1 U14739 ( .A1(n13230), .A2(n13481), .ZN(n13088) );
  OAI211_X1 U14740 ( .C1(n13449), .C2(n13217), .A(n13089), .B(n13088), .ZN(
        n13090) );
  AOI21_X1 U14741 ( .B1(n13480), .B2(n13190), .A(n13090), .ZN(n13091) );
  OAI21_X1 U14742 ( .B1(n13092), .B2(n13196), .A(n13091), .ZN(P3_U3163) );
  INV_X1 U14743 ( .A(n13093), .ZN(n13094) );
  NOR2_X1 U14744 ( .A1(n13095), .A2(n13094), .ZN(n13096) );
  XNOR2_X1 U14745 ( .A(n13097), .B(n13096), .ZN(n13104) );
  NOR2_X1 U14746 ( .A1(n13234), .A2(n15971), .ZN(n13101) );
  NAND2_X1 U14747 ( .A1(n13215), .A2(n13244), .ZN(n13099) );
  OAI211_X1 U14748 ( .C1(n13581), .C2(n13217), .A(n13099), .B(n13098), .ZN(
        n13100) );
  AOI211_X1 U14749 ( .C1(n13102), .C2(n13230), .A(n13101), .B(n13100), .ZN(
        n13103) );
  OAI21_X1 U14750 ( .B1(n13104), .B2(n13196), .A(n13103), .ZN(P3_U3164) );
  INV_X1 U14751 ( .A(n13107), .ZN(n13147) );
  INV_X1 U14752 ( .A(n13108), .ZN(n13110) );
  NOR3_X1 U14753 ( .A1(n13147), .A2(n13110), .A3(n13109), .ZN(n13113) );
  INV_X1 U14754 ( .A(n13111), .ZN(n13112) );
  OAI21_X1 U14755 ( .B1(n13113), .B2(n13112), .A(n13223), .ZN(n13117) );
  NOR2_X1 U14756 ( .A1(n13450), .A2(n13227), .ZN(n13115) );
  OAI22_X1 U14757 ( .A1(n13396), .A2(n13217), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15267), .ZN(n13114) );
  AOI211_X1 U14758 ( .C1(n13429), .C2(n13230), .A(n13115), .B(n13114), .ZN(
        n13116) );
  OAI211_X1 U14759 ( .C1(n13671), .C2(n13234), .A(n13117), .B(n13116), .ZN(
        P3_U3165) );
  NOR2_X1 U14760 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15264), .ZN(n13284) );
  NOR2_X1 U14761 ( .A1(n13217), .A2(n13524), .ZN(n13118) );
  AOI211_X1 U14762 ( .C1(n13215), .C2(n13551), .A(n13284), .B(n13118), .ZN(
        n13119) );
  OAI21_X1 U14763 ( .B1(n13554), .B2(n13175), .A(n13119), .ZN(n13123) );
  AOI211_X1 U14764 ( .C1(n13121), .C2(n13120), .A(n13196), .B(n7272), .ZN(
        n13122) );
  AOI211_X1 U14765 ( .C1(n13644), .C2(n13190), .A(n13123), .B(n13122), .ZN(
        n13124) );
  INV_X1 U14766 ( .A(n13124), .ZN(P3_U3166) );
  XNOR2_X1 U14767 ( .A(n13126), .B(n13125), .ZN(n13127) );
  NAND2_X1 U14768 ( .A1(n13127), .A2(n13223), .ZN(n13135) );
  AOI21_X1 U14769 ( .B1(n13190), .B2(n13129), .A(n13128), .ZN(n13134) );
  AOI22_X1 U14770 ( .A1(n13225), .A2(n13249), .B1(n13215), .B2(n13251), .ZN(
        n13133) );
  INV_X1 U14771 ( .A(n13130), .ZN(n13131) );
  NAND2_X1 U14772 ( .A1(n13230), .A2(n13131), .ZN(n13132) );
  NAND4_X1 U14773 ( .A1(n13135), .A2(n13134), .A3(n13133), .A4(n13132), .ZN(
        P3_U3167) );
  XNOR2_X1 U14774 ( .A(n13136), .B(n13552), .ZN(n13137) );
  XNOR2_X1 U14775 ( .A(n13138), .B(n13137), .ZN(n13143) );
  NAND2_X1 U14776 ( .A1(n13215), .A2(n13565), .ZN(n13139) );
  NAND2_X1 U14777 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13306)
         );
  OAI211_X1 U14778 ( .C1(n13536), .C2(n13217), .A(n13139), .B(n13306), .ZN(
        n13141) );
  NOR2_X1 U14779 ( .A1(n13700), .A2(n13234), .ZN(n13140) );
  AOI211_X1 U14780 ( .C1(n13540), .C2(n13230), .A(n13141), .B(n13140), .ZN(
        n13142) );
  OAI21_X1 U14781 ( .B1(n13143), .B2(n13196), .A(n13142), .ZN(P3_U3168) );
  INV_X1 U14782 ( .A(n13144), .ZN(n13146) );
  NOR3_X1 U14783 ( .A1(n7187), .A2(n13146), .A3(n13145), .ZN(n13148) );
  OAI21_X1 U14784 ( .B1(n13148), .B2(n13147), .A(n13223), .ZN(n13152) );
  NOR2_X1 U14785 ( .A1(n13227), .A2(n13462), .ZN(n13150) );
  INV_X1 U14786 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n15354) );
  OAI22_X1 U14787 ( .A1(n13437), .A2(n13217), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15354), .ZN(n13149) );
  AOI211_X1 U14788 ( .C1(n13442), .C2(n13230), .A(n13150), .B(n13149), .ZN(
        n13151) );
  OAI211_X1 U14789 ( .C1(n13234), .C2(n13675), .A(n13152), .B(n13151), .ZN(
        P3_U3169) );
  OAI21_X1 U14790 ( .B1(n13155), .B2(n13154), .A(n13153), .ZN(n13156) );
  NAND2_X1 U14791 ( .A1(n13156), .A2(n13223), .ZN(n13162) );
  AOI21_X1 U14792 ( .B1(n13190), .B2(n15906), .A(n13157), .ZN(n13161) );
  AOI22_X1 U14793 ( .A1(n13225), .A2(n13250), .B1(n13215), .B2(n15847), .ZN(
        n13160) );
  NAND2_X1 U14794 ( .A1(n13230), .A2(n13158), .ZN(n13159) );
  NAND4_X1 U14795 ( .A1(n13162), .A2(n13161), .A3(n13160), .A4(n13159), .ZN(
        P3_U3170) );
  OAI211_X1 U14796 ( .C1(n13165), .C2(n13164), .A(n7303), .B(n13223), .ZN(
        n13169) );
  OAI22_X1 U14797 ( .A1(n13217), .A2(n13461), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15261), .ZN(n13167) );
  NOR2_X1 U14798 ( .A1(n13227), .A2(n13525), .ZN(n13166) );
  AOI211_X1 U14799 ( .C1(n13497), .C2(n13230), .A(n13167), .B(n13166), .ZN(
        n13168) );
  OAI211_X1 U14800 ( .C1(n13691), .C2(n13234), .A(n13169), .B(n13168), .ZN(
        P3_U3173) );
  XOR2_X1 U14801 ( .A(n13171), .B(n13170), .Z(n13179) );
  NOR2_X1 U14802 ( .A1(n13217), .A2(n13228), .ZN(n13172) );
  AOI211_X1 U14803 ( .C1(n13215), .C2(n13243), .A(n13173), .B(n13172), .ZN(
        n13174) );
  OAI21_X1 U14804 ( .B1(n13176), .B2(n13175), .A(n13174), .ZN(n13177) );
  AOI21_X1 U14805 ( .B1(n13657), .B2(n13190), .A(n13177), .ZN(n13178) );
  OAI21_X1 U14806 ( .B1(n13179), .B2(n13196), .A(n13178), .ZN(P3_U3174) );
  INV_X1 U14807 ( .A(n13181), .ZN(n13182) );
  AOI21_X1 U14808 ( .B1(n13474), .B2(n13180), .A(n13182), .ZN(n13188) );
  AOI22_X1 U14809 ( .A1(n13215), .A2(n13493), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13184) );
  NAND2_X1 U14810 ( .A1(n13230), .A2(n13467), .ZN(n13183) );
  OAI211_X1 U14811 ( .C1(n13462), .C2(n13217), .A(n13184), .B(n13183), .ZN(
        n13185) );
  AOI21_X1 U14812 ( .B1(n13186), .B2(n13190), .A(n13185), .ZN(n13187) );
  OAI21_X1 U14813 ( .B1(n13188), .B2(n13196), .A(n13187), .ZN(P3_U3175) );
  INV_X1 U14814 ( .A(n13189), .ZN(n13201) );
  AOI22_X1 U14815 ( .A1(n13215), .A2(n13245), .B1(n13191), .B2(n13190), .ZN(
        n13192) );
  NAND2_X1 U14816 ( .A1(P3_REG3_REG_11__SCAN_IN), .A2(P3_U3151), .ZN(n15821)
         );
  OAI211_X1 U14817 ( .C1(n13193), .C2(n13217), .A(n13192), .B(n15821), .ZN(
        n13200) );
  INV_X1 U14818 ( .A(n13194), .ZN(n13195) );
  AOI211_X1 U14819 ( .C1(n13201), .C2(n13230), .A(n13200), .B(n13199), .ZN(
        n13202) );
  INV_X1 U14820 ( .A(n13202), .ZN(P3_U3176) );
  INV_X1 U14821 ( .A(n13636), .ZN(n13210) );
  OAI211_X1 U14822 ( .C1(n13205), .C2(n13204), .A(n13203), .B(n13223), .ZN(
        n13209) );
  NOR2_X1 U14823 ( .A1(n15253), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13327) );
  AOI21_X1 U14824 ( .B1(n13225), .B2(n13492), .A(n13327), .ZN(n13206) );
  OAI21_X1 U14825 ( .B1(n13524), .B2(n13227), .A(n13206), .ZN(n13207) );
  AOI21_X1 U14826 ( .B1(n13526), .B2(n13230), .A(n13207), .ZN(n13208) );
  OAI211_X1 U14827 ( .C1(n13210), .C2(n13234), .A(n13209), .B(n13208), .ZN(
        P3_U3178) );
  OAI21_X1 U14828 ( .B1(n13213), .B2(n13211), .A(n13212), .ZN(n13214) );
  AOI22_X1 U14829 ( .A1(n13238), .A2(n13215), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13216) );
  OAI21_X1 U14830 ( .B1(n13412), .B2(n13217), .A(n13216), .ZN(n13218) );
  AOI21_X1 U14831 ( .B1(n13416), .B2(n13230), .A(n13218), .ZN(n13219) );
  OAI21_X1 U14832 ( .B1(n13222), .B2(n13221), .A(n13220), .ZN(n13224) );
  NAND2_X1 U14833 ( .A1(n13224), .A2(n13223), .ZN(n13233) );
  INV_X1 U14834 ( .A(n13570), .ZN(n13231) );
  INV_X1 U14835 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n15259) );
  NOR2_X1 U14836 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15259), .ZN(n13260) );
  AOI21_X1 U14837 ( .B1(n13225), .B2(n13565), .A(n13260), .ZN(n13226) );
  OAI21_X1 U14838 ( .B1(n13228), .B2(n13227), .A(n13226), .ZN(n13229) );
  AOI21_X1 U14839 ( .B1(n13231), .B2(n13230), .A(n13229), .ZN(n13232) );
  OAI211_X1 U14840 ( .C1(n13234), .C2(n13651), .A(n13233), .B(n13232), .ZN(
        P3_U3181) );
  MUX2_X1 U14841 ( .A(n13235), .B(P3_DATAO_REG_31__SCAN_IN), .S(n13240), .Z(
        P3_U3522) );
  MUX2_X1 U14842 ( .A(n13236), .B(P3_DATAO_REG_30__SCAN_IN), .S(n13240), .Z(
        P3_U3521) );
  MUX2_X1 U14843 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n13237), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14844 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n7563), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14845 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n13238), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14846 ( .A(n13423), .B(P3_DATAO_REG_24__SCAN_IN), .S(n13240), .Z(
        P3_U3515) );
  MUX2_X1 U14847 ( .A(n13239), .B(P3_DATAO_REG_23__SCAN_IN), .S(n13240), .Z(
        P3_U3514) );
  MUX2_X1 U14848 ( .A(n13474), .B(P3_DATAO_REG_22__SCAN_IN), .S(n13240), .Z(
        P3_U3513) );
  MUX2_X1 U14849 ( .A(n13493), .B(P3_DATAO_REG_21__SCAN_IN), .S(n13240), .Z(
        P3_U3512) );
  MUX2_X1 U14850 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13473), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14851 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n13492), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14852 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13241), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14853 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n13552), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14854 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n13565), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14855 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n13551), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14856 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n13564), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14857 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n13242), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14858 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n13243), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14859 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n13244), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14860 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n13245), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14861 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n13246), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U14862 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n13247), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14863 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n13248), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14864 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n13249), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14865 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n13250), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14866 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n13251), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14867 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n15847), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14868 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n13252), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14869 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n7349), .S(P3_U3897), .Z(
        P3_U3492) );
  AND2_X1 U14870 ( .A1(n13263), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n13253) );
  AOI21_X1 U14871 ( .B1(n13256), .B2(n13265), .A(n13274), .ZN(n13272) );
  NAND2_X1 U14872 ( .A1(P3_REG2_REG_14__SCAN_IN), .A2(n13263), .ZN(n13258) );
  OAI21_X1 U14873 ( .B1(n13259), .B2(P3_REG2_REG_15__SCAN_IN), .A(n13287), 
        .ZN(n13270) );
  AOI21_X1 U14874 ( .B1(n15806), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n13260), 
        .ZN(n13261) );
  OAI21_X1 U14875 ( .B1(n13362), .B2(n13285), .A(n13261), .ZN(n13269) );
  XOR2_X1 U14876 ( .A(n13285), .B(n13279), .Z(n13267) );
  MUX2_X1 U14877 ( .A(n13571), .B(n13265), .S(n13728), .Z(n13266) );
  NOR2_X1 U14878 ( .A1(n13267), .A2(n13266), .ZN(n13280) );
  AOI211_X1 U14879 ( .C1(n13267), .C2(n13266), .A(n15763), .B(n13280), .ZN(
        n13268) );
  AOI211_X1 U14880 ( .C1(n15815), .C2(n13270), .A(n13269), .B(n13268), .ZN(
        n13271) );
  OAI21_X1 U14881 ( .B1(n13272), .B2(n15800), .A(n13271), .ZN(P3_U3197) );
  INV_X1 U14882 ( .A(n13273), .ZN(n13275) );
  NAND2_X1 U14883 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n13309), .ZN(n13276) );
  OAI21_X1 U14884 ( .B1(P3_REG1_REG_16__SCAN_IN), .B2(n13309), .A(n13276), 
        .ZN(n13277) );
  NOR2_X1 U14885 ( .A1(n13278), .A2(n13277), .ZN(n13299) );
  AOI21_X1 U14886 ( .B1(n13278), .B2(n13277), .A(n13299), .ZN(n13298) );
  INV_X1 U14887 ( .A(n13279), .ZN(n13281) );
  AOI21_X1 U14888 ( .B1(n13285), .B2(n13281), .A(n13280), .ZN(n13283) );
  MUX2_X1 U14889 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n13728), .Z(n13310) );
  XNOR2_X1 U14890 ( .A(n13309), .B(n13310), .ZN(n13282) );
  NOR2_X1 U14891 ( .A1(n13283), .A2(n13282), .ZN(n13308) );
  AOI211_X1 U14892 ( .C1(n13283), .C2(n13282), .A(n15763), .B(n13308), .ZN(
        n13296) );
  AOI21_X1 U14893 ( .B1(n15806), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n13284), 
        .ZN(n13294) );
  NAND2_X1 U14894 ( .A1(n13286), .A2(n13285), .ZN(n13288) );
  AOI22_X1 U14895 ( .A1(n13289), .A2(n13555), .B1(P3_REG2_REG_16__SCAN_IN), 
        .B2(n13309), .ZN(n13290) );
  OAI21_X1 U14896 ( .B1(n13291), .B2(n13290), .A(n13301), .ZN(n13292) );
  NAND2_X1 U14897 ( .A1(n15815), .A2(n13292), .ZN(n13293) );
  OAI211_X1 U14898 ( .C1(n13362), .C2(n13309), .A(n13294), .B(n13293), .ZN(
        n13295) );
  NOR2_X1 U14899 ( .A1(n13296), .A2(n13295), .ZN(n13297) );
  OAI21_X1 U14900 ( .B1(n13298), .B2(n15800), .A(n13297), .ZN(P3_U3198) );
  AOI21_X1 U14901 ( .B1(n13642), .B2(n13300), .A(n13331), .ZN(n13316) );
  INV_X1 U14902 ( .A(n13318), .ZN(n13332) );
  NAND2_X1 U14903 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n13309), .ZN(n13302) );
  OAI21_X1 U14904 ( .B1(P3_REG2_REG_17__SCAN_IN), .B2(n13303), .A(n13323), 
        .ZN(n13304) );
  INV_X1 U14905 ( .A(n13304), .ZN(n13307) );
  NAND2_X1 U14906 ( .A1(n15806), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n13305) );
  OAI211_X1 U14907 ( .C1(n15742), .C2(n13307), .A(n13306), .B(n13305), .ZN(
        n13314) );
  AOI21_X1 U14908 ( .B1(n13310), .B2(n13309), .A(n13308), .ZN(n13312) );
  MUX2_X1 U14909 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13728), .Z(n13319) );
  XNOR2_X1 U14910 ( .A(n13318), .B(n13319), .ZN(n13311) );
  NOR2_X1 U14911 ( .A1(n13312), .A2(n13311), .ZN(n13317) );
  AOI211_X1 U14912 ( .C1(n13312), .C2(n13311), .A(n15763), .B(n13317), .ZN(
        n13313) );
  AOI211_X1 U14913 ( .C1(n15808), .C2(n13332), .A(n13314), .B(n13313), .ZN(
        n13315) );
  OAI21_X1 U14914 ( .B1(n13316), .B2(n15800), .A(n13315), .ZN(P3_U3199) );
  MUX2_X1 U14915 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n13728), .Z(n13321) );
  XNOR2_X1 U14916 ( .A(n13351), .B(n13350), .ZN(n13320) );
  NOR2_X1 U14917 ( .A1(n13320), .A2(n13321), .ZN(n13349) );
  AOI21_X1 U14918 ( .B1(n13321), .B2(n13320), .A(n13349), .ZN(n13343) );
  INV_X1 U14919 ( .A(n13322), .ZN(n13324) );
  NOR2_X1 U14920 ( .A1(n13350), .A2(n13528), .ZN(n13356) );
  NAND2_X1 U14921 ( .A1(n13350), .A2(n13528), .ZN(n13355) );
  INV_X1 U14922 ( .A(n13355), .ZN(n13325) );
  NOR2_X1 U14923 ( .A1(n13356), .A2(n13325), .ZN(n13326) );
  XNOR2_X1 U14924 ( .A(n13357), .B(n13326), .ZN(n13330) );
  AOI21_X1 U14925 ( .B1(n15806), .B2(P3_ADDR_REG_18__SCAN_IN), .A(n13327), 
        .ZN(n13328) );
  OAI21_X1 U14926 ( .B1(n13362), .B2(n13334), .A(n13328), .ZN(n13329) );
  AOI21_X1 U14927 ( .B1(n13330), .B2(n15815), .A(n13329), .ZN(n13342) );
  OR2_X1 U14928 ( .A1(n13333), .A2(n13332), .ZN(n13338) );
  NAND2_X1 U14929 ( .A1(n13334), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n13344) );
  NAND2_X1 U14930 ( .A1(n13350), .A2(n13335), .ZN(n13336) );
  NAND2_X1 U14931 ( .A1(n13344), .A2(n13336), .ZN(n13337) );
  AND3_X1 U14932 ( .A1(n13339), .A2(n13338), .A3(n13337), .ZN(n13340) );
  OAI21_X1 U14933 ( .B1(n13346), .B2(n13340), .A(n15819), .ZN(n13341) );
  OAI211_X1 U14934 ( .C1(n13343), .C2(n15763), .A(n13342), .B(n13341), .ZN(
        P3_U3200) );
  INV_X1 U14935 ( .A(n13344), .ZN(n13345) );
  NOR2_X1 U14936 ( .A1(n13346), .A2(n13345), .ZN(n13348) );
  XNOR2_X1 U14937 ( .A(n13361), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13352) );
  INV_X1 U14938 ( .A(n13352), .ZN(n13347) );
  XNOR2_X1 U14939 ( .A(n13348), .B(n13347), .ZN(n13370) );
  AOI21_X1 U14940 ( .B1(n13351), .B2(n13350), .A(n13349), .ZN(n13354) );
  XNOR2_X1 U14941 ( .A(n13361), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n13358) );
  MUX2_X1 U14942 ( .A(n13358), .B(n13352), .S(n13728), .Z(n13353) );
  XNOR2_X1 U14943 ( .A(n13354), .B(n13353), .ZN(n13368) );
  INV_X1 U14944 ( .A(n13358), .ZN(n13359) );
  XNOR2_X1 U14945 ( .A(n13360), .B(n13359), .ZN(n13366) );
  NOR2_X1 U14946 ( .A1(n13362), .A2(n13361), .ZN(n13363) );
  AOI211_X1 U14947 ( .C1(P3_ADDR_REG_19__SCAN_IN), .C2(n15806), .A(n13364), 
        .B(n13363), .ZN(n13365) );
  OAI21_X1 U14948 ( .B1(n13366), .B2(n15742), .A(n13365), .ZN(n13367) );
  AOI21_X1 U14949 ( .B1(n13368), .B2(n15814), .A(n13367), .ZN(n13369) );
  OAI21_X1 U14950 ( .B1(n13370), .B2(n15800), .A(n13369), .ZN(P3_U3201) );
  INV_X1 U14951 ( .A(n13371), .ZN(n13372) );
  NAND2_X1 U14952 ( .A1(n13372), .A2(n13541), .ZN(n13382) );
  NAND3_X1 U14953 ( .A1(n13382), .A2(n15867), .A3(n16038), .ZN(n13377) );
  OAI21_X1 U14954 ( .B1(n15867), .B2(P3_REG2_REG_31__SCAN_IN), .A(n13377), 
        .ZN(n13375) );
  OAI21_X1 U14955 ( .B1(n13376), .B2(n13587), .A(n13375), .ZN(P3_U3202) );
  OAI21_X1 U14956 ( .B1(n15867), .B2(P3_REG2_REG_30__SCAN_IN), .A(n13377), 
        .ZN(n13378) );
  OAI21_X1 U14957 ( .B1(n13379), .B2(n13587), .A(n13378), .ZN(P3_U3203) );
  INV_X1 U14958 ( .A(n13380), .ZN(n13387) );
  NAND2_X1 U14959 ( .A1(n15869), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n13381) );
  OAI211_X1 U14960 ( .C1(n13383), .C2(n13587), .A(n13382), .B(n13381), .ZN(
        n13384) );
  AOI21_X1 U14961 ( .B1(n13385), .B2(n13592), .A(n13384), .ZN(n13386) );
  OAI21_X1 U14962 ( .B1(n13387), .B2(n15869), .A(n13386), .ZN(P3_U3204) );
  AOI22_X1 U14963 ( .A1(n13388), .A2(n13541), .B1(n15869), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n13389) );
  OAI21_X1 U14964 ( .B1(n13597), .B2(n13587), .A(n13389), .ZN(n13390) );
  AOI21_X1 U14965 ( .B1(n13391), .B2(n13592), .A(n13390), .ZN(n13392) );
  OAI21_X1 U14966 ( .B1(n13393), .B2(n15869), .A(n13392), .ZN(P3_U3205) );
  OAI22_X1 U14967 ( .A1(n13397), .A2(n13580), .B1(n13396), .B2(n13582), .ZN(
        n13403) );
  NAND2_X1 U14968 ( .A1(n13399), .A2(n13398), .ZN(n13400) );
  AOI21_X1 U14969 ( .B1(n13401), .B2(n13400), .A(n13578), .ZN(n13402) );
  NAND2_X1 U14970 ( .A1(n13599), .A2(n13500), .ZN(n13407) );
  AOI22_X1 U14971 ( .A1(n13405), .A2(n13541), .B1(n15869), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n13406) );
  OAI211_X1 U14972 ( .C1(n13664), .C2(n13587), .A(n13407), .B(n13406), .ZN(
        n13408) );
  AOI21_X1 U14973 ( .B1(n13598), .B2(n15867), .A(n13408), .ZN(n13409) );
  INV_X1 U14974 ( .A(n13409), .ZN(P3_U3206) );
  XNOR2_X1 U14975 ( .A(n13410), .B(n13413), .ZN(n13411) );
  OAI222_X1 U14976 ( .A1(n13580), .A2(n13412), .B1(n13582), .B2(n13437), .C1(
        n13578), .C2(n13411), .ZN(n13601) );
  INV_X1 U14977 ( .A(n13601), .ZN(n13420) );
  NAND2_X1 U14978 ( .A1(n13414), .A2(n13413), .ZN(n13415) );
  AOI22_X1 U14979 ( .A1(n13416), .A2(n13541), .B1(n15869), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n13417) );
  OAI21_X1 U14980 ( .B1(n7564), .B2(n13587), .A(n13417), .ZN(n13418) );
  AOI21_X1 U14981 ( .B1(n13602), .B2(n13592), .A(n13418), .ZN(n13419) );
  OAI21_X1 U14982 ( .B1(n13420), .B2(n15869), .A(n13419), .ZN(P3_U3207) );
  OAI211_X1 U14983 ( .C1(n7230), .C2(n13422), .A(n15851), .B(n13421), .ZN(
        n13425) );
  AOI22_X1 U14984 ( .A1(n7563), .A2(n15846), .B1(n15848), .B2(n13423), .ZN(
        n13424) );
  NAND2_X1 U14985 ( .A1(n13425), .A2(n13424), .ZN(n13605) );
  INV_X1 U14986 ( .A(n13605), .ZN(n13433) );
  OAI21_X1 U14987 ( .B1(n13428), .B2(n13427), .A(n13426), .ZN(n13606) );
  AOI22_X1 U14988 ( .A1(n15869), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n13429), 
        .B2(n13541), .ZN(n13430) );
  OAI21_X1 U14989 ( .B1(n13671), .B2(n13587), .A(n13430), .ZN(n13431) );
  AOI21_X1 U14990 ( .B1(n13606), .B2(n13592), .A(n13431), .ZN(n13432) );
  OAI21_X1 U14991 ( .B1(n13433), .B2(n15869), .A(n13432), .ZN(P3_U3208) );
  XNOR2_X1 U14992 ( .A(n13434), .B(n13435), .ZN(n13441) );
  XNOR2_X1 U14993 ( .A(n13436), .B(n13435), .ZN(n13439) );
  OAI22_X1 U14994 ( .A1(n13437), .A2(n13580), .B1(n13462), .B2(n13582), .ZN(
        n13438) );
  AOI21_X1 U14995 ( .B1(n13439), .B2(n15851), .A(n13438), .ZN(n13440) );
  OAI21_X1 U14996 ( .B1(n15855), .B2(n13441), .A(n13440), .ZN(n13609) );
  INV_X1 U14997 ( .A(n13609), .ZN(n13446) );
  INV_X1 U14998 ( .A(n13441), .ZN(n13610) );
  AOI22_X1 U14999 ( .A1(n15869), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n13541), 
        .B2(n13442), .ZN(n13443) );
  OAI21_X1 U15000 ( .B1(n13675), .B2(n13587), .A(n13443), .ZN(n13444) );
  AOI21_X1 U15001 ( .B1(n13610), .B2(n13500), .A(n13444), .ZN(n13445) );
  OAI21_X1 U15002 ( .B1(n13446), .B2(n15869), .A(n13445), .ZN(P3_U3209) );
  XNOR2_X1 U15003 ( .A(n13447), .B(n13452), .ZN(n13448) );
  OAI222_X1 U15004 ( .A1(n13580), .A2(n13450), .B1(n13582), .B2(n13449), .C1(
        n13578), .C2(n13448), .ZN(n13613) );
  INV_X1 U15005 ( .A(n13613), .ZN(n13457) );
  XNOR2_X1 U15006 ( .A(n13451), .B(n13452), .ZN(n13614) );
  AOI22_X1 U15007 ( .A1(n15869), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n13541), 
        .B2(n13453), .ZN(n13454) );
  OAI21_X1 U15008 ( .B1(n13679), .B2(n13587), .A(n13454), .ZN(n13455) );
  AOI21_X1 U15009 ( .B1(n13614), .B2(n13592), .A(n13455), .ZN(n13456) );
  OAI21_X1 U15010 ( .B1(n13457), .B2(n15869), .A(n13456), .ZN(P3_U3210) );
  XNOR2_X1 U15011 ( .A(n13458), .B(n13460), .ZN(n13466) );
  XNOR2_X1 U15012 ( .A(n13459), .B(n13460), .ZN(n13464) );
  OAI22_X1 U15013 ( .A1(n13462), .A2(n13580), .B1(n13461), .B2(n13582), .ZN(
        n13463) );
  AOI21_X1 U15014 ( .B1(n13464), .B2(n15851), .A(n13463), .ZN(n13465) );
  OAI21_X1 U15015 ( .B1(n15855), .B2(n13466), .A(n13465), .ZN(n13617) );
  INV_X1 U15016 ( .A(n13617), .ZN(n13471) );
  INV_X1 U15017 ( .A(n13466), .ZN(n13618) );
  AOI22_X1 U15018 ( .A1(n15869), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n13541), 
        .B2(n13467), .ZN(n13468) );
  OAI21_X1 U15019 ( .B1(n13683), .B2(n13587), .A(n13468), .ZN(n13469) );
  AOI21_X1 U15020 ( .B1(n13618), .B2(n13500), .A(n13469), .ZN(n13470) );
  OAI21_X1 U15021 ( .B1(n13471), .B2(n15869), .A(n13470), .ZN(P3_U3211) );
  XNOR2_X1 U15022 ( .A(n13472), .B(n13475), .ZN(n13479) );
  AOI22_X1 U15023 ( .A1(n13474), .A2(n15846), .B1(n15848), .B2(n13473), .ZN(
        n13478) );
  XNOR2_X1 U15024 ( .A(n13476), .B(n13475), .ZN(n13622) );
  NAND2_X1 U15025 ( .A1(n13622), .A2(n15977), .ZN(n13477) );
  OAI211_X1 U15026 ( .C1(n13479), .C2(n13578), .A(n13478), .B(n13477), .ZN(
        n13621) );
  INV_X1 U15027 ( .A(n13621), .ZN(n13485) );
  INV_X1 U15028 ( .A(n13480), .ZN(n13687) );
  AOI22_X1 U15029 ( .A1(n15869), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n13541), 
        .B2(n13481), .ZN(n13482) );
  OAI21_X1 U15030 ( .B1(n13687), .B2(n13587), .A(n13482), .ZN(n13483) );
  AOI21_X1 U15031 ( .B1(n13622), .B2(n13500), .A(n13483), .ZN(n13484) );
  OAI21_X1 U15032 ( .B1(n13485), .B2(n15869), .A(n13484), .ZN(P3_U3212) );
  OR2_X1 U15033 ( .A1(n13486), .A2(n13489), .ZN(n13487) );
  NAND2_X1 U15034 ( .A1(n13488), .A2(n13487), .ZN(n13496) );
  XNOR2_X1 U15035 ( .A(n13490), .B(n13489), .ZN(n13491) );
  NAND2_X1 U15036 ( .A1(n13491), .A2(n15851), .ZN(n13495) );
  AOI22_X1 U15037 ( .A1(n13493), .A2(n15846), .B1(n15848), .B2(n13492), .ZN(
        n13494) );
  OAI211_X1 U15038 ( .C1(n15855), .C2(n13496), .A(n13495), .B(n13494), .ZN(
        n13625) );
  INV_X1 U15039 ( .A(n13625), .ZN(n13502) );
  INV_X1 U15040 ( .A(n13496), .ZN(n13626) );
  AOI22_X1 U15041 ( .A1(n15869), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n13541), 
        .B2(n13497), .ZN(n13498) );
  OAI21_X1 U15042 ( .B1(n13691), .B2(n13587), .A(n13498), .ZN(n13499) );
  AOI21_X1 U15043 ( .B1(n13626), .B2(n13500), .A(n13499), .ZN(n13501) );
  OAI21_X1 U15044 ( .B1(n13502), .B2(n15869), .A(n13501), .ZN(P3_U3213) );
  XOR2_X1 U15045 ( .A(n13509), .B(n13503), .Z(n13504) );
  OAI222_X1 U15046 ( .A1(n13582), .A2(n13536), .B1(n13580), .B2(n13505), .C1(
        n13578), .C2(n13504), .ZN(n13630) );
  INV_X1 U15047 ( .A(n13630), .ZN(n13516) );
  INV_X1 U15048 ( .A(n13506), .ZN(n13507) );
  OAI22_X1 U15049 ( .A1(n15867), .A2(n13508), .B1(n13507), .B2(n15860), .ZN(
        n13513) );
  INV_X1 U15050 ( .A(n13631), .ZN(n13511) );
  AND2_X1 U15051 ( .A1(n13510), .A2(n13509), .ZN(n13629) );
  NOR3_X1 U15052 ( .A1(n13511), .A2(n13629), .A3(n13532), .ZN(n13512) );
  AOI211_X1 U15053 ( .C1(n13557), .C2(n13514), .A(n13513), .B(n13512), .ZN(
        n13515) );
  OAI21_X1 U15054 ( .B1(n13516), .B2(n15869), .A(n13515), .ZN(P3_U3214) );
  INV_X1 U15055 ( .A(n13522), .ZN(n13517) );
  XNOR2_X1 U15056 ( .A(n13518), .B(n13517), .ZN(n13638) );
  INV_X1 U15057 ( .A(n13519), .ZN(n13520) );
  AOI21_X1 U15058 ( .B1(n13522), .B2(n13521), .A(n13520), .ZN(n13523) );
  OAI222_X1 U15059 ( .A1(n13580), .A2(n13525), .B1(n13582), .B2(n13524), .C1(
        n13578), .C2(n13523), .ZN(n13635) );
  NAND2_X1 U15060 ( .A1(n13635), .A2(n15867), .ZN(n13531) );
  INV_X1 U15061 ( .A(n13526), .ZN(n13527) );
  OAI22_X1 U15062 ( .A1(n15867), .A2(n13528), .B1(n13527), .B2(n15860), .ZN(
        n13529) );
  AOI21_X1 U15063 ( .B1(n13636), .B2(n13557), .A(n13529), .ZN(n13530) );
  OAI211_X1 U15064 ( .C1(n13638), .C2(n13532), .A(n13531), .B(n13530), .ZN(
        P3_U3215) );
  XNOR2_X1 U15065 ( .A(n13533), .B(n13538), .ZN(n13534) );
  OAI222_X1 U15066 ( .A1(n13580), .A2(n13536), .B1(n13582), .B2(n13535), .C1(
        n13578), .C2(n13534), .ZN(n13640) );
  INV_X1 U15067 ( .A(n13640), .ZN(n13545) );
  OAI21_X1 U15068 ( .B1(n13539), .B2(n13538), .A(n13537), .ZN(n13641) );
  AOI22_X1 U15069 ( .A1(n15869), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n13541), 
        .B2(n13540), .ZN(n13542) );
  OAI21_X1 U15070 ( .B1(n13700), .B2(n13587), .A(n13542), .ZN(n13543) );
  AOI21_X1 U15071 ( .B1(n13641), .B2(n13592), .A(n13543), .ZN(n13544) );
  OAI21_X1 U15072 ( .B1(n13545), .B2(n15869), .A(n13544), .ZN(P3_U3216) );
  NAND2_X1 U15073 ( .A1(n13563), .A2(n13567), .ZN(n13562) );
  NAND2_X1 U15074 ( .A1(n13562), .A2(n13548), .ZN(n13550) );
  XNOR2_X1 U15075 ( .A(n13550), .B(n13549), .ZN(n13553) );
  AOI222_X1 U15076 ( .A1(n15851), .A2(n13553), .B1(n13552), .B2(n15846), .C1(
        n13551), .C2(n15848), .ZN(n13647) );
  OAI22_X1 U15077 ( .A1(n15867), .A2(n13555), .B1(n13554), .B2(n15860), .ZN(
        n13556) );
  AOI21_X1 U15078 ( .B1(n13644), .B2(n13557), .A(n13556), .ZN(n13561) );
  XNOR2_X1 U15079 ( .A(n13559), .B(n13558), .ZN(n13645) );
  NAND2_X1 U15080 ( .A1(n13645), .A2(n13592), .ZN(n13560) );
  OAI211_X1 U15081 ( .C1(n13647), .C2(n15869), .A(n13561), .B(n13560), .ZN(
        P3_U3217) );
  OAI21_X1 U15082 ( .B1(n13563), .B2(n13567), .A(n13562), .ZN(n13566) );
  AOI222_X1 U15083 ( .A1(n15851), .A2(n13566), .B1(n13565), .B2(n15846), .C1(
        n13564), .C2(n15848), .ZN(n13650) );
  OAI21_X1 U15084 ( .B1(n13569), .B2(n8437), .A(n13568), .ZN(n13648) );
  NOR2_X1 U15085 ( .A1(n13651), .A2(n13587), .ZN(n13573) );
  OAI22_X1 U15086 ( .A1(n15867), .A2(n13571), .B1(n13570), .B2(n15860), .ZN(
        n13572) );
  AOI211_X1 U15087 ( .C1(n13648), .C2(n13592), .A(n13573), .B(n13572), .ZN(
        n13574) );
  OAI21_X1 U15088 ( .B1(n13650), .B2(n15869), .A(n13574), .ZN(P3_U3218) );
  XNOR2_X1 U15089 ( .A(n13576), .B(n13575), .ZN(n13577) );
  OAI222_X1 U15090 ( .A1(n13582), .A2(n13581), .B1(n13580), .B2(n13579), .C1(
        n13578), .C2(n13577), .ZN(n13652) );
  INV_X1 U15091 ( .A(n13652), .ZN(n13594) );
  INV_X1 U15092 ( .A(n13583), .ZN(n13584) );
  AOI21_X1 U15093 ( .B1(n13586), .B2(n13585), .A(n13584), .ZN(n13653) );
  NOR2_X1 U15094 ( .A1(n13706), .A2(n13587), .ZN(n13591) );
  OAI22_X1 U15095 ( .A1(n15867), .A2(n13589), .B1(n13588), .B2(n15860), .ZN(
        n13590) );
  AOI211_X1 U15096 ( .C1(n13653), .C2(n13592), .A(n13591), .B(n13590), .ZN(
        n13593) );
  OAI21_X1 U15097 ( .B1(n13594), .B2(n15869), .A(n13593), .ZN(P3_U3219) );
  OAI21_X1 U15098 ( .B1(n13597), .B2(n13656), .A(n13596), .ZN(P3_U3487) );
  INV_X1 U15099 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n13600) );
  INV_X1 U15100 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13603) );
  AOI21_X1 U15101 ( .B1(n13602), .B2(n13658), .A(n13601), .ZN(n13665) );
  MUX2_X1 U15102 ( .A(n13603), .B(n13665), .S(n16039), .Z(n13604) );
  OAI21_X1 U15103 ( .B1(n7564), .B2(n13656), .A(n13604), .ZN(P3_U3485) );
  INV_X1 U15104 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13607) );
  AOI21_X1 U15105 ( .B1(n13658), .B2(n13606), .A(n13605), .ZN(n13668) );
  MUX2_X1 U15106 ( .A(n13607), .B(n13668), .S(n16039), .Z(n13608) );
  OAI21_X1 U15107 ( .B1(n13671), .B2(n13656), .A(n13608), .ZN(P3_U3484) );
  INV_X1 U15108 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13611) );
  AOI21_X1 U15109 ( .B1(n15857), .B2(n13610), .A(n13609), .ZN(n13672) );
  MUX2_X1 U15110 ( .A(n13611), .B(n13672), .S(n16039), .Z(n13612) );
  OAI21_X1 U15111 ( .B1(n13656), .B2(n13675), .A(n13612), .ZN(P3_U3483) );
  INV_X1 U15112 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13615) );
  AOI21_X1 U15113 ( .B1(n13614), .B2(n13658), .A(n13613), .ZN(n13676) );
  MUX2_X1 U15114 ( .A(n13615), .B(n13676), .S(n16039), .Z(n13616) );
  OAI21_X1 U15115 ( .B1(n13679), .B2(n13656), .A(n13616), .ZN(P3_U3482) );
  INV_X1 U15116 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13619) );
  AOI21_X1 U15117 ( .B1(n15857), .B2(n13618), .A(n13617), .ZN(n13680) );
  MUX2_X1 U15118 ( .A(n13619), .B(n13680), .S(n16039), .Z(n13620) );
  OAI21_X1 U15119 ( .B1(n13683), .B2(n13656), .A(n13620), .ZN(P3_U3481) );
  INV_X1 U15120 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13623) );
  AOI21_X1 U15121 ( .B1(n15857), .B2(n13622), .A(n13621), .ZN(n13684) );
  MUX2_X1 U15122 ( .A(n13623), .B(n13684), .S(n16039), .Z(n13624) );
  OAI21_X1 U15123 ( .B1(n13687), .B2(n13656), .A(n13624), .ZN(P3_U3480) );
  INV_X1 U15124 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13627) );
  AOI21_X1 U15125 ( .B1(n15857), .B2(n13626), .A(n13625), .ZN(n13688) );
  MUX2_X1 U15126 ( .A(n13627), .B(n13688), .S(n16039), .Z(n13628) );
  OAI21_X1 U15127 ( .B1(n13691), .B2(n13656), .A(n13628), .ZN(P3_U3479) );
  NOR2_X1 U15128 ( .A1(n13629), .A2(n13639), .ZN(n13632) );
  AOI21_X1 U15129 ( .B1(n13632), .B2(n13631), .A(n13630), .ZN(n13692) );
  MUX2_X1 U15130 ( .A(n13633), .B(n13692), .S(n16039), .Z(n13634) );
  OAI21_X1 U15131 ( .B1(n13695), .B2(n13656), .A(n13634), .ZN(P3_U3478) );
  AOI21_X1 U15132 ( .B1(n15907), .B2(n13636), .A(n13635), .ZN(n13637) );
  OAI21_X1 U15133 ( .B1(n13639), .B2(n13638), .A(n13637), .ZN(n13696) );
  MUX2_X1 U15134 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n13696), .S(n16039), .Z(
        P3_U3477) );
  AOI21_X1 U15135 ( .B1(n13658), .B2(n13641), .A(n13640), .ZN(n13697) );
  MUX2_X1 U15136 ( .A(n13642), .B(n13697), .S(n16039), .Z(n13643) );
  OAI21_X1 U15137 ( .B1(n13656), .B2(n13700), .A(n13643), .ZN(P3_U3476) );
  AOI22_X1 U15138 ( .A1(n13645), .A2(n13658), .B1(n15907), .B2(n13644), .ZN(
        n13646) );
  NAND2_X1 U15139 ( .A1(n13647), .A2(n13646), .ZN(n13701) );
  MUX2_X1 U15140 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n13701), .S(n16039), .Z(
        P3_U3475) );
  NAND2_X1 U15141 ( .A1(n13648), .A2(n13658), .ZN(n13649) );
  OAI211_X1 U15142 ( .C1(n15970), .C2(n13651), .A(n13650), .B(n13649), .ZN(
        n13702) );
  MUX2_X1 U15143 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n13702), .S(n16039), .Z(
        P3_U3474) );
  AOI21_X1 U15144 ( .B1(n13653), .B2(n13658), .A(n13652), .ZN(n13703) );
  MUX2_X1 U15145 ( .A(n13654), .B(n13703), .S(n16039), .Z(n13655) );
  OAI21_X1 U15146 ( .B1(n13656), .B2(n13706), .A(n13655), .ZN(P3_U3473) );
  AOI22_X1 U15147 ( .A1(n13659), .A2(n13658), .B1(n13657), .B2(n15907), .ZN(
        n13660) );
  NAND2_X1 U15148 ( .A1(n13661), .A2(n13660), .ZN(n13708) );
  MUX2_X1 U15149 ( .A(P3_REG1_REG_13__SCAN_IN), .B(n13708), .S(n16039), .Z(
        P3_U3472) );
  MUX2_X1 U15150 ( .A(n13666), .B(n13665), .S(n16042), .Z(n13667) );
  OAI21_X1 U15151 ( .B1(n7564), .B2(n13707), .A(n13667), .ZN(P3_U3453) );
  MUX2_X1 U15152 ( .A(n13669), .B(n13668), .S(n16042), .Z(n13670) );
  OAI21_X1 U15153 ( .B1(n13671), .B2(n13707), .A(n13670), .ZN(P3_U3452) );
  MUX2_X1 U15154 ( .A(n13673), .B(n13672), .S(n16042), .Z(n13674) );
  OAI21_X1 U15155 ( .B1(n13707), .B2(n13675), .A(n13674), .ZN(P3_U3451) );
  MUX2_X1 U15156 ( .A(n13677), .B(n13676), .S(n16042), .Z(n13678) );
  OAI21_X1 U15157 ( .B1(n13679), .B2(n13707), .A(n13678), .ZN(P3_U3450) );
  MUX2_X1 U15158 ( .A(n13681), .B(n13680), .S(n16042), .Z(n13682) );
  OAI21_X1 U15159 ( .B1(n13683), .B2(n13707), .A(n13682), .ZN(P3_U3449) );
  MUX2_X1 U15160 ( .A(n13685), .B(n13684), .S(n16042), .Z(n13686) );
  OAI21_X1 U15161 ( .B1(n13687), .B2(n13707), .A(n13686), .ZN(P3_U3448) );
  INV_X1 U15162 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13689) );
  MUX2_X1 U15163 ( .A(n13689), .B(n13688), .S(n16042), .Z(n13690) );
  OAI21_X1 U15164 ( .B1(n13691), .B2(n13707), .A(n13690), .ZN(P3_U3447) );
  INV_X1 U15165 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13693) );
  MUX2_X1 U15166 ( .A(n13693), .B(n13692), .S(n16042), .Z(n13694) );
  OAI21_X1 U15167 ( .B1(n13695), .B2(n13707), .A(n13694), .ZN(P3_U3446) );
  MUX2_X1 U15168 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n13696), .S(n16042), .Z(
        P3_U3444) );
  MUX2_X1 U15169 ( .A(n13698), .B(n13697), .S(n16042), .Z(n13699) );
  OAI21_X1 U15170 ( .B1(n13707), .B2(n13700), .A(n13699), .ZN(P3_U3441) );
  MUX2_X1 U15171 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n13701), .S(n16042), .Z(
        P3_U3438) );
  MUX2_X1 U15172 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n13702), .S(n16042), .Z(
        P3_U3435) );
  INV_X1 U15173 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13704) );
  MUX2_X1 U15174 ( .A(n13704), .B(n13703), .S(n16042), .Z(n13705) );
  OAI21_X1 U15175 ( .B1(n13707), .B2(n13706), .A(n13705), .ZN(P3_U3432) );
  MUX2_X1 U15176 ( .A(P3_REG0_REG_13__SCAN_IN), .B(n13708), .S(n16042), .Z(
        P3_U3429) );
  MUX2_X1 U15177 ( .A(P3_D_REG_1__SCAN_IN), .B(n13709), .S(n13710), .Z(
        P3_U3377) );
  MUX2_X1 U15178 ( .A(P3_D_REG_0__SCAN_IN), .B(n13711), .S(n13710), .Z(
        P3_U3376) );
  INV_X1 U15179 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13712) );
  NAND3_X1 U15180 ( .A1(n13712), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n13714) );
  OAI22_X1 U15181 ( .A1(n13715), .A2(n13714), .B1(n13713), .B2(n13723), .ZN(
        n13716) );
  AOI21_X1 U15182 ( .B1(n13718), .B2(n13717), .A(n13716), .ZN(n13719) );
  INV_X1 U15183 ( .A(n13719), .ZN(P3_U3264) );
  OAI222_X1 U15184 ( .A1(P3_U3151), .A2(n13721), .B1(n13730), .B2(n13720), 
        .C1(n15284), .C2(n13723), .ZN(P3_U3265) );
  INV_X1 U15185 ( .A(n13722), .ZN(n13726) );
  OAI222_X1 U15186 ( .A1(n13730), .A2(n13726), .B1(P3_U3151), .B2(n13725), 
        .C1(n13724), .C2(n13723), .ZN(P3_U3266) );
  INV_X1 U15187 ( .A(n13727), .ZN(n13729) );
  OAI222_X1 U15188 ( .A1(n13730), .A2(n13729), .B1(n13723), .B2(n15289), .C1(
        P3_U3151), .C2(n13728), .ZN(P3_U3268) );
  XNOR2_X1 U15189 ( .A(n14195), .B(n13773), .ZN(n13748) );
  INV_X1 U15190 ( .A(n13748), .ZN(n13853) );
  XNOR2_X1 U15191 ( .A(n16030), .B(n13805), .ZN(n13733) );
  NAND2_X1 U15192 ( .A1(n14276), .A2(n14282), .ZN(n13734) );
  NAND2_X1 U15193 ( .A1(n13733), .A2(n13734), .ZN(n13738) );
  INV_X1 U15194 ( .A(n13733), .ZN(n13736) );
  INV_X1 U15195 ( .A(n13734), .ZN(n13735) );
  NAND2_X1 U15196 ( .A1(n13736), .A2(n13735), .ZN(n13737) );
  AND2_X1 U15197 ( .A1(n13738), .A2(n13737), .ZN(n13837) );
  NAND2_X1 U15198 ( .A1(n14250), .A2(n14282), .ZN(n13740) );
  XNOR2_X1 U15199 ( .A(n13739), .B(n13740), .ZN(n13885) );
  INV_X1 U15200 ( .A(n13739), .ZN(n13742) );
  INV_X1 U15201 ( .A(n13740), .ZN(n13741) );
  NAND2_X1 U15202 ( .A1(n13742), .A2(n13741), .ZN(n13743) );
  XNOR2_X1 U15203 ( .A(n14355), .B(n13764), .ZN(n13744) );
  NOR2_X1 U15204 ( .A1(n14238), .A2(n14348), .ZN(n13745) );
  XNOR2_X1 U15205 ( .A(n13744), .B(n13745), .ZN(n13794) );
  INV_X1 U15206 ( .A(n13744), .ZN(n13746) );
  NAND2_X1 U15207 ( .A1(n13746), .A2(n13745), .ZN(n13747) );
  INV_X1 U15208 ( .A(n13855), .ZN(n13750) );
  NOR2_X1 U15209 ( .A1(n14210), .A2(n14348), .ZN(n13852) );
  XNOR2_X1 U15210 ( .A(n14182), .B(n13764), .ZN(n13751) );
  NAND2_X1 U15211 ( .A1(n14189), .A2(n14282), .ZN(n13752) );
  XNOR2_X1 U15212 ( .A(n13751), .B(n13752), .ZN(n13815) );
  INV_X1 U15213 ( .A(n13752), .ZN(n13753) );
  NAND2_X1 U15214 ( .A1(n13814), .A2(n13754), .ZN(n13755) );
  NAND2_X1 U15215 ( .A1(n13917), .A2(n8098), .ZN(n13864) );
  NOR2_X1 U15216 ( .A1(n13865), .A2(n13864), .ZN(n13863) );
  AND2_X1 U15217 ( .A1(n13755), .A2(n8101), .ZN(n13756) );
  NOR2_X1 U15218 ( .A1(n13868), .A2(n14348), .ZN(n13785) );
  XNOR2_X1 U15219 ( .A(n14134), .B(n13805), .ZN(n13761) );
  OR2_X1 U15220 ( .A1(n13828), .A2(n14151), .ZN(n13760) );
  NOR2_X1 U15221 ( .A1(n13761), .A2(n13760), .ZN(n13762) );
  AOI21_X1 U15222 ( .B1(n13761), .B2(n13760), .A(n13762), .ZN(n13845) );
  INV_X1 U15223 ( .A(n13762), .ZN(n13763) );
  XNOR2_X1 U15224 ( .A(n14384), .B(n13764), .ZN(n13766) );
  NAND2_X1 U15225 ( .A1(n13914), .A2(n14282), .ZN(n13765) );
  NOR2_X1 U15226 ( .A1(n13766), .A2(n13765), .ZN(n13767) );
  AOI21_X1 U15227 ( .B1(n13766), .B2(n13765), .A(n13767), .ZN(n13826) );
  INV_X1 U15228 ( .A(n13767), .ZN(n13768) );
  XNOR2_X1 U15229 ( .A(n14314), .B(n13805), .ZN(n13769) );
  NOR2_X1 U15230 ( .A1(n13829), .A2(n14348), .ZN(n13770) );
  XNOR2_X1 U15231 ( .A(n13769), .B(n13770), .ZN(n13897) );
  INV_X1 U15232 ( .A(n13769), .ZN(n13772) );
  INV_X1 U15233 ( .A(n13770), .ZN(n13771) );
  XNOR2_X1 U15234 ( .A(n14309), .B(n13773), .ZN(n13775) );
  NAND2_X1 U15235 ( .A1(n13912), .A2(n14282), .ZN(n13774) );
  NOR2_X1 U15236 ( .A1(n13775), .A2(n13774), .ZN(n13802) );
  AOI21_X1 U15237 ( .B1(n13775), .B2(n13774), .A(n13802), .ZN(n13776) );
  NAND2_X1 U15238 ( .A1(n13777), .A2(n13776), .ZN(n13804) );
  OAI211_X1 U15239 ( .C1(n13777), .C2(n13776), .A(n13804), .B(n13881), .ZN(
        n13783) );
  OAI22_X1 U15240 ( .A1(n13778), .A2(n14237), .B1(n13829), .B2(n14235), .ZN(
        n14084) );
  INV_X1 U15241 ( .A(n14090), .ZN(n13780) );
  OAI22_X1 U15242 ( .A1(n13780), .A2(n13902), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13779), .ZN(n13781) );
  AOI21_X1 U15243 ( .B1(n14084), .B2(n13872), .A(n13781), .ZN(n13782) );
  OAI211_X1 U15244 ( .C1(n14093), .C2(n13889), .A(n13783), .B(n13782), .ZN(
        P2_U3186) );
  OAI211_X1 U15245 ( .C1(n13786), .C2(n13785), .A(n13784), .B(n13881), .ZN(
        n13792) );
  OR2_X1 U15246 ( .A1(n13828), .A2(n14237), .ZN(n13788) );
  OR2_X1 U15247 ( .A1(n13817), .A2(n14235), .ZN(n13787) );
  NAND2_X1 U15248 ( .A1(n13788), .A2(n13787), .ZN(n14142) );
  OAI22_X1 U15249 ( .A1(n14147), .A2(n13902), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13789), .ZN(n13790) );
  AOI21_X1 U15250 ( .B1(n14142), .B2(n13872), .A(n13790), .ZN(n13791) );
  OAI211_X1 U15251 ( .C1(n14149), .C2(n13889), .A(n13792), .B(n13791), .ZN(
        P2_U3188) );
  XNOR2_X1 U15252 ( .A(n13793), .B(n13794), .ZN(n13801) );
  NAND2_X1 U15253 ( .A1(n13856), .A2(n13795), .ZN(n13797) );
  OAI211_X1 U15254 ( .C1(n13859), .C2(n14210), .A(n13797), .B(n13796), .ZN(
        n13799) );
  NOR2_X1 U15255 ( .A1(n14355), .A2(n13889), .ZN(n13798) );
  AOI211_X1 U15256 ( .C1(n13892), .C2(n14250), .A(n13799), .B(n13798), .ZN(
        n13800) );
  OAI21_X1 U15257 ( .B1(n13801), .B2(n13907), .A(n13800), .ZN(P2_U3191) );
  INV_X1 U15258 ( .A(n13802), .ZN(n13803) );
  NAND2_X1 U15259 ( .A1(n13804), .A2(n13803), .ZN(n13808) );
  MUX2_X1 U15260 ( .A(n14078), .B(n14305), .S(n14151), .Z(n13806) );
  XNOR2_X1 U15261 ( .A(n13806), .B(n13805), .ZN(n13807) );
  XNOR2_X1 U15262 ( .A(n13808), .B(n13807), .ZN(n13813) );
  AOI22_X1 U15263 ( .A1(n14275), .A2(n13910), .B1(n13912), .B2(n14274), .ZN(
        n14073) );
  INV_X1 U15264 ( .A(n14069), .ZN(n13809) );
  AOI22_X1 U15265 ( .A1(n13809), .A2(n13856), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13810) );
  OAI21_X1 U15266 ( .B1(n14073), .B2(n13900), .A(n13810), .ZN(n13811) );
  AOI21_X1 U15267 ( .B1(n14305), .B2(n13905), .A(n13811), .ZN(n13812) );
  OAI21_X1 U15268 ( .B1(n13813), .B2(n13907), .A(n13812), .ZN(P2_U3192) );
  OAI211_X1 U15269 ( .C1(n13816), .C2(n13815), .A(n13814), .B(n13881), .ZN(
        n13824) );
  OR2_X1 U15270 ( .A1(n13817), .A2(n14237), .ZN(n13819) );
  OR2_X1 U15271 ( .A1(n14210), .A2(n14235), .ZN(n13818) );
  AND2_X1 U15272 ( .A1(n13819), .A2(n13818), .ZN(n14172) );
  INV_X1 U15273 ( .A(n14172), .ZN(n13822) );
  OAI22_X1 U15274 ( .A1(n13902), .A2(n14180), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13820), .ZN(n13821) );
  AOI21_X1 U15275 ( .B1(n13822), .B2(n13872), .A(n13821), .ZN(n13823) );
  OAI211_X1 U15276 ( .C1(n14391), .C2(n13889), .A(n13824), .B(n13823), .ZN(
        P2_U3195) );
  OAI211_X1 U15277 ( .C1(n13827), .C2(n13826), .A(n13825), .B(n13881), .ZN(
        n13834) );
  OAI22_X1 U15278 ( .A1(n13829), .A2(n14237), .B1(n13828), .B2(n14235), .ZN(
        n14112) );
  INV_X1 U15279 ( .A(n14120), .ZN(n13831) );
  OAI22_X1 U15280 ( .A1(n13831), .A2(n13902), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13830), .ZN(n13832) );
  AOI21_X1 U15281 ( .B1(n14112), .B2(n13872), .A(n13832), .ZN(n13833) );
  OAI211_X1 U15282 ( .C1(n14384), .C2(n13889), .A(n13834), .B(n13833), .ZN(
        P2_U3197) );
  OAI21_X1 U15283 ( .B1(n13837), .B2(n13836), .A(n13835), .ZN(n13838) );
  NAND2_X1 U15284 ( .A1(n13838), .A2(n13881), .ZN(n13843) );
  NAND2_X1 U15285 ( .A1(n13887), .A2(n14250), .ZN(n13840) );
  OAI211_X1 U15286 ( .C1(n13902), .C2(n14256), .A(n13840), .B(n13839), .ZN(
        n13841) );
  AOI21_X1 U15287 ( .B1(n13892), .B2(n14249), .A(n13841), .ZN(n13842) );
  OAI211_X1 U15288 ( .C1(n16030), .C2(n13889), .A(n13843), .B(n13842), .ZN(
        P2_U3200) );
  OAI211_X1 U15289 ( .C1(n13846), .C2(n13845), .A(n13844), .B(n13881), .ZN(
        n13851) );
  OAI22_X1 U15290 ( .A1(n13898), .A2(n14237), .B1(n13868), .B2(n14235), .ZN(
        n14128) );
  INV_X1 U15291 ( .A(n14132), .ZN(n13848) );
  OAI22_X1 U15292 ( .A1(n13848), .A2(n13902), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13847), .ZN(n13849) );
  AOI21_X1 U15293 ( .B1(n14128), .B2(n13872), .A(n13849), .ZN(n13850) );
  OAI211_X1 U15294 ( .C1(n14134), .C2(n13889), .A(n13851), .B(n13850), .ZN(
        P2_U3201) );
  XNOR2_X1 U15295 ( .A(n13853), .B(n13852), .ZN(n13854) );
  XNOR2_X1 U15296 ( .A(n13855), .B(n13854), .ZN(n13862) );
  NAND2_X1 U15297 ( .A1(n13892), .A2(n14188), .ZN(n13858) );
  AOI22_X1 U15298 ( .A1(n13856), .A2(n14193), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13857) );
  OAI211_X1 U15299 ( .C1(n13859), .C2(n13867), .A(n13858), .B(n13857), .ZN(
        n13860) );
  AOI21_X1 U15300 ( .B1(n14346), .B2(n13905), .A(n13860), .ZN(n13861) );
  OAI21_X1 U15301 ( .B1(n13862), .B2(n13907), .A(n13861), .ZN(P2_U3205) );
  AOI211_X1 U15302 ( .C1(n13865), .C2(n13864), .A(n13907), .B(n13863), .ZN(
        n13866) );
  INV_X1 U15303 ( .A(n13866), .ZN(n13874) );
  OAI22_X1 U15304 ( .A1(n13868), .A2(n14237), .B1(n13867), .B2(n14235), .ZN(
        n14158) );
  INV_X1 U15305 ( .A(n14160), .ZN(n13870) );
  OAI22_X1 U15306 ( .A1(n13870), .A2(n13902), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13869), .ZN(n13871) );
  AOI21_X1 U15307 ( .B1(n14158), .B2(n13872), .A(n13871), .ZN(n13873) );
  OAI211_X1 U15308 ( .C1(n14162), .C2(n13889), .A(n13874), .B(n13873), .ZN(
        P2_U3207) );
  AOI22_X1 U15309 ( .A1(n13887), .A2(n13929), .B1(n13892), .B2(n13932), .ZN(
        n13884) );
  AOI22_X1 U15310 ( .A1(n13905), .A2(n13876), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n13875), .ZN(n13883) );
  OAI21_X1 U15311 ( .B1(n13879), .B2(n13878), .A(n13877), .ZN(n13880) );
  NAND2_X1 U15312 ( .A1(n13881), .A2(n13880), .ZN(n13882) );
  NAND3_X1 U15313 ( .A1(n13884), .A2(n13883), .A3(n13882), .ZN(P2_U3209) );
  XNOR2_X1 U15314 ( .A(n13886), .B(n13885), .ZN(n13894) );
  NAND2_X1 U15315 ( .A1(n13887), .A2(n14188), .ZN(n13888) );
  NAND2_X1 U15316 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n15498)
         );
  OAI211_X1 U15317 ( .C1(n13902), .C2(n14229), .A(n13888), .B(n15498), .ZN(
        n13891) );
  NOR2_X1 U15318 ( .A1(n14397), .A2(n13889), .ZN(n13890) );
  AOI211_X1 U15319 ( .C1(n13892), .C2(n14276), .A(n13891), .B(n13890), .ZN(
        n13893) );
  OAI21_X1 U15320 ( .B1(n13894), .B2(n13907), .A(n13893), .ZN(P2_U3210) );
  NOR2_X1 U15321 ( .A1(n13898), .A2(n14235), .ZN(n13899) );
  AOI21_X1 U15322 ( .B1(n13912), .B2(n14275), .A(n13899), .ZN(n14099) );
  NOR2_X1 U15323 ( .A1(n14099), .A2(n13900), .ZN(n13904) );
  OAI22_X1 U15324 ( .A1(n14103), .A2(n13902), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13901), .ZN(n13903) );
  AOI211_X1 U15325 ( .C1(n14314), .C2(n13905), .A(n13904), .B(n13903), .ZN(
        n13906) );
  OAI21_X1 U15326 ( .B1(n13908), .B2(n13907), .A(n13906), .ZN(P2_U3212) );
  MUX2_X1 U15327 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n14046), .S(P2_U3947), .Z(
        P2_U3562) );
  INV_X2 U15328 ( .A(P2_U3947), .ZN(n13930) );
  MUX2_X1 U15329 ( .A(n13909), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13930), .Z(
        P2_U3561) );
  MUX2_X1 U15330 ( .A(n13910), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13930), .Z(
        P2_U3560) );
  MUX2_X1 U15331 ( .A(n13911), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13930), .Z(
        P2_U3559) );
  MUX2_X1 U15332 ( .A(n13912), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13930), .Z(
        P2_U3558) );
  MUX2_X1 U15333 ( .A(n13913), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13930), .Z(
        P2_U3557) );
  MUX2_X1 U15334 ( .A(n13914), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13930), .Z(
        P2_U3556) );
  MUX2_X1 U15335 ( .A(n13915), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13930), .Z(
        P2_U3555) );
  MUX2_X1 U15336 ( .A(n13916), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13930), .Z(
        P2_U3554) );
  MUX2_X1 U15337 ( .A(n13917), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13930), .Z(
        P2_U3553) );
  MUX2_X1 U15338 ( .A(n14189), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13930), .Z(
        P2_U3552) );
  MUX2_X1 U15339 ( .A(n13918), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13930), .Z(
        P2_U3551) );
  MUX2_X1 U15340 ( .A(n14188), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13930), .Z(
        P2_U3550) );
  MUX2_X1 U15341 ( .A(n14250), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13930), .Z(
        P2_U3549) );
  MUX2_X1 U15342 ( .A(n14276), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13930), .Z(
        P2_U3548) );
  MUX2_X1 U15343 ( .A(n14249), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13930), .Z(
        P2_U3547) );
  MUX2_X1 U15344 ( .A(n14273), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13930), .Z(
        P2_U3546) );
  MUX2_X1 U15345 ( .A(n13919), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13930), .Z(
        P2_U3545) );
  MUX2_X1 U15346 ( .A(n13920), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13930), .Z(
        P2_U3543) );
  MUX2_X1 U15347 ( .A(n13921), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13930), .Z(
        P2_U3542) );
  MUX2_X1 U15348 ( .A(n13922), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13930), .Z(
        P2_U3541) );
  MUX2_X1 U15349 ( .A(n13923), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13930), .Z(
        P2_U3540) );
  MUX2_X1 U15350 ( .A(n13924), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13930), .Z(
        P2_U3539) );
  MUX2_X1 U15351 ( .A(n13925), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13930), .Z(
        P2_U3538) );
  MUX2_X1 U15352 ( .A(n13926), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13930), .Z(
        P2_U3537) );
  MUX2_X1 U15353 ( .A(n13927), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13930), .Z(
        P2_U3536) );
  MUX2_X1 U15354 ( .A(n13928), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13930), .Z(
        P2_U3535) );
  MUX2_X1 U15355 ( .A(n13929), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13930), .Z(
        P2_U3534) );
  MUX2_X1 U15356 ( .A(n13931), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13930), .Z(
        P2_U3533) );
  MUX2_X1 U15357 ( .A(n13932), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13930), .Z(
        P2_U3532) );
  INV_X1 U15358 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n13934) );
  OAI21_X1 U15359 ( .B1(n15534), .B2(n13934), .A(n13933), .ZN(n13935) );
  AOI21_X1 U15360 ( .B1(n13936), .B2(n15521), .A(n13935), .ZN(n13946) );
  MUX2_X1 U15361 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n11522), .S(n13940), .Z(
        n13938) );
  NAND3_X1 U15362 ( .A1(n13938), .A2(n15480), .A3(n13937), .ZN(n13939) );
  NAND3_X1 U15363 ( .A1(n15523), .A2(n13952), .A3(n13939), .ZN(n13945) );
  MUX2_X1 U15364 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10500), .S(n13940), .Z(
        n13942) );
  NAND3_X1 U15365 ( .A1(n13942), .A2(n15477), .A3(n13941), .ZN(n13943) );
  NAND3_X1 U15366 ( .A1(n15527), .A2(n13957), .A3(n13943), .ZN(n13944) );
  NAND3_X1 U15367 ( .A1(n13946), .A2(n13945), .A3(n13944), .ZN(P2_U3218) );
  INV_X1 U15368 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n13948) );
  OAI21_X1 U15369 ( .B1(n15534), .B2(n13948), .A(n13947), .ZN(n13949) );
  AOI21_X1 U15370 ( .B1(n13954), .B2(n15521), .A(n13949), .ZN(n13961) );
  MUX2_X1 U15371 ( .A(n11533), .B(P2_REG2_REG_5__SCAN_IN), .S(n13954), .Z(
        n13950) );
  NAND3_X1 U15372 ( .A1(n13952), .A2(n13951), .A3(n13950), .ZN(n13953) );
  NAND3_X1 U15373 ( .A1(n15523), .A2(n13972), .A3(n13953), .ZN(n13960) );
  MUX2_X1 U15374 ( .A(n10503), .B(P2_REG1_REG_5__SCAN_IN), .S(n13954), .Z(
        n13955) );
  NAND3_X1 U15375 ( .A1(n13957), .A2(n13956), .A3(n13955), .ZN(n13958) );
  NAND3_X1 U15376 ( .A1(n15527), .A2(n13967), .A3(n13958), .ZN(n13959) );
  NAND3_X1 U15377 ( .A1(n13961), .A2(n13960), .A3(n13959), .ZN(P2_U3219) );
  INV_X1 U15378 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n13963) );
  OAI21_X1 U15379 ( .B1(n15534), .B2(n13963), .A(n13962), .ZN(n13964) );
  AOI21_X1 U15380 ( .B1(n13969), .B2(n15521), .A(n13964), .ZN(n13976) );
  MUX2_X1 U15381 ( .A(n10506), .B(P2_REG1_REG_6__SCAN_IN), .S(n13969), .Z(
        n13965) );
  NAND3_X1 U15382 ( .A1(n13967), .A2(n13966), .A3(n13965), .ZN(n13968) );
  NAND3_X1 U15383 ( .A1(n15527), .A2(n13982), .A3(n13968), .ZN(n13975) );
  MUX2_X1 U15384 ( .A(n10481), .B(P2_REG2_REG_6__SCAN_IN), .S(n13969), .Z(
        n13970) );
  NAND3_X1 U15385 ( .A1(n13972), .A2(n13971), .A3(n13970), .ZN(n13973) );
  NAND3_X1 U15386 ( .A1(n15523), .A2(n13987), .A3(n13973), .ZN(n13974) );
  NAND3_X1 U15387 ( .A1(n13976), .A2(n13975), .A3(n13974), .ZN(P2_U3220) );
  INV_X1 U15388 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n13978) );
  OAI21_X1 U15389 ( .B1(n15534), .B2(n13978), .A(n13977), .ZN(n13979) );
  AOI21_X1 U15390 ( .B1(n13984), .B2(n15521), .A(n13979), .ZN(n13991) );
  MUX2_X1 U15391 ( .A(n10509), .B(P2_REG1_REG_7__SCAN_IN), .S(n13984), .Z(
        n13980) );
  NAND3_X1 U15392 ( .A1(n13982), .A2(n13981), .A3(n13980), .ZN(n13983) );
  NAND3_X1 U15393 ( .A1(n15527), .A2(n13997), .A3(n13983), .ZN(n13990) );
  MUX2_X1 U15394 ( .A(n11551), .B(P2_REG2_REG_7__SCAN_IN), .S(n13984), .Z(
        n13985) );
  NAND3_X1 U15395 ( .A1(n13987), .A2(n13986), .A3(n13985), .ZN(n13988) );
  NAND3_X1 U15396 ( .A1(n15523), .A2(n14003), .A3(n13988), .ZN(n13989) );
  NAND3_X1 U15397 ( .A1(n13991), .A2(n13990), .A3(n13989), .ZN(P2_U3221) );
  INV_X1 U15398 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n13993) );
  OAI21_X1 U15399 ( .B1(n15534), .B2(n13993), .A(n13992), .ZN(n13994) );
  AOI21_X1 U15400 ( .B1(n14000), .B2(n15521), .A(n13994), .ZN(n14008) );
  MUX2_X1 U15401 ( .A(n10512), .B(P2_REG1_REG_8__SCAN_IN), .S(n14000), .Z(
        n13995) );
  NAND3_X1 U15402 ( .A1(n13997), .A2(n13996), .A3(n13995), .ZN(n13998) );
  NAND3_X1 U15403 ( .A1(n13999), .A2(n15527), .A3(n13998), .ZN(n14007) );
  MUX2_X1 U15404 ( .A(n11400), .B(P2_REG2_REG_8__SCAN_IN), .S(n14000), .Z(
        n14001) );
  NAND3_X1 U15405 ( .A1(n14003), .A2(n14002), .A3(n14001), .ZN(n14004) );
  NAND3_X1 U15406 ( .A1(n14005), .A2(n15523), .A3(n14004), .ZN(n14006) );
  NAND3_X1 U15407 ( .A1(n14008), .A2(n14007), .A3(n14006), .ZN(P2_U3222) );
  OAI21_X1 U15408 ( .B1(n14010), .B2(n14009), .A(n15518), .ZN(n14011) );
  NAND2_X1 U15409 ( .A1(n14011), .A2(n15523), .ZN(n14023) );
  OAI21_X1 U15410 ( .B1(n15534), .B2(n7617), .A(n14012), .ZN(n14013) );
  AOI21_X1 U15411 ( .B1(n14014), .B2(n15521), .A(n14013), .ZN(n14022) );
  MUX2_X1 U15412 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n11138), .S(n14015), .Z(
        n14016) );
  NAND3_X1 U15413 ( .A1(n14018), .A2(n14017), .A3(n14016), .ZN(n14019) );
  NAND3_X1 U15414 ( .A1(n14020), .A2(n15527), .A3(n14019), .ZN(n14021) );
  NAND3_X1 U15415 ( .A1(n14023), .A2(n14022), .A3(n14021), .ZN(P2_U3225) );
  NOR2_X1 U15416 ( .A1(n14032), .A2(n14024), .ZN(n14026) );
  AOI211_X1 U15417 ( .C1(n14032), .C2(n14024), .A(n14026), .B(n14025), .ZN(
        n14029) );
  INV_X1 U15418 ( .A(n14027), .ZN(n14028) );
  OAI21_X1 U15419 ( .B1(n14029), .B2(n14028), .A(n15523), .ZN(n14041) );
  OAI21_X1 U15420 ( .B1(n15534), .B2(n7610), .A(n14030), .ZN(n14031) );
  AOI21_X1 U15421 ( .B1(n14032), .B2(n15521), .A(n14031), .ZN(n14040) );
  INV_X1 U15422 ( .A(n15508), .ZN(n14038) );
  NAND2_X1 U15423 ( .A1(n14035), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n14033) );
  OAI211_X1 U15424 ( .C1(P2_REG1_REG_14__SCAN_IN), .C2(n14035), .A(n14034), 
        .B(n14033), .ZN(n14037) );
  OAI211_X1 U15425 ( .C1(n14038), .C2(n14037), .A(n14036), .B(n15527), .ZN(
        n14039) );
  NAND3_X1 U15426 ( .A1(n14041), .A2(n14040), .A3(n14039), .ZN(P2_U3228) );
  INV_X1 U15427 ( .A(n14049), .ZN(n14042) );
  INV_X1 U15428 ( .A(n14299), .ZN(n14377) );
  NAND2_X1 U15429 ( .A1(n14042), .A2(n14377), .ZN(n14051) );
  XNOR2_X1 U15430 ( .A(n14051), .B(n14373), .ZN(n14043) );
  NAND2_X1 U15431 ( .A1(n14043), .A2(n14151), .ZN(n14294) );
  INV_X1 U15432 ( .A(n14044), .ZN(n14045) );
  NAND2_X1 U15433 ( .A1(n14046), .A2(n14045), .ZN(n14296) );
  NOR2_X1 U15434 ( .A1(n14265), .A2(n14296), .ZN(n14054) );
  NOR2_X1 U15435 ( .A1(n14373), .A2(n14288), .ZN(n14047) );
  AOI211_X1 U15436 ( .C1(P2_REG2_REG_31__SCAN_IN), .C2(n14265), .A(n14054), 
        .B(n14047), .ZN(n14048) );
  OAI21_X1 U15437 ( .B1(n14261), .B2(n14294), .A(n14048), .ZN(P2_U3234) );
  AOI21_X1 U15438 ( .B1(n14049), .B2(n14299), .A(n14282), .ZN(n14050) );
  NAND2_X1 U15439 ( .A1(n14051), .A2(n14050), .ZN(n14297) );
  NOR2_X1 U15440 ( .A1(n14280), .A2(n14052), .ZN(n14053) );
  AOI211_X1 U15441 ( .C1(n14299), .C2(n14258), .A(n14054), .B(n14053), .ZN(
        n14055) );
  OAI21_X1 U15442 ( .B1(n14297), .B2(n14261), .A(n14055), .ZN(P2_U3235) );
  NAND2_X1 U15443 ( .A1(n14056), .A2(n14280), .ZN(n14066) );
  INV_X1 U15444 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n14057) );
  OAI22_X1 U15445 ( .A1(n14058), .A2(n14255), .B1(n14057), .B2(n14280), .ZN(
        n14059) );
  AOI21_X1 U15446 ( .B1(n14060), .B2(n14258), .A(n14059), .ZN(n14065) );
  NAND2_X1 U15447 ( .A1(n14061), .A2(n14263), .ZN(n14064) );
  NAND2_X1 U15448 ( .A1(n14062), .A2(n14290), .ZN(n14063) );
  NAND4_X1 U15449 ( .A1(n14066), .A2(n14065), .A3(n14064), .A4(n14063), .ZN(
        P2_U3236) );
  AOI21_X1 U15450 ( .B1(n14089), .B2(n14305), .A(n14282), .ZN(n14068) );
  NOR2_X1 U15451 ( .A1(n14069), .A2(n14255), .ZN(n14075) );
  OAI211_X1 U15452 ( .C1(n14072), .C2(n14071), .A(n14070), .B(n14271), .ZN(
        n14074) );
  NAND2_X1 U15453 ( .A1(n14074), .A2(n14073), .ZN(n14303) );
  AOI211_X1 U15454 ( .C1(n14304), .C2(n14076), .A(n14075), .B(n14303), .ZN(
        n14082) );
  AOI22_X1 U15455 ( .A1(n14305), .A2(n14258), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n14265), .ZN(n14081) );
  OAI21_X1 U15456 ( .B1(n14079), .B2(n14078), .A(n14077), .ZN(n14302) );
  NAND2_X1 U15457 ( .A1(n14302), .A2(n14263), .ZN(n14080) );
  OAI211_X1 U15458 ( .C1(n14082), .C2(n14265), .A(n14081), .B(n14080), .ZN(
        P2_U3237) );
  XNOR2_X1 U15459 ( .A(n14083), .B(n7327), .ZN(n14085) );
  AOI21_X1 U15460 ( .B1(n14085), .B2(n14271), .A(n14084), .ZN(n14311) );
  XNOR2_X1 U15461 ( .A(n14087), .B(n14086), .ZN(n14312) );
  INV_X1 U15462 ( .A(n14312), .ZN(n14095) );
  OR2_X1 U15463 ( .A1(n14093), .A2(n14102), .ZN(n14088) );
  AND3_X1 U15464 ( .A1(n14089), .A2(n14151), .A3(n14088), .ZN(n14308) );
  NAND2_X1 U15465 ( .A1(n14308), .A2(n14290), .ZN(n14092) );
  AOI22_X1 U15466 ( .A1(n14090), .A2(n14285), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n14265), .ZN(n14091) );
  OAI211_X1 U15467 ( .C1(n14093), .C2(n14288), .A(n14092), .B(n14091), .ZN(
        n14094) );
  AOI21_X1 U15468 ( .B1(n14095), .B2(n14263), .A(n14094), .ZN(n14096) );
  OAI21_X1 U15469 ( .B1(n14311), .B2(n14265), .A(n14096), .ZN(P2_U3238) );
  XNOR2_X1 U15470 ( .A(n14098), .B(n14097), .ZN(n14101) );
  INV_X1 U15471 ( .A(n14099), .ZN(n14100) );
  AOI21_X1 U15472 ( .B1(n14101), .B2(n14271), .A(n14100), .ZN(n14319) );
  AOI211_X1 U15473 ( .C1(n14314), .C2(n14117), .A(n14282), .B(n14102), .ZN(
        n14313) );
  INV_X1 U15474 ( .A(n14103), .ZN(n14104) );
  AOI22_X1 U15475 ( .A1(n14104), .A2(n14285), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14265), .ZN(n14105) );
  OAI21_X1 U15476 ( .B1(n14106), .B2(n14288), .A(n14105), .ZN(n14107) );
  AOI21_X1 U15477 ( .B1(n14313), .B2(n14290), .A(n14107), .ZN(n14110) );
  NAND2_X1 U15478 ( .A1(n14108), .A2(n7483), .ZN(n14315) );
  NAND3_X1 U15479 ( .A1(n14316), .A2(n14315), .A3(n14263), .ZN(n14109) );
  OAI211_X1 U15480 ( .C1(n14319), .C2(n14265), .A(n14110), .B(n14109), .ZN(
        P2_U3239) );
  XNOR2_X1 U15481 ( .A(n14111), .B(n14116), .ZN(n14114) );
  INV_X1 U15482 ( .A(n14112), .ZN(n14113) );
  OAI21_X1 U15483 ( .B1(n14114), .B2(n14243), .A(n14113), .ZN(n14320) );
  INV_X1 U15484 ( .A(n14320), .ZN(n14125) );
  OAI21_X1 U15485 ( .B1(n7217), .B2(n14116), .A(n14115), .ZN(n14322) );
  INV_X1 U15486 ( .A(n14117), .ZN(n14118) );
  AOI211_X1 U15487 ( .C1(n14119), .C2(n14130), .A(n14282), .B(n14118), .ZN(
        n14321) );
  NAND2_X1 U15488 ( .A1(n14321), .A2(n14290), .ZN(n14122) );
  AOI22_X1 U15489 ( .A1(n14120), .A2(n14285), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n14265), .ZN(n14121) );
  OAI211_X1 U15490 ( .C1(n14384), .C2(n14288), .A(n14122), .B(n14121), .ZN(
        n14123) );
  AOI21_X1 U15491 ( .B1(n14263), .B2(n14322), .A(n14123), .ZN(n14124) );
  OAI21_X1 U15492 ( .B1(n14125), .B2(n14265), .A(n14124), .ZN(P2_U3240) );
  OAI21_X1 U15493 ( .B1(n7212), .B2(n14127), .A(n14126), .ZN(n14129) );
  AOI21_X1 U15494 ( .B1(n14129), .B2(n14271), .A(n14128), .ZN(n14328) );
  AOI21_X1 U15495 ( .B1(n14152), .B2(n14326), .A(n14282), .ZN(n14131) );
  AND2_X1 U15496 ( .A1(n14131), .A2(n14130), .ZN(n14325) );
  AOI22_X1 U15497 ( .A1(n14132), .A2(n14285), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n14265), .ZN(n14133) );
  OAI21_X1 U15498 ( .B1(n14134), .B2(n14288), .A(n14133), .ZN(n14138) );
  OAI21_X1 U15499 ( .B1(n14136), .B2(n8034), .A(n14135), .ZN(n14329) );
  NOR2_X1 U15500 ( .A1(n14329), .A2(n14198), .ZN(n14137) );
  AOI211_X1 U15501 ( .C1(n14325), .C2(n14290), .A(n14138), .B(n14137), .ZN(
        n14139) );
  OAI21_X1 U15502 ( .B1(n14328), .B2(n14265), .A(n14139), .ZN(P2_U3241) );
  AOI211_X1 U15503 ( .C1(n7200), .C2(n14141), .A(n14243), .B(n14140), .ZN(
        n14143) );
  NOR2_X1 U15504 ( .A1(n14143), .A2(n14142), .ZN(n14333) );
  OAI21_X1 U15505 ( .B1(n7200), .B2(n14145), .A(n14144), .ZN(n14334) );
  INV_X1 U15506 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n14146) );
  OAI22_X1 U15507 ( .A1(n14147), .A2(n14255), .B1(n14146), .B2(n14280), .ZN(
        n14148) );
  AOI21_X1 U15508 ( .B1(n14331), .B2(n14258), .A(n14148), .ZN(n14154) );
  OR2_X1 U15509 ( .A1(n7180), .A2(n14149), .ZN(n14150) );
  AND3_X1 U15510 ( .A1(n14152), .A2(n14151), .A3(n14150), .ZN(n14330) );
  NAND2_X1 U15511 ( .A1(n14330), .A2(n14290), .ZN(n14153) );
  OAI211_X1 U15512 ( .C1(n14334), .C2(n14198), .A(n14154), .B(n14153), .ZN(
        n14155) );
  INV_X1 U15513 ( .A(n14155), .ZN(n14156) );
  OAI21_X1 U15514 ( .B1(n14333), .B2(n14265), .A(n14156), .ZN(P2_U3242) );
  XOR2_X1 U15515 ( .A(n14157), .B(n14164), .Z(n14159) );
  AOI21_X1 U15516 ( .B1(n14159), .B2(n14271), .A(n14158), .ZN(n14337) );
  AOI211_X1 U15517 ( .C1(n14336), .C2(n7589), .A(n8098), .B(n7180), .ZN(n14335) );
  AOI22_X1 U15518 ( .A1(n14160), .A2(n14285), .B1(P2_REG2_REG_22__SCAN_IN), 
        .B2(n14265), .ZN(n14161) );
  OAI21_X1 U15519 ( .B1(n14162), .B2(n14288), .A(n14161), .ZN(n14168) );
  OR2_X1 U15520 ( .A1(n14164), .A2(n14163), .ZN(n14165) );
  NAND2_X1 U15521 ( .A1(n14166), .A2(n14165), .ZN(n14339) );
  NOR2_X1 U15522 ( .A1(n14339), .A2(n14198), .ZN(n14167) );
  AOI211_X1 U15523 ( .C1(n14335), .C2(n14290), .A(n14168), .B(n14167), .ZN(
        n14169) );
  OAI21_X1 U15524 ( .B1(n14265), .B2(n14337), .A(n14169), .ZN(P2_U3243) );
  OAI211_X1 U15525 ( .C1(n14175), .C2(n14171), .A(n14170), .B(n14271), .ZN(
        n14173) );
  AND2_X1 U15526 ( .A1(n14173), .A2(n14172), .ZN(n14343) );
  NAND2_X1 U15527 ( .A1(n14175), .A2(n14174), .ZN(n14176) );
  AND2_X1 U15528 ( .A1(n14177), .A2(n14176), .ZN(n14340) );
  AND2_X1 U15529 ( .A1(n14182), .A2(n14191), .ZN(n14179) );
  OR3_X1 U15530 ( .A1(n14179), .A2(n14178), .A3(n8098), .ZN(n14341) );
  INV_X1 U15531 ( .A(n14180), .ZN(n14181) );
  AOI22_X1 U15532 ( .A1(n14181), .A2(n14285), .B1(P2_REG2_REG_21__SCAN_IN), 
        .B2(n14265), .ZN(n14184) );
  NAND2_X1 U15533 ( .A1(n14182), .A2(n14258), .ZN(n14183) );
  OAI211_X1 U15534 ( .C1(n14341), .C2(n14261), .A(n14184), .B(n14183), .ZN(
        n14185) );
  AOI21_X1 U15535 ( .B1(n14263), .B2(n14340), .A(n14185), .ZN(n14186) );
  OAI21_X1 U15536 ( .B1(n14265), .B2(n14343), .A(n14186), .ZN(P2_U3244) );
  XNOR2_X1 U15537 ( .A(n14197), .B(n14187), .ZN(n14190) );
  AOI222_X1 U15538 ( .A1(n14271), .A2(n14190), .B1(n14189), .B2(n14275), .C1(
        n14188), .C2(n14274), .ZN(n14350) );
  OR2_X1 U15539 ( .A1(n14195), .A2(n14216), .ZN(n14192) );
  AND2_X1 U15540 ( .A1(n14192), .A2(n14191), .ZN(n14349) );
  AOI22_X1 U15541 ( .A1(P2_REG2_REG_20__SCAN_IN), .A2(n14265), .B1(n14193), 
        .B2(n14285), .ZN(n14194) );
  OAI21_X1 U15542 ( .B1(n14195), .B2(n14288), .A(n14194), .ZN(n14200) );
  XNOR2_X1 U15543 ( .A(n14197), .B(n14196), .ZN(n14352) );
  NOR2_X1 U15544 ( .A1(n14352), .A2(n14198), .ZN(n14199) );
  AOI211_X1 U15545 ( .C1(n14349), .C2(n14201), .A(n14200), .B(n14199), .ZN(
        n14202) );
  OAI21_X1 U15546 ( .B1(n14265), .B2(n14350), .A(n14202), .ZN(P2_U3245) );
  OR2_X1 U15547 ( .A1(n14203), .A2(n14206), .ZN(n14204) );
  NAND2_X1 U15548 ( .A1(n14205), .A2(n14204), .ZN(n14357) );
  INV_X1 U15549 ( .A(n14279), .ZN(n14240) );
  NAND2_X1 U15550 ( .A1(n14357), .A2(n14240), .ZN(n14214) );
  XNOR2_X1 U15551 ( .A(n14207), .B(n14206), .ZN(n14208) );
  NAND2_X1 U15552 ( .A1(n14208), .A2(n14271), .ZN(n14213) );
  OAI22_X1 U15553 ( .A1(n14210), .A2(n14237), .B1(n14209), .B2(n14235), .ZN(
        n14211) );
  INV_X1 U15554 ( .A(n14211), .ZN(n14212) );
  INV_X1 U15555 ( .A(n14293), .ZN(n14223) );
  OAI21_X1 U15556 ( .B1(n14355), .B2(n14227), .A(n14348), .ZN(n14215) );
  OR2_X1 U15557 ( .A1(n14216), .A2(n14215), .ZN(n14354) );
  OAI22_X1 U15558 ( .A1(n14280), .A2(n14218), .B1(n14217), .B2(n14255), .ZN(
        n14219) );
  AOI21_X1 U15559 ( .B1(n14220), .B2(n14258), .A(n14219), .ZN(n14221) );
  OAI21_X1 U15560 ( .B1(n14354), .B2(n14261), .A(n14221), .ZN(n14222) );
  AOI21_X1 U15561 ( .B1(n14223), .B2(n14357), .A(n14222), .ZN(n14224) );
  OAI21_X1 U15562 ( .B1(n14359), .B2(n14265), .A(n14224), .ZN(P2_U3246) );
  OAI21_X1 U15563 ( .B1(n14233), .B2(n14226), .A(n14225), .ZN(n14362) );
  INV_X1 U15564 ( .A(n14362), .ZN(n14246) );
  AOI211_X1 U15565 ( .C1(n14228), .C2(n14254), .A(n14282), .B(n14227), .ZN(
        n14361) );
  INV_X1 U15566 ( .A(n14229), .ZN(n14230) );
  AOI22_X1 U15567 ( .A1(n14265), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14230), 
        .B2(n14285), .ZN(n14231) );
  OAI21_X1 U15568 ( .B1(n14397), .B2(n14288), .A(n14231), .ZN(n14232) );
  AOI21_X1 U15569 ( .B1(n14361), .B2(n14290), .A(n14232), .ZN(n14245) );
  XNOR2_X1 U15570 ( .A(n14234), .B(n14233), .ZN(n14242) );
  OAI22_X1 U15571 ( .A1(n14238), .A2(n14237), .B1(n14236), .B2(n14235), .ZN(
        n14239) );
  AOI21_X1 U15572 ( .B1(n14362), .B2(n14240), .A(n14239), .ZN(n14241) );
  OAI21_X1 U15573 ( .B1(n14243), .B2(n14242), .A(n14241), .ZN(n14360) );
  NAND2_X1 U15574 ( .A1(n14360), .A2(n14280), .ZN(n14244) );
  OAI211_X1 U15575 ( .C1(n14246), .C2(n14293), .A(n14245), .B(n14244), .ZN(
        P2_U3247) );
  XNOR2_X1 U15576 ( .A(n14248), .B(n14247), .ZN(n14251) );
  AOI222_X1 U15577 ( .A1(n14271), .A2(n14251), .B1(n14250), .B2(n14275), .C1(
        n14249), .C2(n14274), .ZN(n16028) );
  XNOR2_X1 U15578 ( .A(n14253), .B(n14252), .ZN(n16032) );
  OAI211_X1 U15579 ( .C1(n16030), .C2(n14281), .A(n14348), .B(n14254), .ZN(
        n16027) );
  OAI22_X1 U15580 ( .A1(n14280), .A2(n12082), .B1(n14256), .B2(n14255), .ZN(
        n14257) );
  AOI21_X1 U15581 ( .B1(n14259), .B2(n14258), .A(n14257), .ZN(n14260) );
  OAI21_X1 U15582 ( .B1(n16027), .B2(n14261), .A(n14260), .ZN(n14262) );
  AOI21_X1 U15583 ( .B1(n16032), .B2(n14263), .A(n14262), .ZN(n14264) );
  OAI21_X1 U15584 ( .B1(n16028), .B2(n14265), .A(n14264), .ZN(P2_U3248) );
  NAND2_X1 U15585 ( .A1(n14266), .A2(n14270), .ZN(n14267) );
  NAND2_X1 U15586 ( .A1(n14268), .A2(n14267), .ZN(n14364) );
  XOR2_X1 U15587 ( .A(n14270), .B(n14269), .Z(n14272) );
  NAND2_X1 U15588 ( .A1(n14272), .A2(n14271), .ZN(n14278) );
  AOI22_X1 U15589 ( .A1(n14276), .A2(n14275), .B1(n14274), .B2(n14273), .ZN(
        n14277) );
  OAI211_X1 U15590 ( .C1(n14364), .C2(n14279), .A(n14278), .B(n14277), .ZN(
        n14365) );
  NAND2_X1 U15591 ( .A1(n14365), .A2(n14280), .ZN(n14292) );
  AOI211_X1 U15592 ( .C1(n14284), .C2(n14283), .A(n14282), .B(n14281), .ZN(
        n14366) );
  AOI22_X1 U15593 ( .A1(n14265), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n14286), 
        .B2(n14285), .ZN(n14287) );
  OAI21_X1 U15594 ( .B1(n14403), .B2(n14288), .A(n14287), .ZN(n14289) );
  AOI21_X1 U15595 ( .B1(n14366), .B2(n14290), .A(n14289), .ZN(n14291) );
  OAI211_X1 U15596 ( .C1(n14364), .C2(n14293), .A(n14292), .B(n14291), .ZN(
        P2_U3249) );
  NAND2_X1 U15597 ( .A1(n14297), .A2(n14296), .ZN(n14374) );
  MUX2_X1 U15598 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n14374), .S(n16035), .Z(
        n14298) );
  AOI21_X1 U15599 ( .B1(n14300), .B2(n14299), .A(n14298), .ZN(n14301) );
  INV_X1 U15600 ( .A(n14301), .ZN(P2_U3529) );
  INV_X1 U15601 ( .A(n14302), .ZN(n14307) );
  OAI21_X1 U15602 ( .B1(n14353), .B2(n14307), .A(n14306), .ZN(n14378) );
  MUX2_X1 U15603 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n14378), .S(n16035), .Z(
        P2_U3527) );
  AOI21_X1 U15604 ( .B1(n14347), .B2(n14309), .A(n14308), .ZN(n14310) );
  OAI211_X1 U15605 ( .C1(n14353), .C2(n14312), .A(n14311), .B(n14310), .ZN(
        n14379) );
  MUX2_X1 U15606 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n14379), .S(n16035), .Z(
        P2_U3526) );
  AOI21_X1 U15607 ( .B1(n14347), .B2(n14314), .A(n14313), .ZN(n14318) );
  NAND3_X1 U15608 ( .A1(n14316), .A2(n14315), .A3(n16033), .ZN(n14317) );
  NAND3_X1 U15609 ( .A1(n14319), .A2(n14318), .A3(n14317), .ZN(n14380) );
  MUX2_X1 U15610 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14380), .S(n16035), .Z(
        P2_U3525) );
  AOI211_X1 U15611 ( .C1(n16033), .C2(n14322), .A(n14321), .B(n14320), .ZN(
        n14381) );
  MUX2_X1 U15612 ( .A(n14323), .B(n14381), .S(n16035), .Z(n14324) );
  OAI21_X1 U15613 ( .B1(n14384), .B2(n14369), .A(n14324), .ZN(P2_U3524) );
  AOI21_X1 U15614 ( .B1(n14347), .B2(n14326), .A(n14325), .ZN(n14327) );
  OAI211_X1 U15615 ( .C1(n14353), .C2(n14329), .A(n14328), .B(n14327), .ZN(
        n14385) );
  MUX2_X1 U15616 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14385), .S(n16035), .Z(
        P2_U3523) );
  AOI21_X1 U15617 ( .B1(n14347), .B2(n14331), .A(n14330), .ZN(n14332) );
  OAI211_X1 U15618 ( .C1(n14353), .C2(n14334), .A(n14333), .B(n14332), .ZN(
        n14386) );
  MUX2_X1 U15619 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14386), .S(n16035), .Z(
        P2_U3522) );
  AOI21_X1 U15620 ( .B1(n14347), .B2(n14336), .A(n14335), .ZN(n14338) );
  OAI211_X1 U15621 ( .C1(n14353), .C2(n14339), .A(n14338), .B(n14337), .ZN(
        n14387) );
  MUX2_X1 U15622 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14387), .S(n16035), .Z(
        P2_U3521) );
  NAND2_X1 U15623 ( .A1(n14340), .A2(n16033), .ZN(n14342) );
  AND3_X1 U15624 ( .A1(n14343), .A2(n14342), .A3(n14341), .ZN(n14389) );
  MUX2_X1 U15625 ( .A(n14389), .B(n14344), .S(n16034), .Z(n14345) );
  OAI21_X1 U15626 ( .B1(n14391), .B2(n14369), .A(n14345), .ZN(P2_U3520) );
  AOI22_X1 U15627 ( .A1(n14349), .A2(n14348), .B1(n14347), .B2(n14346), .ZN(
        n14351) );
  OAI211_X1 U15628 ( .C1(n14353), .C2(n14352), .A(n14351), .B(n14350), .ZN(
        n14392) );
  MUX2_X1 U15629 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14392), .S(n16035), .Z(
        P2_U3519) );
  OAI21_X1 U15630 ( .B1(n14355), .B2(n16029), .A(n14354), .ZN(n14356) );
  AOI21_X1 U15631 ( .B1(n16024), .B2(n14357), .A(n14356), .ZN(n14358) );
  NAND2_X1 U15632 ( .A1(n14359), .A2(n14358), .ZN(n14393) );
  MUX2_X1 U15633 ( .A(n14393), .B(P2_REG1_REG_19__SCAN_IN), .S(n16034), .Z(
        P2_U3518) );
  AOI211_X1 U15634 ( .C1(n16024), .C2(n14362), .A(n14361), .B(n14360), .ZN(
        n14394) );
  MUX2_X1 U15635 ( .A(n15490), .B(n14394), .S(n16035), .Z(n14363) );
  OAI21_X1 U15636 ( .B1(n14397), .B2(n14369), .A(n14363), .ZN(P2_U3517) );
  INV_X1 U15637 ( .A(n14364), .ZN(n14367) );
  AOI211_X1 U15638 ( .C1(n14367), .C2(n16024), .A(n14366), .B(n14365), .ZN(
        n14399) );
  MUX2_X1 U15639 ( .A(n11616), .B(n14399), .S(n16035), .Z(n14368) );
  OAI21_X1 U15640 ( .B1(n14403), .B2(n14369), .A(n14368), .ZN(P2_U3515) );
  MUX2_X1 U15641 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n14370), .S(n16035), .Z(
        P2_U3499) );
  MUX2_X1 U15642 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n14374), .S(n14398), .Z(
        n14375) );
  INV_X1 U15643 ( .A(n14375), .ZN(n14376) );
  OAI21_X1 U15644 ( .B1(n14377), .B2(n14402), .A(n14376), .ZN(P2_U3497) );
  MUX2_X1 U15645 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n14378), .S(n14398), .Z(
        P2_U3495) );
  MUX2_X1 U15646 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n14379), .S(n14398), .Z(
        P2_U3494) );
  MUX2_X1 U15647 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14380), .S(n14398), .Z(
        P2_U3493) );
  INV_X1 U15648 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n14382) );
  MUX2_X1 U15649 ( .A(n14382), .B(n14381), .S(n14398), .Z(n14383) );
  OAI21_X1 U15650 ( .B1(n14384), .B2(n14402), .A(n14383), .ZN(P2_U3492) );
  MUX2_X1 U15651 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14385), .S(n14398), .Z(
        P2_U3491) );
  MUX2_X1 U15652 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14386), .S(n14398), .Z(
        P2_U3490) );
  MUX2_X1 U15653 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14387), .S(n14398), .Z(
        P2_U3489) );
  INV_X1 U15654 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n14388) );
  MUX2_X1 U15655 ( .A(n14389), .B(n14388), .S(n16001), .Z(n14390) );
  OAI21_X1 U15656 ( .B1(n14391), .B2(n14402), .A(n14390), .ZN(P2_U3488) );
  MUX2_X1 U15657 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14392), .S(n14398), .Z(
        P2_U3487) );
  MUX2_X1 U15658 ( .A(n14393), .B(P2_REG0_REG_19__SCAN_IN), .S(n16001), .Z(
        P2_U3486) );
  INV_X1 U15659 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n14395) );
  MUX2_X1 U15660 ( .A(n14395), .B(n14394), .S(n14398), .Z(n14396) );
  OAI21_X1 U15661 ( .B1(n14397), .B2(n14402), .A(n14396), .ZN(P2_U3484) );
  INV_X1 U15662 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n14400) );
  MUX2_X1 U15663 ( .A(n14400), .B(n14399), .S(n14398), .Z(n14401) );
  OAI21_X1 U15664 ( .B1(n14403), .B2(n14402), .A(n14401), .ZN(P2_U3478) );
  OAI222_X1 U15665 ( .A1(n14416), .A2(n14406), .B1(P2_U3088), .B2(n14405), 
        .C1(n14404), .C2(n14422), .ZN(P2_U3298) );
  NAND2_X1 U15666 ( .A1(n15428), .A2(n14419), .ZN(n14408) );
  OAI211_X1 U15667 ( .C1(n14422), .C2(n14409), .A(n14408), .B(n14407), .ZN(
        P2_U3299) );
  INV_X1 U15668 ( .A(n14410), .ZN(n15433) );
  OAI222_X1 U15669 ( .A1(n14422), .A2(n14413), .B1(n14416), .B2(n15433), .C1(
        P2_U3088), .C2(n14411), .ZN(P2_U3300) );
  INV_X1 U15670 ( .A(n14414), .ZN(n15436) );
  OAI222_X1 U15671 ( .A1(P2_U3088), .A2(n14417), .B1(n14416), .B2(n15436), 
        .C1(n14415), .C2(n14422), .ZN(P2_U3301) );
  NAND2_X1 U15672 ( .A1(n14418), .A2(n14419), .ZN(n14421) );
  OAI211_X1 U15673 ( .C1(n14423), .C2(n14422), .A(n14421), .B(n14420), .ZN(
        P2_U3304) );
  MUX2_X1 U15674 ( .A(n14424), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  INV_X1 U15675 ( .A(n14870), .ZN(n15387) );
  NAND2_X1 U15676 ( .A1(n14870), .A2(n14532), .ZN(n14426) );
  NAND2_X1 U15677 ( .A1(n14442), .A2(n14716), .ZN(n14425) );
  NAND2_X1 U15678 ( .A1(n14426), .A2(n14425), .ZN(n14427) );
  XNOR2_X1 U15679 ( .A(n14427), .B(n14586), .ZN(n14431) );
  NAND2_X1 U15680 ( .A1(n14870), .A2(n14509), .ZN(n14429) );
  NAND2_X1 U15681 ( .A1(n14537), .A2(n14716), .ZN(n14428) );
  NAND2_X1 U15682 ( .A1(n14429), .A2(n14428), .ZN(n14430) );
  NOR2_X1 U15683 ( .A1(n14431), .A2(n14430), .ZN(n14582) );
  AOI21_X1 U15684 ( .B1(n14431), .B2(n14430), .A(n14582), .ZN(n14545) );
  OAI22_X1 U15685 ( .A1(n14686), .A2(n14590), .B1(n14432), .B2(n14588), .ZN(
        n14478) );
  NAND2_X1 U15686 ( .A1(n15407), .A2(n14532), .ZN(n14434) );
  NAND2_X1 U15687 ( .A1(n14725), .A2(n14442), .ZN(n14433) );
  NAND2_X1 U15688 ( .A1(n14434), .A2(n14433), .ZN(n14435) );
  XNOR2_X1 U15689 ( .A(n14435), .B(n14586), .ZN(n14477) );
  INV_X1 U15690 ( .A(n14438), .ZN(n14439) );
  NAND2_X1 U15691 ( .A1(n14440), .A2(n14439), .ZN(n14441) );
  NAND2_X1 U15692 ( .A1(n14561), .A2(n14532), .ZN(n14444) );
  NAND2_X1 U15693 ( .A1(n14442), .A2(n14730), .ZN(n14443) );
  NAND2_X1 U15694 ( .A1(n14444), .A2(n14443), .ZN(n14445) );
  XNOR2_X1 U15695 ( .A(n14445), .B(n14522), .ZN(n14448) );
  NOR2_X1 U15696 ( .A1(n14588), .A2(n14446), .ZN(n14447) );
  AOI21_X1 U15697 ( .B1(n14561), .B2(n14509), .A(n14447), .ZN(n14449) );
  NAND2_X1 U15698 ( .A1(n14448), .A2(n14449), .ZN(n14453) );
  INV_X1 U15699 ( .A(n14448), .ZN(n14451) );
  INV_X1 U15700 ( .A(n14449), .ZN(n14450) );
  NAND2_X1 U15701 ( .A1(n14451), .A2(n14450), .ZN(n14452) );
  NAND2_X1 U15702 ( .A1(n14453), .A2(n14452), .ZN(n14556) );
  OAI22_X1 U15703 ( .A1(n15050), .A2(n14585), .B1(n14455), .B2(n14590), .ZN(
        n14454) );
  XNOR2_X1 U15704 ( .A(n14454), .B(n14586), .ZN(n14457) );
  OAI22_X1 U15705 ( .A1(n15050), .A2(n14590), .B1(n14455), .B2(n14588), .ZN(
        n14699) );
  INV_X1 U15706 ( .A(n14456), .ZN(n14458) );
  NAND2_X1 U15707 ( .A1(n15150), .A2(n14492), .ZN(n14460) );
  NAND2_X1 U15708 ( .A1(n14728), .A2(n14509), .ZN(n14459) );
  NAND2_X1 U15709 ( .A1(n14460), .A2(n14459), .ZN(n14461) );
  XNOR2_X1 U15710 ( .A(n14461), .B(n14586), .ZN(n14465) );
  NAND2_X1 U15711 ( .A1(n15150), .A2(n14509), .ZN(n14463) );
  NAND2_X1 U15712 ( .A1(n14728), .A2(n14537), .ZN(n14462) );
  NAND2_X1 U15713 ( .A1(n14463), .A2(n14462), .ZN(n14464) );
  NOR2_X1 U15714 ( .A1(n14465), .A2(n14464), .ZN(n14466) );
  AOI21_X1 U15715 ( .B1(n14465), .B2(n14464), .A(n14466), .ZN(n14628) );
  NAND2_X1 U15716 ( .A1(n14627), .A2(n14628), .ZN(n14626) );
  INV_X1 U15717 ( .A(n14466), .ZN(n14467) );
  NAND2_X1 U15718 ( .A1(n14626), .A2(n14467), .ZN(n14635) );
  NAND2_X1 U15719 ( .A1(n15142), .A2(n14532), .ZN(n14469) );
  NAND2_X1 U15720 ( .A1(n14726), .A2(n14509), .ZN(n14468) );
  NAND2_X1 U15721 ( .A1(n14469), .A2(n14468), .ZN(n14470) );
  XNOR2_X1 U15722 ( .A(n14470), .B(n14586), .ZN(n14473) );
  NAND2_X1 U15723 ( .A1(n15142), .A2(n14509), .ZN(n14472) );
  NAND2_X1 U15724 ( .A1(n14726), .A2(n14537), .ZN(n14471) );
  NAND2_X1 U15725 ( .A1(n14472), .A2(n14471), .ZN(n14474) );
  NAND2_X1 U15726 ( .A1(n14473), .A2(n14474), .ZN(n14636) );
  INV_X1 U15727 ( .A(n14473), .ZN(n14476) );
  INV_X1 U15728 ( .A(n14474), .ZN(n14475) );
  NAND2_X1 U15729 ( .A1(n14476), .A2(n14475), .ZN(n14638) );
  XOR2_X1 U15730 ( .A(n14478), .B(n14477), .Z(n14678) );
  NAND2_X1 U15731 ( .A1(n14980), .A2(n14532), .ZN(n14480) );
  NAND2_X1 U15732 ( .A1(n14724), .A2(n14509), .ZN(n14479) );
  NAND2_X1 U15733 ( .A1(n14480), .A2(n14479), .ZN(n14481) );
  XNOR2_X1 U15734 ( .A(n14481), .B(n14586), .ZN(n14574) );
  NAND2_X1 U15735 ( .A1(n14980), .A2(n14509), .ZN(n14483) );
  NAND2_X1 U15736 ( .A1(n14724), .A2(n14537), .ZN(n14482) );
  NAND2_X1 U15737 ( .A1(n14483), .A2(n14482), .ZN(n14573) );
  NOR2_X1 U15738 ( .A1(n14574), .A2(n14573), .ZN(n14486) );
  INV_X1 U15739 ( .A(n14574), .ZN(n14485) );
  INV_X1 U15740 ( .A(n14573), .ZN(n14484) );
  OAI22_X1 U15741 ( .A1(n15403), .A2(n14585), .B1(n14606), .B2(n14590), .ZN(
        n14487) );
  XNOR2_X1 U15742 ( .A(n14487), .B(n14586), .ZN(n14490) );
  AND2_X1 U15743 ( .A1(n14723), .A2(n14537), .ZN(n14488) );
  AOI21_X1 U15744 ( .B1(n14967), .B2(n14442), .A(n14488), .ZN(n14489) );
  XNOR2_X1 U15745 ( .A(n14490), .B(n14489), .ZN(n14655) );
  INV_X1 U15746 ( .A(n14489), .ZN(n14491) );
  AOI22_X1 U15747 ( .A1(n15115), .A2(n14509), .B1(n14537), .B2(n14722), .ZN(
        n14497) );
  AOI22_X1 U15748 ( .A1(n15115), .A2(n14492), .B1(n14509), .B2(n14722), .ZN(
        n14493) );
  XNOR2_X1 U15749 ( .A(n14493), .B(n14586), .ZN(n14498) );
  XOR2_X1 U15750 ( .A(n14497), .B(n14498), .Z(n14603) );
  OR2_X1 U15751 ( .A1(n15108), .A2(n14590), .ZN(n14495) );
  NAND2_X1 U15752 ( .A1(n14721), .A2(n14537), .ZN(n14494) );
  NAND2_X1 U15753 ( .A1(n14495), .A2(n14494), .ZN(n14506) );
  OAI22_X1 U15754 ( .A1(n15108), .A2(n14585), .B1(n14608), .B2(n14590), .ZN(
        n14496) );
  XNOR2_X1 U15755 ( .A(n14496), .B(n14586), .ZN(n14507) );
  XOR2_X1 U15756 ( .A(n14506), .B(n14507), .Z(n14664) );
  NAND2_X1 U15757 ( .A1(n14498), .A2(n14497), .ZN(n14665) );
  NAND2_X1 U15758 ( .A1(n15100), .A2(n14532), .ZN(n14500) );
  NAND2_X1 U15759 ( .A1(n14509), .A2(n14720), .ZN(n14499) );
  NAND2_X1 U15760 ( .A1(n14500), .A2(n14499), .ZN(n14501) );
  XNOR2_X1 U15761 ( .A(n14501), .B(n14586), .ZN(n14505) );
  NAND2_X1 U15762 ( .A1(n15100), .A2(n14509), .ZN(n14503) );
  NAND2_X1 U15763 ( .A1(n14537), .A2(n14720), .ZN(n14502) );
  NAND2_X1 U15764 ( .A1(n14503), .A2(n14502), .ZN(n14504) );
  NOR2_X1 U15765 ( .A1(n14505), .A2(n14504), .ZN(n14508) );
  AOI21_X1 U15766 ( .B1(n14505), .B2(n14504), .A(n14508), .ZN(n14564) );
  NAND2_X1 U15767 ( .A1(n14507), .A2(n14506), .ZN(n14565) );
  INV_X1 U15768 ( .A(n14508), .ZN(n14646) );
  NAND2_X1 U15769 ( .A1(n14905), .A2(n14532), .ZN(n14511) );
  NAND2_X1 U15770 ( .A1(n14509), .A2(n14719), .ZN(n14510) );
  NAND2_X1 U15771 ( .A1(n14511), .A2(n14510), .ZN(n14512) );
  XNOR2_X1 U15772 ( .A(n14512), .B(n14522), .ZN(n14514) );
  NOR2_X1 U15773 ( .A1(n14588), .A2(n14568), .ZN(n14513) );
  AOI21_X1 U15774 ( .B1(n14905), .B2(n14509), .A(n14513), .ZN(n14515) );
  NAND2_X1 U15775 ( .A1(n14514), .A2(n14515), .ZN(n14519) );
  INV_X1 U15776 ( .A(n14514), .ZN(n14517) );
  INV_X1 U15777 ( .A(n14515), .ZN(n14516) );
  NAND2_X1 U15778 ( .A1(n14517), .A2(n14516), .ZN(n14518) );
  NAND2_X1 U15779 ( .A1(n14519), .A2(n14518), .ZN(n14645) );
  INV_X1 U15780 ( .A(n14519), .ZN(n14616) );
  NAND2_X1 U15781 ( .A1(n14897), .A2(n14532), .ZN(n14521) );
  NAND2_X1 U15782 ( .A1(n14533), .A2(n14718), .ZN(n14520) );
  NAND2_X1 U15783 ( .A1(n14521), .A2(n14520), .ZN(n14523) );
  XNOR2_X1 U15784 ( .A(n14523), .B(n14522), .ZN(n14526) );
  NOR2_X1 U15785 ( .A1(n14588), .A2(n14524), .ZN(n14525) );
  AOI21_X1 U15786 ( .B1(n14897), .B2(n14442), .A(n14525), .ZN(n14527) );
  NAND2_X1 U15787 ( .A1(n14526), .A2(n14527), .ZN(n14531) );
  INV_X1 U15788 ( .A(n14526), .ZN(n14529) );
  INV_X1 U15789 ( .A(n14527), .ZN(n14528) );
  NAND2_X1 U15790 ( .A1(n14529), .A2(n14528), .ZN(n14530) );
  AND2_X1 U15791 ( .A1(n14531), .A2(n14530), .ZN(n14615) );
  NAND2_X1 U15792 ( .A1(n15079), .A2(n14532), .ZN(n14535) );
  NAND2_X1 U15793 ( .A1(n14533), .A2(n14717), .ZN(n14534) );
  NAND2_X1 U15794 ( .A1(n14535), .A2(n14534), .ZN(n14536) );
  XNOR2_X1 U15795 ( .A(n14536), .B(n14586), .ZN(n14541) );
  NAND2_X1 U15796 ( .A1(n15079), .A2(n14509), .ZN(n14539) );
  NAND2_X1 U15797 ( .A1(n14537), .A2(n14717), .ZN(n14538) );
  NAND2_X1 U15798 ( .A1(n14539), .A2(n14538), .ZN(n14540) );
  NOR2_X1 U15799 ( .A1(n14541), .A2(n14540), .ZN(n14542) );
  AOI21_X1 U15800 ( .B1(n14541), .B2(n14540), .A(n14542), .ZN(n14689) );
  NAND2_X1 U15801 ( .A1(n14688), .A2(n14689), .ZN(n14687) );
  INV_X1 U15802 ( .A(n14542), .ZN(n14543) );
  NAND2_X1 U15803 ( .A1(n14687), .A2(n14543), .ZN(n14544) );
  NAND2_X1 U15804 ( .A1(n14544), .A2(n14545), .ZN(n14584) );
  OAI21_X1 U15805 ( .B1(n14545), .B2(n14544), .A(n14584), .ZN(n14546) );
  NAND2_X1 U15806 ( .A1(n14546), .A2(n14690), .ZN(n14554) );
  INV_X1 U15807 ( .A(n14867), .ZN(n14552) );
  NAND2_X1 U15808 ( .A1(n14704), .A2(n14715), .ZN(n14548) );
  NAND2_X1 U15809 ( .A1(n14702), .A2(n14717), .ZN(n14547) );
  NAND2_X1 U15810 ( .A1(n14548), .A2(n14547), .ZN(n14863) );
  INV_X1 U15811 ( .A(n14863), .ZN(n14550) );
  OAI22_X1 U15812 ( .A1(n14706), .A2(n14550), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14549), .ZN(n14551) );
  AOI21_X1 U15813 ( .B1(n14695), .B2(n14552), .A(n14551), .ZN(n14553) );
  OAI211_X1 U15814 ( .C1(n15387), .C2(n14698), .A(n14554), .B(n14553), .ZN(
        P1_U3214) );
  AOI21_X1 U15815 ( .B1(n14556), .B2(n14555), .A(n7276), .ZN(n14563) );
  NOR2_X1 U15816 ( .A1(n14701), .A2(n14557), .ZN(n14560) );
  OAI21_X1 U15817 ( .B1(n14706), .B2(n16004), .A(n14558), .ZN(n14559) );
  AOI211_X1 U15818 ( .C1(n14561), .C2(n14709), .A(n14560), .B(n14559), .ZN(
        n14562) );
  OAI21_X1 U15819 ( .B1(n14563), .B2(n14711), .A(n14562), .ZN(P1_U3215) );
  INV_X1 U15820 ( .A(n15100), .ZN(n14924) );
  INV_X1 U15821 ( .A(n14647), .ZN(n14567) );
  AOI21_X1 U15822 ( .B1(n14663), .B2(n14565), .A(n14564), .ZN(n14566) );
  OAI21_X1 U15823 ( .B1(n14567), .B2(n14566), .A(n14690), .ZN(n14572) );
  OAI22_X1 U15824 ( .A1(n14608), .A2(n14605), .B1(n14568), .B2(n14607), .ZN(
        n15099) );
  INV_X1 U15825 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n14569) );
  OAI22_X1 U15826 ( .A1(n14701), .A2(n14919), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14569), .ZN(n14570) );
  AOI21_X1 U15827 ( .B1(n15099), .B2(n14671), .A(n14570), .ZN(n14571) );
  OAI211_X1 U15828 ( .C1(n14924), .C2(n14698), .A(n14572), .B(n14571), .ZN(
        P1_U3216) );
  XNOR2_X1 U15829 ( .A(n14574), .B(n14573), .ZN(n14575) );
  XNOR2_X1 U15830 ( .A(n14576), .B(n14575), .ZN(n14581) );
  NOR2_X1 U15831 ( .A1(n14701), .A2(n14984), .ZN(n14579) );
  AND2_X1 U15832 ( .A1(n14725), .A2(n14702), .ZN(n14577) );
  AOI21_X1 U15833 ( .B1(n14723), .B2(n14704), .A(n14577), .ZN(n15126) );
  NAND2_X1 U15834 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14819)
         );
  OAI21_X1 U15835 ( .B1(n15126), .B2(n14706), .A(n14819), .ZN(n14578) );
  AOI211_X1 U15836 ( .C1(n14980), .C2(n14709), .A(n14579), .B(n14578), .ZN(
        n14580) );
  OAI21_X1 U15837 ( .B1(n14581), .B2(n14711), .A(n14580), .ZN(P1_U3219) );
  INV_X1 U15838 ( .A(n14582), .ZN(n14583) );
  NAND2_X1 U15839 ( .A1(n14584), .A2(n14583), .ZN(n14594) );
  OAI22_X1 U15840 ( .A1(n14849), .A2(n14585), .B1(n14589), .B2(n14590), .ZN(
        n14587) );
  XNOR2_X1 U15841 ( .A(n14587), .B(n14586), .ZN(n14592) );
  OAI22_X1 U15842 ( .A1(n14849), .A2(n14590), .B1(n14589), .B2(n14588), .ZN(
        n14591) );
  XNOR2_X1 U15843 ( .A(n14592), .B(n14591), .ZN(n14593) );
  XNOR2_X1 U15844 ( .A(n14594), .B(n14593), .ZN(n14601) );
  NOR2_X1 U15845 ( .A1(n14701), .A2(n14850), .ZN(n14598) );
  OAI22_X1 U15846 ( .A1(n14706), .A2(n14596), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14595), .ZN(n14597) );
  AOI211_X1 U15847 ( .C1(n14599), .C2(n14709), .A(n14598), .B(n14597), .ZN(
        n14600) );
  OAI21_X1 U15848 ( .B1(n14601), .B2(n14711), .A(n14600), .ZN(P1_U3220) );
  INV_X1 U15849 ( .A(n15115), .ZN(n14613) );
  OAI21_X1 U15850 ( .B1(n14603), .B2(n14602), .A(n14666), .ZN(n14604) );
  NAND2_X1 U15851 ( .A1(n14604), .A2(n14690), .ZN(n14612) );
  OAI22_X1 U15852 ( .A1(n14608), .A2(n14607), .B1(n14606), .B2(n14605), .ZN(
        n15114) );
  INV_X1 U15853 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n14609) );
  OAI22_X1 U15854 ( .A1(n14701), .A2(n14950), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14609), .ZN(n14610) );
  AOI21_X1 U15855 ( .B1(n15114), .B2(n14671), .A(n14610), .ZN(n14611) );
  OAI211_X1 U15856 ( .C1(n14613), .C2(n14698), .A(n14612), .B(n14611), .ZN(
        P1_U3223) );
  INV_X1 U15857 ( .A(n14614), .ZN(n14618) );
  NOR3_X1 U15858 ( .A1(n14649), .A2(n14616), .A3(n14615), .ZN(n14617) );
  OAI21_X1 U15859 ( .B1(n14618), .B2(n14617), .A(n14690), .ZN(n14625) );
  INV_X1 U15860 ( .A(n14894), .ZN(n14623) );
  NAND2_X1 U15861 ( .A1(n14704), .A2(n14717), .ZN(n14620) );
  NAND2_X1 U15862 ( .A1(n14702), .A2(n14719), .ZN(n14619) );
  AND2_X1 U15863 ( .A1(n14620), .A2(n14619), .ZN(n15085) );
  OAI22_X1 U15864 ( .A1(n14706), .A2(n15085), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14621), .ZN(n14622) );
  AOI21_X1 U15865 ( .B1(n14695), .B2(n14623), .A(n14622), .ZN(n14624) );
  OAI211_X1 U15866 ( .C1(n15392), .C2(n14698), .A(n14625), .B(n14624), .ZN(
        P1_U3225) );
  OAI21_X1 U15867 ( .B1(n14628), .B2(n14627), .A(n14626), .ZN(n14629) );
  NAND2_X1 U15868 ( .A1(n14629), .A2(n14690), .ZN(n14633) );
  AND2_X1 U15869 ( .A1(n14729), .A2(n14702), .ZN(n14630) );
  AOI21_X1 U15870 ( .B1(n14726), .B2(n14704), .A(n14630), .ZN(n15031) );
  NAND2_X1 U15871 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n15568)
         );
  OAI21_X1 U15872 ( .B1(n15031), .B2(n14706), .A(n15568), .ZN(n14631) );
  AOI21_X1 U15873 ( .B1(n14695), .B2(n15037), .A(n14631), .ZN(n14632) );
  OAI211_X1 U15874 ( .C1(n7673), .C2(n14698), .A(n14633), .B(n14632), .ZN(
        P1_U3226) );
  INV_X1 U15875 ( .A(n14634), .ZN(n14639) );
  AOI21_X1 U15876 ( .B1(n14636), .B2(n14638), .A(n14635), .ZN(n14637) );
  AOI21_X1 U15877 ( .B1(n14639), .B2(n14638), .A(n14637), .ZN(n14644) );
  NOR2_X1 U15878 ( .A1(n14701), .A2(n15017), .ZN(n14642) );
  AND2_X1 U15879 ( .A1(n14728), .A2(n14702), .ZN(n14640) );
  AOI21_X1 U15880 ( .B1(n14725), .B2(n14704), .A(n14640), .ZN(n15143) );
  NAND2_X1 U15881 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n15542)
         );
  OAI21_X1 U15882 ( .B1(n15143), .B2(n14706), .A(n15542), .ZN(n14641) );
  AOI211_X1 U15883 ( .C1(n15142), .C2(n14709), .A(n14642), .B(n14641), .ZN(
        n14643) );
  OAI21_X1 U15884 ( .B1(n14644), .B2(n14711), .A(n14643), .ZN(P1_U3228) );
  AND3_X1 U15885 ( .A1(n14647), .A2(n14646), .A3(n14645), .ZN(n14648) );
  OAI21_X1 U15886 ( .B1(n14649), .B2(n14648), .A(n14690), .ZN(n14654) );
  INV_X1 U15887 ( .A(n14906), .ZN(n14652) );
  AOI22_X1 U15888 ( .A1(n14704), .A2(n14718), .B1(n14702), .B2(n14720), .ZN(
        n14903) );
  OAI22_X1 U15889 ( .A1(n14706), .A2(n14903), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14650), .ZN(n14651) );
  AOI21_X1 U15890 ( .B1(n14695), .B2(n14652), .A(n14651), .ZN(n14653) );
  OAI211_X1 U15891 ( .C1(n7668), .C2(n14698), .A(n14654), .B(n14653), .ZN(
        P1_U3229) );
  XNOR2_X1 U15892 ( .A(n14656), .B(n14655), .ZN(n14662) );
  AND2_X1 U15893 ( .A1(n14724), .A2(n14702), .ZN(n14657) );
  AOI21_X1 U15894 ( .B1(n14722), .B2(n14704), .A(n14657), .ZN(n14959) );
  OAI22_X1 U15895 ( .A1(n14959), .A2(n14706), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14658), .ZN(n14660) );
  NOR2_X1 U15896 ( .A1(n15403), .A2(n14698), .ZN(n14659) );
  AOI211_X1 U15897 ( .C1(n14968), .C2(n14695), .A(n14660), .B(n14659), .ZN(
        n14661) );
  OAI21_X1 U15898 ( .B1(n14662), .B2(n14711), .A(n14661), .ZN(P1_U3233) );
  INV_X1 U15899 ( .A(n14663), .ZN(n14668) );
  AOI21_X1 U15900 ( .B1(n14666), .B2(n14665), .A(n14664), .ZN(n14667) );
  NOR3_X1 U15901 ( .A1(n14668), .A2(n14667), .A3(n14711), .ZN(n14675) );
  NAND2_X1 U15902 ( .A1(n14722), .A2(n14702), .ZN(n14670) );
  NAND2_X1 U15903 ( .A1(n14704), .A2(n14720), .ZN(n14669) );
  NAND2_X1 U15904 ( .A1(n14670), .A2(n14669), .ZN(n15105) );
  AOI22_X1 U15905 ( .A1(n15105), .A2(n14671), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14673) );
  NAND2_X1 U15906 ( .A1(n14695), .A2(n14936), .ZN(n14672) );
  OAI211_X1 U15907 ( .C1(n15108), .C2(n14698), .A(n14673), .B(n14672), .ZN(
        n14674) );
  OR2_X1 U15908 ( .A1(n14675), .A2(n14674), .ZN(P1_U3235) );
  OAI21_X1 U15909 ( .B1(n14678), .B2(n14677), .A(n14676), .ZN(n14679) );
  NAND2_X1 U15910 ( .A1(n14679), .A2(n14690), .ZN(n14685) );
  INV_X1 U15911 ( .A(n15001), .ZN(n14683) );
  AND2_X1 U15912 ( .A1(n14726), .A2(n14702), .ZN(n14680) );
  AOI21_X1 U15913 ( .B1(n14724), .B2(n14704), .A(n14680), .ZN(n15138) );
  OAI22_X1 U15914 ( .A1(n15138), .A2(n14706), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14681), .ZN(n14682) );
  AOI21_X1 U15915 ( .B1(n14683), .B2(n14695), .A(n14682), .ZN(n14684) );
  OAI211_X1 U15916 ( .C1(n14686), .C2(n14698), .A(n14685), .B(n14684), .ZN(
        P1_U3238) );
  INV_X1 U15917 ( .A(n15079), .ZN(n14883) );
  OAI21_X1 U15918 ( .B1(n14689), .B2(n14688), .A(n14687), .ZN(n14691) );
  NAND2_X1 U15919 ( .A1(n14691), .A2(n14690), .ZN(n14697) );
  INV_X1 U15920 ( .A(n14880), .ZN(n14694) );
  AOI22_X1 U15921 ( .A1(n14704), .A2(n14716), .B1(n14702), .B2(n14718), .ZN(
        n15076) );
  OAI22_X1 U15922 ( .A1(n14706), .A2(n15076), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14692), .ZN(n14693) );
  AOI21_X1 U15923 ( .B1(n14695), .B2(n14694), .A(n14693), .ZN(n14696) );
  OAI211_X1 U15924 ( .C1(n14883), .C2(n14698), .A(n14697), .B(n14696), .ZN(
        P1_U3240) );
  XNOR2_X1 U15925 ( .A(n14700), .B(n14699), .ZN(n14712) );
  NOR2_X1 U15926 ( .A1(n14701), .A2(n15052), .ZN(n14708) );
  AND2_X1 U15927 ( .A1(n14730), .A2(n14702), .ZN(n14703) );
  AOI21_X1 U15928 ( .B1(n14728), .B2(n14704), .A(n14703), .ZN(n15047) );
  OAI22_X1 U15929 ( .A1(n14706), .A2(n15047), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14705), .ZN(n14707) );
  AOI211_X1 U15930 ( .C1(n15413), .C2(n14709), .A(n14708), .B(n14707), .ZN(
        n14710) );
  OAI21_X1 U15931 ( .B1(n14712), .B2(n14711), .A(n14710), .ZN(P1_U3241) );
  MUX2_X1 U15932 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14713), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15933 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14714), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15934 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14715), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15935 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14716), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15936 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14717), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15937 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14718), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15938 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14719), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15939 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14720), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15940 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14721), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15941 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14722), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15942 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14723), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15943 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14724), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15944 ( .A(n14725), .B(P1_DATAO_REG_18__SCAN_IN), .S(n14727), .Z(
        P1_U3578) );
  MUX2_X1 U15945 ( .A(n14726), .B(P1_DATAO_REG_17__SCAN_IN), .S(n14727), .Z(
        P1_U3577) );
  MUX2_X1 U15946 ( .A(n14728), .B(P1_DATAO_REG_16__SCAN_IN), .S(n14727), .Z(
        P1_U3576) );
  MUX2_X1 U15947 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14729), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15948 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14730), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15949 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14731), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U15950 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14732), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U15951 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14733), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U15952 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14734), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U15953 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14735), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U15954 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14736), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U15955 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14737), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U15956 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14738), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U15957 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14739), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U15958 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14740), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U15959 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14741), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U15960 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14742), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U15961 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14743), .S(P1_U4016), .Z(
        P1_U3561) );
  INV_X1 U15962 ( .A(n14744), .ZN(n14749) );
  MUX2_X1 U15963 ( .A(n11159), .B(P1_REG2_REG_1__SCAN_IN), .S(n14745), .Z(
        n14748) );
  INV_X1 U15964 ( .A(n14746), .ZN(n14747) );
  OAI211_X1 U15965 ( .C1(n14749), .C2(n14748), .A(n15558), .B(n14747), .ZN(
        n14757) );
  OAI211_X1 U15966 ( .C1(n14752), .C2(n14751), .A(n15566), .B(n14750), .ZN(
        n14756) );
  AOI22_X1 U15967 ( .A1(n15544), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14755) );
  NAND2_X1 U15968 ( .A1(n15548), .A2(n14753), .ZN(n14754) );
  NAND4_X1 U15969 ( .A1(n14757), .A2(n14756), .A3(n14755), .A4(n14754), .ZN(
        P1_U3244) );
  OAI22_X1 U15970 ( .A1(n15570), .A2(n15589), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14758), .ZN(n14759) );
  AOI21_X1 U15971 ( .B1(n14760), .B2(n15548), .A(n14759), .ZN(n14774) );
  MUX2_X1 U15972 ( .A(n10344), .B(P1_REG1_REG_3__SCAN_IN), .S(n14760), .Z(
        n14761) );
  NAND3_X1 U15973 ( .A1(n14763), .A2(n14762), .A3(n14761), .ZN(n14764) );
  NAND3_X1 U15974 ( .A1(n15566), .A2(n14765), .A3(n14764), .ZN(n14773) );
  INV_X1 U15975 ( .A(n14766), .ZN(n14771) );
  NAND3_X1 U15976 ( .A1(n14769), .A2(n14768), .A3(n14767), .ZN(n14770) );
  NAND3_X1 U15977 ( .A1(n15558), .A2(n14771), .A3(n14770), .ZN(n14772) );
  NAND3_X1 U15978 ( .A1(n14774), .A2(n14773), .A3(n14772), .ZN(P1_U3246) );
  NOR2_X1 U15979 ( .A1(n15564), .A2(n14775), .ZN(n14776) );
  AOI211_X1 U15980 ( .C1(n15544), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n14777), .B(
        n14776), .ZN(n14788) );
  OAI211_X1 U15981 ( .C1(n14780), .C2(n14779), .A(n15566), .B(n14778), .ZN(
        n14787) );
  OR3_X1 U15982 ( .A1(n14783), .A2(n14782), .A3(n14781), .ZN(n14784) );
  NAND3_X1 U15983 ( .A1(n15558), .A2(n14785), .A3(n14784), .ZN(n14786) );
  NAND3_X1 U15984 ( .A1(n14788), .A2(n14787), .A3(n14786), .ZN(P1_U3249) );
  NOR2_X1 U15985 ( .A1(n14790), .A2(n14789), .ZN(n14792) );
  NOR2_X1 U15986 ( .A1(n14792), .A2(n14791), .ZN(n15555) );
  XNOR2_X1 U15987 ( .A(n15563), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n15556) );
  AOI22_X1 U15988 ( .A1(n15555), .A2(n15556), .B1(P1_REG1_REG_16__SCAN_IN), 
        .B2(n14793), .ZN(n15535) );
  XNOR2_X1 U15989 ( .A(n15540), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n15536) );
  INV_X1 U15990 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14795) );
  OAI22_X1 U15991 ( .A1(n15535), .A2(n15536), .B1(n14795), .B2(n14794), .ZN(
        n14796) );
  XOR2_X1 U15992 ( .A(n15547), .B(n14796), .Z(n15550) );
  NAND2_X1 U15993 ( .A1(n15550), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n15549) );
  NAND2_X1 U15994 ( .A1(n14796), .A2(n15547), .ZN(n14797) );
  NAND2_X1 U15995 ( .A1(n15549), .A2(n14797), .ZN(n14799) );
  XNOR2_X1 U15996 ( .A(n14799), .B(n14798), .ZN(n14815) );
  INV_X1 U15997 ( .A(n14815), .ZN(n14813) );
  NAND2_X1 U15998 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n15540), .ZN(n14807) );
  INV_X1 U15999 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n14804) );
  AOI21_X1 U16000 ( .B1(n14802), .B2(n14801), .A(n14800), .ZN(n15561) );
  NAND2_X1 U16001 ( .A1(n15563), .A2(n14804), .ZN(n14803) );
  OAI211_X1 U16002 ( .C1(n15563), .C2(n14804), .A(n15561), .B(n14803), .ZN(
        n15559) );
  OAI21_X1 U16003 ( .B1(n14804), .B2(n15563), .A(n15559), .ZN(n15538) );
  MUX2_X1 U16004 ( .A(n15016), .B(P1_REG2_REG_17__SCAN_IN), .S(n15540), .Z(
        n15537) );
  INV_X1 U16005 ( .A(n15537), .ZN(n14805) );
  NAND2_X1 U16006 ( .A1(n15538), .A2(n14805), .ZN(n14806) );
  NAND2_X1 U16007 ( .A1(n14807), .A2(n14806), .ZN(n14808) );
  XOR2_X1 U16008 ( .A(n15547), .B(n14808), .Z(n15546) );
  NAND2_X1 U16009 ( .A1(n15546), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n15545) );
  NAND2_X1 U16010 ( .A1(n14808), .A2(n15547), .ZN(n14809) );
  NAND2_X1 U16011 ( .A1(n15545), .A2(n14809), .ZN(n14810) );
  XOR2_X1 U16012 ( .A(n14810), .B(P1_REG2_REG_19__SCAN_IN), .Z(n14814) );
  OAI21_X1 U16013 ( .B1(n14814), .B2(n14811), .A(n15564), .ZN(n14812) );
  AOI21_X1 U16014 ( .B1(n14813), .B2(n15566), .A(n14812), .ZN(n14818) );
  AOI22_X1 U16015 ( .A1(n14815), .A2(n15566), .B1(n15558), .B2(n14814), .ZN(
        n14817) );
  MUX2_X1 U16016 ( .A(n14818), .B(n14817), .S(n14816), .Z(n14820) );
  OAI211_X1 U16017 ( .C1(n8155), .C2(n15570), .A(n14820), .B(n14819), .ZN(
        P1_U3262) );
  INV_X1 U16018 ( .A(n15064), .ZN(n14825) );
  NAND2_X1 U16019 ( .A1(n15062), .A2(n15935), .ZN(n14824) );
  NOR2_X1 U16020 ( .A1(n14822), .A2(n14821), .ZN(n15063) );
  INV_X1 U16021 ( .A(n15063), .ZN(n15066) );
  NOR2_X1 U16022 ( .A1(n15895), .A2(n15066), .ZN(n14830) );
  AOI21_X1 U16023 ( .B1(n15895), .B2(P1_REG2_REG_31__SCAN_IN), .A(n14830), 
        .ZN(n14823) );
  OAI211_X1 U16024 ( .C1(n14825), .C2(n15942), .A(n14824), .B(n14823), .ZN(
        P1_U3263) );
  NAND2_X1 U16025 ( .A1(n14826), .A2(n15382), .ZN(n14827) );
  NAND2_X1 U16026 ( .A1(n14827), .A2(n15878), .ZN(n14828) );
  OR2_X1 U16027 ( .A1(n14829), .A2(n14828), .ZN(n15067) );
  AOI21_X1 U16028 ( .B1(n15895), .B2(P1_REG2_REG_30__SCAN_IN), .A(n14830), 
        .ZN(n14832) );
  NAND2_X1 U16029 ( .A1(n15382), .A2(n15887), .ZN(n14831) );
  OAI211_X1 U16030 ( .C1(n15067), .C2(n15057), .A(n14832), .B(n14831), .ZN(
        P1_U3264) );
  INV_X1 U16031 ( .A(n14833), .ZN(n14847) );
  NOR2_X1 U16032 ( .A1(n14834), .A2(n15057), .ZN(n14844) );
  OAI22_X1 U16033 ( .A1(n14837), .A2(n14836), .B1(n14835), .B2(n15051), .ZN(
        n14840) );
  NOR2_X1 U16034 ( .A1(n15895), .A2(n14838), .ZN(n14839) );
  AOI211_X1 U16035 ( .C1(n15895), .C2(P1_REG2_REG_29__SCAN_IN), .A(n14840), 
        .B(n14839), .ZN(n14841) );
  OAI21_X1 U16036 ( .B1(n14842), .B2(n15942), .A(n14841), .ZN(n14843) );
  AOI211_X1 U16037 ( .C1(n14845), .C2(n15000), .A(n14844), .B(n14843), .ZN(
        n14846) );
  OAI21_X1 U16038 ( .B1(n14847), .B2(n15061), .A(n14846), .ZN(P1_U3356) );
  NAND2_X1 U16039 ( .A1(n14848), .A2(n15054), .ZN(n14856) );
  NOR2_X1 U16040 ( .A1(n14849), .A2(n15942), .ZN(n14853) );
  OAI22_X1 U16041 ( .A1(n15054), .A2(n14851), .B1(n14850), .B2(n15051), .ZN(
        n14852) );
  AOI211_X1 U16042 ( .C1(n14854), .C2(n15935), .A(n14853), .B(n14852), .ZN(
        n14855) );
  OAI211_X1 U16043 ( .C1(n14858), .C2(n14857), .A(n14856), .B(n14855), .ZN(
        P1_U3265) );
  XNOR2_X1 U16044 ( .A(n14859), .B(n14861), .ZN(n15070) );
  INV_X1 U16045 ( .A(n15070), .ZN(n14875) );
  AOI21_X1 U16046 ( .B1(n14864), .B2(n16013), .A(n14863), .ZN(n15073) );
  INV_X1 U16047 ( .A(n15073), .ZN(n14873) );
  AOI21_X1 U16048 ( .B1(n14878), .B2(n14870), .A(n15985), .ZN(n14866) );
  NAND2_X1 U16049 ( .A1(n14866), .A2(n14865), .ZN(n15071) );
  OAI22_X1 U16050 ( .A1(n15054), .A2(n14868), .B1(n14867), .B2(n15051), .ZN(
        n14869) );
  AOI21_X1 U16051 ( .B1(n14870), .B2(n15887), .A(n14869), .ZN(n14871) );
  OAI21_X1 U16052 ( .B1(n15071), .B2(n15057), .A(n14871), .ZN(n14872) );
  AOI21_X1 U16053 ( .B1(n14873), .B2(n15054), .A(n14872), .ZN(n14874) );
  OAI21_X1 U16054 ( .B1(n14875), .B2(n15061), .A(n14874), .ZN(P1_U3266) );
  OAI21_X1 U16055 ( .B1(n14877), .B2(n14885), .A(n14876), .ZN(n15083) );
  INV_X1 U16056 ( .A(n14878), .ZN(n14879) );
  AOI211_X1 U16057 ( .C1(n15079), .C2(n14892), .A(n15985), .B(n14879), .ZN(
        n15077) );
  OAI22_X1 U16058 ( .A1(n15895), .A2(n15076), .B1(n14880), .B2(n15051), .ZN(
        n14881) );
  AOI21_X1 U16059 ( .B1(P1_REG2_REG_26__SCAN_IN), .B2(n15895), .A(n14881), 
        .ZN(n14882) );
  OAI21_X1 U16060 ( .B1(n14883), .B2(n15942), .A(n14882), .ZN(n14884) );
  AOI21_X1 U16061 ( .B1(n15077), .B2(n15935), .A(n14884), .ZN(n14888) );
  XNOR2_X1 U16062 ( .A(n14886), .B(n14885), .ZN(n15080) );
  NAND2_X1 U16063 ( .A1(n15080), .A2(n15022), .ZN(n14887) );
  OAI211_X1 U16064 ( .C1(n15083), .C2(n15024), .A(n14888), .B(n14887), .ZN(
        P1_U3267) );
  XNOR2_X1 U16065 ( .A(n14889), .B(n14890), .ZN(n15084) );
  INV_X1 U16066 ( .A(n15084), .ZN(n14901) );
  XNOR2_X1 U16067 ( .A(n14891), .B(n14890), .ZN(n15088) );
  OAI211_X1 U16068 ( .C1(n7188), .C2(n15392), .A(n15878), .B(n14892), .ZN(
        n15086) );
  NOR2_X1 U16069 ( .A1(n15054), .A2(n14893), .ZN(n14896) );
  OAI22_X1 U16070 ( .A1(n15895), .A2(n15085), .B1(n14894), .B2(n15051), .ZN(
        n14895) );
  AOI211_X1 U16071 ( .C1(n14897), .C2(n15887), .A(n14896), .B(n14895), .ZN(
        n14898) );
  OAI21_X1 U16072 ( .B1(n15086), .B2(n15057), .A(n14898), .ZN(n14899) );
  AOI21_X1 U16073 ( .B1(n15088), .B2(n15000), .A(n14899), .ZN(n14900) );
  OAI21_X1 U16074 ( .B1(n14901), .B2(n15061), .A(n14900), .ZN(P1_U3268) );
  XNOR2_X1 U16075 ( .A(n14902), .B(n14911), .ZN(n14904) );
  OAI21_X1 U16076 ( .B1(n14904), .B2(n15987), .A(n14903), .ZN(n15093) );
  INV_X1 U16077 ( .A(n15093), .ZN(n14914) );
  AOI211_X1 U16078 ( .C1(n14905), .C2(n14917), .A(n15985), .B(n7188), .ZN(
        n15094) );
  NOR2_X1 U16079 ( .A1(n7668), .A2(n15942), .ZN(n14909) );
  OAI22_X1 U16080 ( .A1(n15054), .A2(n14907), .B1(n14906), .B2(n15051), .ZN(
        n14908) );
  AOI211_X1 U16081 ( .C1(n15094), .C2(n15935), .A(n14909), .B(n14908), .ZN(
        n14913) );
  OAI21_X1 U16082 ( .B1(n7252), .B2(n14911), .A(n14910), .ZN(n15095) );
  NAND2_X1 U16083 ( .A1(n15095), .A2(n15022), .ZN(n14912) );
  OAI211_X1 U16084 ( .C1(n14914), .C2(n15895), .A(n14913), .B(n14912), .ZN(
        P1_U3269) );
  XNOR2_X1 U16085 ( .A(n14916), .B(n14915), .ZN(n15101) );
  AOI21_X1 U16086 ( .B1(n15100), .B2(n14939), .A(n15985), .ZN(n14918) );
  AND2_X1 U16087 ( .A1(n14918), .A2(n14917), .ZN(n15098) );
  NAND2_X1 U16088 ( .A1(n15098), .A2(n15935), .ZN(n14923) );
  OAI22_X1 U16089 ( .A1(n15054), .A2(n14920), .B1(n14919), .B2(n15051), .ZN(
        n14921) );
  AOI21_X1 U16090 ( .B1(n15099), .B2(n15054), .A(n14921), .ZN(n14922) );
  OAI211_X1 U16091 ( .C1(n14924), .C2(n15942), .A(n14923), .B(n14922), .ZN(
        n14929) );
  OAI21_X1 U16092 ( .B1(n14927), .B2(n14926), .A(n14925), .ZN(n15104) );
  NOR2_X1 U16093 ( .A1(n15104), .A2(n15061), .ZN(n14928) );
  AOI211_X1 U16094 ( .C1(n15000), .C2(n15101), .A(n14929), .B(n14928), .ZN(
        n14930) );
  INV_X1 U16095 ( .A(n14930), .ZN(P1_U3270) );
  OAI21_X1 U16096 ( .B1(n14934), .B2(n14932), .A(n14931), .ZN(n14933) );
  INV_X1 U16097 ( .A(n14933), .ZN(n15112) );
  OAI21_X1 U16098 ( .B1(n7864), .B2(n7241), .A(n14935), .ZN(n15110) );
  AOI22_X1 U16099 ( .A1(n14936), .A2(n15938), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n15895), .ZN(n14938) );
  NAND2_X1 U16100 ( .A1(n15105), .A2(n15054), .ZN(n14937) );
  OAI211_X1 U16101 ( .C1(n15108), .C2(n15942), .A(n14938), .B(n14937), .ZN(
        n14941) );
  OAI211_X1 U16102 ( .C1(n15108), .C2(n14953), .A(n15878), .B(n14939), .ZN(
        n15107) );
  NOR2_X1 U16103 ( .A1(n15107), .A2(n15057), .ZN(n14940) );
  AOI211_X1 U16104 ( .C1(n15110), .C2(n15022), .A(n14941), .B(n14940), .ZN(
        n14942) );
  OAI21_X1 U16105 ( .B1(n15112), .B2(n15024), .A(n14942), .ZN(P1_U3271) );
  XNOR2_X1 U16106 ( .A(n14944), .B(n14943), .ZN(n15116) );
  OAI21_X1 U16107 ( .B1(n14947), .B2(n14946), .A(n14945), .ZN(n15119) );
  NAND2_X1 U16108 ( .A1(n15114), .A2(n15054), .ZN(n14949) );
  NAND2_X1 U16109 ( .A1(n15895), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n14948) );
  OAI211_X1 U16110 ( .C1(n15051), .C2(n14950), .A(n14949), .B(n14948), .ZN(
        n14951) );
  AOI21_X1 U16111 ( .B1(n15115), .B2(n15887), .A(n14951), .ZN(n14955) );
  AND2_X1 U16112 ( .A1(n15115), .A2(n14964), .ZN(n14952) );
  NOR3_X1 U16113 ( .A1(n14953), .A2(n14952), .A3(n15985), .ZN(n15113) );
  NAND2_X1 U16114 ( .A1(n15113), .A2(n15935), .ZN(n14954) );
  OAI211_X1 U16115 ( .C1(n15119), .C2(n15024), .A(n14955), .B(n14954), .ZN(
        n14956) );
  AOI21_X1 U16116 ( .B1(n15022), .B2(n15116), .A(n14956), .ZN(n14957) );
  INV_X1 U16117 ( .A(n14957), .ZN(P1_U3272) );
  OAI211_X1 U16118 ( .C1(n7234), .C2(n7952), .A(n16013), .B(n14958), .ZN(
        n14960) );
  NAND2_X1 U16119 ( .A1(n14960), .A2(n14959), .ZN(n15121) );
  INV_X1 U16120 ( .A(n15121), .ZN(n14973) );
  NAND2_X1 U16121 ( .A1(n7952), .A2(n14961), .ZN(n14962) );
  INV_X1 U16122 ( .A(n14983), .ZN(n14966) );
  INV_X1 U16123 ( .A(n14964), .ZN(n14965) );
  AOI211_X1 U16124 ( .C1(n14967), .C2(n14966), .A(n15985), .B(n14965), .ZN(
        n15120) );
  NAND2_X1 U16125 ( .A1(n15120), .A2(n15935), .ZN(n14970) );
  AOI22_X1 U16126 ( .A1(P1_REG2_REG_20__SCAN_IN), .A2(n15895), .B1(n14968), 
        .B2(n15938), .ZN(n14969) );
  OAI211_X1 U16127 ( .C1(n15403), .C2(n15942), .A(n14970), .B(n14969), .ZN(
        n14971) );
  AOI21_X1 U16128 ( .B1(n15022), .B2(n15122), .A(n14971), .ZN(n14972) );
  OAI21_X1 U16129 ( .B1(n15895), .B2(n14973), .A(n14972), .ZN(P1_U3273) );
  INV_X1 U16130 ( .A(n14974), .ZN(n14975) );
  AOI21_X1 U16131 ( .B1(n14978), .B2(n14976), .A(n14975), .ZN(n15132) );
  OAI21_X1 U16132 ( .B1(n14979), .B2(n14978), .A(n14977), .ZN(n15130) );
  INV_X1 U16133 ( .A(n14980), .ZN(n15127) );
  NAND2_X1 U16134 ( .A1(n14980), .A2(n14997), .ZN(n14981) );
  NAND2_X1 U16135 ( .A1(n14981), .A2(n15878), .ZN(n14982) );
  NOR2_X1 U16136 ( .A1(n14983), .A2(n14982), .ZN(n15128) );
  NAND2_X1 U16137 ( .A1(n15128), .A2(n15935), .ZN(n14989) );
  INV_X1 U16138 ( .A(n15126), .ZN(n14987) );
  INV_X1 U16139 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14985) );
  OAI22_X1 U16140 ( .A1(n15054), .A2(n14985), .B1(n14984), .B2(n15051), .ZN(
        n14986) );
  AOI21_X1 U16141 ( .B1(n14987), .B2(n15054), .A(n14986), .ZN(n14988) );
  OAI211_X1 U16142 ( .C1(n15127), .C2(n15942), .A(n14989), .B(n14988), .ZN(
        n14990) );
  AOI21_X1 U16143 ( .B1(n15022), .B2(n15130), .A(n14990), .ZN(n14991) );
  OAI21_X1 U16144 ( .B1(n15132), .B2(n15024), .A(n14991), .ZN(P1_U3274) );
  OAI21_X1 U16145 ( .B1(n14994), .B2(n14993), .A(n14992), .ZN(n15133) );
  INV_X1 U16146 ( .A(n15015), .ZN(n14995) );
  AOI21_X1 U16147 ( .B1(n15407), .B2(n14995), .A(n15985), .ZN(n14996) );
  NAND2_X1 U16148 ( .A1(n14997), .A2(n14996), .ZN(n15136) );
  OR2_X1 U16149 ( .A1(n14999), .A2(n14998), .ZN(n15135) );
  NAND3_X1 U16150 ( .A1(n15135), .A2(n15134), .A3(n15000), .ZN(n15007) );
  INV_X1 U16151 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n15002) );
  OAI22_X1 U16152 ( .A1(n15054), .A2(n15002), .B1(n15001), .B2(n15051), .ZN(
        n15003) );
  INV_X1 U16153 ( .A(n15003), .ZN(n15004) );
  OAI21_X1 U16154 ( .B1(n15138), .B2(n15895), .A(n15004), .ZN(n15005) );
  AOI21_X1 U16155 ( .B1(n15407), .B2(n15887), .A(n15005), .ZN(n15006) );
  OAI211_X1 U16156 ( .C1(n15136), .C2(n15057), .A(n15007), .B(n15006), .ZN(
        n15008) );
  AOI21_X1 U16157 ( .B1(n15022), .B2(n15133), .A(n15008), .ZN(n15009) );
  INV_X1 U16158 ( .A(n15009), .ZN(P1_U3275) );
  XOR2_X1 U16159 ( .A(n15010), .B(n15013), .Z(n15149) );
  AOI21_X1 U16160 ( .B1(n15013), .B2(n15012), .A(n7908), .ZN(n15147) );
  AND2_X1 U16161 ( .A1(n15142), .A2(n15035), .ZN(n15014) );
  OR3_X1 U16162 ( .A1(n15015), .A2(n15014), .A3(n15985), .ZN(n15144) );
  NOR2_X1 U16163 ( .A1(n15054), .A2(n15016), .ZN(n15019) );
  OAI22_X1 U16164 ( .A1(n15143), .A2(n15895), .B1(n15017), .B2(n15051), .ZN(
        n15018) );
  AOI211_X1 U16165 ( .C1(n15142), .C2(n15887), .A(n15019), .B(n15018), .ZN(
        n15020) );
  OAI21_X1 U16166 ( .B1(n15144), .B2(n15057), .A(n15020), .ZN(n15021) );
  AOI21_X1 U16167 ( .B1(n15147), .B2(n15022), .A(n15021), .ZN(n15023) );
  OAI21_X1 U16168 ( .B1(n15149), .B2(n15024), .A(n15023), .ZN(P1_U3276) );
  OAI21_X1 U16169 ( .B1(n15027), .B2(n15026), .A(n15025), .ZN(n15028) );
  INV_X1 U16170 ( .A(n15028), .ZN(n15154) );
  OAI21_X1 U16171 ( .B1(n7274), .B2(n15030), .A(n15029), .ZN(n15033) );
  INV_X1 U16172 ( .A(n15031), .ZN(n15032) );
  AOI21_X1 U16173 ( .B1(n15033), .B2(n16013), .A(n15032), .ZN(n15153) );
  NAND2_X1 U16174 ( .A1(n15049), .A2(n15150), .ZN(n15034) );
  AND2_X1 U16175 ( .A1(n15035), .A2(n15034), .ZN(n15151) );
  AOI22_X1 U16176 ( .A1(n15151), .A2(n7785), .B1(n15037), .B2(n15938), .ZN(
        n15038) );
  AOI21_X1 U16177 ( .B1(n15153), .B2(n15038), .A(n15895), .ZN(n15039) );
  INV_X1 U16178 ( .A(n15039), .ZN(n15041) );
  AOI22_X1 U16179 ( .A1(n15150), .A2(n15887), .B1(P1_REG2_REG_16__SCAN_IN), 
        .B2(n15895), .ZN(n15040) );
  OAI211_X1 U16180 ( .C1(n15154), .C2(n15061), .A(n15041), .B(n15040), .ZN(
        P1_U3277) );
  XNOR2_X1 U16181 ( .A(n15043), .B(n15042), .ZN(n15157) );
  OAI211_X1 U16182 ( .C1(n15046), .C2(n15045), .A(n15044), .B(n16013), .ZN(
        n15048) );
  AND2_X1 U16183 ( .A1(n15048), .A2(n15047), .ZN(n15156) );
  INV_X1 U16184 ( .A(n15156), .ZN(n15059) );
  OAI211_X1 U16185 ( .C1(n15050), .C2(n7270), .A(n15878), .B(n15049), .ZN(
        n15155) );
  OAI22_X1 U16186 ( .A1(n15054), .A2(n15053), .B1(n15052), .B2(n15051), .ZN(
        n15055) );
  AOI21_X1 U16187 ( .B1(n15413), .B2(n15887), .A(n15055), .ZN(n15056) );
  OAI21_X1 U16188 ( .B1(n15155), .B2(n15057), .A(n15056), .ZN(n15058) );
  AOI21_X1 U16189 ( .B1(n15059), .B2(n15054), .A(n15058), .ZN(n15060) );
  OAI21_X1 U16190 ( .B1(n15157), .B2(n15061), .A(n15060), .ZN(P1_U3278) );
  NAND2_X1 U16191 ( .A1(n7362), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n15065) );
  OAI21_X1 U16192 ( .B1(n15160), .B2(n7362), .A(n15065), .ZN(P1_U3559) );
  NAND2_X1 U16193 ( .A1(n15067), .A2(n15066), .ZN(n15380) );
  MUX2_X1 U16194 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15380), .S(n16014), .Z(
        n15068) );
  AOI21_X1 U16195 ( .B1(n10229), .B2(n15382), .A(n15068), .ZN(n15069) );
  INV_X1 U16196 ( .A(n15069), .ZN(P1_U3558) );
  NAND2_X1 U16197 ( .A1(n15070), .A2(n15992), .ZN(n15072) );
  MUX2_X1 U16198 ( .A(n15074), .B(n15384), .S(n16014), .Z(n15075) );
  INV_X1 U16199 ( .A(n15076), .ZN(n15078) );
  AOI211_X1 U16200 ( .C1(n15079), .C2(n15982), .A(n15078), .B(n15077), .ZN(
        n15082) );
  NAND2_X1 U16201 ( .A1(n15080), .A2(n15992), .ZN(n15081) );
  OAI211_X1 U16202 ( .C1(n15987), .C2(n15083), .A(n15082), .B(n15081), .ZN(
        n15388) );
  MUX2_X1 U16203 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15388), .S(n16014), .Z(
        P1_U3554) );
  INV_X1 U16204 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n15091) );
  NAND2_X1 U16205 ( .A1(n15084), .A2(n15992), .ZN(n15090) );
  NAND2_X1 U16206 ( .A1(n15086), .A2(n15085), .ZN(n15087) );
  AOI21_X1 U16207 ( .B1(n15088), .B2(n16013), .A(n15087), .ZN(n15089) );
  AND2_X1 U16208 ( .A1(n15090), .A2(n15089), .ZN(n15389) );
  MUX2_X1 U16209 ( .A(n15091), .B(n15389), .S(n16014), .Z(n15092) );
  OAI21_X1 U16210 ( .B1(n15392), .B2(n15125), .A(n15092), .ZN(P1_U3553) );
  INV_X1 U16211 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n15096) );
  AOI211_X1 U16212 ( .C1(n15992), .C2(n15095), .A(n15094), .B(n15093), .ZN(
        n15393) );
  MUX2_X1 U16213 ( .A(n15096), .B(n15393), .S(n16014), .Z(n15097) );
  OAI21_X1 U16214 ( .B1(n7668), .B2(n15125), .A(n15097), .ZN(P1_U3552) );
  AOI211_X1 U16215 ( .C1(n15100), .C2(n15982), .A(n15099), .B(n15098), .ZN(
        n15103) );
  NAND2_X1 U16216 ( .A1(n15101), .A2(n16013), .ZN(n15102) );
  OAI211_X1 U16217 ( .C1(n16008), .C2(n15104), .A(n15103), .B(n15102), .ZN(
        n15396) );
  MUX2_X1 U16218 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15396), .S(n16014), .Z(
        P1_U3551) );
  INV_X1 U16219 ( .A(n15105), .ZN(n15106) );
  OAI211_X1 U16220 ( .C1(n16006), .C2(n15108), .A(n15107), .B(n15106), .ZN(
        n15109) );
  AOI21_X1 U16221 ( .B1(n15110), .B2(n15992), .A(n15109), .ZN(n15111) );
  OAI21_X1 U16222 ( .B1(n15987), .B2(n15112), .A(n15111), .ZN(n15397) );
  MUX2_X1 U16223 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15397), .S(n16014), .Z(
        P1_U3550) );
  AOI211_X1 U16224 ( .C1(n15115), .C2(n15982), .A(n15114), .B(n15113), .ZN(
        n15118) );
  NAND2_X1 U16225 ( .A1(n15116), .A2(n15992), .ZN(n15117) );
  OAI211_X1 U16226 ( .C1(n15987), .C2(n15119), .A(n15118), .B(n15117), .ZN(
        n15398) );
  MUX2_X1 U16227 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15398), .S(n16014), .Z(
        P1_U3549) );
  INV_X1 U16228 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n15123) );
  AOI211_X1 U16229 ( .C1(n15122), .C2(n15992), .A(n15121), .B(n15120), .ZN(
        n15399) );
  MUX2_X1 U16230 ( .A(n15123), .B(n15399), .S(n16014), .Z(n15124) );
  OAI21_X1 U16231 ( .B1(n15403), .B2(n15125), .A(n15124), .ZN(P1_U3548) );
  OAI21_X1 U16232 ( .B1(n15127), .B2(n16006), .A(n15126), .ZN(n15129) );
  AOI211_X1 U16233 ( .C1(n15130), .C2(n15992), .A(n15129), .B(n15128), .ZN(
        n15131) );
  OAI21_X1 U16234 ( .B1(n15132), .B2(n15987), .A(n15131), .ZN(n15404) );
  MUX2_X1 U16235 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15404), .S(n16014), .Z(
        P1_U3547) );
  NAND2_X1 U16236 ( .A1(n15133), .A2(n15992), .ZN(n15139) );
  NAND3_X1 U16237 ( .A1(n15135), .A2(n15134), .A3(n16013), .ZN(n15137) );
  NAND4_X1 U16238 ( .A1(n15139), .A2(n15138), .A3(n15137), .A4(n15136), .ZN(
        n15405) );
  MUX2_X1 U16239 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15405), .S(n16014), .Z(
        n15140) );
  AOI21_X1 U16240 ( .B1(n10229), .B2(n15407), .A(n15140), .ZN(n15141) );
  INV_X1 U16241 ( .A(n15141), .ZN(P1_U3546) );
  INV_X1 U16242 ( .A(n15142), .ZN(n15145) );
  OAI211_X1 U16243 ( .C1(n15145), .C2(n16006), .A(n15144), .B(n15143), .ZN(
        n15146) );
  AOI21_X1 U16244 ( .B1(n15147), .B2(n15992), .A(n15146), .ZN(n15148) );
  OAI21_X1 U16245 ( .B1(n15987), .B2(n15149), .A(n15148), .ZN(n15409) );
  MUX2_X1 U16246 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15409), .S(n16014), .Z(
        P1_U3545) );
  AOI22_X1 U16247 ( .A1(n15151), .A2(n15878), .B1(n15150), .B2(n15982), .ZN(
        n15152) );
  OAI211_X1 U16248 ( .C1(n16008), .C2(n15154), .A(n15153), .B(n15152), .ZN(
        n15410) );
  MUX2_X1 U16249 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15410), .S(n16014), .Z(
        P1_U3544) );
  OAI211_X1 U16250 ( .C1(n16008), .C2(n15157), .A(n15156), .B(n15155), .ZN(
        n15411) );
  MUX2_X1 U16251 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15411), .S(n16014), .Z(
        n15158) );
  AOI21_X1 U16252 ( .B1(n10229), .B2(n15413), .A(n15158), .ZN(n15159) );
  INV_X1 U16253 ( .A(n15159), .ZN(P1_U3543) );
  XNOR2_X1 U16254 ( .A(n15162), .B(keyinput_126), .ZN(n15378) );
  INV_X1 U16255 ( .A(keyinput_117), .ZN(n15245) );
  INV_X1 U16256 ( .A(keyinput_116), .ZN(n15243) );
  INV_X1 U16257 ( .A(keyinput_115), .ZN(n15241) );
  OAI22_X1 U16258 ( .A1(P3_REG3_REG_21__SCAN_IN), .A2(keyinput_109), .B1(
        P3_REG3_REG_17__SCAN_IN), .B2(keyinput_114), .ZN(n15163) );
  AOI221_X1 U16259 ( .B1(P3_REG3_REG_21__SCAN_IN), .B2(keyinput_109), .C1(
        keyinput_114), .C2(P3_REG3_REG_17__SCAN_IN), .A(n15163), .ZN(n15239)
         );
  OAI22_X1 U16260 ( .A1(n15165), .A2(keyinput_110), .B1(keyinput_112), .B2(
        P3_REG3_REG_16__SCAN_IN), .ZN(n15164) );
  AOI221_X1 U16261 ( .B1(n15165), .B2(keyinput_110), .C1(
        P3_REG3_REG_16__SCAN_IN), .C2(keyinput_112), .A(n15164), .ZN(n15238)
         );
  OAI22_X1 U16262 ( .A1(P3_REG3_REG_25__SCAN_IN), .A2(keyinput_111), .B1(
        keyinput_113), .B2(P3_REG3_REG_5__SCAN_IN), .ZN(n15166) );
  AOI221_X1 U16263 ( .B1(P3_REG3_REG_25__SCAN_IN), .B2(keyinput_111), .C1(
        P3_REG3_REG_5__SCAN_IN), .C2(keyinput_113), .A(n15166), .ZN(n15237) );
  AOI22_X1 U16264 ( .A1(n15269), .A2(keyinput_107), .B1(n8181), .B2(
        keyinput_106), .ZN(n15167) );
  OAI221_X1 U16265 ( .B1(n15269), .B2(keyinput_107), .C1(n8181), .C2(
        keyinput_106), .A(n15167), .ZN(n15235) );
  AOI22_X1 U16266 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(keyinput_103), .B1(
        n15169), .B2(keyinput_104), .ZN(n15168) );
  OAI221_X1 U16267 ( .B1(P3_REG3_REG_10__SCAN_IN), .B2(keyinput_103), .C1(
        n15169), .C2(keyinput_104), .A(n15168), .ZN(n15230) );
  AOI22_X1 U16268 ( .A1(P3_RD_REG_SCAN_IN), .A2(keyinput_97), .B1(n9657), .B2(
        keyinput_96), .ZN(n15170) );
  OAI221_X1 U16269 ( .B1(P3_RD_REG_SCAN_IN), .B2(keyinput_97), .C1(n9657), 
        .C2(keyinput_96), .A(n15170), .ZN(n15222) );
  OAI22_X1 U16270 ( .A1(n15318), .A2(keyinput_83), .B1(n15172), .B2(
        keyinput_84), .ZN(n15171) );
  AOI221_X1 U16271 ( .B1(n15318), .B2(keyinput_83), .C1(keyinput_84), .C2(
        n15172), .A(n15171), .ZN(n15220) );
  INV_X1 U16272 ( .A(keyinput_82), .ZN(n15202) );
  INV_X1 U16273 ( .A(keyinput_81), .ZN(n15200) );
  INV_X1 U16274 ( .A(keyinput_80), .ZN(n15198) );
  INV_X1 U16275 ( .A(keyinput_74), .ZN(n15189) );
  INV_X1 U16276 ( .A(keyinput_73), .ZN(n15187) );
  AOI22_X1 U16277 ( .A1(SI_26_), .A2(keyinput_70), .B1(n15174), .B2(
        keyinput_71), .ZN(n15173) );
  OAI221_X1 U16278 ( .B1(SI_26_), .B2(keyinput_70), .C1(n15174), .C2(
        keyinput_71), .A(n15173), .ZN(n15183) );
  AOI22_X1 U16279 ( .A1(SI_28_), .A2(keyinput_68), .B1(SI_29_), .B2(
        keyinput_67), .ZN(n15175) );
  OAI221_X1 U16280 ( .B1(SI_28_), .B2(keyinput_68), .C1(SI_29_), .C2(
        keyinput_67), .A(n15175), .ZN(n15180) );
  INV_X1 U16281 ( .A(keyinput_66), .ZN(n15178) );
  OAI22_X1 U16282 ( .A1(SI_31_), .A2(keyinput_65), .B1(P3_WR_REG_SCAN_IN), 
        .B2(keyinput_64), .ZN(n15176) );
  AOI221_X1 U16283 ( .B1(SI_31_), .B2(keyinput_65), .C1(keyinput_64), .C2(
        P3_WR_REG_SCAN_IN), .A(n15176), .ZN(n15177) );
  AOI221_X1 U16284 ( .B1(SI_30_), .B2(n15178), .C1(n15284), .C2(keyinput_66), 
        .A(n15177), .ZN(n15179) );
  OAI22_X1 U16285 ( .A1(keyinput_69), .A2(n15289), .B1(n15180), .B2(n15179), 
        .ZN(n15181) );
  AOI21_X1 U16286 ( .B1(keyinput_69), .B2(n15289), .A(n15181), .ZN(n15182) );
  OAI22_X1 U16287 ( .A1(keyinput_72), .A2(n15185), .B1(n15183), .B2(n15182), 
        .ZN(n15184) );
  AOI21_X1 U16288 ( .B1(keyinput_72), .B2(n15185), .A(n15184), .ZN(n15186) );
  AOI221_X1 U16289 ( .B1(SI_23_), .B2(keyinput_73), .C1(n15294), .C2(n15187), 
        .A(n15186), .ZN(n15188) );
  AOI221_X1 U16290 ( .B1(SI_22_), .B2(keyinput_74), .C1(n15297), .C2(n15189), 
        .A(n15188), .ZN(n15196) );
  XNOR2_X1 U16291 ( .A(SI_21_), .B(keyinput_75), .ZN(n15195) );
  OAI22_X1 U16292 ( .A1(n15191), .A2(keyinput_76), .B1(n15301), .B2(
        keyinput_79), .ZN(n15190) );
  AOI221_X1 U16293 ( .B1(n15191), .B2(keyinput_76), .C1(keyinput_79), .C2(
        n15301), .A(n15190), .ZN(n15194) );
  OAI22_X1 U16294 ( .A1(SI_19_), .A2(keyinput_77), .B1(keyinput_78), .B2(
        SI_18_), .ZN(n15192) );
  AOI221_X1 U16295 ( .B1(SI_19_), .B2(keyinput_77), .C1(SI_18_), .C2(
        keyinput_78), .A(n15192), .ZN(n15193) );
  OAI211_X1 U16296 ( .C1(n15196), .C2(n15195), .A(n15194), .B(n15193), .ZN(
        n15197) );
  OAI221_X1 U16297 ( .B1(SI_16_), .B2(n15198), .C1(n15310), .C2(keyinput_80), 
        .A(n15197), .ZN(n15199) );
  OAI221_X1 U16298 ( .B1(SI_15_), .B2(n15200), .C1(n15313), .C2(keyinput_81), 
        .A(n15199), .ZN(n15201) );
  OAI221_X1 U16299 ( .B1(SI_14_), .B2(n15202), .C1(n15315), .C2(keyinput_82), 
        .A(n15201), .ZN(n15219) );
  OAI22_X1 U16300 ( .A1(n15320), .A2(keyinput_87), .B1(keyinput_92), .B2(SI_4_), .ZN(n15203) );
  AOI221_X1 U16301 ( .B1(n15320), .B2(keyinput_87), .C1(SI_4_), .C2(
        keyinput_92), .A(n15203), .ZN(n15212) );
  OAI22_X1 U16302 ( .A1(SI_10_), .A2(keyinput_86), .B1(keyinput_90), .B2(SI_6_), .ZN(n15204) );
  AOI221_X1 U16303 ( .B1(SI_10_), .B2(keyinput_86), .C1(SI_6_), .C2(
        keyinput_90), .A(n15204), .ZN(n15211) );
  OAI22_X1 U16304 ( .A1(n15207), .A2(keyinput_88), .B1(n15206), .B2(
        keyinput_91), .ZN(n15205) );
  AOI221_X1 U16305 ( .B1(n15207), .B2(keyinput_88), .C1(keyinput_91), .C2(
        n15206), .A(n15205), .ZN(n15210) );
  OAI22_X1 U16306 ( .A1(SI_11_), .A2(keyinput_85), .B1(keyinput_94), .B2(SI_2_), .ZN(n15208) );
  AOI221_X1 U16307 ( .B1(SI_11_), .B2(keyinput_85), .C1(SI_2_), .C2(
        keyinput_94), .A(n15208), .ZN(n15209) );
  NAND4_X1 U16308 ( .A1(n15212), .A2(n15211), .A3(n15210), .A4(n15209), .ZN(
        n15216) );
  XOR2_X1 U16309 ( .A(SI_3_), .B(keyinput_93), .Z(n15215) );
  AND2_X1 U16310 ( .A1(SI_7_), .A2(keyinput_89), .ZN(n15214) );
  XNOR2_X1 U16311 ( .A(SI_1_), .B(keyinput_95), .ZN(n15213) );
  NOR4_X1 U16312 ( .A1(n15216), .A2(n15215), .A3(n15214), .A4(n15213), .ZN(
        n15217) );
  OAI21_X1 U16313 ( .B1(keyinput_89), .B2(SI_7_), .A(n15217), .ZN(n15218) );
  AOI21_X1 U16314 ( .B1(n15220), .B2(n15219), .A(n15218), .ZN(n15221) );
  OAI22_X1 U16315 ( .A1(n15222), .A2(n15221), .B1(P3_U3151), .B2(keyinput_98), 
        .ZN(n15223) );
  AOI21_X1 U16316 ( .B1(P3_U3151), .B2(keyinput_98), .A(n15223), .ZN(n15228)
         );
  OAI22_X1 U16317 ( .A1(n15272), .A2(keyinput_100), .B1(keyinput_99), .B2(
        P3_REG3_REG_7__SCAN_IN), .ZN(n15224) );
  AOI221_X1 U16318 ( .B1(n15272), .B2(keyinput_100), .C1(
        P3_REG3_REG_7__SCAN_IN), .C2(keyinput_99), .A(n15224), .ZN(n15227) );
  INV_X1 U16319 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n15338) );
  AOI22_X1 U16320 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(keyinput_101), .B1(
        n15338), .B2(keyinput_102), .ZN(n15225) );
  OAI221_X1 U16321 ( .B1(P3_REG3_REG_14__SCAN_IN), .B2(keyinput_101), .C1(
        n15338), .C2(keyinput_102), .A(n15225), .ZN(n15226) );
  AOI21_X1 U16322 ( .B1(n15228), .B2(n15227), .A(n15226), .ZN(n15229) );
  OAI22_X1 U16323 ( .A1(keyinput_105), .A2(n15232), .B1(n15230), .B2(n15229), 
        .ZN(n15231) );
  AOI21_X1 U16324 ( .B1(keyinput_105), .B2(n15232), .A(n15231), .ZN(n15234) );
  NAND2_X1 U16325 ( .A1(n8223), .A2(keyinput_108), .ZN(n15233) );
  OAI221_X1 U16326 ( .B1(n15235), .B2(n15234), .C1(n8223), .C2(keyinput_108), 
        .A(n15233), .ZN(n15236) );
  NAND4_X1 U16327 ( .A1(n15239), .A2(n15238), .A3(n15237), .A4(n15236), .ZN(
        n15240) );
  OAI221_X1 U16328 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(keyinput_115), .C1(
        n15354), .C2(n15241), .A(n15240), .ZN(n15242) );
  OAI221_X1 U16329 ( .B1(P3_REG3_REG_4__SCAN_IN), .B2(keyinput_116), .C1(
        n15356), .C2(n15243), .A(n15242), .ZN(n15244) );
  OAI221_X1 U16330 ( .B1(P3_REG3_REG_9__SCAN_IN), .B2(n15245), .C1(n15360), 
        .C2(keyinput_117), .A(n15244), .ZN(n15249) );
  OAI22_X1 U16331 ( .A1(n15261), .A2(keyinput_119), .B1(n8216), .B2(
        keyinput_118), .ZN(n15246) );
  AOI221_X1 U16332 ( .B1(n15261), .B2(keyinput_119), .C1(keyinput_118), .C2(
        n8216), .A(n15246), .ZN(n15248) );
  NOR2_X1 U16333 ( .A1(P3_REG3_REG_13__SCAN_IN), .A2(keyinput_120), .ZN(n15247) );
  AOI221_X1 U16334 ( .B1(n15249), .B2(n15248), .C1(keyinput_120), .C2(
        P3_REG3_REG_13__SCAN_IN), .A(n15247), .ZN(n15257) );
  XOR2_X1 U16335 ( .A(P3_REG3_REG_22__SCAN_IN), .B(keyinput_121), .Z(n15256)
         );
  OAI22_X1 U16336 ( .A1(P3_REG3_REG_11__SCAN_IN), .A2(keyinput_122), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(keyinput_123), .ZN(n15250) );
  AOI221_X1 U16337 ( .B1(P3_REG3_REG_11__SCAN_IN), .B2(keyinput_122), .C1(
        keyinput_123), .C2(P3_REG3_REG_2__SCAN_IN), .A(n15250), .ZN(n15255) );
  OAI22_X1 U16338 ( .A1(n15253), .A2(keyinput_124), .B1(n15252), .B2(
        keyinput_125), .ZN(n15251) );
  AOI221_X1 U16339 ( .B1(n15253), .B2(keyinput_124), .C1(keyinput_125), .C2(
        n15252), .A(n15251), .ZN(n15254) );
  OAI211_X1 U16340 ( .C1(n15257), .C2(n15256), .A(n15255), .B(n15254), .ZN(
        n15377) );
  NAND2_X1 U16341 ( .A1(keyinput_127), .A2(n15259), .ZN(n15258) );
  OAI21_X1 U16342 ( .B1(n15259), .B2(keyinput_127), .A(n15258), .ZN(n15376) );
  INV_X1 U16343 ( .A(keyinput_62), .ZN(n15372) );
  XOR2_X1 U16344 ( .A(P3_REG3_REG_22__SCAN_IN), .B(keyinput_57), .Z(n15370) );
  OAI22_X1 U16345 ( .A1(n15261), .A2(keyinput_55), .B1(P3_REG3_REG_0__SCAN_IN), 
        .B2(keyinput_54), .ZN(n15260) );
  AOI221_X1 U16346 ( .B1(n15261), .B2(keyinput_55), .C1(keyinput_54), .C2(
        P3_REG3_REG_0__SCAN_IN), .A(n15260), .ZN(n15362) );
  INV_X1 U16347 ( .A(keyinput_53), .ZN(n15359) );
  INV_X1 U16348 ( .A(keyinput_52), .ZN(n15357) );
  INV_X1 U16349 ( .A(keyinput_51), .ZN(n15353) );
  OAI22_X1 U16350 ( .A1(P3_REG3_REG_21__SCAN_IN), .A2(keyinput_45), .B1(
        keyinput_46), .B2(P3_REG3_REG_12__SCAN_IN), .ZN(n15262) );
  AOI221_X1 U16351 ( .B1(P3_REG3_REG_21__SCAN_IN), .B2(keyinput_45), .C1(
        P3_REG3_REG_12__SCAN_IN), .C2(keyinput_46), .A(n15262), .ZN(n15351) );
  OAI22_X1 U16352 ( .A1(n15264), .A2(keyinput_48), .B1(keyinput_49), .B2(
        P3_REG3_REG_5__SCAN_IN), .ZN(n15263) );
  AOI221_X1 U16353 ( .B1(n15264), .B2(keyinput_48), .C1(P3_REG3_REG_5__SCAN_IN), .C2(keyinput_49), .A(n15263), .ZN(n15350) );
  INV_X1 U16354 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n15266) );
  OAI22_X1 U16355 ( .A1(n15267), .A2(keyinput_47), .B1(n15266), .B2(
        keyinput_50), .ZN(n15265) );
  AOI221_X1 U16356 ( .B1(n15267), .B2(keyinput_47), .C1(keyinput_50), .C2(
        n15266), .A(n15265), .ZN(n15349) );
  OAI22_X1 U16357 ( .A1(n8181), .A2(keyinput_42), .B1(n15269), .B2(keyinput_43), .ZN(n15268) );
  AOI221_X1 U16358 ( .B1(n8181), .B2(keyinput_42), .C1(keyinput_43), .C2(
        n15269), .A(n15268), .ZN(n15346) );
  OAI22_X1 U16359 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(keyinput_39), .B1(
        keyinput_40), .B2(P3_REG3_REG_3__SCAN_IN), .ZN(n15270) );
  AOI221_X1 U16360 ( .B1(P3_REG3_REG_10__SCAN_IN), .B2(keyinput_39), .C1(
        P3_REG3_REG_3__SCAN_IN), .C2(keyinput_40), .A(n15270), .ZN(n15343) );
  AOI22_X1 U16361 ( .A1(n15272), .A2(keyinput_36), .B1(keyinput_34), .B2(
        P3_U3151), .ZN(n15271) );
  OAI221_X1 U16362 ( .B1(n15272), .B2(keyinput_36), .C1(P3_U3151), .C2(
        keyinput_34), .A(n15271), .ZN(n15341) );
  INV_X1 U16363 ( .A(P3_RD_REG_SCAN_IN), .ZN(n15824) );
  AOI22_X1 U16364 ( .A1(n15824), .A2(keyinput_33), .B1(n9657), .B2(keyinput_32), .ZN(n15273) );
  OAI221_X1 U16365 ( .B1(n15824), .B2(keyinput_33), .C1(n9657), .C2(
        keyinput_32), .A(n15273), .ZN(n15336) );
  AOI22_X1 U16366 ( .A1(SI_5_), .A2(keyinput_27), .B1(n15275), .B2(keyinput_21), .ZN(n15274) );
  OAI221_X1 U16367 ( .B1(SI_5_), .B2(keyinput_27), .C1(n15275), .C2(
        keyinput_21), .A(n15274), .ZN(n15333) );
  AOI22_X1 U16368 ( .A1(SI_2_), .A2(keyinput_30), .B1(SI_3_), .B2(keyinput_29), 
        .ZN(n15276) );
  OAI221_X1 U16369 ( .B1(SI_2_), .B2(keyinput_30), .C1(SI_3_), .C2(keyinput_29), .A(n15276), .ZN(n15332) );
  AOI22_X1 U16370 ( .A1(SI_7_), .A2(keyinput_25), .B1(n15278), .B2(keyinput_26), .ZN(n15277) );
  OAI221_X1 U16371 ( .B1(SI_7_), .B2(keyinput_25), .C1(n15278), .C2(
        keyinput_26), .A(n15277), .ZN(n15329) );
  INV_X1 U16372 ( .A(keyinput_18), .ZN(n15316) );
  INV_X1 U16373 ( .A(keyinput_17), .ZN(n15312) );
  INV_X1 U16374 ( .A(keyinput_16), .ZN(n15309) );
  XNOR2_X1 U16375 ( .A(SI_21_), .B(keyinput_11), .ZN(n15307) );
  INV_X1 U16376 ( .A(keyinput_10), .ZN(n15298) );
  INV_X1 U16377 ( .A(keyinput_9), .ZN(n15295) );
  OAI22_X1 U16378 ( .A1(SI_26_), .A2(keyinput_6), .B1(keyinput_7), .B2(SI_25_), 
        .ZN(n15279) );
  AOI221_X1 U16379 ( .B1(SI_26_), .B2(keyinput_6), .C1(SI_25_), .C2(keyinput_7), .A(n15279), .ZN(n15291) );
  OAI22_X1 U16380 ( .A1(n15281), .A2(keyinput_4), .B1(SI_29_), .B2(keyinput_3), 
        .ZN(n15280) );
  AOI221_X1 U16381 ( .B1(n15281), .B2(keyinput_4), .C1(keyinput_3), .C2(SI_29_), .A(n15280), .ZN(n15287) );
  INV_X1 U16382 ( .A(keyinput_2), .ZN(n15285) );
  AOI22_X1 U16383 ( .A1(P3_WR_REG_SCAN_IN), .A2(keyinput_0), .B1(SI_31_), .B2(
        keyinput_1), .ZN(n15282) );
  OAI221_X1 U16384 ( .B1(P3_WR_REG_SCAN_IN), .B2(keyinput_0), .C1(SI_31_), 
        .C2(keyinput_1), .A(n15282), .ZN(n15283) );
  OAI221_X1 U16385 ( .B1(SI_30_), .B2(n15285), .C1(n15284), .C2(keyinput_2), 
        .A(n15283), .ZN(n15286) );
  AOI22_X1 U16386 ( .A1(keyinput_5), .A2(n15289), .B1(n15287), .B2(n15286), 
        .ZN(n15288) );
  OAI21_X1 U16387 ( .B1(n15289), .B2(keyinput_5), .A(n15288), .ZN(n15290) );
  AOI22_X1 U16388 ( .A1(n15291), .A2(n15290), .B1(keyinput_8), .B2(SI_24_), 
        .ZN(n15292) );
  OAI21_X1 U16389 ( .B1(keyinput_8), .B2(SI_24_), .A(n15292), .ZN(n15293) );
  OAI221_X1 U16390 ( .B1(SI_23_), .B2(n15295), .C1(n15294), .C2(keyinput_9), 
        .A(n15293), .ZN(n15296) );
  OAI221_X1 U16391 ( .B1(SI_22_), .B2(n15298), .C1(n15297), .C2(keyinput_10), 
        .A(n15296), .ZN(n15306) );
  AOI22_X1 U16392 ( .A1(n15301), .A2(keyinput_15), .B1(n15300), .B2(
        keyinput_14), .ZN(n15299) );
  OAI221_X1 U16393 ( .B1(n15301), .B2(keyinput_15), .C1(n15300), .C2(
        keyinput_14), .A(n15299), .ZN(n15305) );
  AOI22_X1 U16394 ( .A1(SI_20_), .A2(keyinput_12), .B1(n15303), .B2(
        keyinput_13), .ZN(n15302) );
  OAI221_X1 U16395 ( .B1(SI_20_), .B2(keyinput_12), .C1(n15303), .C2(
        keyinput_13), .A(n15302), .ZN(n15304) );
  AOI211_X1 U16396 ( .C1(n15307), .C2(n15306), .A(n15305), .B(n15304), .ZN(
        n15308) );
  AOI221_X1 U16397 ( .B1(SI_16_), .B2(keyinput_16), .C1(n15310), .C2(n15309), 
        .A(n15308), .ZN(n15311) );
  AOI221_X1 U16398 ( .B1(SI_15_), .B2(keyinput_17), .C1(n15313), .C2(n15312), 
        .A(n15311), .ZN(n15314) );
  AOI221_X1 U16399 ( .B1(SI_14_), .B2(n15316), .C1(n15315), .C2(keyinput_18), 
        .A(n15314), .ZN(n15327) );
  AOI22_X1 U16400 ( .A1(SI_12_), .A2(keyinput_20), .B1(n15318), .B2(
        keyinput_19), .ZN(n15317) );
  OAI221_X1 U16401 ( .B1(SI_12_), .B2(keyinput_20), .C1(n15318), .C2(
        keyinput_19), .A(n15317), .ZN(n15326) );
  OAI22_X1 U16402 ( .A1(n15321), .A2(keyinput_22), .B1(n15320), .B2(
        keyinput_23), .ZN(n15319) );
  AOI221_X1 U16403 ( .B1(n15321), .B2(keyinput_22), .C1(keyinput_23), .C2(
        n15320), .A(n15319), .ZN(n15325) );
  OAI22_X1 U16404 ( .A1(n15323), .A2(keyinput_28), .B1(n8049), .B2(keyinput_31), .ZN(n15322) );
  AOI221_X1 U16405 ( .B1(n15323), .B2(keyinput_28), .C1(keyinput_31), .C2(
        n8049), .A(n15322), .ZN(n15324) );
  OAI211_X1 U16406 ( .C1(n15327), .C2(n15326), .A(n15325), .B(n15324), .ZN(
        n15328) );
  AOI211_X1 U16407 ( .C1(keyinput_24), .C2(SI_8_), .A(n15329), .B(n15328), 
        .ZN(n15330) );
  OAI21_X1 U16408 ( .B1(keyinput_24), .B2(SI_8_), .A(n15330), .ZN(n15331) );
  NOR3_X1 U16409 ( .A1(n15333), .A2(n15332), .A3(n15331), .ZN(n15335) );
  NAND2_X1 U16410 ( .A1(keyinput_35), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n15334)
         );
  OAI221_X1 U16411 ( .B1(n15336), .B2(n15335), .C1(keyinput_35), .C2(
        P3_REG3_REG_7__SCAN_IN), .A(n15334), .ZN(n15340) );
  OAI22_X1 U16412 ( .A1(n15338), .A2(keyinput_38), .B1(keyinput_37), .B2(
        P3_REG3_REG_14__SCAN_IN), .ZN(n15337) );
  AOI221_X1 U16413 ( .B1(n15338), .B2(keyinput_38), .C1(
        P3_REG3_REG_14__SCAN_IN), .C2(keyinput_37), .A(n15337), .ZN(n15339) );
  OAI21_X1 U16414 ( .B1(n15341), .B2(n15340), .A(n15339), .ZN(n15342) );
  AOI22_X1 U16415 ( .A1(n15343), .A2(n15342), .B1(keyinput_41), .B2(
        P3_REG3_REG_19__SCAN_IN), .ZN(n15344) );
  OAI21_X1 U16416 ( .B1(keyinput_41), .B2(P3_REG3_REG_19__SCAN_IN), .A(n15344), 
        .ZN(n15345) );
  AOI22_X1 U16417 ( .A1(n15346), .A2(n15345), .B1(keyinput_44), .B2(
        P3_REG3_REG_1__SCAN_IN), .ZN(n15347) );
  OAI21_X1 U16418 ( .B1(keyinput_44), .B2(P3_REG3_REG_1__SCAN_IN), .A(n15347), 
        .ZN(n15348) );
  NAND4_X1 U16419 ( .A1(n15351), .A2(n15350), .A3(n15349), .A4(n15348), .ZN(
        n15352) );
  OAI221_X1 U16420 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(keyinput_51), .C1(
        n15354), .C2(n15353), .A(n15352), .ZN(n15355) );
  OAI221_X1 U16421 ( .B1(P3_REG3_REG_4__SCAN_IN), .B2(n15357), .C1(n15356), 
        .C2(keyinput_52), .A(n15355), .ZN(n15358) );
  OAI221_X1 U16422 ( .B1(P3_REG3_REG_9__SCAN_IN), .B2(keyinput_53), .C1(n15360), .C2(n15359), .A(n15358), .ZN(n15361) );
  AOI22_X1 U16423 ( .A1(n15362), .A2(n15361), .B1(keyinput_56), .B2(
        P3_REG3_REG_13__SCAN_IN), .ZN(n15363) );
  OAI21_X1 U16424 ( .B1(keyinput_56), .B2(P3_REG3_REG_13__SCAN_IN), .A(n15363), 
        .ZN(n15369) );
  INV_X1 U16425 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n15365) );
  AOI22_X1 U16426 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(keyinput_60), .B1(n15365), .B2(keyinput_58), .ZN(n15364) );
  OAI221_X1 U16427 ( .B1(P3_REG3_REG_18__SCAN_IN), .B2(keyinput_60), .C1(
        n15365), .C2(keyinput_58), .A(n15364), .ZN(n15368) );
  AOI22_X1 U16428 ( .A1(P3_REG3_REG_2__SCAN_IN), .A2(keyinput_59), .B1(
        P3_REG3_REG_6__SCAN_IN), .B2(keyinput_61), .ZN(n15366) );
  OAI221_X1 U16429 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(keyinput_59), .C1(
        P3_REG3_REG_6__SCAN_IN), .C2(keyinput_61), .A(n15366), .ZN(n15367) );
  AOI211_X1 U16430 ( .C1(n15370), .C2(n15369), .A(n15368), .B(n15367), .ZN(
        n15371) );
  AOI221_X1 U16431 ( .B1(P3_REG3_REG_26__SCAN_IN), .B2(n15372), .C1(n15162), 
        .C2(keyinput_62), .A(n15371), .ZN(n15374) );
  XOR2_X1 U16432 ( .A(keyinput_127), .B(keyinput_63), .Z(n15373) );
  NOR2_X1 U16433 ( .A1(n15374), .A2(n15373), .ZN(n15375) );
  AOI211_X1 U16434 ( .C1(n15378), .C2(n15377), .A(n15376), .B(n15375), .ZN(
        n15379) );
  MUX2_X1 U16435 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15380), .S(n16017), .Z(
        n15381) );
  AOI21_X1 U16436 ( .B1(n10105), .B2(n15382), .A(n15381), .ZN(n15383) );
  INV_X1 U16437 ( .A(n15383), .ZN(P1_U3526) );
  INV_X1 U16438 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n15385) );
  MUX2_X1 U16439 ( .A(n15385), .B(n15384), .S(n16017), .Z(n15386) );
  MUX2_X1 U16440 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15388), .S(n16017), .Z(
        P1_U3522) );
  MUX2_X1 U16441 ( .A(n15390), .B(n15389), .S(n16017), .Z(n15391) );
  OAI21_X1 U16442 ( .B1(n15392), .B2(n15402), .A(n15391), .ZN(P1_U3521) );
  MUX2_X1 U16443 ( .A(n15394), .B(n15393), .S(n16017), .Z(n15395) );
  OAI21_X1 U16444 ( .B1(n7668), .B2(n15402), .A(n15395), .ZN(P1_U3520) );
  MUX2_X1 U16445 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15396), .S(n16017), .Z(
        P1_U3519) );
  MUX2_X1 U16446 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15397), .S(n16017), .Z(
        P1_U3518) );
  MUX2_X1 U16447 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15398), .S(n16017), .Z(
        P1_U3517) );
  MUX2_X1 U16448 ( .A(n15400), .B(n15399), .S(n16017), .Z(n15401) );
  OAI21_X1 U16449 ( .B1(n15403), .B2(n15402), .A(n15401), .ZN(P1_U3516) );
  MUX2_X1 U16450 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15404), .S(n16017), .Z(
        P1_U3515) );
  MUX2_X1 U16451 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15405), .S(n16017), .Z(
        n15406) );
  AOI21_X1 U16452 ( .B1(n10105), .B2(n15407), .A(n15406), .ZN(n15408) );
  INV_X1 U16453 ( .A(n15408), .ZN(P1_U3513) );
  MUX2_X1 U16454 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15409), .S(n16017), .Z(
        P1_U3510) );
  MUX2_X1 U16455 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15410), .S(n16017), .Z(
        P1_U3507) );
  MUX2_X1 U16456 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15411), .S(n16017), .Z(
        n15412) );
  AOI21_X1 U16457 ( .B1(n10105), .B2(n15413), .A(n15412), .ZN(n15414) );
  INV_X1 U16458 ( .A(n15414), .ZN(P1_U3504) );
  INV_X1 U16459 ( .A(n15415), .ZN(n15417) );
  MUX2_X1 U16461 ( .A(n15418), .B(P1_D_REG_1__SCAN_IN), .S(n7155), .Z(P1_U3446) );
  MUX2_X1 U16462 ( .A(n15419), .B(P1_D_REG_0__SCAN_IN), .S(n7155), .Z(P1_U3445) );
  INV_X1 U16463 ( .A(n12861), .ZN(n15425) );
  NOR4_X1 U16464 ( .A1(n15421), .A2(P1_IR_REG_30__SCAN_IN), .A3(n15420), .A4(
        P1_U3086), .ZN(n15422) );
  AOI21_X1 U16465 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n15423), .A(n15422), 
        .ZN(n15424) );
  OAI21_X1 U16466 ( .B1(n15425), .B2(n15437), .A(n15424), .ZN(P1_U3324) );
  OAI222_X1 U16467 ( .A1(n15437), .A2(n15427), .B1(P1_U3086), .B2(n9610), .C1(
        n15426), .C2(n15435), .ZN(P1_U3325) );
  INV_X1 U16468 ( .A(n15428), .ZN(n15430) );
  OAI222_X1 U16469 ( .A1(n15435), .A2(n15431), .B1(n15437), .B2(n15430), .C1(
        P1_U3086), .C2(n15429), .ZN(P1_U3327) );
  OAI222_X1 U16470 ( .A1(n15435), .A2(n15434), .B1(n15437), .B2(n15433), .C1(
        P1_U3086), .C2(n15432), .ZN(P1_U3328) );
  OAI222_X1 U16471 ( .A1(P1_U3086), .A2(n15438), .B1(n15437), .B2(n15436), 
        .C1(n8134), .C2(n15435), .ZN(P1_U3329) );
  NAND2_X1 U16472 ( .A1(n14418), .A2(n15439), .ZN(n15441) );
  OAI211_X1 U16473 ( .C1(n15442), .C2(n15435), .A(n15441), .B(n15440), .ZN(
        P1_U3332) );
  MUX2_X1 U16474 ( .A(n15444), .B(n15443), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16475 ( .A(n15445), .ZN(n15446) );
  MUX2_X1 U16476 ( .A(n15446), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AND2_X1 U16477 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n7155), .ZN(P1_U3323) );
  AND2_X1 U16478 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n7155), .ZN(P1_U3322) );
  AND2_X1 U16479 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n7155), .ZN(P1_U3321) );
  AND2_X1 U16480 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n7155), .ZN(P1_U3320) );
  AND2_X1 U16481 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n7155), .ZN(P1_U3319) );
  AND2_X1 U16482 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n7155), .ZN(P1_U3318) );
  AND2_X1 U16483 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n7155), .ZN(P1_U3317) );
  AND2_X1 U16484 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n7155), .ZN(P1_U3316) );
  AND2_X1 U16485 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n7155), .ZN(P1_U3315) );
  AND2_X1 U16486 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n7155), .ZN(P1_U3314) );
  AND2_X1 U16487 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n7155), .ZN(P1_U3313) );
  AND2_X1 U16488 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n7155), .ZN(P1_U3312) );
  AND2_X1 U16489 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n7155), .ZN(P1_U3311) );
  AND2_X1 U16490 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n7155), .ZN(P1_U3310) );
  AND2_X1 U16491 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n7155), .ZN(P1_U3309) );
  AND2_X1 U16492 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n7155), .ZN(P1_U3308) );
  AND2_X1 U16493 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n7155), .ZN(P1_U3307) );
  AND2_X1 U16494 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n7155), .ZN(P1_U3306) );
  AND2_X1 U16495 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n7155), .ZN(P1_U3305) );
  AND2_X1 U16496 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n7155), .ZN(P1_U3304) );
  AND2_X1 U16497 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n7155), .ZN(P1_U3303) );
  AND2_X1 U16498 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n7155), .ZN(P1_U3302) );
  AND2_X1 U16499 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n7155), .ZN(P1_U3301) );
  AND2_X1 U16500 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n7155), .ZN(P1_U3300) );
  AND2_X1 U16501 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n7155), .ZN(P1_U3299) );
  AND2_X1 U16502 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n7155), .ZN(P1_U3298) );
  AND2_X1 U16503 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n7155), .ZN(P1_U3297) );
  AND2_X1 U16504 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n7155), .ZN(P1_U3296) );
  AND2_X1 U16505 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n7155), .ZN(P1_U3295) );
  AND2_X1 U16506 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n7155), .ZN(P1_U3294) );
  AOI21_X1 U16507 ( .B1(n15449), .B2(n15452), .A(n15448), .ZN(P2_U3417) );
  AND2_X1 U16508 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15451), .ZN(P2_U3295) );
  AND2_X1 U16509 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15451), .ZN(P2_U3294) );
  AND2_X1 U16510 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15451), .ZN(P2_U3293) );
  AND2_X1 U16511 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15451), .ZN(P2_U3292) );
  AND2_X1 U16512 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15451), .ZN(P2_U3291) );
  AND2_X1 U16513 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15451), .ZN(P2_U3290) );
  AND2_X1 U16514 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15451), .ZN(P2_U3289) );
  AND2_X1 U16515 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15451), .ZN(P2_U3288) );
  AND2_X1 U16516 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15451), .ZN(P2_U3287) );
  AND2_X1 U16517 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15451), .ZN(P2_U3286) );
  AND2_X1 U16518 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15451), .ZN(P2_U3285) );
  AND2_X1 U16519 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15451), .ZN(P2_U3284) );
  AND2_X1 U16520 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15451), .ZN(P2_U3283) );
  AND2_X1 U16521 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15451), .ZN(P2_U3282) );
  AND2_X1 U16522 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15451), .ZN(P2_U3281) );
  AND2_X1 U16523 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15451), .ZN(P2_U3280) );
  AND2_X1 U16524 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15451), .ZN(P2_U3279) );
  AND2_X1 U16525 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15451), .ZN(P2_U3278) );
  AND2_X1 U16526 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15451), .ZN(P2_U3277) );
  AND2_X1 U16527 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15451), .ZN(P2_U3276) );
  AND2_X1 U16528 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15451), .ZN(P2_U3275) );
  AND2_X1 U16529 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15451), .ZN(P2_U3274) );
  AND2_X1 U16530 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15451), .ZN(P2_U3273) );
  AND2_X1 U16531 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15451), .ZN(P2_U3272) );
  AND2_X1 U16532 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15451), .ZN(P2_U3271) );
  AND2_X1 U16533 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15451), .ZN(P2_U3270) );
  AND2_X1 U16534 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15451), .ZN(P2_U3269) );
  AND2_X1 U16535 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15451), .ZN(P2_U3268) );
  AND2_X1 U16536 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15451), .ZN(P2_U3267) );
  AND2_X1 U16537 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15451), .ZN(P2_U3266) );
  NOR2_X1 U16538 ( .A1(n15501), .A2(P2_U3947), .ZN(P2_U3087) );
  NOR2_X1 U16539 ( .A1(P3_U3897), .A2(n15806), .ZN(P3_U3150) );
  INV_X1 U16540 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15453) );
  AOI22_X1 U16541 ( .A1(n15455), .A2(n15454), .B1(n15453), .B2(n15452), .ZN(
        P2_U3416) );
  AOI22_X1 U16542 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n15527), .B1(n15523), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n15459) );
  AOI22_X1 U16543 ( .A1(n15501), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n15458) );
  OAI22_X1 U16544 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n15502), .B1(n15488), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n15456) );
  OAI21_X1 U16545 ( .B1(n15456), .B2(n15521), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n15457) );
  OAI211_X1 U16546 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n15459), .A(n15458), .B(
        n15457), .ZN(P2_U3214) );
  INV_X1 U16547 ( .A(n15460), .ZN(n15475) );
  OAI21_X1 U16548 ( .B1(n15475), .B2(n15461), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15462) );
  OAI21_X1 U16549 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15462), .ZN(n15472) );
  OAI211_X1 U16550 ( .C1(n15465), .C2(n15464), .A(n15523), .B(n15463), .ZN(
        n15471) );
  OAI211_X1 U16551 ( .C1(n15468), .C2(n15467), .A(n15527), .B(n15466), .ZN(
        n15470) );
  NAND2_X1 U16552 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n15501), .ZN(n15469) );
  NAND4_X1 U16553 ( .A1(n15472), .A2(n15471), .A3(n15470), .A4(n15469), .ZN(
        P2_U3215) );
  INV_X1 U16554 ( .A(n15473), .ZN(n15474) );
  OAI21_X1 U16555 ( .B1(n15475), .B2(n15474), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15476) );
  OAI21_X1 U16556 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15476), .ZN(n15486) );
  OAI211_X1 U16557 ( .C1(n15479), .C2(n15478), .A(n15527), .B(n15477), .ZN(
        n15485) );
  OAI211_X1 U16558 ( .C1(n15482), .C2(n15481), .A(n15523), .B(n15480), .ZN(
        n15484) );
  NAND2_X1 U16559 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(n15501), .ZN(n15483) );
  NAND4_X1 U16560 ( .A1(n15486), .A2(n15485), .A3(n15484), .A4(n15483), .ZN(
        P2_U3217) );
  INV_X1 U16561 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n15500) );
  INV_X1 U16562 ( .A(n15487), .ZN(n15491) );
  AOI211_X1 U16563 ( .C1(n15491), .C2(n15490), .A(n15489), .B(n15488), .ZN(
        n15496) );
  AOI21_X1 U16564 ( .B1(n15493), .B2(P2_REG2_REG_18__SCAN_IN), .A(n15492), 
        .ZN(n15494) );
  NOR2_X1 U16565 ( .A1(n15494), .A2(n15502), .ZN(n15495) );
  AOI211_X1 U16566 ( .C1(n15497), .C2(n15521), .A(n15496), .B(n15495), .ZN(
        n15499) );
  OAI211_X1 U16567 ( .C1(n15500), .C2(n15534), .A(n15499), .B(n15498), .ZN(
        P2_U3232) );
  AOI22_X1 U16568 ( .A1(n15501), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3088), .ZN(n15514) );
  AOI21_X1 U16569 ( .B1(n15504), .B2(n15503), .A(n15502), .ZN(n15506) );
  NAND2_X1 U16570 ( .A1(n15506), .A2(n15505), .ZN(n15513) );
  NAND2_X1 U16571 ( .A1(n15521), .A2(n15507), .ZN(n15512) );
  OAI211_X1 U16572 ( .C1(n15510), .C2(n15509), .A(n15508), .B(n15527), .ZN(
        n15511) );
  NAND4_X1 U16573 ( .A1(n15514), .A2(n15513), .A3(n15512), .A4(n15511), .ZN(
        P2_U3227) );
  INV_X1 U16574 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15664) );
  INV_X1 U16575 ( .A(n15515), .ZN(n15517) );
  NAND3_X1 U16576 ( .A1(n15518), .A2(n15517), .A3(n15516), .ZN(n15519) );
  NAND2_X1 U16577 ( .A1(n15520), .A2(n15519), .ZN(n15524) );
  AOI22_X1 U16578 ( .A1(n15524), .A2(n15523), .B1(n15522), .B2(n15521), .ZN(
        n15531) );
  AND2_X1 U16579 ( .A1(n15526), .A2(n15525), .ZN(n15528) );
  OAI21_X1 U16580 ( .B1(n15529), .B2(n15528), .A(n15527), .ZN(n15530) );
  AND2_X1 U16581 ( .A1(n15531), .A2(n15530), .ZN(n15533) );
  OAI211_X1 U16582 ( .C1(n15664), .C2(n15534), .A(n15533), .B(n15532), .ZN(
        P2_U3226) );
  INV_X1 U16583 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n15718) );
  XOR2_X1 U16584 ( .A(n15536), .B(n15535), .Z(n15541) );
  XNOR2_X1 U16585 ( .A(n15538), .B(n15537), .ZN(n15539) );
  AOI222_X1 U16586 ( .A1(n15541), .A2(n15566), .B1(n15540), .B2(n15548), .C1(
        n15539), .C2(n15558), .ZN(n15543) );
  OAI211_X1 U16587 ( .C1(n15718), .C2(n15570), .A(n15543), .B(n15542), .ZN(
        P1_U3260) );
  AOI22_X1 U16588 ( .A1(n15544), .A2(P1_ADDR_REG_18__SCAN_IN), .B1(
        P1_REG3_REG_18__SCAN_IN), .B2(P1_U3086), .ZN(n15554) );
  OAI211_X1 U16589 ( .C1(n15546), .C2(P1_REG2_REG_18__SCAN_IN), .A(n15545), 
        .B(n15558), .ZN(n15553) );
  NAND2_X1 U16590 ( .A1(n15548), .A2(n15547), .ZN(n15552) );
  OAI211_X1 U16591 ( .C1(n15550), .C2(P1_REG1_REG_18__SCAN_IN), .A(n15549), 
        .B(n15566), .ZN(n15551) );
  NAND4_X1 U16592 ( .A1(n15554), .A2(n15553), .A3(n15552), .A4(n15551), .ZN(
        P1_U3261) );
  INV_X1 U16593 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n15705) );
  XOR2_X1 U16594 ( .A(n15556), .B(n15555), .Z(n15567) );
  NAND2_X1 U16595 ( .A1(n15563), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n15557) );
  OAI21_X1 U16596 ( .B1(n15563), .B2(P1_REG2_REG_16__SCAN_IN), .A(n15557), 
        .ZN(n15560) );
  OAI211_X1 U16597 ( .C1(n15561), .C2(n15560), .A(n15559), .B(n15558), .ZN(
        n15562) );
  OAI21_X1 U16598 ( .B1(n15564), .B2(n15563), .A(n15562), .ZN(n15565) );
  AOI21_X1 U16599 ( .B1(n15567), .B2(n15566), .A(n15565), .ZN(n15569) );
  OAI211_X1 U16600 ( .C1(n15705), .C2(n15570), .A(n15569), .B(n15568), .ZN(
        P1_U3259) );
  XNOR2_X1 U16601 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15571), .ZN(SUB_1596_U53)
         );
  NAND2_X1 U16602 ( .A1(n15740), .A2(n15739), .ZN(n15572) );
  AOI21_X1 U16603 ( .B1(P2_ADDR_REG_1__SCAN_IN), .B2(n15572), .A(n15738), .ZN(
        n15579) );
  NAND2_X1 U16604 ( .A1(n15574), .A2(n15573), .ZN(n15575) );
  OAI21_X1 U16605 ( .B1(P1_ADDR_REG_1__SCAN_IN), .B2(n15576), .A(n15575), .ZN(
        n15582) );
  XNOR2_X1 U16606 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n15583) );
  XOR2_X1 U16607 ( .A(n15582), .B(n15583), .Z(n15578) );
  NAND2_X1 U16608 ( .A1(n15579), .A2(n15578), .ZN(n15580) );
  OAI21_X1 U16609 ( .B1(n15579), .B2(n15578), .A(n15580), .ZN(n15577) );
  XNOR2_X1 U16610 ( .A(n15577), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  NOR2_X1 U16611 ( .A1(n15579), .A2(n15578), .ZN(n15581) );
  OAI21_X1 U16612 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n15581), .A(n15580), .ZN(
        n15594) );
  NAND2_X1 U16613 ( .A1(n15583), .A2(n15582), .ZN(n15584) );
  XOR2_X1 U16614 ( .A(P3_ADDR_REG_3__SCAN_IN), .B(n15588), .Z(n15590) );
  XNOR2_X1 U16615 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n15590), .ZN(n15595) );
  INV_X1 U16616 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15586) );
  OAI21_X1 U16617 ( .B1(n15587), .B2(n15586), .A(n15596), .ZN(SUB_1596_U60) );
  NAND2_X1 U16618 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n15588), .ZN(n15592) );
  NAND2_X1 U16619 ( .A1(n15590), .A2(n15589), .ZN(n15591) );
  NAND2_X1 U16620 ( .A1(n15592), .A2(n15591), .ZN(n15602) );
  XNOR2_X1 U16621 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P3_ADDR_REG_4__SCAN_IN), 
        .ZN(n15593) );
  XNOR2_X1 U16622 ( .A(n15602), .B(n15593), .ZN(n15600) );
  XNOR2_X1 U16623 ( .A(n15600), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15599) );
  NAND2_X1 U16624 ( .A1(n15595), .A2(n15594), .ZN(n15597) );
  NAND2_X1 U16625 ( .A1(n15597), .A2(n15596), .ZN(n15598) );
  AOI21_X1 U16626 ( .B1(n15599), .B2(n15598), .A(n15601), .ZN(SUB_1596_U59) );
  XNOR2_X1 U16627 ( .A(P3_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n15605) );
  AND2_X1 U16628 ( .A1(n15604), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n15603) );
  XNOR2_X1 U16629 ( .A(n15605), .B(n15611), .ZN(n15607) );
  AOI21_X1 U16630 ( .B1(n15608), .B2(n15607), .A(n15609), .ZN(n15606) );
  XOR2_X1 U16631 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n15606), .Z(SUB_1596_U58) );
  XNOR2_X1 U16632 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n15613) );
  XOR2_X1 U16633 ( .A(n15613), .B(n15616), .Z(n15735) );
  NAND2_X1 U16634 ( .A1(n15736), .A2(n15735), .ZN(n15614) );
  NOR2_X1 U16635 ( .A1(n15736), .A2(n15735), .ZN(n15734) );
  XNOR2_X1 U16636 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n15625), .ZN(n15619) );
  INV_X1 U16637 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n15621) );
  AND2_X1 U16638 ( .A1(n15615), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n15617) );
  XNOR2_X1 U16639 ( .A(n15621), .B(n15620), .ZN(n15622) );
  XOR2_X1 U16640 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n15622), .Z(n15618) );
  NAND2_X1 U16641 ( .A1(n15619), .A2(n15618), .ZN(n15626) );
  OAI21_X1 U16642 ( .B1(n15619), .B2(n15618), .A(n15626), .ZN(SUB_1596_U56) );
  XNOR2_X1 U16643 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n15635) );
  NOR2_X1 U16644 ( .A1(n15621), .A2(n15620), .ZN(n15624) );
  NOR2_X1 U16645 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n15622), .ZN(n15623) );
  XOR2_X1 U16646 ( .A(n15635), .B(n15634), .Z(n15629) );
  NAND2_X1 U16647 ( .A1(n15625), .A2(n13978), .ZN(n15627) );
  NAND2_X1 U16648 ( .A1(n15629), .A2(n15628), .ZN(n15631) );
  OAI222_X1 U16649 ( .A1(n13993), .A2(n15631), .B1(n13993), .B2(n15633), .C1(
        n15630), .C2(n15632), .ZN(SUB_1596_U55) );
  NAND2_X1 U16650 ( .A1(n15635), .A2(n15634), .ZN(n15636) );
  XOR2_X1 U16651 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(n15642), .Z(n15640) );
  XNOR2_X1 U16652 ( .A(n15639), .B(n15640), .ZN(n15643) );
  AOI21_X1 U16653 ( .B1(n15644), .B2(n15643), .A(n15645), .ZN(n15638) );
  XOR2_X1 U16654 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n15638), .Z(SUB_1596_U54) );
  NAND2_X1 U16655 ( .A1(n15640), .A2(n15639), .ZN(n15641) );
  XOR2_X1 U16656 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n15648) );
  XOR2_X1 U16657 ( .A(n15649), .B(n15648), .Z(n15654) );
  NAND2_X1 U16658 ( .A1(n15644), .A2(n15643), .ZN(n15646) );
  NOR2_X1 U16659 ( .A1(n15654), .A2(n15653), .ZN(n15655) );
  AOI21_X1 U16660 ( .B1(n15654), .B2(n15653), .A(n15655), .ZN(n15647) );
  XOR2_X1 U16661 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n15647), .Z(SUB_1596_U70)
         );
  XNOR2_X1 U16662 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n15652) );
  INV_X1 U16663 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n15651) );
  XNOR2_X1 U16664 ( .A(n15652), .B(n15663), .ZN(n15658) );
  NAND2_X1 U16665 ( .A1(n15654), .A2(n15653), .ZN(n15656) );
  OAI21_X1 U16666 ( .B1(n15658), .B2(n15659), .A(n15660), .ZN(n15657) );
  XNOR2_X1 U16667 ( .A(n15657), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  XNOR2_X1 U16668 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n15667) );
  INV_X1 U16669 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n15661) );
  OR2_X1 U16670 ( .A1(n15661), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n15662) );
  XOR2_X1 U16671 ( .A(n15667), .B(n15666), .Z(n15671) );
  NAND2_X1 U16672 ( .A1(n15665), .A2(n15664), .ZN(n15672) );
  OAI21_X1 U16673 ( .B1(n15665), .B2(n15664), .A(n15672), .ZN(SUB_1596_U68) );
  NAND2_X1 U16674 ( .A1(n15667), .A2(n15666), .ZN(n15668) );
  XNOR2_X1 U16675 ( .A(n15682), .B(P1_ADDR_REG_13__SCAN_IN), .ZN(n15679) );
  XNOR2_X1 U16676 ( .A(n15680), .B(n15679), .ZN(n15676) );
  NAND2_X1 U16677 ( .A1(n15671), .A2(n15670), .ZN(n15673) );
  NAND2_X1 U16678 ( .A1(n15673), .A2(n15672), .ZN(n15675) );
  NAND2_X1 U16679 ( .A1(n15676), .A2(n15675), .ZN(n15677) );
  OAI21_X1 U16680 ( .B1(n15676), .B2(n15675), .A(n15677), .ZN(n15674) );
  XNOR2_X1 U16681 ( .A(n15674), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  NOR2_X1 U16682 ( .A1(n15676), .A2(n15675), .ZN(n15678) );
  NOR2_X1 U16683 ( .A1(n15680), .A2(n15679), .ZN(n15681) );
  AOI21_X1 U16684 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(n15682), .A(n15681), 
        .ZN(n15689) );
  NAND2_X1 U16685 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(n15691), .ZN(n15683) );
  OAI21_X1 U16686 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n15691), .A(n15683), 
        .ZN(n15688) );
  XNOR2_X1 U16687 ( .A(n15689), .B(n15688), .ZN(n15685) );
  OAI21_X1 U16688 ( .B1(n15686), .B2(n15685), .A(n15687), .ZN(n15684) );
  XNOR2_X1 U16689 ( .A(n15684), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  NOR2_X1 U16690 ( .A1(n15689), .A2(n15688), .ZN(n15690) );
  AOI21_X1 U16691 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n15691), .A(n15690), 
        .ZN(n15701) );
  INV_X1 U16692 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n15703) );
  NAND2_X1 U16693 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n15703), .ZN(n15692) );
  OAI21_X1 U16694 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n15703), .A(n15692), 
        .ZN(n15700) );
  XOR2_X1 U16695 ( .A(n15701), .B(n15700), .Z(n15693) );
  NAND2_X1 U16696 ( .A1(n15694), .A2(n15693), .ZN(n15696) );
  INV_X1 U16697 ( .A(n15695), .ZN(n15699) );
  NAND2_X1 U16698 ( .A1(n15697), .A2(n15696), .ZN(n15698) );
  OAI222_X1 U16699 ( .A1(n15697), .A2(n15696), .B1(n15697), .B2(n15699), .C1(
        n15695), .C2(n15698), .ZN(SUB_1596_U65) );
  NOR2_X1 U16700 ( .A1(n15701), .A2(n15700), .ZN(n15702) );
  AOI21_X1 U16701 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n15703), .A(n15702), 
        .ZN(n15706) );
  XOR2_X1 U16702 ( .A(n15706), .B(P1_ADDR_REG_16__SCAN_IN), .Z(n15707) );
  XNOR2_X1 U16703 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n15707), .ZN(n15710) );
  NAND2_X1 U16704 ( .A1(n15711), .A2(n15710), .ZN(n15712) );
  OAI21_X1 U16705 ( .B1(n15711), .B2(n15710), .A(n15712), .ZN(n15704) );
  XNOR2_X1 U16706 ( .A(n15704), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  NOR2_X1 U16707 ( .A1(n15706), .A2(n15705), .ZN(n15709) );
  NOR2_X1 U16708 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n15707), .ZN(n15708) );
  NOR2_X1 U16709 ( .A1(n15709), .A2(n15708), .ZN(n15719) );
  XNOR2_X1 U16710 ( .A(n15718), .B(n15719), .ZN(n15720) );
  XOR2_X1 U16711 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n15720), .Z(n15715) );
  XNOR2_X1 U16712 ( .A(n15715), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(n15714) );
  AOI21_X1 U16713 ( .B1(n15714), .B2(n15713), .A(n15716), .ZN(SUB_1596_U63) );
  AND2_X1 U16714 ( .A1(n15715), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n15717) );
  NOR2_X1 U16715 ( .A1(n15719), .A2(n15718), .ZN(n15722) );
  NOR2_X1 U16716 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n15720), .ZN(n15721) );
  NOR2_X1 U16717 ( .A1(n15722), .A2(n15721), .ZN(n15730) );
  INV_X1 U16718 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15732) );
  NAND2_X1 U16719 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n15732), .ZN(n15723) );
  OAI21_X1 U16720 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n15732), .A(n15723), 
        .ZN(n15729) );
  XNOR2_X1 U16721 ( .A(n15730), .B(n15729), .ZN(n15725) );
  NOR2_X1 U16722 ( .A1(n15726), .A2(n15725), .ZN(n15727) );
  AOI21_X1 U16723 ( .B1(n15726), .B2(n15725), .A(n15727), .ZN(n15724) );
  XOR2_X1 U16724 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n15724), .Z(SUB_1596_U62)
         );
  NAND2_X1 U16725 ( .A1(n15726), .A2(n15725), .ZN(n15728) );
  NOR2_X1 U16726 ( .A1(n15730), .A2(n15729), .ZN(n15731) );
  AOI21_X1 U16727 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n15732), .A(n15731), 
        .ZN(n15733) );
  AOI21_X1 U16728 ( .B1(n15736), .B2(n15735), .A(n15734), .ZN(n15737) );
  XOR2_X1 U16729 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n15737), .Z(SUB_1596_U57) );
  AOI21_X1 U16730 ( .B1(n15740), .B2(n15739), .A(n15738), .ZN(n15741) );
  XOR2_X1 U16731 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n15741), .Z(SUB_1596_U5) );
  NAND3_X1 U16732 ( .A1(n15800), .A2(n15742), .A3(n15763), .ZN(n15746) );
  OAI21_X1 U16733 ( .B1(P3_IR_REG_0__SCAN_IN), .B2(n15744), .A(n15743), .ZN(
        n15745) );
  NAND2_X1 U16734 ( .A1(n15746), .A2(n15745), .ZN(n15748) );
  AOI22_X1 U16735 ( .A1(n15808), .A2(P3_IR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n15747) );
  OAI211_X1 U16736 ( .C1(n15749), .C2(n15787), .A(n15748), .B(n15747), .ZN(
        P3_U3182) );
  INV_X1 U16737 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15768) );
  XOR2_X1 U16738 ( .A(n15751), .B(n15750), .Z(n15764) );
  OAI21_X1 U16739 ( .B1(n15754), .B2(n15753), .A(n15752), .ZN(n15756) );
  AOI22_X1 U16740 ( .A1(n15756), .A2(n15815), .B1(n15755), .B2(n15808), .ZN(
        n15762) );
  OAI21_X1 U16741 ( .B1(n15759), .B2(n15758), .A(n15757), .ZN(n15760) );
  NAND2_X1 U16742 ( .A1(n15760), .A2(n15819), .ZN(n15761) );
  OAI211_X1 U16743 ( .C1(n15764), .C2(n15763), .A(n15762), .B(n15761), .ZN(
        n15765) );
  INV_X1 U16744 ( .A(n15765), .ZN(n15767) );
  OAI211_X1 U16745 ( .C1(n15768), .C2(n15787), .A(n15767), .B(n15766), .ZN(
        P3_U3190) );
  INV_X1 U16746 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n15788) );
  XNOR2_X1 U16747 ( .A(n15770), .B(n15769), .ZN(n15771) );
  NAND2_X1 U16748 ( .A1(n15771), .A2(n15814), .ZN(n15784) );
  OAI21_X1 U16749 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n15773), .A(n15772), .ZN(
        n15774) );
  NAND2_X1 U16750 ( .A1(n15774), .A2(n15815), .ZN(n15783) );
  INV_X1 U16751 ( .A(n15775), .ZN(n15776) );
  NAND2_X1 U16752 ( .A1(n15776), .A2(n8331), .ZN(n15777) );
  NAND2_X1 U16753 ( .A1(n15778), .A2(n15777), .ZN(n15779) );
  NAND2_X1 U16754 ( .A1(n15779), .A2(n15819), .ZN(n15782) );
  NAND2_X1 U16755 ( .A1(n15808), .A2(n15780), .ZN(n15781) );
  AND4_X1 U16756 ( .A1(n15784), .A2(n15783), .A3(n15782), .A4(n15781), .ZN(
        n15786) );
  OAI211_X1 U16757 ( .C1(n15788), .C2(n15787), .A(n15786), .B(n15785), .ZN(
        P3_U3191) );
  AOI22_X1 U16758 ( .A1(n15808), .A2(n15789), .B1(n15806), .B2(
        P3_ADDR_REG_10__SCAN_IN), .ZN(n15805) );
  XNOR2_X1 U16759 ( .A(n15791), .B(n15790), .ZN(n15796) );
  OAI21_X1 U16760 ( .B1(n15794), .B2(n15793), .A(n15792), .ZN(n15795) );
  AOI22_X1 U16761 ( .A1(n15796), .A2(n15814), .B1(n15795), .B2(n15815), .ZN(
        n15804) );
  AOI21_X1 U16762 ( .B1(n15799), .B2(n15798), .A(n15797), .ZN(n15801) );
  OR2_X1 U16763 ( .A1(n15801), .A2(n15800), .ZN(n15802) );
  NAND4_X1 U16764 ( .A1(n15805), .A2(n15804), .A3(n15803), .A4(n15802), .ZN(
        P3_U3192) );
  AOI22_X1 U16765 ( .A1(n15808), .A2(n15807), .B1(n15806), .B2(
        P3_ADDR_REG_11__SCAN_IN), .ZN(n15823) );
  OAI21_X1 U16766 ( .B1(n15810), .B2(P3_REG2_REG_11__SCAN_IN), .A(n15809), 
        .ZN(n15816) );
  XNOR2_X1 U16767 ( .A(n15812), .B(n15811), .ZN(n15813) );
  AOI22_X1 U16768 ( .A1(n15816), .A2(n15815), .B1(n15814), .B2(n15813), .ZN(
        n15822) );
  XOR2_X1 U16769 ( .A(n15817), .B(n11799), .Z(n15818) );
  NAND2_X1 U16770 ( .A1(n15819), .A2(n15818), .ZN(n15820) );
  NAND4_X1 U16771 ( .A1(n15823), .A2(n15822), .A3(n15821), .A4(n15820), .ZN(
        P3_U3193) );
  OAI221_X1 U16772 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(n8157), .C2(n8154), .A(n15824), .ZN(U29) );
  INV_X1 U16773 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15825) );
  AOI22_X1 U16774 ( .A1(n16017), .A2(n15826), .B1(n15825), .B2(n7917), .ZN(
        P1_U3459) );
  NAND2_X1 U16775 ( .A1(n10000), .A2(n15827), .ZN(n15829) );
  AOI21_X1 U16776 ( .B1(n15830), .B2(n15829), .A(n15828), .ZN(n15833) );
  AOI22_X1 U16777 ( .A1(n15946), .A2(n15831), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n15938), .ZN(n15832) );
  OAI221_X1 U16778 ( .B1(n15895), .B2(n15833), .C1(n15054), .C2(n10356), .A(
        n15832), .ZN(P1_U3293) );
  AOI21_X1 U16779 ( .B1(n15835), .B2(n15982), .A(n15834), .ZN(n15839) );
  OAI21_X1 U16780 ( .B1(n15926), .B2(n15837), .A(n15836), .ZN(n15838) );
  AND3_X1 U16781 ( .A1(n15840), .A2(n15839), .A3(n15838), .ZN(n15841) );
  AOI22_X1 U16782 ( .A1(n16014), .A2(n15841), .B1(n9632), .B2(n7362), .ZN(
        P1_U3529) );
  AOI22_X1 U16783 ( .A1(n16017), .A2(n15841), .B1(n9637), .B2(n7917), .ZN(
        P1_U3462) );
  INV_X1 U16784 ( .A(n15842), .ZN(n15843) );
  AOI21_X1 U16785 ( .B1(n15844), .B2(n15849), .A(n15843), .ZN(n15856) );
  INV_X1 U16786 ( .A(n15856), .ZN(n15865) );
  NOR2_X1 U16787 ( .A1(n15845), .A2(n15970), .ZN(n15859) );
  AOI22_X1 U16788 ( .A1(n15848), .A2(n7349), .B1(n15847), .B2(n15846), .ZN(
        n15854) );
  XNOR2_X1 U16789 ( .A(n15850), .B(n15849), .ZN(n15852) );
  NAND2_X1 U16790 ( .A1(n15852), .A2(n15851), .ZN(n15853) );
  OAI211_X1 U16791 ( .C1(n15856), .C2(n15855), .A(n15854), .B(n15853), .ZN(
        n15863) );
  AOI211_X1 U16792 ( .C1(n15857), .C2(n15865), .A(n15859), .B(n15863), .ZN(
        n15858) );
  AOI22_X1 U16793 ( .A1(n16039), .A2(n15858), .B1(n8201), .B2(n8727), .ZN(
        P3_U3461) );
  AOI22_X1 U16794 ( .A1(n16042), .A2(n15858), .B1(n8202), .B2(n16048), .ZN(
        P3_U3396) );
  INV_X1 U16795 ( .A(n15859), .ZN(n15862) );
  OAI22_X1 U16796 ( .A1(n15862), .A2(n15861), .B1(n8203), .B2(n15860), .ZN(
        n15864) );
  AOI211_X1 U16797 ( .C1(n15866), .C2(n15865), .A(n15864), .B(n15863), .ZN(
        n15868) );
  AOI22_X1 U16798 ( .A1(n15869), .A2(n10884), .B1(n15868), .B2(n15867), .ZN(
        P3_U3231) );
  XOR2_X1 U16799 ( .A(n15870), .B(n15873), .Z(n15889) );
  OAI21_X1 U16800 ( .B1(n15873), .B2(n15872), .A(n15871), .ZN(n15877) );
  NOR2_X1 U16801 ( .A1(n15889), .A2(n15874), .ZN(n15875) );
  AOI211_X1 U16802 ( .C1(n16013), .C2(n15877), .A(n15876), .B(n15875), .ZN(
        n15894) );
  OAI21_X1 U16803 ( .B1(n15880), .B2(n15879), .A(n15878), .ZN(n15882) );
  NOR2_X1 U16804 ( .A1(n15882), .A2(n15881), .ZN(n15890) );
  AOI21_X1 U16805 ( .B1(n15888), .B2(n15982), .A(n15890), .ZN(n15883) );
  OAI211_X1 U16806 ( .C1(n15889), .C2(n15884), .A(n15894), .B(n15883), .ZN(
        n15885) );
  INV_X1 U16807 ( .A(n15885), .ZN(n15886) );
  AOI22_X1 U16808 ( .A1(n16014), .A2(n15886), .B1(n10342), .B2(n7362), .ZN(
        P1_U3530) );
  AOI22_X1 U16809 ( .A1(n16017), .A2(n15886), .B1(n9619), .B2(n7917), .ZN(
        P1_U3465) );
  AOI222_X1 U16810 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n15895), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n15938), .C1(n15888), .C2(n15887), .ZN(
        n15893) );
  INV_X1 U16811 ( .A(n15889), .ZN(n15891) );
  AOI22_X1 U16812 ( .A1(n15891), .A2(n15946), .B1(n15935), .B2(n15890), .ZN(
        n15892) );
  OAI211_X1 U16813 ( .C1(n15895), .C2(n15894), .A(n15893), .B(n15892), .ZN(
        P1_U3291) );
  INV_X1 U16814 ( .A(n15896), .ZN(n15901) );
  OAI21_X1 U16815 ( .B1(n15898), .B2(n16006), .A(n15897), .ZN(n15900) );
  AOI211_X1 U16816 ( .C1(n15926), .C2(n15901), .A(n15900), .B(n15899), .ZN(
        n15903) );
  AOI22_X1 U16817 ( .A1(n16014), .A2(n15903), .B1(n10344), .B2(n7362), .ZN(
        P1_U3531) );
  INV_X1 U16818 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n15902) );
  AOI22_X1 U16819 ( .A1(n16017), .A2(n15903), .B1(n15902), .B2(n7917), .ZN(
        P1_U3468) );
  AOI211_X1 U16820 ( .C1(n15907), .C2(n15906), .A(n15905), .B(n15904), .ZN(
        n15908) );
  OR2_X1 U16821 ( .A1(n15908), .A2(n8727), .ZN(n15909) );
  OAI21_X1 U16822 ( .B1(n16039), .B2(n15910), .A(n15909), .ZN(P3_U3463) );
  NAND2_X1 U16823 ( .A1(n15911), .A2(n15935), .ZN(n15915) );
  INV_X1 U16824 ( .A(n15912), .ZN(n15913) );
  AOI22_X1 U16825 ( .A1(n15895), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n15913), 
        .B2(n15938), .ZN(n15914) );
  OAI211_X1 U16826 ( .C1(n15916), .C2(n15942), .A(n15915), .B(n15914), .ZN(
        n15917) );
  AOI21_X1 U16827 ( .B1(n15946), .B2(n15918), .A(n15917), .ZN(n15919) );
  OAI21_X1 U16828 ( .B1(n15895), .B2(n15920), .A(n15919), .ZN(P1_U3288) );
  INV_X1 U16829 ( .A(n15921), .ZN(n15922) );
  OAI21_X1 U16830 ( .B1(n7659), .B2(n16006), .A(n15922), .ZN(n15923) );
  AOI211_X1 U16831 ( .C1(n15926), .C2(n15925), .A(n15924), .B(n15923), .ZN(
        n15928) );
  AOI22_X1 U16832 ( .A1(n16014), .A2(n15928), .B1(n10383), .B2(n7362), .ZN(
        P1_U3536) );
  INV_X1 U16833 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15927) );
  AOI22_X1 U16834 ( .A1(n16017), .A2(n15928), .B1(n15927), .B2(n7917), .ZN(
        P1_U3483) );
  OAI22_X1 U16835 ( .A1(n15930), .A2(n15972), .B1(n15929), .B2(n15970), .ZN(
        n15931) );
  NOR2_X1 U16836 ( .A1(n15932), .A2(n15931), .ZN(n15934) );
  AOI22_X1 U16837 ( .A1(n16039), .A2(n15934), .B1(n8331), .B2(n8727), .ZN(
        P3_U3468) );
  INV_X1 U16838 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15933) );
  AOI22_X1 U16839 ( .A1(n16042), .A2(n15934), .B1(n15933), .B2(n16048), .ZN(
        P3_U3417) );
  NAND2_X1 U16840 ( .A1(n15936), .A2(n15935), .ZN(n15941) );
  INV_X1 U16841 ( .A(n15937), .ZN(n15939) );
  AOI22_X1 U16842 ( .A1(n15895), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n15939), 
        .B2(n15938), .ZN(n15940) );
  OAI211_X1 U16843 ( .C1(n15943), .C2(n15942), .A(n15941), .B(n15940), .ZN(
        n15944) );
  AOI21_X1 U16844 ( .B1(n15946), .B2(n15945), .A(n15944), .ZN(n15947) );
  OAI21_X1 U16845 ( .B1(n15895), .B2(n15948), .A(n15947), .ZN(P1_U3284) );
  INV_X1 U16846 ( .A(n15949), .ZN(n15954) );
  OAI21_X1 U16847 ( .B1(n15951), .B2(n16029), .A(n15950), .ZN(n15953) );
  AOI211_X1 U16848 ( .C1(n16024), .C2(n15954), .A(n15953), .B(n15952), .ZN(
        n15956) );
  AOI22_X1 U16849 ( .A1(n16035), .A2(n15956), .B1(n10516), .B2(n16034), .ZN(
        P2_U3508) );
  INV_X1 U16850 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n15955) );
  AOI22_X1 U16851 ( .A1(n14398), .A2(n15956), .B1(n15955), .B2(n16001), .ZN(
        P2_U3457) );
  OAI22_X1 U16852 ( .A1(n15958), .A2(n15972), .B1(n15957), .B2(n15970), .ZN(
        n15959) );
  NOR2_X1 U16853 ( .A1(n15960), .A2(n15959), .ZN(n15962) );
  AOI22_X1 U16854 ( .A1(n16039), .A2(n15962), .B1(n8356), .B2(n8727), .ZN(
        P3_U3469) );
  INV_X1 U16855 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15961) );
  AOI22_X1 U16856 ( .A1(n16042), .A2(n15962), .B1(n15961), .B2(n16048), .ZN(
        P3_U3420) );
  AND2_X1 U16857 ( .A1(n15963), .A2(n16033), .ZN(n15967) );
  OAI21_X1 U16858 ( .B1(n15965), .B2(n16029), .A(n15964), .ZN(n15966) );
  NOR3_X1 U16859 ( .A1(n15968), .A2(n15967), .A3(n15966), .ZN(n15969) );
  AOI22_X1 U16860 ( .A1(n16035), .A2(n15969), .B1(n11138), .B2(n16034), .ZN(
        P2_U3510) );
  AOI22_X1 U16861 ( .A1(n14398), .A2(n15969), .B1(n9042), .B2(n16001), .ZN(
        P2_U3463) );
  OAI22_X1 U16862 ( .A1(n15973), .A2(n15972), .B1(n15971), .B2(n15970), .ZN(
        n15975) );
  AOI211_X1 U16863 ( .C1(n15977), .C2(n15976), .A(n15975), .B(n15974), .ZN(
        n15979) );
  AOI22_X1 U16864 ( .A1(n16039), .A2(n15979), .B1(n15978), .B2(n8727), .ZN(
        P3_U3471) );
  AOI22_X1 U16865 ( .A1(n16042), .A2(n15979), .B1(n8383), .B2(n16048), .ZN(
        P3_U3426) );
  INV_X1 U16866 ( .A(n15980), .ZN(n15981) );
  AOI21_X1 U16867 ( .B1(n15983), .B2(n15982), .A(n15981), .ZN(n15984) );
  OAI21_X1 U16868 ( .B1(n15986), .B2(n15985), .A(n15984), .ZN(n15990) );
  NOR2_X1 U16869 ( .A1(n15988), .A2(n15987), .ZN(n15989) );
  AOI211_X1 U16870 ( .C1(n15992), .C2(n15991), .A(n15990), .B(n15989), .ZN(
        n15994) );
  AOI22_X1 U16871 ( .A1(n16014), .A2(n15994), .B1(n9805), .B2(n7362), .ZN(
        P1_U3541) );
  INV_X1 U16872 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n15993) );
  AOI22_X1 U16873 ( .A1(n16017), .A2(n15994), .B1(n15993), .B2(n7917), .ZN(
        P1_U3498) );
  INV_X1 U16874 ( .A(n15995), .ZN(n16000) );
  OAI21_X1 U16875 ( .B1(n15997), .B2(n16029), .A(n15996), .ZN(n15999) );
  AOI211_X1 U16876 ( .C1(n16024), .C2(n16000), .A(n15999), .B(n15998), .ZN(
        n16003) );
  AOI22_X1 U16877 ( .A1(n16035), .A2(n16003), .B1(n11144), .B2(n16034), .ZN(
        P2_U3512) );
  INV_X1 U16878 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n16002) );
  AOI22_X1 U16879 ( .A1(n14398), .A2(n16003), .B1(n16002), .B2(n16001), .ZN(
        P2_U3469) );
  OAI211_X1 U16880 ( .C1(n16007), .C2(n16006), .A(n16005), .B(n16004), .ZN(
        n16011) );
  NOR2_X1 U16881 ( .A1(n16009), .A2(n16008), .ZN(n16010) );
  AOI211_X1 U16882 ( .C1(n16013), .C2(n16012), .A(n16011), .B(n16010), .ZN(
        n16016) );
  AOI22_X1 U16883 ( .A1(n16014), .A2(n16016), .B1(n11894), .B2(n7362), .ZN(
        P1_U3542) );
  INV_X1 U16884 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n16015) );
  AOI22_X1 U16885 ( .A1(n16017), .A2(n16016), .B1(n16015), .B2(n7917), .ZN(
        P1_U3501) );
  INV_X1 U16886 ( .A(n16018), .ZN(n16023) );
  OAI21_X1 U16887 ( .B1(n16020), .B2(n16029), .A(n16019), .ZN(n16022) );
  AOI211_X1 U16888 ( .C1(n16024), .C2(n16023), .A(n16022), .B(n16021), .ZN(
        n16026) );
  AOI22_X1 U16889 ( .A1(n16035), .A2(n16026), .B1(n9144), .B2(n16034), .ZN(
        P2_U3514) );
  INV_X1 U16890 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n16025) );
  AOI22_X1 U16891 ( .A1(n14398), .A2(n16026), .B1(n16025), .B2(n16001), .ZN(
        P2_U3475) );
  OAI211_X1 U16892 ( .C1(n16030), .C2(n16029), .A(n16028), .B(n16027), .ZN(
        n16031) );
  AOI21_X1 U16893 ( .B1(n16033), .B2(n16032), .A(n16031), .ZN(n16037) );
  AOI22_X1 U16894 ( .A1(n16035), .A2(n16037), .B1(n11682), .B2(n16034), .ZN(
        P2_U3516) );
  INV_X1 U16895 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n16036) );
  AOI22_X1 U16896 ( .A1(n14398), .A2(n16037), .B1(n16036), .B2(n16001), .ZN(
        P2_U3481) );
  AOI22_X1 U16897 ( .A1(n16045), .A2(n16041), .B1(P3_REG1_REG_30__SCAN_IN), 
        .B2(n8727), .ZN(n16040) );
  INV_X1 U16898 ( .A(n16038), .ZN(n16043) );
  NAND2_X1 U16899 ( .A1(n16043), .A2(n16039), .ZN(n16046) );
  NAND2_X1 U16900 ( .A1(n16040), .A2(n16046), .ZN(P3_U3489) );
  AOI22_X1 U16901 ( .A1(n16049), .A2(n16041), .B1(P3_REG0_REG_30__SCAN_IN), 
        .B2(n16048), .ZN(n16044) );
  NAND2_X1 U16902 ( .A1(n16043), .A2(n16042), .ZN(n16051) );
  NAND2_X1 U16903 ( .A1(n16044), .A2(n16051), .ZN(P3_U3457) );
  AOI22_X1 U16904 ( .A1(n16050), .A2(n16045), .B1(P3_REG1_REG_31__SCAN_IN), 
        .B2(n8727), .ZN(n16047) );
  NAND2_X1 U16905 ( .A1(n16047), .A2(n16046), .ZN(P3_U3490) );
  AOI22_X1 U16906 ( .A1(n16050), .A2(n16049), .B1(P3_REG0_REG_31__SCAN_IN), 
        .B2(n16048), .ZN(n16052) );
  NAND2_X1 U16907 ( .A1(n16052), .A2(n16051), .ZN(P3_U3458) );
  AOI21_X1 U16908 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n16053) );
  OAI21_X1 U16909 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n16053), 
        .ZN(U28) );
  CLKBUF_X1 U7273 ( .A(n10784), .Z(n13764) );
  CLKBUF_X1 U7280 ( .A(n8215), .Z(n8567) );
  INV_X1 U7539 ( .A(n9679), .ZN(n10335) );
  AND2_X1 U8404 ( .A1(n15417), .A2(n15416), .ZN(n16058) );
endmodule

