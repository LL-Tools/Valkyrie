

module b21_C_AntiSAT_k_256_6 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, 
        keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, 
        keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, 
        keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, 
        keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, 
        keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, 
        keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, 
        keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, 
        keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, 
        keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, 
        keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, 
        keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, 
        keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, 
        keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, 
        keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, 
        keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, 
        keyinput205, keyinput206, keyinput207, keyinput208, keyinput209, 
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214, 
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219, 
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224, 
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229, 
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234, 
        keyinput235, keyinput236, keyinput237, keyinput238, keyinput239, 
        keyinput240, keyinput241, keyinput242, keyinput243, keyinput244, 
        keyinput245, keyinput246, keyinput247, keyinput248, keyinput249, 
        keyinput250, keyinput251, keyinput252, keyinput253, keyinput254, 
        keyinput255, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, 
        ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, 
        ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, 
        ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, 
        ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, 
        P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, 
        P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, 
        P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, 
        P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, 
        P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, 
        P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, 
        P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, 
        P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, 
        P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, 
        P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, 
        P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, 
        P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, 
        P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, 
        P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, 
        P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, 
        P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, 
        P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, 
        P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, 
        P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, 
        P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348;

  INV_X2 U4966 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X2 U4967 ( .A(n9840), .ZN(n9842) );
  NAND2_X1 U4968 ( .A1(n6236), .A2(n8149), .ZN(n8159) );
  INV_X1 U4969 ( .A(n5747), .ZN(n7785) );
  XNOR2_X1 U4970 ( .A(n6209), .B(P2_IR_REG_22__SCAN_IN), .ZN(n5747) );
  XNOR2_X1 U4971 ( .A(n5390), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5395) );
  INV_X1 U4972 ( .A(n8112), .ZN(n8103) );
  NAND2_X1 U4973 ( .A1(n7785), .A2(n4475), .ZN(n8112) );
  INV_X1 U4974 ( .A(n7233), .ZN(n7680) );
  OR2_X1 U4975 ( .A1(n7332), .A2(n8004), .ZN(n9798) );
  INV_X1 U4976 ( .A(n7233), .ZN(n7695) );
  OAI211_X1 U4977 ( .C1(n5241), .C2(n6323), .A(n5260), .B(n5259), .ZN(n6879)
         );
  INV_X2 U4979 ( .A(n7966), .ZN(n5791) );
  NOR2_X1 U4980 ( .A1(n7141), .A2(n4561), .ZN(n8180) );
  INV_X1 U4981 ( .A(n7302), .ZN(n6803) );
  INV_X1 U4982 ( .A(n7326), .ZN(n9866) );
  INV_X1 U4983 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5721) );
  AND2_X2 U4984 ( .A1(n6387), .A2(n6359), .ZN(n7693) );
  OR2_X1 U4985 ( .A1(n9264), .A2(n9402), .ZN(n9253) );
  AND2_X1 U4986 ( .A1(n6358), .A2(n6390), .ZN(n7616) );
  NAND2_X1 U4987 ( .A1(n5154), .A2(n5153), .ZN(n5352) );
  INV_X2 U4988 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9451) );
  AOI21_X1 U4989 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n6984), .A(n7129), .ZN(
        n7093) );
  AOI21_X1 U4990 ( .B1(n6986), .B2(P2_REG2_REG_6__SCAN_IN), .A(n7091), .ZN(
        n7159) );
  AOI21_X1 U4991 ( .B1(n6993), .B2(P2_REG2_REG_9__SCAN_IN), .A(n7181), .ZN(
        n7143) );
  OAI211_X1 U4992 ( .C1(n5792), .C2(n6326), .A(n5854), .B(n5853), .ZN(n7326)
         );
  AND4_X1 U4993 ( .A1(n5402), .A2(n5401), .A3(n5400), .A4(n5399), .ZN(n5644)
         );
  INV_X1 U4994 ( .A(n8273), .ZN(n8149) );
  OAI21_X2 U4995 ( .B1(n5225), .B2(n4877), .A(n5073), .ZN(n5233) );
  AOI21_X2 U4996 ( .B1(n6889), .B2(n6888), .A(n5802), .ZN(n6867) );
  OAI21_X2 U4997 ( .B1(n6832), .B2(n6833), .A(n5784), .ZN(n6889) );
  NOR2_X2 U4998 ( .A1(n5099), .A2(n4636), .ZN(n4635) );
  NAND2_X2 U4999 ( .A1(n4767), .A2(n4768), .ZN(n8286) );
  NAND2_X2 U5000 ( .A1(n7735), .A2(n7734), .ZN(n9144) );
  NOR2_X2 U5001 ( .A1(n7169), .A2(n4694), .ZN(n7183) );
  NOR2_X2 U5002 ( .A1(n5251), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5257) );
  NAND2_X2 U5003 ( .A1(n7387), .A2(n7386), .ZN(n7395) );
  OAI211_X2 U5004 ( .C1(n5792), .C2(n6321), .A(n5815), .B(n5814), .ZN(n7322)
         );
  INV_X8 U5005 ( .A(n6401), .ZN(n7694) );
  INV_X2 U5006 ( .A(n6407), .ZN(n6401) );
  OAI21_X2 U5007 ( .B1(n6738), .B2(n5428), .A(n8854), .ZN(n8937) );
  XNOR2_X2 U5008 ( .A(n4792), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5727) );
  BUF_X2 U5009 ( .A(n9471), .Z(n4461) );
  XNOR2_X1 U5010 ( .A(n4704), .B(P2_IR_REG_1__SCAN_IN), .ZN(n9471) );
  AND2_X1 U5011 ( .A1(n4698), .A2(n4697), .ZN(n8255) );
  AND2_X1 U5012 ( .A1(n4806), .A2(n4804), .ZN(n7347) );
  OR2_X1 U5013 ( .A1(n7070), .A2(n4544), .ZN(n4806) );
  OAI21_X1 U5014 ( .B1(n6800), .B2(n8119), .A(n6631), .ZN(n6632) );
  NAND2_X1 U5015 ( .A1(n6803), .A2(n8175), .ZN(n7984) );
  INV_X4 U5016 ( .A(n7616), .ZN(n7696) );
  CLKBUF_X3 U5017 ( .A(n5851), .Z(n7753) );
  INV_X1 U5018 ( .A(n8767), .ZN(n9732) );
  CLKBUF_X2 U5019 ( .A(n5244), .Z(n6270) );
  NOR2_X1 U5020 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n7442) );
  OR2_X1 U5021 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n5752) );
  NOR2_X2 U5022 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5235) );
  OAI22_X1 U5023 ( .A1(n9070), .A2(n9069), .B1(n5632), .B2(n5043), .ZN(n9081)
         );
  NAND2_X1 U5024 ( .A1(n4959), .A2(n4958), .ZN(n4964) );
  AOI21_X1 U5025 ( .B1(n8362), .B2(n8361), .A(n8360), .ZN(n8364) );
  AOI21_X1 U5026 ( .B1(n4779), .B2(n4781), .A(n4493), .ZN(n4777) );
  OR2_X1 U5027 ( .A1(n9167), .A2(n9168), .ZN(n9165) );
  NAND2_X1 U5028 ( .A1(n5024), .A2(n5022), .ZN(n8351) );
  NAND2_X1 U5029 ( .A1(n8398), .A2(n8088), .ZN(n8375) );
  AOI21_X1 U5030 ( .B1(n9226), .B2(n4744), .A(n4743), .ZN(n9192) );
  NOR2_X1 U5031 ( .A1(n8255), .A2(n8254), .ZN(n8264) );
  NAND2_X1 U5032 ( .A1(n5381), .A2(n5380), .ZN(n9382) );
  OR2_X1 U5033 ( .A1(n7461), .A2(n4943), .ZN(n4940) );
  NAND2_X1 U5034 ( .A1(n4622), .A2(n4993), .ZN(n8488) );
  NAND2_X1 U5035 ( .A1(n4884), .A2(n4883), .ZN(n9325) );
  NAND2_X1 U5036 ( .A1(n7606), .A2(n8045), .ZN(n8520) );
  AOI21_X1 U5037 ( .B1(n4473), .B2(n4948), .A(n4525), .ZN(n4947) );
  AND2_X1 U5038 ( .A1(n5842), .A2(n5841), .ZN(n7070) );
  NAND2_X1 U5039 ( .A1(n4680), .A2(n9879), .ZN(n9800) );
  NAND2_X2 U5040 ( .A1(n7280), .A2(n8345), .ZN(n9840) );
  AOI21_X1 U5041 ( .B1(n7337), .B2(n8120), .A(n7336), .ZN(n7338) );
  NOR2_X1 U5042 ( .A1(n9512), .A2(n9555), .ZN(n7482) );
  AND2_X1 U5043 ( .A1(n8006), .A2(n8000), .ZN(n8120) );
  NAND2_X1 U5044 ( .A1(n5286), .A2(n5285), .ZN(n5112) );
  AND2_X1 U5045 ( .A1(n4696), .A2(n4695), .ZN(n7169) );
  AOI21_X1 U5046 ( .B1(n6628), .B2(n7966), .A(n5773), .ZN(n6826) );
  OR2_X1 U5047 ( .A1(n7157), .A2(n4547), .ZN(n4696) );
  AND2_X1 U5048 ( .A1(n4833), .A2(n4690), .ZN(n6802) );
  OAI21_X1 U5049 ( .B1(n6326), .B2(n5241), .A(n4521), .ZN(n9742) );
  XNOR2_X1 U5050 ( .A(n4662), .B(n5265), .ZN(n6326) );
  NAND2_X1 U5051 ( .A1(n5749), .A2(n8151), .ZN(n4834) );
  NOR2_X1 U5052 ( .A1(n6231), .A2(n5748), .ZN(n5749) );
  INV_X1 U5053 ( .A(n6387), .ZN(n7233) );
  AND4_X1 U5054 ( .A1(n5808), .A2(n5807), .A3(n5806), .A4(n5805), .ZN(n7262)
         );
  INV_X2 U5055 ( .A(n6627), .ZN(n6625) );
  NAND2_X1 U5056 ( .A1(n4569), .A2(n5406), .ZN(n9102) );
  AND4_X1 U5057 ( .A1(n5778), .A2(n5777), .A3(n5776), .A4(n5775), .ZN(n6794)
         );
  OR2_X1 U5058 ( .A1(n5412), .A2(n4468), .ZN(n9099) );
  NAND4_X1 U5059 ( .A1(n5427), .A2(n5426), .A3(n5425), .A4(n5424), .ZN(n9097)
         );
  INV_X1 U5060 ( .A(n5644), .ZN(n9101) );
  NOR2_X2 U5061 ( .A1(n6358), .A2(n6363), .ZN(n6407) );
  OAI211_X1 U5062 ( .C1(n5793), .C2(n5074), .A(n4988), .B(n4987), .ZN(n7302)
         );
  AND4_X1 U5063 ( .A1(n5790), .A2(n5789), .A3(n5788), .A4(n5787), .ZN(n6806)
         );
  NAND2_X1 U5064 ( .A1(n4482), .A2(n5420), .ZN(n9098) );
  CLKBUF_X3 U5065 ( .A(n5809), .Z(n4467) );
  NAND2_X1 U5066 ( .A1(n5671), .A2(n5670), .ZN(n6358) );
  OAI211_X1 U5067 ( .C1(n5241), .C2(n6318), .A(n5248), .B(n5247), .ZN(n6587)
         );
  INV_X1 U5068 ( .A(n5793), .ZN(n5851) );
  NAND2_X1 U5069 ( .A1(n4835), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5740) );
  INV_X2 U5070 ( .A(n5804), .ZN(n4464) );
  NAND2_X1 U5071 ( .A1(n5745), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5746) );
  OAI211_X2 U5072 ( .C1(n5241), .C2(n6314), .A(n5227), .B(n5226), .ZN(n9042)
         );
  OAI211_X1 U5073 ( .C1(n5241), .C2(n6316), .A(n5240), .B(n5239), .ZN(n8767)
         );
  OAI21_X1 U5074 ( .B1(n5228), .B2(n6494), .A(n5231), .ZN(n6597) );
  NAND2_X1 U5075 ( .A1(n5744), .A2(n5036), .ZN(n5745) );
  INV_X1 U5076 ( .A(n6382), .ZN(n6363) );
  NAND2_X1 U5077 ( .A1(n5727), .A2(n5726), .ZN(n5804) );
  INV_X1 U5078 ( .A(n5396), .ZN(n9458) );
  AND2_X2 U5079 ( .A1(n5228), .A2(n7727), .ZN(n5234) );
  INV_X1 U5080 ( .A(n5726), .ZN(n8655) );
  NAND2_X1 U5081 ( .A1(n5724), .A2(n4793), .ZN(n5726) );
  NAND2_X1 U5082 ( .A1(n5057), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5059) );
  XNOR2_X1 U5083 ( .A(n5066), .B(n5067), .ZN(n5670) );
  MUX2_X1 U5084 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5723), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5724) );
  OR2_X1 U5085 ( .A1(n5950), .A2(n5734), .ZN(n6007) );
  OR2_X1 U5086 ( .A1(n5393), .A2(n9451), .ZN(n5390) );
  NOR2_X1 U5087 ( .A1(n9467), .A2(n6978), .ZN(n9480) );
  AND2_X1 U5088 ( .A1(n5679), .A2(n4927), .ZN(n5393) );
  NAND2_X1 U5089 ( .A1(n5387), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5678) );
  NAND2_X2 U5090 ( .A1(n7717), .A2(P1_U3084), .ZN(n9460) );
  AND2_X1 U5091 ( .A1(n4675), .A2(n4676), .ZN(n4674) );
  NOR2_X1 U5092 ( .A1(n5041), .A2(n5833), .ZN(n4476) );
  CLKBUF_X3 U5093 ( .A(n5094), .Z(n5770) );
  OR2_X1 U5094 ( .A1(n4970), .A2(n9451), .ZN(n4969) );
  AND2_X1 U5095 ( .A1(n4764), .A2(n4677), .ZN(n4676) );
  INV_X1 U5096 ( .A(n7727), .ZN(n5094) );
  NAND2_X1 U5097 ( .A1(n4494), .A2(n4474), .ZN(n5041) );
  AND2_X1 U5098 ( .A1(n5025), .A2(n4765), .ZN(n4764) );
  AND2_X1 U5099 ( .A1(n10237), .A2(n4762), .ZN(n4761) );
  AND2_X1 U5100 ( .A1(n5714), .A2(n5715), .ZN(n5025) );
  AND4_X1 U5101 ( .A1(n5743), .A2(n10206), .A3(n6229), .A4(n6212), .ZN(n4474)
         );
  AND2_X1 U5102 ( .A1(n5047), .A2(n5046), .ZN(n4974) );
  AND2_X1 U5103 ( .A1(n5713), .A2(n4766), .ZN(n4763) );
  AND2_X1 U5104 ( .A1(n5048), .A2(n5049), .ZN(n4986) );
  OR2_X1 U5105 ( .A1(n5752), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n5722) );
  AND2_X1 U5106 ( .A1(n4880), .A2(n4879), .ZN(n5055) );
  NOR2_X1 U5107 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4879) );
  NOR2_X1 U5108 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4880) );
  NOR2_X2 U5109 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5779) );
  NOR2_X1 U5110 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5053) );
  NOR2_X1 U5111 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5052) );
  NOR2_X1 U5112 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5054) );
  INV_X1 U5113 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n10206) );
  INV_X1 U5114 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5048) );
  INV_X1 U5115 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6229) );
  NOR2_X1 U5116 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5743) );
  NOR2_X1 U5117 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5690) );
  INV_X1 U5118 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5692) );
  NOR2_X1 U5119 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5716) );
  INV_X1 U5120 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5714) );
  INV_X1 U5121 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5046) );
  AND2_X1 U5122 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n7441) );
  INV_X2 U5123 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n10237) );
  NAND2_X1 U5124 ( .A1(n4797), .A2(n4796), .ZN(n6136) );
  OAI21_X2 U5125 ( .B1(n8753), .B2(n8754), .A(n8751), .ZN(n7667) );
  NOR2_X1 U5126 ( .A1(n9144), .A2(n9143), .ZN(n9142) );
  XNOR2_X2 U5127 ( .A(n7730), .B(n7729), .ZN(n7749) );
  NAND2_X2 U5128 ( .A1(n5751), .A2(n5037), .ZN(n6975) );
  AND2_X1 U5129 ( .A1(n5727), .A2(n8655), .ZN(n4462) );
  OAI22_X2 U5130 ( .A1(n7395), .A2(n7396), .B1(n9891), .B2(n7910), .ZN(n7388)
         );
  NOR2_X2 U5131 ( .A1(n7548), .A2(n8835), .ZN(n7549) );
  OAI211_X2 U5132 ( .C1(n5792), .C2(n6318), .A(n5798), .B(n5797), .ZN(n6892)
         );
  AND2_X4 U5133 ( .A1(n5725), .A2(n5726), .ZN(n5785) );
  NOR2_X1 U5134 ( .A1(n9468), .A2(n4703), .ZN(n9467) );
  INV_X2 U5135 ( .A(n5804), .ZN(n4463) );
  AND2_X1 U5136 ( .A1(n5228), .A2(n7727), .ZN(n4465) );
  AND2_X1 U5137 ( .A1(n5228), .A2(n7727), .ZN(n4466) );
  INV_X1 U5138 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n4677) );
  OR2_X1 U5139 ( .A1(n7485), .A2(n7528), .ZN(n8964) );
  INV_X1 U5140 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5140) );
  INV_X1 U5141 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5139) );
  INV_X1 U5142 ( .A(n4904), .ZN(n4903) );
  NAND2_X1 U5143 ( .A1(n9417), .A2(n10326), .ZN(n4661) );
  INV_X1 U5144 ( .A(n4986), .ZN(n4736) );
  OR2_X1 U5145 ( .A1(n8562), .A2(n8404), .ZN(n7972) );
  XNOR2_X1 U5146 ( .A(n8570), .B(n8436), .ZN(n8422) );
  NAND2_X1 U5147 ( .A1(n4918), .A2(n4481), .ZN(n4917) );
  NAND2_X1 U5148 ( .A1(n9168), .A2(n4919), .ZN(n4918) );
  INV_X1 U5149 ( .A(n8905), .ZN(n4919) );
  AOI21_X1 U5150 ( .B1(n9191), .B2(n9193), .A(n5666), .ZN(n9175) );
  NOR2_X1 U5151 ( .A1(n9382), .A2(n9185), .ZN(n5666) );
  NOR2_X1 U5152 ( .A1(n4652), .A2(n4552), .ZN(n4650) );
  INV_X2 U5153 ( .A(n5241), .ZN(n7739) );
  NAND2_X1 U5154 ( .A1(n7441), .A2(n5069), .ZN(n4669) );
  NAND2_X1 U5155 ( .A1(n7442), .A2(n5068), .ZN(n4670) );
  INV_X1 U5156 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5069) );
  OR2_X1 U5157 ( .A1(n6107), .A2(n6106), .ZN(n6108) );
  INV_X1 U5158 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5713) );
  NAND2_X1 U5159 ( .A1(n4878), .A2(n7722), .ZN(n7725) );
  OR2_X1 U5160 ( .A1(n7736), .A2(n7723), .ZN(n4878) );
  INV_X1 U5161 ( .A(n5279), .ZN(n4630) );
  INV_X1 U5162 ( .A(n5093), .ZN(n4636) );
  NAND2_X1 U5163 ( .A1(n7829), .A2(n7906), .ZN(n8035) );
  NAND2_X1 U5164 ( .A1(n5747), .A2(n8273), .ZN(n8151) );
  AOI21_X1 U5165 ( .B1(n9843), .B2(n10076), .A(n9849), .ZN(n7252) );
  INV_X1 U5166 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5735) );
  INV_X1 U5167 ( .A(n8735), .ZN(n4965) );
  NAND2_X1 U5168 ( .A1(n4584), .A2(n4505), .ZN(n9032) );
  NAND2_X1 U5169 ( .A1(n4586), .A2(n4585), .ZN(n4584) );
  NAND2_X1 U5170 ( .A1(n4756), .A2(n9252), .ZN(n4908) );
  INV_X1 U5171 ( .A(n8982), .ZN(n4722) );
  OR2_X1 U5172 ( .A1(n9328), .A2(n5523), .ZN(n5524) );
  OR2_X1 U5173 ( .A1(n7477), .A2(n5492), .ZN(n5493) );
  NOR2_X1 U5174 ( .A1(n4477), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4929) );
  NOR2_X1 U5175 ( .A1(n5251), .A2(n4740), .ZN(n4739) );
  NAND2_X1 U5176 ( .A1(n5211), .A2(n4741), .ZN(n4740) );
  INV_X1 U5177 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4741) );
  OAI21_X1 U5178 ( .B1(n5352), .B2(n5351), .A(n5159), .ZN(n5356) );
  AND2_X1 U5179 ( .A1(n5145), .A2(n5144), .ZN(n5330) );
  AOI21_X1 U5180 ( .B1(n4863), .B2(n4483), .A(n4862), .ZN(n4861) );
  AND2_X1 U5181 ( .A1(n5128), .A2(n5127), .ZN(n5308) );
  INV_X1 U5182 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5049) );
  NOR2_X1 U5183 ( .A1(n7077), .A2(n4812), .ZN(n4811) );
  INV_X1 U5184 ( .A(n5860), .ZN(n4812) );
  NAND2_X1 U5185 ( .A1(n8116), .A2(n6236), .ZN(n8155) );
  NAND2_X1 U5186 ( .A1(n4594), .A2(n8110), .ZN(n8115) );
  AND4_X1 U5187 ( .A1(n6092), .A2(n6091), .A3(n6090), .A4(n6089), .ZN(n8296)
         );
  OR3_X1 U5188 ( .A1(n7571), .A2(n7595), .A3(n7589), .ZN(n6974) );
  NOR2_X1 U5189 ( .A1(n8362), .A2(n5023), .ZN(n5022) );
  INV_X1 U5190 ( .A(n7972), .ZN(n5023) );
  AND3_X1 U5191 ( .A1(n6128), .A2(n6127), .A3(n6126), .ZN(n8377) );
  OR2_X1 U5192 ( .A1(n8394), .A2(n6178), .ZN(n6127) );
  INV_X1 U5193 ( .A(n4642), .ZN(n4641) );
  OAI21_X1 U5194 ( .B1(n4645), .B2(n4643), .A(n8422), .ZN(n4642) );
  INV_X1 U5195 ( .A(n4644), .ZN(n4643) );
  AOI21_X1 U5196 ( .B1(n4527), .B2(n4771), .A(n4769), .ZN(n4768) );
  NOR2_X1 U5197 ( .A1(n8603), .A2(n8503), .ZN(n4769) );
  NOR2_X2 U5198 ( .A1(n8516), .A2(n8606), .ZN(n8505) );
  INV_X1 U5199 ( .A(n5899), .ZN(n5809) );
  INV_X1 U5200 ( .A(n8482), .ZN(n8593) );
  NAND2_X1 U5201 ( .A1(n4674), .A2(n4476), .ZN(n6206) );
  NAND2_X1 U5202 ( .A1(n6210), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6230) );
  INV_X1 U5203 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6208) );
  XNOR2_X1 U5204 ( .A(n6230), .B(n6229), .ZN(n6352) );
  NOR2_X1 U5205 ( .A1(n4965), .A2(n4958), .ZN(n4957) );
  NOR2_X1 U5206 ( .A1(n4965), .A2(n8685), .ZN(n4963) );
  AND2_X1 U5207 ( .A1(n4969), .A2(n5067), .ZN(n4968) );
  NAND2_X1 U5208 ( .A1(n8917), .A2(n8918), .ZN(n9028) );
  AOI21_X1 U5209 ( .B1(n4917), .B2(n4921), .A(n4915), .ZN(n4914) );
  INV_X1 U5210 ( .A(n4917), .ZN(n4916) );
  AOI21_X1 U5211 ( .B1(n4898), .B2(n4899), .A(n4530), .ZN(n4896) );
  INV_X1 U5212 ( .A(n9242), .ZN(n9209) );
  OR2_X1 U5213 ( .A1(n9390), .A2(n9209), .ZN(n8926) );
  NAND2_X1 U5214 ( .A1(n4478), .A2(n4660), .ZN(n4652) );
  NAND2_X1 U5215 ( .A1(n9283), .A2(n9304), .ZN(n4660) );
  AOI21_X1 U5216 ( .B1(n4664), .B2(n4663), .A(n4885), .ZN(n9346) );
  AND2_X1 U5217 ( .A1(n8835), .A2(n9087), .ZN(n4885) );
  NAND2_X1 U5218 ( .A1(n9537), .A2(n9344), .ZN(n4663) );
  INV_X1 U5219 ( .A(n7546), .ZN(n4664) );
  OR2_X1 U5220 ( .A1(n9365), .A2(n9762), .ZN(n4667) );
  OR2_X1 U5221 ( .A1(n9004), .A2(n5632), .ZN(n9756) );
  AND2_X1 U5222 ( .A1(n5688), .A2(n5687), .ZN(n6520) );
  XNOR2_X1 U5223 ( .A(n4638), .B(n5299), .ZN(n6345) );
  NAND2_X1 U5224 ( .A1(n4639), .A2(n5116), .ZN(n4638) );
  NAND2_X1 U5225 ( .A1(n5112), .A2(n4866), .ZN(n4639) );
  NAND2_X1 U5226 ( .A1(n4849), .A2(n4850), .ZN(n5268) );
  AOI21_X1 U5227 ( .B1(n4852), .B2(n4854), .A(n4522), .ZN(n4850) );
  INV_X1 U5228 ( .A(n4853), .ZN(n4852) );
  NAND2_X1 U5229 ( .A1(n7004), .A2(n7001), .ZN(n9786) );
  NAND2_X1 U5230 ( .A1(n5217), .A2(n5216), .ZN(n7763) );
  NAND2_X1 U5231 ( .A1(n7741), .A2(n7740), .ZN(n9367) );
  NAND2_X1 U5232 ( .A1(n7996), .A2(n8000), .ZN(n4593) );
  OAI21_X1 U5233 ( .B1(n4602), .B2(n4601), .A(n5010), .ZN(n4600) );
  INV_X1 U5234 ( .A(n8039), .ZN(n4601) );
  AOI21_X1 U5235 ( .B1(n8024), .B2(n8023), .A(n4603), .ZN(n4602) );
  OAI21_X1 U5236 ( .B1(n4582), .B2(n4581), .A(n8995), .ZN(n4580) );
  INV_X1 U5237 ( .A(n8992), .ZN(n4581) );
  AOI21_X1 U5238 ( .B1(n8991), .B2(n8990), .A(n8998), .ZN(n4582) );
  AOI21_X1 U5239 ( .B1(n4578), .B2(n4470), .A(n4515), .ZN(n4576) );
  OR2_X1 U5240 ( .A1(n4574), .A2(n9011), .ZN(n4577) );
  AOI21_X1 U5241 ( .B1(n4800), .B2(n4799), .A(n4526), .ZN(n4798) );
  INV_X1 U5242 ( .A(n4563), .ZN(n4799) );
  AND2_X1 U5243 ( .A1(n5002), .A2(n8102), .ZN(n5001) );
  NAND2_X1 U5244 ( .A1(n5003), .A2(n5005), .ZN(n5002) );
  INV_X1 U5245 ( .A(n5006), .ZN(n5003) );
  INV_X1 U5246 ( .A(n5005), .ZN(n5004) );
  INV_X1 U5247 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n4765) );
  NAND2_X1 U5248 ( .A1(n4945), .A2(n4944), .ZN(n4943) );
  INV_X1 U5249 ( .A(n7463), .ZN(n4944) );
  INV_X1 U5250 ( .A(n7611), .ZN(n4945) );
  AND2_X1 U5251 ( .A1(n8704), .A2(n4938), .ZN(n4937) );
  OR2_X1 U5252 ( .A1(n4939), .A2(n8743), .ZN(n4938) );
  INV_X1 U5253 ( .A(n7655), .ZN(n4939) );
  NOR2_X1 U5254 ( .A1(n8727), .A2(n4981), .ZN(n4980) );
  INV_X1 U5255 ( .A(n4982), .ZN(n4981) );
  INV_X1 U5256 ( .A(n5382), .ZN(n4870) );
  INV_X1 U5257 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5146) );
  INV_X1 U5258 ( .A(SI_15_), .ZN(n5134) );
  INV_X1 U5259 ( .A(SI_12_), .ZN(n5118) );
  NOR2_X1 U5260 ( .A1(n4822), .A2(n4819), .ZN(n4818) );
  INV_X1 U5261 ( .A(n5949), .ZN(n4819) );
  INV_X1 U5262 ( .A(n4823), .ZN(n4822) );
  AND2_X1 U5263 ( .A1(n5963), .A2(n4824), .ZN(n4823) );
  INV_X1 U5264 ( .A(n7880), .ZN(n4824) );
  OAI211_X1 U5265 ( .C1(n4834), .C2(n7312), .A(n4830), .B(n4829), .ZN(n5758)
         );
  NAND2_X1 U5266 ( .A1(n4833), .A2(n4832), .ZN(n4829) );
  NAND2_X1 U5267 ( .A1(n4834), .A2(n4831), .ZN(n4830) );
  NOR2_X1 U5268 ( .A1(n4833), .A2(n4832), .ZN(n4831) );
  AND2_X1 U5269 ( .A1(n7968), .A2(n8098), .ZN(n5006) );
  OR2_X1 U5270 ( .A1(n8550), .A2(n8309), .ZN(n8098) );
  OR2_X1 U5271 ( .A1(n8557), .A2(n8378), .ZN(n8094) );
  OR2_X1 U5272 ( .A1(n8565), .A2(n8377), .ZN(n8088) );
  OR2_X1 U5273 ( .A1(n8581), .A2(n8294), .ZN(n8078) );
  NOR2_X1 U5274 ( .A1(n4692), .A2(n8586), .ZN(n4691) );
  INV_X1 U5275 ( .A(n4693), .ZN(n4692) );
  OR2_X1 U5276 ( .A1(n8586), .A2(n8475), .ZN(n8079) );
  OR2_X1 U5277 ( .A1(n8596), .A2(n8492), .ZN(n8064) );
  OR2_X1 U5278 ( .A1(n8603), .A2(n7918), .ZN(n8059) );
  AND2_X1 U5279 ( .A1(n5012), .A2(n5010), .ZN(n5009) );
  NOR2_X1 U5280 ( .A1(n8136), .A2(n4791), .ZN(n4790) );
  NOR2_X1 U5281 ( .A1(n9804), .A2(n5030), .ZN(n5029) );
  INV_X1 U5282 ( .A(n5031), .ZN(n5030) );
  NAND2_X1 U5283 ( .A1(n7281), .A2(n9866), .ZN(n7332) );
  OAI211_X1 U5284 ( .C1(n5793), .C2(n10091), .A(n5757), .B(n5756), .ZN(n6627)
         );
  NOR2_X1 U5285 ( .A1(n9878), .A2(n5748), .ZN(n6622) );
  INV_X1 U5286 ( .A(n5395), .ZN(n5397) );
  OR2_X1 U5287 ( .A1(n7763), .A2(n7764), .ZN(n9020) );
  OR2_X1 U5288 ( .A1(n9370), .A2(n7705), .ZN(n9018) );
  OR2_X1 U5289 ( .A1(n9206), .A2(n4746), .ZN(n4745) );
  INV_X1 U5290 ( .A(n8926), .ZN(n4746) );
  NOR2_X1 U5291 ( .A1(n9427), .A2(n9430), .ZN(n4750) );
  INV_X1 U5292 ( .A(n8939), .ZN(n5652) );
  NAND2_X1 U5293 ( .A1(n4881), .A2(n4882), .ZN(n9047) );
  NOR2_X1 U5294 ( .A1(n4468), .A2(n9732), .ZN(n4881) );
  NAND2_X1 U5295 ( .A1(n9078), .A2(n9135), .ZN(n6390) );
  NOR2_X1 U5296 ( .A1(n9042), .A2(n6597), .ZN(n6613) );
  XNOR2_X1 U5297 ( .A(n7725), .B(n7724), .ZN(n7733) );
  NAND2_X1 U5298 ( .A1(n7716), .A2(n7715), .ZN(n7736) );
  NAND2_X1 U5299 ( .A1(n7712), .A2(n7711), .ZN(n7716) );
  OAI21_X1 U5300 ( .B1(n5360), .B2(n5166), .A(n5169), .ZN(n5364) );
  INV_X1 U5301 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5058) );
  AND2_X1 U5302 ( .A1(n5164), .A2(n5163), .ZN(n5355) );
  AND2_X1 U5303 ( .A1(n4543), .A2(n5056), .ZN(n4970) );
  NAND2_X1 U5304 ( .A1(n4838), .A2(n4836), .ZN(n5338) );
  AOI21_X1 U5305 ( .B1(n4840), .B2(n4843), .A(n4837), .ZN(n4836) );
  INV_X1 U5306 ( .A(n5145), .ZN(n4837) );
  NOR2_X1 U5307 ( .A1(n5117), .A2(n4867), .ZN(n4866) );
  INV_X1 U5308 ( .A(n5111), .ZN(n4867) );
  AND2_X1 U5309 ( .A1(n5105), .A2(n5104), .ZN(n5279) );
  AOI21_X1 U5310 ( .B1(n4635), .B2(n4633), .A(n4632), .ZN(n4631) );
  INV_X1 U5311 ( .A(n5100), .ZN(n4632) );
  INV_X1 U5312 ( .A(n5267), .ZN(n4633) );
  INV_X1 U5313 ( .A(n4635), .ZN(n4634) );
  INV_X1 U5314 ( .A(n4811), .ZN(n4810) );
  INV_X1 U5315 ( .A(n6323), .ZN(n4991) );
  INV_X1 U5316 ( .A(n7268), .ZN(n4807) );
  NAND2_X1 U5317 ( .A1(n6070), .A2(n4563), .ZN(n4802) );
  NAND2_X1 U5318 ( .A1(n4802), .A2(n4800), .ZN(n7872) );
  AND2_X1 U5319 ( .A1(n5930), .A2(n7344), .ZN(n4828) );
  NAND2_X1 U5320 ( .A1(n4816), .A2(n6158), .ZN(n4815) );
  INV_X1 U5321 ( .A(n7836), .ZN(n4816) );
  NAND3_X1 U5322 ( .A1(n6143), .A2(n6142), .A3(n4503), .ZN(n4814) );
  INV_X1 U5323 ( .A(n5987), .ZN(n5985) );
  OAI21_X2 U5324 ( .B1(n5745), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6209) );
  AND4_X1 U5325 ( .A1(n5883), .A2(n5882), .A3(n5881), .A4(n5880), .ZN(n7369)
         );
  AND4_X1 U5326 ( .A1(n5850), .A2(n5849), .A3(n5848), .A4(n5847), .ZN(n7276)
         );
  AND2_X1 U5327 ( .A1(n5725), .A2(n8655), .ZN(n5786) );
  XNOR2_X1 U5328 ( .A(n4461), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n9468) );
  INV_X1 U5329 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5980) );
  OR2_X1 U5330 ( .A1(n8229), .A2(n8228), .ZN(n4698) );
  NAND2_X1 U5331 ( .A1(n4859), .A2(n4858), .ZN(n4856) );
  NAND2_X1 U5332 ( .A1(n7753), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n4858) );
  NOR2_X1 U5333 ( .A1(n8365), .A2(n4686), .ZN(n8279) );
  OR3_X1 U5334 ( .A1(n8545), .A2(n4687), .A3(n8280), .ZN(n4686) );
  NAND2_X1 U5335 ( .A1(n8331), .A2(n7968), .ZN(n5005) );
  OR2_X1 U5336 ( .A1(n6161), .A2(n7928), .ZN(n6176) );
  NAND2_X1 U5337 ( .A1(n8375), .A2(n8374), .ZN(n5024) );
  NAND2_X1 U5338 ( .A1(n8094), .A2(n8350), .ZN(n8362) );
  INV_X1 U5339 ( .A(n8303), .ZN(n8374) );
  NAND2_X1 U5340 ( .A1(n8390), .A2(n8302), .ZN(n8373) );
  AND3_X1 U5341 ( .A1(n6152), .A2(n6151), .A3(n6150), .ZN(n8404) );
  OR2_X1 U5342 ( .A1(n8383), .A2(n6178), .ZN(n6152) );
  AND2_X1 U5343 ( .A1(n8088), .A2(n8089), .ZN(n8399) );
  AND2_X1 U5344 ( .A1(n4469), .A2(n8070), .ZN(n4645) );
  NAND2_X1 U5345 ( .A1(n4519), .A2(n8070), .ZN(n4644) );
  OR3_X1 U5346 ( .A1(n6013), .A2(n6012), .A3(n6011), .ZN(n6032) );
  AND2_X1 U5347 ( .A1(n4994), .A2(n8056), .ZN(n4993) );
  NAND2_X1 U5348 ( .A1(n8520), .A2(n4992), .ZN(n4622) );
  NAND2_X1 U5349 ( .A1(n8055), .A2(n4995), .ZN(n4994) );
  INV_X1 U5350 ( .A(n4774), .ZN(n4773) );
  AOI21_X1 U5351 ( .B1(n4774), .B2(n4772), .A(n4518), .ZN(n4771) );
  AND2_X1 U5352 ( .A1(n8510), .A2(n4488), .ZN(n4774) );
  OR2_X1 U5353 ( .A1(n8612), .A2(n7849), .ZN(n8051) );
  NAND2_X1 U5354 ( .A1(n8520), .A2(n4772), .ZN(n8519) );
  OR2_X1 U5355 ( .A1(n7601), .A2(n8521), .ZN(n7602) );
  AOI21_X1 U5356 ( .B1(n5014), .B2(n7514), .A(n5013), .ZN(n5012) );
  INV_X1 U5357 ( .A(n8034), .ZN(n5013) );
  NAND2_X1 U5358 ( .A1(n7515), .A2(n5014), .ZN(n5011) );
  AND2_X1 U5359 ( .A1(n5011), .A2(n5009), .ZN(n7577) );
  NAND2_X1 U5360 ( .A1(n7512), .A2(n4790), .ZN(n4789) );
  AND2_X1 U5361 ( .A1(n8034), .A2(n8035), .ZN(n8136) );
  AND2_X1 U5362 ( .A1(n8015), .A2(n8010), .ZN(n9793) );
  INV_X1 U5363 ( .A(n8491), .ZN(n9807) );
  AND2_X1 U5364 ( .A1(n6972), .A2(n6245), .ZN(n9806) );
  AND4_X1 U5365 ( .A1(n5830), .A2(n5829), .A3(n5828), .A4(n5827), .ZN(n7287)
         );
  INV_X1 U5366 ( .A(n9806), .ZN(n8474) );
  AND2_X1 U5367 ( .A1(n7965), .A2(n8151), .ZN(n9813) );
  OR2_X1 U5368 ( .A1(n6634), .A2(n6245), .ZN(n8491) );
  NAND2_X1 U5369 ( .A1(n6145), .A2(n6144), .ZN(n8562) );
  NAND2_X1 U5370 ( .A1(n6115), .A2(n6114), .ZN(n8570) );
  INV_X1 U5371 ( .A(n8444), .ZN(n8581) );
  NAND2_X1 U5372 ( .A1(n8493), .A2(n8284), .ZN(n8478) );
  INV_X1 U5373 ( .A(n7246), .ZN(n9860) );
  AND2_X1 U5374 ( .A1(n6216), .A2(n6215), .ZN(n9843) );
  INV_X1 U5375 ( .A(n7595), .ZN(n6216) );
  NAND2_X1 U5376 ( .A1(n6974), .A2(n9850), .ZN(n9844) );
  NOR2_X1 U5377 ( .A1(n4679), .A2(n5041), .ZN(n5033) );
  NOR2_X1 U5378 ( .A1(n5041), .A2(n5034), .ZN(n5032) );
  INV_X1 U5379 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U5380 ( .A1(n6043), .A2(n5742), .ZN(n4835) );
  AND2_X1 U5381 ( .A1(n5834), .A2(n5833), .ZN(n6984) );
  NAND2_X1 U5382 ( .A1(n9102), .A2(n6407), .ZN(n6365) );
  AND2_X1 U5383 ( .A1(n6362), .A2(n6361), .ZN(n6366) );
  INV_X1 U5384 ( .A(n7039), .ZN(n4948) );
  INV_X1 U5385 ( .A(n7044), .ZN(n4949) );
  NAND2_X1 U5386 ( .A1(n4953), .A2(n4512), .ZN(n4952) );
  INV_X1 U5387 ( .A(n4961), .ZN(n4953) );
  AND2_X1 U5388 ( .A1(n4963), .A2(n4962), .ZN(n4961) );
  AND2_X1 U5389 ( .A1(n9135), .A2(n5670), .ZN(n6535) );
  NAND2_X1 U5390 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n10082), .ZN(n4934) );
  NOR2_X1 U5391 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(n5058), .ZN(n4933) );
  AND2_X1 U5392 ( .A1(n6469), .A2(n4485), .ZN(n4617) );
  NOR2_X1 U5393 ( .A1(n6817), .A2(n4606), .ZN(n6511) );
  AND2_X1 U5394 ( .A1(n6510), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4606) );
  NAND2_X1 U5395 ( .A1(n6511), .A2(n6512), .ZN(n9104) );
  NAND2_X1 U5396 ( .A1(n9618), .A2(n9106), .ZN(n9632) );
  NAND2_X1 U5397 ( .A1(n9632), .A2(n9633), .ZN(n4614) );
  OAI21_X1 U5398 ( .B1(n9664), .B2(n4608), .A(n4607), .ZN(n9672) );
  NAND2_X1 U5399 ( .A1(n4611), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4608) );
  NAND2_X1 U5400 ( .A1(n9111), .A2(n4611), .ZN(n4607) );
  INV_X1 U5401 ( .A(n9673), .ZN(n4611) );
  OR2_X1 U5402 ( .A1(n9664), .A2(n9663), .ZN(n4610) );
  NOR2_X1 U5403 ( .A1(n9683), .A2(n4621), .ZN(n9704) );
  AND2_X1 U5404 ( .A1(n9116), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4621) );
  NAND2_X1 U5405 ( .A1(n6363), .A2(n7473), .ZN(n6307) );
  OR2_X1 U5406 ( .A1(n9375), .A2(n9164), .ZN(n8904) );
  AND2_X1 U5407 ( .A1(n9375), .A2(n9164), .ZN(n8905) );
  NAND2_X1 U5408 ( .A1(n5582), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5593) );
  INV_X1 U5409 ( .A(n4745), .ZN(n4744) );
  OR2_X1 U5410 ( .A1(n9226), .A2(n9219), .ZN(n9227) );
  NAND2_X1 U5411 ( .A1(n4532), .A2(n4908), .ZN(n4904) );
  AND2_X1 U5412 ( .A1(n4908), .A2(n9248), .ZN(n4905) );
  AND2_X1 U5413 ( .A1(n8831), .A2(n8993), .ZN(n9241) );
  NOR2_X1 U5414 ( .A1(n4721), .A2(n4718), .ZN(n4717) );
  OAI21_X1 U5415 ( .B1(n4487), .B2(n4718), .A(n4716), .ZN(n4715) );
  INV_X1 U5416 ( .A(n8990), .ZN(n4718) );
  NOR2_X1 U5417 ( .A1(n4546), .A2(n4656), .ZN(n4655) );
  NOR2_X1 U5418 ( .A1(n9292), .A2(n9410), .ZN(n9280) );
  NAND2_X1 U5419 ( .A1(n4533), .A2(n4661), .ZN(n4657) );
  NAND2_X1 U5420 ( .A1(n4484), .A2(n5661), .ZN(n4659) );
  NAND2_X1 U5421 ( .A1(n4484), .A2(n4661), .ZN(n4656) );
  NAND2_X1 U5422 ( .A1(n7549), .A2(n4748), .ZN(n9292) );
  AND2_X1 U5423 ( .A1(n4472), .A2(n4749), .ZN(n4748) );
  AOI21_X1 U5424 ( .B1(n9318), .B2(n9427), .A(n9324), .ZN(n9307) );
  NOR2_X1 U5425 ( .A1(n9325), .A2(n9327), .ZN(n9324) );
  INV_X1 U5426 ( .A(n4729), .ZN(n4728) );
  AOI21_X1 U5427 ( .B1(n4729), .B2(n4727), .A(n4726), .ZN(n4725) );
  NOR2_X1 U5428 ( .A1(n7545), .A2(n4730), .ZN(n4729) );
  NAND2_X1 U5429 ( .A1(n7527), .A2(n8895), .ZN(n7526) );
  NAND2_X1 U5430 ( .A1(n4887), .A2(n4886), .ZN(n7546) );
  NOR2_X1 U5431 ( .A1(n4890), .A2(n4549), .ZN(n4886) );
  NAND2_X1 U5432 ( .A1(n4531), .A2(n4471), .ZN(n4893) );
  NAND2_X1 U5433 ( .A1(n5659), .A2(n5658), .ZN(n4895) );
  NAND2_X1 U5434 ( .A1(n4471), .A2(n5658), .ZN(n4892) );
  AND2_X1 U5435 ( .A1(n7482), .A2(n9549), .ZN(n7533) );
  AND2_X1 U5436 ( .A1(n8933), .A2(n8942), .ZN(n8939) );
  AND2_X1 U5437 ( .A1(n8885), .A2(n5649), .ZN(n4922) );
  INV_X1 U5438 ( .A(n9097), .ZN(n6732) );
  INV_X1 U5439 ( .A(n9098), .ZN(n6741) );
  AND2_X1 U5440 ( .A1(n9102), .A2(n6597), .ZN(n6604) );
  OR2_X1 U5441 ( .A1(n9036), .A2(n9572), .ZN(n9501) );
  AND2_X1 U5442 ( .A1(n7763), .A2(n9750), .ZN(n4732) );
  OAI211_X1 U5443 ( .C1(n7573), .C2(n5686), .A(n7591), .B(n5685), .ZN(n9717)
         );
  NAND2_X1 U5444 ( .A1(n7591), .A2(n5694), .ZN(n6382) );
  AND2_X1 U5445 ( .A1(n7573), .A2(n5696), .ZN(n5694) );
  NAND2_X1 U5446 ( .A1(n5394), .A2(n9452), .ZN(n5396) );
  XNOR2_X1 U5447 ( .A(n5383), .B(n5382), .ZN(n7590) );
  NAND2_X1 U5448 ( .A1(n4868), .A2(n4872), .ZN(n5383) );
  NAND2_X1 U5449 ( .A1(n5375), .A2(n4875), .ZN(n4868) );
  AND2_X1 U5450 ( .A1(n5055), .A2(n4986), .ZN(n4738) );
  INV_X1 U5451 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n10241) );
  NAND2_X1 U5452 ( .A1(n4839), .A2(n4845), .ZN(n5331) );
  NAND2_X1 U5453 ( .A1(n5314), .A2(n4847), .ZN(n4839) );
  OAI21_X1 U5454 ( .B1(n5112), .B2(n4483), .A(n4863), .ZN(n5309) );
  AND2_X1 U5455 ( .A1(n5100), .A2(n5098), .ZN(n5272) );
  AND2_X1 U5456 ( .A1(n4986), .A2(n5050), .ZN(n4985) );
  INV_X1 U5457 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5050) );
  NAND2_X1 U5458 ( .A1(n5085), .A2(n5084), .ZN(n5256) );
  INV_X1 U5459 ( .A(n5224), .ZN(n4877) );
  NAND2_X1 U5460 ( .A1(n5094), .A2(n5071), .ZN(n5229) );
  AND4_X1 U5461 ( .A1(n5973), .A2(n5972), .A3(n5971), .A4(n5970), .ZN(n8040)
         );
  AND4_X1 U5462 ( .A1(n5943), .A2(n5942), .A3(n5941), .A4(n5940), .ZN(n7828)
         );
  AOI21_X1 U5463 ( .B1(n4809), .B2(n4811), .A(n4524), .ZN(n4808) );
  INV_X1 U5464 ( .A(n7071), .ZN(n4809) );
  OR2_X1 U5465 ( .A1(n7070), .A2(n4810), .ZN(n4803) );
  NAND2_X1 U5466 ( .A1(n5953), .A2(n5952), .ZN(n7829) );
  NAND2_X1 U5467 ( .A1(n6250), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7909) );
  NAND2_X1 U5468 ( .A1(n7070), .A2(n7071), .ZN(n7069) );
  OR2_X1 U5469 ( .A1(n7929), .A2(n8491), .ZN(n7938) );
  OR2_X1 U5470 ( .A1(n8155), .A2(n5035), .ZN(n4605) );
  NAND2_X1 U5471 ( .A1(n8158), .A2(n8157), .ZN(n4626) );
  INV_X1 U5472 ( .A(n7369), .ZN(n8170) );
  INV_X1 U5473 ( .A(n7170), .ZN(n4695) );
  AOI21_X1 U5474 ( .B1(n8272), .B2(n9783), .A(n9483), .ZN(n4710) );
  OAI21_X1 U5475 ( .B1(n8277), .B2(n8278), .A(n8276), .ZN(n4712) );
  OR2_X1 U5476 ( .A1(n6206), .A2(n5752), .ZN(n5037) );
  OR2_X1 U5477 ( .A1(n6201), .A2(n5721), .ZN(n5750) );
  INV_X1 U5478 ( .A(n9086), .ZN(n9330) );
  NAND2_X1 U5479 ( .A1(n5373), .A2(n5372), .ZN(n9390) );
  XOR2_X1 U5480 ( .A(n7699), .B(n7698), .Z(n7700) );
  INV_X1 U5481 ( .A(n9088), .ZN(n7542) );
  NAND2_X1 U5482 ( .A1(n5377), .A2(n5376), .ZN(n9387) );
  INV_X1 U5483 ( .A(n6597), .ZN(n6614) );
  NAND2_X1 U5484 ( .A1(n5298), .A2(n5297), .ZN(n9555) );
  NAND2_X1 U5485 ( .A1(n6378), .A2(n9294), .ZN(n8807) );
  OR2_X1 U5486 ( .A1(n5042), .A2(n5670), .ZN(n9069) );
  NAND2_X1 U5487 ( .A1(n5581), .A2(n5580), .ZN(n9242) );
  NAND2_X1 U5488 ( .A1(n9143), .A2(n7777), .ZN(n9365) );
  AOI21_X1 U5489 ( .B1(n4914), .B2(n4916), .A(n4506), .ZN(n4911) );
  NAND2_X1 U5490 ( .A1(n4747), .A2(n7775), .ZN(n9366) );
  NAND2_X1 U5491 ( .A1(n7769), .A2(n9351), .ZN(n4747) );
  NAND2_X1 U5492 ( .A1(n4734), .A2(n5643), .ZN(n9154) );
  AOI21_X1 U5493 ( .B1(n9186), .B2(n9317), .A(n5642), .ZN(n5643) );
  NAND2_X1 U5494 ( .A1(n4735), .A2(n9351), .ZN(n4734) );
  NOR2_X1 U5495 ( .A1(n7766), .A2(n9501), .ZN(n5642) );
  INV_X1 U5496 ( .A(n9135), .ZN(n9257) );
  OAI21_X1 U5497 ( .B1(n4592), .B2(n4510), .A(n8129), .ZN(n8009) );
  AOI21_X1 U5498 ( .B1(n7991), .B2(n7990), .A(n4593), .ZN(n4592) );
  NAND2_X1 U5499 ( .A1(n8030), .A2(n8136), .ZN(n4603) );
  OAI211_X1 U5500 ( .C1(n4573), .C2(n4572), .A(n4511), .B(n4571), .ZN(n8935)
         );
  NAND2_X1 U5501 ( .A1(n8885), .A2(n6908), .ZN(n4571) );
  INV_X1 U5502 ( .A(n6908), .ZN(n4572) );
  OAI21_X1 U5503 ( .B1(n8950), .B2(n8954), .A(n8949), .ZN(n4591) );
  NAND2_X1 U5504 ( .A1(n4600), .A2(n4599), .ZN(n8048) );
  NOR2_X1 U5505 ( .A1(n8043), .A2(n8044), .ZN(n4599) );
  AOI21_X1 U5506 ( .B1(n4590), .B2(n9030), .A(n4587), .ZN(n8961) );
  NAND2_X1 U5507 ( .A1(n4589), .A2(n4588), .ZN(n4587) );
  NAND2_X1 U5508 ( .A1(n4591), .A2(n8964), .ZN(n4590) );
  NAND2_X1 U5509 ( .A1(n8952), .A2(n9004), .ZN(n4589) );
  NAND2_X1 U5510 ( .A1(n4583), .A2(n4579), .ZN(n9007) );
  NAND2_X1 U5511 ( .A1(n4580), .A2(n4502), .ZN(n4579) );
  NAND2_X1 U5512 ( .A1(n9005), .A2(n9004), .ZN(n4583) );
  NAND2_X1 U5513 ( .A1(n4470), .A2(n4575), .ZN(n4574) );
  INV_X1 U5514 ( .A(n9015), .ZN(n4575) );
  OAI21_X1 U5515 ( .B1(n9015), .B2(n9010), .A(n4517), .ZN(n4578) );
  INV_X1 U5516 ( .A(n7265), .ZN(n4832) );
  NOR2_X1 U5517 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5717) );
  AOI21_X1 U5518 ( .B1(n9027), .B2(n9004), .A(n9028), .ZN(n4586) );
  NAND2_X1 U5519 ( .A1(n9026), .A2(n9030), .ZN(n4585) );
  NAND2_X1 U5520 ( .A1(n9216), .A2(n4754), .ZN(n4753) );
  INV_X1 U5521 ( .A(n4755), .ZN(n4754) );
  NOR2_X1 U5522 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5389) );
  AOI21_X1 U5523 ( .B1(n4845), .B2(n4842), .A(n4841), .ZN(n4840) );
  INV_X1 U5524 ( .A(n5330), .ZN(n4841) );
  INV_X1 U5525 ( .A(n4847), .ZN(n4842) );
  INV_X1 U5526 ( .A(n4845), .ZN(n4843) );
  INV_X1 U5527 ( .A(SI_16_), .ZN(n5141) );
  INV_X1 U5528 ( .A(n5308), .ZN(n4862) );
  INV_X1 U5529 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5123) );
  INV_X1 U5530 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5113) );
  AOI21_X1 U5531 ( .B1(n4798), .B2(n4801), .A(n4516), .ZN(n4796) );
  INV_X1 U5532 ( .A(n6196), .ZN(n6118) );
  AOI21_X1 U5533 ( .B1(n5001), .B2(n5004), .A(n4999), .ZN(n4998) );
  INV_X1 U5534 ( .A(n8105), .ZN(n4999) );
  NAND2_X1 U5535 ( .A1(n4597), .A2(n4595), .ZN(n4594) );
  NOR2_X1 U5536 ( .A1(n8111), .A2(n4596), .ZN(n4595) );
  NAND2_X1 U5537 ( .A1(n8107), .A2(n8106), .ZN(n4596) );
  NAND2_X1 U5538 ( .A1(n8191), .A2(n4700), .ZN(n8214) );
  NAND2_X1 U5539 ( .A1(n8199), .A2(n4701), .ZN(n4700) );
  INV_X1 U5540 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n4701) );
  NAND2_X1 U5541 ( .A1(n8539), .A2(n8344), .ZN(n4687) );
  OR2_X1 U5542 ( .A1(n6190), .A2(n6251), .ZN(n6238) );
  NOR2_X1 U5543 ( .A1(n8593), .A2(n8596), .ZN(n4693) );
  INV_X1 U5544 ( .A(n8051), .ZN(n4995) );
  NOR2_X1 U5545 ( .A1(n8140), .A2(n4996), .ZN(n4992) );
  INV_X1 U5546 ( .A(n8055), .ZN(n4996) );
  NAND2_X1 U5547 ( .A1(n4684), .A2(n8617), .ZN(n4683) );
  INV_X1 U5548 ( .A(n8035), .ZN(n4647) );
  INV_X1 U5549 ( .A(n8031), .ZN(n5016) );
  NOR2_X1 U5550 ( .A1(n8623), .A2(n7829), .ZN(n4684) );
  NAND2_X1 U5551 ( .A1(n9805), .A2(n9872), .ZN(n5031) );
  NAND2_X1 U5552 ( .A1(n8172), .A2(n9860), .ZN(n7999) );
  AND3_X1 U5553 ( .A1(n5832), .A2(n4671), .A3(n4673), .ZN(n4672) );
  INV_X1 U5554 ( .A(n5752), .ZN(n4673) );
  INV_X1 U5555 ( .A(n5716), .ZN(n5034) );
  INV_X1 U5556 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5742) );
  INV_X1 U5557 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5715) );
  AND2_X1 U5558 ( .A1(n10237), .A2(n10247), .ZN(n4825) );
  NAND2_X1 U5559 ( .A1(n4945), .A2(n4942), .ZN(n4941) );
  NAND2_X1 U5560 ( .A1(n7612), .A2(n7493), .ZN(n4942) );
  NAND2_X1 U5561 ( .A1(n4936), .A2(n4935), .ZN(n7664) );
  AOI21_X1 U5562 ( .B1(n4937), .B2(n4939), .A(n4514), .ZN(n4935) );
  AOI21_X1 U5563 ( .B1(n4980), .B2(n4983), .A(n4978), .ZN(n4977) );
  INV_X1 U5564 ( .A(n4980), .ZN(n4979) );
  NOR2_X1 U5565 ( .A1(n7634), .A2(n7635), .ZN(n4978) );
  INV_X1 U5566 ( .A(n6652), .ZN(n4973) );
  INV_X1 U5567 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5494) );
  AND2_X1 U5568 ( .A1(n4614), .A2(n4613), .ZN(n9108) );
  NAND2_X1 U5569 ( .A1(n9638), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4613) );
  OR2_X1 U5570 ( .A1(n9367), .A2(n7766), .ZN(n8917) );
  NAND2_X1 U5571 ( .A1(n9225), .A2(n4756), .ZN(n4755) );
  NAND2_X1 U5572 ( .A1(n5548), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5565) );
  OR2_X1 U5573 ( .A1(n5509), .A2(n5508), .ZN(n5517) );
  INV_X1 U5574 ( .A(n8836), .ZN(n4730) );
  INV_X1 U5575 ( .A(n8846), .ZN(n4726) );
  OR2_X1 U5576 ( .A1(n5495), .A2(n5494), .ZN(n5502) );
  NAND2_X1 U5577 ( .A1(n5501), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5509) );
  INV_X1 U5578 ( .A(n5502), .ZN(n5501) );
  NOR2_X1 U5579 ( .A1(n5660), .A2(n4892), .ZN(n4891) );
  NOR2_X1 U5580 ( .A1(n4893), .A2(n5660), .ZN(n4890) );
  OAI21_X1 U5581 ( .B1(n6842), .B2(n4925), .A(n4923), .ZN(n7194) );
  INV_X1 U5582 ( .A(n4926), .ZN(n4925) );
  AOI21_X1 U5583 ( .B1(n4926), .B2(n4924), .A(n4492), .ZN(n4923) );
  AND2_X1 U5584 ( .A1(n6919), .A2(n4760), .ZN(n4759) );
  INV_X1 U5585 ( .A(n8937), .ZN(n4573) );
  NAND2_X1 U5586 ( .A1(n6741), .A2(n6587), .ZN(n9048) );
  INV_X1 U5587 ( .A(n4872), .ZN(n4871) );
  AOI21_X1 U5588 ( .B1(n4872), .B2(n4874), .A(n4870), .ZN(n4869) );
  AND2_X1 U5589 ( .A1(n5206), .A2(n5205), .ZN(n5218) );
  AND2_X1 U5590 ( .A1(n5199), .A2(n5198), .ZN(n5382) );
  INV_X1 U5591 ( .A(n5186), .ZN(n4876) );
  AOI21_X1 U5592 ( .B1(n5187), .B2(n4875), .A(n4873), .ZN(n4872) );
  INV_X1 U5593 ( .A(n5193), .ZN(n4873) );
  OR2_X1 U5594 ( .A1(n5364), .A2(n5363), .ZN(n5175) );
  OAI21_X1 U5595 ( .B1(n5338), .B2(n5150), .A(n5149), .ZN(n5346) );
  NOR2_X1 U5596 ( .A1(n5323), .A2(n4848), .ZN(n4847) );
  INV_X1 U5597 ( .A(n5132), .ZN(n4848) );
  AOI21_X1 U5598 ( .B1(n5133), .B2(n4847), .A(n4846), .ZN(n4845) );
  INV_X1 U5599 ( .A(n5138), .ZN(n4846) );
  AND2_X1 U5600 ( .A1(n5316), .A2(n5315), .ZN(n5333) );
  INV_X1 U5601 ( .A(n5116), .ZN(n4865) );
  INV_X1 U5602 ( .A(n4864), .ZN(n4863) );
  OAI21_X1 U5603 ( .B1(n4866), .B2(n4483), .A(n5122), .ZN(n4864) );
  INV_X1 U5604 ( .A(SI_10_), .ZN(n5107) );
  AOI21_X1 U5605 ( .B1(n4631), .B2(n4634), .A(n4630), .ZN(n4629) );
  OAI21_X1 U5606 ( .B1(n5255), .B2(n4854), .A(n5265), .ZN(n4853) );
  INV_X1 U5607 ( .A(n5089), .ZN(n4854) );
  INV_X1 U5608 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5047) );
  NAND2_X1 U5609 ( .A1(n5772), .A2(n5229), .ZN(n5072) );
  AND2_X1 U5610 ( .A1(n5235), .A2(n5046), .ZN(n5237) );
  XNOR2_X1 U5611 ( .A(n5072), .B(SI_1_), .ZN(n5225) );
  INV_X1 U5612 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5068) );
  AOI21_X1 U5613 ( .B1(n4823), .B2(n4821), .A(n4560), .ZN(n4820) );
  INV_X1 U5614 ( .A(n7826), .ZN(n4821) );
  INV_X1 U5615 ( .A(n5758), .ZN(n5760) );
  OR2_X1 U5616 ( .A1(n6097), .A2(n7820), .ZN(n6099) );
  NAND2_X1 U5617 ( .A1(n7903), .A2(n5949), .ZN(n7827) );
  OR2_X1 U5618 ( .A1(n6099), .A2(n10204), .ZN(n6129) );
  NAND2_X1 U5619 ( .A1(n6073), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6097) );
  INV_X1 U5620 ( .A(n6075), .ZN(n6073) );
  NAND2_X1 U5621 ( .A1(n7827), .A2(n7826), .ZN(n7825) );
  OR2_X1 U5622 ( .A1(n5968), .A2(n5967), .ZN(n5987) );
  OR2_X1 U5623 ( .A1(n5954), .A2(n10132), .ZN(n5968) );
  NOR2_X1 U5624 ( .A1(n6858), .A2(n4827), .ZN(n4826) );
  INV_X1 U5625 ( .A(n5821), .ZN(n4827) );
  AND2_X1 U5626 ( .A1(n6183), .A2(n6182), .ZN(n8309) );
  OR2_X1 U5627 ( .A1(n8346), .A2(n6178), .ZN(n6183) );
  AND4_X1 U5628 ( .A1(n6103), .A2(n6102), .A3(n6101), .A4(n6100), .ZN(n8294)
         );
  AND4_X1 U5629 ( .A1(n6065), .A2(n6064), .A3(n6063), .A4(n6062), .ZN(n8287)
         );
  AND4_X1 U5630 ( .A1(n6018), .A2(n6017), .A3(n6016), .A4(n6015), .ZN(n8166)
         );
  AND4_X1 U5631 ( .A1(n5992), .A2(n5991), .A3(n5990), .A4(n5989), .ZN(n7936)
         );
  NAND2_X1 U5632 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n4703) );
  AOI21_X1 U5633 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7062), .A(n7056), .ZN(
        n6997) );
  NAND2_X1 U5634 ( .A1(n7028), .A2(n4702), .ZN(n7030) );
  OR2_X1 U5635 ( .A1(n7029), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4702) );
  NAND2_X1 U5636 ( .A1(n7030), .A2(n7031), .ZN(n8191) );
  NAND2_X1 U5637 ( .A1(n8253), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4697) );
  NAND2_X1 U5638 ( .A1(n7755), .A2(n7754), .ZN(n8280) );
  AND2_X1 U5639 ( .A1(n8331), .A2(n4780), .ZN(n4779) );
  NAND2_X1 U5640 ( .A1(n8352), .A2(n8310), .ZN(n4780) );
  INV_X1 U5641 ( .A(n8310), .ZN(n4781) );
  OR2_X1 U5642 ( .A1(n8365), .A2(n8550), .ZN(n8342) );
  AND3_X1 U5643 ( .A1(n6165), .A2(n6164), .A3(n6163), .ZN(n8378) );
  AOI21_X1 U5644 ( .B1(n4489), .B2(n8471), .A(n5020), .ZN(n5019) );
  INV_X1 U5645 ( .A(n8079), .ZN(n5020) );
  NAND2_X1 U5646 ( .A1(n5021), .A2(n4469), .ZN(n8446) );
  NAND2_X1 U5647 ( .A1(n8493), .A2(n4693), .ZN(n8476) );
  AND2_X1 U5648 ( .A1(n8493), .A2(n4691), .ZN(n8455) );
  OR2_X1 U5649 ( .A1(n8472), .A2(n8471), .ZN(n8459) );
  INV_X1 U5650 ( .A(n6032), .ZN(n6031) );
  NAND2_X1 U5651 ( .A1(n8515), .A2(n8140), .ZN(n4775) );
  AND2_X1 U5652 ( .A1(n5007), .A2(n5008), .ZN(n7578) );
  AOI21_X1 U5653 ( .B1(n5009), .B2(n5015), .A(n5018), .ZN(n5008) );
  NAND2_X1 U5654 ( .A1(n4648), .A2(n5009), .ZN(n5007) );
  AND2_X1 U5655 ( .A1(n8623), .A2(n8040), .ZN(n5018) );
  NAND2_X1 U5656 ( .A1(n7578), .A2(n8137), .ZN(n7606) );
  NAND2_X1 U5657 ( .A1(n4788), .A2(n4786), .ZN(n7576) );
  NAND2_X1 U5658 ( .A1(n4787), .A2(n4486), .ZN(n4786) );
  NAND2_X1 U5659 ( .A1(n4490), .A2(n8135), .ZN(n4787) );
  NOR2_X1 U5660 ( .A1(n7519), .A2(n4682), .ZN(n7581) );
  INV_X1 U5661 ( .A(n4684), .ZN(n4682) );
  AND4_X1 U5662 ( .A1(n5919), .A2(n5918), .A3(n5917), .A4(n5916), .ZN(n7910)
         );
  AND2_X1 U5663 ( .A1(n8026), .A2(n8025), .ZN(n7396) );
  CLKBUF_X1 U5664 ( .A(n5899), .Z(n6998) );
  NAND2_X1 U5665 ( .A1(n5027), .A2(n8015), .ZN(n5026) );
  INV_X1 U5666 ( .A(n5029), .ZN(n5027) );
  NOR2_X1 U5667 ( .A1(n9793), .A2(n4785), .ZN(n4784) );
  INV_X1 U5668 ( .A(n9798), .ZN(n4680) );
  NAND2_X1 U5669 ( .A1(n7372), .A2(n5031), .ZN(n9803) );
  NAND2_X1 U5670 ( .A1(n7338), .A2(n8129), .ZN(n7372) );
  INV_X1 U5671 ( .A(n7285), .ZN(n8122) );
  AND2_X1 U5672 ( .A1(n7255), .A2(n9860), .ZN(n7281) );
  NOR2_X1 U5673 ( .A1(n6719), .A2(n7322), .ZN(n7255) );
  NAND2_X1 U5674 ( .A1(n4689), .A2(n9826), .ZN(n6719) );
  INV_X1 U5675 ( .A(n6801), .ZN(n4689) );
  NAND2_X1 U5676 ( .A1(n6802), .A2(n6803), .ZN(n6801) );
  AND2_X1 U5677 ( .A1(n8127), .A2(n8124), .ZN(n6804) );
  NAND2_X1 U5678 ( .A1(n6770), .A2(n7993), .ZN(n8127) );
  AND2_X1 U5679 ( .A1(n9843), .A2(n9846), .ZN(n6227) );
  NAND2_X1 U5680 ( .A1(n6160), .A2(n6159), .ZN(n8557) );
  NAND2_X1 U5681 ( .A1(n6117), .A2(n6116), .ZN(n8565) );
  INV_X1 U5682 ( .A(n7384), .ZN(n7385) );
  OR2_X1 U5683 ( .A1(n6643), .A2(n8152), .ZN(n9907) );
  NAND2_X1 U5684 ( .A1(n7289), .A2(n7288), .ZN(n7290) );
  INV_X1 U5685 ( .A(n9905), .ZN(n8624) );
  NAND2_X1 U5686 ( .A1(n7402), .A2(n9878), .ZN(n9912) );
  INV_X1 U5687 ( .A(n6704), .ZN(n7251) );
  AND2_X1 U5688 ( .A1(n6624), .A2(n6623), .ZN(n6705) );
  XNOR2_X1 U5689 ( .A(n5754), .B(n5753), .ZN(n7003) );
  INV_X1 U5690 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U5691 ( .A1(n4678), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5754) );
  NAND2_X1 U5692 ( .A1(n4674), .A2(n4672), .ZN(n4678) );
  INV_X1 U5693 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n10077) );
  INV_X1 U5694 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5733) );
  INV_X1 U5695 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5732) );
  AND2_X1 U5696 ( .A1(n5922), .A2(n5932), .ZN(n7146) );
  AND2_X1 U5697 ( .A1(n5904), .A2(n5903), .ZN(n6993) );
  AND2_X1 U5698 ( .A1(n5832), .A2(n5714), .ZN(n5861) );
  OR2_X1 U5699 ( .A1(n5540), .A2(n8699), .ZN(n5550) );
  NAND2_X1 U5700 ( .A1(n8718), .A2(n4984), .ZN(n4982) );
  NOR2_X1 U5701 ( .A1(n8718), .A2(n4984), .ZN(n4983) );
  INV_X1 U5702 ( .A(n4964), .ZN(n8684) );
  NAND2_X1 U5703 ( .A1(n8742), .A2(n8743), .ZN(n8741) );
  OR2_X1 U5704 ( .A1(n9036), .A2(n6535), .ZN(n6522) );
  INV_X1 U5705 ( .A(n7693), .ZN(n7677) );
  NAND2_X1 U5706 ( .A1(n8911), .A2(n5062), .ZN(n9035) );
  OR3_X1 U5707 ( .A1(n8910), .A2(n9066), .A3(n8909), .ZN(n8911) );
  OR2_X1 U5708 ( .A1(n5419), .A2(n5408), .ZN(n5410) );
  NAND2_X1 U5709 ( .A1(n5404), .A2(n5405), .ZN(n4570) );
  OR2_X1 U5710 ( .A1(n6578), .A2(n6577), .ZN(n4618) );
  NOR2_X1 U5711 ( .A1(n6819), .A2(n6818), .ZN(n6817) );
  AND2_X1 U5712 ( .A1(n9104), .A2(n9105), .ZN(n9619) );
  XNOR2_X1 U5713 ( .A(n9108), .B(n9653), .ZN(n9648) );
  NOR2_X1 U5714 ( .A1(n9704), .A2(n9703), .ZN(n9702) );
  XNOR2_X1 U5715 ( .A(n4619), .B(n5544), .ZN(n9134) );
  OR2_X1 U5716 ( .A1(n9702), .A2(n4620), .ZN(n4619) );
  AND2_X1 U5717 ( .A1(n9708), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4620) );
  XNOR2_X1 U5718 ( .A(n5631), .B(n5667), .ZN(n4735) );
  AND2_X1 U5719 ( .A1(n5622), .A2(n5614), .ZN(n9161) );
  OR2_X1 U5720 ( .A1(n9382), .A2(n9208), .ZN(n9181) );
  OR2_X1 U5721 ( .A1(n8906), .A2(n8905), .ZN(n9184) );
  OAI21_X1 U5722 ( .B1(n4745), .B2(n4567), .A(n8925), .ZN(n4743) );
  NAND2_X1 U5723 ( .A1(n4902), .A2(n4910), .ZN(n4898) );
  OR2_X1 U5724 ( .A1(n4903), .A2(n4900), .ZN(n4899) );
  INV_X1 U5725 ( .A(n4910), .ZN(n4900) );
  NOR2_X1 U5726 ( .A1(n9253), .A2(n4755), .ZN(n9221) );
  NOR2_X1 U5727 ( .A1(n9253), .A2(n9395), .ZN(n9237) );
  OR2_X1 U5728 ( .A1(n8931), .A2(n5539), .ZN(n4724) );
  NAND2_X1 U5729 ( .A1(n5524), .A2(n4720), .ZN(n4719) );
  NAND2_X1 U5730 ( .A1(n4719), .A2(n4487), .ZN(n9285) );
  NAND2_X1 U5731 ( .A1(n5525), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5540) );
  INV_X1 U5732 ( .A(n5534), .ZN(n5525) );
  NAND2_X1 U5733 ( .A1(n5524), .A2(n8982), .ZN(n9316) );
  NAND2_X1 U5734 ( .A1(n7549), .A2(n4472), .ZN(n9308) );
  AND2_X1 U5735 ( .A1(n9299), .A2(n9298), .ZN(n9315) );
  OR2_X1 U5736 ( .A1(n9430), .A2(n9086), .ZN(n4883) );
  NAND2_X1 U5737 ( .A1(n9346), .A2(n4501), .ZN(n4884) );
  NAND2_X1 U5738 ( .A1(n7549), .A2(n5329), .ZN(n9352) );
  INV_X1 U5739 ( .A(n9089), .ZN(n7528) );
  INV_X1 U5740 ( .A(n9087), .ZN(n9344) );
  NAND2_X1 U5741 ( .A1(n5476), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5486) );
  INV_X1 U5742 ( .A(n5478), .ZN(n5476) );
  INV_X1 U5743 ( .A(n9090), .ZN(n9500) );
  NAND2_X1 U5744 ( .A1(n4713), .A2(n4509), .ZN(n9495) );
  NAND2_X1 U5745 ( .A1(n8934), .A2(n8887), .ZN(n4714) );
  OR2_X1 U5746 ( .A1(n9510), .A2(n7356), .ZN(n9498) );
  INV_X1 U5747 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5469) );
  OR2_X1 U5748 ( .A1(n5470), .A2(n5469), .ZN(n5478) );
  OR2_X1 U5749 ( .A1(n5462), .A2(n5461), .ZN(n5470) );
  NAND2_X1 U5750 ( .A1(n7211), .A2(n8934), .ZN(n7196) );
  INV_X1 U5751 ( .A(n9091), .ZN(n7356) );
  AND3_X1 U5752 ( .A1(n6914), .A2(n4759), .A3(n4758), .ZN(n7221) );
  AND2_X1 U5753 ( .A1(n7215), .A2(n5654), .ZN(n4926) );
  NAND2_X1 U5754 ( .A1(n6914), .A2(n4759), .ZN(n7219) );
  NAND2_X1 U5755 ( .A1(n6842), .A2(n8887), .ZN(n6841) );
  OR2_X1 U5756 ( .A1(n6848), .A2(n8887), .ZN(n7211) );
  NAND2_X1 U5757 ( .A1(n6914), .A2(n6919), .ZN(n6915) );
  NAND2_X1 U5758 ( .A1(n4573), .A2(n5650), .ZN(n6909) );
  AND2_X1 U5759 ( .A1(n6762), .A2(n5651), .ZN(n6906) );
  NAND2_X1 U5760 ( .A1(n9048), .A2(n8853), .ZN(n6526) );
  NAND2_X1 U5761 ( .A1(n6605), .A2(n5407), .ZN(n9046) );
  XNOR2_X1 U5762 ( .A(n5644), .B(n9042), .ZN(n8884) );
  INV_X1 U5763 ( .A(n9099), .ZN(n6608) );
  INV_X1 U5764 ( .A(n9501), .ZN(n9319) );
  NAND2_X1 U5765 ( .A1(n5358), .A2(n5357), .ZN(n9405) );
  NAND2_X1 U5766 ( .A1(n5354), .A2(n5353), .ZN(n9410) );
  INV_X1 U5767 ( .A(n9760), .ZN(n9750) );
  INV_X1 U5768 ( .A(n9762), .ZN(n9751) );
  OR2_X1 U5769 ( .A1(n6536), .A2(n6535), .ZN(n9760) );
  XNOR2_X1 U5770 ( .A(n5693), .B(n5692), .ZN(n7473) );
  OAI21_X1 U5771 ( .B1(n7733), .B2(n10152), .A(n7726), .ZN(n7730) );
  AND2_X1 U5772 ( .A1(n4929), .A2(n4928), .ZN(n4927) );
  INV_X1 U5773 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4928) );
  XNOR2_X1 U5774 ( .A(n7733), .B(SI_30_), .ZN(n8651) );
  XNOR2_X1 U5775 ( .A(n7736), .B(n7738), .ZN(n8653) );
  NAND2_X1 U5776 ( .A1(n5221), .A2(n5206), .ZN(n7712) );
  OAI21_X1 U5777 ( .B1(n5375), .B2(n5187), .A(n5186), .ZN(n5379) );
  XNOR2_X1 U5778 ( .A(n5681), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5696) );
  INV_X1 U5779 ( .A(n5679), .ZN(n5680) );
  XNOR2_X1 U5780 ( .A(n5375), .B(n5374), .ZN(n7556) );
  INV_X1 U5781 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5067) );
  NAND2_X1 U5782 ( .A1(n4844), .A2(n5132), .ZN(n5324) );
  OR2_X1 U5783 ( .A1(n5314), .A2(n5133), .ZN(n4844) );
  INV_X1 U5784 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5317) );
  OR3_X1 U5785 ( .A1(n5300), .A2(P1_IR_REG_10__SCAN_IN), .A3(
        P1_IR_REG_11__SCAN_IN), .ZN(n5302) );
  NOR2_X1 U5786 ( .A1(n5302), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5316) );
  NAND2_X1 U5787 ( .A1(n4628), .A2(n4631), .ZN(n5280) );
  OR2_X1 U5788 ( .A1(n5268), .A2(n4634), .ZN(n4628) );
  INV_X1 U5789 ( .A(n7409), .ZN(n9891) );
  NAND2_X1 U5790 ( .A1(n5912), .A2(n7344), .ZN(n6261) );
  AND4_X1 U5791 ( .A1(n6080), .A2(n6079), .A3(n6078), .A4(n6077), .ZN(n8475)
         );
  NAND2_X1 U5792 ( .A1(n4794), .A2(n5774), .ZN(n6825) );
  INV_X1 U5793 ( .A(n4795), .ZN(n4794) );
  AND2_X1 U5794 ( .A1(n5774), .A2(n5762), .ZN(n6827) );
  NAND2_X1 U5795 ( .A1(n7837), .A2(n7836), .ZN(n7835) );
  NAND2_X1 U5796 ( .A1(n6010), .A2(n6009), .ZN(n8606) );
  NAND2_X1 U5797 ( .A1(n5905), .A2(n4991), .ZN(n4990) );
  NAND2_X1 U5798 ( .A1(n6865), .A2(n5821), .ZN(n6859) );
  NAND2_X1 U5799 ( .A1(n6030), .A2(n6029), .ZN(n8603) );
  INV_X1 U5800 ( .A(n4805), .ZN(n4804) );
  OAI21_X1 U5801 ( .B1(n4808), .B2(n4807), .A(n4523), .ZN(n4805) );
  NAND2_X1 U5802 ( .A1(n6072), .A2(n6071), .ZN(n8586) );
  AND2_X1 U5803 ( .A1(n4802), .A2(n7810), .ZN(n7874) );
  NAND2_X1 U5804 ( .A1(n7825), .A2(n5963), .ZN(n7882) );
  INV_X1 U5805 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10204) );
  NAND2_X1 U5806 ( .A1(n6087), .A2(n6086), .ZN(n8576) );
  NAND2_X1 U5807 ( .A1(n6259), .A2(n5931), .ZN(n7905) );
  AND2_X1 U5808 ( .A1(n4815), .A2(n7926), .ZN(n4813) );
  AND2_X1 U5809 ( .A1(n4814), .A2(n4815), .ZN(n7927) );
  INV_X1 U5810 ( .A(n7909), .ZN(n7940) );
  INV_X1 U5811 ( .A(n7933), .ZN(n7941) );
  INV_X1 U5812 ( .A(n8162), .ZN(n4625) );
  AND4_X1 U5813 ( .A1(n6049), .A2(n6048), .A3(n6047), .A4(n6046), .ZN(n8492)
         );
  INV_X1 U5814 ( .A(n7276), .ZN(n8171) );
  NAND2_X1 U5815 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4704) );
  AOI21_X1 U5816 ( .B1(n6981), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7104), .ZN(
        n7118) );
  AOI21_X1 U5817 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(n6982), .A(n7116), .ZN(
        n7131) );
  AND2_X1 U5818 ( .A1(n6991), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4694) );
  NAND2_X1 U5819 ( .A1(n8178), .A2(n4705), .ZN(n7058) );
  NAND2_X1 U5820 ( .A1(n4707), .A2(n4706), .ZN(n4705) );
  INV_X1 U5821 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n4706) );
  INV_X1 U5822 ( .A(n8183), .ZN(n4707) );
  NOR2_X1 U5823 ( .A1(n8226), .A2(n4699), .ZN(n8229) );
  AND2_X1 U5824 ( .A1(n8232), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4699) );
  INV_X1 U5825 ( .A(n4698), .ZN(n8252) );
  INV_X1 U5826 ( .A(n4856), .ZN(n8532) );
  INV_X1 U5827 ( .A(n7953), .ZN(n8539) );
  NAND2_X1 U5828 ( .A1(n5000), .A2(n5005), .ZN(n8314) );
  AOI21_X1 U5829 ( .B1(n8338), .B2(n9857), .A(n8337), .ZN(n8548) );
  NAND2_X1 U5830 ( .A1(n8336), .A2(n8335), .ZN(n8337) );
  NAND2_X1 U5831 ( .A1(n5024), .A2(n7972), .ZN(n8361) );
  INV_X1 U5832 ( .A(n8565), .ZN(n8397) );
  NAND2_X1 U5833 ( .A1(n8420), .A2(n8301), .ZN(n8393) );
  CLKBUF_X1 U5834 ( .A(n8390), .Z(n8391) );
  NAND2_X1 U5835 ( .A1(n4640), .A2(n4644), .ZN(n8411) );
  NAND2_X1 U5836 ( .A1(n5021), .A2(n4645), .ZN(n4640) );
  INV_X1 U5837 ( .A(n8576), .ZN(n8432) );
  AND2_X1 U5838 ( .A1(n6096), .A2(n6095), .ZN(n8444) );
  AND2_X1 U5839 ( .A1(n6056), .A2(n6055), .ZN(n8482) );
  OAI21_X1 U5840 ( .B1(n8515), .B2(n4773), .A(n4771), .ZN(n8485) );
  NAND2_X1 U5841 ( .A1(n8519), .A2(n8051), .ZN(n8502) );
  NAND2_X1 U5842 ( .A1(n5011), .A2(n5012), .ZN(n7562) );
  AND2_X1 U5843 ( .A1(n4789), .A2(n4490), .ZN(n7575) );
  NAND2_X1 U5844 ( .A1(n5017), .A2(n8031), .ZN(n7561) );
  OR2_X1 U5845 ( .A1(n7515), .A2(n7514), .ZN(n5017) );
  AND2_X1 U5846 ( .A1(n7291), .A2(n7288), .ZN(n4782) );
  NAND2_X1 U5847 ( .A1(n5809), .A2(n9482), .ZN(n4987) );
  INV_X1 U5848 ( .A(n6316), .ZN(n4989) );
  OR2_X1 U5849 ( .A1(n9844), .A2(n6247), .ZN(n8345) );
  INV_X1 U5850 ( .A(n8529), .ZN(n8512) );
  INV_X1 U5851 ( .A(n9835), .ZN(n7410) );
  AND2_X2 U5852 ( .A1(n6705), .A2(n6704), .ZN(n9927) );
  AND2_X2 U5853 ( .A1(n6705), .A2(n7251), .ZN(n9915) );
  AND2_X1 U5854 ( .A1(n6352), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9850) );
  INV_X1 U5855 ( .A(n9845), .ZN(n9848) );
  NAND2_X1 U5856 ( .A1(n4793), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4792) );
  NAND2_X1 U5857 ( .A1(n6203), .A2(n6202), .ZN(n7595) );
  INV_X1 U5858 ( .A(n6205), .ZN(n6207) );
  INV_X1 U5859 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n10120) );
  NAND2_X1 U5860 ( .A1(n6211), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6213) );
  INV_X1 U5861 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n10128) );
  INV_X1 U5862 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7090) );
  INV_X1 U5863 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7086) );
  INV_X1 U5864 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5737) );
  INV_X1 U5865 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7600) );
  INV_X1 U5866 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6710) );
  INV_X1 U5867 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10095) );
  INV_X1 U5868 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6351) );
  INV_X1 U5869 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6347) );
  INV_X1 U5870 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10246) );
  INV_X1 U5871 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6337) );
  INV_X1 U5872 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6330) );
  INV_X1 U5873 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6324) );
  NAND2_X1 U5874 ( .A1(n5223), .A2(n5222), .ZN(n9370) );
  NAND2_X1 U5875 ( .A1(n5322), .A2(n5321), .ZN(n8835) );
  NAND2_X1 U5876 ( .A1(n4950), .A2(n7044), .ZN(n7232) );
  NAND2_X1 U5877 ( .A1(n7040), .A2(n7039), .ZN(n4950) );
  NAND2_X1 U5878 ( .A1(n8741), .A2(n7655), .ZN(n8705) );
  NAND2_X1 U5879 ( .A1(n5307), .A2(n5306), .ZN(n7485) );
  NAND2_X1 U5880 ( .A1(n4964), .A2(n4963), .ZN(n4960) );
  NAND2_X1 U5881 ( .A1(n4975), .A2(n4982), .ZN(n8728) );
  NAND2_X1 U5882 ( .A1(n8720), .A2(n4976), .ZN(n4975) );
  INV_X1 U5883 ( .A(n4983), .ZN(n4976) );
  NAND2_X1 U5884 ( .A1(n6450), .A2(n6449), .ZN(n6653) );
  INV_X1 U5885 ( .A(n9273), .ZN(n8758) );
  NAND2_X1 U5886 ( .A1(n4946), .A2(n4947), .ZN(n7455) );
  INV_X1 U5887 ( .A(n8778), .ZN(n8801) );
  AND2_X1 U5888 ( .A1(n6420), .A2(n5635), .ZN(n8789) );
  INV_X1 U5889 ( .A(n8782), .ZN(n8765) );
  NAND2_X1 U5890 ( .A1(n4951), .A2(n4954), .ZN(n8788) );
  OAI21_X1 U5891 ( .B1(n8711), .B2(n4966), .A(n4528), .ZN(n4955) );
  NAND2_X1 U5892 ( .A1(n5385), .A2(n5384), .ZN(n9375) );
  NAND3_X1 U5893 ( .A1(n4931), .A2(n4930), .A3(n4932), .ZN(n9078) );
  OAI22_X1 U5894 ( .A1(n9451), .A2(n4933), .B1(P1_IR_REG_22__SCAN_IN), .B2(
        P1_IR_REG_31__SCAN_IN), .ZN(n4932) );
  OR2_X1 U5895 ( .A1(n7702), .A2(n5636), .ZN(n5630) );
  NAND2_X1 U5896 ( .A1(n5610), .A2(n5609), .ZN(n9164) );
  OR2_X1 U5897 ( .A1(n9212), .A2(n5636), .ZN(n5591) );
  NAND2_X1 U5898 ( .A1(n6496), .A2(n4548), .ZN(n6495) );
  XNOR2_X1 U5899 ( .A(n4612), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6493) );
  NAND2_X1 U5900 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4612) );
  NAND2_X1 U5901 ( .A1(n4618), .A2(n4617), .ZN(n6468) );
  AOI21_X1 U5902 ( .B1(n4617), .B2(n6577), .A(n4553), .ZN(n4616) );
  NAND2_X1 U5903 ( .A1(n9131), .A2(n5635), .ZN(n9691) );
  INV_X1 U5904 ( .A(n4614), .ZN(n9635) );
  INV_X1 U5905 ( .A(n4610), .ZN(n9662) );
  INV_X1 U5906 ( .A(n9111), .ZN(n4609) );
  NAND2_X1 U5907 ( .A1(n4913), .A2(n4917), .ZN(n5668) );
  AND2_X1 U5908 ( .A1(n5603), .A2(n5594), .ZN(n9197) );
  NAND2_X1 U5909 ( .A1(n9227), .A2(n8926), .ZN(n9205) );
  INV_X1 U5910 ( .A(n9390), .ZN(n9225) );
  NAND2_X1 U5911 ( .A1(n4901), .A2(n4904), .ZN(n9220) );
  NAND2_X1 U5912 ( .A1(n9247), .A2(n4905), .ZN(n4901) );
  AND2_X1 U5913 ( .A1(n4906), .A2(n4909), .ZN(n9236) );
  NAND2_X1 U5914 ( .A1(n9247), .A2(n9248), .ZN(n4906) );
  NAND2_X1 U5915 ( .A1(n5362), .A2(n5361), .ZN(n9402) );
  INV_X1 U5916 ( .A(n9405), .ZN(n9269) );
  AND2_X1 U5917 ( .A1(n4651), .A2(n4649), .ZN(n9263) );
  INV_X1 U5918 ( .A(n4652), .ZN(n4649) );
  NAND2_X1 U5919 ( .A1(n4653), .A2(n4657), .ZN(n9279) );
  NAND2_X1 U5920 ( .A1(n9307), .A2(n4654), .ZN(n4653) );
  INV_X1 U5921 ( .A(n4656), .ZN(n4654) );
  NAND2_X1 U5922 ( .A1(n4658), .A2(n4484), .ZN(n9291) );
  OR2_X1 U5923 ( .A1(n9307), .A2(n5661), .ZN(n4658) );
  NAND2_X1 U5924 ( .A1(n5336), .A2(n5335), .ZN(n9427) );
  NAND2_X1 U5925 ( .A1(n7526), .A2(n8836), .ZN(n7541) );
  NAND2_X1 U5926 ( .A1(n4888), .A2(n4893), .ZN(n7525) );
  NAND2_X1 U5927 ( .A1(n7354), .A2(n4889), .ZN(n4888) );
  INV_X1 U5928 ( .A(n4892), .ZN(n4889) );
  NAND2_X1 U5929 ( .A1(n5312), .A2(n5311), .ZN(n7537) );
  NAND2_X1 U5930 ( .A1(n4894), .A2(n5658), .ZN(n7475) );
  OR2_X1 U5931 ( .A1(n7354), .A2(n5659), .ZN(n4894) );
  AND2_X1 U5932 ( .A1(n6739), .A2(n5649), .ZN(n6763) );
  OR2_X1 U5933 ( .A1(n9519), .A2(n6537), .ZN(n7782) );
  OR2_X1 U5934 ( .A1(n9519), .A2(n6538), .ZN(n9357) );
  OR2_X1 U5935 ( .A1(n9756), .A2(n6377), .ZN(n9294) );
  NAND2_X1 U5936 ( .A1(n6758), .A2(n9294), .ZN(n9338) );
  NAND2_X1 U5937 ( .A1(n5228), .A2(n9466), .ZN(n5231) );
  INV_X1 U5938 ( .A(n9294), .ZN(n9508) );
  INV_X1 U5939 ( .A(n9357), .ZN(n9509) );
  INV_X1 U5940 ( .A(n7782), .ZN(n9361) );
  AND2_X1 U5941 ( .A1(n4667), .A2(n4556), .ZN(n4666) );
  OR2_X1 U5942 ( .A1(n9368), .A2(n9534), .ZN(n4665) );
  INV_X1 U5943 ( .A(n9366), .ZN(n4668) );
  NAND2_X1 U5944 ( .A1(n4733), .A2(n4508), .ZN(n9369) );
  INV_X1 U5945 ( .A(n9154), .ZN(n4733) );
  NOR2_X1 U5946 ( .A1(n9148), .A2(n4732), .ZN(n4731) );
  INV_X1 U5947 ( .A(n9718), .ZN(n9719) );
  XNOR2_X1 U5948 ( .A(n7712), .B(n7711), .ZN(n9462) );
  XNOR2_X1 U5949 ( .A(n5684), .B(P1_IR_REG_26__SCAN_IN), .ZN(n7591) );
  INV_X1 U5950 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7471) );
  INV_X1 U5951 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7761) );
  CLKBUF_X1 U5952 ( .A(n5669), .Z(n5062) );
  INV_X1 U5953 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10222) );
  INV_X1 U5954 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6924) );
  NAND2_X1 U5955 ( .A1(n5065), .A2(n5064), .ZN(n9135) );
  AND2_X1 U5956 ( .A1(n5342), .A2(n5347), .ZN(n9116) );
  INV_X1 U5957 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10102) );
  INV_X1 U5958 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10266) );
  INV_X1 U5959 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6344) );
  INV_X1 U5960 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6341) );
  INV_X1 U5961 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6332) );
  NAND2_X1 U5962 ( .A1(n4637), .A2(n5093), .ZN(n5273) );
  INV_X1 U5963 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10185) );
  OR2_X1 U5964 ( .A1(n5264), .A2(n5051), .ZN(n6465) );
  INV_X1 U5965 ( .A(n5263), .ZN(n5051) );
  NAND2_X1 U5966 ( .A1(n4851), .A2(n5089), .ZN(n4662) );
  NAND2_X1 U5967 ( .A1(n5256), .A2(n5255), .ZN(n4851) );
  INV_X1 U5968 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10226) );
  NOR2_X1 U5969 ( .A1(n7436), .A2(n10340), .ZN(n9957) );
  AOI21_X1 U5970 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9955), .ZN(n9954) );
  NOR2_X1 U5971 ( .A1(n9954), .A2(n9953), .ZN(n9952) );
  AOI21_X1 U5972 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9952), .ZN(n9951) );
  OAI21_X1 U5973 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9949), .ZN(n9947) );
  NAND2_X1 U5974 ( .A1(n7069), .A2(n5860), .ZN(n7078) );
  NAND2_X1 U5975 ( .A1(n4803), .A2(n4808), .ZN(n7269) );
  NAND2_X1 U5976 ( .A1(n4624), .A2(n4623), .ZN(P2_U3244) );
  OR2_X1 U5977 ( .A1(n8161), .A2(n8160), .ZN(n4623) );
  NAND2_X1 U5978 ( .A1(n4604), .A2(n4625), .ZN(n4624) );
  INV_X1 U5979 ( .A(n4696), .ZN(n7171) );
  INV_X1 U5980 ( .A(n4712), .ZN(n4711) );
  NAND2_X1 U5981 ( .A1(n4709), .A2(n8273), .ZN(n4708) );
  INV_X1 U5982 ( .A(n5905), .ZN(n5792) );
  AND2_X1 U5983 ( .A1(n5422), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n4468) );
  AND2_X1 U5984 ( .A1(n5019), .A2(n4646), .ZN(n4469) );
  INV_X1 U5985 ( .A(n9078), .ZN(n5672) );
  INV_X1 U5986 ( .A(n8471), .ZN(n7948) );
  OR2_X1 U5987 ( .A1(n8545), .A2(n8311), .ZN(n7968) );
  INV_X1 U5988 ( .A(n8998), .ZN(n4716) );
  NAND2_X1 U5989 ( .A1(n9016), .A2(n8924), .ZN(n4470) );
  INV_X1 U5990 ( .A(n8887), .ZN(n4924) );
  NAND2_X1 U5991 ( .A1(n7485), .A2(n9089), .ZN(n4471) );
  OR2_X1 U5992 ( .A1(n8576), .A2(n8296), .ZN(n8070) );
  AND2_X1 U5993 ( .A1(n4750), .A2(n9314), .ZN(n4472) );
  INV_X1 U5994 ( .A(n8140), .ZN(n4772) );
  NOR2_X1 U5995 ( .A1(n7231), .A2(n4949), .ZN(n4473) );
  INV_X1 U5996 ( .A(n4857), .ZN(n4855) );
  AND2_X1 U5997 ( .A1(n5748), .A2(n8273), .ZN(n4475) );
  INV_X1 U5998 ( .A(n5667), .ZN(n4915) );
  AOI21_X1 U5999 ( .B1(n4961), .B2(n7666), .A(n4955), .ZN(n4954) );
  INV_X1 U6000 ( .A(n4801), .ZN(n4800) );
  NAND2_X1 U6001 ( .A1(n7873), .A2(n7810), .ZN(n4801) );
  NAND2_X1 U6002 ( .A1(n5389), .A2(n5388), .ZN(n4477) );
  AND2_X1 U6003 ( .A1(n6358), .A2(n6382), .ZN(n6387) );
  OR2_X1 U6004 ( .A1(n4657), .A2(n4546), .ZN(n4478) );
  NAND2_X1 U6005 ( .A1(n8170), .A2(n9797), .ZN(n4479) );
  INV_X1 U6006 ( .A(n9284), .ZN(n4723) );
  OR2_X1 U6007 ( .A1(n7519), .A2(n4683), .ZN(n4480) );
  NAND2_X1 U6008 ( .A1(n6841), .A2(n4926), .ZN(n7214) );
  INV_X1 U6009 ( .A(n4463), .ZN(n7959) );
  INV_X1 U6010 ( .A(n5786), .ZN(n6241) );
  OR2_X1 U6011 ( .A1(n9370), .A2(n9186), .ZN(n4481) );
  AND3_X1 U6012 ( .A1(n5418), .A2(n5417), .A3(n5416), .ZN(n4482) );
  OR2_X1 U6013 ( .A1(n5299), .A2(n4865), .ZN(n4483) );
  OR2_X1 U6014 ( .A1(n9314), .A2(n9331), .ZN(n4484) );
  INV_X1 U6015 ( .A(n8711), .ZN(n4962) );
  INV_X1 U6016 ( .A(n8545), .ZN(n4688) );
  NAND2_X1 U6017 ( .A1(n6234), .A2(n6233), .ZN(n8545) );
  INV_X1 U6018 ( .A(n5234), .ZN(n5319) );
  OR2_X1 U6019 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6583), .ZN(n4485) );
  AND2_X1 U6020 ( .A1(n8059), .A2(n8060), .ZN(n8487) );
  INV_X1 U6021 ( .A(n8487), .ZN(n4770) );
  NAND2_X1 U6022 ( .A1(n8623), .A2(n8167), .ZN(n4486) );
  AND2_X1 U6023 ( .A1(n4723), .A2(n4724), .ZN(n4487) );
  NAND2_X1 U6024 ( .A1(n4856), .A2(n7954), .ZN(n4857) );
  OR2_X1 U6025 ( .A1(n8612), .A2(n7604), .ZN(n4488) );
  INV_X1 U6026 ( .A(n9852), .ZN(n4690) );
  AND2_X1 U6027 ( .A1(n8461), .A2(n8460), .ZN(n4489) );
  OR2_X1 U6028 ( .A1(n7829), .A2(n7558), .ZN(n4490) );
  AND3_X1 U6029 ( .A1(n5054), .A2(n5052), .A3(n5053), .ZN(n4491) );
  NAND2_X1 U6030 ( .A1(n5366), .A2(n5365), .ZN(n9395) );
  INV_X1 U6031 ( .A(n9395), .ZN(n4756) );
  AND2_X1 U6032 ( .A1(n9749), .A2(n9093), .ZN(n4492) );
  INV_X1 U6033 ( .A(n9219), .ZN(n4567) );
  NAND2_X1 U6034 ( .A1(n6173), .A2(n6172), .ZN(n8550) );
  AND2_X1 U6035 ( .A1(n4688), .A2(n8311), .ZN(n4493) );
  AND4_X1 U6036 ( .A1(n5720), .A2(n5719), .A3(n5718), .A4(n5717), .ZN(n4494)
         );
  NAND2_X1 U6037 ( .A1(n5328), .A2(n5327), .ZN(n9430) );
  AND2_X1 U6038 ( .A1(n5395), .A2(n5396), .ZN(n5415) );
  AND2_X1 U6039 ( .A1(n5257), .A2(n5048), .ZN(n5261) );
  OR3_X1 U6040 ( .A1(n8365), .A2(n8545), .A3(n4687), .ZN(n4495) );
  AND2_X1 U6041 ( .A1(n9395), .A2(n9229), .ZN(n4496) );
  NAND2_X1 U6042 ( .A1(n4764), .A2(n5832), .ZN(n5901) );
  OR2_X1 U6043 ( .A1(n9899), .A2(n7828), .ZN(n4497) );
  AND2_X1 U6044 ( .A1(n5422), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n4498) );
  AND2_X1 U6045 ( .A1(n5021), .A2(n5019), .ZN(n4499) );
  AND3_X1 U6046 ( .A1(n8921), .A2(n8920), .A3(n8919), .ZN(n4500) );
  NOR3_X1 U6047 ( .A1(n9253), .A2(n4753), .A3(n9382), .ZN(n4757) );
  NAND2_X1 U6048 ( .A1(n5966), .A2(n5965), .ZN(n8623) );
  NAND2_X1 U6049 ( .A1(n6045), .A2(n6044), .ZN(n8596) );
  INV_X1 U6050 ( .A(n8308), .ZN(n8352) );
  OR2_X1 U6051 ( .A1(n5329), .A2(n9330), .ZN(n4501) );
  NOR2_X1 U6052 ( .A1(n8994), .A2(n9004), .ZN(n4502) );
  AND2_X1 U6053 ( .A1(n6141), .A2(n6158), .ZN(n4503) );
  NAND2_X1 U6054 ( .A1(n5344), .A2(n5343), .ZN(n9420) );
  AND2_X1 U6055 ( .A1(n8015), .A2(n8129), .ZN(n4504) );
  AND2_X1 U6056 ( .A1(n9029), .A2(n4500), .ZN(n4505) );
  NAND2_X1 U6057 ( .A1(n5064), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5066) );
  INV_X1 U6058 ( .A(n5015), .ZN(n5014) );
  OR2_X1 U6059 ( .A1(n5016), .A2(n4647), .ZN(n5015) );
  INV_X1 U6060 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n10082) );
  INV_X1 U6061 ( .A(n4752), .ZN(n9210) );
  NOR2_X1 U6062 ( .A1(n9253), .A2(n4753), .ZN(n4752) );
  AND2_X1 U6063 ( .A1(n7763), .A2(n9171), .ZN(n4506) );
  OR2_X1 U6064 ( .A1(n5228), .A2(n6465), .ZN(n4507) );
  AND2_X1 U6065 ( .A1(n5677), .A2(n4731), .ZN(n4508) );
  AND2_X1 U6066 ( .A1(n4714), .A2(n8948), .ZN(n4509) );
  AND2_X1 U6067 ( .A1(n8003), .A2(n8103), .ZN(n4510) );
  INV_X1 U6068 ( .A(n4921), .ZN(n4920) );
  NAND2_X1 U6069 ( .A1(n4481), .A2(n8904), .ZN(n4921) );
  AND2_X1 U6070 ( .A1(n8944), .A2(n8933), .ZN(n4511) );
  NAND2_X1 U6071 ( .A1(n4957), .A2(n4962), .ZN(n4512) );
  AND2_X1 U6072 ( .A1(n9227), .A2(n4744), .ZN(n4513) );
  NOR2_X1 U6073 ( .A1(n7661), .A2(n7660), .ZN(n4514) );
  NOR2_X1 U6074 ( .A1(n9017), .A2(n9016), .ZN(n4515) );
  NOR2_X1 U6075 ( .A1(n6113), .A2(n6112), .ZN(n4516) );
  INV_X1 U6076 ( .A(n4721), .ZN(n4720) );
  OR2_X1 U6077 ( .A1(n8930), .A2(n4722), .ZN(n4721) );
  AND2_X1 U6078 ( .A1(n9013), .A2(n9014), .ZN(n4517) );
  NOR2_X1 U6079 ( .A1(n8508), .A2(n8166), .ZN(n4518) );
  OR2_X1 U6080 ( .A1(n8435), .A2(n7949), .ZN(n4519) );
  NAND2_X1 U6081 ( .A1(n5281), .A2(n4543), .ZN(n4520) );
  AND2_X1 U6082 ( .A1(n5266), .A2(n4507), .ZN(n4521) );
  AND2_X1 U6083 ( .A1(n5090), .A2(SI_6_), .ZN(n4522) );
  OR2_X1 U6084 ( .A1(n5890), .A2(n5889), .ZN(n4523) );
  INV_X1 U6085 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5211) );
  AND2_X1 U6086 ( .A1(n5876), .A2(n5875), .ZN(n4524) );
  AND2_X1 U6087 ( .A1(n7230), .A2(n7229), .ZN(n4525) );
  NAND2_X1 U6088 ( .A1(n7817), .A2(n6108), .ZN(n4526) );
  AND2_X1 U6089 ( .A1(n4773), .A2(n4770), .ZN(n4527) );
  OR2_X1 U6090 ( .A1(n7679), .A2(n7678), .ZN(n4528) );
  INV_X1 U6091 ( .A(n7312), .ZN(n4833) );
  INV_X1 U6092 ( .A(n6625), .ZN(n7312) );
  INV_X1 U6093 ( .A(n8331), .ZN(n8325) );
  NAND2_X1 U6094 ( .A1(n7968), .A2(n7969), .ZN(n8331) );
  AND2_X1 U6095 ( .A1(n4956), .A2(n4966), .ZN(n4529) );
  NOR2_X1 U6096 ( .A1(n9216), .A2(n9196), .ZN(n4530) );
  OAI21_X1 U6097 ( .B1(n4905), .B2(n4903), .A(n5663), .ZN(n4902) );
  NAND2_X1 U6098 ( .A1(n8893), .A2(n4895), .ZN(n4531) );
  OR2_X1 U6099 ( .A1(n4496), .A2(n4907), .ZN(n4532) );
  NAND2_X1 U6100 ( .A1(n9302), .A2(n4659), .ZN(n4533) );
  AND2_X1 U6101 ( .A1(n4771), .A2(n4770), .ZN(n4534) );
  AND2_X1 U6102 ( .A1(n4529), .A2(n4960), .ZN(n4535) );
  NAND2_X1 U6103 ( .A1(n5257), .A2(n4986), .ZN(n5263) );
  AND2_X1 U6104 ( .A1(n8131), .A2(n4479), .ZN(n4536) );
  AND2_X1 U6105 ( .A1(n4790), .A2(n4486), .ZN(n4537) );
  AND2_X1 U6106 ( .A1(n4691), .A2(n8444), .ZN(n4538) );
  NOR2_X1 U6107 ( .A1(n5722), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n4539) );
  AND2_X1 U6108 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(n5058), .ZN(n4540) );
  AND2_X1 U6109 ( .A1(n5213), .A2(n5039), .ZN(n4541) );
  AND2_X1 U6110 ( .A1(n7950), .A2(n8301), .ZN(n4542) );
  AND2_X1 U6111 ( .A1(n4491), .A2(n5055), .ZN(n4543) );
  NOR2_X1 U6112 ( .A1(n5034), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4675) );
  AND3_X1 U6113 ( .A1(n5257), .A2(n4543), .A3(n4742), .ZN(n5679) );
  OR2_X1 U6114 ( .A1(n4810), .A2(n4807), .ZN(n4544) );
  INV_X1 U6115 ( .A(n8135), .ZN(n5010) );
  INV_X1 U6116 ( .A(n8953), .ZN(n4588) );
  INV_X1 U6117 ( .A(n7666), .ZN(n4958) );
  NAND2_X1 U6118 ( .A1(n5350), .A2(n5349), .ZN(n9417) );
  INV_X1 U6119 ( .A(n9417), .ZN(n4749) );
  OR2_X1 U6120 ( .A1(n7519), .A2(n7829), .ZN(n4545) );
  NAND2_X1 U6121 ( .A1(n4775), .A2(n4774), .ZN(n8511) );
  INV_X2 U6122 ( .A(n5468), .ZN(n7770) );
  INV_X1 U6123 ( .A(n5415), .ZN(n5468) );
  AND2_X1 U6124 ( .A1(n9410), .A2(n9274), .ZN(n4546) );
  NAND2_X1 U6125 ( .A1(n5900), .A2(n5716), .ZN(n5950) );
  INV_X1 U6126 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5739) );
  INV_X1 U6127 ( .A(n8445), .ZN(n4646) );
  AND2_X1 U6128 ( .A1(n6989), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4547) );
  NOR3_X1 U6129 ( .A1(n7519), .A2(n4683), .A3(n8612), .ZN(n4681) );
  NAND2_X1 U6130 ( .A1(n5025), .A2(n5832), .ZN(n5884) );
  AND2_X1 U6131 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n4548) );
  NOR2_X1 U6132 ( .A1(n7537), .A2(n9088), .ZN(n4549) );
  NAND2_X1 U6133 ( .A1(n7549), .A2(n4750), .ZN(n4751) );
  AND2_X1 U6134 ( .A1(n4719), .A2(n4724), .ZN(n4550) );
  AND2_X1 U6135 ( .A1(n4610), .A2(n4609), .ZN(n4551) );
  NOR2_X1 U6136 ( .A1(n9405), .A2(n9286), .ZN(n4552) );
  INV_X1 U6137 ( .A(n7398), .ZN(n9808) );
  AND4_X1 U6138 ( .A1(n5898), .A2(n5897), .A3(n5896), .A4(n5895), .ZN(n7398)
         );
  AND2_X1 U6139 ( .A1(n6298), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4553) );
  AND2_X1 U6140 ( .A1(n4783), .A2(n4479), .ZN(n4554) );
  AND2_X1 U6141 ( .A1(n6255), .A2(n6254), .ZN(n4555) );
  NAND2_X1 U6142 ( .A1(n9367), .A2(n9750), .ZN(n4556) );
  INV_X1 U6143 ( .A(n4909), .ZN(n4907) );
  NAND2_X1 U6144 ( .A1(n9402), .A2(n9273), .ZN(n4909) );
  AND2_X1 U6145 ( .A1(n4775), .A2(n4488), .ZN(n4557) );
  AND2_X1 U6146 ( .A1(n6653), .A2(n6652), .ZN(n4558) );
  NOR2_X1 U6147 ( .A1(n6206), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n6201) );
  AND2_X1 U6148 ( .A1(n4676), .A2(n5832), .ZN(n5900) );
  NAND2_X1 U6149 ( .A1(n6244), .A2(n6232), .ZN(n7944) );
  INV_X1 U6150 ( .A(n7944), .ZN(n7924) );
  AND2_X1 U6151 ( .A1(n7785), .A2(n7967), .ZN(n6231) );
  NAND2_X1 U6152 ( .A1(n6006), .A2(n6005), .ZN(n8612) );
  INV_X1 U6153 ( .A(n8612), .ZN(n4685) );
  NAND2_X1 U6154 ( .A1(n6937), .A2(n7011), .ZN(n7040) );
  AND2_X1 U6155 ( .A1(n7494), .A2(n7493), .ZN(n7613) );
  INV_X1 U6156 ( .A(n8895), .ZN(n4727) );
  NAND2_X1 U6157 ( .A1(n4922), .A2(n6739), .ZN(n6762) );
  OR2_X1 U6158 ( .A1(n7461), .A2(n7463), .ZN(n7494) );
  AND2_X1 U6159 ( .A1(n6909), .A2(n6908), .ZN(n4559) );
  AND2_X1 U6160 ( .A1(n5977), .A2(n5976), .ZN(n4560) );
  INV_X1 U6161 ( .A(n4875), .ZN(n4874) );
  NOR2_X1 U6162 ( .A1(n5378), .A2(n4876), .ZN(n4875) );
  AND2_X1 U6163 ( .A1(n7146), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4561) );
  AND2_X1 U6164 ( .A1(n7372), .A2(n5029), .ZN(n4562) );
  NAND2_X1 U6165 ( .A1(n6066), .A2(n6067), .ZN(n4563) );
  AND2_X1 U6166 ( .A1(n6841), .A2(n5654), .ZN(n4564) );
  AND2_X1 U6167 ( .A1(n5900), .A2(n5032), .ZN(n4565) );
  INV_X1 U6168 ( .A(n6236), .ZN(n8152) );
  XNOR2_X1 U6169 ( .A(n5738), .B(n5737), .ZN(n6236) );
  NAND2_X1 U6170 ( .A1(n5634), .A2(n5633), .ZN(n9351) );
  INV_X1 U6171 ( .A(n6897), .ZN(n4760) );
  INV_X1 U6172 ( .A(n9749), .ZN(n4758) );
  NAND2_X1 U6173 ( .A1(n5672), .A2(n9257), .ZN(n9004) );
  OAI211_X1 U6174 ( .C1(n7233), .C2(n6614), .A(n6365), .B(n6364), .ZN(n6394)
         );
  INV_X1 U6175 ( .A(n5646), .ZN(n8882) );
  AND2_X1 U6176 ( .A1(n4618), .A2(n4485), .ZN(n4566) );
  NAND2_X2 U6177 ( .A1(n7388), .A2(n8133), .ZN(n7512) );
  NAND2_X2 U6178 ( .A1(n7603), .A2(n7602), .ZN(n8515) );
  NAND2_X1 U6179 ( .A1(n4778), .A2(n8310), .ZN(n8326) );
  AND2_X2 U6180 ( .A1(n5899), .A2(n7727), .ZN(n5905) );
  NAND2_X2 U6181 ( .A1(n6975), .A2(n7003), .ZN(n5899) );
  NAND2_X1 U6182 ( .A1(n4783), .A2(n4536), .ZN(n7387) );
  NAND2_X1 U6183 ( .A1(n8292), .A2(n8291), .ZN(n8441) );
  NAND2_X1 U6184 ( .A1(n8425), .A2(n8435), .ZN(n8298) );
  NOR2_X1 U6185 ( .A1(n8257), .A2(n8258), .ZN(n8263) );
  NAND2_X1 U6186 ( .A1(n6997), .A2(n6996), .ZN(n7028) );
  NAND2_X1 U6187 ( .A1(n8180), .A2(n8179), .ZN(n8178) );
  OAI21_X1 U6188 ( .B1(n8271), .B2(n9786), .A(n4710), .ZN(n4709) );
  NOR2_X1 U6189 ( .A1(n7058), .A2(n7057), .ZN(n7056) );
  NOR2_X1 U6190 ( .A1(n7159), .A2(n7158), .ZN(n7157) );
  OAI211_X1 U6191 ( .C1(n8274), .C2(n8273), .A(n4711), .B(n4708), .ZN(P2_U3264) );
  XNOR2_X2 U6192 ( .A(n5794), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9482) );
  NAND2_X1 U6193 ( .A1(n5175), .A2(n5174), .ZN(n5367) );
  NAND2_X1 U6194 ( .A1(n5165), .A2(n5164), .ZN(n5360) );
  NAND2_X1 U6195 ( .A1(n5611), .A2(n9014), .ZN(n9167) );
  AOI211_X2 U6196 ( .C1(n9319), .C2(n9171), .A(n9170), .B(n9169), .ZN(n9373)
         );
  NAND3_X1 U6197 ( .A1(n6257), .A2(n4568), .A3(n4555), .ZN(P2_U3222) );
  NAND2_X1 U6198 ( .A1(n6256), .A2(n8545), .ZN(n4568) );
  NAND2_X4 U6199 ( .A1(n4834), .A2(n7265), .ZN(n6196) );
  OAI21_X2 U6200 ( .B1(n5021), .B2(n4643), .A(n4641), .ZN(n8410) );
  INV_X1 U6201 ( .A(n7515), .ZN(n4648) );
  OAI21_X1 U6202 ( .B1(n6714), .B2(n8126), .A(n7979), .ZN(n6715) );
  NAND2_X2 U6203 ( .A1(n6625), .A2(n6626), .ZN(n8124) );
  NOR2_X1 U6204 ( .A1(n4570), .A2(n4498), .ZN(n4569) );
  NAND2_X1 U6205 ( .A1(n4577), .A2(n4576), .ZN(n9019) );
  NAND3_X1 U6206 ( .A1(n4598), .A2(n8102), .A3(n8101), .ZN(n4597) );
  NAND3_X1 U6207 ( .A1(n8100), .A2(n8325), .A3(n8099), .ZN(n4598) );
  NAND3_X1 U6208 ( .A1(n8156), .A2(n4626), .A3(n4605), .ZN(n4604) );
  XNOR2_X2 U6209 ( .A(n5740), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8273) );
  XNOR2_X1 U6210 ( .A(n9110), .B(n9122), .ZN(n9664) );
  MUX2_X1 U6211 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6272), .S(n6493), .Z(n6496)
         );
  NAND2_X1 U6212 ( .A1(n6578), .A2(n4617), .ZN(n4615) );
  NAND2_X1 U6213 ( .A1(n4615), .A2(n4616), .ZN(n6566) );
  INV_X1 U6214 ( .A(n4618), .ZN(n6576) );
  NAND2_X1 U6215 ( .A1(n4627), .A2(n4629), .ZN(n5106) );
  NAND2_X1 U6216 ( .A1(n5268), .A2(n4631), .ZN(n4627) );
  NAND2_X1 U6217 ( .A1(n5268), .A2(n5267), .ZN(n4637) );
  NAND2_X1 U6218 ( .A1(n9307), .A2(n4655), .ZN(n4651) );
  NAND2_X1 U6219 ( .A1(n4651), .A2(n4650), .ZN(n5662) );
  NAND2_X1 U6220 ( .A1(n6905), .A2(n5653), .ZN(n6842) );
  NAND3_X1 U6221 ( .A1(n6762), .A2(n5652), .A3(n5651), .ZN(n6905) );
  NAND3_X1 U6222 ( .A1(n4668), .A2(n4666), .A3(n4665), .ZN(n9436) );
  INV_X2 U6223 ( .A(n7727), .ZN(n7717) );
  MUX2_X1 U6224 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n7727), .Z(n5079) );
  AND2_X4 U6225 ( .A1(n4670), .A2(n4669), .ZN(n7727) );
  INV_X1 U6226 ( .A(n5041), .ZN(n4671) );
  INV_X1 U6227 ( .A(n4675), .ZN(n4679) );
  INV_X1 U6228 ( .A(n4681), .ZN(n8516) );
  NOR3_X1 U6229 ( .A1(n8365), .A2(n8545), .A3(n8550), .ZN(n8327) );
  AND2_X2 U6230 ( .A1(n8493), .A2(n4538), .ZN(n8426) );
  INV_X1 U6231 ( .A(n8884), .ZN(n6607) );
  NAND2_X1 U6232 ( .A1(n6604), .A2(n8884), .ZN(n6603) );
  NAND2_X1 U6233 ( .A1(n6848), .A2(n8934), .ZN(n4713) );
  NAND2_X1 U6234 ( .A1(n9495), .A2(n8949), .ZN(n9491) );
  AOI21_X1 U6235 ( .B1(n5524), .B2(n4717), .A(n4715), .ZN(n9249) );
  OAI21_X1 U6236 ( .B1(n7527), .B2(n4728), .A(n4725), .ZN(n9342) );
  NOR2_X1 U6237 ( .A1(n4736), .A2(n5210), .ZN(n4742) );
  INV_X1 U6238 ( .A(n5210), .ZN(n4737) );
  NAND4_X1 U6239 ( .A1(n4739), .A2(n4491), .A3(n4738), .A4(n4737), .ZN(n5387)
         );
  INV_X1 U6240 ( .A(n4751), .ZN(n9332) );
  NAND2_X1 U6241 ( .A1(n5678), .A2(n5213), .ZN(n5215) );
  NAND2_X1 U6242 ( .A1(n5678), .A2(n4541), .ZN(n5214) );
  INV_X1 U6243 ( .A(n4757), .ZN(n5045) );
  NAND4_X1 U6244 ( .A1(n6914), .A2(n4759), .A3(n4758), .A4(n9761), .ZN(n9511)
         );
  INV_X1 U6245 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4766) );
  INV_X1 U6246 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4762) );
  AND3_X2 U6247 ( .A1(n4763), .A2(n5779), .A3(n4761), .ZN(n5832) );
  NAND3_X1 U6248 ( .A1(n4763), .A2(n10237), .A3(n5779), .ZN(n5810) );
  NAND2_X1 U6249 ( .A1(n8515), .A2(n4534), .ZN(n4767) );
  NAND2_X1 U6250 ( .A1(n8341), .A2(n4779), .ZN(n4776) );
  NAND2_X1 U6251 ( .A1(n4776), .A2(n4777), .ZN(n8312) );
  NAND2_X1 U6252 ( .A1(n8341), .A2(n8308), .ZN(n4778) );
  AND2_X1 U6253 ( .A1(n7328), .A2(n7327), .ZN(n7330) );
  NAND2_X1 U6254 ( .A1(n4782), .A2(n7289), .ZN(n7328) );
  NAND2_X1 U6255 ( .A1(n8420), .A2(n4542), .ZN(n8390) );
  OAI21_X2 U6256 ( .B1(n8441), .B2(n8293), .A(n8295), .ZN(n8425) );
  NAND2_X1 U6257 ( .A1(n7368), .A2(n4784), .ZN(n4783) );
  NAND2_X1 U6258 ( .A1(n7368), .A2(n7367), .ZN(n9794) );
  INV_X1 U6259 ( .A(n4783), .ZN(n9796) );
  INV_X1 U6260 ( .A(n7367), .ZN(n4785) );
  NAND2_X1 U6261 ( .A1(n7512), .A2(n4537), .ZN(n4788) );
  NAND2_X1 U6262 ( .A1(n7512), .A2(n4497), .ZN(n7513) );
  INV_X1 U6263 ( .A(n4789), .ZN(n7559) );
  INV_X1 U6264 ( .A(n4497), .ZN(n4791) );
  NAND3_X1 U6265 ( .A1(n5900), .A2(n5033), .A3(n4539), .ZN(n4793) );
  AND2_X4 U6266 ( .A1(n5727), .A2(n8655), .ZN(n5822) );
  NAND2_X1 U6267 ( .A1(n4466), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5226) );
  NAND2_X1 U6268 ( .A1(n5774), .A2(n4795), .ZN(n6833) );
  NAND2_X1 U6269 ( .A1(n5762), .A2(n6826), .ZN(n4795) );
  NAND2_X1 U6270 ( .A1(n6070), .A2(n4798), .ZN(n4797) );
  NAND2_X1 U6271 ( .A1(n4814), .A2(n4813), .ZN(n7925) );
  NAND3_X1 U6272 ( .A1(n6143), .A2(n6142), .A3(n6141), .ZN(n7837) );
  NAND2_X1 U6273 ( .A1(n7903), .A2(n4818), .ZN(n4817) );
  NAND2_X1 U6274 ( .A1(n4817), .A2(n4820), .ZN(n7795) );
  NAND2_X1 U6275 ( .A1(n4825), .A2(n5779), .ZN(n5811) );
  NAND2_X1 U6276 ( .A1(n6867), .A2(n6866), .ZN(n6865) );
  NAND2_X1 U6277 ( .A1(n6865), .A2(n4826), .ZN(n5842) );
  NAND2_X1 U6278 ( .A1(n5912), .A2(n4828), .ZN(n6259) );
  NOR2_X2 U6279 ( .A1(n6007), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n6026) );
  NAND2_X1 U6280 ( .A1(n5314), .A2(n4840), .ZN(n4838) );
  NAND2_X1 U6281 ( .A1(n5256), .A2(n4852), .ZN(n4849) );
  NOR2_X1 U6282 ( .A1(n8111), .A2(n4855), .ZN(n8109) );
  NAND2_X1 U6283 ( .A1(n7749), .A2(n7752), .ZN(n4859) );
  NAND2_X1 U6284 ( .A1(n4860), .A2(n4861), .ZN(n5129) );
  NAND2_X1 U6285 ( .A1(n5112), .A2(n4863), .ZN(n4860) );
  NAND2_X1 U6286 ( .A1(n5112), .A2(n5111), .ZN(n5294) );
  OAI21_X1 U6287 ( .B1(n5375), .B2(n4871), .A(n4869), .ZN(n5200) );
  MUX2_X1 U6288 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n7727), .Z(n5224) );
  INV_X1 U6289 ( .A(n5412), .ZN(n4882) );
  NAND2_X1 U6290 ( .A1(n7354), .A2(n4891), .ZN(n4887) );
  OAI21_X1 U6291 ( .B1(n9247), .B2(n4899), .A(n4898), .ZN(n9204) );
  NAND2_X1 U6292 ( .A1(n4897), .A2(n4896), .ZN(n5665) );
  NAND2_X1 U6293 ( .A1(n9247), .A2(n4898), .ZN(n4897) );
  NAND2_X1 U6294 ( .A1(n9390), .A2(n9242), .ZN(n4910) );
  NAND2_X1 U6295 ( .A1(n9175), .A2(n4920), .ZN(n4913) );
  AOI21_X1 U6296 ( .B1(n9175), .B2(n8904), .A(n8905), .ZN(n9157) );
  OAI21_X1 U6297 ( .B1(n9175), .B2(n4916), .A(n4914), .ZN(n7765) );
  NAND2_X1 U6298 ( .A1(n4912), .A2(n4911), .ZN(n7767) );
  NAND2_X1 U6299 ( .A1(n9175), .A2(n4914), .ZN(n4912) );
  NAND2_X1 U6300 ( .A1(n5679), .A2(n4929), .ZN(n5391) );
  NAND2_X1 U6301 ( .A1(n5059), .A2(n4540), .ZN(n4930) );
  OR2_X1 U6302 ( .A1(n5059), .A2(n4934), .ZN(n4931) );
  NAND2_X1 U6303 ( .A1(n5059), .A2(n5058), .ZN(n5060) );
  NAND2_X1 U6304 ( .A1(n8742), .A2(n4937), .ZN(n4936) );
  NAND2_X1 U6305 ( .A1(n4940), .A2(n4941), .ZN(n7620) );
  NAND3_X1 U6306 ( .A1(n6937), .A2(n4473), .A3(n7011), .ZN(n4946) );
  NAND2_X1 U6307 ( .A1(n7667), .A2(n4952), .ZN(n4951) );
  NAND2_X1 U6308 ( .A1(n7667), .A2(n4957), .ZN(n4956) );
  INV_X1 U6309 ( .A(n7667), .ZN(n4959) );
  NAND2_X1 U6310 ( .A1(n7667), .A2(n7666), .ZN(n8682) );
  OAI21_X1 U6311 ( .B1(n8684), .B2(n8685), .A(n8682), .ZN(n8734) );
  NAND2_X1 U6312 ( .A1(n7673), .A2(n7672), .ZN(n4966) );
  OR2_X1 U6313 ( .A1(n5281), .A2(n9451), .ZN(n4967) );
  NAND2_X1 U6314 ( .A1(n4967), .A2(n4968), .ZN(n5057) );
  NAND2_X1 U6315 ( .A1(n5281), .A2(n4970), .ZN(n5064) );
  NAND2_X1 U6316 ( .A1(n6417), .A2(n4971), .ZN(n4972) );
  AND2_X1 U6317 ( .A1(n6652), .A2(n6418), .ZN(n4971) );
  NAND2_X1 U6318 ( .A1(n6417), .A2(n6418), .ZN(n6450) );
  OAI211_X1 U6319 ( .C1(n6449), .C2(n4973), .A(n6659), .B(n4972), .ZN(n6669)
         );
  NAND2_X1 U6320 ( .A1(n4974), .A2(n5235), .ZN(n5251) );
  OAI21_X2 U6321 ( .B1(n8720), .B2(n4979), .A(n4977), .ZN(n7639) );
  NOR2_X2 U6322 ( .A1(n7639), .A2(n7638), .ZN(n8774) );
  INV_X1 U6323 ( .A(n8717), .ZN(n4984) );
  NAND2_X1 U6324 ( .A1(n5257), .A2(n4985), .ZN(n5274) );
  NAND2_X1 U6325 ( .A1(n5905), .A2(n4989), .ZN(n4988) );
  NAND2_X1 U6326 ( .A1(n5899), .A2(n5770), .ZN(n5793) );
  NAND3_X1 U6327 ( .A1(n5835), .A2(n5836), .A3(n4990), .ZN(n7246) );
  NAND2_X1 U6328 ( .A1(n7999), .A2(n7981), .ZN(n7285) );
  NAND2_X1 U6329 ( .A1(n7952), .A2(n5001), .ZN(n4997) );
  NAND2_X1 U6330 ( .A1(n4997), .A2(n4998), .ZN(n7961) );
  NAND2_X1 U6331 ( .A1(n7952), .A2(n5006), .ZN(n5000) );
  NAND2_X1 U6332 ( .A1(n7952), .A2(n8098), .ZN(n8332) );
  NAND2_X1 U6333 ( .A1(n8472), .A2(n4489), .ZN(n5021) );
  INV_X1 U6334 ( .A(n8351), .ZN(n8360) );
  NAND2_X1 U6335 ( .A1(n7338), .A2(n4504), .ZN(n5028) );
  NAND2_X1 U6336 ( .A1(n5028), .A2(n5026), .ZN(n7389) );
  NAND2_X1 U6337 ( .A1(n5676), .A2(n5675), .ZN(n5677) );
  INV_X1 U6338 ( .A(n9156), .ZN(n5676) );
  CLKBUF_X1 U6339 ( .A(n6786), .Z(n6791) );
  NAND2_X1 U6340 ( .A1(n6235), .A2(n4688), .ZN(n6257) );
  INV_X1 U6341 ( .A(n6026), .ZN(n6027) );
  INV_X1 U6342 ( .A(n5421), .ZN(n5627) );
  AND2_X1 U6343 ( .A1(n6237), .A2(n7924), .ZN(n6235) );
  OR2_X1 U6344 ( .A1(n5059), .A2(n5058), .ZN(n5061) );
  AND2_X1 U6345 ( .A1(n7004), .A2(n7003), .ZN(n9483) );
  NAND2_X1 U6346 ( .A1(n9078), .A2(n5671), .ZN(n9036) );
  OAI211_X1 U6347 ( .C1(n7961), .C2(n8280), .A(n5748), .B(n7954), .ZN(n7963)
         );
  AOI22_X1 U6348 ( .A1(n8286), .A2(n8285), .B1(n8284), .B2(n8492), .ZN(n8469)
         );
  INV_X1 U6349 ( .A(n6933), .ZN(n6936) );
  AND4_X2 U6350 ( .A1(n5731), .A2(n5730), .A3(n5729), .A4(n5728), .ZN(n6807)
         );
  NAND2_X1 U6351 ( .A1(n6535), .A2(n5672), .ZN(n6359) );
  AND2_X4 U6352 ( .A1(n5395), .A2(n9458), .ZN(n5422) );
  NOR2_X1 U6353 ( .A1(n6715), .A2(n8118), .ZN(n7277) );
  OR2_X1 U6354 ( .A1(n8117), .A2(n6231), .ZN(n5035) );
  AND2_X1 U6355 ( .A1(n5743), .A2(n5742), .ZN(n5036) );
  NAND2_X2 U6356 ( .A1(n6258), .A2(n9850), .ZN(n8176) );
  AND2_X1 U6357 ( .A1(n8352), .A2(n8350), .ZN(n5038) );
  NAND2_X1 U6358 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n5039) );
  OR2_X1 U6359 ( .A1(n9269), .A2(n9251), .ZN(n5040) );
  NAND2_X1 U6360 ( .A1(n5630), .A2(n5629), .ZN(n9171) );
  NAND2_X1 U6361 ( .A1(n5619), .A2(n5618), .ZN(n9186) );
  OR2_X1 U6362 ( .A1(n9036), .A2(n5635), .ZN(n9502) );
  AND4_X1 U6363 ( .A1(n6002), .A2(n6001), .A3(n6000), .A4(n5999), .ZN(n7849)
         );
  INV_X1 U6364 ( .A(n9185), .ZN(n9208) );
  NAND2_X1 U6365 ( .A1(n5600), .A2(n5599), .ZN(n9185) );
  XNOR2_X1 U6366 ( .A(n5746), .B(P2_IR_REG_21__SCAN_IN), .ZN(n5748) );
  NAND2_X1 U6367 ( .A1(n6694), .A2(n5646), .ZN(n6693) );
  AND4_X1 U6368 ( .A1(n5959), .A2(n5958), .A3(n5957), .A4(n5956), .ZN(n7906)
         );
  INV_X1 U6369 ( .A(n5670), .ZN(n5632) );
  AND4_X1 U6370 ( .A1(n9039), .A2(n5671), .A3(n9067), .A4(n5672), .ZN(n5042)
         );
  NAND2_X1 U6371 ( .A1(n9073), .A2(n9257), .ZN(n5043) );
  INV_X1 U6372 ( .A(n8422), .ZN(n8299) );
  NOR3_X1 U6373 ( .A1(n9193), .A2(n8903), .A3(n8902), .ZN(n5044) );
  INV_X1 U6374 ( .A(n9430), .ZN(n5329) );
  INV_X1 U6375 ( .A(n9534), .ZN(n5675) );
  INV_X2 U6376 ( .A(n9768), .ZN(n9759) );
  INV_X1 U6377 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5877) );
  NOR2_X1 U6378 ( .A1(n9541), .A2(n7542), .ZN(n5660) );
  INV_X1 U6379 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5913) );
  INV_X1 U6380 ( .A(n7849), .ZN(n7604) );
  OR2_X1 U6381 ( .A1(n5878), .A2(n5877), .ZN(n5893) );
  INV_X1 U6382 ( .A(n8120), .ZN(n7291) );
  OAI21_X1 U6383 ( .B1(n6206), .B2(n5722), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5723) );
  INV_X1 U6384 ( .A(n6934), .ZN(n6935) );
  INV_X1 U6385 ( .A(n5550), .ZN(n5548) );
  INV_X1 U6386 ( .A(n5517), .ZN(n5516) );
  INV_X1 U6387 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5508) );
  INV_X1 U6388 ( .A(SI_23_), .ZN(n5178) );
  INV_X1 U6389 ( .A(SI_20_), .ZN(n5160) );
  OR2_X1 U6390 ( .A1(n5339), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n5340) );
  INV_X1 U6391 ( .A(SI_13_), .ZN(n5124) );
  OR2_X1 U6392 ( .A1(n5914), .A2(n5913), .ZN(n5938) );
  INV_X1 U6393 ( .A(n6788), .ZN(n6628) );
  INV_X1 U6394 ( .A(n8177), .ZN(n6639) );
  INV_X1 U6395 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5967) );
  INV_X1 U6396 ( .A(n6262), .ZN(n5930) );
  INV_X1 U6397 ( .A(n5822), .ZN(n6178) );
  INV_X1 U6398 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10132) );
  INV_X1 U6399 ( .A(n7906), .ZN(n7558) );
  AOI21_X1 U6400 ( .B1(n8119), .B2(n6804), .A(n6640), .ZN(n6714) );
  NAND2_X1 U6401 ( .A1(n8333), .A2(n9807), .ZN(n8336) );
  NAND2_X1 U6402 ( .A1(n8486), .A2(n8059), .ZN(n7946) );
  NAND2_X1 U6403 ( .A1(n6209), .A2(n6208), .ZN(n6210) );
  INV_X1 U6404 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U6405 ( .A1(n6936), .A2(n6935), .ZN(n7011) );
  OR2_X1 U6406 ( .A1(n5613), .A2(n5612), .ZN(n5622) );
  OR2_X1 U6407 ( .A1(n5593), .A2(n5592), .ZN(n5603) );
  OR3_X1 U6408 ( .A1(n5565), .A2(n5564), .A3(n5563), .ZN(n5574) );
  INV_X1 U6409 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U6410 ( .A1(n5516), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5532) );
  INV_X1 U6411 ( .A(n9171), .ZN(n7764) );
  AND2_X1 U6412 ( .A1(n8842), .A2(n8836), .ZN(n8895) );
  INV_X1 U6413 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5056) );
  OR2_X1 U6414 ( .A1(n6060), .A2(n6059), .ZN(n6075) );
  OR2_X1 U6415 ( .A1(n7863), .A2(n7867), .ZN(n6141) );
  NAND2_X1 U6416 ( .A1(n6639), .A2(n9852), .ZN(n6770) );
  NAND2_X1 U6417 ( .A1(n6031), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U6418 ( .A1(n5985), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6013) );
  AND2_X1 U6419 ( .A1(n6238), .A2(n6191), .ZN(n8328) );
  INV_X1 U6420 ( .A(n6972), .ZN(n6634) );
  AND2_X1 U6421 ( .A1(n5747), .A2(n5748), .ZN(n6972) );
  NAND2_X1 U6422 ( .A1(n7398), .A2(n7385), .ZN(n7386) );
  NAND2_X1 U6423 ( .A1(n9823), .A2(n8625), .ZN(n9836) );
  INV_X1 U6424 ( .A(n9907), .ZN(n8625) );
  NAND2_X1 U6425 ( .A1(n7330), .A2(n7329), .ZN(n7368) );
  OR3_X1 U6426 ( .A1(n8152), .A2(n5747), .A3(n8149), .ZN(n9878) );
  INV_X1 U6427 ( .A(n9186), .ZN(n7705) );
  INV_X1 U6428 ( .A(n9093), .ZN(n7198) );
  AND2_X1 U6429 ( .A1(n6416), .A2(n6415), .ZN(n8764) );
  OR2_X1 U6430 ( .A1(n6421), .A2(n5635), .ZN(n8778) );
  INV_X1 U6431 ( .A(n8789), .ZN(n8805) );
  OR2_X1 U6432 ( .A1(n5532), .A2(n5531), .ZN(n5534) );
  OR2_X1 U6433 ( .A1(n5419), .A2(n5398), .ZN(n5399) );
  INV_X1 U6434 ( .A(n9116), .ZN(n9690) );
  INV_X1 U6435 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8699) );
  INV_X1 U6436 ( .A(n9230), .ZN(n9196) );
  INV_X1 U6437 ( .A(n9286), .ZN(n9251) );
  AND2_X1 U6438 ( .A1(n8983), .A2(n8982), .ZN(n9327) );
  AND2_X1 U6439 ( .A1(n8978), .A2(n8979), .ZN(n9345) );
  INV_X1 U6440 ( .A(n9351), .ZN(n9497) );
  AND2_X1 U6441 ( .A1(n5674), .A2(n5673), .ZN(n9347) );
  NAND2_X1 U6442 ( .A1(n5219), .A2(n5218), .ZN(n5221) );
  AND2_X1 U6443 ( .A1(n5111), .A2(n5110), .ZN(n5285) );
  OR2_X1 U6444 ( .A1(n7929), .A2(n8474), .ZN(n7937) );
  AND2_X1 U6445 ( .A1(n6176), .A2(n6162), .ZN(n8367) );
  NOR2_X1 U6446 ( .A1(n6248), .A2(n9844), .ZN(n6244) );
  AOI21_X1 U6447 ( .B1(n8328), .B2(n5822), .A(n6195), .ZN(n8311) );
  AND4_X1 U6448 ( .A1(n6037), .A2(n6036), .A3(n6035), .A4(n6034), .ZN(n7918)
         );
  INV_X1 U6449 ( .A(n9786), .ZN(n9782) );
  AND2_X1 U6450 ( .A1(n6999), .A2(n6976), .ZN(n9783) );
  INV_X1 U6451 ( .A(n9836), .ZN(n8527) );
  NOR2_X1 U6452 ( .A1(n9847), .A2(n6227), .ZN(n6704) );
  NAND2_X1 U6453 ( .A1(n8159), .A2(n6231), .ZN(n9905) );
  INV_X1 U6454 ( .A(n9912), .ZN(n9864) );
  INV_X1 U6455 ( .A(n9813), .ZN(n9857) );
  AND2_X1 U6456 ( .A1(n6003), .A2(n5982), .ZN(n8192) );
  NAND2_X1 U6457 ( .A1(n6386), .A2(n6385), .ZN(n8802) );
  OR2_X1 U6458 ( .A1(n9177), .A2(n5636), .ZN(n5610) );
  INV_X1 U6459 ( .A(n5422), .ZN(n5636) );
  NOR2_X1 U6460 ( .A1(n6284), .A2(n5635), .ZN(n9687) );
  INV_X1 U6461 ( .A(n9712), .ZN(n9693) );
  INV_X1 U6462 ( .A(n9691), .ZN(n9707) );
  OR2_X1 U6463 ( .A1(n8998), .A2(n8878), .ZN(n9262) );
  INV_X1 U6464 ( .A(n9347), .ZN(n9506) );
  INV_X1 U6465 ( .A(n9502), .ZN(n9317) );
  INV_X1 U6466 ( .A(n6432), .ZN(n6433) );
  OR2_X1 U6467 ( .A1(n6536), .A2(n5632), .ZN(n9762) );
  AND2_X1 U6468 ( .A1(n9347), .A2(n9756), .ZN(n9534) );
  OR2_X1 U6469 ( .A1(n5695), .A2(n6369), .ZN(n6434) );
  INV_X1 U6470 ( .A(n9756), .ZN(n9767) );
  AND2_X1 U6471 ( .A1(n5295), .A2(n5290), .ZN(n6510) );
  INV_X1 U6472 ( .A(n8277), .ZN(n9788) );
  INV_X1 U6473 ( .A(n8562), .ZN(n8387) );
  INV_X1 U6474 ( .A(n8287), .ZN(n8464) );
  INV_X1 U6475 ( .A(n9783), .ZN(n8224) );
  AND2_X1 U6476 ( .A1(n6355), .A2(n6354), .ZN(n8277) );
  NAND2_X1 U6477 ( .A1(n9840), .A2(n9833), .ZN(n8529) );
  INV_X1 U6478 ( .A(n9927), .ZN(n9924) );
  INV_X1 U6479 ( .A(n9915), .ZN(n9913) );
  NOR2_X1 U6480 ( .A1(n9844), .A2(n9843), .ZN(n9845) );
  AND2_X1 U6481 ( .A1(n7571), .A2(n7595), .ZN(n9847) );
  XNOR2_X1 U6482 ( .A(n6213), .B(n6212), .ZN(n7571) );
  INV_X1 U6483 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6458) );
  INV_X1 U6484 ( .A(n8654), .ZN(n8661) );
  INV_X1 U6485 ( .A(n8807), .ZN(n8750) );
  OR3_X1 U6486 ( .A1(n6376), .A2(n9750), .A3(n6368), .ZN(n8782) );
  NAND2_X1 U6487 ( .A1(n5591), .A2(n5590), .ZN(n9230) );
  INV_X1 U6488 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9617) );
  INV_X1 U6489 ( .A(n9687), .ZN(n9701) );
  NAND2_X1 U6490 ( .A1(n6308), .A2(n6307), .ZN(n9716) );
  AND2_X1 U6491 ( .A1(n7532), .A2(n7531), .ZN(n9546) );
  OR2_X1 U6492 ( .A1(n9519), .A2(n6764), .ZN(n9340) );
  INV_X1 U6493 ( .A(n9338), .ZN(n9312) );
  OR2_X1 U6494 ( .A1(n6434), .A2(n6433), .ZN(n9779) );
  AND2_X1 U6495 ( .A1(n9546), .A2(n9545), .ZN(n9567) );
  OR2_X1 U6496 ( .A1(n6434), .A2(n6521), .ZN(n9768) );
  AND2_X1 U6497 ( .A1(n9722), .A2(n9717), .ZN(n9718) );
  AND3_X1 U6498 ( .A1(n7473), .A2(P1_STATE_REG_SCAN_IN), .A3(n6382), .ZN(n9722) );
  INV_X1 U6499 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10223) );
  INV_X1 U6500 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6459) );
  INV_X1 U6501 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6334) );
  INV_X1 U6502 ( .A(n9463), .ZN(n7760) );
  NOR2_X1 U6503 ( .A1(n9957), .A2(n9956), .ZN(n9955) );
  INV_X1 U6504 ( .A(n8176), .ZN(P2_U3966) );
  INV_X1 U6505 ( .A(n9100), .ZN(P1_U4006) );
  NAND2_X1 U6506 ( .A1(n5712), .A2(n5711), .ZN(P1_U3519) );
  NOR2_X2 U6507 ( .A1(n5274), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5281) );
  NAND2_X1 U6508 ( .A1(n5061), .A2(n5060), .ZN(n5669) );
  NAND2_X1 U6509 ( .A1(n5672), .A2(n5062), .ZN(n6536) );
  NAND2_X1 U6510 ( .A1(n4520), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5063) );
  MUX2_X1 U6511 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5063), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n5065) );
  AND2_X1 U6512 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5070) );
  NAND2_X1 U6513 ( .A1(n7727), .A2(n5070), .ZN(n5772) );
  AND2_X1 U6514 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n5071) );
  NAND2_X1 U6515 ( .A1(n5072), .A2(SI_1_), .ZN(n5073) );
  INV_X1 U6516 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5074) );
  INV_X1 U6517 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6317) );
  MUX2_X1 U6518 ( .A(n5074), .B(n6317), .S(n5094), .Z(n5075) );
  XNOR2_X1 U6519 ( .A(n5075), .B(SI_2_), .ZN(n5232) );
  NAND2_X1 U6520 ( .A1(n5233), .A2(n5232), .ZN(n5078) );
  INV_X1 U6521 ( .A(n5075), .ZN(n5076) );
  NAND2_X1 U6522 ( .A1(n5076), .A2(SI_2_), .ZN(n5077) );
  NAND2_X1 U6523 ( .A1(n5078), .A2(n5077), .ZN(n5243) );
  INV_X1 U6524 ( .A(SI_3_), .ZN(n10193) );
  XNOR2_X1 U6525 ( .A(n5079), .B(n10193), .ZN(n5242) );
  NAND2_X1 U6526 ( .A1(n5243), .A2(n5242), .ZN(n5081) );
  NAND2_X1 U6527 ( .A1(n5079), .A2(SI_3_), .ZN(n5080) );
  NAND2_X1 U6528 ( .A1(n5081), .A2(n5080), .ZN(n5250) );
  INV_X1 U6529 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6320) );
  MUX2_X1 U6530 ( .A(n6320), .B(n10226), .S(n7717), .Z(n5082) );
  XNOR2_X1 U6531 ( .A(n5082), .B(SI_4_), .ZN(n5249) );
  NAND2_X1 U6532 ( .A1(n5250), .A2(n5249), .ZN(n5085) );
  INV_X1 U6533 ( .A(n5082), .ZN(n5083) );
  NAND2_X1 U6534 ( .A1(n5083), .A2(SI_4_), .ZN(n5084) );
  INV_X1 U6535 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n5086) );
  MUX2_X1 U6536 ( .A(n6324), .B(n5086), .S(n7717), .Z(n5087) );
  XNOR2_X1 U6537 ( .A(n5087), .B(SI_5_), .ZN(n5255) );
  INV_X1 U6538 ( .A(n5087), .ZN(n5088) );
  NAND2_X1 U6539 ( .A1(n5088), .A2(SI_5_), .ZN(n5089) );
  MUX2_X1 U6540 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7717), .Z(n5090) );
  INV_X1 U6541 ( .A(SI_6_), .ZN(n10154) );
  XNOR2_X1 U6542 ( .A(n5090), .B(n10154), .ZN(n5265) );
  INV_X1 U6543 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6329) );
  MUX2_X1 U6544 ( .A(n6329), .B(n10185), .S(n7717), .Z(n5091) );
  XNOR2_X1 U6545 ( .A(n5091), .B(SI_7_), .ZN(n5267) );
  INV_X1 U6546 ( .A(n5091), .ZN(n5092) );
  NAND2_X1 U6547 ( .A1(n5092), .A2(SI_7_), .ZN(n5093) );
  MUX2_X1 U6548 ( .A(n6330), .B(n6332), .S(n5770), .Z(n5096) );
  INV_X1 U6549 ( .A(SI_8_), .ZN(n5095) );
  NAND2_X1 U6550 ( .A1(n5096), .A2(n5095), .ZN(n5100) );
  INV_X1 U6551 ( .A(n5096), .ZN(n5097) );
  NAND2_X1 U6552 ( .A1(n5097), .A2(SI_8_), .ZN(n5098) );
  INV_X1 U6553 ( .A(n5272), .ZN(n5099) );
  MUX2_X1 U6554 ( .A(n6337), .B(n6334), .S(n7717), .Z(n5102) );
  INV_X1 U6555 ( .A(SI_9_), .ZN(n5101) );
  NAND2_X1 U6556 ( .A1(n5102), .A2(n5101), .ZN(n5105) );
  INV_X1 U6557 ( .A(n5102), .ZN(n5103) );
  NAND2_X1 U6558 ( .A1(n5103), .A2(SI_9_), .ZN(n5104) );
  NAND2_X1 U6559 ( .A1(n5106), .A2(n5105), .ZN(n5286) );
  MUX2_X1 U6560 ( .A(n10246), .B(n6341), .S(n7717), .Z(n5108) );
  NAND2_X1 U6561 ( .A1(n5108), .A2(n5107), .ZN(n5111) );
  INV_X1 U6562 ( .A(n5108), .ZN(n5109) );
  NAND2_X1 U6563 ( .A1(n5109), .A2(SI_10_), .ZN(n5110) );
  MUX2_X1 U6564 ( .A(n5113), .B(n6344), .S(n5770), .Z(n5114) );
  XNOR2_X1 U6565 ( .A(n5114), .B(SI_11_), .ZN(n5293) );
  INV_X1 U6566 ( .A(n5293), .ZN(n5117) );
  INV_X1 U6567 ( .A(n5114), .ZN(n5115) );
  NAND2_X1 U6568 ( .A1(n5115), .A2(SI_11_), .ZN(n5116) );
  MUX2_X1 U6569 ( .A(n6347), .B(n10266), .S(n7717), .Z(n5119) );
  NAND2_X1 U6570 ( .A1(n5119), .A2(n5118), .ZN(n5122) );
  INV_X1 U6571 ( .A(n5119), .ZN(n5120) );
  NAND2_X1 U6572 ( .A1(n5120), .A2(SI_12_), .ZN(n5121) );
  NAND2_X1 U6573 ( .A1(n5122), .A2(n5121), .ZN(n5299) );
  MUX2_X1 U6574 ( .A(n6351), .B(n5123), .S(n5770), .Z(n5125) );
  NAND2_X1 U6575 ( .A1(n5125), .A2(n5124), .ZN(n5128) );
  INV_X1 U6576 ( .A(n5125), .ZN(n5126) );
  NAND2_X1 U6577 ( .A1(n5126), .A2(SI_13_), .ZN(n5127) );
  NAND2_X1 U6578 ( .A1(n5129), .A2(n5128), .ZN(n5314) );
  MUX2_X1 U6579 ( .A(n10095), .B(n10102), .S(n5770), .Z(n5130) );
  XNOR2_X1 U6580 ( .A(n5130), .B(SI_14_), .ZN(n5313) );
  INV_X1 U6581 ( .A(n5313), .ZN(n5133) );
  INV_X1 U6582 ( .A(n5130), .ZN(n5131) );
  NAND2_X1 U6583 ( .A1(n5131), .A2(SI_14_), .ZN(n5132) );
  MUX2_X1 U6584 ( .A(n6458), .B(n6459), .S(n7717), .Z(n5135) );
  NAND2_X1 U6585 ( .A1(n5135), .A2(n5134), .ZN(n5138) );
  INV_X1 U6586 ( .A(n5135), .ZN(n5136) );
  NAND2_X1 U6587 ( .A1(n5136), .A2(SI_15_), .ZN(n5137) );
  NAND2_X1 U6588 ( .A1(n5138), .A2(n5137), .ZN(n5323) );
  MUX2_X1 U6589 ( .A(n5140), .B(n5139), .S(n5770), .Z(n5142) );
  NAND2_X1 U6590 ( .A1(n5142), .A2(n5141), .ZN(n5145) );
  INV_X1 U6591 ( .A(n5142), .ZN(n5143) );
  NAND2_X1 U6592 ( .A1(n5143), .A2(SI_16_), .ZN(n5144) );
  MUX2_X1 U6593 ( .A(n6710), .B(n5146), .S(n5770), .Z(n5147) );
  XNOR2_X1 U6594 ( .A(n5147), .B(SI_17_), .ZN(n5337) );
  INV_X1 U6595 ( .A(n5337), .ZN(n5150) );
  INV_X1 U6596 ( .A(n5147), .ZN(n5148) );
  NAND2_X1 U6597 ( .A1(n5148), .A2(SI_17_), .ZN(n5149) );
  MUX2_X1 U6598 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5770), .Z(n5152) );
  XNOR2_X1 U6599 ( .A(n5152), .B(SI_18_), .ZN(n5345) );
  INV_X1 U6600 ( .A(n5345), .ZN(n5151) );
  NAND2_X1 U6601 ( .A1(n5346), .A2(n5151), .ZN(n5154) );
  NAND2_X1 U6602 ( .A1(n5152), .A2(SI_18_), .ZN(n5153) );
  MUX2_X1 U6603 ( .A(n7600), .B(n6924), .S(n7717), .Z(n5156) );
  INV_X1 U6604 ( .A(SI_19_), .ZN(n5155) );
  NAND2_X1 U6605 ( .A1(n5156), .A2(n5155), .ZN(n5159) );
  INV_X1 U6606 ( .A(n5156), .ZN(n5157) );
  NAND2_X1 U6607 ( .A1(n5157), .A2(SI_19_), .ZN(n5158) );
  NAND2_X1 U6608 ( .A1(n5159), .A2(n5158), .ZN(n5351) );
  MUX2_X1 U6609 ( .A(n7086), .B(n10222), .S(n5770), .Z(n5161) );
  NAND2_X1 U6610 ( .A1(n5161), .A2(n5160), .ZN(n5164) );
  INV_X1 U6611 ( .A(n5161), .ZN(n5162) );
  NAND2_X1 U6612 ( .A1(n5162), .A2(SI_20_), .ZN(n5163) );
  NAND2_X1 U6613 ( .A1(n5356), .A2(n5355), .ZN(n5165) );
  MUX2_X1 U6614 ( .A(n7090), .B(n7761), .S(n7717), .Z(n5167) );
  XNOR2_X1 U6615 ( .A(n5167), .B(SI_21_), .ZN(n5359) );
  INV_X1 U6616 ( .A(n5359), .ZN(n5166) );
  INV_X1 U6617 ( .A(n5167), .ZN(n5168) );
  NAND2_X1 U6618 ( .A1(n5168), .A2(SI_21_), .ZN(n5169) );
  MUX2_X1 U6619 ( .A(n10128), .B(n7471), .S(n5770), .Z(n5171) );
  INV_X1 U6620 ( .A(SI_22_), .ZN(n5170) );
  NAND2_X1 U6621 ( .A1(n5171), .A2(n5170), .ZN(n5174) );
  INV_X1 U6622 ( .A(n5171), .ZN(n5172) );
  NAND2_X1 U6623 ( .A1(n5172), .A2(SI_22_), .ZN(n5173) );
  NAND2_X1 U6624 ( .A1(n5174), .A2(n5173), .ZN(n5363) );
  INV_X1 U6625 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5177) );
  INV_X1 U6626 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5176) );
  MUX2_X1 U6627 ( .A(n5177), .B(n5176), .S(n5770), .Z(n5179) );
  NAND2_X1 U6628 ( .A1(n5179), .A2(n5178), .ZN(n5183) );
  INV_X1 U6629 ( .A(n5179), .ZN(n5180) );
  NAND2_X1 U6630 ( .A1(n5180), .A2(SI_23_), .ZN(n5181) );
  NAND2_X1 U6631 ( .A1(n5183), .A2(n5181), .ZN(n5368) );
  INV_X1 U6632 ( .A(n5368), .ZN(n5182) );
  NAND2_X1 U6633 ( .A1(n5367), .A2(n5182), .ZN(n5370) );
  NAND2_X1 U6634 ( .A1(n5370), .A2(n5183), .ZN(n5375) );
  MUX2_X1 U6635 ( .A(n10120), .B(n10223), .S(n7717), .Z(n5184) );
  XNOR2_X1 U6636 ( .A(n5184), .B(SI_24_), .ZN(n5374) );
  INV_X1 U6637 ( .A(n5374), .ZN(n5187) );
  INV_X1 U6638 ( .A(n5184), .ZN(n5185) );
  NAND2_X1 U6639 ( .A1(n5185), .A2(SI_24_), .ZN(n5186) );
  INV_X1 U6640 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n10104) );
  INV_X1 U6641 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n5188) );
  MUX2_X1 U6642 ( .A(n10104), .B(n5188), .S(n7717), .Z(n5190) );
  INV_X1 U6643 ( .A(SI_25_), .ZN(n5189) );
  NAND2_X1 U6644 ( .A1(n5190), .A2(n5189), .ZN(n5193) );
  INV_X1 U6645 ( .A(n5190), .ZN(n5191) );
  NAND2_X1 U6646 ( .A1(n5191), .A2(SI_25_), .ZN(n5192) );
  NAND2_X1 U6647 ( .A1(n5193), .A2(n5192), .ZN(n5378) );
  INV_X1 U6648 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7594) );
  INV_X1 U6649 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n5194) );
  MUX2_X1 U6650 ( .A(n7594), .B(n5194), .S(n5770), .Z(n5196) );
  INV_X1 U6651 ( .A(SI_26_), .ZN(n5195) );
  NAND2_X1 U6652 ( .A1(n5196), .A2(n5195), .ZN(n5199) );
  INV_X1 U6653 ( .A(n5196), .ZN(n5197) );
  NAND2_X1 U6654 ( .A1(n5197), .A2(SI_26_), .ZN(n5198) );
  NAND2_X1 U6655 ( .A1(n5200), .A2(n5199), .ZN(n5219) );
  INV_X1 U6656 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7710) );
  INV_X1 U6657 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5201) );
  MUX2_X1 U6658 ( .A(n7710), .B(n5201), .S(n7717), .Z(n5203) );
  INV_X1 U6659 ( .A(SI_27_), .ZN(n5202) );
  NAND2_X1 U6660 ( .A1(n5203), .A2(n5202), .ZN(n5206) );
  INV_X1 U6661 ( .A(n5203), .ZN(n5204) );
  NAND2_X1 U6662 ( .A1(n5204), .A2(SI_27_), .ZN(n5205) );
  INV_X1 U6663 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n10118) );
  INV_X1 U6664 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5207) );
  MUX2_X1 U6665 ( .A(n10118), .B(n5207), .S(n5770), .Z(n7714) );
  XNOR2_X1 U6666 ( .A(n7714), .B(SI_28_), .ZN(n7711) );
  NOR2_X1 U6667 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5209) );
  NOR2_X1 U6668 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5208) );
  NAND4_X1 U6669 ( .A1(n5690), .A2(n5209), .A3(n5208), .A4(n5692), .ZN(n5210)
         );
  INV_X1 U6670 ( .A(n5389), .ZN(n5212) );
  NAND2_X1 U6671 ( .A1(n5212), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5213) );
  XNOR2_X2 U6672 ( .A(n5214), .B(P1_IR_REG_28__SCAN_IN), .ZN(n5635) );
  XNOR2_X2 U6673 ( .A(n5215), .B(P1_IR_REG_27__SCAN_IN), .ZN(n9074) );
  NAND2_X2 U6674 ( .A1(n5635), .A2(n9074), .ZN(n5228) );
  NAND2_X2 U6675 ( .A1(n5228), .A2(n7717), .ZN(n5241) );
  NAND2_X1 U6676 ( .A1(n9462), .A2(n7739), .ZN(n5217) );
  NAND2_X1 U6677 ( .A1(n5234), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5216) );
  OR2_X1 U6678 ( .A1(n5219), .A2(n5218), .ZN(n5220) );
  NAND2_X1 U6679 ( .A1(n5221), .A2(n5220), .ZN(n7596) );
  NAND2_X1 U6680 ( .A1(n7596), .A2(n7739), .ZN(n5223) );
  NAND2_X1 U6681 ( .A1(n5234), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5222) );
  INV_X1 U6682 ( .A(n9370), .ZN(n9163) );
  XNOR2_X1 U6683 ( .A(n5225), .B(n5224), .ZN(n5755) );
  INV_X1 U6684 ( .A(n5755), .ZN(n6314) );
  INV_X1 U6685 ( .A(n5228), .ZN(n5244) );
  NAND2_X1 U6686 ( .A1(n5244), .A2(n6493), .ZN(n5227) );
  INV_X1 U6687 ( .A(SI_0_), .ZN(n5769) );
  INV_X1 U6688 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n10106) );
  OAI21_X1 U6689 ( .B1(n7727), .B2(n5769), .A(n10106), .ZN(n5230) );
  AND2_X1 U6690 ( .A1(n5230), .A2(n5229), .ZN(n9466) );
  XNOR2_X1 U6691 ( .A(n5233), .B(n5232), .ZN(n6316) );
  NAND2_X1 U6692 ( .A1(n4465), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5240) );
  NOR2_X1 U6693 ( .A1(n5235), .A2(n9451), .ZN(n5236) );
  MUX2_X1 U6694 ( .A(n9451), .B(n5236), .S(P1_IR_REG_2__SCAN_IN), .Z(n5238) );
  NOR2_X1 U6695 ( .A1(n5238), .A2(n5237), .ZN(n6292) );
  NAND2_X1 U6696 ( .A1(n5244), .A2(n6292), .ZN(n5239) );
  NAND2_X1 U6697 ( .A1(n6613), .A2(n9732), .ZN(n9729) );
  XNOR2_X1 U6698 ( .A(n5243), .B(n5242), .ZN(n6318) );
  NAND2_X1 U6699 ( .A1(n5234), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5248) );
  INV_X1 U6700 ( .A(n5237), .ZN(n5245) );
  NAND2_X1 U6701 ( .A1(n5245), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5246) );
  XNOR2_X1 U6702 ( .A(n5246), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6481) );
  NAND2_X1 U6703 ( .A1(n6270), .A2(n6481), .ZN(n5247) );
  OR2_X1 U6704 ( .A1(n9729), .A2(n6587), .ZN(n6745) );
  XNOR2_X1 U6705 ( .A(n5250), .B(n5249), .ZN(n6321) );
  NAND2_X1 U6706 ( .A1(n5234), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U6707 ( .A1(n5251), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5252) );
  XNOR2_X1 U6708 ( .A(n5252), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U6709 ( .A1(n6270), .A2(n6296), .ZN(n5253) );
  OAI211_X1 U6710 ( .C1(n5241), .C2(n6321), .A(n5254), .B(n5253), .ZN(n6747)
         );
  OR2_X1 U6711 ( .A1(n6745), .A2(n6747), .ZN(n6755) );
  XNOR2_X1 U6712 ( .A(n5256), .B(n5255), .ZN(n6323) );
  NAND2_X1 U6713 ( .A1(n5234), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5260) );
  OR2_X1 U6714 ( .A1(n5257), .A2(n9451), .ZN(n5258) );
  XNOR2_X1 U6715 ( .A(n5258), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6583) );
  NAND2_X1 U6716 ( .A1(n6270), .A2(n6583), .ZN(n5259) );
  NOR2_X2 U6717 ( .A1(n6755), .A2(n6879), .ZN(n6914) );
  NOR2_X1 U6718 ( .A1(n5261), .A2(n9451), .ZN(n5262) );
  MUX2_X1 U6719 ( .A(n9451), .B(n5262), .S(P1_IR_REG_6__SCAN_IN), .Z(n5264) );
  NAND2_X1 U6720 ( .A1(n5234), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n5266) );
  INV_X1 U6721 ( .A(n9742), .ZN(n6919) );
  XNOR2_X1 U6722 ( .A(n5268), .B(n5267), .ZN(n6328) );
  OR2_X1 U6723 ( .A1(n6328), .A2(n5241), .ZN(n5271) );
  NAND2_X1 U6724 ( .A1(n5263), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5269) );
  XNOR2_X1 U6725 ( .A(n5269), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6300) );
  AOI22_X1 U6726 ( .A1(n5234), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6270), .B2(
        n6300), .ZN(n5270) );
  NAND2_X1 U6727 ( .A1(n5271), .A2(n5270), .ZN(n6897) );
  XNOR2_X1 U6728 ( .A(n5273), .B(n5272), .ZN(n6331) );
  OR2_X1 U6729 ( .A1(n6331), .A2(n5241), .ZN(n5278) );
  NAND2_X1 U6730 ( .A1(n5274), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5276) );
  INV_X1 U6731 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5275) );
  XNOR2_X1 U6732 ( .A(n5276), .B(n5275), .ZN(n6560) );
  INV_X1 U6733 ( .A(n6560), .ZN(n6282) );
  AOI22_X1 U6734 ( .A1(n5234), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6270), .B2(
        n6282), .ZN(n5277) );
  NAND2_X1 U6735 ( .A1(n5278), .A2(n5277), .ZN(n9749) );
  XNOR2_X1 U6736 ( .A(n5280), .B(n5279), .ZN(n6333) );
  NAND2_X1 U6737 ( .A1(n6333), .A2(n7739), .ZN(n5284) );
  OR2_X1 U6738 ( .A1(n5281), .A2(n9451), .ZN(n5282) );
  XNOR2_X1 U6739 ( .A(n5282), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6508) );
  AOI22_X1 U6740 ( .A1(n5234), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6270), .B2(
        n6508), .ZN(n5283) );
  NAND2_X1 U6741 ( .A1(n5284), .A2(n5283), .ZN(n7205) );
  INV_X1 U6742 ( .A(n7205), .ZN(n9761) );
  XNOR2_X1 U6743 ( .A(n5286), .B(n5285), .ZN(n6340) );
  NAND2_X1 U6744 ( .A1(n6340), .A2(n7739), .ZN(n5292) );
  INV_X1 U6745 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5287) );
  NAND2_X1 U6746 ( .A1(n5281), .A2(n5287), .ZN(n5300) );
  NAND2_X1 U6747 ( .A1(n5300), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5289) );
  INV_X1 U6748 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5288) );
  NAND2_X1 U6749 ( .A1(n5289), .A2(n5288), .ZN(n5295) );
  OR2_X1 U6750 ( .A1(n5289), .A2(n5288), .ZN(n5290) );
  AOI22_X1 U6751 ( .A1(n5234), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6270), .B2(
        n6510), .ZN(n5291) );
  NAND2_X1 U6752 ( .A1(n5292), .A2(n5291), .ZN(n9510) );
  OR2_X1 U6753 ( .A1(n9511), .A2(n9510), .ZN(n9512) );
  XNOR2_X1 U6754 ( .A(n5294), .B(n5293), .ZN(n6338) );
  NAND2_X1 U6755 ( .A1(n6338), .A2(n7739), .ZN(n5298) );
  NAND2_X1 U6756 ( .A1(n5295), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5296) );
  XNOR2_X1 U6757 ( .A(n5296), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9103) );
  AOI22_X1 U6758 ( .A1(n5234), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6270), .B2(
        n9103), .ZN(n5297) );
  NAND2_X1 U6759 ( .A1(n6345), .A2(n7739), .ZN(n5307) );
  NAND2_X1 U6760 ( .A1(n5302), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5301) );
  MUX2_X1 U6761 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5301), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n5304) );
  INV_X1 U6762 ( .A(n5316), .ZN(n5303) );
  NAND2_X1 U6763 ( .A1(n5304), .A2(n5303), .ZN(n9119) );
  OAI22_X1 U6764 ( .A1(n5319), .A2(n10266), .B1(n9119), .B2(n5228), .ZN(n5305)
         );
  INV_X1 U6765 ( .A(n5305), .ZN(n5306) );
  INV_X1 U6766 ( .A(n7485), .ZN(n9549) );
  XNOR2_X1 U6767 ( .A(n5309), .B(n5308), .ZN(n6348) );
  NAND2_X1 U6768 ( .A1(n6348), .A2(n7739), .ZN(n5312) );
  OR2_X1 U6769 ( .A1(n5316), .A2(n9451), .ZN(n5310) );
  XNOR2_X1 U6770 ( .A(n5310), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9638) );
  AOI22_X1 U6771 ( .A1(n5234), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n9638), .B2(
        n6270), .ZN(n5311) );
  INV_X1 U6772 ( .A(n7537), .ZN(n9541) );
  NAND2_X1 U6773 ( .A1(n7533), .A2(n9541), .ZN(n7548) );
  XNOR2_X1 U6774 ( .A(n5314), .B(n5313), .ZN(n6356) );
  NAND2_X1 U6775 ( .A1(n6356), .A2(n7739), .ZN(n5322) );
  INV_X1 U6776 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5315) );
  OR2_X1 U6777 ( .A1(n5333), .A2(n9451), .ZN(n5318) );
  NAND2_X1 U6778 ( .A1(n5318), .A2(n5317), .ZN(n5325) );
  OAI21_X1 U6779 ( .B1(n5318), .B2(n5317), .A(n5325), .ZN(n9653) );
  OAI22_X1 U6780 ( .A1(n9653), .A2(n5228), .B1(n5319), .B2(n10102), .ZN(n5320)
         );
  INV_X1 U6781 ( .A(n5320), .ZN(n5321) );
  XNOR2_X1 U6782 ( .A(n5324), .B(n5323), .ZN(n6457) );
  NAND2_X1 U6783 ( .A1(n6457), .A2(n7739), .ZN(n5328) );
  NAND2_X1 U6784 ( .A1(n5325), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5326) );
  XNOR2_X1 U6785 ( .A(n5326), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9667) );
  AOI22_X1 U6786 ( .A1(n9667), .A2(n6270), .B1(n5234), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n5327) );
  XNOR2_X1 U6787 ( .A(n5331), .B(n5330), .ZN(n6543) );
  NAND2_X1 U6788 ( .A1(n6543), .A2(n7739), .ZN(n5336) );
  NOR2_X1 U6789 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5332) );
  NAND2_X1 U6790 ( .A1(n5333), .A2(n5332), .ZN(n5339) );
  NAND2_X1 U6791 ( .A1(n5339), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5334) );
  XNOR2_X1 U6792 ( .A(n5334), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9676) );
  AOI22_X1 U6793 ( .A1(n9676), .A2(n6270), .B1(n5234), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n5335) );
  XNOR2_X1 U6794 ( .A(n5338), .B(n5337), .ZN(n6601) );
  NAND2_X1 U6795 ( .A1(n6601), .A2(n7739), .ZN(n5344) );
  NAND2_X1 U6796 ( .A1(n5340), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5341) );
  OR2_X1 U6797 ( .A1(n5341), .A2(n10241), .ZN(n5342) );
  NAND2_X1 U6798 ( .A1(n5341), .A2(n10241), .ZN(n5347) );
  AOI22_X1 U6799 ( .A1(n9116), .A2(n6270), .B1(n5234), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n5343) );
  INV_X1 U6800 ( .A(n9420), .ZN(n9314) );
  XNOR2_X1 U6801 ( .A(n5346), .B(n5345), .ZN(n6839) );
  NAND2_X1 U6802 ( .A1(n6839), .A2(n7739), .ZN(n5350) );
  NAND2_X1 U6803 ( .A1(n5347), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5348) );
  XNOR2_X1 U6804 ( .A(n5348), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9708) );
  AOI22_X1 U6805 ( .A1(n9708), .A2(n6270), .B1(n5234), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n5349) );
  XNOR2_X1 U6806 ( .A(n5352), .B(n5351), .ZN(n6923) );
  NAND2_X1 U6807 ( .A1(n6923), .A2(n7739), .ZN(n5354) );
  AOI22_X1 U6808 ( .A1(n5234), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9257), .B2(
        n6270), .ZN(n5353) );
  XNOR2_X1 U6809 ( .A(n5356), .B(n5355), .ZN(n7085) );
  NAND2_X1 U6810 ( .A1(n7085), .A2(n7739), .ZN(n5358) );
  NAND2_X1 U6811 ( .A1(n5234), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5357) );
  NAND2_X1 U6812 ( .A1(n9280), .A2(n9269), .ZN(n9264) );
  XNOR2_X1 U6813 ( .A(n5360), .B(n5359), .ZN(n7089) );
  NAND2_X1 U6814 ( .A1(n7089), .A2(n7739), .ZN(n5362) );
  NAND2_X1 U6815 ( .A1(n5234), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5361) );
  XNOR2_X1 U6816 ( .A(n5364), .B(n5363), .ZN(n7470) );
  NAND2_X1 U6817 ( .A1(n7470), .A2(n7739), .ZN(n5366) );
  NAND2_X1 U6818 ( .A1(n5234), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5365) );
  INV_X1 U6819 ( .A(n5367), .ZN(n5369) );
  NAND2_X1 U6820 ( .A1(n5369), .A2(n5368), .ZN(n5371) );
  NAND2_X1 U6821 ( .A1(n5371), .A2(n5370), .ZN(n7472) );
  NAND2_X1 U6822 ( .A1(n7472), .A2(n7739), .ZN(n5373) );
  NAND2_X1 U6823 ( .A1(n5234), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5372) );
  NAND2_X1 U6824 ( .A1(n7556), .A2(n7739), .ZN(n5377) );
  NAND2_X1 U6825 ( .A1(n5234), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5376) );
  INV_X1 U6826 ( .A(n9387), .ZN(n9216) );
  XNOR2_X1 U6827 ( .A(n5379), .B(n5378), .ZN(n7572) );
  NAND2_X1 U6828 ( .A1(n7572), .A2(n7739), .ZN(n5381) );
  NAND2_X1 U6829 ( .A1(n5234), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5380) );
  NAND2_X1 U6830 ( .A1(n7590), .A2(n7739), .ZN(n5385) );
  NAND2_X1 U6831 ( .A1(n5234), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5384) );
  NOR2_X2 U6832 ( .A1(n5045), .A2(n9375), .ZN(n9176) );
  NAND2_X1 U6833 ( .A1(n9163), .A2(n9176), .ZN(n9158) );
  OR2_X2 U6834 ( .A1(n7763), .A2(n9158), .ZN(n7776) );
  INV_X1 U6835 ( .A(n7776), .ZN(n5386) );
  AOI211_X1 U6836 ( .C1(n7763), .C2(n9158), .A(n9762), .B(n5386), .ZN(n9148)
         );
  NOR2_X1 U6837 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5388) );
  NAND2_X1 U6838 ( .A1(n5391), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5392) );
  MUX2_X1 U6839 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5392), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5394) );
  INV_X1 U6840 ( .A(n5393), .ZN(n9452) );
  NAND2_X1 U6841 ( .A1(n5415), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5402) );
  NAND2_X1 U6842 ( .A1(n5422), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5401) );
  AND2_X4 U6843 ( .A1(n9458), .A2(n5397), .ZN(n5421) );
  NAND2_X1 U6844 ( .A1(n5421), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5400) );
  NAND2_X2 U6845 ( .A1(n5397), .A2(n5396), .ZN(n5419) );
  INV_X1 U6846 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5398) );
  NAND2_X1 U6847 ( .A1(n5421), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U6848 ( .A1(n5415), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5405) );
  INV_X1 U6849 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5403) );
  OR2_X1 U6850 ( .A1(n5419), .A2(n5403), .ZN(n5404) );
  INV_X1 U6851 ( .A(n9102), .ZN(n6609) );
  AND2_X1 U6852 ( .A1(n6609), .A2(n6597), .ZN(n6606) );
  NAND2_X1 U6853 ( .A1(n6607), .A2(n6606), .ZN(n6605) );
  NAND2_X1 U6854 ( .A1(n5644), .A2(n9042), .ZN(n5407) );
  NAND2_X1 U6855 ( .A1(n5415), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5411) );
  INV_X1 U6856 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5408) );
  NAND2_X1 U6857 ( .A1(n5421), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5409) );
  NAND3_X1 U6858 ( .A1(n5411), .A2(n5410), .A3(n5409), .ZN(n5412) );
  NAND2_X1 U6859 ( .A1(n9732), .A2(n9099), .ZN(n9044) );
  NAND2_X1 U6860 ( .A1(n9047), .A2(n9044), .ZN(n5646) );
  NAND2_X1 U6861 ( .A1(n9046), .A2(n8882), .ZN(n5413) );
  NAND2_X1 U6862 ( .A1(n5413), .A2(n9047), .ZN(n8860) );
  INV_X1 U6863 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5414) );
  NAND2_X1 U6864 ( .A1(n5422), .A2(n5414), .ZN(n5418) );
  NAND2_X1 U6865 ( .A1(n5415), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5417) );
  NAND2_X1 U6866 ( .A1(n5421), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5416) );
  INV_X2 U6867 ( .A(n5419), .ZN(n5431) );
  NAND2_X1 U6868 ( .A1(n5431), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5420) );
  INV_X1 U6869 ( .A(n6587), .ZN(n6539) );
  NAND2_X1 U6870 ( .A1(n6539), .A2(n9098), .ZN(n8853) );
  INV_X1 U6871 ( .A(n6526), .ZN(n8880) );
  NAND2_X1 U6872 ( .A1(n8860), .A2(n8880), .ZN(n6528) );
  NAND2_X1 U6873 ( .A1(n6528), .A2(n9048), .ZN(n6738) );
  NAND2_X1 U6874 ( .A1(n7770), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5427) );
  NAND2_X1 U6875 ( .A1(n5421), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5426) );
  INV_X1 U6876 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5423) );
  XNOR2_X1 U6877 ( .A(n5423), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n6748) );
  NAND2_X1 U6878 ( .A1(n5422), .A2(n6748), .ZN(n5425) );
  NAND2_X1 U6879 ( .A1(n5431), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5424) );
  NAND2_X1 U6880 ( .A1(n6732), .A2(n6747), .ZN(n9052) );
  INV_X1 U6881 ( .A(n9052), .ZN(n5428) );
  INV_X1 U6882 ( .A(n6747), .ZN(n9736) );
  NAND2_X1 U6883 ( .A1(n9736), .A2(n9097), .ZN(n8854) );
  NAND2_X1 U6884 ( .A1(n7770), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U6885 ( .A1(n5421), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5434) );
  NAND3_X1 U6886 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5439) );
  INV_X1 U6887 ( .A(n5439), .ZN(n5429) );
  NAND2_X1 U6888 ( .A1(n5429), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5448) );
  INV_X1 U6889 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6464) );
  NAND2_X1 U6890 ( .A1(n5439), .A2(n6464), .ZN(n5430) );
  AND2_X1 U6891 ( .A1(n5448), .A2(n5430), .ZN(n6774) );
  NAND2_X1 U6892 ( .A1(n5422), .A2(n6774), .ZN(n5433) );
  NAND2_X1 U6893 ( .A1(n5431), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5432) );
  NAND4_X1 U6894 ( .A1(n5435), .A2(n5434), .A3(n5433), .A4(n5432), .ZN(n9095)
         );
  INV_X1 U6895 ( .A(n9095), .ZN(n6850) );
  NAND2_X1 U6896 ( .A1(n6850), .A2(n9742), .ZN(n8942) );
  NAND2_X1 U6897 ( .A1(n7770), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5443) );
  NAND2_X1 U6898 ( .A1(n5421), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5442) );
  INV_X1 U6899 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5437) );
  NAND2_X1 U6900 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5436) );
  NAND2_X1 U6901 ( .A1(n5437), .A2(n5436), .ZN(n5438) );
  AND2_X1 U6902 ( .A1(n5439), .A2(n5438), .ZN(n6759) );
  NAND2_X1 U6903 ( .A1(n5422), .A2(n6759), .ZN(n5441) );
  NAND2_X1 U6904 ( .A1(n5431), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5440) );
  NAND4_X1 U6905 ( .A1(n5443), .A2(n5442), .A3(n5441), .A4(n5440), .ZN(n9096)
         );
  INV_X1 U6906 ( .A(n9096), .ZN(n6907) );
  NAND2_X1 U6907 ( .A1(n6907), .A2(n6879), .ZN(n8936) );
  AND2_X1 U6908 ( .A1(n8942), .A2(n8936), .ZN(n9053) );
  NAND2_X1 U6909 ( .A1(n8937), .A2(n9053), .ZN(n5445) );
  NAND2_X1 U6910 ( .A1(n6919), .A2(n9095), .ZN(n8933) );
  INV_X1 U6911 ( .A(n6879), .ZN(n6761) );
  NAND2_X1 U6912 ( .A1(n6761), .A2(n9096), .ZN(n8938) );
  NAND2_X1 U6913 ( .A1(n8933), .A2(n8938), .ZN(n5444) );
  NAND2_X1 U6914 ( .A1(n5444), .A2(n8942), .ZN(n9055) );
  NAND2_X1 U6915 ( .A1(n5445), .A2(n9055), .ZN(n6848) );
  NAND2_X1 U6916 ( .A1(n5421), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5453) );
  NAND2_X1 U6917 ( .A1(n7770), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5452) );
  INV_X1 U6918 ( .A(n5448), .ZN(n5446) );
  NAND2_X1 U6919 ( .A1(n5446), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5455) );
  INV_X1 U6920 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U6921 ( .A1(n5448), .A2(n5447), .ZN(n5449) );
  AND2_X1 U6922 ( .A1(n5455), .A2(n5449), .ZN(n6845) );
  NAND2_X1 U6923 ( .A1(n5422), .A2(n6845), .ZN(n5451) );
  NAND2_X1 U6924 ( .A1(n5431), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5450) );
  NAND4_X1 U6925 ( .A1(n5453), .A2(n5452), .A3(n5451), .A4(n5450), .ZN(n9094)
         );
  INV_X1 U6926 ( .A(n9094), .ZN(n7213) );
  OR2_X1 U6927 ( .A1(n7213), .A2(n6897), .ZN(n8944) );
  NAND2_X1 U6928 ( .A1(n6897), .A2(n7213), .ZN(n8941) );
  NAND2_X1 U6929 ( .A1(n8944), .A2(n8941), .ZN(n8887) );
  NAND2_X1 U6930 ( .A1(n5421), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U6931 ( .A1(n7770), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5459) );
  INV_X1 U6932 ( .A(n5455), .ZN(n5454) );
  NAND2_X1 U6933 ( .A1(n5454), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5462) );
  INV_X1 U6934 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6557) );
  NAND2_X1 U6935 ( .A1(n5455), .A2(n6557), .ZN(n5456) );
  AND2_X1 U6936 ( .A1(n5462), .A2(n5456), .ZN(n7222) );
  NAND2_X1 U6937 ( .A1(n5422), .A2(n7222), .ZN(n5458) );
  NAND2_X1 U6938 ( .A1(n5431), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5457) );
  NAND4_X1 U6939 ( .A1(n5460), .A2(n5459), .A3(n5458), .A4(n5457), .ZN(n9093)
         );
  NAND2_X1 U6940 ( .A1(n9749), .A2(n7198), .ZN(n8955) );
  AND2_X1 U6941 ( .A1(n8955), .A2(n8941), .ZN(n8934) );
  NAND2_X1 U6942 ( .A1(n5462), .A2(n5461), .ZN(n5463) );
  AND2_X1 U6943 ( .A1(n5470), .A2(n5463), .ZN(n7204) );
  NAND2_X1 U6944 ( .A1(n5422), .A2(n7204), .ZN(n5467) );
  NAND2_X1 U6945 ( .A1(n7770), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5466) );
  NAND2_X1 U6946 ( .A1(n5431), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5465) );
  NAND2_X1 U6947 ( .A1(n5421), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5464) );
  NAND4_X1 U6948 ( .A1(n5467), .A2(n5466), .A3(n5465), .A4(n5464), .ZN(n9092)
         );
  INV_X1 U6949 ( .A(n9092), .ZN(n9503) );
  OR2_X1 U6950 ( .A1(n7205), .A2(n9503), .ZN(n7193) );
  OR2_X1 U6951 ( .A1(n9749), .A2(n7198), .ZN(n7195) );
  AND2_X1 U6952 ( .A1(n7193), .A2(n7195), .ZN(n8948) );
  NAND2_X1 U6953 ( .A1(n7770), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U6954 ( .A1(n5421), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U6955 ( .A1(n5470), .A2(n5469), .ZN(n5471) );
  AND2_X1 U6956 ( .A1(n5478), .A2(n5471), .ZN(n9507) );
  NAND2_X1 U6957 ( .A1(n5422), .A2(n9507), .ZN(n5473) );
  NAND2_X1 U6958 ( .A1(n5431), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5472) );
  NAND4_X1 U6959 ( .A1(n5475), .A2(n5474), .A3(n5473), .A4(n5472), .ZN(n9091)
         );
  NAND2_X1 U6960 ( .A1(n9510), .A2(n7356), .ZN(n8951) );
  NAND2_X1 U6961 ( .A1(n7205), .A2(n9503), .ZN(n9494) );
  AND2_X1 U6962 ( .A1(n8951), .A2(n9494), .ZN(n8949) );
  NAND2_X1 U6963 ( .A1(n9491), .A2(n9498), .ZN(n7355) );
  NAND2_X1 U6964 ( .A1(n7770), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5483) );
  NAND2_X1 U6965 ( .A1(n5421), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5482) );
  INV_X1 U6966 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U6967 ( .A1(n5478), .A2(n5477), .ZN(n5479) );
  AND2_X1 U6968 ( .A1(n5486), .A2(n5479), .ZN(n7362) );
  NAND2_X1 U6969 ( .A1(n5422), .A2(n7362), .ZN(n5481) );
  NAND2_X1 U6970 ( .A1(n5431), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5480) );
  NAND4_X1 U6971 ( .A1(n5483), .A2(n5482), .A3(n5481), .A4(n5480), .ZN(n9090)
         );
  NAND2_X1 U6972 ( .A1(n9555), .A2(n9500), .ZN(n8962) );
  NAND2_X1 U6973 ( .A1(n7355), .A2(n8962), .ZN(n5484) );
  OR2_X1 U6974 ( .A1(n9555), .A2(n9500), .ZN(n8843) );
  NAND2_X1 U6975 ( .A1(n5484), .A2(n8843), .ZN(n7477) );
  NAND2_X1 U6976 ( .A1(n7770), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5491) );
  NAND2_X1 U6977 ( .A1(n5421), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5490) );
  INV_X1 U6978 ( .A(n5486), .ZN(n5485) );
  NAND2_X1 U6979 ( .A1(n5485), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5495) );
  INV_X1 U6980 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7464) );
  NAND2_X1 U6981 ( .A1(n5486), .A2(n7464), .ZN(n5487) );
  AND2_X1 U6982 ( .A1(n5495), .A2(n5487), .ZN(n7484) );
  NAND2_X1 U6983 ( .A1(n5422), .A2(n7484), .ZN(n5489) );
  NAND2_X1 U6984 ( .A1(n5431), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5488) );
  NAND4_X1 U6985 ( .A1(n5491), .A2(n5490), .A3(n5489), .A4(n5488), .ZN(n9089)
         );
  INV_X1 U6986 ( .A(n8964), .ZN(n5492) );
  NAND2_X1 U6987 ( .A1(n7485), .A2(n7528), .ZN(n8963) );
  NAND2_X1 U6988 ( .A1(n5493), .A2(n8963), .ZN(n7527) );
  NAND2_X1 U6989 ( .A1(n5421), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U6990 ( .A1(n7770), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5499) );
  NAND2_X1 U6991 ( .A1(n5495), .A2(n5494), .ZN(n5496) );
  AND2_X1 U6992 ( .A1(n5502), .A2(n5496), .ZN(n7506) );
  NAND2_X1 U6993 ( .A1(n5422), .A2(n7506), .ZN(n5498) );
  NAND2_X1 U6994 ( .A1(n5431), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5497) );
  NAND4_X1 U6995 ( .A1(n5500), .A2(n5499), .A3(n5498), .A4(n5497), .ZN(n9088)
         );
  OR2_X1 U6996 ( .A1(n7537), .A2(n7542), .ZN(n8842) );
  NAND2_X1 U6997 ( .A1(n7537), .A2(n7542), .ZN(n8836) );
  NAND2_X1 U6998 ( .A1(n7770), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U6999 ( .A1(n5431), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5506) );
  INV_X1 U7000 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8675) );
  NAND2_X1 U7001 ( .A1(n5502), .A2(n8675), .ZN(n5503) );
  AND2_X1 U7002 ( .A1(n5509), .A2(n5503), .ZN(n8676) );
  NAND2_X1 U7003 ( .A1(n5422), .A2(n8676), .ZN(n5505) );
  NAND2_X1 U7004 ( .A1(n5421), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5504) );
  NAND4_X1 U7005 ( .A1(n5507), .A2(n5506), .A3(n5505), .A4(n5504), .ZN(n9087)
         );
  XNOR2_X1 U7006 ( .A(n8835), .B(n9344), .ZN(n7545) );
  OR2_X1 U7007 ( .A1(n8835), .A2(n9344), .ZN(n8846) );
  NAND2_X1 U7008 ( .A1(n7770), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5514) );
  NAND2_X1 U7009 ( .A1(n5421), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5513) );
  NAND2_X1 U7010 ( .A1(n5509), .A2(n5508), .ZN(n5510) );
  AND2_X1 U7011 ( .A1(n5517), .A2(n5510), .ZN(n9355) );
  NAND2_X1 U7012 ( .A1(n5422), .A2(n9355), .ZN(n5512) );
  NAND2_X1 U7013 ( .A1(n5431), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5511) );
  NAND4_X1 U7014 ( .A1(n5514), .A2(n5513), .A3(n5512), .A4(n5511), .ZN(n9086)
         );
  NAND2_X1 U7015 ( .A1(n9430), .A2(n9330), .ZN(n8979) );
  NAND2_X1 U7016 ( .A1(n9342), .A2(n8979), .ZN(n5515) );
  OR2_X1 U7017 ( .A1(n9430), .A2(n9330), .ZN(n8978) );
  NAND2_X1 U7018 ( .A1(n5515), .A2(n8978), .ZN(n9328) );
  INV_X1 U7019 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8721) );
  NAND2_X1 U7020 ( .A1(n5517), .A2(n8721), .ZN(n5518) );
  AND2_X1 U7021 ( .A1(n5532), .A2(n5518), .ZN(n9333) );
  NAND2_X1 U7022 ( .A1(n9333), .A2(n5422), .ZN(n5522) );
  NAND2_X1 U7023 ( .A1(n5421), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U7024 ( .A1(n7770), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U7025 ( .A1(n5431), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5519) );
  NAND4_X1 U7026 ( .A1(n5522), .A2(n5521), .A3(n5520), .A4(n5519), .ZN(n9318)
         );
  INV_X1 U7027 ( .A(n9318), .ZN(n9343) );
  OR2_X1 U7028 ( .A1(n9427), .A2(n9343), .ZN(n8983) );
  INV_X1 U7029 ( .A(n8983), .ZN(n5523) );
  NAND2_X1 U7030 ( .A1(n9427), .A2(n9343), .ZN(n8982) );
  INV_X1 U7031 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n5530) );
  INV_X1 U7032 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U7033 ( .A1(n5534), .A2(n5526), .ZN(n5527) );
  NAND2_X1 U7034 ( .A1(n5540), .A2(n5527), .ZN(n9295) );
  OR2_X1 U7035 ( .A1(n9295), .A2(n5636), .ZN(n5529) );
  AOI22_X1 U7036 ( .A1(n5421), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n7770), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n5528) );
  OAI211_X1 U7037 ( .C1(n5419), .C2(n5530), .A(n5529), .B(n5528), .ZN(n10326)
         );
  INV_X1 U7038 ( .A(n10326), .ZN(n7637) );
  NAND2_X1 U7039 ( .A1(n9417), .A2(n7637), .ZN(n8824) );
  NAND2_X1 U7040 ( .A1(n5532), .A2(n5531), .ZN(n5533) );
  NAND2_X1 U7041 ( .A1(n5534), .A2(n5533), .ZN(n9310) );
  NAND2_X1 U7042 ( .A1(n7770), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5536) );
  NAND2_X1 U7043 ( .A1(n5421), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5535) );
  AND2_X1 U7044 ( .A1(n5536), .A2(n5535), .ZN(n5538) );
  NAND2_X1 U7045 ( .A1(n5431), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5537) );
  OAI211_X1 U7046 ( .C1(n9310), .C2(n5636), .A(n5538), .B(n5537), .ZN(n9085)
         );
  INV_X1 U7047 ( .A(n9085), .ZN(n9331) );
  NAND2_X1 U7048 ( .A1(n9420), .A2(n9331), .ZN(n9298) );
  NAND2_X1 U7049 ( .A1(n8824), .A2(n9298), .ZN(n8930) );
  OR2_X1 U7050 ( .A1(n9417), .A2(n7637), .ZN(n8988) );
  OR2_X1 U7051 ( .A1(n9420), .A2(n9331), .ZN(n9299) );
  AND2_X1 U7052 ( .A1(n8988), .A2(n9299), .ZN(n8931) );
  INV_X1 U7053 ( .A(n8824), .ZN(n5539) );
  NAND2_X1 U7054 ( .A1(n5540), .A2(n8699), .ZN(n5541) );
  AND2_X1 U7055 ( .A1(n5550), .A2(n5541), .ZN(n9281) );
  NAND2_X1 U7056 ( .A1(n9281), .A2(n5422), .ZN(n5547) );
  INV_X1 U7057 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U7058 ( .A1(n5421), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5543) );
  NAND2_X1 U7059 ( .A1(n5431), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5542) );
  OAI211_X1 U7060 ( .C1(n5468), .C2(n5544), .A(n5543), .B(n5542), .ZN(n5545)
         );
  INV_X1 U7061 ( .A(n5545), .ZN(n5546) );
  NAND2_X1 U7062 ( .A1(n5547), .A2(n5546), .ZN(n9274) );
  INV_X1 U7063 ( .A(n9274), .ZN(n9304) );
  OR2_X1 U7064 ( .A1(n9410), .A2(n9304), .ZN(n8989) );
  NAND2_X1 U7065 ( .A1(n9410), .A2(n9304), .ZN(n9270) );
  NAND2_X1 U7066 ( .A1(n8989), .A2(n9270), .ZN(n9284) );
  INV_X1 U7067 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5549) );
  NAND2_X1 U7068 ( .A1(n5550), .A2(n5549), .ZN(n5551) );
  NAND2_X1 U7069 ( .A1(n5565), .A2(n5551), .ZN(n8745) );
  OR2_X1 U7070 ( .A1(n8745), .A2(n5636), .ZN(n5556) );
  INV_X1 U7071 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10209) );
  NAND2_X1 U7072 ( .A1(n5421), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5553) );
  NAND2_X1 U7073 ( .A1(n7770), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5552) );
  OAI211_X1 U7074 ( .C1(n10209), .C2(n5419), .A(n5553), .B(n5552), .ZN(n5554)
         );
  INV_X1 U7075 ( .A(n5554), .ZN(n5555) );
  NAND2_X1 U7076 ( .A1(n5556), .A2(n5555), .ZN(n9286) );
  NAND2_X1 U7077 ( .A1(n9405), .A2(n9251), .ZN(n8827) );
  AND2_X1 U7078 ( .A1(n8827), .A2(n9270), .ZN(n8990) );
  NOR2_X1 U7079 ( .A1(n9405), .A2(n9251), .ZN(n8998) );
  XNOR2_X1 U7080 ( .A(n5565), .B(P1_REG3_REG_21__SCAN_IN), .ZN(n9255) );
  NAND2_X1 U7081 ( .A1(n9255), .A2(n5422), .ZN(n5561) );
  INV_X1 U7082 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10122) );
  NAND2_X1 U7083 ( .A1(n7770), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5558) );
  NAND2_X1 U7084 ( .A1(n5421), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5557) );
  OAI211_X1 U7085 ( .C1(n10122), .C2(n5419), .A(n5558), .B(n5557), .ZN(n5559)
         );
  INV_X1 U7086 ( .A(n5559), .ZN(n5560) );
  NAND2_X1 U7087 ( .A1(n5561), .A2(n5560), .ZN(n9273) );
  OR2_X1 U7088 ( .A1(n9402), .A2(n8758), .ZN(n8828) );
  NAND2_X1 U7089 ( .A1(n9402), .A2(n8758), .ZN(n8992) );
  NAND2_X1 U7090 ( .A1(n8828), .A2(n8992), .ZN(n9248) );
  INV_X1 U7091 ( .A(n9248), .ZN(n8901) );
  NAND2_X1 U7092 ( .A1(n9249), .A2(n8901), .ZN(n5562) );
  NAND2_X1 U7093 ( .A1(n5562), .A2(n8992), .ZN(n9240) );
  INV_X1 U7094 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5563) );
  INV_X1 U7095 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5564) );
  OAI21_X1 U7096 ( .B1(n5565), .B2(n5563), .A(n5564), .ZN(n5566) );
  AND2_X1 U7097 ( .A1(n5566), .A2(n5574), .ZN(n9238) );
  NAND2_X1 U7098 ( .A1(n9238), .A2(n5422), .ZN(n5571) );
  INV_X1 U7099 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n10134) );
  NAND2_X1 U7100 ( .A1(n5421), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U7101 ( .A1(n7770), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5567) );
  OAI211_X1 U7102 ( .C1(n10134), .C2(n5419), .A(n5568), .B(n5567), .ZN(n5569)
         );
  INV_X1 U7103 ( .A(n5569), .ZN(n5570) );
  NAND2_X1 U7104 ( .A1(n5571), .A2(n5570), .ZN(n9229) );
  INV_X1 U7105 ( .A(n9229), .ZN(n9252) );
  OR2_X1 U7106 ( .A1(n9395), .A2(n9252), .ZN(n8831) );
  NAND2_X1 U7107 ( .A1(n9395), .A2(n9252), .ZN(n8993) );
  NAND2_X1 U7108 ( .A1(n9240), .A2(n9241), .ZN(n5572) );
  NAND2_X1 U7109 ( .A1(n5572), .A2(n8993), .ZN(n9226) );
  INV_X1 U7110 ( .A(n5574), .ZN(n5573) );
  NAND2_X1 U7111 ( .A1(n5573), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5584) );
  INV_X1 U7112 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n10116) );
  NAND2_X1 U7113 ( .A1(n5574), .A2(n10116), .ZN(n5575) );
  AND2_X1 U7114 ( .A1(n5584), .A2(n5575), .ZN(n9223) );
  NAND2_X1 U7115 ( .A1(n9223), .A2(n5422), .ZN(n5581) );
  INV_X1 U7116 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U7117 ( .A1(n7770), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5577) );
  NAND2_X1 U7118 ( .A1(n5431), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5576) );
  OAI211_X1 U7119 ( .C1(n5578), .C2(n5627), .A(n5577), .B(n5576), .ZN(n5579)
         );
  INV_X1 U7120 ( .A(n5579), .ZN(n5580) );
  NAND2_X1 U7121 ( .A1(n9390), .A2(n9209), .ZN(n9001) );
  NAND2_X1 U7122 ( .A1(n8926), .A2(n9001), .ZN(n9219) );
  INV_X1 U7123 ( .A(n5584), .ZN(n5582) );
  INV_X1 U7124 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U7125 ( .A1(n5584), .A2(n5583), .ZN(n5585) );
  NAND2_X1 U7126 ( .A1(n5593), .A2(n5585), .ZN(n9212) );
  INV_X1 U7127 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7128 ( .A1(n7770), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U7129 ( .A1(n5431), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5586) );
  OAI211_X1 U7130 ( .C1(n5627), .C2(n5588), .A(n5587), .B(n5586), .ZN(n5589)
         );
  INV_X1 U7131 ( .A(n5589), .ZN(n5590) );
  XNOR2_X1 U7132 ( .A(n9387), .B(n9196), .ZN(n9206) );
  NAND2_X1 U7133 ( .A1(n9387), .A2(n9196), .ZN(n8925) );
  INV_X1 U7134 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U7135 ( .A1(n5593), .A2(n5592), .ZN(n5594) );
  NAND2_X1 U7136 ( .A1(n9197), .A2(n5422), .ZN(n5600) );
  INV_X1 U7137 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U7138 ( .A1(n5421), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5596) );
  NAND2_X1 U7139 ( .A1(n7770), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5595) );
  OAI211_X1 U7140 ( .C1(n5597), .C2(n5419), .A(n5596), .B(n5595), .ZN(n5598)
         );
  INV_X1 U7141 ( .A(n5598), .ZN(n5599) );
  NAND2_X1 U7142 ( .A1(n9382), .A2(n9208), .ZN(n9012) );
  NAND2_X1 U7143 ( .A1(n9192), .A2(n9012), .ZN(n9182) );
  INV_X1 U7144 ( .A(n5603), .ZN(n5601) );
  NAND2_X1 U7145 ( .A1(n5601), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5613) );
  INV_X1 U7146 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5602) );
  NAND2_X1 U7147 ( .A1(n5603), .A2(n5602), .ZN(n5604) );
  NAND2_X1 U7148 ( .A1(n5613), .A2(n5604), .ZN(n9177) );
  INV_X1 U7149 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n5607) );
  NAND2_X1 U7150 ( .A1(n7770), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U7151 ( .A1(n5431), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5605) );
  OAI211_X1 U7152 ( .C1(n5627), .C2(n5607), .A(n5606), .B(n5605), .ZN(n5608)
         );
  INV_X1 U7153 ( .A(n5608), .ZN(n5609) );
  INV_X1 U7154 ( .A(n9164), .ZN(n9195) );
  OR2_X1 U7155 ( .A1(n9375), .A2(n9195), .ZN(n8923) );
  AND2_X1 U7156 ( .A1(n8923), .A2(n9181), .ZN(n9017) );
  NAND2_X1 U7157 ( .A1(n9182), .A2(n9017), .ZN(n5611) );
  NAND2_X1 U7158 ( .A1(n9375), .A2(n9195), .ZN(n9014) );
  INV_X1 U7159 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5612) );
  NAND2_X1 U7160 ( .A1(n5613), .A2(n5612), .ZN(n5614) );
  NAND2_X1 U7161 ( .A1(n9161), .A2(n5422), .ZN(n5619) );
  INV_X1 U7162 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10228) );
  NAND2_X1 U7163 ( .A1(n7770), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5616) );
  NAND2_X1 U7164 ( .A1(n5431), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5615) );
  OAI211_X1 U7165 ( .C1(n5627), .C2(n10228), .A(n5616), .B(n5615), .ZN(n5617)
         );
  INV_X1 U7166 ( .A(n5617), .ZN(n5618) );
  NAND2_X1 U7167 ( .A1(n9370), .A2(n7705), .ZN(n8922) );
  NAND2_X1 U7168 ( .A1(n9018), .A2(n8922), .ZN(n9168) );
  NAND2_X1 U7169 ( .A1(n9165), .A2(n9018), .ZN(n5631) );
  INV_X1 U7170 ( .A(n5622), .ZN(n5620) );
  NAND2_X1 U7171 ( .A1(n5620), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n7779) );
  INV_X1 U7172 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5621) );
  NAND2_X1 U7173 ( .A1(n5622), .A2(n5621), .ZN(n5623) );
  NAND2_X1 U7174 ( .A1(n7779), .A2(n5623), .ZN(n7702) );
  INV_X1 U7175 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U7176 ( .A1(n7770), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U7177 ( .A1(n5431), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5624) );
  OAI211_X1 U7178 ( .C1(n5627), .C2(n5626), .A(n5625), .B(n5624), .ZN(n5628)
         );
  INV_X1 U7179 ( .A(n5628), .ZN(n5629) );
  NAND2_X1 U7180 ( .A1(n7763), .A2(n7764), .ZN(n8810) );
  NAND2_X1 U7181 ( .A1(n9020), .A2(n8810), .ZN(n5667) );
  OR2_X1 U7182 ( .A1(n5672), .A2(n9135), .ZN(n5634) );
  OR2_X1 U7183 ( .A1(n5062), .A2(n5670), .ZN(n5633) );
  OR2_X1 U7184 ( .A1(n7779), .A2(n5636), .ZN(n5641) );
  INV_X1 U7185 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n7778) );
  NAND2_X1 U7186 ( .A1(n5421), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U7187 ( .A1(n5431), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5637) );
  OAI211_X1 U7188 ( .C1(n5468), .C2(n7778), .A(n5638), .B(n5637), .ZN(n5639)
         );
  INV_X1 U7189 ( .A(n5639), .ZN(n5640) );
  NAND2_X1 U7190 ( .A1(n5641), .A2(n5640), .ZN(n9084) );
  INV_X1 U7191 ( .A(n9084), .ZN(n7766) );
  INV_X1 U7192 ( .A(n5635), .ZN(n9572) );
  INV_X1 U7193 ( .A(n8835), .ZN(n9537) );
  NAND2_X1 U7194 ( .A1(n9042), .A2(n9101), .ZN(n5645) );
  AND2_X1 U7195 ( .A1(n6603), .A2(n5645), .ZN(n6694) );
  NAND2_X1 U7196 ( .A1(n9732), .A2(n6608), .ZN(n5647) );
  NAND2_X1 U7197 ( .A1(n6693), .A2(n5647), .ZN(n6519) );
  NAND2_X1 U7198 ( .A1(n6519), .A2(n6526), .ZN(n6518) );
  NAND2_X1 U7199 ( .A1(n6539), .A2(n6741), .ZN(n5648) );
  NAND2_X1 U7200 ( .A1(n6518), .A2(n5648), .ZN(n6740) );
  NAND2_X1 U7201 ( .A1(n8854), .A2(n9052), .ZN(n8879) );
  NAND2_X1 U7202 ( .A1(n6740), .A2(n8879), .ZN(n6739) );
  NAND2_X1 U7203 ( .A1(n9736), .A2(n6732), .ZN(n5649) );
  AND2_X1 U7204 ( .A1(n8938), .A2(n8936), .ZN(n5650) );
  INV_X1 U7205 ( .A(n5650), .ZN(n8885) );
  NAND2_X1 U7206 ( .A1(n6879), .A2(n9096), .ZN(n5651) );
  NAND2_X1 U7207 ( .A1(n6919), .A2(n6850), .ZN(n5653) );
  OR2_X1 U7208 ( .A1(n6897), .A2(n9094), .ZN(n5654) );
  NAND2_X1 U7209 ( .A1(n7195), .A2(n8955), .ZN(n7215) );
  AND2_X1 U7210 ( .A1(n7205), .A2(n9092), .ZN(n5655) );
  OAI22_X1 U7211 ( .A1(n7194), .A2(n5655), .B1(n9092), .B2(n7205), .ZN(n9490)
         );
  NAND2_X1 U7212 ( .A1(n9498), .A2(n8951), .ZN(n9492) );
  NAND2_X1 U7213 ( .A1(n9490), .A2(n9492), .ZN(n5657) );
  OR2_X1 U7214 ( .A1(n9510), .A2(n9091), .ZN(n5656) );
  NAND2_X1 U7215 ( .A1(n5657), .A2(n5656), .ZN(n7354) );
  NOR2_X1 U7216 ( .A1(n9555), .A2(n9090), .ZN(n5659) );
  NAND2_X1 U7217 ( .A1(n9555), .A2(n9090), .ZN(n5658) );
  NAND2_X1 U7218 ( .A1(n8964), .A2(n8963), .ZN(n8893) );
  NOR2_X1 U7219 ( .A1(n9420), .A2(n9085), .ZN(n5661) );
  NAND2_X1 U7220 ( .A1(n8988), .A2(n8824), .ZN(n9302) );
  INV_X1 U7221 ( .A(n9410), .ZN(n9283) );
  NAND2_X1 U7222 ( .A1(n5662), .A2(n5040), .ZN(n9247) );
  NAND2_X1 U7223 ( .A1(n9225), .A2(n9209), .ZN(n5663) );
  NAND2_X1 U7224 ( .A1(n9216), .A2(n9196), .ZN(n5664) );
  NAND2_X1 U7225 ( .A1(n5665), .A2(n5664), .ZN(n9191) );
  NAND2_X1 U7226 ( .A1(n9181), .A2(n9012), .ZN(n9193) );
  INV_X1 U7227 ( .A(n9382), .ZN(n9200) );
  OAI21_X1 U7228 ( .B1(n5668), .B2(n5667), .A(n7765), .ZN(n9156) );
  INV_X1 U7229 ( .A(n5669), .ZN(n5671) );
  INV_X1 U7230 ( .A(n6358), .ZN(n6524) );
  OR2_X1 U7231 ( .A1(n6524), .A2(n6390), .ZN(n5674) );
  OR2_X1 U7232 ( .A1(n6359), .A2(n5062), .ZN(n5673) );
  XNOR2_X1 U7233 ( .A(n5678), .B(P1_IR_REG_25__SCAN_IN), .ZN(n7573) );
  NAND2_X1 U7234 ( .A1(n5680), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5681) );
  INV_X1 U7235 ( .A(n5696), .ZN(n7557) );
  NAND2_X1 U7236 ( .A1(n7557), .A2(P1_B_REG_SCAN_IN), .ZN(n5686) );
  INV_X1 U7237 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5682) );
  NAND2_X1 U7238 ( .A1(n5678), .A2(n5682), .ZN(n5683) );
  NAND2_X1 U7239 ( .A1(n5683), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5684) );
  INV_X1 U7240 ( .A(P1_B_REG_SCAN_IN), .ZN(n7742) );
  NAND2_X1 U7241 ( .A1(n5696), .A2(n7742), .ZN(n5685) );
  OR2_X1 U7242 ( .A1(n9717), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5688) );
  OR2_X1 U7243 ( .A1(n7591), .A2(n7573), .ZN(n5687) );
  INV_X1 U7244 ( .A(n6520), .ZN(n5689) );
  OAI21_X1 U7245 ( .B1(n9756), .B2(n5671), .A(n5689), .ZN(n5695) );
  NAND2_X1 U7246 ( .A1(n5690), .A2(n10082), .ZN(n5691) );
  OAI21_X1 U7247 ( .B1(n5064), .B2(n5691), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5693) );
  NAND2_X1 U7248 ( .A1(n6522), .A2(n9722), .ZN(n6369) );
  OR2_X1 U7249 ( .A1(n9717), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5698) );
  OR2_X1 U7250 ( .A1(n7591), .A2(n5696), .ZN(n5697) );
  AND2_X1 U7251 ( .A1(n5698), .A2(n5697), .ZN(n9450) );
  INV_X1 U7252 ( .A(n9450), .ZN(n5710) );
  NOR2_X1 U7253 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .ZN(
        n5702) );
  NOR4_X1 U7254 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5701) );
  NOR4_X1 U7255 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n5700) );
  NOR4_X1 U7256 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n5699) );
  NAND4_X1 U7257 ( .A1(n5702), .A2(n5701), .A3(n5700), .A4(n5699), .ZN(n5708)
         );
  NOR4_X1 U7258 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5706) );
  NOR4_X1 U7259 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5705) );
  NOR4_X1 U7260 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5704) );
  NOR4_X1 U7261 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5703) );
  NAND4_X1 U7262 ( .A1(n5706), .A2(n5705), .A3(n5704), .A4(n5703), .ZN(n5707)
         );
  NOR2_X1 U7263 ( .A1(n5708), .A2(n5707), .ZN(n5709) );
  OR2_X1 U7264 ( .A1(n9717), .A2(n5709), .ZN(n6367) );
  NAND2_X1 U7265 ( .A1(n5710), .A2(n6367), .ZN(n6521) );
  NAND2_X1 U7266 ( .A1(n9369), .A2(n9759), .ZN(n5712) );
  NAND2_X1 U7267 ( .A1(n9768), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5711) );
  NOR2_X1 U7268 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5720) );
  NOR2_X1 U7269 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5719) );
  NOR2_X1 U7270 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5718) );
  INV_X1 U7271 ( .A(n5727), .ZN(n5725) );
  NAND2_X1 U7272 ( .A1(n5786), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5731) );
  NAND2_X1 U7273 ( .A1(n5785), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5730) );
  NAND2_X1 U7274 ( .A1(n4463), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5729) );
  NAND2_X1 U7275 ( .A1(n4462), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5728) );
  NAND4_X1 U7276 ( .A1(n10206), .A2(n5733), .A3(n5980), .A4(n5732), .ZN(n5734)
         );
  NAND2_X1 U7277 ( .A1(n6026), .A2(n5735), .ZN(n5741) );
  NAND2_X1 U7278 ( .A1(n5741), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U7279 ( .A1(n5740), .A2(n5739), .ZN(n5736) );
  NAND2_X1 U7280 ( .A1(n5736), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5738) );
  INV_X1 U7281 ( .A(n8159), .ZN(n6243) );
  INV_X1 U7282 ( .A(n5741), .ZN(n5744) );
  INV_X1 U7283 ( .A(n5748), .ZN(n7967) );
  NAND2_X2 U7284 ( .A1(n6243), .A2(n6231), .ZN(n7966) );
  NOR2_X1 U7285 ( .A1(n6807), .A2(n5791), .ZN(n5761) );
  INV_X1 U7286 ( .A(n5761), .ZN(n5759) );
  NAND2_X1 U7287 ( .A1(n6236), .A2(n5748), .ZN(n7265) );
  MUX2_X2 U7288 ( .A(n5750), .B(P2_IR_REG_31__SCAN_IN), .S(n10077), .Z(n5751)
         );
  INV_X1 U7289 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10091) );
  INV_X1 U7290 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9791) );
  NAND2_X1 U7291 ( .A1(n5809), .A2(n4461), .ZN(n5757) );
  NAND2_X1 U7292 ( .A1(n5905), .A2(n5755), .ZN(n5756) );
  NAND2_X1 U7293 ( .A1(n5759), .A2(n5758), .ZN(n5774) );
  NAND2_X1 U7294 ( .A1(n5761), .A2(n5760), .ZN(n5762) );
  NAND2_X1 U7295 ( .A1(n5786), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5765) );
  NAND2_X1 U7296 ( .A1(n4464), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5764) );
  NAND2_X1 U7297 ( .A1(n5785), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5763) );
  AND3_X1 U7298 ( .A1(n5765), .A2(n5764), .A3(n5763), .ZN(n5767) );
  NAND2_X1 U7299 ( .A1(n5822), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5766) );
  NAND2_X1 U7300 ( .A1(n5767), .A2(n5766), .ZN(n8177) );
  INV_X1 U7301 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5768) );
  OAI21_X1 U7302 ( .B1(n5770), .B2(n5769), .A(n5768), .ZN(n5771) );
  AND2_X1 U7303 ( .A1(n5772), .A2(n5771), .ZN(n8662) );
  MUX2_X1 U7304 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8662), .S(n5899), .Z(n9852) );
  NAND2_X1 U7305 ( .A1(n8177), .A2(n9852), .ZN(n6788) );
  NOR2_X1 U7306 ( .A1(n6196), .A2(n9852), .ZN(n5773) );
  NAND2_X1 U7307 ( .A1(n5785), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5778) );
  NAND2_X1 U7308 ( .A1(n5822), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5777) );
  NAND2_X1 U7309 ( .A1(n4463), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5776) );
  NAND2_X1 U7310 ( .A1(n5786), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5775) );
  OR2_X1 U7311 ( .A1(n6794), .A2(n5791), .ZN(n5780) );
  OR2_X1 U7312 ( .A1(n5779), .A2(n5721), .ZN(n5794) );
  XNOR2_X1 U7313 ( .A(n6803), .B(n6196), .ZN(n5781) );
  XNOR2_X1 U7314 ( .A(n5780), .B(n5781), .ZN(n6832) );
  INV_X1 U7315 ( .A(n5780), .ZN(n5783) );
  INV_X1 U7316 ( .A(n5781), .ZN(n5782) );
  NAND2_X1 U7317 ( .A1(n5783), .A2(n5782), .ZN(n5784) );
  INV_X1 U7318 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10240) );
  NAND2_X1 U7319 ( .A1(n5822), .A2(n10240), .ZN(n5790) );
  NAND2_X1 U7320 ( .A1(n5785), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U7321 ( .A1(n4464), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5788) );
  NAND2_X1 U7322 ( .A1(n5786), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5787) );
  OR2_X1 U7323 ( .A1(n6806), .A2(n5791), .ZN(n5801) );
  NAND2_X1 U7324 ( .A1(n5851), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5798) );
  NAND2_X1 U7325 ( .A1(n5794), .A2(n10237), .ZN(n5795) );
  NAND2_X1 U7326 ( .A1(n5795), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5796) );
  XNOR2_X1 U7327 ( .A(n5796), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6981) );
  NAND2_X1 U7328 ( .A1(n5809), .A2(n6981), .ZN(n5797) );
  XNOR2_X1 U7329 ( .A(n6196), .B(n6892), .ZN(n5799) );
  XNOR2_X1 U7330 ( .A(n5801), .B(n5799), .ZN(n6888) );
  INV_X1 U7331 ( .A(n5799), .ZN(n5800) );
  NOR2_X1 U7332 ( .A1(n5801), .A2(n5800), .ZN(n5802) );
  NAND2_X1 U7333 ( .A1(n5785), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5808) );
  INV_X2 U7334 ( .A(n6241), .ZN(n7955) );
  NAND2_X1 U7335 ( .A1(n7955), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5807) );
  NAND2_X1 U7336 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5825) );
  OAI21_X1 U7337 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5825), .ZN(n7316) );
  INV_X1 U7338 ( .A(n7316), .ZN(n5803) );
  NAND2_X1 U7339 ( .A1(n5822), .A2(n5803), .ZN(n5806) );
  NAND2_X1 U7340 ( .A1(n4463), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5805) );
  NOR2_X1 U7341 ( .A1(n7262), .A2(n5791), .ZN(n5816) );
  NAND2_X1 U7342 ( .A1(n5851), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5815) );
  NAND2_X1 U7343 ( .A1(n5811), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5812) );
  MUX2_X1 U7344 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5812), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5813) );
  AND2_X1 U7345 ( .A1(n5810), .A2(n5813), .ZN(n6982) );
  NAND2_X1 U7346 ( .A1(n4467), .A2(n6982), .ZN(n5814) );
  XNOR2_X1 U7347 ( .A(n6196), .B(n7322), .ZN(n5817) );
  NAND2_X1 U7348 ( .A1(n5816), .A2(n5817), .ZN(n5820) );
  INV_X1 U7349 ( .A(n5816), .ZN(n5819) );
  INV_X1 U7350 ( .A(n5817), .ZN(n5818) );
  NAND2_X1 U7351 ( .A1(n5819), .A2(n5818), .ZN(n5821) );
  AND2_X1 U7352 ( .A1(n5820), .A2(n5821), .ZN(n6866) );
  NAND2_X1 U7353 ( .A1(n7955), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5830) );
  NAND2_X1 U7354 ( .A1(n5785), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5829) );
  INV_X1 U7355 ( .A(n5825), .ZN(n5823) );
  NAND2_X1 U7356 ( .A1(n5823), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5845) );
  INV_X1 U7357 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5824) );
  NAND2_X1 U7358 ( .A1(n5825), .A2(n5824), .ZN(n5826) );
  AND2_X1 U7359 ( .A1(n5845), .A2(n5826), .ZN(n7257) );
  NAND2_X1 U7360 ( .A1(n5822), .A2(n7257), .ZN(n5828) );
  NAND2_X1 U7361 ( .A1(n4463), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5827) );
  OR2_X1 U7362 ( .A1(n7287), .A2(n5791), .ZN(n5837) );
  NAND2_X1 U7363 ( .A1(n5851), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5836) );
  NAND2_X1 U7364 ( .A1(n5810), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5831) );
  MUX2_X1 U7365 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5831), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5834) );
  INV_X1 U7366 ( .A(n5832), .ZN(n5833) );
  NAND2_X1 U7367 ( .A1(n4467), .A2(n6984), .ZN(n5835) );
  XNOR2_X1 U7368 ( .A(n9860), .B(n6196), .ZN(n5838) );
  XNOR2_X1 U7369 ( .A(n5837), .B(n5838), .ZN(n6858) );
  INV_X1 U7370 ( .A(n5837), .ZN(n5840) );
  INV_X1 U7371 ( .A(n5838), .ZN(n5839) );
  NAND2_X1 U7372 ( .A1(n5840), .A2(n5839), .ZN(n5841) );
  NAND2_X1 U7373 ( .A1(n5785), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5850) );
  NAND2_X1 U7374 ( .A1(n7955), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5849) );
  INV_X1 U7375 ( .A(n5845), .ZN(n5843) );
  NAND2_X1 U7376 ( .A1(n5843), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5867) );
  INV_X1 U7377 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5844) );
  NAND2_X1 U7378 ( .A1(n5845), .A2(n5844), .ZN(n5846) );
  AND2_X1 U7379 ( .A1(n5867), .A2(n5846), .ZN(n7282) );
  NAND2_X1 U7380 ( .A1(n5822), .A2(n7282), .ZN(n5848) );
  NAND2_X1 U7381 ( .A1(n4464), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5847) );
  NOR2_X1 U7382 ( .A1(n7276), .A2(n5791), .ZN(n5855) );
  NAND2_X1 U7383 ( .A1(n7753), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n5854) );
  OR2_X1 U7384 ( .A1(n5832), .A2(n5721), .ZN(n5852) );
  XNOR2_X1 U7385 ( .A(n5852), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6986) );
  NAND2_X1 U7386 ( .A1(n4467), .A2(n6986), .ZN(n5853) );
  XNOR2_X1 U7387 ( .A(n6196), .B(n7326), .ZN(n5856) );
  NAND2_X1 U7388 ( .A1(n5855), .A2(n5856), .ZN(n5859) );
  INV_X1 U7389 ( .A(n5855), .ZN(n5858) );
  INV_X1 U7390 ( .A(n5856), .ZN(n5857) );
  NAND2_X1 U7391 ( .A1(n5858), .A2(n5857), .ZN(n5860) );
  AND2_X1 U7392 ( .A1(n5859), .A2(n5860), .ZN(n7071) );
  NAND2_X1 U7393 ( .A1(n7753), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n5864) );
  OR2_X1 U7394 ( .A1(n5861), .A2(n5721), .ZN(n5862) );
  XNOR2_X1 U7395 ( .A(n5862), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6989) );
  NAND2_X1 U7396 ( .A1(n4467), .A2(n6989), .ZN(n5863) );
  OAI211_X1 U7397 ( .C1(n5792), .C2(n6328), .A(n5864), .B(n5863), .ZN(n8004)
         );
  INV_X1 U7398 ( .A(n8004), .ZN(n9872) );
  XNOR2_X1 U7399 ( .A(n9872), .B(n6196), .ZN(n5874) );
  NAND2_X1 U7400 ( .A1(n7955), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5872) );
  NAND2_X1 U7401 ( .A1(n5785), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5871) );
  INV_X1 U7402 ( .A(n5867), .ZN(n5865) );
  NAND2_X1 U7403 ( .A1(n5865), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5878) );
  INV_X1 U7404 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5866) );
  NAND2_X1 U7405 ( .A1(n5867), .A2(n5866), .ZN(n5868) );
  AND2_X1 U7406 ( .A1(n5878), .A2(n5868), .ZN(n7079) );
  NAND2_X1 U7407 ( .A1(n5822), .A2(n7079), .ZN(n5870) );
  NAND2_X1 U7408 ( .A1(n4464), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5869) );
  NAND4_X1 U7409 ( .A1(n5872), .A2(n5871), .A3(n5870), .A4(n5869), .ZN(n9805)
         );
  NAND2_X1 U7410 ( .A1(n9805), .A2(n7966), .ZN(n5873) );
  XNOR2_X1 U7411 ( .A(n5874), .B(n5873), .ZN(n7077) );
  INV_X1 U7412 ( .A(n5873), .ZN(n5876) );
  INV_X1 U7413 ( .A(n5874), .ZN(n5875) );
  NAND2_X1 U7414 ( .A1(n5878), .A2(n5877), .ZN(n5879) );
  AND2_X1 U7415 ( .A1(n5893), .A2(n5879), .ZN(n9815) );
  NAND2_X1 U7416 ( .A1(n5822), .A2(n9815), .ZN(n5883) );
  NAND2_X1 U7417 ( .A1(n5785), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5882) );
  NAND2_X1 U7418 ( .A1(n4463), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5881) );
  NAND2_X1 U7419 ( .A1(n7955), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5880) );
  OR2_X1 U7420 ( .A1(n7369), .A2(n5791), .ZN(n5890) );
  NAND2_X1 U7421 ( .A1(n7753), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n5887) );
  NAND2_X1 U7422 ( .A1(n5884), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5885) );
  XNOR2_X1 U7423 ( .A(n5885), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6991) );
  NAND2_X1 U7424 ( .A1(n4467), .A2(n6991), .ZN(n5886) );
  OAI211_X1 U7425 ( .C1(n5792), .C2(n6331), .A(n5887), .B(n5886), .ZN(n9797)
         );
  XNOR2_X1 U7426 ( .A(n6196), .B(n9797), .ZN(n5888) );
  XNOR2_X1 U7427 ( .A(n5890), .B(n5888), .ZN(n7268) );
  INV_X1 U7428 ( .A(n5888), .ZN(n5889) );
  NAND2_X1 U7429 ( .A1(n7955), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5898) );
  NAND2_X1 U7430 ( .A1(n5785), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5897) );
  INV_X1 U7431 ( .A(n5893), .ZN(n5891) );
  NAND2_X1 U7432 ( .A1(n5891), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5914) );
  INV_X1 U7433 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U7434 ( .A1(n5893), .A2(n5892), .ZN(n5894) );
  AND2_X1 U7435 ( .A1(n5914), .A2(n5894), .ZN(n7378) );
  NAND2_X1 U7436 ( .A1(n5822), .A2(n7378), .ZN(n5896) );
  NAND2_X1 U7437 ( .A1(n4463), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5895) );
  NOR2_X1 U7438 ( .A1(n7398), .A2(n5791), .ZN(n5908) );
  INV_X1 U7439 ( .A(n5900), .ZN(n5904) );
  NAND2_X1 U7440 ( .A1(n5901), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5902) );
  MUX2_X1 U7441 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5902), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n5903) );
  INV_X1 U7442 ( .A(n6993), .ZN(n7190) );
  NAND2_X1 U7443 ( .A1(n6333), .A2(n7752), .ZN(n5907) );
  NAND2_X1 U7444 ( .A1(n7753), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n5906) );
  OAI211_X1 U7445 ( .C1(n6998), .C2(n7190), .A(n5907), .B(n5906), .ZN(n7384)
         );
  XNOR2_X1 U7446 ( .A(n7384), .B(n6196), .ZN(n5909) );
  NAND2_X1 U7447 ( .A1(n5908), .A2(n5909), .ZN(n7345) );
  NAND2_X1 U7448 ( .A1(n7347), .A2(n7345), .ZN(n5912) );
  INV_X1 U7449 ( .A(n5908), .ZN(n5911) );
  INV_X1 U7450 ( .A(n5909), .ZN(n5910) );
  NAND2_X1 U7451 ( .A1(n5911), .A2(n5910), .ZN(n7344) );
  NAND2_X1 U7452 ( .A1(n7955), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U7453 ( .A1(n5785), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5918) );
  NAND2_X1 U7454 ( .A1(n5914), .A2(n5913), .ZN(n5915) );
  AND2_X1 U7455 ( .A1(n5938), .A2(n5915), .ZN(n6263) );
  NAND2_X1 U7456 ( .A1(n5822), .A2(n6263), .ZN(n5917) );
  NAND2_X1 U7457 ( .A1(n4463), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5916) );
  NOR2_X1 U7458 ( .A1(n7910), .A2(n5791), .ZN(n5925) );
  NAND2_X1 U7459 ( .A1(n6340), .A2(n7752), .ZN(n5924) );
  OR2_X1 U7460 ( .A1(n5900), .A2(n5721), .ZN(n5921) );
  INV_X1 U7461 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5920) );
  OR2_X1 U7462 ( .A1(n5921), .A2(n5920), .ZN(n5922) );
  NAND2_X1 U7463 ( .A1(n5921), .A2(n5920), .ZN(n5932) );
  AOI22_X1 U7464 ( .A1(n7753), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n4467), .B2(
        n7146), .ZN(n5923) );
  NAND2_X1 U7465 ( .A1(n5924), .A2(n5923), .ZN(n7409) );
  XNOR2_X1 U7466 ( .A(n7409), .B(n6196), .ZN(n5926) );
  NAND2_X1 U7467 ( .A1(n5925), .A2(n5926), .ZN(n5931) );
  INV_X1 U7468 ( .A(n5925), .ZN(n5928) );
  INV_X1 U7469 ( .A(n5926), .ZN(n5927) );
  NAND2_X1 U7470 ( .A1(n5928), .A2(n5927), .ZN(n5929) );
  NAND2_X1 U7471 ( .A1(n5931), .A2(n5929), .ZN(n6262) );
  NAND2_X1 U7472 ( .A1(n6338), .A2(n7752), .ZN(n5935) );
  NAND2_X1 U7473 ( .A1(n5932), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5933) );
  XNOR2_X1 U7474 ( .A(n5933), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8183) );
  AOI22_X1 U7475 ( .A1(n7753), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n4467), .B2(
        n8183), .ZN(n5934) );
  NAND2_X1 U7476 ( .A1(n5935), .A2(n5934), .ZN(n7517) );
  XNOR2_X1 U7477 ( .A(n7517), .B(n6196), .ZN(n5944) );
  NAND2_X1 U7478 ( .A1(n7955), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5943) );
  NAND2_X1 U7479 ( .A1(n5785), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5942) );
  INV_X1 U7480 ( .A(n5938), .ZN(n5936) );
  NAND2_X1 U7481 ( .A1(n5936), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5954) );
  INV_X1 U7482 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5937) );
  NAND2_X1 U7483 ( .A1(n5938), .A2(n5937), .ZN(n5939) );
  AND2_X1 U7484 ( .A1(n5954), .A2(n5939), .ZN(n7907) );
  NAND2_X1 U7485 ( .A1(n5822), .A2(n7907), .ZN(n5941) );
  NAND2_X1 U7486 ( .A1(n4464), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5940) );
  NOR2_X1 U7487 ( .A1(n7828), .A2(n5791), .ZN(n5945) );
  NAND2_X1 U7488 ( .A1(n5944), .A2(n5945), .ZN(n5949) );
  INV_X1 U7489 ( .A(n5944), .ZN(n5947) );
  INV_X1 U7490 ( .A(n5945), .ZN(n5946) );
  NAND2_X1 U7491 ( .A1(n5947), .A2(n5946), .ZN(n5948) );
  AND2_X1 U7492 ( .A1(n5949), .A2(n5948), .ZN(n7904) );
  NAND2_X1 U7493 ( .A1(n7905), .A2(n7904), .ZN(n7903) );
  NAND2_X1 U7494 ( .A1(n6345), .A2(n7752), .ZN(n5953) );
  NAND2_X1 U7495 ( .A1(n5950), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5951) );
  XNOR2_X1 U7496 ( .A(n5951), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7062) );
  AOI22_X1 U7497 ( .A1(n7753), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n4467), .B2(
        n7062), .ZN(n5952) );
  XNOR2_X1 U7498 ( .A(n7829), .B(n6118), .ZN(n5960) );
  NAND2_X1 U7499 ( .A1(n7955), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U7500 ( .A1(n5785), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5958) );
  NAND2_X1 U7501 ( .A1(n5954), .A2(n10132), .ZN(n5955) );
  AND2_X1 U7502 ( .A1(n5968), .A2(n5955), .ZN(n7830) );
  NAND2_X1 U7503 ( .A1(n5822), .A2(n7830), .ZN(n5957) );
  NAND2_X1 U7504 ( .A1(n4464), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5956) );
  NOR2_X1 U7505 ( .A1(n7906), .A2(n5791), .ZN(n5961) );
  XNOR2_X1 U7506 ( .A(n5960), .B(n5961), .ZN(n7826) );
  INV_X1 U7507 ( .A(n5960), .ZN(n5962) );
  NAND2_X1 U7508 ( .A1(n5962), .A2(n5961), .ZN(n5963) );
  NAND2_X1 U7509 ( .A1(n6348), .A2(n7752), .ZN(n5966) );
  OR2_X1 U7510 ( .A1(n5950), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U7511 ( .A1(n5964), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5978) );
  XNOR2_X1 U7512 ( .A(n5978), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7029) );
  AOI22_X1 U7513 ( .A1(n7753), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n4467), .B2(
        n7029), .ZN(n5965) );
  XNOR2_X1 U7514 ( .A(n8623), .B(n6196), .ZN(n5974) );
  NAND2_X1 U7515 ( .A1(n7955), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5973) );
  NAND2_X1 U7516 ( .A1(n5785), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U7517 ( .A1(n5968), .A2(n5967), .ZN(n5969) );
  AND2_X1 U7518 ( .A1(n5987), .A2(n5969), .ZN(n7889) );
  NAND2_X1 U7519 ( .A1(n5822), .A2(n7889), .ZN(n5971) );
  NAND2_X1 U7520 ( .A1(n4464), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5970) );
  NOR2_X1 U7521 ( .A1(n8040), .A2(n5791), .ZN(n5975) );
  AND2_X1 U7522 ( .A1(n5974), .A2(n5975), .ZN(n7880) );
  INV_X1 U7523 ( .A(n5974), .ZN(n5977) );
  INV_X1 U7524 ( .A(n5975), .ZN(n5976) );
  NAND2_X1 U7525 ( .A1(n6356), .A2(n7752), .ZN(n5984) );
  NAND2_X1 U7526 ( .A1(n5978), .A2(n10206), .ZN(n5979) );
  NAND2_X1 U7527 ( .A1(n5979), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7528 ( .A1(n5981), .A2(n5980), .ZN(n6003) );
  OR2_X1 U7529 ( .A1(n5981), .A2(n5980), .ZN(n5982) );
  AOI22_X1 U7530 ( .A1(n7753), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n4467), .B2(
        n8192), .ZN(n5983) );
  NAND2_X1 U7531 ( .A1(n5984), .A2(n5983), .ZN(n7601) );
  XNOR2_X1 U7532 ( .A(n7601), .B(n6118), .ZN(n5993) );
  NAND2_X1 U7533 ( .A1(n7955), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5992) );
  NAND2_X1 U7534 ( .A1(n5785), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5991) );
  INV_X1 U7535 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7536 ( .A1(n5987), .A2(n5986), .ZN(n5988) );
  AND2_X1 U7537 ( .A1(n6013), .A2(n5988), .ZN(n7800) );
  NAND2_X1 U7538 ( .A1(n5822), .A2(n7800), .ZN(n5990) );
  NAND2_X1 U7539 ( .A1(n4464), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5989) );
  OR2_X1 U7540 ( .A1(n7936), .A2(n5791), .ZN(n5994) );
  NAND2_X1 U7541 ( .A1(n5993), .A2(n5994), .ZN(n5998) );
  INV_X1 U7542 ( .A(n5993), .ZN(n5996) );
  INV_X1 U7543 ( .A(n5994), .ZN(n5995) );
  NAND2_X1 U7544 ( .A1(n5996), .A2(n5995), .ZN(n5997) );
  AND2_X1 U7545 ( .A1(n5998), .A2(n5997), .ZN(n7796) );
  NAND2_X1 U7546 ( .A1(n7795), .A2(n7796), .ZN(n7794) );
  NAND2_X2 U7547 ( .A1(n7794), .A2(n5998), .ZN(n7842) );
  NAND2_X1 U7548 ( .A1(n7955), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U7549 ( .A1(n5785), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6001) );
  XNOR2_X1 U7550 ( .A(n6013), .B(P2_REG3_REG_15__SCAN_IN), .ZN(n8517) );
  NAND2_X1 U7551 ( .A1(n5822), .A2(n8517), .ZN(n6000) );
  NAND2_X1 U7552 ( .A1(n4463), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5999) );
  NOR2_X1 U7553 ( .A1(n7849), .A2(n5791), .ZN(n7934) );
  NAND2_X1 U7554 ( .A1(n6457), .A2(n7752), .ZN(n6006) );
  NAND2_X1 U7555 ( .A1(n6003), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6004) );
  XNOR2_X1 U7556 ( .A(n6004), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8206) );
  AOI22_X1 U7557 ( .A1(n7753), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n4467), .B2(
        n8206), .ZN(n6005) );
  XNOR2_X1 U7558 ( .A(n8612), .B(n6196), .ZN(n7843) );
  NAND2_X1 U7559 ( .A1(n6543), .A2(n7752), .ZN(n6010) );
  NAND2_X1 U7560 ( .A1(n6007), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6008) );
  XNOR2_X1 U7561 ( .A(n6008), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8232) );
  AOI22_X1 U7562 ( .A1(n7753), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n4467), .B2(
        n8232), .ZN(n6009) );
  XNOR2_X1 U7563 ( .A(n8606), .B(n6118), .ZN(n6019) );
  NAND2_X1 U7564 ( .A1(n5785), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U7565 ( .A1(n4464), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6017) );
  INV_X1 U7566 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6011) );
  INV_X1 U7567 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6012) );
  OAI21_X1 U7568 ( .B1(n6013), .B2(n6011), .A(n6012), .ZN(n6014) );
  AND2_X1 U7569 ( .A1(n6014), .A2(n6032), .ZN(n8506) );
  NAND2_X1 U7570 ( .A1(n5822), .A2(n8506), .ZN(n6016) );
  NAND2_X1 U7571 ( .A1(n7955), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6015) );
  OR2_X1 U7572 ( .A1(n8166), .A2(n5791), .ZN(n6020) );
  NAND2_X1 U7573 ( .A1(n6019), .A2(n6020), .ZN(n7846) );
  OAI21_X1 U7574 ( .B1(n7934), .B2(n7843), .A(n7846), .ZN(n6025) );
  NAND3_X1 U7575 ( .A1(n7846), .A2(n7934), .A3(n7843), .ZN(n6023) );
  INV_X1 U7576 ( .A(n6019), .ZN(n6022) );
  INV_X1 U7577 ( .A(n6020), .ZN(n6021) );
  NAND2_X1 U7578 ( .A1(n6022), .A2(n6021), .ZN(n7845) );
  AND2_X1 U7579 ( .A1(n6023), .A2(n7845), .ZN(n6024) );
  OAI21_X2 U7580 ( .B1(n7842), .B2(n6025), .A(n6024), .ZN(n7855) );
  NAND2_X1 U7581 ( .A1(n6601), .A2(n7752), .ZN(n6030) );
  NAND2_X1 U7582 ( .A1(n6027), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6028) );
  XNOR2_X1 U7583 ( .A(n6028), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8253) );
  AOI22_X1 U7584 ( .A1(n7753), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n4467), .B2(
        n8253), .ZN(n6029) );
  XNOR2_X1 U7585 ( .A(n8603), .B(n6118), .ZN(n6038) );
  NAND2_X1 U7586 ( .A1(n7955), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U7587 ( .A1(n5785), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6036) );
  INV_X1 U7588 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8230) );
  NAND2_X1 U7589 ( .A1(n6032), .A2(n8230), .ZN(n6033) );
  AND2_X1 U7590 ( .A1(n6060), .A2(n6033), .ZN(n8496) );
  NAND2_X1 U7591 ( .A1(n5822), .A2(n8496), .ZN(n6035) );
  NAND2_X1 U7592 ( .A1(n4463), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6034) );
  NOR2_X1 U7593 ( .A1(n7918), .A2(n5791), .ZN(n6039) );
  XNOR2_X1 U7594 ( .A(n6038), .B(n6039), .ZN(n7854) );
  NAND2_X1 U7595 ( .A1(n7855), .A2(n7854), .ZN(n6042) );
  INV_X1 U7596 ( .A(n6038), .ZN(n6040) );
  NAND2_X1 U7597 ( .A1(n6040), .A2(n6039), .ZN(n6041) );
  NAND2_X1 U7598 ( .A1(n6042), .A2(n6041), .ZN(n7917) );
  NAND2_X1 U7599 ( .A1(n6839), .A2(n7752), .ZN(n6045) );
  XNOR2_X1 U7600 ( .A(n6043), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8261) );
  AOI22_X1 U7601 ( .A1(n7753), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n4467), .B2(
        n8261), .ZN(n6044) );
  XNOR2_X1 U7602 ( .A(n8596), .B(n6118), .ZN(n6050) );
  NAND2_X1 U7603 ( .A1(n5785), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U7604 ( .A1(n7955), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6048) );
  XNOR2_X1 U7605 ( .A(n6060), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n7920) );
  NAND2_X1 U7606 ( .A1(n5822), .A2(n7920), .ZN(n6047) );
  NAND2_X1 U7607 ( .A1(n4464), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6046) );
  NOR2_X1 U7608 ( .A1(n8492), .A2(n5791), .ZN(n6051) );
  XNOR2_X1 U7609 ( .A(n6050), .B(n6051), .ZN(n7916) );
  NAND2_X1 U7610 ( .A1(n7917), .A2(n7916), .ZN(n6054) );
  INV_X1 U7611 ( .A(n6050), .ZN(n6052) );
  NAND2_X1 U7612 ( .A1(n6052), .A2(n6051), .ZN(n6053) );
  NAND2_X1 U7613 ( .A1(n6054), .A2(n6053), .ZN(n7812) );
  INV_X1 U7614 ( .A(n7812), .ZN(n6070) );
  NAND2_X1 U7615 ( .A1(n6923), .A2(n7752), .ZN(n6056) );
  AOI22_X1 U7616 ( .A1(n7753), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n4467), .B2(
        n8273), .ZN(n6055) );
  XNOR2_X1 U7617 ( .A(n8482), .B(n6118), .ZN(n6066) );
  NAND2_X1 U7618 ( .A1(n7955), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7619 ( .A1(n5785), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6064) );
  INV_X1 U7620 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6058) );
  INV_X1 U7621 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6057) );
  OAI21_X1 U7622 ( .B1(n6060), .B2(n6058), .A(n6057), .ZN(n6061) );
  NAND2_X1 U7623 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n6059) );
  AND2_X1 U7624 ( .A1(n6061), .A2(n6075), .ZN(n8479) );
  NAND2_X1 U7625 ( .A1(n5822), .A2(n8479), .ZN(n6063) );
  NAND2_X1 U7626 ( .A1(n4464), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6062) );
  NOR2_X1 U7627 ( .A1(n8287), .A2(n5791), .ZN(n6067) );
  INV_X1 U7628 ( .A(n6066), .ZN(n6069) );
  INV_X1 U7629 ( .A(n6067), .ZN(n6068) );
  NAND2_X1 U7630 ( .A1(n6069), .A2(n6068), .ZN(n7810) );
  NAND2_X1 U7631 ( .A1(n7085), .A2(n7752), .ZN(n6072) );
  NAND2_X1 U7632 ( .A1(n7753), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6071) );
  XNOR2_X1 U7633 ( .A(n8586), .B(n6196), .ZN(n6081) );
  NAND2_X1 U7634 ( .A1(n7955), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7635 ( .A1(n5785), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6079) );
  INV_X1 U7636 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U7637 ( .A1(n6075), .A2(n6074), .ZN(n6076) );
  AND2_X1 U7638 ( .A1(n6097), .A2(n6076), .ZN(n8456) );
  NAND2_X1 U7639 ( .A1(n5822), .A2(n8456), .ZN(n6078) );
  NAND2_X1 U7640 ( .A1(n4463), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6077) );
  NOR2_X1 U7641 ( .A1(n8475), .A2(n5791), .ZN(n6082) );
  NAND2_X1 U7642 ( .A1(n6081), .A2(n6082), .ZN(n7817) );
  INV_X1 U7643 ( .A(n6081), .ZN(n6084) );
  INV_X1 U7644 ( .A(n6082), .ZN(n6083) );
  NAND2_X1 U7645 ( .A1(n6084), .A2(n6083), .ZN(n6085) );
  AND2_X1 U7646 ( .A1(n7817), .A2(n6085), .ZN(n7873) );
  NAND2_X1 U7647 ( .A1(n7470), .A2(n7752), .ZN(n6087) );
  NAND2_X1 U7648 ( .A1(n7753), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6086) );
  XNOR2_X1 U7649 ( .A(n8576), .B(n6196), .ZN(n7895) );
  INV_X1 U7650 ( .A(n7895), .ZN(n6093) );
  NAND2_X1 U7651 ( .A1(n7955), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U7652 ( .A1(n5785), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6091) );
  INV_X1 U7653 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n7820) );
  NAND2_X1 U7654 ( .A1(n6099), .A2(n10204), .ZN(n6088) );
  AND2_X1 U7655 ( .A1(n6129), .A2(n6088), .ZN(n8430) );
  NAND2_X1 U7656 ( .A1(n5822), .A2(n8430), .ZN(n6090) );
  NAND2_X1 U7657 ( .A1(n4463), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6089) );
  NOR2_X1 U7658 ( .A1(n8296), .A2(n5791), .ZN(n6094) );
  INV_X1 U7659 ( .A(n6094), .ZN(n7894) );
  NAND2_X1 U7660 ( .A1(n6093), .A2(n7894), .ZN(n6111) );
  INV_X1 U7661 ( .A(n6111), .ZN(n6107) );
  NAND2_X1 U7662 ( .A1(n7895), .A2(n6094), .ZN(n6105) );
  NAND2_X1 U7663 ( .A1(n7089), .A2(n7752), .ZN(n6096) );
  NAND2_X1 U7664 ( .A1(n7753), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6095) );
  XNOR2_X1 U7665 ( .A(n8444), .B(n6196), .ZN(n6110) );
  INV_X1 U7666 ( .A(n6110), .ZN(n6104) );
  NAND2_X1 U7667 ( .A1(n7955), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7668 ( .A1(n5785), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6102) );
  NAND2_X1 U7669 ( .A1(n6097), .A2(n7820), .ZN(n6098) );
  AND2_X1 U7670 ( .A1(n6099), .A2(n6098), .ZN(n8442) );
  NAND2_X1 U7671 ( .A1(n5822), .A2(n8442), .ZN(n6101) );
  NAND2_X1 U7672 ( .A1(n4463), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6100) );
  NOR2_X1 U7673 ( .A1(n8294), .A2(n5791), .ZN(n6109) );
  NAND2_X1 U7674 ( .A1(n6104), .A2(n6109), .ZN(n7892) );
  AND2_X1 U7675 ( .A1(n6105), .A2(n7892), .ZN(n6106) );
  INV_X1 U7676 ( .A(n6108), .ZN(n6113) );
  XNOR2_X1 U7677 ( .A(n6110), .B(n6109), .ZN(n7819) );
  AND2_X1 U7678 ( .A1(n7819), .A2(n6111), .ZN(n6112) );
  NAND2_X1 U7679 ( .A1(n7472), .A2(n7752), .ZN(n6115) );
  NAND2_X1 U7680 ( .A1(n7753), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6114) );
  XNOR2_X1 U7681 ( .A(n8570), .B(n6196), .ZN(n6137) );
  XNOR2_X1 U7682 ( .A(n6136), .B(n6137), .ZN(n7803) );
  NAND2_X1 U7683 ( .A1(n7556), .A2(n7752), .ZN(n6117) );
  NAND2_X1 U7684 ( .A1(n7753), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6116) );
  XNOR2_X1 U7685 ( .A(n8565), .B(n6118), .ZN(n7863) );
  NAND2_X1 U7686 ( .A1(n7955), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U7687 ( .A1(n5785), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6119) );
  AND2_X1 U7688 ( .A1(n6120), .A2(n6119), .ZN(n6128) );
  INV_X1 U7689 ( .A(n6129), .ZN(n6122) );
  AND2_X1 U7690 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(P2_REG3_REG_24__SCAN_IN), 
        .ZN(n6121) );
  NAND2_X1 U7691 ( .A1(n6122), .A2(n6121), .ZN(n6148) );
  INV_X1 U7692 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n6124) );
  INV_X1 U7693 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6123) );
  OAI21_X1 U7694 ( .B1(n6129), .B2(n6124), .A(n6123), .ZN(n6125) );
  NAND2_X1 U7695 ( .A1(n6148), .A2(n6125), .ZN(n8394) );
  NAND2_X1 U7696 ( .A1(n4464), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6126) );
  NAND2_X1 U7697 ( .A1(n7955), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6133) );
  XNOR2_X1 U7698 ( .A(n6129), .B(P2_REG3_REG_23__SCAN_IN), .ZN(n8416) );
  NAND2_X1 U7699 ( .A1(n8416), .A2(n5822), .ZN(n6132) );
  NAND2_X1 U7700 ( .A1(n5785), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6131) );
  NAND2_X1 U7701 ( .A1(n4464), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6130) );
  NAND4_X1 U7702 ( .A1(n6133), .A2(n6132), .A3(n6131), .A4(n6130), .ZN(n8436)
         );
  NAND2_X1 U7703 ( .A1(n8436), .A2(n7966), .ZN(n7804) );
  AOI21_X1 U7704 ( .B1(n7863), .B2(n8377), .A(n7804), .ZN(n6134) );
  NAND2_X1 U7705 ( .A1(n7803), .A2(n6134), .ZN(n6143) );
  NOR2_X1 U7706 ( .A1(n8377), .A2(n5791), .ZN(n6140) );
  INV_X1 U7707 ( .A(n7863), .ZN(n6135) );
  OR2_X1 U7708 ( .A1(n6140), .A2(n6135), .ZN(n6139) );
  INV_X1 U7709 ( .A(n6136), .ZN(n6138) );
  AND2_X1 U7710 ( .A1(n6138), .A2(n6137), .ZN(n7861) );
  NAND2_X1 U7711 ( .A1(n6139), .A2(n7861), .ZN(n6142) );
  INV_X1 U7712 ( .A(n6140), .ZN(n7867) );
  NAND2_X1 U7713 ( .A1(n7572), .A2(n7752), .ZN(n6145) );
  NAND2_X1 U7714 ( .A1(n7753), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6144) );
  XNOR2_X1 U7715 ( .A(n8562), .B(n6196), .ZN(n6153) );
  INV_X1 U7716 ( .A(n6148), .ZN(n6146) );
  NAND2_X1 U7717 ( .A1(n6146), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6161) );
  INV_X1 U7718 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7719 ( .A1(n6148), .A2(n6147), .ZN(n6149) );
  NAND2_X1 U7720 ( .A1(n6161), .A2(n6149), .ZN(n8383) );
  AOI22_X1 U7721 ( .A1(n7955), .A2(P2_REG1_REG_25__SCAN_IN), .B1(n5785), .B2(
        P2_REG0_REG_25__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7722 ( .A1(n4464), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6150) );
  NOR2_X1 U7723 ( .A1(n8404), .A2(n5791), .ZN(n6154) );
  NAND2_X1 U7724 ( .A1(n6153), .A2(n6154), .ZN(n6158) );
  INV_X1 U7725 ( .A(n6153), .ZN(n6156) );
  INV_X1 U7726 ( .A(n6154), .ZN(n6155) );
  NAND2_X1 U7727 ( .A1(n6156), .A2(n6155), .ZN(n6157) );
  AND2_X1 U7728 ( .A1(n6158), .A2(n6157), .ZN(n7836) );
  NAND2_X1 U7729 ( .A1(n7590), .A2(n7752), .ZN(n6160) );
  NAND2_X1 U7730 ( .A1(n7753), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6159) );
  XNOR2_X1 U7731 ( .A(n8557), .B(n6196), .ZN(n6166) );
  INV_X1 U7732 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n7928) );
  NAND2_X1 U7733 ( .A1(n6161), .A2(n7928), .ZN(n6162) );
  NAND2_X1 U7734 ( .A1(n8367), .A2(n5822), .ZN(n6165) );
  AOI22_X1 U7735 ( .A1(n7955), .A2(P2_REG1_REG_26__SCAN_IN), .B1(n5785), .B2(
        P2_REG0_REG_26__SCAN_IN), .ZN(n6164) );
  NAND2_X1 U7736 ( .A1(n4463), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6163) );
  NOR2_X1 U7737 ( .A1(n8378), .A2(n5791), .ZN(n6167) );
  NAND2_X1 U7738 ( .A1(n6166), .A2(n6167), .ZN(n6171) );
  INV_X1 U7739 ( .A(n6166), .ZN(n6169) );
  INV_X1 U7740 ( .A(n6167), .ZN(n6168) );
  NAND2_X1 U7741 ( .A1(n6169), .A2(n6168), .ZN(n6170) );
  AND2_X1 U7742 ( .A1(n6171), .A2(n6170), .ZN(n7926) );
  NAND2_X1 U7743 ( .A1(n7925), .A2(n6171), .ZN(n7789) );
  NAND2_X1 U7744 ( .A1(n7596), .A2(n7752), .ZN(n6173) );
  NAND2_X1 U7745 ( .A1(n7753), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6172) );
  XNOR2_X1 U7746 ( .A(n8550), .B(n6196), .ZN(n6184) );
  INV_X1 U7747 ( .A(n6176), .ZN(n6174) );
  NAND2_X1 U7748 ( .A1(n6174), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6190) );
  INV_X1 U7749 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U7750 ( .A1(n6176), .A2(n6175), .ZN(n6177) );
  NAND2_X1 U7751 ( .A1(n6190), .A2(n6177), .ZN(n8346) );
  INV_X1 U7752 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8347) );
  NAND2_X1 U7753 ( .A1(n7955), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U7754 ( .A1(n5785), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6179) );
  OAI211_X1 U7755 ( .C1(n8347), .C2(n7959), .A(n6180), .B(n6179), .ZN(n6181)
         );
  INV_X1 U7756 ( .A(n6181), .ZN(n6182) );
  NOR2_X1 U7757 ( .A1(n8309), .A2(n5791), .ZN(n6185) );
  NAND2_X1 U7758 ( .A1(n6184), .A2(n6185), .ZN(n6189) );
  INV_X1 U7759 ( .A(n6184), .ZN(n6187) );
  INV_X1 U7760 ( .A(n6185), .ZN(n6186) );
  NAND2_X1 U7761 ( .A1(n6187), .A2(n6186), .ZN(n6188) );
  AND2_X1 U7762 ( .A1(n6189), .A2(n6188), .ZN(n7788) );
  NAND2_X1 U7763 ( .A1(n7789), .A2(n7788), .ZN(n7787) );
  NAND2_X1 U7764 ( .A1(n7787), .A2(n6189), .ZN(n6199) );
  INV_X1 U7765 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6251) );
  NAND2_X1 U7766 ( .A1(n6190), .A2(n6251), .ZN(n6191) );
  INV_X1 U7767 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7768 ( .A1(n7955), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6193) );
  NAND2_X1 U7769 ( .A1(n5785), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6192) );
  OAI211_X1 U7770 ( .C1(n6194), .C2(n7959), .A(n6193), .B(n6192), .ZN(n6195)
         );
  OR2_X1 U7771 ( .A1(n8311), .A2(n5791), .ZN(n6197) );
  XNOR2_X1 U7772 ( .A(n6197), .B(n6196), .ZN(n6198) );
  XNOR2_X1 U7773 ( .A(n6199), .B(n6198), .ZN(n6237) );
  NAND2_X1 U7774 ( .A1(n6206), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6200) );
  MUX2_X1 U7775 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6200), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6203) );
  INV_X1 U7776 ( .A(n6201), .ZN(n6202) );
  NOR2_X1 U7777 ( .A1(n4565), .A2(n5721), .ZN(n6204) );
  MUX2_X1 U7778 ( .A(n5721), .B(n6204), .S(P2_IR_REG_25__SCAN_IN), .Z(n6205)
         );
  NAND2_X1 U7779 ( .A1(n6207), .A2(n6206), .ZN(n7589) );
  NAND2_X1 U7780 ( .A1(n6230), .A2(n6229), .ZN(n6211) );
  XNOR2_X1 U7781 ( .A(n7571), .B(P2_B_REG_SCAN_IN), .ZN(n6214) );
  NAND2_X1 U7782 ( .A1(n7589), .A2(n6214), .ZN(n6215) );
  INV_X1 U7783 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10076) );
  AND2_X1 U7784 ( .A1(n7589), .A2(n7595), .ZN(n9849) );
  NOR4_X1 U7785 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6220) );
  NOR4_X1 U7786 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n6219) );
  NOR4_X1 U7787 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6218) );
  NOR4_X1 U7788 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6217) );
  NAND4_X1 U7789 ( .A1(n6220), .A2(n6219), .A3(n6218), .A4(n6217), .ZN(n6226)
         );
  NOR2_X1 U7790 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .ZN(
        n6224) );
  NOR4_X1 U7791 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6223) );
  NOR4_X1 U7792 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n6222) );
  NOR4_X1 U7793 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n6221) );
  NAND4_X1 U7794 ( .A1(n6224), .A2(n6223), .A3(n6222), .A4(n6221), .ZN(n6225)
         );
  OAI21_X1 U7795 ( .B1(n6226), .B2(n6225), .A(n9843), .ZN(n6621) );
  INV_X1 U7796 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9846) );
  AND2_X1 U7797 ( .A1(n6621), .A2(n6704), .ZN(n6228) );
  NAND2_X1 U7798 ( .A1(n7252), .A2(n6228), .ZN(n6248) );
  AND2_X1 U7799 ( .A1(n9905), .A2(n6634), .ZN(n6232) );
  NAND2_X1 U7800 ( .A1(n9462), .A2(n7752), .ZN(n6234) );
  NAND2_X1 U7801 ( .A1(n7753), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6233) );
  AND2_X1 U7802 ( .A1(n8152), .A2(n6231), .ZN(n7256) );
  INV_X1 U7803 ( .A(n6622), .ZN(n6247) );
  INV_X2 U7804 ( .A(n8345), .ZN(n9838) );
  AOI21_X2 U7805 ( .B1(n6244), .B2(n7256), .A(n9838), .ZN(n7933) );
  OAI21_X1 U7806 ( .B1(n6237), .B2(n7944), .A(n7933), .ZN(n6256) );
  INV_X1 U7807 ( .A(n6238), .ZN(n8319) );
  INV_X1 U7808 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n10271) );
  NAND2_X1 U7809 ( .A1(n4464), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6240) );
  NAND2_X1 U7810 ( .A1(n5785), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6239) );
  OAI211_X1 U7811 ( .C1(n6241), .C2(n10271), .A(n6240), .B(n6239), .ZN(n6242)
         );
  AOI21_X1 U7812 ( .B1(n8319), .B2(n5822), .A(n6242), .ZN(n8164) );
  NAND2_X1 U7813 ( .A1(n6244), .A2(n6243), .ZN(n7929) );
  INV_X1 U7814 ( .A(n7003), .ZN(n6245) );
  OAI22_X1 U7815 ( .A1(n8164), .A2(n7938), .B1(n7937), .B2(n8309), .ZN(n6246)
         );
  INV_X1 U7816 ( .A(n6246), .ZN(n6255) );
  NAND2_X1 U7817 ( .A1(n6248), .A2(n6247), .ZN(n6769) );
  AND2_X1 U7818 ( .A1(n8159), .A2(n6972), .ZN(n6620) );
  INV_X1 U7819 ( .A(n6620), .ZN(n6249) );
  NAND4_X1 U7820 ( .A1(n6769), .A2(n6974), .A3(n6352), .A4(n6249), .ZN(n6250)
         );
  INV_X1 U7821 ( .A(n8328), .ZN(n6252) );
  OAI22_X1 U7822 ( .A1(n7909), .A2(n6252), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6251), .ZN(n6253) );
  INV_X1 U7823 ( .A(n6253), .ZN(n6254) );
  INV_X2 U7824 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  OR2_X2 U7825 ( .A1(n6307), .A2(P1_U3084), .ZN(n9100) );
  INV_X1 U7826 ( .A(n6974), .ZN(n6258) );
  INV_X1 U7827 ( .A(n6259), .ZN(n6260) );
  AOI211_X1 U7828 ( .C1(n6262), .C2(n6261), .A(n7944), .B(n6260), .ZN(n6267)
         );
  NOR2_X1 U7829 ( .A1(n7938), .A2(n7828), .ZN(n6266) );
  OAI22_X1 U7830 ( .A1(n9891), .A2(n7933), .B1(n7937), .B2(n7398), .ZN(n6265)
         );
  INV_X1 U7831 ( .A(n6263), .ZN(n7403) );
  NAND2_X1 U7832 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n7144) );
  OAI21_X1 U7833 ( .B1(n7909), .B2(n7403), .A(n7144), .ZN(n6264) );
  OR4_X1 U7834 ( .A1(n6267), .A2(n6266), .A3(n6265), .A4(n6264), .ZN(P2_U3219)
         );
  INV_X1 U7835 ( .A(n7473), .ZN(n6268) );
  OR2_X1 U7836 ( .A1(n9036), .A2(n6268), .ZN(n6269) );
  NAND2_X1 U7837 ( .A1(n6269), .A2(n6307), .ZN(n6305) );
  OR2_X1 U7838 ( .A1(n6305), .A2(n6270), .ZN(n6271) );
  NAND2_X1 U7839 ( .A1(n6271), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  AND2_X1 U7840 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6942) );
  INV_X1 U7841 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6281) );
  INV_X1 U7842 ( .A(n6300), .ZN(n6570) );
  INV_X1 U7843 ( .A(n6465), .ZN(n6298) );
  NOR2_X1 U7844 ( .A1(n6296), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6277) );
  NAND2_X1 U7845 ( .A1(n6481), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6275) );
  XNOR2_X1 U7846 ( .A(n6292), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n9582) );
  INV_X1 U7847 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6272) );
  INV_X1 U7848 ( .A(n6493), .ZN(n6313) );
  OAI21_X1 U7849 ( .B1(n6272), .B2(n6313), .A(n6495), .ZN(n9581) );
  INV_X1 U7850 ( .A(n9581), .ZN(n6274) );
  INV_X1 U7851 ( .A(n6292), .ZN(n9588) );
  INV_X1 U7852 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6273) );
  OAI22_X1 U7853 ( .A1(n9582), .A2(n6274), .B1(n9588), .B2(n6273), .ZN(n6484)
         );
  OAI211_X1 U7854 ( .C1(n6481), .C2(P1_REG2_REG_3__SCAN_IN), .A(n6484), .B(
        n6275), .ZN(n6482) );
  NAND2_X1 U7855 ( .A1(n6275), .A2(n6482), .ZN(n9603) );
  INV_X1 U7856 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6276) );
  INV_X1 U7857 ( .A(n6296), .ZN(n9613) );
  AOI22_X1 U7858 ( .A1(n6296), .A2(n6276), .B1(P1_REG2_REG_4__SCAN_IN), .B2(
        n9613), .ZN(n9602) );
  NOR2_X1 U7859 ( .A1(n9603), .A2(n9602), .ZN(n9601) );
  NOR2_X1 U7860 ( .A1(n6277), .A2(n9601), .ZN(n6578) );
  INV_X1 U7861 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6278) );
  MUX2_X1 U7862 ( .A(n6278), .B(P1_REG2_REG_5__SCAN_IN), .S(n6583), .Z(n6577)
         );
  INV_X1 U7863 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6279) );
  MUX2_X1 U7864 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6279), .S(n6465), .Z(n6280)
         );
  INV_X1 U7865 ( .A(n6280), .ZN(n6469) );
  MUX2_X1 U7866 ( .A(n6281), .B(P1_REG2_REG_7__SCAN_IN), .S(n6300), .Z(n6565)
         );
  NOR2_X1 U7867 ( .A1(n6566), .A2(n6565), .ZN(n6564) );
  AOI21_X1 U7868 ( .B1(n6281), .B2(n6570), .A(n6564), .ZN(n6549) );
  INV_X1 U7869 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6548) );
  NAND2_X1 U7870 ( .A1(n6560), .A2(n6548), .ZN(n6547) );
  AOI22_X1 U7871 ( .A1(n6549), .A2(n6547), .B1(n6282), .B2(
        P1_REG2_REG_8__SCAN_IN), .ZN(n6286) );
  NAND2_X1 U7872 ( .A1(n6508), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6283) );
  OAI21_X1 U7873 ( .B1(n6508), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6283), .ZN(
        n6285) );
  NOR2_X1 U7874 ( .A1(n6286), .A2(n6285), .ZN(n6507) );
  OR2_X1 U7875 ( .A1(n9074), .A2(P1_U3084), .ZN(n7597) );
  NOR2_X1 U7876 ( .A1(n6305), .A2(n7597), .ZN(n9131) );
  INV_X1 U7877 ( .A(n9131), .ZN(n6284) );
  AOI211_X1 U7878 ( .C1(n6286), .C2(n6285), .A(n6507), .B(n9701), .ZN(n6311)
         );
  INV_X1 U7879 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6287) );
  MUX2_X1 U7880 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n6287), .S(n6300), .Z(n6569)
         );
  INV_X1 U7881 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U7882 ( .A1(n6465), .A2(n6288), .ZN(n6299) );
  NAND2_X1 U7883 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6583), .ZN(n6289) );
  OAI21_X1 U7884 ( .B1(n6583), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6289), .ZN(
        n6580) );
  NOR2_X1 U7885 ( .A1(n6296), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6290) );
  AOI21_X1 U7886 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n6296), .A(n6290), .ZN(
        n9608) );
  XNOR2_X1 U7887 ( .A(n6292), .B(n9772), .ZN(n9585) );
  INV_X1 U7888 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9770) );
  MUX2_X1 U7889 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9770), .S(n6493), .Z(n6490)
         );
  AND2_X1 U7890 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6489) );
  NAND2_X1 U7891 ( .A1(n6490), .A2(n6489), .ZN(n6488) );
  NAND2_X1 U7892 ( .A1(n6493), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6291) );
  NAND2_X1 U7893 ( .A1(n6488), .A2(n6291), .ZN(n9584) );
  NAND2_X1 U7894 ( .A1(n9585), .A2(n9584), .ZN(n9583) );
  NAND2_X1 U7895 ( .A1(n6292), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6293) );
  NAND2_X1 U7896 ( .A1(n9583), .A2(n6293), .ZN(n6475) );
  INV_X1 U7897 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6294) );
  XNOR2_X1 U7898 ( .A(n6481), .B(n6294), .ZN(n6476) );
  NAND2_X1 U7899 ( .A1(n6475), .A2(n6476), .ZN(n6474) );
  NAND2_X1 U7900 ( .A1(n6481), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6295) );
  AND2_X1 U7901 ( .A1(n6474), .A2(n6295), .ZN(n9607) );
  NAND2_X1 U7902 ( .A1(n9608), .A2(n9607), .ZN(n9606) );
  OAI21_X1 U7903 ( .B1(n6296), .B2(P1_REG1_REG_4__SCAN_IN), .A(n9606), .ZN(
        n6581) );
  NOR2_X1 U7904 ( .A1(n6580), .A2(n6581), .ZN(n6579) );
  AOI21_X1 U7905 ( .B1(n6583), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6579), .ZN(
        n6462) );
  INV_X1 U7906 ( .A(n6299), .ZN(n6297) );
  AOI21_X1 U7907 ( .B1(n6298), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6297), .ZN(
        n6463) );
  NAND2_X1 U7908 ( .A1(n6462), .A2(n6463), .ZN(n6461) );
  NAND2_X1 U7909 ( .A1(n6299), .A2(n6461), .ZN(n6568) );
  NAND2_X1 U7910 ( .A1(n6569), .A2(n6568), .ZN(n6567) );
  OR2_X1 U7911 ( .A1(n6300), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U7912 ( .A1(n6567), .A2(n6301), .ZN(n6554) );
  INV_X1 U7913 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9777) );
  OR2_X1 U7914 ( .A1(n6560), .A2(n9777), .ZN(n6553) );
  NAND2_X1 U7915 ( .A1(n6554), .A2(n6553), .ZN(n6302) );
  NAND2_X1 U7916 ( .A1(n6560), .A2(n9777), .ZN(n6551) );
  AND2_X1 U7917 ( .A1(n6302), .A2(n6551), .ZN(n6556) );
  INV_X1 U7918 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10207) );
  INV_X1 U7919 ( .A(n6508), .ZN(n6335) );
  AOI22_X1 U7920 ( .A1(n6508), .A2(n10207), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6335), .ZN(n6303) );
  NOR2_X1 U7921 ( .A1(n6556), .A2(n6303), .ZN(n6500) );
  AOI21_X1 U7922 ( .B1(n6556), .B2(n6303), .A(n6500), .ZN(n6306) );
  INV_X1 U7923 ( .A(n9074), .ZN(n9574) );
  NOR2_X1 U7924 ( .A1(n9574), .A2(n5635), .ZN(n9589) );
  NAND2_X1 U7925 ( .A1(n9589), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6304) );
  OR2_X1 U7926 ( .A1(n6305), .A2(n6304), .ZN(n9712) );
  NOR2_X1 U7927 ( .A1(n6306), .A2(n9712), .ZN(n6310) );
  INV_X1 U7928 ( .A(P1_U3083), .ZN(n6308) );
  INV_X1 U7929 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10342) );
  OAI22_X1 U7930 ( .A1(n9716), .A2(n10342), .B1(n9691), .B2(n6335), .ZN(n6309)
         );
  OR4_X1 U7931 ( .A1(n6942), .A2(n6311), .A3(n6310), .A4(n6309), .ZN(P1_U3250)
         );
  XNOR2_X1 U7932 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AND2_X1 U7933 ( .A1(n7727), .A2(P2_U3152), .ZN(n8658) );
  INV_X2 U7934 ( .A(n8658), .ZN(n8657) );
  NOR2_X1 U7935 ( .A1(n7727), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8654) );
  AOI22_X1 U7936 ( .A1(n8654), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n9482), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6312) );
  OAI21_X1 U7937 ( .B1(n6316), .B2(n8657), .A(n6312), .ZN(P2_U3356) );
  INV_X1 U7938 ( .A(n4461), .ZN(n6956) );
  OAI222_X1 U7939 ( .A1(n8661), .A2(n10091), .B1(n8657), .B2(n6314), .C1(
        P2_U3152), .C2(n6956), .ZN(P2_U3357) );
  AND2_X1 U7940 ( .A1(n7727), .A2(P1_U3084), .ZN(n9463) );
  INV_X1 U7941 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6315) );
  OAI222_X1 U7942 ( .A1(n7760), .A2(n6315), .B1(n9460), .B2(n6314), .C1(n6313), 
        .C2(P1_U3084), .ZN(P1_U3352) );
  OAI222_X1 U7943 ( .A1(n7760), .A2(n6317), .B1(n9460), .B2(n6316), .C1(n9588), 
        .C2(P1_U3084), .ZN(P1_U3351) );
  INV_X1 U7944 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10229) );
  INV_X1 U7945 ( .A(n6481), .ZN(n6479) );
  OAI222_X1 U7946 ( .A1(n7760), .A2(n10229), .B1(n9460), .B2(n6318), .C1(n6479), .C2(P1_U3084), .ZN(P1_U3350) );
  INV_X1 U7947 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6319) );
  INV_X1 U7948 ( .A(n6981), .ZN(n7113) );
  OAI222_X1 U7949 ( .A1(n8661), .A2(n6319), .B1(n8657), .B2(n6318), .C1(
        P2_U3152), .C2(n7113), .ZN(P2_U3355) );
  INV_X1 U7950 ( .A(n6982), .ZN(n7126) );
  OAI222_X1 U7951 ( .A1(n8661), .A2(n6320), .B1(n8657), .B2(n6321), .C1(
        P2_U3152), .C2(n7126), .ZN(P2_U3354) );
  OAI222_X1 U7952 ( .A1(n9613), .A2(P1_U3084), .B1(n9460), .B2(n6321), .C1(
        n10226), .C2(n7760), .ZN(P1_U3349) );
  AOI22_X1 U7953 ( .A1(n6583), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9463), .ZN(n6322) );
  OAI21_X1 U7954 ( .B1(n6323), .B2(n9460), .A(n6322), .ZN(P1_U3348) );
  INV_X1 U7955 ( .A(n6984), .ZN(n7138) );
  OAI222_X1 U7956 ( .A1(n8661), .A2(n6324), .B1(n8657), .B2(n6323), .C1(
        P2_U3152), .C2(n7138), .ZN(P2_U3353) );
  INV_X1 U7957 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6325) );
  INV_X1 U7958 ( .A(n6986), .ZN(n7101) );
  OAI222_X1 U7959 ( .A1(n8661), .A2(n6325), .B1(n8657), .B2(n6326), .C1(
        P2_U3152), .C2(n7101), .ZN(P2_U3352) );
  INV_X1 U7960 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6327) );
  OAI222_X1 U7961 ( .A1(n7760), .A2(n6327), .B1(n9460), .B2(n6326), .C1(n6465), 
        .C2(P1_U3084), .ZN(P1_U3347) );
  OAI222_X1 U7962 ( .A1(n7760), .A2(n10185), .B1(n9460), .B2(n6328), .C1(n6570), .C2(P1_U3084), .ZN(P1_U3346) );
  INV_X1 U7963 ( .A(n6989), .ZN(n7166) );
  OAI222_X1 U7964 ( .A1(n8661), .A2(n6329), .B1(n8657), .B2(n6328), .C1(
        P2_U3152), .C2(n7166), .ZN(P2_U3351) );
  INV_X1 U7965 ( .A(n6991), .ZN(n7178) );
  OAI222_X1 U7966 ( .A1(n8661), .A2(n6330), .B1(n8657), .B2(n6331), .C1(
        P2_U3152), .C2(n7178), .ZN(P2_U3350) );
  OAI222_X1 U7967 ( .A1(n7760), .A2(n6332), .B1(n9460), .B2(n6331), .C1(n6560), 
        .C2(P1_U3084), .ZN(P1_U3345) );
  INV_X1 U7968 ( .A(n6333), .ZN(n6336) );
  OAI222_X1 U7969 ( .A1(P1_U3084), .A2(n6335), .B1(n9460), .B2(n6336), .C1(
        n6334), .C2(n7760), .ZN(P1_U3344) );
  OAI222_X1 U7970 ( .A1(n8661), .A2(n6337), .B1(n8657), .B2(n6336), .C1(n7190), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U7971 ( .A(n6338), .ZN(n6343) );
  AOI22_X1 U7972 ( .A1(n8183), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n8654), .ZN(n6339) );
  OAI21_X1 U7973 ( .B1(n6343), .B2(n8657), .A(n6339), .ZN(P2_U3347) );
  INV_X1 U7974 ( .A(n6510), .ZN(n6816) );
  INV_X1 U7975 ( .A(n6340), .ZN(n6342) );
  OAI222_X1 U7976 ( .A1(P1_U3084), .A2(n6816), .B1(n9460), .B2(n6342), .C1(
        n6341), .C2(n7760), .ZN(P1_U3343) );
  INV_X1 U7977 ( .A(n7146), .ZN(n7154) );
  OAI222_X1 U7978 ( .A1(n8661), .A2(n10246), .B1(n8657), .B2(n6342), .C1(n7154), .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U7979 ( .A(n9103), .ZN(n9118) );
  OAI222_X1 U7980 ( .A1(n7760), .A2(n6344), .B1(n9460), .B2(n6343), .C1(
        P1_U3084), .C2(n9118), .ZN(P1_U3342) );
  INV_X1 U7981 ( .A(n6345), .ZN(n6346) );
  OAI222_X1 U7982 ( .A1(n7760), .A2(n10266), .B1(n9460), .B2(n6346), .C1(n9119), .C2(P1_U3084), .ZN(P1_U3341) );
  INV_X1 U7983 ( .A(n7062), .ZN(n6969) );
  OAI222_X1 U7984 ( .A1(n8661), .A2(n6347), .B1(n8657), .B2(n6346), .C1(
        P2_U3152), .C2(n6969), .ZN(P2_U3346) );
  INV_X1 U7985 ( .A(n6348), .ZN(n6350) );
  AOI22_X1 U7986 ( .A1(n9638), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9463), .ZN(n6349) );
  OAI21_X1 U7987 ( .B1(n6350), .B2(n9460), .A(n6349), .ZN(P1_U3340) );
  INV_X1 U7988 ( .A(n7029), .ZN(n7024) );
  OAI222_X1 U7989 ( .A1(n8661), .A2(n6351), .B1(n8657), .B2(n6350), .C1(n7024), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  OR2_X1 U7990 ( .A1(n6352), .A2(P2_U3152), .ZN(n8162) );
  NAND2_X1 U7991 ( .A1(n9844), .A2(n8162), .ZN(n6353) );
  NAND2_X1 U7992 ( .A1(n6353), .A2(n4467), .ZN(n6355) );
  OR2_X1 U7993 ( .A1(n9844), .A2(n6634), .ZN(n6354) );
  NOR2_X1 U7994 ( .A1(n9788), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7995 ( .A(n6356), .ZN(n6357) );
  INV_X1 U7996 ( .A(n8192), .ZN(n8199) );
  OAI222_X1 U7997 ( .A1(n8661), .A2(n10095), .B1(n8657), .B2(n6357), .C1(n8199), .C2(P2_U3152), .ZN(P2_U3344) );
  OAI222_X1 U7998 ( .A1(P1_U3084), .A2(n9653), .B1(n9460), .B2(n6357), .C1(
        n10102), .C2(n7760), .ZN(P1_U3339) );
  NAND2_X1 U7999 ( .A1(n7693), .A2(n9102), .ZN(n6362) );
  INV_X1 U8000 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6494) );
  NOR2_X1 U8001 ( .A1(n6382), .A2(n6494), .ZN(n6360) );
  AOI21_X1 U8002 ( .B1(n6407), .B2(n6597), .A(n6360), .ZN(n6361) );
  NAND2_X1 U8003 ( .A1(n6363), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6364) );
  NAND2_X1 U8004 ( .A1(n6366), .A2(n6394), .ZN(n6397) );
  OAI21_X1 U8005 ( .B1(n6366), .B2(n6394), .A(n6397), .ZN(n9595) );
  INV_X1 U8006 ( .A(n9595), .ZN(n6381) );
  AND2_X1 U8007 ( .A1(n9450), .A2(n6367), .ZN(n6432) );
  NAND2_X1 U8008 ( .A1(n6432), .A2(n6520), .ZN(n6372) );
  INV_X1 U8009 ( .A(n6372), .ZN(n6371) );
  AND2_X1 U8010 ( .A1(n6371), .A2(n9722), .ZN(n6375) );
  INV_X1 U8011 ( .A(n6375), .ZN(n6376) );
  INV_X1 U8012 ( .A(n9036), .ZN(n6368) );
  INV_X1 U8013 ( .A(n6369), .ZN(n6373) );
  OR2_X1 U8014 ( .A1(n6536), .A2(n5670), .ZN(n6538) );
  INV_X1 U8015 ( .A(n9722), .ZN(n6370) );
  OR3_X1 U8016 ( .A1(n6538), .A2(n6371), .A3(n6370), .ZN(n6385) );
  NAND2_X1 U8017 ( .A1(n9760), .A2(n6372), .ZN(n6383) );
  NAND3_X1 U8018 ( .A1(n6373), .A2(n6385), .A3(n6383), .ZN(n8768) );
  INV_X1 U8019 ( .A(n6390), .ZN(n6374) );
  AND2_X1 U8020 ( .A1(n6374), .A2(n6524), .ZN(n9075) );
  AND2_X1 U8021 ( .A1(n6375), .A2(n9075), .ZN(n6420) );
  OR2_X1 U8022 ( .A1(n6376), .A2(n6538), .ZN(n6378) );
  NAND2_X1 U8023 ( .A1(n9722), .A2(n5062), .ZN(n6377) );
  OAI22_X1 U8024 ( .A1(n8805), .A2(n5644), .B1(n8750), .B2(n6614), .ZN(n6379)
         );
  AOI21_X1 U8025 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n8768), .A(n6379), .ZN(
        n6380) );
  OAI21_X1 U8026 ( .B1(n6381), .B2(n8782), .A(n6380), .ZN(P1_U3230) );
  NAND4_X1 U8027 ( .A1(n6383), .A2(n6382), .A3(n7473), .A4(n6522), .ZN(n6384)
         );
  NAND2_X1 U8028 ( .A1(n6384), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6386) );
  INV_X1 U8029 ( .A(n8802), .ZN(n8792) );
  NAND2_X1 U8030 ( .A1(n6407), .A2(n9098), .ZN(n6389) );
  NAND2_X1 U8031 ( .A1(n6587), .A2(n7695), .ZN(n6388) );
  NAND2_X1 U8032 ( .A1(n6389), .A2(n6388), .ZN(n6391) );
  XNOR2_X1 U8033 ( .A(n6391), .B(n7696), .ZN(n6440) );
  NAND2_X1 U8034 ( .A1(n7693), .A2(n9098), .ZN(n6393) );
  NAND2_X1 U8035 ( .A1(n6407), .A2(n6587), .ZN(n6392) );
  AND2_X1 U8036 ( .A1(n6393), .A2(n6392), .ZN(n6441) );
  XNOR2_X1 U8037 ( .A(n6440), .B(n6441), .ZN(n6418) );
  INV_X1 U8038 ( .A(n6394), .ZN(n6395) );
  NAND2_X1 U8039 ( .A1(n6395), .A2(n7696), .ZN(n6396) );
  AND2_X1 U8040 ( .A1(n6397), .A2(n6396), .ZN(n6402) );
  NAND2_X1 U8041 ( .A1(n6407), .A2(n9101), .ZN(n6399) );
  NAND2_X1 U8042 ( .A1(n9042), .A2(n7695), .ZN(n6398) );
  NAND2_X1 U8043 ( .A1(n6399), .A2(n6398), .ZN(n6400) );
  XNOR2_X1 U8044 ( .A(n6400), .B(n7696), .ZN(n6403) );
  NAND2_X1 U8045 ( .A1(n6402), .A2(n6403), .ZN(n6425) );
  AOI22_X1 U8046 ( .A1(n7693), .A2(n9101), .B1(n7694), .B2(n9042), .ZN(n6427)
         );
  NAND2_X1 U8047 ( .A1(n6425), .A2(n6427), .ZN(n6406) );
  INV_X1 U8048 ( .A(n6402), .ZN(n6405) );
  INV_X1 U8049 ( .A(n6403), .ZN(n6404) );
  NAND2_X1 U8050 ( .A1(n6405), .A2(n6404), .ZN(n6426) );
  NAND2_X1 U8051 ( .A1(n6406), .A2(n6426), .ZN(n8763) );
  NAND2_X1 U8052 ( .A1(n9099), .A2(n6407), .ZN(n6409) );
  NAND2_X1 U8053 ( .A1(n8767), .A2(n6387), .ZN(n6408) );
  NAND2_X1 U8054 ( .A1(n6409), .A2(n6408), .ZN(n6410) );
  XNOR2_X1 U8055 ( .A(n6410), .B(n7616), .ZN(n6411) );
  AOI22_X1 U8056 ( .A1(n7693), .A2(n9099), .B1(n6407), .B2(n8767), .ZN(n6412)
         );
  NAND2_X1 U8057 ( .A1(n6411), .A2(n6412), .ZN(n6416) );
  INV_X1 U8058 ( .A(n6411), .ZN(n6414) );
  INV_X1 U8059 ( .A(n6412), .ZN(n6413) );
  NAND2_X1 U8060 ( .A1(n6414), .A2(n6413), .ZN(n6415) );
  NAND2_X1 U8061 ( .A1(n8763), .A2(n8764), .ZN(n8762) );
  NAND2_X1 U8062 ( .A1(n8762), .A2(n6416), .ZN(n6417) );
  OAI21_X1 U8063 ( .B1(n6418), .B2(n6417), .A(n6450), .ZN(n6419) );
  NAND2_X1 U8064 ( .A1(n6419), .A2(n8765), .ZN(n6424) );
  AND2_X1 U8065 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6473) );
  INV_X1 U8066 ( .A(n6420), .ZN(n6421) );
  OAI22_X1 U8067 ( .A1(n6539), .A2(n8750), .B1(n8778), .B2(n6608), .ZN(n6422)
         );
  AOI211_X1 U8068 ( .C1(n8789), .C2(n9097), .A(n6473), .B(n6422), .ZN(n6423)
         );
  OAI211_X1 U8069 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n8792), .A(n6424), .B(
        n6423), .ZN(P1_U3216) );
  NAND2_X1 U8070 ( .A1(n6425), .A2(n6426), .ZN(n6428) );
  XNOR2_X1 U8071 ( .A(n6428), .B(n6427), .ZN(n6431) );
  AOI22_X1 U8072 ( .A1(n8801), .A2(n9102), .B1(n8789), .B2(n9099), .ZN(n6430)
         );
  AOI22_X1 U8073 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(n8768), .B1(n8807), .B2(
        n9042), .ZN(n6429) );
  OAI211_X1 U8074 ( .C1(n6431), .C2(n8782), .A(n6430), .B(n6429), .ZN(P1_U3220) );
  INV_X2 U8075 ( .A(n9779), .ZN(n9781) );
  INV_X1 U8076 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9578) );
  AND2_X1 U8077 ( .A1(n6614), .A2(n9102), .ZN(n9040) );
  NOR2_X1 U8078 ( .A1(n9040), .A2(n6606), .ZN(n8883) );
  INV_X1 U8079 ( .A(n6536), .ZN(n6435) );
  NOR3_X1 U8080 ( .A1(n8883), .A2(n9075), .A3(n6435), .ZN(n6436) );
  AOI21_X1 U8081 ( .B1(n9319), .B2(n9101), .A(n6436), .ZN(n6600) );
  OAI21_X1 U8082 ( .B1(n6614), .B2(n6536), .A(n6600), .ZN(n6438) );
  NAND2_X1 U8083 ( .A1(n6438), .A2(n9781), .ZN(n6437) );
  OAI21_X1 U8084 ( .B1(n9781), .B2(n9578), .A(n6437), .ZN(P1_U3523) );
  NAND2_X1 U8085 ( .A1(n6438), .A2(n9759), .ZN(n6439) );
  OAI21_X1 U8086 ( .B1(n9759), .B2(n5403), .A(n6439), .ZN(P1_U3454) );
  INV_X1 U8087 ( .A(n6748), .ZN(n6456) );
  INV_X1 U8088 ( .A(n6440), .ZN(n6442) );
  NAND2_X1 U8089 ( .A1(n6442), .A2(n6441), .ZN(n6448) );
  AND2_X1 U8090 ( .A1(n6450), .A2(n6448), .ZN(n6452) );
  NAND2_X1 U8091 ( .A1(n6407), .A2(n9097), .ZN(n6444) );
  NAND2_X1 U8092 ( .A1(n6747), .A2(n7695), .ZN(n6443) );
  NAND2_X1 U8093 ( .A1(n6444), .A2(n6443), .ZN(n6445) );
  XNOR2_X1 U8094 ( .A(n6445), .B(n7696), .ZN(n6651) );
  NAND2_X1 U8095 ( .A1(n7693), .A2(n9097), .ZN(n6447) );
  NAND2_X1 U8096 ( .A1(n6407), .A2(n6747), .ZN(n6446) );
  AND2_X1 U8097 ( .A1(n6447), .A2(n6446), .ZN(n6649) );
  XNOR2_X1 U8098 ( .A(n6651), .B(n6649), .ZN(n6451) );
  AND2_X1 U8099 ( .A1(n6451), .A2(n6448), .ZN(n6449) );
  OAI211_X1 U8100 ( .C1(n6452), .C2(n6451), .A(n8765), .B(n6653), .ZN(n6455)
         );
  AND2_X1 U8101 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9609) );
  OAI22_X1 U8102 ( .A1(n8805), .A2(n6907), .B1(n9736), .B2(n8750), .ZN(n6453)
         );
  AOI211_X1 U8103 ( .C1(n8801), .C2(n9098), .A(n9609), .B(n6453), .ZN(n6454)
         );
  OAI211_X1 U8104 ( .C1(n8792), .C2(n6456), .A(n6455), .B(n6454), .ZN(P1_U3228) );
  INV_X1 U8105 ( .A(n6457), .ZN(n6460) );
  INV_X1 U8106 ( .A(n8206), .ZN(n8215) );
  OAI222_X1 U8107 ( .A1(n8661), .A2(n6458), .B1(n8657), .B2(n6460), .C1(
        P2_U3152), .C2(n8215), .ZN(P2_U3343) );
  INV_X1 U8108 ( .A(n9667), .ZN(n9122) );
  OAI222_X1 U8109 ( .A1(n9122), .A2(P1_U3084), .B1(n9460), .B2(n6460), .C1(
        n6459), .C2(n7760), .ZN(P1_U3338) );
  INV_X1 U8110 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6472) );
  OAI21_X1 U8111 ( .B1(n6463), .B2(n6462), .A(n6461), .ZN(n6467) );
  NOR2_X1 U8112 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6464), .ZN(n6783) );
  NOR2_X1 U8113 ( .A1(n9691), .A2(n6465), .ZN(n6466) );
  AOI211_X1 U8114 ( .C1(n9693), .C2(n6467), .A(n6783), .B(n6466), .ZN(n6471)
         );
  OAI211_X1 U8115 ( .C1(n4566), .C2(n6469), .A(n9687), .B(n6468), .ZN(n6470)
         );
  OAI211_X1 U8116 ( .C1(n6472), .C2(n9716), .A(n6471), .B(n6470), .ZN(P1_U3247) );
  INV_X1 U8117 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6487) );
  INV_X1 U8118 ( .A(n6473), .ZN(n6478) );
  OAI211_X1 U8119 ( .C1(n6476), .C2(n6475), .A(n9693), .B(n6474), .ZN(n6477)
         );
  OAI211_X1 U8120 ( .C1(n9691), .C2(n6479), .A(n6478), .B(n6477), .ZN(n6480)
         );
  INV_X1 U8121 ( .A(n6480), .ZN(n6486) );
  INV_X1 U8122 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6533) );
  MUX2_X1 U8123 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6533), .S(n6481), .Z(n6483)
         );
  OAI211_X1 U8124 ( .C1(n6484), .C2(n6483), .A(n9687), .B(n6482), .ZN(n6485)
         );
  OAI211_X1 U8125 ( .C1(n6487), .C2(n9716), .A(n6486), .B(n6485), .ZN(P1_U3244) );
  INV_X1 U8126 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6499) );
  INV_X1 U8127 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6615) );
  OAI211_X1 U8128 ( .C1(n6490), .C2(n6489), .A(n9693), .B(n6488), .ZN(n6491)
         );
  OAI21_X1 U8129 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6615), .A(n6491), .ZN(n6492) );
  AOI21_X1 U8130 ( .B1(n6493), .B2(n9707), .A(n6492), .ZN(n6498) );
  INV_X1 U8131 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6596) );
  NOR2_X1 U8132 ( .A1(n6494), .A2(n6596), .ZN(n9591) );
  OAI211_X1 U8133 ( .C1(n9591), .C2(n6496), .A(n9687), .B(n6495), .ZN(n6497)
         );
  OAI211_X1 U8134 ( .C1(n6499), .C2(n9716), .A(n6498), .B(n6497), .ZN(P1_U3242) );
  NOR2_X1 U8135 ( .A1(n6508), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6501) );
  NOR2_X1 U8136 ( .A1(n6501), .A2(n6500), .ZN(n6815) );
  INV_X1 U8137 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9527) );
  AOI22_X1 U8138 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n6816), .B1(n6510), .B2(
        n9527), .ZN(n6814) );
  NOR2_X1 U8139 ( .A1(n6815), .A2(n6814), .ZN(n6813) );
  NOR2_X1 U8140 ( .A1(n6510), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6502) );
  NOR2_X1 U8141 ( .A1(n6813), .A2(n6502), .ZN(n6505) );
  INV_X1 U8142 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6503) );
  MUX2_X1 U8143 ( .A(n6503), .B(P1_REG1_REG_11__SCAN_IN), .S(n9103), .Z(n6504)
         );
  NOR2_X1 U8144 ( .A1(n6505), .A2(n6504), .ZN(n9117) );
  AOI21_X1 U8145 ( .B1(n6505), .B2(n6504), .A(n9117), .ZN(n6517) );
  INV_X1 U8146 ( .A(n9716), .ZN(n6822) );
  NOR2_X1 U8147 ( .A1(n9103), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6506) );
  AOI21_X1 U8148 ( .B1(n9103), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6506), .ZN(
        n6512) );
  AOI21_X1 U8149 ( .B1(n6508), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6507), .ZN(
        n6819) );
  NAND2_X1 U8150 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n6510), .ZN(n6509) );
  OAI21_X1 U8151 ( .B1(n6510), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6509), .ZN(
        n6818) );
  OAI21_X1 U8152 ( .B1(n6512), .B2(n6511), .A(n9104), .ZN(n6513) );
  NAND2_X1 U8153 ( .A1(n9687), .A2(n6513), .ZN(n6514) );
  NAND2_X1 U8154 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7238) );
  OAI211_X1 U8155 ( .C1(n9691), .C2(n9118), .A(n6514), .B(n7238), .ZN(n6515)
         );
  AOI21_X1 U8156 ( .B1(n6822), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n6515), .ZN(
        n6516) );
  OAI21_X1 U8157 ( .B1(n6517), .B2(n9712), .A(n6516), .ZN(P1_U3252) );
  OAI21_X1 U8158 ( .B1(n6519), .B2(n6526), .A(n6518), .ZN(n6532) );
  INV_X1 U8159 ( .A(n6532), .ZN(n6591) );
  NAND2_X1 U8160 ( .A1(n9722), .A2(n6520), .ZN(n9720) );
  NOR2_X1 U8161 ( .A1(n6521), .A2(n9720), .ZN(n6523) );
  NAND2_X1 U8162 ( .A1(n6523), .A2(n6522), .ZN(n6758) );
  INV_X2 U8163 ( .A(n9338), .ZN(n9519) );
  NAND2_X1 U8164 ( .A1(n6524), .A2(n9257), .ZN(n6525) );
  OR2_X1 U8165 ( .A1(n9519), .A2(n6525), .ZN(n9358) );
  OAI22_X1 U8166 ( .A1(n6732), .A2(n9501), .B1(n9502), .B2(n6608), .ZN(n6531)
         );
  INV_X1 U8167 ( .A(n8860), .ZN(n6527) );
  NAND2_X1 U8168 ( .A1(n6527), .A2(n6526), .ZN(n6529) );
  AOI21_X1 U8169 ( .B1(n6529), .B2(n6528), .A(n9497), .ZN(n6530) );
  AOI211_X1 U8170 ( .C1(n9506), .C2(n6532), .A(n6531), .B(n6530), .ZN(n6590)
         );
  MUX2_X1 U8171 ( .A(n6533), .B(n6590), .S(n9338), .Z(n6542) );
  INV_X1 U8172 ( .A(n6745), .ZN(n6534) );
  AOI21_X1 U8173 ( .B1(n6587), .B2(n9729), .A(n6534), .ZN(n6588) );
  INV_X1 U8174 ( .A(n6535), .ZN(n9072) );
  OR2_X1 U8175 ( .A1(n6536), .A2(n9072), .ZN(n6537) );
  OAI22_X1 U8176 ( .A1(n9357), .A2(n6539), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9294), .ZN(n6540) );
  AOI21_X1 U8177 ( .B1(n6588), .B2(n9361), .A(n6540), .ZN(n6541) );
  OAI211_X1 U8178 ( .C1(n6591), .C2(n9358), .A(n6542), .B(n6541), .ZN(P1_U3288) );
  INV_X1 U8179 ( .A(n6543), .ZN(n6546) );
  AOI22_X1 U8180 ( .A1(n9676), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9463), .ZN(n6544) );
  OAI21_X1 U8181 ( .B1(n6546), .B2(n9460), .A(n6544), .ZN(P1_U3337) );
  AOI22_X1 U8182 ( .A1(n8232), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n8654), .ZN(n6545) );
  OAI21_X1 U8183 ( .B1(n6546), .B2(n8657), .A(n6545), .ZN(P2_U3342) );
  OAI21_X1 U8184 ( .B1(n6548), .B2(n6560), .A(n6547), .ZN(n6550) );
  XOR2_X1 U8185 ( .A(n6550), .B(n6549), .Z(n6563) );
  INV_X1 U8186 ( .A(n6551), .ZN(n6552) );
  AND2_X1 U8187 ( .A1(n6554), .A2(n6552), .ZN(n6555) );
  OAI22_X1 U8188 ( .A1(n6556), .A2(n6555), .B1(n6554), .B2(n6553), .ZN(n6558)
         );
  NOR2_X1 U8189 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6557), .ZN(n7014) );
  AOI21_X1 U8190 ( .B1(n9693), .B2(n6558), .A(n7014), .ZN(n6559) );
  OAI21_X1 U8191 ( .B1(n9691), .B2(n6560), .A(n6559), .ZN(n6561) );
  AOI21_X1 U8192 ( .B1(n6822), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n6561), .ZN(
        n6562) );
  OAI21_X1 U8193 ( .B1(n6563), .B2(n9701), .A(n6562), .ZN(P1_U3249) );
  AOI21_X1 U8194 ( .B1(n6566), .B2(n6565), .A(n6564), .ZN(n6575) );
  OAI21_X1 U8195 ( .B1(n6569), .B2(n6568), .A(n6567), .ZN(n6572) );
  AND2_X1 U8196 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6685) );
  NOR2_X1 U8197 ( .A1(n9691), .A2(n6570), .ZN(n6571) );
  AOI211_X1 U8198 ( .C1(n9693), .C2(n6572), .A(n6685), .B(n6571), .ZN(n6574)
         );
  NAND2_X1 U8199 ( .A1(n6822), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n6573) );
  OAI211_X1 U8200 ( .C1(n6575), .C2(n9701), .A(n6574), .B(n6573), .ZN(P1_U3248) );
  AOI21_X1 U8201 ( .B1(n6578), .B2(n6577), .A(n6576), .ZN(n6586) );
  AND2_X1 U8202 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6734) );
  AOI211_X1 U8203 ( .C1(n6581), .C2(n6580), .A(n6579), .B(n9712), .ZN(n6582)
         );
  AOI211_X1 U8204 ( .C1(n9707), .C2(n6583), .A(n6734), .B(n6582), .ZN(n6585)
         );
  NAND2_X1 U8205 ( .A1(n6822), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n6584) );
  OAI211_X1 U8206 ( .C1(n6586), .C2(n9701), .A(n6585), .B(n6584), .ZN(P1_U3246) );
  INV_X1 U8207 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6593) );
  AOI22_X1 U8208 ( .A1(n6588), .A2(n9751), .B1(n9750), .B2(n6587), .ZN(n6589)
         );
  OAI211_X1 U8209 ( .C1(n6591), .C2(n9756), .A(n6590), .B(n6589), .ZN(n6594)
         );
  NAND2_X1 U8210 ( .A1(n6594), .A2(n9759), .ZN(n6592) );
  OAI21_X1 U8211 ( .B1(n9759), .B2(n6593), .A(n6592), .ZN(P1_U3463) );
  NAND2_X1 U8212 ( .A1(n6594), .A2(n9781), .ZN(n6595) );
  OAI21_X1 U8213 ( .B1(n9781), .B2(n6294), .A(n6595), .ZN(P1_U3526) );
  AOI22_X1 U8214 ( .A1(n9312), .A2(P1_REG2_REG_0__SCAN_IN), .B1(n9508), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n6599) );
  OAI21_X1 U8215 ( .B1(n9361), .B2(n9509), .A(n6597), .ZN(n6598) );
  OAI211_X1 U8216 ( .C1(n6600), .C2(n9519), .A(n6599), .B(n6598), .ZN(P1_U3291) );
  INV_X1 U8217 ( .A(n6601), .ZN(n6709) );
  AOI22_X1 U8218 ( .A1(n9116), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9463), .ZN(n6602) );
  OAI21_X1 U8219 ( .B1(n6709), .B2(n9460), .A(n6602), .ZN(P1_U3336) );
  OAI21_X1 U8220 ( .B1(n8884), .B2(n6604), .A(n6603), .ZN(n9723) );
  OAI21_X1 U8221 ( .B1(n6607), .B2(n6606), .A(n6605), .ZN(n6611) );
  OAI22_X1 U8222 ( .A1(n6609), .A2(n9502), .B1(n9501), .B2(n6608), .ZN(n6610)
         );
  AOI21_X1 U8223 ( .B1(n6611), .B2(n9351), .A(n6610), .ZN(n6612) );
  OAI21_X1 U8224 ( .B1(n9347), .B2(n9723), .A(n6612), .ZN(n9726) );
  INV_X1 U8225 ( .A(n9042), .ZN(n9725) );
  INV_X1 U8226 ( .A(n6613), .ZN(n6698) );
  OAI211_X1 U8227 ( .C1(n9725), .C2(n6614), .A(n6698), .B(n9751), .ZN(n9724)
         );
  OAI22_X1 U8228 ( .A1(n9724), .A2(n9257), .B1(n9294), .B2(n6615), .ZN(n6616)
         );
  OAI21_X1 U8229 ( .B1(n9726), .B2(n6616), .A(n9338), .ZN(n6618) );
  AOI22_X1 U8230 ( .A1(n9509), .A2(n9042), .B1(n9519), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n6617) );
  OAI211_X1 U8231 ( .C1(n9723), .C2(n9358), .A(n6618), .B(n6617), .ZN(P1_U3290) );
  NAND2_X1 U8232 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n8176), .ZN(n6619) );
  OAI21_X1 U8233 ( .B1(n8492), .B2(n8176), .A(n6619), .ZN(P2_U3570) );
  NOR2_X1 U8234 ( .A1(n9844), .A2(n6620), .ZN(n6768) );
  NAND2_X1 U8235 ( .A1(n6621), .A2(n6768), .ZN(n7250) );
  NOR2_X1 U8236 ( .A1(n7250), .A2(n6622), .ZN(n6624) );
  INV_X1 U8237 ( .A(n7252), .ZN(n6623) );
  INV_X1 U8238 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6648) );
  INV_X1 U8239 ( .A(n6807), .ZN(n6626) );
  NAND2_X1 U8240 ( .A1(n6807), .A2(n6627), .ZN(n7993) );
  NAND2_X1 U8241 ( .A1(n8124), .A2(n7993), .ZN(n6786) );
  NAND2_X1 U8242 ( .A1(n6786), .A2(n6788), .ZN(n6787) );
  NAND2_X1 U8243 ( .A1(n6787), .A2(n6626), .ZN(n6630) );
  NAND2_X1 U8244 ( .A1(n6628), .A2(n7312), .ZN(n6629) );
  NAND2_X1 U8245 ( .A1(n6630), .A2(n6629), .ZN(n6800) );
  INV_X1 U8246 ( .A(n6794), .ZN(n8175) );
  NAND2_X1 U8247 ( .A1(n6794), .A2(n7302), .ZN(n7994) );
  AND2_X2 U8248 ( .A1(n7984), .A2(n7994), .ZN(n8119) );
  NAND2_X1 U8249 ( .A1(n6794), .A2(n6803), .ZN(n6631) );
  INV_X1 U8250 ( .A(n6806), .ZN(n8174) );
  INV_X1 U8251 ( .A(n6892), .ZN(n9826) );
  NAND2_X1 U8252 ( .A1(n8174), .A2(n9826), .ZN(n7998) );
  NAND2_X1 U8253 ( .A1(n6806), .A2(n6892), .ZN(n7979) );
  NAND2_X1 U8254 ( .A1(n7998), .A2(n7979), .ZN(n8126) );
  NAND2_X1 U8255 ( .A1(n6632), .A2(n8126), .ZN(n6712) );
  OR2_X1 U8256 ( .A1(n6632), .A2(n8126), .ZN(n6633) );
  NAND2_X1 U8257 ( .A1(n6712), .A2(n6633), .ZN(n9820) );
  INV_X1 U8258 ( .A(n9820), .ZN(n6646) );
  AND2_X1 U8259 ( .A1(n6634), .A2(n8149), .ZN(n6636) );
  NAND2_X1 U8260 ( .A1(n7265), .A2(n7785), .ZN(n6635) );
  NAND2_X1 U8261 ( .A1(n6636), .A2(n6635), .ZN(n7402) );
  INV_X1 U8262 ( .A(n7402), .ZN(n9810) );
  OR2_X1 U8263 ( .A1(n7262), .A2(n8491), .ZN(n6638) );
  OR2_X1 U8264 ( .A1(n6794), .A2(n8474), .ZN(n6637) );
  NAND2_X1 U8265 ( .A1(n6638), .A2(n6637), .ZN(n6890) );
  INV_X1 U8266 ( .A(n7994), .ZN(n6640) );
  INV_X1 U8267 ( .A(n8126), .ZN(n7988) );
  XNOR2_X1 U8268 ( .A(n6714), .B(n7988), .ZN(n6641) );
  NAND2_X1 U8269 ( .A1(n8152), .A2(n5748), .ZN(n7965) );
  NOR2_X1 U8270 ( .A1(n6641), .A2(n9813), .ZN(n6642) );
  AOI211_X1 U8271 ( .C1(n9810), .C2(n9820), .A(n6890), .B(n6642), .ZN(n9830)
         );
  INV_X1 U8272 ( .A(n6231), .ZN(n6643) );
  AOI21_X1 U8273 ( .B1(n6801), .B2(n6892), .A(n9907), .ZN(n6644) );
  AND2_X1 U8274 ( .A1(n6644), .A2(n6719), .ZN(n9822) );
  AOI21_X1 U8275 ( .B1(n8624), .B2(n6892), .A(n9822), .ZN(n6645) );
  OAI211_X1 U8276 ( .C1(n6646), .C2(n9878), .A(n9830), .B(n6645), .ZN(n6706)
         );
  NAND2_X1 U8277 ( .A1(n6706), .A2(n9927), .ZN(n6647) );
  OAI21_X1 U8278 ( .B1(n9927), .B2(n6648), .A(n6647), .ZN(P2_U3523) );
  INV_X1 U8279 ( .A(n6649), .ZN(n6650) );
  NAND2_X1 U8280 ( .A1(n6651), .A2(n6650), .ZN(n6652) );
  NAND2_X1 U8281 ( .A1(n7694), .A2(n9096), .ZN(n6655) );
  NAND2_X1 U8282 ( .A1(n6879), .A2(n7680), .ZN(n6654) );
  NAND2_X1 U8283 ( .A1(n6655), .A2(n6654), .ZN(n6656) );
  XNOR2_X1 U8284 ( .A(n6656), .B(n7616), .ZN(n6729) );
  NAND2_X1 U8285 ( .A1(n7693), .A2(n9096), .ZN(n6658) );
  NAND2_X1 U8286 ( .A1(n7694), .A2(n6879), .ZN(n6657) );
  AND2_X1 U8287 ( .A1(n6658), .A2(n6657), .ZN(n6665) );
  NAND2_X1 U8288 ( .A1(n6729), .A2(n6665), .ZN(n6659) );
  NAND2_X1 U8289 ( .A1(n6407), .A2(n9095), .ZN(n6661) );
  NAND2_X1 U8290 ( .A1(n9742), .A2(n7680), .ZN(n6660) );
  NAND2_X1 U8291 ( .A1(n6661), .A2(n6660), .ZN(n6662) );
  XNOR2_X1 U8292 ( .A(n6662), .B(n7696), .ZN(n6670) );
  NAND2_X1 U8293 ( .A1(n7693), .A2(n9095), .ZN(n6664) );
  NAND2_X1 U8294 ( .A1(n7694), .A2(n9742), .ZN(n6663) );
  AND2_X1 U8295 ( .A1(n6664), .A2(n6663), .ZN(n6671) );
  XNOR2_X1 U8296 ( .A(n6670), .B(n6671), .ZN(n6777) );
  INV_X1 U8297 ( .A(n6729), .ZN(n6666) );
  INV_X1 U8298 ( .A(n6665), .ZN(n6731) );
  NAND2_X1 U8299 ( .A1(n6666), .A2(n6731), .ZN(n6667) );
  AND2_X1 U8300 ( .A1(n6777), .A2(n6667), .ZN(n6668) );
  NAND2_X1 U8301 ( .A1(n6669), .A2(n6668), .ZN(n6779) );
  INV_X1 U8302 ( .A(n6670), .ZN(n6672) );
  NAND2_X1 U8303 ( .A1(n6672), .A2(n6671), .ZN(n6673) );
  NAND2_X1 U8304 ( .A1(n6779), .A2(n6673), .ZN(n6927) );
  NAND2_X1 U8305 ( .A1(n6897), .A2(n7680), .ZN(n6675) );
  NAND2_X1 U8306 ( .A1(n7694), .A2(n9094), .ZN(n6674) );
  NAND2_X1 U8307 ( .A1(n6675), .A2(n6674), .ZN(n6676) );
  XNOR2_X1 U8308 ( .A(n6676), .B(n7616), .ZN(n6682) );
  INV_X1 U8309 ( .A(n6682), .ZN(n6680) );
  NAND2_X1 U8310 ( .A1(n7693), .A2(n9094), .ZN(n6678) );
  NAND2_X1 U8311 ( .A1(n6897), .A2(n7694), .ZN(n6677) );
  AND2_X1 U8312 ( .A1(n6678), .A2(n6677), .ZN(n6681) );
  INV_X1 U8313 ( .A(n6681), .ZN(n6679) );
  NAND2_X1 U8314 ( .A1(n6680), .A2(n6679), .ZN(n6925) );
  INV_X1 U8315 ( .A(n6925), .ZN(n6683) );
  AND2_X1 U8316 ( .A1(n6682), .A2(n6681), .ZN(n6926) );
  NOR2_X1 U8317 ( .A1(n6683), .A2(n6926), .ZN(n6684) );
  XNOR2_X1 U8318 ( .A(n6927), .B(n6684), .ZN(n6691) );
  AOI21_X1 U8319 ( .B1(n8789), .B2(n9093), .A(n6685), .ZN(n6689) );
  NAND2_X1 U8320 ( .A1(n8807), .A2(n6897), .ZN(n6688) );
  NAND2_X1 U8321 ( .A1(n8802), .A2(n6845), .ZN(n6687) );
  OR2_X1 U8322 ( .A1(n8778), .A2(n6850), .ZN(n6686) );
  NAND4_X1 U8323 ( .A1(n6689), .A2(n6688), .A3(n6687), .A4(n6686), .ZN(n6690)
         );
  AOI21_X1 U8324 ( .B1(n6691), .B2(n8765), .A(n6690), .ZN(n6692) );
  INV_X1 U8325 ( .A(n6692), .ZN(P1_U3211) );
  XOR2_X1 U8326 ( .A(n8882), .B(n9046), .Z(n6697) );
  OAI21_X1 U8327 ( .B1(n6694), .B2(n5646), .A(n6693), .ZN(n9735) );
  OAI22_X1 U8328 ( .A1(n6741), .A2(n9501), .B1(n9502), .B2(n5644), .ZN(n6695)
         );
  AOI21_X1 U8329 ( .B1(n9735), .B2(n9506), .A(n6695), .ZN(n6696) );
  OAI21_X1 U8330 ( .B1(n9497), .B2(n6697), .A(n6696), .ZN(n9733) );
  INV_X1 U8331 ( .A(n9733), .ZN(n6703) );
  INV_X1 U8332 ( .A(n9358), .ZN(n9516) );
  NAND2_X1 U8333 ( .A1(n6698), .A2(n8767), .ZN(n9730) );
  NAND3_X1 U8334 ( .A1(n9361), .A2(n9729), .A3(n9730), .ZN(n6700) );
  AOI22_X1 U8335 ( .A1(n9312), .A2(P1_REG2_REG_2__SCAN_IN), .B1(n9508), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n6699) );
  OAI211_X1 U8336 ( .C1(n9732), .C2(n9357), .A(n6700), .B(n6699), .ZN(n6701)
         );
  AOI21_X1 U8337 ( .B1(n9516), .B2(n9735), .A(n6701), .ZN(n6702) );
  OAI21_X1 U8338 ( .B1(n6703), .B2(n9312), .A(n6702), .ZN(P1_U3289) );
  INV_X1 U8339 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6708) );
  NAND2_X1 U8340 ( .A1(n6706), .A2(n9915), .ZN(n6707) );
  OAI21_X1 U8341 ( .B1(n9915), .B2(n6708), .A(n6707), .ZN(P2_U3460) );
  INV_X1 U8342 ( .A(n8253), .ZN(n8244) );
  OAI222_X1 U8343 ( .A1(n8661), .A2(n6710), .B1(n8657), .B2(n6709), .C1(n8244), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U8344 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6725) );
  NAND2_X1 U8345 ( .A1(n6806), .A2(n9826), .ZN(n6711) );
  NAND2_X1 U8346 ( .A1(n6712), .A2(n6711), .ZN(n6713) );
  NAND2_X1 U8347 ( .A1(n7262), .A2(n7322), .ZN(n7980) );
  INV_X1 U8348 ( .A(n7262), .ZN(n8173) );
  INV_X1 U8349 ( .A(n7322), .ZN(n7261) );
  NAND2_X1 U8350 ( .A1(n8173), .A2(n7261), .ZN(n7997) );
  NAND2_X1 U8351 ( .A1(n7980), .A2(n7997), .ZN(n8118) );
  NAND2_X1 U8352 ( .A1(n6713), .A2(n8118), .ZN(n7264) );
  OAI21_X1 U8353 ( .B1(n6713), .B2(n8118), .A(n7264), .ZN(n7323) );
  INV_X1 U8354 ( .A(n7323), .ZN(n6723) );
  AOI211_X1 U8355 ( .C1(n8118), .C2(n6715), .A(n9813), .B(n7277), .ZN(n6718)
         );
  OR2_X1 U8356 ( .A1(n7287), .A2(n8491), .ZN(n6717) );
  OR2_X1 U8357 ( .A1(n6806), .A2(n8474), .ZN(n6716) );
  NAND2_X1 U8358 ( .A1(n6717), .A2(n6716), .ZN(n6868) );
  NOR2_X1 U8359 ( .A1(n6718), .A2(n6868), .ZN(n7318) );
  NAND2_X1 U8360 ( .A1(n6719), .A2(n7322), .ZN(n6720) );
  NAND2_X1 U8361 ( .A1(n6720), .A2(n8625), .ZN(n6721) );
  NOR2_X1 U8362 ( .A1(n7255), .A2(n6721), .ZN(n7321) );
  AOI21_X1 U8363 ( .B1(n8624), .B2(n7322), .A(n7321), .ZN(n6722) );
  OAI211_X1 U8364 ( .C1(n9864), .C2(n6723), .A(n7318), .B(n6722), .ZN(n6726)
         );
  NAND2_X1 U8365 ( .A1(n6726), .A2(n9927), .ZN(n6724) );
  OAI21_X1 U8366 ( .B1(n9927), .B2(n6725), .A(n6724), .ZN(P2_U3524) );
  INV_X1 U8367 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6728) );
  NAND2_X1 U8368 ( .A1(n6726), .A2(n9915), .ZN(n6727) );
  OAI21_X1 U8369 ( .B1(n9915), .B2(n6728), .A(n6727), .ZN(P2_U3463) );
  NAND2_X1 U8370 ( .A1(n4558), .A2(n6729), .ZN(n6775) );
  OAI21_X1 U8371 ( .B1(n4558), .B2(n6729), .A(n6775), .ZN(n6730) );
  NOR2_X1 U8372 ( .A1(n6730), .A2(n6731), .ZN(n6778) );
  AOI21_X1 U8373 ( .B1(n6731), .B2(n6730), .A(n6778), .ZN(n6737) );
  OAI22_X1 U8374 ( .A1(n6761), .A2(n8750), .B1(n8778), .B2(n6732), .ZN(n6733)
         );
  AOI211_X1 U8375 ( .C1(n8789), .C2(n9095), .A(n6734), .B(n6733), .ZN(n6736)
         );
  NAND2_X1 U8376 ( .A1(n8802), .A2(n6759), .ZN(n6735) );
  OAI211_X1 U8377 ( .C1(n6737), .C2(n8782), .A(n6736), .B(n6735), .ZN(P1_U3225) );
  XNOR2_X1 U8378 ( .A(n8879), .B(n6738), .ZN(n6744) );
  OAI21_X1 U8379 ( .B1(n6740), .B2(n8879), .A(n6739), .ZN(n9740) );
  OAI22_X1 U8380 ( .A1(n6741), .A2(n9502), .B1(n9501), .B2(n6907), .ZN(n6742)
         );
  AOI21_X1 U8381 ( .B1(n9740), .B2(n9506), .A(n6742), .ZN(n6743) );
  OAI21_X1 U8382 ( .B1(n9497), .B2(n6744), .A(n6743), .ZN(n9738) );
  INV_X1 U8383 ( .A(n9738), .ZN(n6753) );
  NAND2_X1 U8384 ( .A1(n6745), .A2(n6747), .ZN(n6746) );
  NAND2_X1 U8385 ( .A1(n6755), .A2(n6746), .ZN(n9737) );
  NAND2_X1 U8386 ( .A1(n9509), .A2(n6747), .ZN(n6750) );
  AOI22_X1 U8387 ( .A1(n9312), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n9508), .B2(
        n6748), .ZN(n6749) );
  OAI211_X1 U8388 ( .C1(n9737), .C2(n7782), .A(n6750), .B(n6749), .ZN(n6751)
         );
  AOI21_X1 U8389 ( .B1(n9740), .B2(n9516), .A(n6751), .ZN(n6752) );
  OAI21_X1 U8390 ( .B1(n6753), .B2(n9312), .A(n6752), .ZN(P1_U3287) );
  XNOR2_X1 U8391 ( .A(n8937), .B(n8885), .ZN(n6754) );
  AOI222_X1 U8392 ( .A1(n9351), .A2(n6754), .B1(n9095), .B2(n9319), .C1(n9097), 
        .C2(n9317), .ZN(n6881) );
  NAND2_X1 U8393 ( .A1(n6755), .A2(n6879), .ZN(n6756) );
  NAND2_X1 U8394 ( .A1(n6756), .A2(n9751), .ZN(n6757) );
  NOR2_X1 U8395 ( .A1(n6914), .A2(n6757), .ZN(n6878) );
  NOR2_X1 U8396 ( .A1(n6758), .A2(n9257), .ZN(n9515) );
  AOI22_X1 U8397 ( .A1(n9519), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n9508), .B2(
        n6759), .ZN(n6760) );
  OAI21_X1 U8398 ( .B1(n9357), .B2(n6761), .A(n6760), .ZN(n6766) );
  OAI21_X1 U8399 ( .B1(n6763), .B2(n8885), .A(n6762), .ZN(n6882) );
  OR2_X1 U8400 ( .A1(n9075), .A2(n7616), .ZN(n6764) );
  NOR2_X1 U8401 ( .A1(n6882), .A2(n9340), .ZN(n6765) );
  AOI211_X1 U8402 ( .C1(n6878), .C2(n9515), .A(n6766), .B(n6765), .ZN(n6767)
         );
  OAI21_X1 U8403 ( .B1(n9519), .B2(n6881), .A(n6767), .ZN(P1_U3286) );
  INV_X1 U8404 ( .A(n7929), .ZN(n6891) );
  NOR2_X1 U8405 ( .A1(n6807), .A2(n8491), .ZN(n9851) );
  NAND2_X1 U8406 ( .A1(n6769), .A2(n6768), .ZN(n6834) );
  AOI22_X1 U8407 ( .A1(n6891), .A2(n9851), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n6834), .ZN(n6773) );
  INV_X1 U8408 ( .A(n6770), .ZN(n9832) );
  NAND2_X1 U8409 ( .A1(n8177), .A2(n4690), .ZN(n8123) );
  INV_X1 U8410 ( .A(n8123), .ZN(n9831) );
  MUX2_X1 U8411 ( .A(n9831), .B(n9852), .S(n5791), .Z(n6771) );
  OAI21_X1 U8412 ( .B1(n9832), .B2(n6771), .A(n7924), .ZN(n6772) );
  OAI211_X1 U8413 ( .C1(n7933), .C2(n4690), .A(n6773), .B(n6772), .ZN(P2_U3234) );
  INV_X1 U8414 ( .A(n6774), .ZN(n6918) );
  INV_X1 U8415 ( .A(n6775), .ZN(n6776) );
  NOR3_X1 U8416 ( .A1(n6778), .A2(n6777), .A3(n6776), .ZN(n6781) );
  INV_X1 U8417 ( .A(n6779), .ZN(n6780) );
  OAI21_X1 U8418 ( .B1(n6781), .B2(n6780), .A(n8765), .ZN(n6785) );
  OAI22_X1 U8419 ( .A1(n6919), .A2(n8750), .B1(n8778), .B2(n6907), .ZN(n6782)
         );
  AOI211_X1 U8420 ( .C1(n8789), .C2(n9094), .A(n6783), .B(n6782), .ZN(n6784)
         );
  OAI211_X1 U8421 ( .C1(n8792), .C2(n6918), .A(n6785), .B(n6784), .ZN(P1_U3237) );
  OAI21_X1 U8422 ( .B1(n6791), .B2(n6788), .A(n6787), .ZN(n7313) );
  NAND2_X1 U8423 ( .A1(n7312), .A2(n9852), .ZN(n6789) );
  NAND2_X1 U8424 ( .A1(n6789), .A2(n8625), .ZN(n6790) );
  OR2_X1 U8425 ( .A1(n6790), .A2(n6802), .ZN(n7307) );
  OAI21_X1 U8426 ( .B1(n6625), .B2(n9905), .A(n7307), .ZN(n6798) );
  INV_X1 U8427 ( .A(n8124), .ZN(n6793) );
  NAND2_X1 U8428 ( .A1(n6791), .A2(n9832), .ZN(n6792) );
  OAI211_X1 U8429 ( .C1(n8127), .C2(n6793), .A(n6792), .B(n9857), .ZN(n6797)
         );
  OR2_X1 U8430 ( .A1(n6794), .A2(n8491), .ZN(n6796) );
  NAND2_X1 U8431 ( .A1(n8177), .A2(n9806), .ZN(n6795) );
  AND2_X1 U8432 ( .A1(n6796), .A2(n6795), .ZN(n6831) );
  NAND2_X1 U8433 ( .A1(n6797), .A2(n6831), .ZN(n7311) );
  AOI211_X1 U8434 ( .C1(n9912), .C2(n7313), .A(n6798), .B(n7311), .ZN(n6855)
         );
  NAND2_X1 U8435 ( .A1(n9924), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6799) );
  OAI21_X1 U8436 ( .B1(n6855), .B2(n9924), .A(n6799), .ZN(P2_U3521) );
  XNOR2_X1 U8437 ( .A(n6800), .B(n8119), .ZN(n7303) );
  OAI211_X1 U8438 ( .C1(n6802), .C2(n6803), .A(n8625), .B(n6801), .ZN(n7298)
         );
  OAI21_X1 U8439 ( .B1(n6803), .B2(n9905), .A(n7298), .ZN(n6811) );
  XNOR2_X1 U8440 ( .A(n6804), .B(n8119), .ZN(n6805) );
  NAND2_X1 U8441 ( .A1(n6805), .A2(n9857), .ZN(n6810) );
  OR2_X1 U8442 ( .A1(n6806), .A2(n8491), .ZN(n6809) );
  OR2_X1 U8443 ( .A1(n6807), .A2(n8474), .ZN(n6808) );
  AND2_X1 U8444 ( .A1(n6809), .A2(n6808), .ZN(n6838) );
  NAND2_X1 U8445 ( .A1(n6810), .A2(n6838), .ZN(n7301) );
  AOI211_X1 U8446 ( .C1(n7303), .C2(n9912), .A(n6811), .B(n7301), .ZN(n6874)
         );
  NAND2_X1 U8447 ( .A1(n9924), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6812) );
  OAI21_X1 U8448 ( .B1(n6874), .B2(n9924), .A(n6812), .ZN(P2_U3522) );
  AOI21_X1 U8449 ( .B1(n6815), .B2(n6814), .A(n6813), .ZN(n6824) );
  NAND2_X1 U8450 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7050) );
  OAI21_X1 U8451 ( .B1(n9691), .B2(n6816), .A(n7050), .ZN(n6821) );
  AOI211_X1 U8452 ( .C1(n6819), .C2(n6818), .A(n6817), .B(n9701), .ZN(n6820)
         );
  AOI211_X1 U8453 ( .C1(P1_ADDR_REG_10__SCAN_IN), .C2(n6822), .A(n6821), .B(
        n6820), .ZN(n6823) );
  OAI21_X1 U8454 ( .B1(n6824), .B2(n9712), .A(n6823), .ZN(P1_U3251) );
  NAND2_X1 U8455 ( .A1(n7941), .A2(n7312), .ZN(n6830) );
  OAI21_X1 U8456 ( .B1(n6827), .B2(n6826), .A(n6825), .ZN(n6828) );
  AOI22_X1 U8457 ( .A1(n7924), .A2(n6828), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n6834), .ZN(n6829) );
  OAI211_X1 U8458 ( .C1(n6831), .C2(n7929), .A(n6830), .B(n6829), .ZN(P2_U3224) );
  NAND2_X1 U8459 ( .A1(n7941), .A2(n7302), .ZN(n6837) );
  XOR2_X1 U8460 ( .A(n6833), .B(n6832), .Z(n6835) );
  AOI22_X1 U8461 ( .A1(n7924), .A2(n6835), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n6834), .ZN(n6836) );
  OAI211_X1 U8462 ( .C1(n6838), .C2(n7929), .A(n6837), .B(n6836), .ZN(P2_U3239) );
  INV_X1 U8463 ( .A(n6839), .ZN(n6877) );
  AOI22_X1 U8464 ( .A1(n8261), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n8654), .ZN(n6840) );
  OAI21_X1 U8465 ( .B1(n6877), .B2(n8657), .A(n6840), .ZN(P2_U3340) );
  OAI21_X1 U8466 ( .B1(n6842), .B2(n8887), .A(n6841), .ZN(n6843) );
  INV_X1 U8467 ( .A(n6843), .ZN(n6900) );
  AOI21_X1 U8468 ( .B1(n6915), .B2(n6897), .A(n9762), .ZN(n6844) );
  AND2_X1 U8469 ( .A1(n6844), .A2(n7219), .ZN(n6896) );
  INV_X1 U8470 ( .A(n6845), .ZN(n6846) );
  OAI22_X1 U8471 ( .A1(n9357), .A2(n4760), .B1(n6846), .B2(n9294), .ZN(n6847)
         );
  AOI21_X1 U8472 ( .B1(n6896), .B2(n9515), .A(n6847), .ZN(n6854) );
  NAND2_X1 U8473 ( .A1(n6848), .A2(n8887), .ZN(n6849) );
  NAND2_X1 U8474 ( .A1(n7211), .A2(n6849), .ZN(n6852) );
  OAI22_X1 U8475 ( .A1(n6850), .A2(n9502), .B1(n9501), .B2(n7198), .ZN(n6851)
         );
  AOI21_X1 U8476 ( .B1(n6852), .B2(n9351), .A(n6851), .ZN(n6899) );
  MUX2_X1 U8477 ( .A(n6899), .B(n6281), .S(n9519), .Z(n6853) );
  OAI211_X1 U8478 ( .C1(n6900), .C2(n9340), .A(n6854), .B(n6853), .ZN(P1_U3284) );
  INV_X1 U8479 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6857) );
  OR2_X1 U8480 ( .A1(n9913), .A2(n6855), .ZN(n6856) );
  OAI21_X1 U8481 ( .B1(n9915), .B2(n6857), .A(n6856), .ZN(P2_U3454) );
  XNOR2_X1 U8482 ( .A(n6859), .B(n6858), .ZN(n6864) );
  OR2_X1 U8483 ( .A1(n7276), .A2(n8491), .ZN(n6861) );
  OR2_X1 U8484 ( .A1(n7262), .A2(n8474), .ZN(n6860) );
  NAND2_X1 U8485 ( .A1(n6861), .A2(n6860), .ZN(n7248) );
  AND2_X1 U8486 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7132) );
  AOI21_X1 U8487 ( .B1(n6891), .B2(n7248), .A(n7132), .ZN(n6863) );
  AOI22_X1 U8488 ( .A1(n7941), .A2(n7246), .B1(n7940), .B2(n7257), .ZN(n6862)
         );
  OAI211_X1 U8489 ( .C1(n6864), .C2(n7944), .A(n6863), .B(n6862), .ZN(P2_U3229) );
  OAI21_X1 U8490 ( .B1(n6867), .B2(n6866), .A(n6865), .ZN(n6872) );
  INV_X1 U8491 ( .A(n6868), .ZN(n6869) );
  INV_X1 U8492 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n7119) );
  OAI22_X1 U8493 ( .A1(n7929), .A2(n6869), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7119), .ZN(n6871) );
  OAI22_X1 U8494 ( .A1(n7933), .A2(n7261), .B1(n7909), .B2(n7316), .ZN(n6870)
         );
  AOI211_X1 U8495 ( .C1(n7924), .C2(n6872), .A(n6871), .B(n6870), .ZN(n6873)
         );
  INV_X1 U8496 ( .A(n6873), .ZN(P2_U3232) );
  INV_X1 U8497 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10273) );
  OR2_X1 U8498 ( .A1(n6874), .A2(n9913), .ZN(n6875) );
  OAI21_X1 U8499 ( .B1(n9915), .B2(n10273), .A(n6875), .ZN(P2_U3457) );
  INV_X1 U8500 ( .A(n9708), .ZN(n9127) );
  INV_X1 U8501 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6876) );
  OAI222_X1 U8502 ( .A1(n9127), .A2(P1_U3084), .B1(n9460), .B2(n6877), .C1(
        n6876), .C2(n7760), .ZN(P1_U3335) );
  INV_X1 U8503 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6884) );
  AOI21_X1 U8504 ( .B1(n9750), .B2(n6879), .A(n6878), .ZN(n6880) );
  OAI211_X1 U8505 ( .C1(n9534), .C2(n6882), .A(n6881), .B(n6880), .ZN(n6885)
         );
  NAND2_X1 U8506 ( .A1(n6885), .A2(n9781), .ZN(n6883) );
  OAI21_X1 U8507 ( .B1(n9781), .B2(n6884), .A(n6883), .ZN(P1_U3528) );
  INV_X1 U8508 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6887) );
  NAND2_X1 U8509 ( .A1(n6885), .A2(n9759), .ZN(n6886) );
  OAI21_X1 U8510 ( .B1(n9759), .B2(n6887), .A(n6886), .ZN(P1_U3469) );
  XNOR2_X1 U8511 ( .A(n6889), .B(n6888), .ZN(n6895) );
  AOI22_X1 U8512 ( .A1(n7941), .A2(n6892), .B1(n6891), .B2(n6890), .ZN(n6894)
         );
  MUX2_X1 U8513 ( .A(n7909), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n6893) );
  OAI211_X1 U8514 ( .C1(n7944), .C2(n6895), .A(n6894), .B(n6893), .ZN(P2_U3220) );
  AOI21_X1 U8515 ( .B1(n9750), .B2(n6897), .A(n6896), .ZN(n6898) );
  OAI211_X1 U8516 ( .C1(n6900), .C2(n9534), .A(n6899), .B(n6898), .ZN(n6902)
         );
  NAND2_X1 U8517 ( .A1(n6902), .A2(n9781), .ZN(n6901) );
  OAI21_X1 U8518 ( .B1(n9781), .B2(n6287), .A(n6901), .ZN(P1_U3530) );
  INV_X1 U8519 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n6904) );
  NAND2_X1 U8520 ( .A1(n6902), .A2(n9759), .ZN(n6903) );
  OAI21_X1 U8521 ( .B1(n9759), .B2(n6904), .A(n6903), .ZN(P1_U3475) );
  OAI21_X1 U8522 ( .B1(n6906), .B2(n5652), .A(n6905), .ZN(n6913) );
  INV_X1 U8523 ( .A(n6913), .ZN(n9746) );
  OAI22_X1 U8524 ( .A1(n6907), .A2(n9502), .B1(n9501), .B2(n7213), .ZN(n6912)
         );
  AND2_X1 U8525 ( .A1(n8939), .A2(n8936), .ZN(n6908) );
  AOI21_X1 U8526 ( .B1(n6909), .B2(n8936), .A(n8939), .ZN(n6910) );
  NOR3_X1 U8527 ( .A1(n4559), .A2(n6910), .A3(n9497), .ZN(n6911) );
  AOI211_X1 U8528 ( .C1(n9506), .C2(n6913), .A(n6912), .B(n6911), .ZN(n9745)
         );
  MUX2_X1 U8529 ( .A(n6279), .B(n9745), .S(n9338), .Z(n6922) );
  INV_X1 U8530 ( .A(n6914), .ZN(n6917) );
  INV_X1 U8531 ( .A(n6915), .ZN(n6916) );
  AOI21_X1 U8532 ( .B1(n9742), .B2(n6917), .A(n6916), .ZN(n9743) );
  OAI22_X1 U8533 ( .A1(n9357), .A2(n6919), .B1(n6918), .B2(n9294), .ZN(n6920)
         );
  AOI21_X1 U8534 ( .B1(n9743), .B2(n9361), .A(n6920), .ZN(n6921) );
  OAI211_X1 U8535 ( .C1(n9746), .C2(n9358), .A(n6922), .B(n6921), .ZN(P1_U3285) );
  INV_X1 U8536 ( .A(n6923), .ZN(n7599) );
  OAI222_X1 U8537 ( .A1(P1_U3084), .A2(n9135), .B1(n9460), .B2(n7599), .C1(
        n6924), .C2(n7760), .ZN(P1_U3334) );
  OAI21_X2 U8538 ( .B1(n6927), .B2(n6926), .A(n6925), .ZN(n6933) );
  NAND2_X1 U8539 ( .A1(n9749), .A2(n7694), .ZN(n6929) );
  NAND2_X1 U8540 ( .A1(n7693), .A2(n9093), .ZN(n6928) );
  NAND2_X1 U8541 ( .A1(n6929), .A2(n6928), .ZN(n6934) );
  NAND2_X1 U8542 ( .A1(n6933), .A2(n6934), .ZN(n7010) );
  NAND2_X1 U8543 ( .A1(n9749), .A2(n7680), .ZN(n6931) );
  NAND2_X1 U8544 ( .A1(n7694), .A2(n9093), .ZN(n6930) );
  NAND2_X1 U8545 ( .A1(n6931), .A2(n6930), .ZN(n6932) );
  XNOR2_X1 U8546 ( .A(n6932), .B(n7616), .ZN(n7013) );
  NAND2_X1 U8547 ( .A1(n7010), .A2(n7013), .ZN(n6937) );
  NAND2_X1 U8548 ( .A1(n7205), .A2(n7680), .ZN(n6939) );
  NAND2_X1 U8549 ( .A1(n7694), .A2(n9092), .ZN(n6938) );
  NAND2_X1 U8550 ( .A1(n6939), .A2(n6938), .ZN(n6940) );
  XNOR2_X1 U8551 ( .A(n6940), .B(n7696), .ZN(n7041) );
  NOR2_X1 U8552 ( .A1(n7677), .A2(n9503), .ZN(n6941) );
  AOI21_X1 U8553 ( .B1(n7205), .B2(n7694), .A(n6941), .ZN(n7042) );
  XNOR2_X1 U8554 ( .A(n7041), .B(n7042), .ZN(n7039) );
  XOR2_X1 U8555 ( .A(n7040), .B(n7039), .Z(n6948) );
  NOR2_X1 U8556 ( .A1(n9761), .A2(n8750), .ZN(n6946) );
  NAND2_X1 U8557 ( .A1(n8789), .A2(n9091), .ZN(n6944) );
  INV_X1 U8558 ( .A(n6942), .ZN(n6943) );
  OAI211_X1 U8559 ( .C1(n7198), .C2(n8778), .A(n6944), .B(n6943), .ZN(n6945)
         );
  AOI211_X1 U8560 ( .C1(n7204), .C2(n8802), .A(n6946), .B(n6945), .ZN(n6947)
         );
  OAI21_X1 U8561 ( .B1(n6948), .B2(n8782), .A(n6947), .ZN(P1_U3229) );
  INV_X1 U8562 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9925) );
  INV_X1 U8563 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6949) );
  MUX2_X1 U8564 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n6949), .S(n7146), .Z(n6965)
         );
  NAND2_X1 U8565 ( .A1(n6993), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6964) );
  INV_X1 U8566 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6950) );
  MUX2_X1 U8567 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n6950), .S(n6993), .Z(n7186)
         );
  NAND2_X1 U8568 ( .A1(n6991), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6963) );
  INV_X1 U8569 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6951) );
  MUX2_X1 U8570 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6951), .S(n6991), .Z(n7174)
         );
  NAND2_X1 U8571 ( .A1(n6989), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6962) );
  INV_X1 U8572 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6952) );
  MUX2_X1 U8573 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6952), .S(n6989), .Z(n7162)
         );
  NAND2_X1 U8574 ( .A1(n6986), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6961) );
  INV_X1 U8575 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6953) );
  MUX2_X1 U8576 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6953), .S(n6986), .Z(n7097)
         );
  NAND2_X1 U8577 ( .A1(n6984), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6960) );
  INV_X1 U8578 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6954) );
  MUX2_X1 U8579 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6954), .S(n6984), .Z(n7135)
         );
  NAND2_X1 U8580 ( .A1(n6981), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6958) );
  MUX2_X1 U8581 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6648), .S(n6981), .Z(n7110)
         );
  NAND2_X1 U8582 ( .A1(n9482), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6957) );
  XOR2_X1 U8583 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n9482), .Z(n9486) );
  INV_X1 U8584 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6955) );
  MUX2_X1 U8585 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6955), .S(n4461), .Z(n9473)
         );
  NAND3_X1 U8586 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n9473), .ZN(n9472) );
  OAI21_X1 U8587 ( .B1(n6956), .B2(n6955), .A(n9472), .ZN(n9485) );
  NAND2_X1 U8588 ( .A1(n9486), .A2(n9485), .ZN(n9484) );
  NAND2_X1 U8589 ( .A1(n6957), .A2(n9484), .ZN(n7109) );
  NAND2_X1 U8590 ( .A1(n7110), .A2(n7109), .ZN(n7108) );
  NAND2_X1 U8591 ( .A1(n6958), .A2(n7108), .ZN(n7123) );
  MUX2_X1 U8592 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6725), .S(n6982), .Z(n7122)
         );
  NAND2_X1 U8593 ( .A1(n7123), .A2(n7122), .ZN(n7121) );
  NAND2_X1 U8594 ( .A1(n6982), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6959) );
  NAND2_X1 U8595 ( .A1(n7121), .A2(n6959), .ZN(n7134) );
  NAND2_X1 U8596 ( .A1(n7135), .A2(n7134), .ZN(n7133) );
  NAND2_X1 U8597 ( .A1(n6960), .A2(n7133), .ZN(n7098) );
  NAND2_X1 U8598 ( .A1(n7097), .A2(n7098), .ZN(n7096) );
  NAND2_X1 U8599 ( .A1(n6961), .A2(n7096), .ZN(n7163) );
  NAND2_X1 U8600 ( .A1(n7162), .A2(n7163), .ZN(n7161) );
  NAND2_X1 U8601 ( .A1(n6962), .A2(n7161), .ZN(n7175) );
  NAND2_X1 U8602 ( .A1(n7174), .A2(n7175), .ZN(n7173) );
  NAND2_X1 U8603 ( .A1(n6963), .A2(n7173), .ZN(n7187) );
  NAND2_X1 U8604 ( .A1(n7186), .A2(n7187), .ZN(n7185) );
  NAND2_X1 U8605 ( .A1(n6964), .A2(n7185), .ZN(n7147) );
  NAND2_X1 U8606 ( .A1(n6965), .A2(n7147), .ZN(n7151) );
  NAND2_X1 U8607 ( .A1(n7146), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6966) );
  NAND2_X1 U8608 ( .A1(n7151), .A2(n6966), .ZN(n8185) );
  INV_X1 U8609 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6967) );
  MUX2_X1 U8610 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n6967), .S(n8183), .Z(n8186)
         );
  NAND2_X1 U8611 ( .A1(n8185), .A2(n8186), .ZN(n8184) );
  NAND2_X1 U8612 ( .A1(n8183), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6968) );
  NAND2_X1 U8613 ( .A1(n8184), .A2(n6968), .ZN(n7061) );
  MUX2_X1 U8614 ( .A(n9925), .B(P2_REG1_REG_12__SCAN_IN), .S(n7062), .Z(n7060)
         );
  NOR2_X1 U8615 ( .A1(n7061), .A2(n7060), .ZN(n7059) );
  AOI21_X1 U8616 ( .B1(n6969), .B2(n9925), .A(n7059), .ZN(n6971) );
  INV_X1 U8617 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7023) );
  AOI22_X1 U8618 ( .A1(n7029), .A2(n7023), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7024), .ZN(n6970) );
  NOR2_X1 U8619 ( .A1(n6971), .A2(n6970), .ZN(n7022) );
  AOI21_X1 U8620 ( .B1(n6971), .B2(n6970), .A(n7022), .ZN(n7009) );
  OR2_X1 U8621 ( .A1(n7003), .A2(P2_U3152), .ZN(n8659) );
  OR2_X1 U8622 ( .A1(n9844), .A2(n6972), .ZN(n6973) );
  OAI211_X1 U8623 ( .C1(n6974), .C2(n8659), .A(n6973), .B(n8162), .ZN(n6999)
         );
  AND2_X1 U8624 ( .A1(n6998), .A2(n6975), .ZN(n6976) );
  NAND2_X1 U8625 ( .A1(n7062), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6977) );
  OAI21_X1 U8626 ( .B1(n7062), .B2(P2_REG2_REG_12__SCAN_IN), .A(n6977), .ZN(
        n7057) );
  XNOR2_X1 U8627 ( .A(n7146), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n7142) );
  INV_X1 U8628 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10075) );
  AND2_X1 U8629 ( .A1(n4461), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6978) );
  NAND2_X1 U8630 ( .A1(n9482), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6979) );
  OAI21_X1 U8631 ( .B1(n9482), .B2(P2_REG2_REG_2__SCAN_IN), .A(n6979), .ZN(
        n9479) );
  NOR2_X1 U8632 ( .A1(n9480), .A2(n9479), .ZN(n9478) );
  AOI21_X1 U8633 ( .B1(n9482), .B2(P2_REG2_REG_2__SCAN_IN), .A(n9478), .ZN(
        n7106) );
  NAND2_X1 U8634 ( .A1(n6981), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6980) );
  OAI21_X1 U8635 ( .B1(n6981), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6980), .ZN(
        n7105) );
  NOR2_X1 U8636 ( .A1(n7106), .A2(n7105), .ZN(n7104) );
  XNOR2_X1 U8637 ( .A(n6982), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n7117) );
  NOR2_X1 U8638 ( .A1(n7118), .A2(n7117), .ZN(n7116) );
  NAND2_X1 U8639 ( .A1(n6984), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6983) );
  OAI21_X1 U8640 ( .B1(n6984), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6983), .ZN(
        n7130) );
  NOR2_X1 U8641 ( .A1(n7131), .A2(n7130), .ZN(n7129) );
  NAND2_X1 U8642 ( .A1(n6986), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6985) );
  OAI21_X1 U8643 ( .B1(n6986), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6985), .ZN(
        n7092) );
  NOR2_X1 U8644 ( .A1(n7093), .A2(n7092), .ZN(n7091) );
  INV_X1 U8645 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6987) );
  MUX2_X1 U8646 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6987), .S(n6989), .Z(n6988)
         );
  INV_X1 U8647 ( .A(n6988), .ZN(n7158) );
  INV_X1 U8648 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6990) );
  MUX2_X1 U8649 ( .A(n6990), .B(P2_REG2_REG_8__SCAN_IN), .S(n6991), .Z(n7170)
         );
  NAND2_X1 U8650 ( .A1(n6993), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6992) );
  OAI21_X1 U8651 ( .B1(n6993), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6992), .ZN(
        n7182) );
  NOR2_X1 U8652 ( .A1(n7183), .A2(n7182), .ZN(n7181) );
  NOR2_X1 U8653 ( .A1(n7142), .A2(n7143), .ZN(n7141) );
  NOR2_X1 U8654 ( .A1(n8183), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6994) );
  AOI21_X1 U8655 ( .B1(n8183), .B2(P2_REG2_REG_11__SCAN_IN), .A(n6994), .ZN(
        n8179) );
  INV_X1 U8656 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6995) );
  AOI22_X1 U8657 ( .A1(n7029), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n6995), .B2(
        n7024), .ZN(n6996) );
  OAI21_X1 U8658 ( .B1(n6997), .B2(n6996), .A(n7028), .ZN(n7002) );
  NAND2_X1 U8659 ( .A1(n6999), .A2(n6998), .ZN(n7000) );
  NAND2_X1 U8660 ( .A1(n7000), .A2(n8176), .ZN(n7004) );
  NOR2_X1 U8661 ( .A1(n7003), .A2(n6975), .ZN(n7001) );
  NAND2_X1 U8662 ( .A1(n7002), .A2(n9782), .ZN(n7008) );
  INV_X1 U8663 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7005) );
  NAND2_X1 U8664 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7884) );
  OAI21_X1 U8665 ( .B1(n8277), .B2(n7005), .A(n7884), .ZN(n7006) );
  AOI21_X1 U8666 ( .B1(n9483), .B2(n7029), .A(n7006), .ZN(n7007) );
  OAI211_X1 U8667 ( .C1(n7009), .C2(n8224), .A(n7008), .B(n7007), .ZN(P2_U3258) );
  NAND2_X1 U8668 ( .A1(n7011), .A2(n7010), .ZN(n7012) );
  XOR2_X1 U8669 ( .A(n7013), .B(n7012), .Z(n7020) );
  AOI21_X1 U8670 ( .B1(n8789), .B2(n9092), .A(n7014), .ZN(n7018) );
  NAND2_X1 U8671 ( .A1(n8807), .A2(n9749), .ZN(n7017) );
  NAND2_X1 U8672 ( .A1(n8802), .A2(n7222), .ZN(n7016) );
  OR2_X1 U8673 ( .A1(n8778), .A2(n7213), .ZN(n7015) );
  NAND4_X1 U8674 ( .A1(n7018), .A2(n7017), .A3(n7016), .A4(n7015), .ZN(n7019)
         );
  AOI21_X1 U8675 ( .B1(n7020), .B2(n8765), .A(n7019), .ZN(n7021) );
  INV_X1 U8676 ( .A(n7021), .ZN(P1_U3219) );
  AOI21_X1 U8677 ( .B1(n7024), .B2(n7023), .A(n7022), .ZN(n7026) );
  INV_X1 U8678 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8198) );
  AOI22_X1 U8679 ( .A1(n8192), .A2(n8198), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n8199), .ZN(n7025) );
  NOR2_X1 U8680 ( .A1(n7026), .A2(n7025), .ZN(n8197) );
  AOI21_X1 U8681 ( .B1(n7026), .B2(n7025), .A(n8197), .ZN(n7038) );
  NOR2_X1 U8682 ( .A1(n8192), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7027) );
  AOI21_X1 U8683 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8192), .A(n7027), .ZN(
        n7031) );
  OAI21_X1 U8684 ( .B1(n7031), .B2(n7030), .A(n8191), .ZN(n7032) );
  NAND2_X1 U8685 ( .A1(n7032), .A2(n9782), .ZN(n7037) );
  INV_X1 U8686 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7034) );
  AND2_X1 U8687 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7799) );
  INV_X1 U8688 ( .A(n7799), .ZN(n7033) );
  OAI21_X1 U8689 ( .B1(n8277), .B2(n7034), .A(n7033), .ZN(n7035) );
  AOI21_X1 U8690 ( .B1(n9483), .B2(n8192), .A(n7035), .ZN(n7036) );
  OAI211_X1 U8691 ( .C1(n7038), .C2(n8224), .A(n7037), .B(n7036), .ZN(P2_U3259) );
  INV_X1 U8692 ( .A(n7041), .ZN(n7043) );
  NAND2_X1 U8693 ( .A1(n7043), .A2(n7042), .ZN(n7044) );
  NAND2_X1 U8694 ( .A1(n9510), .A2(n7680), .ZN(n7046) );
  NAND2_X1 U8695 ( .A1(n7694), .A2(n9091), .ZN(n7045) );
  NAND2_X1 U8696 ( .A1(n7046), .A2(n7045), .ZN(n7047) );
  XNOR2_X1 U8697 ( .A(n7047), .B(n7616), .ZN(n7227) );
  NOR2_X1 U8698 ( .A1(n7677), .A2(n7356), .ZN(n7048) );
  AOI21_X1 U8699 ( .B1(n9510), .B2(n7694), .A(n7048), .ZN(n7228) );
  XNOR2_X1 U8700 ( .A(n7227), .B(n7228), .ZN(n7049) );
  XNOR2_X1 U8701 ( .A(n7232), .B(n7049), .ZN(n7055) );
  NAND2_X1 U8702 ( .A1(n8789), .A2(n9090), .ZN(n7051) );
  OAI211_X1 U8703 ( .C1(n9503), .C2(n8778), .A(n7051), .B(n7050), .ZN(n7053)
         );
  INV_X1 U8704 ( .A(n9510), .ZN(n9521) );
  NOR2_X1 U8705 ( .A1(n9521), .A2(n8750), .ZN(n7052) );
  AOI211_X1 U8706 ( .C1(n9507), .C2(n8802), .A(n7053), .B(n7052), .ZN(n7054)
         );
  OAI21_X1 U8707 ( .B1(n7055), .B2(n8782), .A(n7054), .ZN(P1_U3215) );
  AOI211_X1 U8708 ( .C1(n7058), .C2(n7057), .A(n7056), .B(n9786), .ZN(n7068)
         );
  AOI21_X1 U8709 ( .B1(n7061), .B2(n7060), .A(n7059), .ZN(n7066) );
  NAND2_X1 U8710 ( .A1(n9483), .A2(n7062), .ZN(n7065) );
  NOR2_X1 U8711 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10132), .ZN(n7063) );
  AOI21_X1 U8712 ( .B1(n9788), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7063), .ZN(
        n7064) );
  OAI211_X1 U8713 ( .C1(n7066), .C2(n8224), .A(n7065), .B(n7064), .ZN(n7067)
         );
  OR2_X1 U8714 ( .A1(n7068), .A2(n7067), .ZN(P2_U3257) );
  OAI21_X1 U8715 ( .B1(n7071), .B2(n7070), .A(n7069), .ZN(n7075) );
  OAI22_X1 U8716 ( .A1(n9866), .A2(n7933), .B1(n7937), .B2(n7287), .ZN(n7074)
         );
  INV_X1 U8717 ( .A(n9805), .ZN(n8005) );
  NAND2_X1 U8718 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7094) );
  NAND2_X1 U8719 ( .A1(n7940), .A2(n7282), .ZN(n7072) );
  OAI211_X1 U8720 ( .C1(n7938), .C2(n8005), .A(n7094), .B(n7072), .ZN(n7073)
         );
  AOI211_X1 U8721 ( .C1(n7075), .C2(n7924), .A(n7074), .B(n7073), .ZN(n7076)
         );
  INV_X1 U8722 ( .A(n7076), .ZN(P2_U3241) );
  XNOR2_X1 U8723 ( .A(n7078), .B(n7077), .ZN(n7084) );
  INV_X1 U8724 ( .A(n7938), .ZN(n7913) );
  INV_X1 U8725 ( .A(n7079), .ZN(n7331) );
  AND2_X1 U8726 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7160) );
  INV_X1 U8727 ( .A(n7160), .ZN(n7080) );
  OAI21_X1 U8728 ( .B1(n7909), .B2(n7331), .A(n7080), .ZN(n7082) );
  OAI22_X1 U8729 ( .A1(n9872), .A2(n7933), .B1(n7937), .B2(n7276), .ZN(n7081)
         );
  AOI211_X1 U8730 ( .C1(n7913), .C2(n8170), .A(n7082), .B(n7081), .ZN(n7083)
         );
  OAI21_X1 U8731 ( .B1(n7084), .B2(n7944), .A(n7083), .ZN(P2_U3215) );
  INV_X1 U8732 ( .A(n7085), .ZN(n7087) );
  OAI222_X1 U8733 ( .A1(n8657), .A2(n7087), .B1(P2_U3152), .B2(n6236), .C1(
        n7086), .C2(n8661), .ZN(P2_U3338) );
  OAI222_X1 U8734 ( .A1(n5670), .A2(P1_U3084), .B1(n9460), .B2(n7087), .C1(
        n10222), .C2(n7760), .ZN(P1_U3333) );
  INV_X1 U8735 ( .A(n7089), .ZN(n7762) );
  OAI222_X1 U8736 ( .A1(n8657), .A2(n7762), .B1(P2_U3152), .B2(n7967), .C1(
        n7090), .C2(n8661), .ZN(P2_U3337) );
  AOI211_X1 U8737 ( .C1(n7093), .C2(n7092), .A(n7091), .B(n9786), .ZN(n7103)
         );
  INV_X1 U8738 ( .A(n9483), .ZN(n9785) );
  INV_X1 U8739 ( .A(n7094), .ZN(n7095) );
  AOI21_X1 U8740 ( .B1(n9788), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n7095), .ZN(
        n7100) );
  OAI211_X1 U8741 ( .C1(n7098), .C2(n7097), .A(n9783), .B(n7096), .ZN(n7099)
         );
  OAI211_X1 U8742 ( .C1(n9785), .C2(n7101), .A(n7100), .B(n7099), .ZN(n7102)
         );
  OR2_X1 U8743 ( .A1(n7103), .A2(n7102), .ZN(P2_U3251) );
  AOI211_X1 U8744 ( .C1(n7106), .C2(n7105), .A(n7104), .B(n9786), .ZN(n7115)
         );
  NOR2_X1 U8745 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10240), .ZN(n7107) );
  AOI21_X1 U8746 ( .B1(n9788), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n7107), .ZN(
        n7112) );
  OAI211_X1 U8747 ( .C1(n7110), .C2(n7109), .A(n9783), .B(n7108), .ZN(n7111)
         );
  OAI211_X1 U8748 ( .C1(n9785), .C2(n7113), .A(n7112), .B(n7111), .ZN(n7114)
         );
  OR2_X1 U8749 ( .A1(n7115), .A2(n7114), .ZN(P2_U3248) );
  AOI211_X1 U8750 ( .C1(n7118), .C2(n7117), .A(n7116), .B(n9786), .ZN(n7128)
         );
  NOR2_X1 U8751 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7119), .ZN(n7120) );
  AOI21_X1 U8752 ( .B1(n9788), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n7120), .ZN(
        n7125) );
  OAI211_X1 U8753 ( .C1(n7123), .C2(n7122), .A(n9783), .B(n7121), .ZN(n7124)
         );
  OAI211_X1 U8754 ( .C1(n9785), .C2(n7126), .A(n7125), .B(n7124), .ZN(n7127)
         );
  OR2_X1 U8755 ( .A1(n7128), .A2(n7127), .ZN(P2_U3249) );
  AOI211_X1 U8756 ( .C1(n7131), .C2(n7130), .A(n7129), .B(n9786), .ZN(n7140)
         );
  AOI21_X1 U8757 ( .B1(n9788), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n7132), .ZN(
        n7137) );
  OAI211_X1 U8758 ( .C1(n7135), .C2(n7134), .A(n9783), .B(n7133), .ZN(n7136)
         );
  OAI211_X1 U8759 ( .C1(n9785), .C2(n7138), .A(n7137), .B(n7136), .ZN(n7139)
         );
  OR2_X1 U8760 ( .A1(n7140), .A2(n7139), .ZN(P2_U3250) );
  AOI211_X1 U8761 ( .C1(n7143), .C2(n7142), .A(n7141), .B(n9786), .ZN(n7156)
         );
  INV_X1 U8762 ( .A(n7144), .ZN(n7145) );
  AOI21_X1 U8763 ( .B1(n9788), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7145), .ZN(
        n7153) );
  MUX2_X1 U8764 ( .A(n6949), .B(P2_REG1_REG_10__SCAN_IN), .S(n7146), .Z(n7149)
         );
  INV_X1 U8765 ( .A(n7147), .ZN(n7148) );
  NAND2_X1 U8766 ( .A1(n7149), .A2(n7148), .ZN(n7150) );
  NAND3_X1 U8767 ( .A1(n9783), .A2(n7151), .A3(n7150), .ZN(n7152) );
  OAI211_X1 U8768 ( .C1(n9785), .C2(n7154), .A(n7153), .B(n7152), .ZN(n7155)
         );
  OR2_X1 U8769 ( .A1(n7156), .A2(n7155), .ZN(P2_U3255) );
  AOI211_X1 U8770 ( .C1(n7159), .C2(n7158), .A(n7157), .B(n9786), .ZN(n7168)
         );
  AOI21_X1 U8771 ( .B1(n9788), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7160), .ZN(
        n7165) );
  OAI211_X1 U8772 ( .C1(n7163), .C2(n7162), .A(n9783), .B(n7161), .ZN(n7164)
         );
  OAI211_X1 U8773 ( .C1(n9785), .C2(n7166), .A(n7165), .B(n7164), .ZN(n7167)
         );
  OR2_X1 U8774 ( .A1(n7168), .A2(n7167), .ZN(P2_U3252) );
  AOI211_X1 U8775 ( .C1(n7171), .C2(n7170), .A(n7169), .B(n9786), .ZN(n7180)
         );
  NAND2_X1 U8776 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n7270) );
  INV_X1 U8777 ( .A(n7270), .ZN(n7172) );
  AOI21_X1 U8778 ( .B1(n9788), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n7172), .ZN(
        n7177) );
  OAI211_X1 U8779 ( .C1(n7175), .C2(n7174), .A(n9783), .B(n7173), .ZN(n7176)
         );
  OAI211_X1 U8780 ( .C1(n9785), .C2(n7178), .A(n7177), .B(n7176), .ZN(n7179)
         );
  OR2_X1 U8781 ( .A1(n7180), .A2(n7179), .ZN(P2_U3253) );
  AOI211_X1 U8782 ( .C1(n7183), .C2(n7182), .A(n7181), .B(n9786), .ZN(n7192)
         );
  NAND2_X1 U8783 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7348) );
  INV_X1 U8784 ( .A(n7348), .ZN(n7184) );
  AOI21_X1 U8785 ( .B1(n9788), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7184), .ZN(
        n7189) );
  OAI211_X1 U8786 ( .C1(n7187), .C2(n7186), .A(n9783), .B(n7185), .ZN(n7188)
         );
  OAI211_X1 U8787 ( .C1(n9785), .C2(n7190), .A(n7189), .B(n7188), .ZN(n7191)
         );
  OR2_X1 U8788 ( .A1(n7192), .A2(n7191), .ZN(P2_U3254) );
  NAND2_X1 U8789 ( .A1(n7193), .A2(n9494), .ZN(n8890) );
  XNOR2_X1 U8790 ( .A(n7194), .B(n8890), .ZN(n7202) );
  NAND2_X1 U8791 ( .A1(n7196), .A2(n7195), .ZN(n7197) );
  XNOR2_X1 U8792 ( .A(n7197), .B(n8890), .ZN(n7200) );
  OAI22_X1 U8793 ( .A1(n7356), .A2(n9501), .B1(n9502), .B2(n7198), .ZN(n7199)
         );
  AOI21_X1 U8794 ( .B1(n7200), .B2(n9351), .A(n7199), .ZN(n7201) );
  OAI21_X1 U8795 ( .B1(n7202), .B2(n9347), .A(n7201), .ZN(n9764) );
  INV_X1 U8796 ( .A(n9764), .ZN(n7210) );
  INV_X1 U8797 ( .A(n7202), .ZN(n9766) );
  OR2_X1 U8798 ( .A1(n7221), .A2(n9761), .ZN(n7203) );
  NAND2_X1 U8799 ( .A1(n9511), .A2(n7203), .ZN(n9763) );
  AOI22_X1 U8800 ( .A1(n9312), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n9508), .B2(
        n7204), .ZN(n7207) );
  NAND2_X1 U8801 ( .A1(n9509), .A2(n7205), .ZN(n7206) );
  OAI211_X1 U8802 ( .C1(n9763), .C2(n7782), .A(n7207), .B(n7206), .ZN(n7208)
         );
  AOI21_X1 U8803 ( .B1(n9766), .B2(n9516), .A(n7208), .ZN(n7209) );
  OAI21_X1 U8804 ( .B1(n7210), .B2(n9312), .A(n7209), .ZN(P1_U3282) );
  NAND2_X1 U8805 ( .A1(n7211), .A2(n8941), .ZN(n7212) );
  INV_X1 U8806 ( .A(n7215), .ZN(n8888) );
  XNOR2_X1 U8807 ( .A(n7212), .B(n8888), .ZN(n7218) );
  OAI22_X1 U8808 ( .A1(n9503), .A2(n9501), .B1(n9502), .B2(n7213), .ZN(n7217)
         );
  OAI21_X1 U8809 ( .B1(n4564), .B2(n7215), .A(n7214), .ZN(n9755) );
  NOR2_X1 U8810 ( .A1(n9755), .A2(n9347), .ZN(n7216) );
  AOI211_X1 U8811 ( .C1(n7218), .C2(n9351), .A(n7217), .B(n7216), .ZN(n9754)
         );
  AND2_X1 U8812 ( .A1(n7219), .A2(n9749), .ZN(n7220) );
  NOR2_X1 U8813 ( .A1(n7221), .A2(n7220), .ZN(n9752) );
  AOI22_X1 U8814 ( .A1(n9519), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n9508), .B2(
        n7222), .ZN(n7223) );
  OAI21_X1 U8815 ( .B1(n9357), .B2(n4758), .A(n7223), .ZN(n7225) );
  NOR2_X1 U8816 ( .A1(n9755), .A2(n9358), .ZN(n7224) );
  AOI211_X1 U8817 ( .C1(n9361), .C2(n9752), .A(n7225), .B(n7224), .ZN(n7226)
         );
  OAI21_X1 U8818 ( .B1(n9754), .B2(n9519), .A(n7226), .ZN(P1_U3283) );
  AND2_X1 U8819 ( .A1(n7227), .A2(n7228), .ZN(n7231) );
  INV_X1 U8820 ( .A(n7227), .ZN(n7230) );
  INV_X1 U8821 ( .A(n7228), .ZN(n7229) );
  NAND2_X1 U8822 ( .A1(n9555), .A2(n7680), .ZN(n7235) );
  NAND2_X1 U8823 ( .A1(n7694), .A2(n9090), .ZN(n7234) );
  NAND2_X1 U8824 ( .A1(n7235), .A2(n7234), .ZN(n7236) );
  XNOR2_X1 U8825 ( .A(n7236), .B(n7696), .ZN(n7458) );
  NOR2_X1 U8826 ( .A1(n7677), .A2(n9500), .ZN(n7237) );
  AOI21_X1 U8827 ( .B1(n9555), .B2(n7694), .A(n7237), .ZN(n7456) );
  XNOR2_X1 U8828 ( .A(n7458), .B(n7456), .ZN(n7454) );
  XNOR2_X1 U8829 ( .A(n7455), .B(n7454), .ZN(n7244) );
  NAND2_X1 U8830 ( .A1(n8789), .A2(n9089), .ZN(n7241) );
  OR2_X1 U8831 ( .A1(n8778), .A2(n7356), .ZN(n7240) );
  NAND2_X1 U8832 ( .A1(n8802), .A2(n7362), .ZN(n7239) );
  NAND4_X1 U8833 ( .A1(n7241), .A2(n7240), .A3(n7239), .A4(n7238), .ZN(n7242)
         );
  AOI21_X1 U8834 ( .B1(n9555), .B2(n8807), .A(n7242), .ZN(n7243) );
  OAI21_X1 U8835 ( .B1(n7244), .B2(n8782), .A(n7243), .ZN(P1_U3234) );
  INV_X1 U8836 ( .A(n7997), .ZN(n7245) );
  NOR2_X1 U8837 ( .A1(n7277), .A2(n7245), .ZN(n7247) );
  NAND2_X1 U8838 ( .A1(n7287), .A2(n7246), .ZN(n7981) );
  INV_X1 U8839 ( .A(n7287), .ZN(n8172) );
  XNOR2_X1 U8840 ( .A(n7247), .B(n8122), .ZN(n7249) );
  AOI21_X1 U8841 ( .B1(n7249), .B2(n9857), .A(n7248), .ZN(n9859) );
  INV_X1 U8842 ( .A(n7250), .ZN(n7253) );
  NAND3_X1 U8843 ( .A1(n7253), .A2(n7252), .A3(n7251), .ZN(n7280) );
  NOR2_X1 U8844 ( .A1(n9842), .A2(n8273), .ZN(n8495) );
  INV_X1 U8845 ( .A(n7281), .ZN(n7254) );
  OAI211_X1 U8846 ( .C1(n9860), .C2(n7255), .A(n7254), .B(n8625), .ZN(n9858)
         );
  INV_X1 U8847 ( .A(n9858), .ZN(n7260) );
  NAND2_X2 U8848 ( .A1(n9840), .A2(n7256), .ZN(n9835) );
  AOI22_X1 U8849 ( .A1(n9842), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n7257), .B2(
        n9838), .ZN(n7258) );
  OAI21_X1 U8850 ( .B1(n9860), .B2(n9835), .A(n7258), .ZN(n7259) );
  AOI21_X1 U8851 ( .B1(n8495), .B2(n7260), .A(n7259), .ZN(n7267) );
  NAND2_X1 U8852 ( .A1(n7262), .A2(n7261), .ZN(n7263) );
  NAND2_X1 U8853 ( .A1(n7264), .A2(n7263), .ZN(n7286) );
  XNOR2_X1 U8854 ( .A(n7286), .B(n7285), .ZN(n9862) );
  OR2_X1 U8855 ( .A1(n7265), .A2(n8149), .ZN(n7370) );
  NAND2_X1 U8856 ( .A1(n7402), .A2(n7370), .ZN(n9833) );
  NAND2_X1 U8857 ( .A1(n9862), .A2(n8512), .ZN(n7266) );
  OAI211_X1 U8858 ( .C1(n9859), .C2(n9842), .A(n7267), .B(n7266), .ZN(P2_U3291) );
  XNOR2_X1 U8859 ( .A(n7269), .B(n7268), .ZN(n7275) );
  INV_X1 U8860 ( .A(n9815), .ZN(n7271) );
  OAI21_X1 U8861 ( .B1(n7909), .B2(n7271), .A(n7270), .ZN(n7273) );
  INV_X1 U8862 ( .A(n9797), .ZN(n9879) );
  OAI22_X1 U8863 ( .A1(n9879), .A2(n7933), .B1(n7937), .B2(n8005), .ZN(n7272)
         );
  AOI211_X1 U8864 ( .C1(n7913), .C2(n9808), .A(n7273), .B(n7272), .ZN(n7274)
         );
  OAI21_X1 U8865 ( .B1(n7275), .B2(n7944), .A(n7274), .ZN(P2_U3223) );
  NAND2_X1 U8866 ( .A1(n7276), .A2(n7326), .ZN(n8006) );
  NAND2_X1 U8867 ( .A1(n8171), .A2(n9866), .ZN(n8000) );
  NAND2_X1 U8868 ( .A1(n8122), .A2(n7997), .ZN(n7278) );
  OAI21_X1 U8869 ( .B1(n7278), .B2(n7277), .A(n7981), .ZN(n7337) );
  XOR2_X1 U8870 ( .A(n8120), .B(n7337), .Z(n7279) );
  OAI222_X1 U8871 ( .A1(n8491), .A2(n8005), .B1(n8474), .B2(n7287), .C1(n7279), 
        .C2(n9813), .ZN(n9868) );
  INV_X1 U8872 ( .A(n9868), .ZN(n7295) );
  OR2_X1 U8873 ( .A1(n7280), .A2(n8273), .ZN(n7308) );
  INV_X1 U8874 ( .A(n7308), .ZN(n9823) );
  OAI21_X1 U8875 ( .B1(n7281), .B2(n9866), .A(n7332), .ZN(n9867) );
  AOI22_X1 U8876 ( .A1(n9842), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n7282), .B2(
        n9838), .ZN(n7283) );
  OAI21_X1 U8877 ( .B1(n9836), .B2(n9867), .A(n7283), .ZN(n7284) );
  AOI21_X1 U8878 ( .B1(n7410), .B2(n7326), .A(n7284), .ZN(n7294) );
  NAND2_X1 U8879 ( .A1(n7286), .A2(n7285), .ZN(n7289) );
  NAND2_X1 U8880 ( .A1(n7287), .A2(n9860), .ZN(n7288) );
  AND2_X1 U8881 ( .A1(n7290), .A2(n8120), .ZN(n9865) );
  INV_X1 U8882 ( .A(n9865), .ZN(n7292) );
  NAND3_X1 U8883 ( .A1(n7292), .A2(n8512), .A3(n7328), .ZN(n7293) );
  OAI211_X1 U8884 ( .C1(n7295), .C2(n9842), .A(n7294), .B(n7293), .ZN(P2_U3290) );
  INV_X1 U8885 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7296) );
  NOR2_X1 U8886 ( .A1(n9840), .A2(n7296), .ZN(n7300) );
  INV_X1 U8887 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7297) );
  OAI22_X1 U8888 ( .A1(n7308), .A2(n7298), .B1(n7297), .B2(n8345), .ZN(n7299)
         );
  AOI211_X1 U8889 ( .C1(n9840), .C2(n7301), .A(n7300), .B(n7299), .ZN(n7305)
         );
  AOI22_X1 U8890 ( .A1(n7303), .A2(n8512), .B1(n7410), .B2(n7302), .ZN(n7304)
         );
  NAND2_X1 U8891 ( .A1(n7305), .A2(n7304), .ZN(P2_U3294) );
  INV_X1 U8892 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10210) );
  NOR2_X1 U8893 ( .A1(n9840), .A2(n10210), .ZN(n7310) );
  INV_X1 U8894 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7306) );
  OAI22_X1 U8895 ( .A1(n7308), .A2(n7307), .B1(n7306), .B2(n8345), .ZN(n7309)
         );
  AOI211_X1 U8896 ( .C1(n9840), .C2(n7311), .A(n7310), .B(n7309), .ZN(n7315)
         );
  AOI22_X1 U8897 ( .A1(n8512), .A2(n7313), .B1(n7410), .B2(n7312), .ZN(n7314)
         );
  NAND2_X1 U8898 ( .A1(n7315), .A2(n7314), .ZN(P2_U3295) );
  NOR2_X1 U8899 ( .A1(n8345), .A2(n7316), .ZN(n7320) );
  NAND2_X1 U8900 ( .A1(n9842), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7317) );
  OAI21_X1 U8901 ( .B1(n7318), .B2(n9842), .A(n7317), .ZN(n7319) );
  AOI211_X1 U8902 ( .C1(n7321), .C2(n9823), .A(n7320), .B(n7319), .ZN(n7325)
         );
  AOI22_X1 U8903 ( .A1(n7323), .A2(n8512), .B1(n7410), .B2(n7322), .ZN(n7324)
         );
  NAND2_X1 U8904 ( .A1(n7325), .A2(n7324), .ZN(P2_U3292) );
  NAND2_X1 U8905 ( .A1(n8171), .A2(n7326), .ZN(n7327) );
  XNOR2_X1 U8906 ( .A(n9805), .B(n8004), .ZN(n8129) );
  INV_X1 U8907 ( .A(n8129), .ZN(n7329) );
  OAI21_X1 U8908 ( .B1(n7330), .B2(n7329), .A(n7368), .ZN(n9876) );
  INV_X1 U8909 ( .A(n9876), .ZN(n7343) );
  OAI22_X1 U8910 ( .A1(n9840), .A2(n6987), .B1(n7331), .B2(n8345), .ZN(n7335)
         );
  INV_X1 U8911 ( .A(n7332), .ZN(n7333) );
  OAI21_X1 U8912 ( .B1(n7333), .B2(n9872), .A(n9798), .ZN(n9873) );
  NOR2_X1 U8913 ( .A1(n9836), .A2(n9873), .ZN(n7334) );
  AOI211_X1 U8914 ( .C1(n7410), .C2(n8004), .A(n7335), .B(n7334), .ZN(n7342)
         );
  INV_X1 U8915 ( .A(n8006), .ZN(n7336) );
  OAI211_X1 U8916 ( .C1(n7338), .C2(n8129), .A(n7372), .B(n9857), .ZN(n7340)
         );
  AOI22_X1 U8917 ( .A1(n9806), .A2(n8171), .B1(n8170), .B2(n9807), .ZN(n7339)
         );
  NAND2_X1 U8918 ( .A1(n7340), .A2(n7339), .ZN(n9874) );
  NAND2_X1 U8919 ( .A1(n9874), .A2(n9840), .ZN(n7341) );
  OAI211_X1 U8920 ( .C1(n7343), .C2(n8529), .A(n7342), .B(n7341), .ZN(P2_U3289) );
  NAND2_X1 U8921 ( .A1(n7345), .A2(n7344), .ZN(n7346) );
  XNOR2_X1 U8922 ( .A(n7347), .B(n7346), .ZN(n7353) );
  INV_X1 U8923 ( .A(n7910), .ZN(n8169) );
  INV_X1 U8924 ( .A(n7378), .ZN(n7349) );
  OAI21_X1 U8925 ( .B1(n7909), .B2(n7349), .A(n7348), .ZN(n7351) );
  OAI22_X1 U8926 ( .A1(n7385), .A2(n7933), .B1(n7937), .B2(n7369), .ZN(n7350)
         );
  AOI211_X1 U8927 ( .C1(n7913), .C2(n8169), .A(n7351), .B(n7350), .ZN(n7352)
         );
  OAI21_X1 U8928 ( .B1(n7353), .B2(n7944), .A(n7352), .ZN(P2_U3233) );
  XNOR2_X1 U8929 ( .A(n9555), .B(n9500), .ZN(n8953) );
  XNOR2_X1 U8930 ( .A(n7354), .B(n8953), .ZN(n9559) );
  XNOR2_X1 U8931 ( .A(n7355), .B(n4588), .ZN(n7359) );
  OAI22_X1 U8932 ( .A1(n7356), .A2(n9502), .B1(n9501), .B2(n7528), .ZN(n7357)
         );
  INV_X1 U8933 ( .A(n7357), .ZN(n7358) );
  OAI21_X1 U8934 ( .B1(n7359), .B2(n9497), .A(n7358), .ZN(n7360) );
  AOI21_X1 U8935 ( .B1(n9559), .B2(n9506), .A(n7360), .ZN(n9561) );
  AND2_X1 U8936 ( .A1(n9512), .A2(n9555), .ZN(n7361) );
  OR2_X1 U8937 ( .A1(n7361), .A2(n7482), .ZN(n9557) );
  AOI22_X1 U8938 ( .A1(n9519), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9508), .B2(
        n7362), .ZN(n7364) );
  NAND2_X1 U8939 ( .A1(n9555), .A2(n9509), .ZN(n7363) );
  OAI211_X1 U8940 ( .C1(n9557), .C2(n7782), .A(n7364), .B(n7363), .ZN(n7365)
         );
  AOI21_X1 U8941 ( .B1(n9559), .B2(n9516), .A(n7365), .ZN(n7366) );
  OAI21_X1 U8942 ( .B1(n9561), .B2(n9519), .A(n7366), .ZN(P1_U3280) );
  NAND2_X1 U8943 ( .A1(n8005), .A2(n9872), .ZN(n7367) );
  NAND2_X1 U8944 ( .A1(n7369), .A2(n9797), .ZN(n8015) );
  NAND2_X1 U8945 ( .A1(n8170), .A2(n9879), .ZN(n8010) );
  NAND2_X1 U8946 ( .A1(n7398), .A2(n7384), .ZN(n8018) );
  NAND2_X1 U8947 ( .A1(n9808), .A2(n7385), .ZN(n8014) );
  NAND2_X1 U8948 ( .A1(n8018), .A2(n8014), .ZN(n8131) );
  OAI21_X1 U8949 ( .B1(n4554), .B2(n8131), .A(n7387), .ZN(n9888) );
  INV_X1 U8950 ( .A(n9888), .ZN(n7383) );
  INV_X1 U8951 ( .A(n7370), .ZN(n7371) );
  AND2_X1 U8952 ( .A1(n9840), .A2(n7371), .ZN(n9821) );
  INV_X1 U8953 ( .A(n9821), .ZN(n9801) );
  INV_X1 U8954 ( .A(n9793), .ZN(n9804) );
  XOR2_X1 U8955 ( .A(n7389), .B(n8131), .Z(n7375) );
  AOI22_X1 U8956 ( .A1(n9806), .A2(n8170), .B1(n8169), .B2(n9807), .ZN(n7374)
         );
  NAND2_X1 U8957 ( .A1(n9888), .A2(n9810), .ZN(n7373) );
  OAI211_X1 U8958 ( .C1(n7375), .C2(n9813), .A(n7374), .B(n7373), .ZN(n9886)
         );
  NAND2_X1 U8959 ( .A1(n9886), .A2(n9840), .ZN(n7382) );
  INV_X1 U8960 ( .A(n9800), .ZN(n7377) );
  NOR2_X2 U8961 ( .A1(n9800), .A2(n7384), .ZN(n7405) );
  INV_X1 U8962 ( .A(n7405), .ZN(n7376) );
  OAI21_X1 U8963 ( .B1(n7385), .B2(n7377), .A(n7376), .ZN(n9885) );
  AOI22_X1 U8964 ( .A1(n9842), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7378), .B2(
        n9838), .ZN(n7379) );
  OAI21_X1 U8965 ( .B1(n9885), .B2(n9836), .A(n7379), .ZN(n7380) );
  AOI21_X1 U8966 ( .B1(n7410), .B2(n7384), .A(n7380), .ZN(n7381) );
  OAI211_X1 U8967 ( .C1(n7383), .C2(n9801), .A(n7382), .B(n7381), .ZN(P2_U3287) );
  NAND2_X1 U8968 ( .A1(n7910), .A2(n7409), .ZN(n8026) );
  NAND2_X1 U8969 ( .A1(n9891), .A2(n8169), .ZN(n8025) );
  OR2_X1 U8970 ( .A1(n7828), .A2(n7517), .ZN(n8033) );
  NAND2_X1 U8971 ( .A1(n7517), .A2(n7828), .ZN(n8031) );
  NAND2_X1 U8972 ( .A1(n8033), .A2(n8031), .ZN(n8133) );
  OAI21_X1 U8973 ( .B1(n7388), .B2(n8133), .A(n7512), .ZN(n9898) );
  INV_X1 U8974 ( .A(n8014), .ZN(n8020) );
  OAI21_X1 U8975 ( .B1(n7389), .B2(n8020), .A(n8018), .ZN(n7397) );
  INV_X1 U8976 ( .A(n7396), .ZN(n8132) );
  OAI21_X1 U8977 ( .B1(n7397), .B2(n8132), .A(n8025), .ZN(n7515) );
  XOR2_X1 U8978 ( .A(n8133), .B(n7515), .Z(n7390) );
  OAI222_X1 U8979 ( .A1(n8474), .A2(n7910), .B1(n8491), .B2(n7906), .C1(n9813), 
        .C2(n7390), .ZN(n9901) );
  NAND2_X1 U8980 ( .A1(n7405), .A2(n9891), .ZN(n7518) );
  XNOR2_X1 U8981 ( .A(n7518), .B(n7517), .ZN(n9900) );
  NOR2_X1 U8982 ( .A1(n9900), .A2(n9836), .ZN(n7393) );
  INV_X1 U8983 ( .A(n7517), .ZN(n9899) );
  AOI22_X1 U8984 ( .A1(n9842), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7907), .B2(
        n9838), .ZN(n7391) );
  OAI21_X1 U8985 ( .B1(n9899), .B2(n9835), .A(n7391), .ZN(n7392) );
  AOI211_X1 U8986 ( .C1(n9901), .C2(n9840), .A(n7393), .B(n7392), .ZN(n7394)
         );
  OAI21_X1 U8987 ( .B1(n8529), .B2(n9898), .A(n7394), .ZN(P2_U3285) );
  XNOR2_X1 U8988 ( .A(n7395), .B(n7396), .ZN(n9890) );
  XNOR2_X1 U8989 ( .A(n7397), .B(n7396), .ZN(n7400) );
  OAI22_X1 U8990 ( .A1(n7398), .A2(n8474), .B1(n7828), .B2(n8491), .ZN(n7399)
         );
  AOI21_X1 U8991 ( .B1(n7400), .B2(n9857), .A(n7399), .ZN(n7401) );
  OAI21_X1 U8992 ( .B1(n9890), .B2(n7402), .A(n7401), .ZN(n9893) );
  NAND2_X1 U8993 ( .A1(n9893), .A2(n9840), .ZN(n7412) );
  INV_X1 U8994 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7404) );
  OAI22_X1 U8995 ( .A1(n9840), .A2(n7404), .B1(n7403), .B2(n8345), .ZN(n7408)
         );
  OR2_X1 U8996 ( .A1(n7405), .A2(n9891), .ZN(n7406) );
  NAND2_X1 U8997 ( .A1(n7518), .A2(n7406), .ZN(n9892) );
  NOR2_X1 U8998 ( .A1(n9892), .A2(n9836), .ZN(n7407) );
  AOI211_X1 U8999 ( .C1(n7410), .C2(n7409), .A(n7408), .B(n7407), .ZN(n7411)
         );
  OAI211_X1 U9000 ( .C1(n9890), .C2(n9801), .A(n7412), .B(n7411), .ZN(P2_U3286) );
  INV_X1 U9001 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10337) );
  NOR2_X1 U9002 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7413) );
  AOI21_X1 U9003 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7413), .ZN(n9936) );
  NOR2_X1 U9004 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7414) );
  AOI21_X1 U9005 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7414), .ZN(n9939) );
  NOR2_X1 U9006 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7415) );
  AOI21_X1 U9007 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7415), .ZN(n9942) );
  NOR2_X1 U9008 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7416) );
  AOI21_X1 U9009 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7416), .ZN(n9945) );
  NOR2_X1 U9010 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7417) );
  AOI21_X1 U9011 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7417), .ZN(n9948) );
  NOR2_X1 U9012 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7423) );
  XOR2_X1 U9013 ( .A(n9617), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10348) );
  NAND2_X1 U9014 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7421) );
  XNOR2_X1 U9015 ( .A(n6487), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(n10346) );
  NAND2_X1 U9016 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7419) );
  INV_X1 U9017 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9600) );
  XNOR2_X1 U9018 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n9600), .ZN(n10331) );
  AOI21_X1 U9019 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9928) );
  INV_X1 U9020 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9932) );
  NAND3_X1 U9021 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9930) );
  OAI21_X1 U9022 ( .B1(n9928), .B2(n9932), .A(n9930), .ZN(n10330) );
  NAND2_X1 U9023 ( .A1(n10331), .A2(n10330), .ZN(n7418) );
  NAND2_X1 U9024 ( .A1(n7419), .A2(n7418), .ZN(n10345) );
  NAND2_X1 U9025 ( .A1(n10346), .A2(n10345), .ZN(n7420) );
  NAND2_X1 U9026 ( .A1(n7421), .A2(n7420), .ZN(n10347) );
  NOR2_X1 U9027 ( .A1(n10348), .A2(n10347), .ZN(n7422) );
  NOR2_X1 U9028 ( .A1(n7423), .A2(n7422), .ZN(n7424) );
  NOR2_X1 U9029 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7424), .ZN(n10333) );
  AND2_X1 U9030 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7424), .ZN(n10332) );
  NOR2_X1 U9031 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10332), .ZN(n7425) );
  NOR2_X1 U9032 ( .A1(n10333), .A2(n7425), .ZN(n7426) );
  NAND2_X1 U9033 ( .A1(n7426), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7428) );
  XOR2_X1 U9034 ( .A(n7426), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10329) );
  NAND2_X1 U9035 ( .A1(n10329), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7427) );
  NAND2_X1 U9036 ( .A1(n7428), .A2(n7427), .ZN(n7429) );
  NAND2_X1 U9037 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7429), .ZN(n7431) );
  XOR2_X1 U9038 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7429), .Z(n10344) );
  NAND2_X1 U9039 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10344), .ZN(n7430) );
  NAND2_X1 U9040 ( .A1(n7431), .A2(n7430), .ZN(n7432) );
  NAND2_X1 U9041 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7432), .ZN(n7434) );
  XOR2_X1 U9042 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7432), .Z(n10343) );
  NAND2_X1 U9043 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10343), .ZN(n7433) );
  NAND2_X1 U9044 ( .A1(n7434), .A2(n7433), .ZN(n7435) );
  AND2_X1 U9045 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7435), .ZN(n7436) );
  XNOR2_X1 U9046 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7435), .ZN(n10341) );
  NOR2_X1 U9047 ( .A1(n10342), .A2(n10341), .ZN(n10340) );
  NAND2_X1 U9048 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7437) );
  OAI21_X1 U9049 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7437), .ZN(n9956) );
  NAND2_X1 U9050 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7438) );
  OAI21_X1 U9051 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7438), .ZN(n9953) );
  NOR2_X1 U9052 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7439) );
  AOI21_X1 U9053 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7439), .ZN(n9950) );
  NAND2_X1 U9054 ( .A1(n9951), .A2(n9950), .ZN(n9949) );
  NAND2_X1 U9055 ( .A1(n9948), .A2(n9947), .ZN(n9946) );
  OAI21_X1 U9056 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9946), .ZN(n9944) );
  NAND2_X1 U9057 ( .A1(n9945), .A2(n9944), .ZN(n9943) );
  OAI21_X1 U9058 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9943), .ZN(n9941) );
  NAND2_X1 U9059 ( .A1(n9942), .A2(n9941), .ZN(n9940) );
  OAI21_X1 U9060 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9940), .ZN(n9938) );
  NAND2_X1 U9061 ( .A1(n9939), .A2(n9938), .ZN(n9937) );
  OAI21_X1 U9062 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9937), .ZN(n9935) );
  NAND2_X1 U9063 ( .A1(n9936), .A2(n9935), .ZN(n9934) );
  OAI21_X1 U9064 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9934), .ZN(n10336) );
  NOR2_X1 U9065 ( .A1(n10337), .A2(n10336), .ZN(n7440) );
  NAND2_X1 U9066 ( .A1(n10337), .A2(n10336), .ZN(n10335) );
  OAI21_X1 U9067 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7440), .A(n10335), .ZN(
        n7444) );
  NOR2_X1 U9068 ( .A1(n7442), .A2(n7441), .ZN(n7443) );
  XNOR2_X1 U9069 ( .A(n7444), .B(n7443), .ZN(ADD_1071_U4) );
  NAND2_X1 U9070 ( .A1(n7485), .A2(n7680), .ZN(n7446) );
  NAND2_X1 U9071 ( .A1(n7694), .A2(n9089), .ZN(n7445) );
  NAND2_X1 U9072 ( .A1(n7446), .A2(n7445), .ZN(n7447) );
  XNOR2_X1 U9073 ( .A(n7447), .B(n7616), .ZN(n7449) );
  NOR2_X1 U9074 ( .A1(n7677), .A2(n7528), .ZN(n7448) );
  AOI21_X1 U9075 ( .B1(n7485), .B2(n7694), .A(n7448), .ZN(n7450) );
  NAND2_X1 U9076 ( .A1(n7449), .A2(n7450), .ZN(n7493) );
  INV_X1 U9077 ( .A(n7449), .ZN(n7452) );
  INV_X1 U9078 ( .A(n7450), .ZN(n7451) );
  NAND2_X1 U9079 ( .A1(n7452), .A2(n7451), .ZN(n7453) );
  NAND2_X1 U9080 ( .A1(n7493), .A2(n7453), .ZN(n7463) );
  NAND2_X1 U9081 ( .A1(n7455), .A2(n7454), .ZN(n7460) );
  INV_X1 U9082 ( .A(n7456), .ZN(n7457) );
  NAND2_X1 U9083 ( .A1(n7458), .A2(n7457), .ZN(n7459) );
  NAND2_X1 U9084 ( .A1(n7460), .A2(n7459), .ZN(n7461) );
  INV_X1 U9085 ( .A(n7494), .ZN(n7462) );
  AOI21_X1 U9086 ( .B1(n7463), .B2(n7461), .A(n7462), .ZN(n7469) );
  NOR2_X1 U9087 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7464), .ZN(n9623) );
  AOI21_X1 U9088 ( .B1(n8801), .B2(n9090), .A(n9623), .ZN(n7466) );
  NAND2_X1 U9089 ( .A1(n8802), .A2(n7484), .ZN(n7465) );
  OAI211_X1 U9090 ( .C1(n8805), .C2(n7542), .A(n7466), .B(n7465), .ZN(n7467)
         );
  AOI21_X1 U9091 ( .B1(n7485), .B2(n8807), .A(n7467), .ZN(n7468) );
  OAI21_X1 U9092 ( .B1(n7469), .B2(n8782), .A(n7468), .ZN(P1_U3222) );
  INV_X1 U9093 ( .A(n7470), .ZN(n7786) );
  OAI222_X1 U9094 ( .A1(P1_U3084), .A2(n5672), .B1(n9460), .B2(n7786), .C1(
        n7471), .C2(n7760), .ZN(P1_U3331) );
  INV_X1 U9095 ( .A(n7472), .ZN(n7492) );
  OR2_X1 U9096 ( .A1(n7473), .A2(P1_U3084), .ZN(n9077) );
  INV_X1 U9097 ( .A(n9077), .ZN(n9071) );
  AOI21_X1 U9098 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9463), .A(n9071), .ZN(
        n7474) );
  OAI21_X1 U9099 ( .B1(n7492), .B2(n9460), .A(n7474), .ZN(P1_U3330) );
  INV_X1 U9100 ( .A(n8893), .ZN(n7476) );
  XNOR2_X1 U9101 ( .A(n7475), .B(n7476), .ZN(n9551) );
  XNOR2_X1 U9102 ( .A(n7477), .B(n7476), .ZN(n7480) );
  OAI22_X1 U9103 ( .A1(n9500), .A2(n9502), .B1(n9501), .B2(n7542), .ZN(n7478)
         );
  INV_X1 U9104 ( .A(n7478), .ZN(n7479) );
  OAI21_X1 U9105 ( .B1(n7480), .B2(n9497), .A(n7479), .ZN(n7481) );
  AOI21_X1 U9106 ( .B1(n9551), .B2(n9506), .A(n7481), .ZN(n9553) );
  OAI21_X1 U9107 ( .B1(n7482), .B2(n9549), .A(n9751), .ZN(n7483) );
  OR2_X1 U9108 ( .A1(n7483), .A2(n7533), .ZN(n9548) );
  INV_X1 U9109 ( .A(n9515), .ZN(n7488) );
  AOI22_X1 U9110 ( .A1(n9519), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n9508), .B2(
        n7484), .ZN(n7487) );
  NAND2_X1 U9111 ( .A1(n7485), .A2(n9509), .ZN(n7486) );
  OAI211_X1 U9112 ( .C1(n9548), .C2(n7488), .A(n7487), .B(n7486), .ZN(n7489)
         );
  AOI21_X1 U9113 ( .B1(n9551), .B2(n9516), .A(n7489), .ZN(n7490) );
  OAI21_X1 U9114 ( .B1(n9553), .B2(n9312), .A(n7490), .ZN(P1_U3279) );
  NAND2_X1 U9115 ( .A1(n8654), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7491) );
  OAI211_X1 U9116 ( .C1(n7492), .C2(n8657), .A(n7491), .B(n8162), .ZN(P2_U3335) );
  NAND2_X1 U9117 ( .A1(n7537), .A2(n7680), .ZN(n7496) );
  NAND2_X1 U9118 ( .A1(n7694), .A2(n9088), .ZN(n7495) );
  NAND2_X1 U9119 ( .A1(n7496), .A2(n7495), .ZN(n7497) );
  XNOR2_X1 U9120 ( .A(n7497), .B(n7696), .ZN(n7503) );
  INV_X1 U9121 ( .A(n7503), .ZN(n7501) );
  NAND2_X1 U9122 ( .A1(n7537), .A2(n7694), .ZN(n7499) );
  NAND2_X1 U9123 ( .A1(n7693), .A2(n9088), .ZN(n7498) );
  NAND2_X1 U9124 ( .A1(n7499), .A2(n7498), .ZN(n7502) );
  INV_X1 U9125 ( .A(n7502), .ZN(n7500) );
  NAND2_X1 U9126 ( .A1(n7501), .A2(n7500), .ZN(n7612) );
  INV_X1 U9127 ( .A(n7612), .ZN(n7504) );
  AND2_X1 U9128 ( .A1(n7503), .A2(n7502), .ZN(n7611) );
  NOR2_X1 U9129 ( .A1(n7504), .A2(n7611), .ZN(n7505) );
  XNOR2_X1 U9130 ( .A(n7613), .B(n7505), .ZN(n7511) );
  INV_X1 U9131 ( .A(n7506), .ZN(n7535) );
  AND2_X1 U9132 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9637) );
  NOR2_X1 U9133 ( .A1(n8778), .A2(n7528), .ZN(n7507) );
  AOI211_X1 U9134 ( .C1(n8789), .C2(n9087), .A(n9637), .B(n7507), .ZN(n7508)
         );
  OAI21_X1 U9135 ( .B1(n8792), .B2(n7535), .A(n7508), .ZN(n7509) );
  AOI21_X1 U9136 ( .B1(n7537), .B2(n8807), .A(n7509), .ZN(n7510) );
  OAI21_X1 U9137 ( .B1(n7511), .B2(n8782), .A(n7510), .ZN(P1_U3232) );
  OR2_X1 U9138 ( .A1(n7829), .A2(n7906), .ZN(n8034) );
  AOI21_X1 U9139 ( .B1(n8136), .B2(n7513), .A(n7559), .ZN(n9904) );
  INV_X1 U9140 ( .A(n8033), .ZN(n7514) );
  XOR2_X1 U9141 ( .A(n7561), .B(n8136), .Z(n7516) );
  OAI222_X1 U9142 ( .A1(n8491), .A2(n8040), .B1(n8474), .B2(n7828), .C1(n7516), 
        .C2(n9813), .ZN(n9909) );
  INV_X1 U9143 ( .A(n7829), .ZN(n9906) );
  OR2_X1 U9144 ( .A1(n7518), .A2(n7517), .ZN(n7519) );
  INV_X1 U9145 ( .A(n7519), .ZN(n7520) );
  OAI21_X1 U9146 ( .B1(n9906), .B2(n7520), .A(n4545), .ZN(n9908) );
  NOR2_X1 U9147 ( .A1(n9908), .A2(n9836), .ZN(n7523) );
  AOI22_X1 U9148 ( .A1(n9842), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7830), .B2(
        n9838), .ZN(n7521) );
  OAI21_X1 U9149 ( .B1(n9906), .B2(n9835), .A(n7521), .ZN(n7522) );
  AOI211_X1 U9150 ( .C1(n9909), .C2(n9840), .A(n7523), .B(n7522), .ZN(n7524)
         );
  OAI21_X1 U9151 ( .B1(n9904), .B2(n8529), .A(n7524), .ZN(P2_U3284) );
  XNOR2_X1 U9152 ( .A(n7525), .B(n4727), .ZN(n9544) );
  NAND2_X1 U9153 ( .A1(n9544), .A2(n9506), .ZN(n7532) );
  OAI21_X1 U9154 ( .B1(n8895), .B2(n7527), .A(n7526), .ZN(n7530) );
  OAI22_X1 U9155 ( .A1(n7528), .A2(n9502), .B1(n9501), .B2(n9344), .ZN(n7529)
         );
  AOI21_X1 U9156 ( .B1(n7530), .B2(n9351), .A(n7529), .ZN(n7531) );
  OR2_X1 U9157 ( .A1(n7533), .A2(n9541), .ZN(n7534) );
  NAND2_X1 U9158 ( .A1(n7548), .A2(n7534), .ZN(n9542) );
  INV_X1 U9159 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9107) );
  OAI22_X1 U9160 ( .A1(n9338), .A2(n9107), .B1(n7535), .B2(n9294), .ZN(n7536)
         );
  AOI21_X1 U9161 ( .B1(n7537), .B2(n9509), .A(n7536), .ZN(n7538) );
  OAI21_X1 U9162 ( .B1(n9542), .B2(n7782), .A(n7538), .ZN(n7539) );
  AOI21_X1 U9163 ( .B1(n9544), .B2(n9516), .A(n7539), .ZN(n7540) );
  OAI21_X1 U9164 ( .B1(n9546), .B2(n9312), .A(n7540), .ZN(P1_U3278) );
  INV_X1 U9165 ( .A(n7545), .ZN(n8897) );
  XNOR2_X1 U9166 ( .A(n7541), .B(n8897), .ZN(n7544) );
  OAI22_X1 U9167 ( .A1(n7542), .A2(n9502), .B1(n9501), .B2(n9330), .ZN(n7543)
         );
  AOI21_X1 U9168 ( .B1(n7544), .B2(n9351), .A(n7543), .ZN(n9536) );
  XNOR2_X1 U9169 ( .A(n7546), .B(n7545), .ZN(n9539) );
  INV_X1 U9170 ( .A(n9340), .ZN(n7547) );
  NAND2_X1 U9171 ( .A1(n9539), .A2(n7547), .ZN(n7555) );
  INV_X1 U9172 ( .A(n7548), .ZN(n7550) );
  INV_X1 U9173 ( .A(n7549), .ZN(n9354) );
  OAI211_X1 U9174 ( .C1(n7550), .C2(n9537), .A(n9751), .B(n9354), .ZN(n9535)
         );
  INV_X1 U9175 ( .A(n9535), .ZN(n7553) );
  AOI22_X1 U9176 ( .A1(n9519), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9508), .B2(
        n8676), .ZN(n7551) );
  OAI21_X1 U9177 ( .B1(n9537), .B2(n9357), .A(n7551), .ZN(n7552) );
  AOI21_X1 U9178 ( .B1(n7553), .B2(n9515), .A(n7552), .ZN(n7554) );
  OAI211_X1 U9179 ( .C1(n9519), .C2(n9536), .A(n7555), .B(n7554), .ZN(P1_U3277) );
  INV_X1 U9180 ( .A(n7556), .ZN(n7570) );
  OAI222_X1 U9181 ( .A1(n7557), .A2(P1_U3084), .B1(n9460), .B2(n7570), .C1(
        n10223), .C2(n7760), .ZN(P1_U3329) );
  XNOR2_X1 U9182 ( .A(n8623), .B(n8040), .ZN(n8135) );
  XNOR2_X1 U9183 ( .A(n7575), .B(n8135), .ZN(n8629) );
  INV_X1 U9184 ( .A(n8623), .ZN(n7886) );
  AOI21_X1 U9185 ( .B1(n8623), .B2(n4545), .A(n7581), .ZN(n8626) );
  AOI22_X1 U9186 ( .A1(n9842), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7889), .B2(
        n9838), .ZN(n7560) );
  OAI21_X1 U9187 ( .B1(n7886), .B2(n9835), .A(n7560), .ZN(n7568) );
  AOI21_X1 U9188 ( .B1(n8135), .B2(n7562), .A(n7577), .ZN(n7563) );
  NOR2_X1 U9189 ( .A1(n7563), .A2(n9813), .ZN(n7566) );
  OR2_X1 U9190 ( .A1(n7936), .A2(n8491), .ZN(n7565) );
  OR2_X1 U9191 ( .A1(n7906), .A2(n8474), .ZN(n7564) );
  NAND2_X1 U9192 ( .A1(n7565), .A2(n7564), .ZN(n7883) );
  NOR2_X1 U9193 ( .A1(n7566), .A2(n7883), .ZN(n8628) );
  NOR2_X1 U9194 ( .A1(n8628), .A2(n9842), .ZN(n7567) );
  AOI211_X1 U9195 ( .C1(n8626), .C2(n8527), .A(n7568), .B(n7567), .ZN(n7569)
         );
  OAI21_X1 U9196 ( .B1(n8529), .B2(n8629), .A(n7569), .ZN(P2_U3283) );
  OAI222_X1 U9197 ( .A1(P2_U3152), .A2(n7571), .B1(n8661), .B2(n10120), .C1(
        n8657), .C2(n7570), .ZN(P2_U3334) );
  INV_X1 U9198 ( .A(n7572), .ZN(n7587) );
  AOI22_X1 U9199 ( .A1(n7573), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n9463), .ZN(n7574) );
  OAI21_X1 U9200 ( .B1(n7587), .B2(n9460), .A(n7574), .ZN(P1_U3328) );
  INV_X1 U9201 ( .A(n8040), .ZN(n8167) );
  OR2_X1 U9202 ( .A1(n7601), .A2(n7936), .ZN(n8045) );
  NAND2_X1 U9203 ( .A1(n7601), .A2(n7936), .ZN(n8046) );
  NAND2_X1 U9204 ( .A1(n8045), .A2(n8046), .ZN(n8043) );
  NAND2_X1 U9205 ( .A1(n7576), .A2(n8043), .ZN(n7603) );
  OAI21_X1 U9206 ( .B1(n7576), .B2(n8043), .A(n7603), .ZN(n8621) );
  INV_X1 U9207 ( .A(n8621), .ZN(n7586) );
  INV_X1 U9208 ( .A(n8043), .ZN(n8137) );
  OAI211_X1 U9209 ( .C1(n7578), .C2(n8137), .A(n7606), .B(n9857), .ZN(n7580)
         );
  AOI22_X1 U9210 ( .A1(n9807), .A2(n7604), .B1(n8167), .B2(n9806), .ZN(n7579)
         );
  NAND2_X1 U9211 ( .A1(n7580), .A2(n7579), .ZN(n8619) );
  INV_X1 U9212 ( .A(n7601), .ZN(n8617) );
  OAI21_X1 U9213 ( .B1(n7581), .B2(n8617), .A(n4480), .ZN(n8618) );
  NOR2_X1 U9214 ( .A1(n8618), .A2(n9836), .ZN(n7584) );
  AOI22_X1 U9215 ( .A1(n9842), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7800), .B2(
        n9838), .ZN(n7582) );
  OAI21_X1 U9216 ( .B1(n8617), .B2(n9835), .A(n7582), .ZN(n7583) );
  AOI211_X1 U9217 ( .C1(n8619), .C2(n9840), .A(n7584), .B(n7583), .ZN(n7585)
         );
  OAI21_X1 U9218 ( .B1(n7586), .B2(n8529), .A(n7585), .ZN(P2_U3282) );
  OAI222_X1 U9219 ( .A1(n7589), .A2(P2_U3152), .B1(n8657), .B2(n7587), .C1(
        n10104), .C2(n8661), .ZN(P2_U3333) );
  INV_X1 U9220 ( .A(n7590), .ZN(n7593) );
  AOI22_X1 U9221 ( .A1(n7591), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n9463), .ZN(n7592) );
  OAI21_X1 U9222 ( .B1(n7593), .B2(n9460), .A(n7592), .ZN(P1_U3327) );
  OAI222_X1 U9223 ( .A1(P2_U3152), .A2(n7595), .B1(n8661), .B2(n7594), .C1(
        n8657), .C2(n7593), .ZN(P2_U3332) );
  INV_X1 U9224 ( .A(n7596), .ZN(n7709) );
  NAND2_X1 U9225 ( .A1(n9463), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n7598) );
  OAI211_X1 U9226 ( .C1(n7709), .C2(n9460), .A(n7598), .B(n7597), .ZN(P1_U3326) );
  OAI222_X1 U9227 ( .A1(n8661), .A2(n7600), .B1(n8657), .B2(n7599), .C1(n8149), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  INV_X1 U9228 ( .A(n7936), .ZN(n8521) );
  NAND2_X1 U9229 ( .A1(n8612), .A2(n7849), .ZN(n8050) );
  NAND2_X1 U9230 ( .A1(n8051), .A2(n8050), .ZN(n8140) );
  OR2_X1 U9231 ( .A1(n8606), .A2(n8166), .ZN(n8056) );
  NAND2_X1 U9232 ( .A1(n8606), .A2(n8166), .ZN(n8055) );
  NAND2_X1 U9233 ( .A1(n8056), .A2(n8055), .ZN(n8510) );
  INV_X1 U9234 ( .A(n8606), .ZN(n8508) );
  NAND2_X1 U9235 ( .A1(n8603), .A2(n7918), .ZN(n8060) );
  INV_X1 U9236 ( .A(n7918), .ZN(n8503) );
  NAND2_X1 U9237 ( .A1(n8596), .A2(n8492), .ZN(n8072) );
  NAND2_X1 U9238 ( .A1(n8064), .A2(n8072), .ZN(n8285) );
  INV_X1 U9239 ( .A(n8285), .ZN(n8142) );
  XNOR2_X1 U9240 ( .A(n8286), .B(n8142), .ZN(n8600) );
  INV_X1 U9241 ( .A(n8603), .ZN(n8499) );
  AND2_X2 U9242 ( .A1(n8505), .A2(n8499), .ZN(n8493) );
  XNOR2_X1 U9243 ( .A(n8493), .B(n8596), .ZN(n8597) );
  INV_X1 U9244 ( .A(n8596), .ZN(n8284) );
  AOI22_X1 U9245 ( .A1(n9842), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n7920), .B2(
        n9838), .ZN(n7605) );
  OAI21_X1 U9246 ( .B1(n8284), .B2(n9835), .A(n7605), .ZN(n7609) );
  NAND2_X1 U9247 ( .A1(n8488), .A2(n8487), .ZN(n8486) );
  XNOR2_X1 U9248 ( .A(n7946), .B(n8285), .ZN(n7607) );
  AOI222_X1 U9249 ( .A1(n9857), .A2(n7607), .B1(n8464), .B2(n9807), .C1(n8503), 
        .C2(n9806), .ZN(n8599) );
  NOR2_X1 U9250 ( .A1(n8599), .A2(n9842), .ZN(n7608) );
  AOI211_X1 U9251 ( .C1(n8597), .C2(n8527), .A(n7609), .B(n7608), .ZN(n7610)
         );
  OAI21_X1 U9252 ( .B1(n8600), .B2(n8529), .A(n7610), .ZN(P2_U3278) );
  AOI22_X1 U9253 ( .A1(n9395), .A2(n7694), .B1(n7693), .B2(n9229), .ZN(n7663)
         );
  AOI22_X1 U9254 ( .A1(n9427), .A2(n7694), .B1(n7693), .B2(n9318), .ZN(n8717)
         );
  NAND2_X1 U9255 ( .A1(n8835), .A2(n7680), .ZN(n7615) );
  NAND2_X1 U9256 ( .A1(n7694), .A2(n9087), .ZN(n7614) );
  NAND2_X1 U9257 ( .A1(n7615), .A2(n7614), .ZN(n7617) );
  XNOR2_X1 U9258 ( .A(n7617), .B(n7616), .ZN(n7621) );
  NAND2_X1 U9259 ( .A1(n7620), .A2(n7621), .ZN(n8671) );
  NAND2_X1 U9260 ( .A1(n8835), .A2(n7694), .ZN(n7619) );
  NAND2_X1 U9261 ( .A1(n7693), .A2(n9087), .ZN(n7618) );
  NAND2_X1 U9262 ( .A1(n7619), .A2(n7618), .ZN(n8674) );
  NAND2_X1 U9263 ( .A1(n8671), .A2(n8674), .ZN(n7624) );
  INV_X1 U9264 ( .A(n7620), .ZN(n7623) );
  INV_X1 U9265 ( .A(n7621), .ZN(n7622) );
  NAND2_X1 U9266 ( .A1(n7623), .A2(n7622), .ZN(n8672) );
  NAND2_X1 U9267 ( .A1(n7624), .A2(n8672), .ZN(n7629) );
  NAND2_X1 U9268 ( .A1(n9430), .A2(n7680), .ZN(n7626) );
  NAND2_X1 U9269 ( .A1(n7694), .A2(n9086), .ZN(n7625) );
  NAND2_X1 U9270 ( .A1(n7626), .A2(n7625), .ZN(n7627) );
  XNOR2_X1 U9271 ( .A(n7627), .B(n7696), .ZN(n7628) );
  NOR2_X1 U9272 ( .A1(n7629), .A2(n7628), .ZN(n8796) );
  AOI22_X1 U9273 ( .A1(n9430), .A2(n7694), .B1(n7693), .B2(n9086), .ZN(n8799)
         );
  NAND2_X1 U9274 ( .A1(n7629), .A2(n7628), .ZN(n8797) );
  OAI21_X2 U9275 ( .B1(n8796), .B2(n8799), .A(n8797), .ZN(n8720) );
  AOI22_X1 U9276 ( .A1(n9427), .A2(n7695), .B1(n7694), .B2(n9318), .ZN(n7630)
         );
  XOR2_X1 U9277 ( .A(n7696), .B(n7630), .Z(n8718) );
  AOI22_X1 U9278 ( .A1(n9420), .A2(n7695), .B1(n7694), .B2(n9085), .ZN(n7631)
         );
  XNOR2_X1 U9279 ( .A(n7631), .B(n7696), .ZN(n7633) );
  AOI22_X1 U9280 ( .A1(n9420), .A2(n7694), .B1(n7693), .B2(n9085), .ZN(n7632)
         );
  XNOR2_X1 U9281 ( .A(n7633), .B(n7632), .ZN(n8727) );
  INV_X1 U9282 ( .A(n7632), .ZN(n7635) );
  INV_X1 U9283 ( .A(n7633), .ZN(n7634) );
  AOI22_X1 U9284 ( .A1(n9417), .A2(n7695), .B1(n7694), .B2(n10326), .ZN(n7636)
         );
  XNOR2_X1 U9285 ( .A(n7636), .B(n7696), .ZN(n7638) );
  OAI22_X1 U9286 ( .A1(n4749), .A2(n6401), .B1(n7637), .B2(n7677), .ZN(n8775)
         );
  NAND2_X1 U9287 ( .A1(n7639), .A2(n7638), .ZN(n8772) );
  OAI21_X1 U9288 ( .B1(n8774), .B2(n8775), .A(n8772), .ZN(n8694) );
  NAND2_X1 U9289 ( .A1(n9410), .A2(n7680), .ZN(n7641) );
  NAND2_X1 U9290 ( .A1(n9274), .A2(n7694), .ZN(n7640) );
  NAND2_X1 U9291 ( .A1(n7641), .A2(n7640), .ZN(n7642) );
  XNOR2_X1 U9292 ( .A(n7642), .B(n7696), .ZN(n7645) );
  NAND2_X1 U9293 ( .A1(n9410), .A2(n7694), .ZN(n7644) );
  NAND2_X1 U9294 ( .A1(n9274), .A2(n7693), .ZN(n7643) );
  NAND2_X1 U9295 ( .A1(n7644), .A2(n7643), .ZN(n7646) );
  NAND2_X1 U9296 ( .A1(n7645), .A2(n7646), .ZN(n8696) );
  NAND2_X1 U9297 ( .A1(n8694), .A2(n8696), .ZN(n8693) );
  INV_X1 U9298 ( .A(n7645), .ZN(n7648) );
  INV_X1 U9299 ( .A(n7646), .ZN(n7647) );
  NAND2_X1 U9300 ( .A1(n7648), .A2(n7647), .ZN(n8695) );
  NAND2_X1 U9301 ( .A1(n8693), .A2(n8695), .ZN(n8742) );
  NAND2_X1 U9302 ( .A1(n9405), .A2(n7680), .ZN(n7650) );
  NAND2_X1 U9303 ( .A1(n9286), .A2(n7694), .ZN(n7649) );
  NAND2_X1 U9304 ( .A1(n7650), .A2(n7649), .ZN(n7651) );
  XNOR2_X1 U9305 ( .A(n7651), .B(n7696), .ZN(n7654) );
  AOI22_X1 U9306 ( .A1(n9405), .A2(n7694), .B1(n7693), .B2(n9286), .ZN(n7652)
         );
  XNOR2_X1 U9307 ( .A(n7654), .B(n7652), .ZN(n8743) );
  INV_X1 U9308 ( .A(n7652), .ZN(n7653) );
  OR2_X1 U9309 ( .A1(n7654), .A2(n7653), .ZN(n7655) );
  INV_X1 U9310 ( .A(n9402), .ZN(n7656) );
  OAI22_X1 U9311 ( .A1(n7656), .A2(n6401), .B1(n8758), .B2(n7677), .ZN(n7660)
         );
  NAND2_X1 U9312 ( .A1(n9402), .A2(n7695), .ZN(n7658) );
  NAND2_X1 U9313 ( .A1(n9273), .A2(n7694), .ZN(n7657) );
  NAND2_X1 U9314 ( .A1(n7658), .A2(n7657), .ZN(n7659) );
  XNOR2_X1 U9315 ( .A(n7659), .B(n7696), .ZN(n7661) );
  XOR2_X1 U9316 ( .A(n7660), .B(n7661), .Z(n8704) );
  NOR2_X1 U9317 ( .A1(n7663), .A2(n7664), .ZN(n8753) );
  AOI22_X1 U9318 ( .A1(n9395), .A2(n7695), .B1(n7694), .B2(n9229), .ZN(n7662)
         );
  XOR2_X1 U9319 ( .A(n7696), .B(n7662), .Z(n8754) );
  NAND2_X1 U9320 ( .A1(n7664), .A2(n7663), .ZN(n8751) );
  AOI22_X1 U9321 ( .A1(n9390), .A2(n7695), .B1(n7694), .B2(n9242), .ZN(n7665)
         );
  XNOR2_X1 U9322 ( .A(n7665), .B(n7696), .ZN(n7666) );
  OAI22_X1 U9323 ( .A1(n9225), .A2(n6401), .B1(n9209), .B2(n7677), .ZN(n8685)
         );
  NAND2_X1 U9324 ( .A1(n9387), .A2(n7680), .ZN(n7669) );
  NAND2_X1 U9325 ( .A1(n9230), .A2(n7694), .ZN(n7668) );
  NAND2_X1 U9326 ( .A1(n7669), .A2(n7668), .ZN(n7670) );
  XNOR2_X1 U9327 ( .A(n7670), .B(n7696), .ZN(n7671) );
  AOI22_X1 U9328 ( .A1(n9387), .A2(n7694), .B1(n7693), .B2(n9230), .ZN(n7672)
         );
  XNOR2_X1 U9329 ( .A(n7671), .B(n7672), .ZN(n8735) );
  INV_X1 U9330 ( .A(n7671), .ZN(n7673) );
  NAND2_X1 U9331 ( .A1(n9382), .A2(n7680), .ZN(n7675) );
  NAND2_X1 U9332 ( .A1(n9185), .A2(n7694), .ZN(n7674) );
  NAND2_X1 U9333 ( .A1(n7675), .A2(n7674), .ZN(n7676) );
  XNOR2_X1 U9334 ( .A(n7676), .B(n7696), .ZN(n7679) );
  OAI22_X1 U9335 ( .A1(n9200), .A2(n6401), .B1(n9208), .B2(n7677), .ZN(n7678)
         );
  XNOR2_X1 U9336 ( .A(n7679), .B(n7678), .ZN(n8711) );
  NAND2_X1 U9337 ( .A1(n9375), .A2(n7680), .ZN(n7682) );
  NAND2_X1 U9338 ( .A1(n9164), .A2(n7694), .ZN(n7681) );
  NAND2_X1 U9339 ( .A1(n7682), .A2(n7681), .ZN(n7683) );
  XNOR2_X1 U9340 ( .A(n7683), .B(n7696), .ZN(n7687) );
  NAND2_X1 U9341 ( .A1(n9375), .A2(n7694), .ZN(n7685) );
  NAND2_X1 U9342 ( .A1(n9164), .A2(n7693), .ZN(n7684) );
  NAND2_X1 U9343 ( .A1(n7685), .A2(n7684), .ZN(n7686) );
  NAND2_X1 U9344 ( .A1(n7687), .A2(n7686), .ZN(n8785) );
  NOR2_X1 U9345 ( .A1(n7687), .A2(n7686), .ZN(n8784) );
  AOI21_X1 U9346 ( .B1(n8788), .B2(n8785), .A(n8784), .ZN(n8665) );
  AOI22_X1 U9347 ( .A1(n9370), .A2(n7695), .B1(n7694), .B2(n9186), .ZN(n7688)
         );
  XNOR2_X1 U9348 ( .A(n7688), .B(n7696), .ZN(n7690) );
  AOI22_X1 U9349 ( .A1(n9370), .A2(n7694), .B1(n7693), .B2(n9186), .ZN(n7689)
         );
  NAND2_X1 U9350 ( .A1(n7690), .A2(n7689), .ZN(n7691) );
  OAI21_X1 U9351 ( .B1(n7690), .B2(n7689), .A(n7691), .ZN(n8664) );
  NOR2_X1 U9352 ( .A1(n8665), .A2(n8664), .ZN(n8663) );
  INV_X1 U9353 ( .A(n7691), .ZN(n7692) );
  NOR2_X1 U9354 ( .A1(n8663), .A2(n7692), .ZN(n7701) );
  AOI22_X1 U9355 ( .A1(n7763), .A2(n7694), .B1(n7693), .B2(n9171), .ZN(n7699)
         );
  AOI22_X1 U9356 ( .A1(n7763), .A2(n7695), .B1(n7694), .B2(n9171), .ZN(n7697)
         );
  XNOR2_X1 U9357 ( .A(n7697), .B(n7696), .ZN(n7698) );
  XNOR2_X1 U9358 ( .A(n7701), .B(n7700), .ZN(n7708) );
  INV_X1 U9359 ( .A(n7702), .ZN(n9149) );
  AOI22_X1 U9360 ( .A1(n9149), .A2(n8802), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n7704) );
  NAND2_X1 U9361 ( .A1(n9084), .A2(n8789), .ZN(n7703) );
  OAI211_X1 U9362 ( .C1(n7705), .C2(n8778), .A(n7704), .B(n7703), .ZN(n7706)
         );
  AOI21_X1 U9363 ( .B1(n7763), .B2(n8807), .A(n7706), .ZN(n7707) );
  OAI21_X1 U9364 ( .B1(n7708), .B2(n8782), .A(n7707), .ZN(P1_U3218) );
  OAI222_X1 U9365 ( .A1(n8661), .A2(n7710), .B1(n8657), .B2(n7709), .C1(n6975), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  INV_X1 U9366 ( .A(SI_28_), .ZN(n7713) );
  NAND2_X1 U9367 ( .A1(n7714), .A2(n7713), .ZN(n7715) );
  INV_X1 U9368 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7719) );
  INV_X1 U9369 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7718) );
  MUX2_X1 U9370 ( .A(n7719), .B(n7718), .S(n7717), .Z(n7737) );
  INV_X1 U9371 ( .A(SI_29_), .ZN(n7720) );
  AND2_X1 U9372 ( .A1(n7737), .A2(n7720), .ZN(n7723) );
  INV_X1 U9373 ( .A(n7737), .ZN(n7721) );
  NAND2_X1 U9374 ( .A1(n7721), .A2(SI_29_), .ZN(n7722) );
  MUX2_X1 U9375 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n7727), .Z(n7724) );
  NAND2_X1 U9376 ( .A1(n7725), .A2(n7724), .ZN(n7726) );
  MUX2_X1 U9377 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7727), .Z(n7728) );
  XNOR2_X1 U9378 ( .A(n7728), .B(SI_31_), .ZN(n7729) );
  NAND2_X1 U9379 ( .A1(n7749), .A2(n7739), .ZN(n7732) );
  NAND2_X1 U9380 ( .A1(n5234), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7731) );
  NAND2_X2 U9381 ( .A1(n7732), .A2(n7731), .ZN(n8876) );
  NAND2_X1 U9382 ( .A1(n8651), .A2(n7739), .ZN(n7735) );
  NAND2_X1 U9383 ( .A1(n5234), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7734) );
  XNOR2_X1 U9384 ( .A(n7737), .B(SI_29_), .ZN(n7738) );
  NAND2_X1 U9385 ( .A1(n8653), .A2(n7739), .ZN(n7741) );
  NAND2_X1 U9386 ( .A1(n5234), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7740) );
  OR2_X2 U9387 ( .A1(n7776), .A2(n9367), .ZN(n9143) );
  XOR2_X1 U9388 ( .A(n8876), .B(n9142), .Z(n9364) );
  NOR2_X1 U9389 ( .A1(n9074), .A2(n7742), .ZN(n7743) );
  NOR2_X1 U9390 ( .A1(n9501), .A2(n7743), .ZN(n7774) );
  NAND2_X1 U9391 ( .A1(n5421), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n7746) );
  NAND2_X1 U9392 ( .A1(n7770), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n7745) );
  NAND2_X1 U9393 ( .A1(n5431), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n7744) );
  AND3_X1 U9394 ( .A1(n7746), .A2(n7745), .A3(n7744), .ZN(n8913) );
  INV_X1 U9395 ( .A(n8913), .ZN(n9082) );
  NAND2_X1 U9396 ( .A1(n7774), .A2(n9082), .ZN(n9529) );
  NOR2_X1 U9397 ( .A1(n9312), .A2(n9529), .ZN(n9145) );
  AOI21_X1 U9398 ( .B1(n9519), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9145), .ZN(
        n7748) );
  NAND2_X1 U9399 ( .A1(n8876), .A2(n9509), .ZN(n7747) );
  OAI211_X1 U9400 ( .C1(n9364), .C2(n7782), .A(n7748), .B(n7747), .ZN(P1_U3261) );
  NAND2_X1 U9401 ( .A1(n8426), .A2(n8432), .ZN(n8427) );
  OR2_X2 U9402 ( .A1(n8427), .A2(n8570), .ZN(n8414) );
  NOR2_X2 U9403 ( .A1(n8414), .A2(n8565), .ZN(n8379) );
  NAND2_X1 U9404 ( .A1(n8379), .A2(n8387), .ZN(n8380) );
  OR2_X2 U9405 ( .A1(n8380), .A2(n8557), .ZN(n8365) );
  NAND2_X1 U9406 ( .A1(n8653), .A2(n7752), .ZN(n7751) );
  NAND2_X1 U9407 ( .A1(n7753), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7750) );
  NAND2_X1 U9408 ( .A1(n7751), .A2(n7750), .ZN(n7953) );
  NAND2_X1 U9409 ( .A1(n8651), .A2(n7752), .ZN(n7755) );
  NAND2_X1 U9410 ( .A1(n7753), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n7754) );
  XOR2_X1 U9411 ( .A(n8532), .B(n8279), .Z(n8530) );
  NAND2_X1 U9412 ( .A1(n8530), .A2(n8527), .ZN(n7759) );
  AOI222_X1 U9413 ( .A1(n4463), .A2(P2_REG2_REG_31__SCAN_IN), .B1(n7955), .B2(
        P2_REG1_REG_31__SCAN_IN), .C1(n5785), .C2(P2_REG0_REG_31__SCAN_IN), 
        .ZN(n7954) );
  INV_X1 U9414 ( .A(n7954), .ZN(n8163) );
  INV_X1 U9415 ( .A(P2_B_REG_SCAN_IN), .ZN(n7756) );
  NOR2_X1 U9416 ( .A1(n6975), .A2(n7756), .ZN(n7757) );
  NOR2_X1 U9417 ( .A1(n8491), .A2(n7757), .ZN(n8316) );
  NAND2_X1 U9418 ( .A1(n8163), .A2(n8316), .ZN(n8535) );
  NOR2_X1 U9419 ( .A1(n9842), .A2(n8535), .ZN(n8281) );
  AOI21_X1 U9420 ( .B1(P2_REG2_REG_31__SCAN_IN), .B2(n9842), .A(n8281), .ZN(
        n7758) );
  OAI211_X1 U9421 ( .C1(n8532), .C2(n9835), .A(n7759), .B(n7758), .ZN(P2_U3265) );
  OAI222_X1 U9422 ( .A1(n5062), .A2(P1_U3084), .B1(n9460), .B2(n7762), .C1(
        n7761), .C2(n7760), .ZN(P1_U3332) );
  INV_X1 U9423 ( .A(n7763), .ZN(n9152) );
  NAND2_X1 U9424 ( .A1(n9367), .A2(n7766), .ZN(n8918) );
  XNOR2_X1 U9425 ( .A(n7767), .B(n9028), .ZN(n9368) );
  AND2_X1 U9426 ( .A1(n9020), .A2(n9018), .ZN(n9024) );
  INV_X1 U9427 ( .A(n8810), .ZN(n9023) );
  AOI21_X1 U9428 ( .B1(n9165), .B2(n9024), .A(n9023), .ZN(n7768) );
  XNOR2_X1 U9429 ( .A(n7768), .B(n9028), .ZN(n7769) );
  NAND2_X1 U9430 ( .A1(n5421), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7773) );
  NAND2_X1 U9431 ( .A1(n7770), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7772) );
  NAND2_X1 U9432 ( .A1(n5431), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7771) );
  NAND3_X1 U9433 ( .A1(n7773), .A2(n7772), .A3(n7771), .ZN(n9083) );
  AOI22_X1 U9434 ( .A1(n9171), .A2(n9317), .B1(n7774), .B2(n9083), .ZN(n7775)
         );
  NAND2_X1 U9435 ( .A1(n9367), .A2(n7776), .ZN(n7777) );
  OAI22_X1 U9436 ( .A1(n7779), .A2(n9294), .B1(n7778), .B2(n9338), .ZN(n7780)
         );
  AOI21_X1 U9437 ( .B1(n9367), .B2(n9509), .A(n7780), .ZN(n7781) );
  OAI21_X1 U9438 ( .B1(n9365), .B2(n7782), .A(n7781), .ZN(n7783) );
  AOI21_X1 U9439 ( .B1(n9366), .B2(n9338), .A(n7783), .ZN(n7784) );
  OAI21_X1 U9440 ( .B1(n9368), .B2(n9340), .A(n7784), .ZN(P1_U3355) );
  OAI222_X1 U9441 ( .A1(n8661), .A2(n10128), .B1(n8657), .B2(n7786), .C1(n7785), .C2(P2_U3152), .ZN(P2_U3336) );
  INV_X1 U9442 ( .A(n8550), .ZN(n8344) );
  OAI211_X1 U9443 ( .C1(n7789), .C2(n7788), .A(n7787), .B(n7924), .ZN(n7793)
         );
  NOR2_X1 U9444 ( .A1(n7909), .A2(n8346), .ZN(n7791) );
  OAI22_X1 U9445 ( .A1(n8311), .A2(n7938), .B1(n7937), .B2(n8378), .ZN(n7790)
         );
  AOI211_X1 U9446 ( .C1(P2_REG3_REG_27__SCAN_IN), .C2(P2_U3152), .A(n7791), 
        .B(n7790), .ZN(n7792) );
  OAI211_X1 U9447 ( .C1(n8344), .C2(n7933), .A(n7793), .B(n7792), .ZN(P2_U3216) );
  OAI21_X1 U9448 ( .B1(n7796), .B2(n7795), .A(n7794), .ZN(n7797) );
  NAND2_X1 U9449 ( .A1(n7797), .A2(n7924), .ZN(n7802) );
  OAI22_X1 U9450 ( .A1(n7849), .A2(n7938), .B1(n7937), .B2(n8040), .ZN(n7798)
         );
  AOI211_X1 U9451 ( .C1(n7940), .C2(n7800), .A(n7799), .B(n7798), .ZN(n7801)
         );
  OAI211_X1 U9452 ( .C1(n8617), .C2(n7933), .A(n7802), .B(n7801), .ZN(P2_U3217) );
  INV_X1 U9453 ( .A(n7803), .ZN(n7805) );
  NOR2_X1 U9454 ( .A1(n7805), .A2(n7804), .ZN(n7862) );
  AOI211_X1 U9455 ( .C1(n7805), .C2(n7804), .A(n7944), .B(n7862), .ZN(n7809)
         );
  INV_X1 U9456 ( .A(n8570), .ZN(n8418) );
  AOI22_X1 U9457 ( .A1(n7940), .A2(n8416), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n7807) );
  INV_X1 U9458 ( .A(n8377), .ZN(n8412) );
  INV_X1 U9459 ( .A(n7937), .ZN(n7875) );
  INV_X1 U9460 ( .A(n8296), .ZN(n8448) );
  AOI22_X1 U9461 ( .A1(n7913), .A2(n8412), .B1(n7875), .B2(n8448), .ZN(n7806)
         );
  OAI211_X1 U9462 ( .C1(n8418), .C2(n7933), .A(n7807), .B(n7806), .ZN(n7808)
         );
  OR2_X1 U9463 ( .A1(n7809), .A2(n7808), .ZN(P2_U3218) );
  NAND2_X1 U9464 ( .A1(n4563), .A2(n7810), .ZN(n7811) );
  XNOR2_X1 U9465 ( .A(n7812), .B(n7811), .ZN(n7813) );
  NAND2_X1 U9466 ( .A1(n7813), .A2(n7924), .ZN(n7816) );
  AND2_X1 U9467 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8275) );
  OAI22_X1 U9468 ( .A1(n8492), .A2(n7937), .B1(n7938), .B2(n8475), .ZN(n7814)
         );
  AOI211_X1 U9469 ( .C1(n7940), .C2(n8479), .A(n8275), .B(n7814), .ZN(n7815)
         );
  OAI211_X1 U9470 ( .C1(n8482), .C2(n7933), .A(n7816), .B(n7815), .ZN(P2_U3221) );
  NAND2_X1 U9471 ( .A1(n7872), .A2(n7817), .ZN(n7818) );
  NAND2_X1 U9472 ( .A1(n7818), .A2(n7819), .ZN(n7893) );
  OAI211_X1 U9473 ( .C1(n7819), .C2(n7818), .A(n7893), .B(n7924), .ZN(n7824)
         );
  NOR2_X1 U9474 ( .A1(n7820), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7822) );
  OAI22_X1 U9475 ( .A1(n8475), .A2(n7937), .B1(n7938), .B2(n8296), .ZN(n7821)
         );
  AOI211_X1 U9476 ( .C1(n7940), .C2(n8442), .A(n7822), .B(n7821), .ZN(n7823)
         );
  OAI211_X1 U9477 ( .C1(n8444), .C2(n7933), .A(n7824), .B(n7823), .ZN(P2_U3225) );
  OAI211_X1 U9478 ( .C1(n7827), .C2(n7826), .A(n7825), .B(n7924), .ZN(n7834)
         );
  INV_X1 U9479 ( .A(n7828), .ZN(n8168) );
  AOI22_X1 U9480 ( .A1(n7829), .A2(n7941), .B1(n7875), .B2(n8168), .ZN(n7833)
         );
  AOI22_X1 U9481 ( .A1(n7940), .A2(n7830), .B1(P2_REG3_REG_12__SCAN_IN), .B2(
        P2_U3152), .ZN(n7832) );
  NAND2_X1 U9482 ( .A1(n7913), .A2(n8167), .ZN(n7831) );
  NAND4_X1 U9483 ( .A1(n7834), .A2(n7833), .A3(n7832), .A4(n7831), .ZN(
        P2_U3226) );
  OAI211_X1 U9484 ( .C1(n7837), .C2(n7836), .A(n7835), .B(n7924), .ZN(n7841)
         );
  NOR2_X1 U9485 ( .A1(n7909), .A2(n8383), .ZN(n7839) );
  OAI22_X1 U9486 ( .A1(n8377), .A2(n7937), .B1(n7938), .B2(n8378), .ZN(n7838)
         );
  AOI211_X1 U9487 ( .C1(P2_REG3_REG_25__SCAN_IN), .C2(P2_U3152), .A(n7839), 
        .B(n7838), .ZN(n7840) );
  OAI211_X1 U9488 ( .C1(n8387), .C2(n7933), .A(n7841), .B(n7840), .ZN(P2_U3227) );
  XNOR2_X1 U9489 ( .A(n7842), .B(n7843), .ZN(n7935) );
  INV_X1 U9490 ( .A(n7842), .ZN(n7844) );
  AOI22_X1 U9491 ( .A1(n7935), .A2(n7934), .B1(n7844), .B2(n7843), .ZN(n7848)
         );
  NAND2_X1 U9492 ( .A1(n7846), .A2(n7845), .ZN(n7847) );
  XNOR2_X1 U9493 ( .A(n7848), .B(n7847), .ZN(n7853) );
  AND2_X1 U9494 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8211) );
  OAI22_X1 U9495 ( .A1(n7849), .A2(n7937), .B1(n7938), .B2(n7918), .ZN(n7850)
         );
  AOI211_X1 U9496 ( .C1(n7940), .C2(n8506), .A(n8211), .B(n7850), .ZN(n7852)
         );
  NAND2_X1 U9497 ( .A1(n7941), .A2(n8606), .ZN(n7851) );
  OAI211_X1 U9498 ( .C1(n7853), .C2(n7944), .A(n7852), .B(n7851), .ZN(P2_U3228) );
  XNOR2_X1 U9499 ( .A(n7855), .B(n7854), .ZN(n7860) );
  INV_X1 U9500 ( .A(n8496), .ZN(n7856) );
  OAI22_X1 U9501 ( .A1(n7909), .A2(n7856), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8230), .ZN(n7858) );
  OAI22_X1 U9502 ( .A1(n8166), .A2(n7937), .B1(n7938), .B2(n8492), .ZN(n7857)
         );
  AOI211_X1 U9503 ( .C1(n8603), .C2(n7941), .A(n7858), .B(n7857), .ZN(n7859)
         );
  OAI21_X1 U9504 ( .B1(n7860), .B2(n7944), .A(n7859), .ZN(P2_U3230) );
  NOR2_X1 U9505 ( .A1(n7862), .A2(n7861), .ZN(n7864) );
  XNOR2_X1 U9506 ( .A(n7864), .B(n7863), .ZN(n7866) );
  AOI21_X1 U9507 ( .B1(n7866), .B2(n7867), .A(n7944), .ZN(n7865) );
  OAI21_X1 U9508 ( .B1(n7867), .B2(n7866), .A(n7865), .ZN(n7871) );
  NOR2_X1 U9509 ( .A1(n7909), .A2(n8394), .ZN(n7869) );
  INV_X1 U9510 ( .A(n8436), .ZN(n8403) );
  OAI22_X1 U9511 ( .A1(n8403), .A2(n7937), .B1(n7938), .B2(n8404), .ZN(n7868)
         );
  AOI211_X1 U9512 ( .C1(P2_REG3_REG_24__SCAN_IN), .C2(P2_U3152), .A(n7869), 
        .B(n7868), .ZN(n7870) );
  OAI211_X1 U9513 ( .C1(n8397), .C2(n7933), .A(n7871), .B(n7870), .ZN(P2_U3231) );
  OAI211_X1 U9514 ( .C1(n7874), .C2(n7873), .A(n7872), .B(n7924), .ZN(n7879)
         );
  AOI22_X1 U9515 ( .A1(n7940), .A2(n8456), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n7878) );
  INV_X1 U9516 ( .A(n8294), .ZN(n8463) );
  AOI22_X1 U9517 ( .A1(n7913), .A2(n8463), .B1(n7875), .B2(n8464), .ZN(n7877)
         );
  NAND2_X1 U9518 ( .A1(n8586), .A2(n7941), .ZN(n7876) );
  NAND4_X1 U9519 ( .A1(n7879), .A2(n7878), .A3(n7877), .A4(n7876), .ZN(
        P2_U3235) );
  NOR2_X1 U9520 ( .A1(n4560), .A2(n7880), .ZN(n7881) );
  XNOR2_X1 U9521 ( .A(n7882), .B(n7881), .ZN(n7891) );
  INV_X1 U9522 ( .A(n7883), .ZN(n7885) );
  OAI21_X1 U9523 ( .B1(n7929), .B2(n7885), .A(n7884), .ZN(n7888) );
  NOR2_X1 U9524 ( .A1(n7933), .A2(n7886), .ZN(n7887) );
  AOI211_X1 U9525 ( .C1(n7940), .C2(n7889), .A(n7888), .B(n7887), .ZN(n7890)
         );
  OAI21_X1 U9526 ( .B1(n7891), .B2(n7944), .A(n7890), .ZN(P2_U3236) );
  NAND2_X1 U9527 ( .A1(n7893), .A2(n7892), .ZN(n7897) );
  XNOR2_X1 U9528 ( .A(n7895), .B(n7894), .ZN(n7896) );
  XNOR2_X1 U9529 ( .A(n7897), .B(n7896), .ZN(n7902) );
  INV_X1 U9530 ( .A(n8430), .ZN(n7898) );
  OAI22_X1 U9531 ( .A1(n7909), .A2(n7898), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10204), .ZN(n7900) );
  OAI22_X1 U9532 ( .A1(n8403), .A2(n7938), .B1(n7937), .B2(n8294), .ZN(n7899)
         );
  AOI211_X1 U9533 ( .C1(n8576), .C2(n7941), .A(n7900), .B(n7899), .ZN(n7901)
         );
  OAI21_X1 U9534 ( .B1(n7902), .B2(n7944), .A(n7901), .ZN(P2_U3237) );
  OAI211_X1 U9535 ( .C1(n7905), .C2(n7904), .A(n7903), .B(n7924), .ZN(n7915)
         );
  INV_X1 U9536 ( .A(n7907), .ZN(n7908) );
  OAI22_X1 U9537 ( .A1(n7909), .A2(n7908), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5937), .ZN(n7912) );
  OAI22_X1 U9538 ( .A1(n9899), .A2(n7933), .B1(n7937), .B2(n7910), .ZN(n7911)
         );
  AOI211_X1 U9539 ( .C1(n7913), .C2(n7558), .A(n7912), .B(n7911), .ZN(n7914)
         );
  NAND2_X1 U9540 ( .A1(n7915), .A2(n7914), .ZN(P2_U3238) );
  XNOR2_X1 U9541 ( .A(n7917), .B(n7916), .ZN(n7923) );
  AND2_X1 U9542 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8249) );
  OAI22_X1 U9543 ( .A1(n7918), .A2(n7937), .B1(n7938), .B2(n8287), .ZN(n7919)
         );
  AOI211_X1 U9544 ( .C1(n7940), .C2(n7920), .A(n8249), .B(n7919), .ZN(n7922)
         );
  NAND2_X1 U9545 ( .A1(n8596), .A2(n7941), .ZN(n7921) );
  OAI211_X1 U9546 ( .C1(n7923), .C2(n7944), .A(n7922), .B(n7921), .ZN(P2_U3240) );
  INV_X1 U9547 ( .A(n8557), .ZN(n8370) );
  OAI211_X1 U9548 ( .C1(n7927), .C2(n7926), .A(n7925), .B(n7924), .ZN(n7932)
         );
  INV_X1 U9549 ( .A(n8309), .ZN(n8334) );
  INV_X1 U9550 ( .A(n8404), .ZN(n8165) );
  AOI22_X1 U9551 ( .A1(n8334), .A2(n9807), .B1(n9806), .B2(n8165), .ZN(n8363)
         );
  OAI22_X1 U9552 ( .A1(n7929), .A2(n8363), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7928), .ZN(n7930) );
  AOI21_X1 U9553 ( .B1(n8367), .B2(n7940), .A(n7930), .ZN(n7931) );
  OAI211_X1 U9554 ( .C1(n8370), .C2(n7933), .A(n7932), .B(n7931), .ZN(P2_U3242) );
  XNOR2_X1 U9555 ( .A(n7935), .B(n7934), .ZN(n7945) );
  AND2_X1 U9556 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8196) );
  OAI22_X1 U9557 ( .A1(n8166), .A2(n7938), .B1(n7937), .B2(n7936), .ZN(n7939)
         );
  AOI211_X1 U9558 ( .C1(n7940), .C2(n8517), .A(n8196), .B(n7939), .ZN(n7943)
         );
  NAND2_X1 U9559 ( .A1(n7941), .A2(n8612), .ZN(n7942) );
  OAI211_X1 U9560 ( .C1(n7945), .C2(n7944), .A(n7943), .B(n7942), .ZN(P2_U3243) );
  NAND2_X1 U9561 ( .A1(n7946), .A2(n8142), .ZN(n7947) );
  NAND2_X1 U9562 ( .A1(n7947), .A2(n8064), .ZN(n8472) );
  OR2_X1 U9563 ( .A1(n8593), .A2(n8287), .ZN(n8074) );
  NAND2_X1 U9564 ( .A1(n8593), .A2(n8287), .ZN(n8460) );
  NAND2_X1 U9565 ( .A1(n8074), .A2(n8460), .ZN(n8471) );
  NAND2_X1 U9566 ( .A1(n8586), .A2(n8475), .ZN(n8076) );
  NAND2_X1 U9567 ( .A1(n8079), .A2(n8076), .ZN(n8454) );
  INV_X1 U9568 ( .A(n8454), .ZN(n8461) );
  NAND2_X1 U9569 ( .A1(n8581), .A2(n8294), .ZN(n8433) );
  NAND2_X1 U9570 ( .A1(n8078), .A2(n8433), .ZN(n8445) );
  NAND2_X1 U9571 ( .A1(n8576), .A2(n8296), .ZN(n8083) );
  NAND2_X1 U9572 ( .A1(n8070), .A2(n8083), .ZN(n8435) );
  INV_X1 U9573 ( .A(n8433), .ZN(n7949) );
  NAND2_X1 U9574 ( .A1(n8565), .A2(n8377), .ZN(n8089) );
  INV_X1 U9575 ( .A(n8399), .ZN(n7950) );
  AND2_X1 U9576 ( .A1(n8570), .A2(n8403), .ZN(n7973) );
  NOR2_X1 U9577 ( .A1(n7950), .A2(n7973), .ZN(n7951) );
  NAND2_X1 U9578 ( .A1(n8410), .A2(n7951), .ZN(n8398) );
  NAND2_X1 U9579 ( .A1(n8562), .A2(n8404), .ZN(n7970) );
  NAND2_X1 U9580 ( .A1(n7972), .A2(n7970), .ZN(n8303) );
  NAND2_X1 U9581 ( .A1(n8557), .A2(n8378), .ZN(n8350) );
  NAND2_X1 U9582 ( .A1(n8550), .A2(n8309), .ZN(n8097) );
  NAND2_X1 U9583 ( .A1(n8098), .A2(n8097), .ZN(n8308) );
  NAND2_X1 U9584 ( .A1(n8351), .A2(n5038), .ZN(n7952) );
  NAND2_X1 U9585 ( .A1(n8545), .A2(n8311), .ZN(n7969) );
  OR2_X1 U9586 ( .A1(n7953), .A2(n8164), .ZN(n8104) );
  NAND2_X1 U9587 ( .A1(n7953), .A2(n8164), .ZN(n8105) );
  NAND2_X1 U9588 ( .A1(n8104), .A2(n8105), .ZN(n8313) );
  INV_X1 U9589 ( .A(n8313), .ZN(n8102) );
  INV_X1 U9590 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n7958) );
  NAND2_X1 U9591 ( .A1(n5785), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n7957) );
  NAND2_X1 U9592 ( .A1(n7955), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n7956) );
  OAI211_X1 U9593 ( .C1(n7959), .C2(n7958), .A(n7957), .B(n7956), .ZN(n8315)
         );
  INV_X1 U9594 ( .A(n8315), .ZN(n7960) );
  OR2_X1 U9595 ( .A1(n8280), .A2(n7960), .ZN(n8146) );
  NAND2_X1 U9596 ( .A1(n8532), .A2(n8163), .ZN(n8113) );
  NAND2_X1 U9597 ( .A1(n8280), .A2(n7960), .ZN(n8107) );
  NAND2_X1 U9598 ( .A1(n8113), .A2(n8107), .ZN(n8108) );
  AOI21_X1 U9599 ( .B1(n7961), .B2(n8146), .A(n8108), .ZN(n7962) );
  AOI21_X1 U9600 ( .B1(n7963), .B2(n7962), .A(n4855), .ZN(n7964) );
  XNOR2_X1 U9601 ( .A(n7964), .B(n8149), .ZN(n8158) );
  NAND2_X1 U9602 ( .A1(n7966), .A2(n7965), .ZN(n8157) );
  INV_X1 U9603 ( .A(n8146), .ZN(n8111) );
  MUX2_X1 U9604 ( .A(n7969), .B(n7968), .S(n8112), .Z(n8101) );
  AND2_X1 U9605 ( .A1(n8350), .A2(n7970), .ZN(n7971) );
  MUX2_X1 U9606 ( .A(n7972), .B(n7971), .S(n8112), .Z(n8093) );
  OAI21_X1 U9607 ( .B1(n8403), .B2(n8570), .A(n8399), .ZN(n7975) );
  INV_X1 U9608 ( .A(n7973), .ZN(n8400) );
  NAND2_X1 U9609 ( .A1(n8089), .A2(n8400), .ZN(n7974) );
  MUX2_X1 U9610 ( .A(n7975), .B(n7974), .S(n8112), .Z(n7976) );
  INV_X1 U9611 ( .A(n7976), .ZN(n8087) );
  NAND2_X1 U9612 ( .A1(n7997), .A2(n7999), .ZN(n7978) );
  NAND2_X1 U9613 ( .A1(n7981), .A2(n7980), .ZN(n7977) );
  MUX2_X1 U9614 ( .A(n7978), .B(n7977), .S(n8103), .Z(n8002) );
  AND2_X1 U9615 ( .A1(n7980), .A2(n7979), .ZN(n7982) );
  OAI211_X1 U9616 ( .C1(n8002), .C2(n7982), .A(n8006), .B(n7981), .ZN(n7983)
         );
  NAND2_X1 U9617 ( .A1(n7983), .A2(n8112), .ZN(n7991) );
  INV_X1 U9618 ( .A(n8002), .ZN(n7989) );
  AND2_X1 U9619 ( .A1(n8123), .A2(n5748), .ZN(n7985) );
  OAI211_X1 U9620 ( .C1(n8127), .C2(n7985), .A(n7984), .B(n8124), .ZN(n7986)
         );
  NAND3_X1 U9621 ( .A1(n7986), .A2(n7994), .A3(n8112), .ZN(n7987) );
  NAND3_X1 U9622 ( .A1(n7989), .A2(n7988), .A3(n7987), .ZN(n7990) );
  NAND2_X1 U9623 ( .A1(n8124), .A2(n8123), .ZN(n7992) );
  NAND3_X1 U9624 ( .A1(n7994), .A2(n7993), .A3(n7992), .ZN(n7995) );
  NAND3_X1 U9625 ( .A1(n7995), .A2(n8103), .A3(n7984), .ZN(n7996) );
  AND2_X1 U9626 ( .A1(n7998), .A2(n7997), .ZN(n8001) );
  OAI211_X1 U9627 ( .C1(n8002), .C2(n8001), .A(n8000), .B(n7999), .ZN(n8003)
         );
  NAND3_X1 U9628 ( .A1(n8005), .A2(n8004), .A3(n8112), .ZN(n8008) );
  NOR2_X1 U9629 ( .A1(n8006), .A2(n8112), .ZN(n8007) );
  AOI21_X1 U9630 ( .B1(n8009), .B2(n8008), .A(n8007), .ZN(n8011) );
  OAI22_X1 U9631 ( .A1(n8011), .A2(n9804), .B1(n8103), .B2(n8010), .ZN(n8013)
         );
  NAND3_X1 U9632 ( .A1(n9805), .A2(n9872), .A3(n8103), .ZN(n8012) );
  NAND2_X1 U9633 ( .A1(n8013), .A2(n8012), .ZN(n8017) );
  MUX2_X1 U9634 ( .A(n8015), .B(n8014), .S(n8112), .Z(n8016) );
  NAND3_X1 U9635 ( .A1(n8017), .A2(n8018), .A3(n8016), .ZN(n8024) );
  NAND2_X1 U9636 ( .A1(n8018), .A2(n8026), .ZN(n8019) );
  MUX2_X1 U9637 ( .A(n8020), .B(n8019), .S(n8112), .Z(n8022) );
  INV_X1 U9638 ( .A(n8025), .ZN(n8021) );
  NOR2_X1 U9639 ( .A1(n8022), .A2(n8021), .ZN(n8023) );
  NAND2_X1 U9640 ( .A1(n8033), .A2(n8025), .ZN(n8028) );
  NAND2_X1 U9641 ( .A1(n8031), .A2(n8026), .ZN(n8027) );
  MUX2_X1 U9642 ( .A(n8028), .B(n8027), .S(n8103), .Z(n8029) );
  INV_X1 U9643 ( .A(n8029), .ZN(n8030) );
  NAND2_X1 U9644 ( .A1(n8035), .A2(n8031), .ZN(n8032) );
  NAND2_X1 U9645 ( .A1(n8032), .A2(n8034), .ZN(n8038) );
  NAND2_X1 U9646 ( .A1(n8034), .A2(n8033), .ZN(n8036) );
  NAND2_X1 U9647 ( .A1(n8036), .A2(n8035), .ZN(n8037) );
  MUX2_X1 U9648 ( .A(n8038), .B(n8037), .S(n8103), .Z(n8039) );
  NOR2_X1 U9649 ( .A1(n8623), .A2(n8112), .ZN(n8042) );
  AND2_X1 U9650 ( .A1(n8623), .A2(n8112), .ZN(n8041) );
  MUX2_X1 U9651 ( .A(n8042), .B(n8041), .S(n8040), .Z(n8044) );
  MUX2_X1 U9652 ( .A(n8046), .B(n8045), .S(n8112), .Z(n8047) );
  NAND2_X1 U9653 ( .A1(n8048), .A2(n8047), .ZN(n8049) );
  NAND2_X1 U9654 ( .A1(n8049), .A2(n4772), .ZN(n8054) );
  INV_X1 U9655 ( .A(n8510), .ZN(n8053) );
  MUX2_X1 U9656 ( .A(n8051), .B(n8050), .S(n8103), .Z(n8052) );
  NAND3_X1 U9657 ( .A1(n8054), .A2(n8053), .A3(n8052), .ZN(n8058) );
  MUX2_X1 U9658 ( .A(n8056), .B(n8055), .S(n8112), .Z(n8057) );
  NAND3_X1 U9659 ( .A1(n8058), .A2(n8487), .A3(n8057), .ZN(n8063) );
  AND2_X1 U9660 ( .A1(n8064), .A2(n8059), .ZN(n8061) );
  MUX2_X1 U9661 ( .A(n8061), .B(n8060), .S(n8103), .Z(n8062) );
  NAND2_X1 U9662 ( .A1(n8063), .A2(n8062), .ZN(n8073) );
  INV_X1 U9663 ( .A(n8072), .ZN(n8065) );
  OAI211_X1 U9664 ( .C1(n8073), .C2(n8065), .A(n8064), .B(n8074), .ZN(n8066)
         );
  NAND2_X1 U9665 ( .A1(n8066), .A2(n8460), .ZN(n8067) );
  NAND2_X1 U9666 ( .A1(n8067), .A2(n8079), .ZN(n8068) );
  NAND3_X1 U9667 ( .A1(n8068), .A2(n8076), .A3(n8433), .ZN(n8069) );
  NAND3_X1 U9668 ( .A1(n8069), .A2(n8103), .A3(n8078), .ZN(n8071) );
  MUX2_X1 U9669 ( .A(n8103), .B(n8071), .S(n8070), .Z(n8085) );
  NAND2_X1 U9670 ( .A1(n8073), .A2(n8072), .ZN(n8075) );
  NAND2_X1 U9671 ( .A1(n8075), .A2(n8074), .ZN(n8077) );
  NAND3_X1 U9672 ( .A1(n8077), .A2(n8076), .A3(n8460), .ZN(n8080) );
  NAND3_X1 U9673 ( .A1(n8080), .A2(n8079), .A3(n8078), .ZN(n8081) );
  NAND3_X1 U9674 ( .A1(n8081), .A2(n8083), .A3(n8433), .ZN(n8082) );
  MUX2_X1 U9675 ( .A(n8083), .B(n8082), .S(n8112), .Z(n8084) );
  NAND3_X1 U9676 ( .A1(n8085), .A2(n8422), .A3(n8084), .ZN(n8086) );
  NAND2_X1 U9677 ( .A1(n8087), .A2(n8086), .ZN(n8091) );
  MUX2_X1 U9678 ( .A(n8089), .B(n8088), .S(n8112), .Z(n8090) );
  NAND3_X1 U9679 ( .A1(n8091), .A2(n8374), .A3(n8090), .ZN(n8092) );
  NAND3_X1 U9680 ( .A1(n8093), .A2(n8094), .A3(n8092), .ZN(n8096) );
  MUX2_X1 U9681 ( .A(n8350), .B(n8094), .S(n8112), .Z(n8095) );
  NAND3_X1 U9682 ( .A1(n8096), .A2(n8352), .A3(n8095), .ZN(n8100) );
  MUX2_X1 U9683 ( .A(n8098), .B(n8097), .S(n8112), .Z(n8099) );
  MUX2_X1 U9684 ( .A(n8105), .B(n8104), .S(n8103), .Z(n8106) );
  INV_X1 U9685 ( .A(n8108), .ZN(n8148) );
  MUX2_X1 U9686 ( .A(n8148), .B(n8109), .S(n8112), .Z(n8110) );
  MUX2_X1 U9687 ( .A(n4857), .B(n8113), .S(n8112), .Z(n8114) );
  NAND2_X1 U9688 ( .A1(n8115), .A2(n8114), .ZN(n8116) );
  INV_X1 U9689 ( .A(n8151), .ZN(n8117) );
  INV_X1 U9690 ( .A(n8118), .ZN(n8121) );
  NAND4_X1 U9691 ( .A1(n8122), .A2(n8121), .A3(n8120), .A4(n8119), .ZN(n8128)
         );
  NAND3_X1 U9692 ( .A1(n8124), .A2(n8123), .A3(n8152), .ZN(n8125) );
  NOR4_X1 U9693 ( .A1(n8128), .A2(n8127), .A3(n8126), .A4(n8125), .ZN(n8130)
         );
  NAND3_X1 U9694 ( .A1(n8130), .A2(n9793), .A3(n8129), .ZN(n8134) );
  NOR4_X1 U9695 ( .A1(n8134), .A2(n8133), .A3(n8132), .A4(n8131), .ZN(n8138)
         );
  NAND4_X1 U9696 ( .A1(n8138), .A2(n8137), .A3(n8136), .A4(n5010), .ZN(n8139)
         );
  NOR4_X1 U9697 ( .A1(n4770), .A2(n8510), .A3(n8140), .A4(n8139), .ZN(n8141)
         );
  NAND4_X1 U9698 ( .A1(n8461), .A2(n8142), .A3(n7948), .A4(n8141), .ZN(n8143)
         );
  NOR4_X1 U9699 ( .A1(n8299), .A2(n8435), .A3(n8445), .A4(n8143), .ZN(n8144)
         );
  NAND4_X1 U9700 ( .A1(n8352), .A2(n8374), .A3(n8399), .A4(n8144), .ZN(n8145)
         );
  NOR4_X1 U9701 ( .A1(n8313), .A2(n8331), .A3(n8145), .A4(n8362), .ZN(n8147)
         );
  NAND4_X1 U9702 ( .A1(n8148), .A2(n8147), .A3(n8146), .A4(n4857), .ZN(n8150)
         );
  XNOR2_X1 U9703 ( .A(n8150), .B(n8149), .ZN(n8153) );
  OAI22_X1 U9704 ( .A1(n8153), .A2(n5748), .B1(n8152), .B2(n8151), .ZN(n8154)
         );
  NAND2_X1 U9705 ( .A1(n8155), .A2(n8154), .ZN(n8156) );
  NOR4_X1 U9706 ( .A1(n9844), .A2(n8474), .A3(n6975), .A4(n8159), .ZN(n8161)
         );
  OAI21_X1 U9707 ( .B1(n8162), .B2(n5747), .A(P2_B_REG_SCAN_IN), .ZN(n8160) );
  MUX2_X1 U9708 ( .A(n8163), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8176), .Z(
        P2_U3583) );
  MUX2_X1 U9709 ( .A(n8315), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8176), .Z(
        P2_U3582) );
  INV_X1 U9710 ( .A(n8164), .ZN(n8333) );
  MUX2_X1 U9711 ( .A(n8333), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8176), .Z(
        P2_U3581) );
  INV_X1 U9712 ( .A(n8311), .ZN(n8354) );
  MUX2_X1 U9713 ( .A(n8354), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8176), .Z(
        P2_U3580) );
  MUX2_X1 U9714 ( .A(n8334), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8176), .Z(
        P2_U3579) );
  INV_X1 U9715 ( .A(n8378), .ZN(n8355) );
  MUX2_X1 U9716 ( .A(n8355), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8176), .Z(
        P2_U3578) );
  MUX2_X1 U9717 ( .A(n8165), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8176), .Z(
        P2_U3577) );
  MUX2_X1 U9718 ( .A(n8412), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8176), .Z(
        P2_U3576) );
  MUX2_X1 U9719 ( .A(n8436), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8176), .Z(
        P2_U3575) );
  MUX2_X1 U9720 ( .A(n8448), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8176), .Z(
        P2_U3574) );
  MUX2_X1 U9721 ( .A(n8463), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8176), .Z(
        P2_U3573) );
  INV_X1 U9722 ( .A(n8475), .ZN(n8447) );
  MUX2_X1 U9723 ( .A(n8447), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8176), .Z(
        P2_U3572) );
  MUX2_X1 U9724 ( .A(n8464), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8176), .Z(
        P2_U3571) );
  MUX2_X1 U9725 ( .A(n8503), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8176), .Z(
        P2_U3569) );
  INV_X1 U9726 ( .A(n8166), .ZN(n8522) );
  MUX2_X1 U9727 ( .A(n8522), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8176), .Z(
        P2_U3568) );
  MUX2_X1 U9728 ( .A(n7604), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8176), .Z(
        P2_U3567) );
  MUX2_X1 U9729 ( .A(n8521), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8176), .Z(
        P2_U3566) );
  MUX2_X1 U9730 ( .A(n8167), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8176), .Z(
        P2_U3565) );
  MUX2_X1 U9731 ( .A(n7558), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8176), .Z(
        P2_U3564) );
  MUX2_X1 U9732 ( .A(n8168), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8176), .Z(
        P2_U3563) );
  MUX2_X1 U9733 ( .A(n8169), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8176), .Z(
        P2_U3562) );
  MUX2_X1 U9734 ( .A(n9808), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8176), .Z(
        P2_U3561) );
  MUX2_X1 U9735 ( .A(n8170), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8176), .Z(
        P2_U3560) );
  MUX2_X1 U9736 ( .A(n9805), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8176), .Z(
        P2_U3559) );
  MUX2_X1 U9737 ( .A(n8171), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8176), .Z(
        P2_U3558) );
  MUX2_X1 U9738 ( .A(n8172), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8176), .Z(
        P2_U3557) );
  MUX2_X1 U9739 ( .A(n8173), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8176), .Z(
        P2_U3556) );
  MUX2_X1 U9740 ( .A(n8174), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8176), .Z(
        P2_U3555) );
  MUX2_X1 U9741 ( .A(n8175), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8176), .Z(
        P2_U3554) );
  MUX2_X1 U9742 ( .A(n6626), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8176), .Z(
        P2_U3553) );
  MUX2_X1 U9743 ( .A(n8177), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8176), .Z(
        P2_U3552) );
  OAI21_X1 U9744 ( .B1(n8180), .B2(n8179), .A(n8178), .ZN(n8181) );
  NAND2_X1 U9745 ( .A1(n9782), .A2(n8181), .ZN(n8190) );
  NOR2_X1 U9746 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5937), .ZN(n8182) );
  AOI21_X1 U9747 ( .B1(n9788), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8182), .ZN(
        n8189) );
  NAND2_X1 U9748 ( .A1(n9483), .A2(n8183), .ZN(n8188) );
  OAI211_X1 U9749 ( .C1(n8186), .C2(n8185), .A(n9783), .B(n8184), .ZN(n8187)
         );
  NAND4_X1 U9750 ( .A1(n8190), .A2(n8189), .A3(n8188), .A4(n8187), .ZN(
        P2_U3256) );
  XNOR2_X1 U9751 ( .A(n8214), .B(n8206), .ZN(n8194) );
  INV_X1 U9752 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8193) );
  NAND2_X1 U9753 ( .A1(n8194), .A2(n8193), .ZN(n8216) );
  OAI21_X1 U9754 ( .B1(n8194), .B2(n8193), .A(n8216), .ZN(n8195) );
  NAND2_X1 U9755 ( .A1(n8195), .A2(n9782), .ZN(n8204) );
  AOI21_X1 U9756 ( .B1(n9788), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8196), .ZN(
        n8203) );
  AOI21_X1 U9757 ( .B1(n8199), .B2(n8198), .A(n8197), .ZN(n8205) );
  XNOR2_X1 U9758 ( .A(n8205), .B(n8215), .ZN(n8200) );
  NAND2_X1 U9759 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8200), .ZN(n8207) );
  OAI211_X1 U9760 ( .C1(n8200), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9783), .B(
        n8207), .ZN(n8202) );
  NAND2_X1 U9761 ( .A1(n9483), .A2(n8206), .ZN(n8201) );
  NAND4_X1 U9762 ( .A1(n8204), .A2(n8203), .A3(n8202), .A4(n8201), .ZN(
        P2_U3260) );
  NAND2_X1 U9763 ( .A1(n8206), .A2(n8205), .ZN(n8208) );
  NAND2_X1 U9764 ( .A1(n8208), .A2(n8207), .ZN(n8210) );
  XNOR2_X1 U9765 ( .A(n8232), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8209) );
  NOR2_X1 U9766 ( .A1(n8209), .A2(n8210), .ZN(n8233) );
  AOI21_X1 U9767 ( .B1(n8210), .B2(n8209), .A(n8233), .ZN(n8225) );
  INV_X1 U9768 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8213) );
  INV_X1 U9769 ( .A(n8211), .ZN(n8212) );
  OAI21_X1 U9770 ( .B1(n8277), .B2(n8213), .A(n8212), .ZN(n8222) );
  NAND2_X1 U9771 ( .A1(n8215), .A2(n8214), .ZN(n8217) );
  NAND2_X1 U9772 ( .A1(n8217), .A2(n8216), .ZN(n8220) );
  NAND2_X1 U9773 ( .A1(n8232), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8218) );
  OAI21_X1 U9774 ( .B1(n8232), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8218), .ZN(
        n8219) );
  NOR2_X1 U9775 ( .A1(n8219), .A2(n8220), .ZN(n8226) );
  AOI211_X1 U9776 ( .C1(n8220), .C2(n8219), .A(n8226), .B(n9786), .ZN(n8221)
         );
  AOI211_X1 U9777 ( .C1(n9483), .C2(n8232), .A(n8222), .B(n8221), .ZN(n8223)
         );
  OAI21_X1 U9778 ( .B1(n8225), .B2(n8224), .A(n8223), .ZN(P2_U3261) );
  NAND2_X1 U9779 ( .A1(n8253), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8227) );
  OAI21_X1 U9780 ( .B1(n8253), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8227), .ZN(
        n8228) );
  AOI211_X1 U9781 ( .C1(n8229), .C2(n8228), .A(n8252), .B(n9786), .ZN(n8241)
         );
  NOR2_X1 U9782 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8230), .ZN(n8231) );
  AOI21_X1 U9783 ( .B1(n9788), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8231), .ZN(
        n8239) );
  INV_X1 U9784 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8245) );
  XNOR2_X1 U9785 ( .A(n8253), .B(n8245), .ZN(n8237) );
  OR2_X1 U9786 ( .A1(n8232), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8235) );
  INV_X1 U9787 ( .A(n8233), .ZN(n8234) );
  AND2_X1 U9788 ( .A1(n8235), .A2(n8234), .ZN(n8236) );
  NAND2_X1 U9789 ( .A1(n8237), .A2(n8236), .ZN(n8243) );
  OAI211_X1 U9790 ( .C1(n8237), .C2(n8236), .A(n9783), .B(n8243), .ZN(n8238)
         );
  OAI211_X1 U9791 ( .C1(n9785), .C2(n8244), .A(n8239), .B(n8238), .ZN(n8240)
         );
  OR2_X1 U9792 ( .A1(n8241), .A2(n8240), .ZN(P2_U3262) );
  OR2_X1 U9793 ( .A1(n8261), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8266) );
  NAND2_X1 U9794 ( .A1(n8261), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8242) );
  NAND2_X1 U9795 ( .A1(n8266), .A2(n8242), .ZN(n8247) );
  OAI21_X1 U9796 ( .B1(n8245), .B2(n8244), .A(n8243), .ZN(n8246) );
  NOR2_X1 U9797 ( .A1(n8247), .A2(n8246), .ZN(n8268) );
  AND2_X1 U9798 ( .A1(n8247), .A2(n8246), .ZN(n8248) );
  OAI21_X1 U9799 ( .B1(n8268), .B2(n8248), .A(n9783), .ZN(n8251) );
  INV_X1 U9800 ( .A(n8249), .ZN(n8250) );
  OAI211_X1 U9801 ( .C1(n8277), .C2(n10337), .A(n8251), .B(n8250), .ZN(n8260)
         );
  INV_X1 U9802 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8258) );
  INV_X1 U9803 ( .A(n8261), .ZN(n8254) );
  AOI21_X1 U9804 ( .B1(n8255), .B2(n8254), .A(n8264), .ZN(n8256) );
  INV_X1 U9805 ( .A(n8256), .ZN(n8257) );
  AOI211_X1 U9806 ( .C1(n8258), .C2(n8257), .A(n8263), .B(n9786), .ZN(n8259)
         );
  AOI211_X1 U9807 ( .C1(n9483), .C2(n8261), .A(n8260), .B(n8259), .ZN(n8262)
         );
  INV_X1 U9808 ( .A(n8262), .ZN(P2_U3263) );
  INV_X1 U9809 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8278) );
  NOR2_X1 U9810 ( .A1(n8264), .A2(n8263), .ZN(n8265) );
  XNOR2_X1 U9811 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8265), .ZN(n8271) );
  INV_X1 U9812 ( .A(n8266), .ZN(n8267) );
  NOR2_X1 U9813 ( .A1(n8268), .A2(n8267), .ZN(n8269) );
  XNOR2_X1 U9814 ( .A(n8269), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8272) );
  INV_X1 U9815 ( .A(n8272), .ZN(n8270) );
  AOI22_X1 U9816 ( .A1(n8271), .A2(n9782), .B1(n8270), .B2(n9783), .ZN(n8274)
         );
  INV_X1 U9817 ( .A(n8275), .ZN(n8276) );
  INV_X1 U9818 ( .A(n8280), .ZN(n8537) );
  INV_X1 U9819 ( .A(n8279), .ZN(n8534) );
  NAND2_X1 U9820 ( .A1(n4495), .A2(n8280), .ZN(n8533) );
  NAND3_X1 U9821 ( .A1(n8534), .A2(n8527), .A3(n8533), .ZN(n8283) );
  AOI21_X1 U9822 ( .B1(n9842), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8281), .ZN(
        n8282) );
  OAI211_X1 U9823 ( .C1(n8537), .C2(n9835), .A(n8283), .B(n8282), .ZN(P2_U3266) );
  NAND2_X1 U9824 ( .A1(n8482), .A2(n8287), .ZN(n8288) );
  NAND2_X1 U9825 ( .A1(n8469), .A2(n8288), .ZN(n8290) );
  NAND2_X1 U9826 ( .A1(n8593), .A2(n8464), .ZN(n8289) );
  NAND2_X1 U9827 ( .A1(n8290), .A2(n8289), .ZN(n8453) );
  NAND2_X1 U9828 ( .A1(n8453), .A2(n8454), .ZN(n8292) );
  NAND2_X1 U9829 ( .A1(n8586), .A2(n8447), .ZN(n8291) );
  NOR2_X1 U9830 ( .A1(n8444), .A2(n8294), .ZN(n8293) );
  NAND2_X1 U9831 ( .A1(n8444), .A2(n8294), .ZN(n8295) );
  NAND2_X1 U9832 ( .A1(n8432), .A2(n8296), .ZN(n8297) );
  NAND2_X1 U9833 ( .A1(n8298), .A2(n8297), .ZN(n8421) );
  INV_X1 U9834 ( .A(n8421), .ZN(n8300) );
  NAND2_X1 U9835 ( .A1(n8300), .A2(n8299), .ZN(n8420) );
  NAND2_X1 U9836 ( .A1(n8570), .A2(n8436), .ZN(n8301) );
  NAND2_X1 U9837 ( .A1(n8397), .A2(n8377), .ZN(n8302) );
  NAND2_X1 U9838 ( .A1(n8373), .A2(n8303), .ZN(n8305) );
  NAND2_X1 U9839 ( .A1(n8387), .A2(n8404), .ZN(n8304) );
  NAND2_X1 U9840 ( .A1(n8305), .A2(n8304), .ZN(n8359) );
  NAND2_X1 U9841 ( .A1(n8359), .A2(n8362), .ZN(n8307) );
  NAND2_X1 U9842 ( .A1(n8370), .A2(n8378), .ZN(n8306) );
  NAND2_X1 U9843 ( .A1(n8307), .A2(n8306), .ZN(n8341) );
  NAND2_X1 U9844 ( .A1(n8344), .A2(n8309), .ZN(n8310) );
  XNOR2_X1 U9845 ( .A(n8312), .B(n8313), .ZN(n8538) );
  INV_X1 U9846 ( .A(n8538), .ZN(n8324) );
  XNOR2_X1 U9847 ( .A(n8314), .B(n8313), .ZN(n8318) );
  AOI22_X1 U9848 ( .A1(n8354), .A2(n9806), .B1(n8316), .B2(n8315), .ZN(n8317)
         );
  OAI21_X1 U9849 ( .B1(n8318), .B2(n9813), .A(n8317), .ZN(n8542) );
  OAI21_X1 U9850 ( .B1(n8327), .B2(n8539), .A(n4495), .ZN(n8540) );
  NOR2_X1 U9851 ( .A1(n8540), .A2(n9836), .ZN(n8322) );
  AOI22_X1 U9852 ( .A1(n9842), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8319), .B2(
        n9838), .ZN(n8320) );
  OAI21_X1 U9853 ( .B1(n8539), .B2(n9835), .A(n8320), .ZN(n8321) );
  AOI211_X1 U9854 ( .C1(n8542), .C2(n9840), .A(n8322), .B(n8321), .ZN(n8323)
         );
  OAI21_X1 U9855 ( .B1(n8324), .B2(n8529), .A(n8323), .ZN(P2_U3267) );
  XNOR2_X1 U9856 ( .A(n8326), .B(n8325), .ZN(n8549) );
  AOI21_X1 U9857 ( .B1(n8545), .B2(n8342), .A(n8327), .ZN(n8546) );
  AOI22_X1 U9858 ( .A1(n9842), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8328), .B2(
        n9838), .ZN(n8329) );
  OAI21_X1 U9859 ( .B1(n4688), .B2(n9835), .A(n8329), .ZN(n8330) );
  AOI21_X1 U9860 ( .B1(n8546), .B2(n8527), .A(n8330), .ZN(n8340) );
  XNOR2_X1 U9861 ( .A(n8332), .B(n8331), .ZN(n8338) );
  NAND2_X1 U9862 ( .A1(n8334), .A2(n9806), .ZN(n8335) );
  OR2_X1 U9863 ( .A1(n8548), .A2(n9842), .ZN(n8339) );
  OAI211_X1 U9864 ( .C1(n8549), .C2(n8529), .A(n8340), .B(n8339), .ZN(P2_U3268) );
  XNOR2_X1 U9865 ( .A(n8341), .B(n8352), .ZN(n8554) );
  INV_X1 U9866 ( .A(n8342), .ZN(n8343) );
  AOI21_X1 U9867 ( .B1(n8550), .B2(n8365), .A(n8343), .ZN(n8551) );
  NOR2_X1 U9868 ( .A1(n8344), .A2(n9835), .ZN(n8349) );
  OAI22_X1 U9869 ( .A1(n9840), .A2(n8347), .B1(n8346), .B2(n8345), .ZN(n8348)
         );
  AOI211_X1 U9870 ( .C1(n8551), .C2(n8527), .A(n8349), .B(n8348), .ZN(n8358)
         );
  NAND2_X1 U9871 ( .A1(n8351), .A2(n8350), .ZN(n8353) );
  XNOR2_X1 U9872 ( .A(n8353), .B(n8352), .ZN(n8356) );
  AOI222_X1 U9873 ( .A1(n9857), .A2(n8356), .B1(n8355), .B2(n9806), .C1(n8354), 
        .C2(n9807), .ZN(n8553) );
  OR2_X1 U9874 ( .A1(n8553), .A2(n9842), .ZN(n8357) );
  OAI211_X1 U9875 ( .C1(n8554), .C2(n8529), .A(n8358), .B(n8357), .ZN(P2_U3269) );
  XOR2_X1 U9876 ( .A(n8362), .B(n8359), .Z(n8559) );
  OAI21_X1 U9877 ( .B1(n8364), .B2(n9813), .A(n8363), .ZN(n8555) );
  INV_X1 U9878 ( .A(n8365), .ZN(n8366) );
  AOI211_X1 U9879 ( .C1(n8557), .C2(n8380), .A(n9907), .B(n8366), .ZN(n8556)
         );
  NAND2_X1 U9880 ( .A1(n8556), .A2(n8495), .ZN(n8369) );
  AOI22_X1 U9881 ( .A1(n9842), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8367), .B2(
        n9838), .ZN(n8368) );
  OAI211_X1 U9882 ( .C1(n8370), .C2(n9835), .A(n8369), .B(n8368), .ZN(n8371)
         );
  AOI21_X1 U9883 ( .B1(n8555), .B2(n9840), .A(n8371), .ZN(n8372) );
  OAI21_X1 U9884 ( .B1(n8559), .B2(n8529), .A(n8372), .ZN(P2_U3270) );
  XNOR2_X1 U9885 ( .A(n8373), .B(n8374), .ZN(n8564) );
  XNOR2_X1 U9886 ( .A(n8375), .B(n8374), .ZN(n8376) );
  OAI222_X1 U9887 ( .A1(n8491), .A2(n8378), .B1(n8474), .B2(n8377), .C1(n9813), 
        .C2(n8376), .ZN(n8560) );
  INV_X1 U9888 ( .A(n8379), .ZN(n8382) );
  INV_X1 U9889 ( .A(n8380), .ZN(n8381) );
  AOI211_X1 U9890 ( .C1(n8562), .C2(n8382), .A(n9907), .B(n8381), .ZN(n8561)
         );
  NAND2_X1 U9891 ( .A1(n8561), .A2(n8495), .ZN(n8386) );
  INV_X1 U9892 ( .A(n8383), .ZN(n8384) );
  AOI22_X1 U9893 ( .A1(n9842), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8384), .B2(
        n9838), .ZN(n8385) );
  OAI211_X1 U9894 ( .C1(n8387), .C2(n9835), .A(n8386), .B(n8385), .ZN(n8388)
         );
  AOI21_X1 U9895 ( .B1(n8560), .B2(n9840), .A(n8388), .ZN(n8389) );
  OAI21_X1 U9896 ( .B1(n8564), .B2(n8529), .A(n8389), .ZN(P2_U3271) );
  INV_X1 U9897 ( .A(n8391), .ZN(n8392) );
  AOI21_X1 U9898 ( .B1(n8399), .B2(n8393), .A(n8392), .ZN(n8569) );
  XNOR2_X1 U9899 ( .A(n8414), .B(n8397), .ZN(n8566) );
  INV_X1 U9900 ( .A(n8394), .ZN(n8395) );
  AOI22_X1 U9901 ( .A1(n9842), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8395), .B2(
        n9838), .ZN(n8396) );
  OAI21_X1 U9902 ( .B1(n8397), .B2(n9835), .A(n8396), .ZN(n8408) );
  INV_X1 U9903 ( .A(n8398), .ZN(n8402) );
  AOI21_X1 U9904 ( .B1(n8410), .B2(n8400), .A(n8399), .ZN(n8401) );
  NOR3_X1 U9905 ( .A1(n8402), .A2(n8401), .A3(n9813), .ZN(n8406) );
  OAI22_X1 U9906 ( .A1(n8404), .A2(n8491), .B1(n8403), .B2(n8474), .ZN(n8405)
         );
  NOR2_X1 U9907 ( .A1(n8406), .A2(n8405), .ZN(n8568) );
  NOR2_X1 U9908 ( .A1(n8568), .A2(n9842), .ZN(n8407) );
  AOI211_X1 U9909 ( .C1(n8566), .C2(n8527), .A(n8408), .B(n8407), .ZN(n8409)
         );
  OAI21_X1 U9910 ( .B1(n8569), .B2(n8529), .A(n8409), .ZN(P2_U3272) );
  OAI21_X1 U9911 ( .B1(n8411), .B2(n8422), .A(n8410), .ZN(n8413) );
  AOI222_X1 U9912 ( .A1(n9857), .A2(n8413), .B1(n8448), .B2(n9806), .C1(n8412), 
        .C2(n9807), .ZN(n8575) );
  INV_X1 U9913 ( .A(n8414), .ZN(n8415) );
  AOI21_X1 U9914 ( .B1(n8570), .B2(n8427), .A(n8415), .ZN(n8571) );
  AOI22_X1 U9915 ( .A1(n9842), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8416), .B2(
        n9838), .ZN(n8417) );
  OAI21_X1 U9916 ( .B1(n8418), .B2(n9835), .A(n8417), .ZN(n8419) );
  AOI21_X1 U9917 ( .B1(n8571), .B2(n8527), .A(n8419), .ZN(n8424) );
  NAND2_X1 U9918 ( .A1(n8421), .A2(n8422), .ZN(n8572) );
  NAND3_X1 U9919 ( .A1(n8420), .A2(n8572), .A3(n8512), .ZN(n8423) );
  OAI211_X1 U9920 ( .C1(n8575), .C2(n9842), .A(n8424), .B(n8423), .ZN(P2_U3273) );
  XOR2_X1 U9921 ( .A(n8425), .B(n8435), .Z(n8580) );
  INV_X1 U9922 ( .A(n8426), .ZN(n8429) );
  INV_X1 U9923 ( .A(n8427), .ZN(n8428) );
  AOI21_X1 U9924 ( .B1(n8576), .B2(n8429), .A(n8428), .ZN(n8577) );
  AOI22_X1 U9925 ( .A1(n9842), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8430), .B2(
        n9838), .ZN(n8431) );
  OAI21_X1 U9926 ( .B1(n8432), .B2(n9835), .A(n8431), .ZN(n8439) );
  NAND2_X1 U9927 ( .A1(n8446), .A2(n8433), .ZN(n8434) );
  XOR2_X1 U9928 ( .A(n8435), .B(n8434), .Z(n8437) );
  AOI222_X1 U9929 ( .A1(n9857), .A2(n8437), .B1(n8463), .B2(n9806), .C1(n8436), 
        .C2(n9807), .ZN(n8579) );
  NOR2_X1 U9930 ( .A1(n8579), .A2(n9842), .ZN(n8438) );
  AOI211_X1 U9931 ( .C1(n8577), .C2(n8527), .A(n8439), .B(n8438), .ZN(n8440)
         );
  OAI21_X1 U9932 ( .B1(n8580), .B2(n8529), .A(n8440), .ZN(P2_U3274) );
  XNOR2_X1 U9933 ( .A(n8441), .B(n8445), .ZN(n8585) );
  XNOR2_X1 U9934 ( .A(n8455), .B(n8581), .ZN(n8582) );
  AOI22_X1 U9935 ( .A1(n9842), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8442), .B2(
        n9838), .ZN(n8443) );
  OAI21_X1 U9936 ( .B1(n8444), .B2(n9835), .A(n8443), .ZN(n8451) );
  OAI21_X1 U9937 ( .B1(n4499), .B2(n4646), .A(n8446), .ZN(n8449) );
  AOI222_X1 U9938 ( .A1(n9857), .A2(n8449), .B1(n8448), .B2(n9807), .C1(n8447), 
        .C2(n9806), .ZN(n8584) );
  NOR2_X1 U9939 ( .A1(n8584), .A2(n9842), .ZN(n8450) );
  AOI211_X1 U9940 ( .C1(n8582), .C2(n8527), .A(n8451), .B(n8450), .ZN(n8452)
         );
  OAI21_X1 U9941 ( .B1(n8529), .B2(n8585), .A(n8452), .ZN(P2_U3275) );
  XNOR2_X1 U9942 ( .A(n8453), .B(n8454), .ZN(n8590) );
  AOI21_X1 U9943 ( .B1(n8586), .B2(n8476), .A(n8455), .ZN(n8587) );
  INV_X1 U9944 ( .A(n8586), .ZN(n8458) );
  AOI22_X1 U9945 ( .A1(n9842), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8456), .B2(
        n9838), .ZN(n8457) );
  OAI21_X1 U9946 ( .B1(n8458), .B2(n9835), .A(n8457), .ZN(n8467) );
  NAND2_X1 U9947 ( .A1(n8459), .A2(n8460), .ZN(n8462) );
  XNOR2_X1 U9948 ( .A(n8462), .B(n8461), .ZN(n8465) );
  AOI222_X1 U9949 ( .A1(n9857), .A2(n8465), .B1(n8464), .B2(n9806), .C1(n8463), 
        .C2(n9807), .ZN(n8589) );
  NOR2_X1 U9950 ( .A1(n8589), .A2(n9842), .ZN(n8466) );
  AOI211_X1 U9951 ( .C1(n8587), .C2(n8527), .A(n8467), .B(n8466), .ZN(n8468)
         );
  OAI21_X1 U9952 ( .B1(n8529), .B2(n8590), .A(n8468), .ZN(P2_U3276) );
  XNOR2_X1 U9953 ( .A(n8469), .B(n8471), .ZN(n8595) );
  INV_X1 U9954 ( .A(n8459), .ZN(n8470) );
  AOI21_X1 U9955 ( .B1(n8472), .B2(n8471), .A(n8470), .ZN(n8473) );
  OAI222_X1 U9956 ( .A1(n8491), .A2(n8475), .B1(n8474), .B2(n8492), .C1(n9813), 
        .C2(n8473), .ZN(n8591) );
  INV_X1 U9957 ( .A(n8476), .ZN(n8477) );
  AOI211_X1 U9958 ( .C1(n8593), .C2(n8478), .A(n9907), .B(n8477), .ZN(n8592)
         );
  NAND2_X1 U9959 ( .A1(n8592), .A2(n8495), .ZN(n8481) );
  AOI22_X1 U9960 ( .A1(n9842), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8479), .B2(
        n9838), .ZN(n8480) );
  OAI211_X1 U9961 ( .C1(n8482), .C2(n9835), .A(n8481), .B(n8480), .ZN(n8483)
         );
  AOI21_X1 U9962 ( .B1(n8591), .B2(n9840), .A(n8483), .ZN(n8484) );
  OAI21_X1 U9963 ( .B1(n8595), .B2(n8529), .A(n8484), .ZN(P2_U3277) );
  XNOR2_X1 U9964 ( .A(n8485), .B(n4770), .ZN(n8605) );
  OAI211_X1 U9965 ( .C1(n8488), .C2(n8487), .A(n8486), .B(n9857), .ZN(n8490)
         );
  NAND2_X1 U9966 ( .A1(n8522), .A2(n9806), .ZN(n8489) );
  OAI211_X1 U9967 ( .C1(n8492), .C2(n8491), .A(n8490), .B(n8489), .ZN(n8601)
         );
  INV_X1 U9968 ( .A(n8505), .ZN(n8494) );
  AOI211_X1 U9969 ( .C1(n8603), .C2(n8494), .A(n9907), .B(n8493), .ZN(n8602)
         );
  NAND2_X1 U9970 ( .A1(n8602), .A2(n8495), .ZN(n8498) );
  AOI22_X1 U9971 ( .A1(n9842), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8496), .B2(
        n9838), .ZN(n8497) );
  OAI211_X1 U9972 ( .C1(n8499), .C2(n9835), .A(n8498), .B(n8497), .ZN(n8500)
         );
  AOI21_X1 U9973 ( .B1(n8601), .B2(n9840), .A(n8500), .ZN(n8501) );
  OAI21_X1 U9974 ( .B1(n8605), .B2(n8529), .A(n8501), .ZN(P2_U3279) );
  XNOR2_X1 U9975 ( .A(n8502), .B(n8510), .ZN(n8504) );
  AOI222_X1 U9976 ( .A1(n9857), .A2(n8504), .B1(n8503), .B2(n9807), .C1(n7604), 
        .C2(n9806), .ZN(n8611) );
  AOI21_X1 U9977 ( .B1(n8606), .B2(n8516), .A(n8505), .ZN(n8607) );
  AOI22_X1 U9978 ( .A1(n9842), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8506), .B2(
        n9838), .ZN(n8507) );
  OAI21_X1 U9979 ( .B1(n8508), .B2(n9835), .A(n8507), .ZN(n8509) );
  AOI21_X1 U9980 ( .B1(n8607), .B2(n8527), .A(n8509), .ZN(n8514) );
  OR2_X1 U9981 ( .A1(n4557), .A2(n8510), .ZN(n8608) );
  NAND3_X1 U9982 ( .A1(n8608), .A2(n8511), .A3(n8512), .ZN(n8513) );
  OAI211_X1 U9983 ( .C1(n8611), .C2(n9842), .A(n8514), .B(n8513), .ZN(P2_U3280) );
  XNOR2_X1 U9984 ( .A(n8515), .B(n4772), .ZN(n8616) );
  AOI21_X1 U9985 ( .B1(n8612), .B2(n4480), .A(n4681), .ZN(n8613) );
  AOI22_X1 U9986 ( .A1(n9842), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8517), .B2(
        n9838), .ZN(n8518) );
  OAI21_X1 U9987 ( .B1(n4685), .B2(n9835), .A(n8518), .ZN(n8526) );
  OAI211_X1 U9988 ( .C1(n8520), .C2(n4772), .A(n8519), .B(n9857), .ZN(n8524)
         );
  AOI22_X1 U9989 ( .A1(n9807), .A2(n8522), .B1(n8521), .B2(n9806), .ZN(n8523)
         );
  AND2_X1 U9990 ( .A1(n8524), .A2(n8523), .ZN(n8615) );
  NOR2_X1 U9991 ( .A1(n8615), .A2(n9842), .ZN(n8525) );
  AOI211_X1 U9992 ( .C1(n8613), .C2(n8527), .A(n8526), .B(n8525), .ZN(n8528)
         );
  OAI21_X1 U9993 ( .B1(n8616), .B2(n8529), .A(n8528), .ZN(P2_U3281) );
  NAND2_X1 U9994 ( .A1(n8530), .A2(n8625), .ZN(n8531) );
  OAI211_X1 U9995 ( .C1(n8532), .C2(n9905), .A(n8531), .B(n8535), .ZN(n8630)
         );
  MUX2_X1 U9996 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8630), .S(n9927), .Z(
        P2_U3551) );
  NAND3_X1 U9997 ( .A1(n8534), .A2(n8625), .A3(n8533), .ZN(n8536) );
  OAI211_X1 U9998 ( .C1(n8537), .C2(n9905), .A(n8536), .B(n8535), .ZN(n8631)
         );
  MUX2_X1 U9999 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8631), .S(n9927), .Z(
        P2_U3550) );
  NAND2_X1 U10000 ( .A1(n8538), .A2(n9912), .ZN(n8544) );
  OAI22_X1 U10001 ( .A1(n8540), .A2(n9907), .B1(n8539), .B2(n9905), .ZN(n8541)
         );
  NOR2_X1 U10002 ( .A1(n8542), .A2(n8541), .ZN(n8543) );
  NAND2_X1 U10003 ( .A1(n8544), .A2(n8543), .ZN(n8632) );
  MUX2_X1 U10004 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8632), .S(n9927), .Z(
        P2_U3549) );
  AOI22_X1 U10005 ( .A1(n8546), .A2(n8625), .B1(n8624), .B2(n8545), .ZN(n8547)
         );
  OAI211_X1 U10006 ( .C1(n8549), .C2(n9864), .A(n8548), .B(n8547), .ZN(n8633)
         );
  MUX2_X1 U10007 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8633), .S(n9927), .Z(
        P2_U3548) );
  AOI22_X1 U10008 ( .A1(n8551), .A2(n8625), .B1(n8624), .B2(n8550), .ZN(n8552)
         );
  OAI211_X1 U10009 ( .C1(n8554), .C2(n9864), .A(n8553), .B(n8552), .ZN(n8634)
         );
  MUX2_X1 U10010 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8634), .S(n9927), .Z(
        P2_U3547) );
  AOI211_X1 U10011 ( .C1(n8624), .C2(n8557), .A(n8556), .B(n8555), .ZN(n8558)
         );
  OAI21_X1 U10012 ( .B1(n9864), .B2(n8559), .A(n8558), .ZN(n8635) );
  MUX2_X1 U10013 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8635), .S(n9927), .Z(
        P2_U3546) );
  AOI211_X1 U10014 ( .C1(n8624), .C2(n8562), .A(n8561), .B(n8560), .ZN(n8563)
         );
  OAI21_X1 U10015 ( .B1(n9864), .B2(n8564), .A(n8563), .ZN(n8636) );
  MUX2_X1 U10016 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8636), .S(n9927), .Z(
        P2_U3545) );
  AOI22_X1 U10017 ( .A1(n8566), .A2(n8625), .B1(n8624), .B2(n8565), .ZN(n8567)
         );
  OAI211_X1 U10018 ( .C1(n8569), .C2(n9864), .A(n8568), .B(n8567), .ZN(n8637)
         );
  MUX2_X1 U10019 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8637), .S(n9927), .Z(
        P2_U3544) );
  AOI22_X1 U10020 ( .A1(n8571), .A2(n8625), .B1(n8624), .B2(n8570), .ZN(n8574)
         );
  NAND3_X1 U10021 ( .A1(n8420), .A2(n8572), .A3(n9912), .ZN(n8573) );
  NAND3_X1 U10022 ( .A1(n8575), .A2(n8574), .A3(n8573), .ZN(n8638) );
  MUX2_X1 U10023 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8638), .S(n9927), .Z(
        P2_U3543) );
  AOI22_X1 U10024 ( .A1(n8577), .A2(n8625), .B1(n8624), .B2(n8576), .ZN(n8578)
         );
  OAI211_X1 U10025 ( .C1(n8580), .C2(n9864), .A(n8579), .B(n8578), .ZN(n8639)
         );
  MUX2_X1 U10026 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8639), .S(n9927), .Z(
        P2_U3542) );
  AOI22_X1 U10027 ( .A1(n8582), .A2(n8625), .B1(n8624), .B2(n8581), .ZN(n8583)
         );
  OAI211_X1 U10028 ( .C1(n9864), .C2(n8585), .A(n8584), .B(n8583), .ZN(n8640)
         );
  MUX2_X1 U10029 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8640), .S(n9927), .Z(
        P2_U3541) );
  AOI22_X1 U10030 ( .A1(n8587), .A2(n8625), .B1(n8624), .B2(n8586), .ZN(n8588)
         );
  OAI211_X1 U10031 ( .C1(n9864), .C2(n8590), .A(n8589), .B(n8588), .ZN(n8641)
         );
  MUX2_X1 U10032 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8641), .S(n9927), .Z(
        P2_U3540) );
  AOI211_X1 U10033 ( .C1(n8624), .C2(n8593), .A(n8592), .B(n8591), .ZN(n8594)
         );
  OAI21_X1 U10034 ( .B1(n9864), .B2(n8595), .A(n8594), .ZN(n8642) );
  MUX2_X1 U10035 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8642), .S(n9927), .Z(
        P2_U3539) );
  AOI22_X1 U10036 ( .A1(n8597), .A2(n8625), .B1(n8624), .B2(n8596), .ZN(n8598)
         );
  OAI211_X1 U10037 ( .C1(n9864), .C2(n8600), .A(n8599), .B(n8598), .ZN(n8643)
         );
  MUX2_X1 U10038 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8643), .S(n9927), .Z(
        P2_U3538) );
  AOI211_X1 U10039 ( .C1(n8624), .C2(n8603), .A(n8602), .B(n8601), .ZN(n8604)
         );
  OAI21_X1 U10040 ( .B1(n9864), .B2(n8605), .A(n8604), .ZN(n8644) );
  MUX2_X1 U10041 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8644), .S(n9927), .Z(
        P2_U3537) );
  AOI22_X1 U10042 ( .A1(n8607), .A2(n8625), .B1(n8624), .B2(n8606), .ZN(n8610)
         );
  NAND3_X1 U10043 ( .A1(n8608), .A2(n8511), .A3(n9912), .ZN(n8609) );
  NAND3_X1 U10044 ( .A1(n8611), .A2(n8610), .A3(n8609), .ZN(n8645) );
  MUX2_X1 U10045 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8645), .S(n9927), .Z(
        P2_U3536) );
  AOI22_X1 U10046 ( .A1(n8613), .A2(n8625), .B1(n8624), .B2(n8612), .ZN(n8614)
         );
  OAI211_X1 U10047 ( .C1(n8616), .C2(n9864), .A(n8615), .B(n8614), .ZN(n8646)
         );
  MUX2_X1 U10048 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8646), .S(n9927), .Z(
        P2_U3535) );
  OAI22_X1 U10049 ( .A1(n8618), .A2(n9907), .B1(n8617), .B2(n9905), .ZN(n8620)
         );
  AOI211_X1 U10050 ( .C1(n9912), .C2(n8621), .A(n8620), .B(n8619), .ZN(n8622)
         );
  INV_X1 U10051 ( .A(n8622), .ZN(n8647) );
  MUX2_X1 U10052 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8647), .S(n9927), .Z(
        P2_U3534) );
  AOI22_X1 U10053 ( .A1(n8626), .A2(n8625), .B1(n8624), .B2(n8623), .ZN(n8627)
         );
  OAI211_X1 U10054 ( .C1(n9864), .C2(n8629), .A(n8628), .B(n8627), .ZN(n8648)
         );
  MUX2_X1 U10055 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8648), .S(n9927), .Z(
        P2_U3533) );
  MUX2_X1 U10056 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8630), .S(n9915), .Z(
        P2_U3519) );
  MUX2_X1 U10057 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8631), .S(n9915), .Z(
        P2_U3518) );
  MUX2_X1 U10058 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8632), .S(n9915), .Z(
        P2_U3517) );
  MUX2_X1 U10059 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8633), .S(n9915), .Z(
        P2_U3516) );
  MUX2_X1 U10060 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8634), .S(n9915), .Z(
        P2_U3515) );
  MUX2_X1 U10061 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8635), .S(n9915), .Z(
        P2_U3514) );
  MUX2_X1 U10062 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8636), .S(n9915), .Z(
        P2_U3513) );
  MUX2_X1 U10063 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8637), .S(n9915), .Z(
        P2_U3512) );
  MUX2_X1 U10064 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8638), .S(n9915), .Z(
        P2_U3511) );
  MUX2_X1 U10065 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8639), .S(n9915), .Z(
        P2_U3510) );
  MUX2_X1 U10066 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8640), .S(n9915), .Z(
        P2_U3509) );
  MUX2_X1 U10067 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8641), .S(n9915), .Z(
        P2_U3508) );
  MUX2_X1 U10068 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8642), .S(n9915), .Z(
        P2_U3507) );
  MUX2_X1 U10069 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8643), .S(n9915), .Z(
        P2_U3505) );
  MUX2_X1 U10070 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8644), .S(n9915), .Z(
        P2_U3502) );
  MUX2_X1 U10071 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8645), .S(n9915), .Z(
        P2_U3499) );
  MUX2_X1 U10072 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8646), .S(n9915), .Z(
        P2_U3496) );
  MUX2_X1 U10073 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8647), .S(n9915), .Z(
        P2_U3493) );
  MUX2_X1 U10074 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8648), .S(n9915), .Z(
        P2_U3490) );
  INV_X1 U10075 ( .A(n7749), .ZN(n9455) );
  NOR4_X1 U10076 ( .A1(n4793), .A2(P2_IR_REG_30__SCAN_IN), .A3(n5721), .A4(
        P2_U3152), .ZN(n8649) );
  AOI21_X1 U10077 ( .B1(n8654), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8649), .ZN(
        n8650) );
  OAI21_X1 U10078 ( .B1(n9455), .B2(n8657), .A(n8650), .ZN(P2_U3327) );
  INV_X1 U10079 ( .A(n8651), .ZN(n9457) );
  AOI22_X1 U10080 ( .A1(n5727), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8654), .ZN(n8652) );
  OAI21_X1 U10081 ( .B1(n9457), .B2(n8657), .A(n8652), .ZN(P2_U3328) );
  INV_X1 U10082 ( .A(n8653), .ZN(n9461) );
  AOI22_X1 U10083 ( .A1(n8655), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n8654), .ZN(n8656) );
  OAI21_X1 U10084 ( .B1(n9461), .B2(n8657), .A(n8656), .ZN(P2_U3329) );
  NAND2_X1 U10085 ( .A1(n9462), .A2(n8658), .ZN(n8660) );
  OAI211_X1 U10086 ( .C1(n8661), .C2(n10118), .A(n8660), .B(n8659), .ZN(
        P2_U3330) );
  MUX2_X1 U10087 ( .A(n8662), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  AOI21_X1 U10088 ( .B1(n8665), .B2(n8664), .A(n8663), .ZN(n8670) );
  NAND2_X1 U10089 ( .A1(n9171), .A2(n8789), .ZN(n8667) );
  AOI22_X1 U10090 ( .A1(n9161), .A2(n8802), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n8666) );
  OAI211_X1 U10091 ( .C1(n9195), .C2(n8778), .A(n8667), .B(n8666), .ZN(n8668)
         );
  AOI21_X1 U10092 ( .B1(n9370), .B2(n8807), .A(n8668), .ZN(n8669) );
  OAI21_X1 U10093 ( .B1(n8670), .B2(n8782), .A(n8669), .ZN(P1_U3212) );
  NAND2_X1 U10094 ( .A1(n8671), .A2(n8672), .ZN(n8673) );
  XOR2_X1 U10095 ( .A(n8674), .B(n8673), .Z(n8681) );
  NOR2_X1 U10096 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8675), .ZN(n9650) );
  AOI21_X1 U10097 ( .B1(n8801), .B2(n9088), .A(n9650), .ZN(n8678) );
  NAND2_X1 U10098 ( .A1(n8802), .A2(n8676), .ZN(n8677) );
  OAI211_X1 U10099 ( .C1(n8805), .C2(n9330), .A(n8678), .B(n8677), .ZN(n8679)
         );
  AOI21_X1 U10100 ( .B1(n8835), .B2(n8807), .A(n8679), .ZN(n8680) );
  OAI21_X1 U10101 ( .B1(n8681), .B2(n8782), .A(n8680), .ZN(P1_U3213) );
  INV_X1 U10102 ( .A(n8682), .ZN(n8683) );
  NOR2_X1 U10103 ( .A1(n8684), .A2(n8683), .ZN(n8686) );
  XNOR2_X1 U10104 ( .A(n8686), .B(n8685), .ZN(n8691) );
  AOI22_X1 U10105 ( .A1(n9229), .A2(n8801), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8688) );
  NAND2_X1 U10106 ( .A1(n9223), .A2(n8802), .ZN(n8687) );
  OAI211_X1 U10107 ( .C1(n9196), .C2(n8805), .A(n8688), .B(n8687), .ZN(n8689)
         );
  AOI21_X1 U10108 ( .B1(n9390), .B2(n8807), .A(n8689), .ZN(n8690) );
  OAI21_X1 U10109 ( .B1(n8691), .B2(n8782), .A(n8690), .ZN(P1_U3214) );
  INV_X1 U10110 ( .A(n8695), .ZN(n8692) );
  NOR2_X1 U10111 ( .A1(n8693), .A2(n8692), .ZN(n8698) );
  AOI21_X1 U10112 ( .B1(n8696), .B2(n8695), .A(n8694), .ZN(n8697) );
  OAI21_X1 U10113 ( .B1(n8698), .B2(n8697), .A(n8765), .ZN(n8703) );
  NOR2_X1 U10114 ( .A1(n8699), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9138) );
  AOI21_X1 U10115 ( .B1(n8801), .B2(n10326), .A(n9138), .ZN(n8700) );
  OAI21_X1 U10116 ( .B1(n8805), .B2(n9251), .A(n8700), .ZN(n8701) );
  AOI21_X1 U10117 ( .B1(n9281), .B2(n8802), .A(n8701), .ZN(n8702) );
  OAI211_X1 U10118 ( .C1(n9283), .C2(n8750), .A(n8703), .B(n8702), .ZN(
        P1_U3217) );
  XOR2_X1 U10119 ( .A(n8705), .B(n8704), .Z(n8710) );
  AOI22_X1 U10120 ( .A1(n9229), .A2(n8789), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8707) );
  NAND2_X1 U10121 ( .A1(n8802), .A2(n9255), .ZN(n8706) );
  OAI211_X1 U10122 ( .C1(n9251), .C2(n8778), .A(n8707), .B(n8706), .ZN(n8708)
         );
  AOI21_X1 U10123 ( .B1(n9402), .B2(n8807), .A(n8708), .ZN(n8709) );
  OAI21_X1 U10124 ( .B1(n8710), .B2(n8782), .A(n8709), .ZN(P1_U3221) );
  XOR2_X1 U10125 ( .A(n8711), .B(n4535), .Z(n8716) );
  AOI22_X1 U10126 ( .A1(n9230), .A2(n8801), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8713) );
  NAND2_X1 U10127 ( .A1(n9197), .A2(n8802), .ZN(n8712) );
  OAI211_X1 U10128 ( .C1(n9195), .C2(n8805), .A(n8713), .B(n8712), .ZN(n8714)
         );
  AOI21_X1 U10129 ( .B1(n9382), .B2(n8807), .A(n8714), .ZN(n8715) );
  OAI21_X1 U10130 ( .B1(n8716), .B2(n8782), .A(n8715), .ZN(P1_U3223) );
  XNOR2_X1 U10131 ( .A(n8718), .B(n8717), .ZN(n8719) );
  XNOR2_X1 U10132 ( .A(n8720), .B(n8719), .ZN(n8726) );
  NOR2_X1 U10133 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8721), .ZN(n9675) );
  AOI21_X1 U10134 ( .B1(n8801), .B2(n9086), .A(n9675), .ZN(n8723) );
  NAND2_X1 U10135 ( .A1(n8802), .A2(n9333), .ZN(n8722) );
  OAI211_X1 U10136 ( .C1(n8805), .C2(n9331), .A(n8723), .B(n8722), .ZN(n8724)
         );
  AOI21_X1 U10137 ( .B1(n9427), .B2(n8807), .A(n8724), .ZN(n8725) );
  OAI21_X1 U10138 ( .B1(n8726), .B2(n8782), .A(n8725), .ZN(P1_U3224) );
  XOR2_X1 U10139 ( .A(n8728), .B(n8727), .Z(n8733) );
  NOR2_X1 U10140 ( .A1(n8792), .A2(n9310), .ZN(n8731) );
  NAND2_X1 U10141 ( .A1(n8789), .A2(n10326), .ZN(n8729) );
  NAND2_X1 U10142 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9688) );
  OAI211_X1 U10143 ( .C1(n9343), .C2(n8778), .A(n8729), .B(n9688), .ZN(n8730)
         );
  AOI211_X1 U10144 ( .C1(n9420), .C2(n8807), .A(n8731), .B(n8730), .ZN(n8732)
         );
  OAI21_X1 U10145 ( .B1(n8733), .B2(n8782), .A(n8732), .ZN(P1_U3226) );
  XOR2_X1 U10146 ( .A(n8735), .B(n8734), .Z(n8740) );
  NAND2_X1 U10147 ( .A1(n9185), .A2(n8789), .ZN(n8737) );
  AOI22_X1 U10148 ( .A1(n9242), .A2(n8801), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8736) );
  OAI211_X1 U10149 ( .C1(n8792), .C2(n9212), .A(n8737), .B(n8736), .ZN(n8738)
         );
  AOI21_X1 U10150 ( .B1(n9387), .B2(n8807), .A(n8738), .ZN(n8739) );
  OAI21_X1 U10151 ( .B1(n8740), .B2(n8782), .A(n8739), .ZN(P1_U3227) );
  OAI21_X1 U10152 ( .B1(n8743), .B2(n8742), .A(n8741), .ZN(n8744) );
  NAND2_X1 U10153 ( .A1(n8744), .A2(n8765), .ZN(n8749) );
  INV_X1 U10154 ( .A(n8745), .ZN(n9267) );
  AOI22_X1 U10155 ( .A1(n8801), .A2(n9274), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8746) );
  OAI21_X1 U10156 ( .B1(n8758), .B2(n8805), .A(n8746), .ZN(n8747) );
  AOI21_X1 U10157 ( .B1(n9267), .B2(n8802), .A(n8747), .ZN(n8748) );
  OAI211_X1 U10158 ( .C1(n9269), .C2(n8750), .A(n8749), .B(n8748), .ZN(
        P1_U3231) );
  INV_X1 U10159 ( .A(n8751), .ZN(n8752) );
  NOR2_X1 U10160 ( .A1(n8753), .A2(n8752), .ZN(n8755) );
  XNOR2_X1 U10161 ( .A(n8755), .B(n8754), .ZN(n8761) );
  AOI22_X1 U10162 ( .A1(n9242), .A2(n8789), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8757) );
  NAND2_X1 U10163 ( .A1(n8802), .A2(n9238), .ZN(n8756) );
  OAI211_X1 U10164 ( .C1(n8758), .C2(n8778), .A(n8757), .B(n8756), .ZN(n8759)
         );
  AOI21_X1 U10165 ( .B1(n9395), .B2(n8807), .A(n8759), .ZN(n8760) );
  OAI21_X1 U10166 ( .B1(n8761), .B2(n8782), .A(n8760), .ZN(P1_U3233) );
  OAI21_X1 U10167 ( .B1(n8764), .B2(n8763), .A(n8762), .ZN(n8766) );
  NAND2_X1 U10168 ( .A1(n8766), .A2(n8765), .ZN(n8771) );
  AOI22_X1 U10169 ( .A1(n8801), .A2(n9101), .B1(n8789), .B2(n9098), .ZN(n8770)
         );
  AOI22_X1 U10170 ( .A1(P1_REG3_REG_2__SCAN_IN), .A2(n8768), .B1(n8807), .B2(
        n8767), .ZN(n8769) );
  NAND3_X1 U10171 ( .A1(n8771), .A2(n8770), .A3(n8769), .ZN(P1_U3235) );
  INV_X1 U10172 ( .A(n8772), .ZN(n8773) );
  NOR2_X1 U10173 ( .A1(n8774), .A2(n8773), .ZN(n8776) );
  XNOR2_X1 U10174 ( .A(n8776), .B(n8775), .ZN(n8783) );
  NOR2_X1 U10175 ( .A1(n8792), .A2(n9295), .ZN(n8780) );
  NAND2_X1 U10176 ( .A1(n8789), .A2(n9274), .ZN(n8777) );
  NAND2_X1 U10177 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9700) );
  OAI211_X1 U10178 ( .C1(n9331), .C2(n8778), .A(n8777), .B(n9700), .ZN(n8779)
         );
  AOI211_X1 U10179 ( .C1(n9417), .C2(n8807), .A(n8780), .B(n8779), .ZN(n8781)
         );
  OAI21_X1 U10180 ( .B1(n8783), .B2(n8782), .A(n8781), .ZN(P1_U3236) );
  INV_X1 U10181 ( .A(n8784), .ZN(n8786) );
  NAND2_X1 U10182 ( .A1(n8786), .A2(n8785), .ZN(n8787) );
  XNOR2_X1 U10183 ( .A(n8788), .B(n8787), .ZN(n8795) );
  NAND2_X1 U10184 ( .A1(n9186), .A2(n8789), .ZN(n8791) );
  AOI22_X1 U10185 ( .A1(n9185), .A2(n8801), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n8790) );
  OAI211_X1 U10186 ( .C1(n8792), .C2(n9177), .A(n8791), .B(n8790), .ZN(n8793)
         );
  AOI21_X1 U10187 ( .B1(n9375), .B2(n8807), .A(n8793), .ZN(n8794) );
  OAI21_X1 U10188 ( .B1(n8795), .B2(n8782), .A(n8794), .ZN(P1_U3238) );
  INV_X1 U10189 ( .A(n8796), .ZN(n8798) );
  NAND2_X1 U10190 ( .A1(n8798), .A2(n8797), .ZN(n8800) );
  XNOR2_X1 U10191 ( .A(n8800), .B(n8799), .ZN(n8809) );
  AND2_X1 U10192 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9666) );
  AOI21_X1 U10193 ( .B1(n8801), .B2(n9087), .A(n9666), .ZN(n8804) );
  NAND2_X1 U10194 ( .A1(n8802), .A2(n9355), .ZN(n8803) );
  OAI211_X1 U10195 ( .C1(n8805), .C2(n9343), .A(n8804), .B(n8803), .ZN(n8806)
         );
  AOI21_X1 U10196 ( .B1(n9430), .B2(n8807), .A(n8806), .ZN(n8808) );
  OAI21_X1 U10197 ( .B1(n8809), .B2(n8782), .A(n8808), .ZN(P1_U3239) );
  INV_X1 U10198 ( .A(n9083), .ZN(n8914) );
  NAND2_X1 U10199 ( .A1(n9144), .A2(n8914), .ZN(n8921) );
  AND2_X1 U10200 ( .A1(n8917), .A2(n9020), .ZN(n8819) );
  AND2_X1 U10201 ( .A1(n8810), .A2(n8922), .ZN(n9022) );
  INV_X1 U10202 ( .A(n9022), .ZN(n8815) );
  NAND2_X1 U10203 ( .A1(n8925), .A2(n9001), .ZN(n8811) );
  OR2_X1 U10204 ( .A1(n9387), .A2(n9196), .ZN(n9006) );
  NAND2_X1 U10205 ( .A1(n8811), .A2(n9006), .ZN(n8812) );
  NAND2_X1 U10206 ( .A1(n9012), .A2(n8812), .ZN(n8928) );
  NAND2_X1 U10207 ( .A1(n9017), .A2(n8928), .ZN(n8813) );
  INV_X1 U10208 ( .A(n9018), .ZN(n8821) );
  AOI21_X1 U10209 ( .B1(n9014), .B2(n8813), .A(n8821), .ZN(n8814) );
  OR2_X1 U10210 ( .A1(n8815), .A2(n8814), .ZN(n8817) );
  INV_X1 U10211 ( .A(n8918), .ZN(n8816) );
  AOI21_X1 U10212 ( .B1(n8819), .B2(n8817), .A(n8816), .ZN(n8818) );
  NAND2_X1 U10213 ( .A1(n8921), .A2(n8818), .ZN(n9064) );
  NAND2_X1 U10214 ( .A1(n9144), .A2(n8913), .ZN(n8920) );
  INV_X1 U10215 ( .A(n8819), .ZN(n8822) );
  INV_X1 U10216 ( .A(n9017), .ZN(n8820) );
  OR3_X1 U10217 ( .A1(n8822), .A2(n8821), .A3(n8820), .ZN(n9062) );
  INV_X1 U10218 ( .A(n9062), .ZN(n8872) );
  NAND2_X1 U10219 ( .A1(n9006), .A2(n8926), .ZN(n9009) );
  INV_X1 U10220 ( .A(n9009), .ZN(n8834) );
  NAND2_X1 U10221 ( .A1(n8831), .A2(n8828), .ZN(n8929) );
  INV_X1 U10222 ( .A(n8989), .ZN(n8823) );
  OR2_X1 U10223 ( .A1(n8929), .A2(n8823), .ZN(n9003) );
  AND2_X1 U10224 ( .A1(n9270), .A2(n8824), .ZN(n8996) );
  INV_X1 U10225 ( .A(n8996), .ZN(n8825) );
  NOR2_X1 U10226 ( .A1(n8825), .A2(n8931), .ZN(n8826) );
  OR2_X1 U10227 ( .A1(n8998), .A2(n8826), .ZN(n8832) );
  INV_X1 U10228 ( .A(n8827), .ZN(n8878) );
  NAND2_X1 U10229 ( .A1(n8828), .A2(n8878), .ZN(n8829) );
  AND2_X1 U10230 ( .A1(n8829), .A2(n8992), .ZN(n8830) );
  NAND2_X1 U10231 ( .A1(n8830), .A2(n8993), .ZN(n8867) );
  NAND2_X1 U10232 ( .A1(n8867), .A2(n8831), .ZN(n9000) );
  OAI21_X1 U10233 ( .B1(n9003), .B2(n8832), .A(n9000), .ZN(n8833) );
  NAND2_X1 U10234 ( .A1(n8834), .A2(n8833), .ZN(n8869) );
  NAND2_X1 U10235 ( .A1(n8835), .A2(n9344), .ZN(n8972) );
  NAND2_X1 U10236 ( .A1(n8972), .A2(n8836), .ZN(n8967) );
  INV_X1 U10237 ( .A(n8967), .ZN(n8840) );
  INV_X1 U10238 ( .A(n9498), .ZN(n8837) );
  OAI211_X1 U10239 ( .C1(n8837), .C2(n8949), .A(n8963), .B(n8962), .ZN(n8838)
         );
  INV_X1 U10240 ( .A(n8838), .ZN(n8839) );
  NAND3_X1 U10241 ( .A1(n8979), .A2(n8840), .A3(n8839), .ZN(n8861) );
  AND2_X1 U10242 ( .A1(n9498), .A2(n8948), .ZN(n8841) );
  OR2_X1 U10243 ( .A1(n8861), .A2(n8841), .ZN(n8849) );
  NAND2_X1 U10244 ( .A1(n8846), .A2(n8842), .ZN(n8973) );
  NAND2_X1 U10245 ( .A1(n8964), .A2(n8843), .ZN(n8844) );
  AND2_X1 U10246 ( .A1(n8844), .A2(n8963), .ZN(n8845) );
  NOR2_X1 U10247 ( .A1(n8973), .A2(n8845), .ZN(n8968) );
  INV_X1 U10248 ( .A(n8968), .ZN(n8847) );
  NAND2_X1 U10249 ( .A1(n8967), .A2(n8846), .ZN(n8974) );
  NAND3_X1 U10250 ( .A1(n8847), .A2(n8974), .A3(n8979), .ZN(n8848) );
  NAND4_X1 U10251 ( .A1(n8849), .A2(n8983), .A3(n8978), .A4(n8848), .ZN(n8850)
         );
  NAND2_X1 U10252 ( .A1(n8850), .A2(n8982), .ZN(n8851) );
  OR2_X1 U10253 ( .A1(n8930), .A2(n8851), .ZN(n8863) );
  NAND2_X1 U10254 ( .A1(n8863), .A2(n8944), .ZN(n8852) );
  OR2_X1 U10255 ( .A1(n8869), .A2(n8852), .ZN(n9059) );
  AND2_X1 U10256 ( .A1(n8854), .A2(n8853), .ZN(n9050) );
  AND2_X1 U10257 ( .A1(n9055), .A2(n9050), .ZN(n8859) );
  NAND2_X1 U10258 ( .A1(n9048), .A2(n9052), .ZN(n8855) );
  NAND3_X1 U10259 ( .A1(n8855), .A2(n8938), .A3(n8854), .ZN(n8857) );
  INV_X1 U10260 ( .A(n8933), .ZN(n8856) );
  AOI21_X1 U10261 ( .B1(n9053), .B2(n8857), .A(n8856), .ZN(n8858) );
  AOI21_X1 U10262 ( .B1(n8860), .B2(n8859), .A(n8858), .ZN(n8870) );
  INV_X1 U10263 ( .A(n8861), .ZN(n8862) );
  NAND3_X1 U10264 ( .A1(n8862), .A2(n8982), .A3(n8934), .ZN(n8864) );
  OAI21_X1 U10265 ( .B1(n8930), .B2(n8864), .A(n8863), .ZN(n8865) );
  NAND2_X1 U10266 ( .A1(n8865), .A2(n9270), .ZN(n8866) );
  NOR2_X1 U10267 ( .A1(n8867), .A2(n8866), .ZN(n8868) );
  OR2_X1 U10268 ( .A1(n8869), .A2(n8868), .ZN(n9057) );
  OAI21_X1 U10269 ( .B1(n9059), .B2(n8870), .A(n9057), .ZN(n8871) );
  NAND2_X1 U10270 ( .A1(n8872), .A2(n8871), .ZN(n8873) );
  NAND2_X1 U10271 ( .A1(n8920), .A2(n8873), .ZN(n8875) );
  NAND2_X1 U10272 ( .A1(n8876), .A2(n8913), .ZN(n8916) );
  OR2_X1 U10273 ( .A1(n9144), .A2(n8914), .ZN(n8874) );
  NAND2_X1 U10274 ( .A1(n8916), .A2(n8874), .ZN(n9066) );
  NAND2_X1 U10275 ( .A1(n9066), .A2(n8876), .ZN(n9029) );
  OAI21_X1 U10276 ( .B1(n9064), .B2(n8875), .A(n9029), .ZN(n8877) );
  OR2_X1 U10277 ( .A1(n8876), .A2(n8913), .ZN(n9067) );
  NAND3_X1 U10278 ( .A1(n8877), .A2(n5671), .A3(n9067), .ZN(n8912) );
  INV_X1 U10279 ( .A(n9067), .ZN(n8910) );
  INV_X1 U10280 ( .A(n9028), .ZN(n8908) );
  INV_X1 U10281 ( .A(n9262), .ZN(n9271) );
  INV_X1 U10282 ( .A(n9345), .ZN(n9341) );
  INV_X1 U10283 ( .A(n8879), .ZN(n8881) );
  NAND4_X1 U10284 ( .A1(n8883), .A2(n8882), .A3(n8881), .A4(n8880), .ZN(n8886)
         );
  NOR3_X1 U10285 ( .A1(n8886), .A2(n8885), .A3(n8884), .ZN(n8889) );
  NAND4_X1 U10286 ( .A1(n8889), .A2(n8939), .A3(n8888), .A4(n4924), .ZN(n8891)
         );
  OR3_X1 U10287 ( .A1(n9492), .A2(n8891), .A3(n8890), .ZN(n8892) );
  NOR2_X1 U10288 ( .A1(n8893), .A2(n8892), .ZN(n8894) );
  NAND3_X1 U10289 ( .A1(n8895), .A2(n8894), .A3(n4588), .ZN(n8896) );
  NOR2_X1 U10290 ( .A1(n9341), .A2(n8896), .ZN(n8898) );
  NAND4_X1 U10291 ( .A1(n9315), .A2(n9327), .A3(n8898), .A4(n8897), .ZN(n8899)
         );
  NOR3_X1 U10292 ( .A1(n9284), .A2(n9302), .A3(n8899), .ZN(n8900) );
  NAND4_X1 U10293 ( .A1(n4567), .A2(n8901), .A3(n9271), .A4(n8900), .ZN(n8903)
         );
  INV_X1 U10294 ( .A(n9241), .ZN(n8902) );
  INV_X1 U10295 ( .A(n9206), .ZN(n9203) );
  INV_X1 U10296 ( .A(n8904), .ZN(n8906) );
  AND4_X1 U10297 ( .A1(n9024), .A2(n5044), .A3(n9203), .A4(n9184), .ZN(n8907)
         );
  NAND4_X1 U10298 ( .A1(n8921), .A2(n9022), .A3(n8908), .A4(n8907), .ZN(n8909)
         );
  AND2_X1 U10299 ( .A1(n8912), .A2(n9035), .ZN(n9038) );
  OAI211_X1 U10300 ( .C1(n8914), .C2(n8913), .A(n9144), .B(n9004), .ZN(n8915)
         );
  AND2_X1 U10301 ( .A1(n9067), .A2(n8915), .ZN(n9034) );
  INV_X1 U10302 ( .A(n8916), .ZN(n9033) );
  MUX2_X1 U10303 ( .A(n8918), .B(n8917), .S(n9004), .Z(n8919) );
  INV_X1 U10304 ( .A(n9004), .ZN(n9030) );
  NAND3_X1 U10305 ( .A1(n8922), .A2(n9030), .A3(n9014), .ZN(n9016) );
  NAND2_X1 U10306 ( .A1(n8923), .A2(n9004), .ZN(n8924) );
  INV_X1 U10307 ( .A(n8925), .ZN(n9008) );
  OAI21_X1 U10308 ( .B1(n9008), .B2(n8926), .A(n9181), .ZN(n8927) );
  MUX2_X1 U10309 ( .A(n8928), .B(n8927), .S(n9004), .Z(n9015) );
  INV_X1 U10310 ( .A(n8929), .ZN(n8995) );
  INV_X1 U10311 ( .A(n8930), .ZN(n8932) );
  MUX2_X1 U10312 ( .A(n8932), .B(n8931), .S(n9004), .Z(n8987) );
  NAND2_X1 U10313 ( .A1(n8935), .A2(n8934), .ZN(n8947) );
  NAND2_X1 U10314 ( .A1(n8937), .A2(n8936), .ZN(n8940) );
  NAND3_X1 U10315 ( .A1(n8940), .A2(n8939), .A3(n8938), .ZN(n8943) );
  NAND3_X1 U10316 ( .A1(n8943), .A2(n8942), .A3(n8941), .ZN(n8945) );
  NAND2_X1 U10317 ( .A1(n8945), .A2(n8944), .ZN(n8946) );
  MUX2_X1 U10318 ( .A(n8947), .B(n8946), .S(n9004), .Z(n8956) );
  INV_X1 U10319 ( .A(n8956), .ZN(n8950) );
  INV_X1 U10320 ( .A(n8948), .ZN(n8954) );
  NAND2_X1 U10321 ( .A1(n8963), .A2(n8951), .ZN(n8952) );
  AOI21_X1 U10322 ( .B1(n8956), .B2(n8955), .A(n8954), .ZN(n8958) );
  INV_X1 U10323 ( .A(n9494), .ZN(n8957) );
  OAI21_X1 U10324 ( .B1(n8958), .B2(n8957), .A(n9498), .ZN(n8959) );
  MUX2_X1 U10325 ( .A(n8959), .B(n9498), .S(n9030), .Z(n8960) );
  NAND2_X1 U10326 ( .A1(n8961), .A2(n8960), .ZN(n8971) );
  NAND2_X1 U10327 ( .A1(n8963), .A2(n8962), .ZN(n8965) );
  AND2_X1 U10328 ( .A1(n8965), .A2(n8964), .ZN(n8966) );
  NOR2_X1 U10329 ( .A1(n8967), .A2(n8966), .ZN(n8969) );
  MUX2_X1 U10330 ( .A(n8969), .B(n8968), .S(n9004), .Z(n8970) );
  NAND2_X1 U10331 ( .A1(n8971), .A2(n8970), .ZN(n8977) );
  NAND2_X1 U10332 ( .A1(n8973), .A2(n8972), .ZN(n8975) );
  MUX2_X1 U10333 ( .A(n8975), .B(n8974), .S(n9004), .Z(n8976) );
  NAND3_X1 U10334 ( .A1(n8977), .A2(n9345), .A3(n8976), .ZN(n8981) );
  MUX2_X1 U10335 ( .A(n8979), .B(n8978), .S(n9004), .Z(n8980) );
  NAND3_X1 U10336 ( .A1(n8981), .A2(n9327), .A3(n8980), .ZN(n8985) );
  MUX2_X1 U10337 ( .A(n8983), .B(n8982), .S(n9004), .Z(n8984) );
  NAND3_X1 U10338 ( .A1(n8985), .A2(n9315), .A3(n8984), .ZN(n8986) );
  NAND2_X1 U10339 ( .A1(n8987), .A2(n8986), .ZN(n8997) );
  NAND3_X1 U10340 ( .A1(n8997), .A2(n8989), .A3(n8988), .ZN(n8991) );
  INV_X1 U10341 ( .A(n8993), .ZN(n8994) );
  NAND2_X1 U10342 ( .A1(n8997), .A2(n8996), .ZN(n8999) );
  NAND2_X1 U10343 ( .A1(n8999), .A2(n4716), .ZN(n9002) );
  OAI211_X1 U10344 ( .C1(n9003), .C2(n9002), .A(n9001), .B(n9000), .ZN(n9005)
         );
  NAND2_X1 U10345 ( .A1(n9007), .A2(n9006), .ZN(n9011) );
  AOI21_X1 U10346 ( .B1(n9030), .B2(n9009), .A(n9008), .ZN(n9010) );
  OR2_X1 U10347 ( .A1(n9012), .A2(n9030), .ZN(n9013) );
  NAND2_X1 U10348 ( .A1(n9019), .A2(n9018), .ZN(n9025) );
  INV_X1 U10349 ( .A(n9020), .ZN(n9021) );
  AOI21_X1 U10350 ( .B1(n9025), .B2(n9022), .A(n9021), .ZN(n9027) );
  AOI21_X1 U10351 ( .B1(n9025), .B2(n9024), .A(n9023), .ZN(n9026) );
  NAND3_X1 U10352 ( .A1(n9066), .A2(n9030), .A3(n8876), .ZN(n9031) );
  OAI211_X1 U10353 ( .C1(n9034), .C2(n9033), .A(n9032), .B(n9031), .ZN(n9039)
         );
  OAI21_X1 U10354 ( .B1(n9039), .B2(n9036), .A(n9035), .ZN(n9037) );
  MUX2_X1 U10355 ( .A(n9038), .B(n9037), .S(n9257), .Z(n9070) );
  INV_X1 U10356 ( .A(n9040), .ZN(n9041) );
  OAI211_X1 U10357 ( .C1(n5644), .C2(n9042), .A(n9041), .B(n5671), .ZN(n9043)
         );
  INV_X1 U10358 ( .A(n9043), .ZN(n9045) );
  OAI21_X1 U10359 ( .B1(n9046), .B2(n9045), .A(n9044), .ZN(n9049) );
  NAND3_X1 U10360 ( .A1(n9049), .A2(n9048), .A3(n9047), .ZN(n9051) );
  NAND2_X1 U10361 ( .A1(n9051), .A2(n9050), .ZN(n9054) );
  NAND3_X1 U10362 ( .A1(n9054), .A2(n9053), .A3(n9052), .ZN(n9056) );
  NAND2_X1 U10363 ( .A1(n9056), .A2(n9055), .ZN(n9058) );
  OAI21_X1 U10364 ( .B1(n9059), .B2(n9058), .A(n9057), .ZN(n9060) );
  INV_X1 U10365 ( .A(n9060), .ZN(n9061) );
  NOR2_X1 U10366 ( .A1(n9062), .A2(n9061), .ZN(n9063) );
  NOR2_X1 U10367 ( .A1(n9064), .A2(n9063), .ZN(n9065) );
  OR2_X1 U10368 ( .A1(n9066), .A2(n9065), .ZN(n9068) );
  NAND2_X1 U10369 ( .A1(n9068), .A2(n9067), .ZN(n9073) );
  OAI21_X1 U10370 ( .B1(n9073), .B2(n9072), .A(n9071), .ZN(n9080) );
  NOR2_X1 U10371 ( .A1(n5635), .A2(n9074), .ZN(n9592) );
  NAND3_X1 U10372 ( .A1(n9075), .A2(n9722), .A3(n9592), .ZN(n9076) );
  OAI211_X1 U10373 ( .C1(n9078), .C2(n9077), .A(n9076), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9079) );
  OAI21_X1 U10374 ( .B1(n9081), .B2(n9080), .A(n9079), .ZN(P1_U3240) );
  MUX2_X1 U10375 ( .A(n9082), .B(P1_DATAO_REG_31__SCAN_IN), .S(n9100), .Z(
        P1_U3586) );
  MUX2_X1 U10376 ( .A(n9083), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9100), .Z(
        P1_U3585) );
  MUX2_X1 U10377 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9084), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10378 ( .A(n9171), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9100), .Z(
        P1_U3583) );
  MUX2_X1 U10379 ( .A(n9186), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9100), .Z(
        P1_U3582) );
  MUX2_X1 U10380 ( .A(n9164), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9100), .Z(
        P1_U3581) );
  MUX2_X1 U10381 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9185), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10382 ( .A(n9230), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9100), .Z(
        P1_U3579) );
  MUX2_X1 U10383 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9242), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10384 ( .A(n9229), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9100), .Z(
        P1_U3577) );
  MUX2_X1 U10385 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9273), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10386 ( .A(n9286), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9100), .Z(
        P1_U3575) );
  MUX2_X1 U10387 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9274), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10388 ( .A(n9085), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9100), .Z(
        P1_U3572) );
  MUX2_X1 U10389 ( .A(n9318), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9100), .Z(
        P1_U3571) );
  MUX2_X1 U10390 ( .A(n9086), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9100), .Z(
        P1_U3570) );
  MUX2_X1 U10391 ( .A(n9087), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9100), .Z(
        P1_U3569) );
  MUX2_X1 U10392 ( .A(n9088), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9100), .Z(
        P1_U3568) );
  MUX2_X1 U10393 ( .A(n9089), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9100), .Z(
        P1_U3567) );
  MUX2_X1 U10394 ( .A(n9090), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9100), .Z(
        P1_U3566) );
  MUX2_X1 U10395 ( .A(n9091), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9100), .Z(
        P1_U3565) );
  MUX2_X1 U10396 ( .A(n9092), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9100), .Z(
        P1_U3564) );
  MUX2_X1 U10397 ( .A(n9093), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9100), .Z(
        P1_U3563) );
  MUX2_X1 U10398 ( .A(n9094), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9100), .Z(
        P1_U3562) );
  MUX2_X1 U10399 ( .A(n9095), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9100), .Z(
        P1_U3561) );
  MUX2_X1 U10400 ( .A(n9096), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9100), .Z(
        P1_U3560) );
  MUX2_X1 U10401 ( .A(n9097), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9100), .Z(
        P1_U3559) );
  MUX2_X1 U10402 ( .A(n9098), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9100), .Z(
        P1_U3558) );
  MUX2_X1 U10403 ( .A(n9099), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9100), .Z(
        P1_U3557) );
  MUX2_X1 U10404 ( .A(n9101), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9100), .Z(
        P1_U3556) );
  MUX2_X1 U10405 ( .A(n9102), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9100), .Z(
        P1_U3555) );
  INV_X1 U10406 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9141) );
  OR2_X1 U10407 ( .A1(n9103), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9105) );
  XNOR2_X1 U10408 ( .A(n9119), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n9620) );
  NAND2_X1 U10409 ( .A1(n9619), .A2(n9620), .ZN(n9618) );
  INV_X1 U10410 ( .A(n9119), .ZN(n9624) );
  NAND2_X1 U10411 ( .A1(n9624), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n9106) );
  MUX2_X1 U10412 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n9107), .S(n9638), .Z(n9633) );
  NOR2_X1 U10413 ( .A1(n9108), .A2(n9653), .ZN(n9109) );
  INV_X1 U10414 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9647) );
  NOR2_X1 U10415 ( .A1(n9647), .A2(n9648), .ZN(n9646) );
  NOR2_X1 U10416 ( .A1(n9109), .A2(n9646), .ZN(n9110) );
  NOR2_X1 U10417 ( .A1(n9110), .A2(n9122), .ZN(n9111) );
  INV_X1 U10418 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9663) );
  NAND2_X1 U10419 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9676), .ZN(n9112) );
  OAI21_X1 U10420 ( .B1(n9676), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9112), .ZN(
        n9673) );
  AOI21_X1 U10421 ( .B1(n9676), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9672), .ZN(
        n9684) );
  NAND2_X1 U10422 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9116), .ZN(n9113) );
  OAI21_X1 U10423 ( .B1(n9116), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9113), .ZN(
        n9685) );
  NOR2_X1 U10424 ( .A1(n9684), .A2(n9685), .ZN(n9683) );
  INV_X1 U10425 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9114) );
  MUX2_X1 U10426 ( .A(P1_REG2_REG_18__SCAN_IN), .B(n9114), .S(n9708), .Z(n9115) );
  INV_X1 U10427 ( .A(n9115), .ZN(n9703) );
  INV_X1 U10428 ( .A(n9134), .ZN(n9132) );
  INV_X1 U10429 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9128) );
  XNOR2_X1 U10430 ( .A(n9708), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9711) );
  INV_X1 U10431 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9126) );
  XNOR2_X1 U10432 ( .A(n9690), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9696) );
  INV_X1 U10433 ( .A(n9676), .ZN(n9125) );
  INV_X1 U10434 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9124) );
  XOR2_X1 U10435 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9676), .Z(n9678) );
  INV_X1 U10436 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9540) );
  INV_X1 U10437 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9547) );
  INV_X1 U10438 ( .A(n9638), .ZN(n9120) );
  INV_X1 U10439 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9554) );
  AOI21_X1 U10440 ( .B1(n9118), .B2(n6503), .A(n9117), .ZN(n9627) );
  MUX2_X1 U10441 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9554), .S(n9119), .Z(n9626) );
  NOR2_X1 U10442 ( .A1(n9627), .A2(n9626), .ZN(n9625) );
  AOI21_X1 U10443 ( .B1(n9554), .B2(n9119), .A(n9625), .ZN(n9641) );
  MUX2_X1 U10444 ( .A(n9547), .B(P1_REG1_REG_13__SCAN_IN), .S(n9638), .Z(n9640) );
  NOR2_X1 U10445 ( .A1(n9641), .A2(n9640), .ZN(n9639) );
  AOI21_X1 U10446 ( .B1(n9547), .B2(n9120), .A(n9639), .ZN(n9657) );
  MUX2_X1 U10447 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9540), .S(n9653), .Z(n9656) );
  NOR2_X1 U10448 ( .A1(n9657), .A2(n9656), .ZN(n9655) );
  AOI21_X1 U10449 ( .B1(n9653), .B2(n9540), .A(n9655), .ZN(n9121) );
  NAND2_X1 U10450 ( .A1(n9667), .A2(n9121), .ZN(n9123) );
  XNOR2_X1 U10451 ( .A(n9122), .B(n9121), .ZN(n9669) );
  NAND2_X1 U10452 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9669), .ZN(n9668) );
  NAND2_X1 U10453 ( .A1(n9123), .A2(n9668), .ZN(n9679) );
  NAND2_X1 U10454 ( .A1(n9678), .A2(n9679), .ZN(n9677) );
  OAI21_X1 U10455 ( .B1(n9125), .B2(n9124), .A(n9677), .ZN(n9695) );
  NAND2_X1 U10456 ( .A1(n9696), .A2(n9695), .ZN(n9694) );
  OAI21_X1 U10457 ( .B1(n9690), .B2(n9126), .A(n9694), .ZN(n9710) );
  NOR2_X1 U10458 ( .A1(n9711), .A2(n9710), .ZN(n9709) );
  AOI21_X1 U10459 ( .B1(n9128), .B2(n9127), .A(n9709), .ZN(n9129) );
  XOR2_X1 U10460 ( .A(n9129), .B(P1_REG1_REG_19__SCAN_IN), .Z(n9133) );
  OAI21_X1 U10461 ( .B1(n9133), .B2(n9712), .A(n9691), .ZN(n9130) );
  AOI21_X1 U10462 ( .B1(n9132), .B2(n9131), .A(n9130), .ZN(n9137) );
  AOI22_X1 U10463 ( .A1(n9134), .A2(n9687), .B1(n9693), .B2(n9133), .ZN(n9136)
         );
  MUX2_X1 U10464 ( .A(n9137), .B(n9136), .S(n9135), .Z(n9140) );
  INV_X1 U10465 ( .A(n9138), .ZN(n9139) );
  OAI211_X1 U10466 ( .C1(n9141), .C2(n9716), .A(n9140), .B(n9139), .ZN(
        P1_U3260) );
  INV_X1 U10467 ( .A(n9144), .ZN(n9530) );
  AOI21_X1 U10468 ( .B1(n9144), .B2(n9143), .A(n9142), .ZN(n9532) );
  NAND2_X1 U10469 ( .A1(n9532), .A2(n9361), .ZN(n9147) );
  AOI21_X1 U10470 ( .B1(n9519), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9145), .ZN(
        n9146) );
  OAI211_X1 U10471 ( .C1(n9530), .C2(n9357), .A(n9147), .B(n9146), .ZN(
        P1_U3262) );
  NAND2_X1 U10472 ( .A1(n9148), .A2(n9515), .ZN(n9151) );
  AOI22_X1 U10473 ( .A1(n9149), .A2(n9508), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9312), .ZN(n9150) );
  OAI211_X1 U10474 ( .C1(n9152), .C2(n9357), .A(n9151), .B(n9150), .ZN(n9153)
         );
  AOI21_X1 U10475 ( .B1(n9154), .B2(n9338), .A(n9153), .ZN(n9155) );
  OAI21_X1 U10476 ( .B1(n9156), .B2(n9340), .A(n9155), .ZN(P1_U3263) );
  XOR2_X1 U10477 ( .A(n9168), .B(n9157), .Z(n9374) );
  INV_X1 U10478 ( .A(n9176), .ZN(n9160) );
  INV_X1 U10479 ( .A(n9158), .ZN(n9159) );
  AOI21_X1 U10480 ( .B1(n9370), .B2(n9160), .A(n9159), .ZN(n9371) );
  AOI22_X1 U10481 ( .A1(n9161), .A2(n9508), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9312), .ZN(n9162) );
  OAI21_X1 U10482 ( .B1(n9163), .B2(n9357), .A(n9162), .ZN(n9173) );
  AND2_X1 U10483 ( .A1(n9164), .A2(n9317), .ZN(n9170) );
  INV_X1 U10484 ( .A(n9165), .ZN(n9166) );
  AOI211_X1 U10485 ( .C1(n9168), .C2(n9167), .A(n9497), .B(n9166), .ZN(n9169)
         );
  NOR2_X1 U10486 ( .A1(n9373), .A2(n9519), .ZN(n9172) );
  AOI211_X1 U10487 ( .C1(n9361), .C2(n9371), .A(n9173), .B(n9172), .ZN(n9174)
         );
  OAI21_X1 U10488 ( .B1(n9374), .B2(n9340), .A(n9174), .ZN(P1_U3264) );
  XOR2_X1 U10489 ( .A(n9184), .B(n9175), .Z(n9379) );
  AOI21_X1 U10490 ( .B1(n9375), .B2(n5045), .A(n9176), .ZN(n9376) );
  INV_X1 U10491 ( .A(n9375), .ZN(n9180) );
  INV_X1 U10492 ( .A(n9177), .ZN(n9178) );
  AOI22_X1 U10493 ( .A1(n9178), .A2(n9508), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9312), .ZN(n9179) );
  OAI21_X1 U10494 ( .B1(n9180), .B2(n9357), .A(n9179), .ZN(n9189) );
  NAND2_X1 U10495 ( .A1(n9182), .A2(n9181), .ZN(n9183) );
  XOR2_X1 U10496 ( .A(n9184), .B(n9183), .Z(n9187) );
  AOI222_X1 U10497 ( .A1(n9351), .A2(n9187), .B1(n9186), .B2(n9319), .C1(n9185), .C2(n9317), .ZN(n9378) );
  NOR2_X1 U10498 ( .A1(n9378), .A2(n9519), .ZN(n9188) );
  AOI211_X1 U10499 ( .C1(n9376), .C2(n9361), .A(n9189), .B(n9188), .ZN(n9190)
         );
  OAI21_X1 U10500 ( .B1(n9379), .B2(n9340), .A(n9190), .ZN(P1_U3265) );
  XOR2_X1 U10501 ( .A(n9191), .B(n9193), .Z(n9384) );
  XOR2_X1 U10502 ( .A(n9193), .B(n9192), .Z(n9194) );
  OAI222_X1 U10503 ( .A1(n9502), .A2(n9196), .B1(n9501), .B2(n9195), .C1(n9194), .C2(n9497), .ZN(n9380) );
  AOI211_X1 U10504 ( .C1(n9382), .C2(n9210), .A(n9762), .B(n4757), .ZN(n9381)
         );
  NAND2_X1 U10505 ( .A1(n9381), .A2(n9515), .ZN(n9199) );
  AOI22_X1 U10506 ( .A1(n9197), .A2(n9508), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9312), .ZN(n9198) );
  OAI211_X1 U10507 ( .C1(n9200), .C2(n9357), .A(n9199), .B(n9198), .ZN(n9201)
         );
  AOI21_X1 U10508 ( .B1(n9380), .B2(n9338), .A(n9201), .ZN(n9202) );
  OAI21_X1 U10509 ( .B1(n9384), .B2(n9340), .A(n9202), .ZN(P1_U3266) );
  XNOR2_X1 U10510 ( .A(n9204), .B(n9203), .ZN(n9389) );
  AOI21_X1 U10511 ( .B1(n9206), .B2(n9205), .A(n4513), .ZN(n9207) );
  OAI222_X1 U10512 ( .A1(n9502), .A2(n9209), .B1(n9501), .B2(n9208), .C1(n9497), .C2(n9207), .ZN(n9385) );
  INV_X1 U10513 ( .A(n9221), .ZN(n9211) );
  AOI211_X1 U10514 ( .C1(n9387), .C2(n9211), .A(n9762), .B(n4752), .ZN(n9386)
         );
  NAND2_X1 U10515 ( .A1(n9386), .A2(n9515), .ZN(n9215) );
  INV_X1 U10516 ( .A(n9212), .ZN(n9213) );
  AOI22_X1 U10517 ( .A1(n9213), .A2(n9508), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9312), .ZN(n9214) );
  OAI211_X1 U10518 ( .C1(n9216), .C2(n9357), .A(n9215), .B(n9214), .ZN(n9217)
         );
  AOI21_X1 U10519 ( .B1(n9385), .B2(n9338), .A(n9217), .ZN(n9218) );
  OAI21_X1 U10520 ( .B1(n9389), .B2(n9340), .A(n9218), .ZN(P1_U3267) );
  XNOR2_X1 U10521 ( .A(n9220), .B(n9219), .ZN(n9394) );
  INV_X1 U10522 ( .A(n9237), .ZN(n9222) );
  AOI21_X1 U10523 ( .B1(n9390), .B2(n9222), .A(n9221), .ZN(n9391) );
  AOI22_X1 U10524 ( .A1(n9223), .A2(n9508), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9312), .ZN(n9224) );
  OAI21_X1 U10525 ( .B1(n9225), .B2(n9357), .A(n9224), .ZN(n9234) );
  INV_X1 U10526 ( .A(n9226), .ZN(n9228) );
  OAI211_X1 U10527 ( .C1(n9228), .C2(n4567), .A(n9227), .B(n9351), .ZN(n9232)
         );
  AOI22_X1 U10528 ( .A1(n9230), .A2(n9319), .B1(n9317), .B2(n9229), .ZN(n9231)
         );
  AND2_X1 U10529 ( .A1(n9232), .A2(n9231), .ZN(n9393) );
  NOR2_X1 U10530 ( .A1(n9393), .A2(n9312), .ZN(n9233) );
  AOI211_X1 U10531 ( .C1(n9391), .C2(n9361), .A(n9234), .B(n9233), .ZN(n9235)
         );
  OAI21_X1 U10532 ( .B1(n9394), .B2(n9340), .A(n9235), .ZN(P1_U3268) );
  XNOR2_X1 U10533 ( .A(n9236), .B(n9241), .ZN(n9399) );
  AOI21_X1 U10534 ( .B1(n9395), .B2(n9253), .A(n9237), .ZN(n9396) );
  AOI22_X1 U10535 ( .A1(n9238), .A2(n9508), .B1(n9312), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9239) );
  OAI21_X1 U10536 ( .B1(n4756), .B2(n9357), .A(n9239), .ZN(n9245) );
  XNOR2_X1 U10537 ( .A(n9240), .B(n9241), .ZN(n9243) );
  AOI222_X1 U10538 ( .A1(n9351), .A2(n9243), .B1(n9273), .B2(n9317), .C1(n9242), .C2(n9319), .ZN(n9398) );
  NOR2_X1 U10539 ( .A1(n9398), .A2(n9312), .ZN(n9244) );
  AOI211_X1 U10540 ( .C1(n9396), .C2(n9361), .A(n9245), .B(n9244), .ZN(n9246)
         );
  OAI21_X1 U10541 ( .B1(n9399), .B2(n9340), .A(n9246), .ZN(P1_U3269) );
  XNOR2_X1 U10542 ( .A(n9247), .B(n9248), .ZN(n9404) );
  AOI22_X1 U10543 ( .A1(n9402), .A2(n9509), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9312), .ZN(n9261) );
  XNOR2_X1 U10544 ( .A(n9249), .B(n9248), .ZN(n9250) );
  OAI222_X1 U10545 ( .A1(n9501), .A2(n9252), .B1(n9502), .B2(n9251), .C1(n9497), .C2(n9250), .ZN(n9400) );
  INV_X1 U10546 ( .A(n9253), .ZN(n9254) );
  AOI211_X1 U10547 ( .C1(n9402), .C2(n9264), .A(n9762), .B(n9254), .ZN(n9401)
         );
  INV_X1 U10548 ( .A(n9401), .ZN(n9258) );
  INV_X1 U10549 ( .A(n9255), .ZN(n9256) );
  OAI22_X1 U10550 ( .A1(n9258), .A2(n9257), .B1(n9294), .B2(n9256), .ZN(n9259)
         );
  OAI21_X1 U10551 ( .B1(n9400), .B2(n9259), .A(n9338), .ZN(n9260) );
  OAI211_X1 U10552 ( .C1(n9404), .C2(n9340), .A(n9261), .B(n9260), .ZN(
        P1_U3270) );
  XNOR2_X1 U10553 ( .A(n9263), .B(n9262), .ZN(n9409) );
  INV_X1 U10554 ( .A(n9280), .ZN(n9266) );
  INV_X1 U10555 ( .A(n9264), .ZN(n9265) );
  AOI21_X1 U10556 ( .B1(n9405), .B2(n9266), .A(n9265), .ZN(n9406) );
  AOI22_X1 U10557 ( .A1(n9312), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9508), .B2(
        n9267), .ZN(n9268) );
  OAI21_X1 U10558 ( .B1(n9269), .B2(n9357), .A(n9268), .ZN(n9277) );
  NAND2_X1 U10559 ( .A1(n9285), .A2(n9270), .ZN(n9272) );
  XNOR2_X1 U10560 ( .A(n9272), .B(n9271), .ZN(n9275) );
  AOI222_X1 U10561 ( .A1(n9351), .A2(n9275), .B1(n9274), .B2(n9317), .C1(n9273), .C2(n9319), .ZN(n9408) );
  NOR2_X1 U10562 ( .A1(n9408), .A2(n9312), .ZN(n9276) );
  AOI211_X1 U10563 ( .C1(n9406), .C2(n9361), .A(n9277), .B(n9276), .ZN(n9278)
         );
  OAI21_X1 U10564 ( .B1(n9409), .B2(n9340), .A(n9278), .ZN(P1_U3271) );
  XOR2_X1 U10565 ( .A(n9279), .B(n9284), .Z(n9414) );
  AOI21_X1 U10566 ( .B1(n9410), .B2(n9292), .A(n9280), .ZN(n9411) );
  AOI22_X1 U10567 ( .A1(n9519), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9508), .B2(
        n9281), .ZN(n9282) );
  OAI21_X1 U10568 ( .B1(n9283), .B2(n9357), .A(n9282), .ZN(n9289) );
  OAI21_X1 U10569 ( .B1(n4550), .B2(n4723), .A(n9285), .ZN(n9287) );
  AOI222_X1 U10570 ( .A1(n9351), .A2(n9287), .B1(n9286), .B2(n9319), .C1(
        n10326), .C2(n9317), .ZN(n9413) );
  NOR2_X1 U10571 ( .A1(n9413), .A2(n9519), .ZN(n9288) );
  AOI211_X1 U10572 ( .C1(n9411), .C2(n9361), .A(n9289), .B(n9288), .ZN(n9290)
         );
  OAI21_X1 U10573 ( .B1(n9414), .B2(n9340), .A(n9290), .ZN(P1_U3272) );
  XNOR2_X1 U10574 ( .A(n9291), .B(n9302), .ZN(n9419) );
  INV_X1 U10575 ( .A(n9292), .ZN(n9293) );
  AOI211_X1 U10576 ( .C1(n9417), .C2(n9308), .A(n9762), .B(n9293), .ZN(n9416)
         );
  NOR2_X1 U10577 ( .A1(n4749), .A2(n9357), .ZN(n9297) );
  OAI22_X1 U10578 ( .A1(n9338), .A2(n9114), .B1(n9295), .B2(n9294), .ZN(n9296)
         );
  AOI211_X1 U10579 ( .C1(n9416), .C2(n9515), .A(n9297), .B(n9296), .ZN(n9306)
         );
  INV_X1 U10580 ( .A(n9298), .ZN(n9300) );
  OAI21_X1 U10581 ( .B1(n9316), .B2(n9300), .A(n9299), .ZN(n9301) );
  XOR2_X1 U10582 ( .A(n9302), .B(n9301), .Z(n9303) );
  OAI222_X1 U10583 ( .A1(n9501), .A2(n9304), .B1(n9502), .B2(n9331), .C1(n9497), .C2(n9303), .ZN(n9415) );
  NAND2_X1 U10584 ( .A1(n9415), .A2(n9338), .ZN(n9305) );
  OAI211_X1 U10585 ( .C1(n9419), .C2(n9340), .A(n9306), .B(n9305), .ZN(
        P1_U3273) );
  XNOR2_X1 U10586 ( .A(n9307), .B(n9315), .ZN(n9424) );
  INV_X1 U10587 ( .A(n9308), .ZN(n9309) );
  AOI21_X1 U10588 ( .B1(n9420), .B2(n4751), .A(n9309), .ZN(n9421) );
  INV_X1 U10589 ( .A(n9310), .ZN(n9311) );
  AOI22_X1 U10590 ( .A1(n9312), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9508), .B2(
        n9311), .ZN(n9313) );
  OAI21_X1 U10591 ( .B1(n9314), .B2(n9357), .A(n9313), .ZN(n9322) );
  XNOR2_X1 U10592 ( .A(n9316), .B(n9315), .ZN(n9320) );
  AOI222_X1 U10593 ( .A1(n9351), .A2(n9320), .B1(n10326), .B2(n9319), .C1(
        n9318), .C2(n9317), .ZN(n9423) );
  NOR2_X1 U10594 ( .A1(n9423), .A2(n9519), .ZN(n9321) );
  AOI211_X1 U10595 ( .C1(n9421), .C2(n9361), .A(n9322), .B(n9321), .ZN(n9323)
         );
  OAI21_X1 U10596 ( .B1(n9424), .B2(n9340), .A(n9323), .ZN(P1_U3274) );
  AOI21_X1 U10597 ( .B1(n9327), .B2(n9325), .A(n9324), .ZN(n9326) );
  INV_X1 U10598 ( .A(n9326), .ZN(n9429) );
  XNOR2_X1 U10599 ( .A(n9328), .B(n9327), .ZN(n9329) );
  OAI222_X1 U10600 ( .A1(n9501), .A2(n9331), .B1(n9502), .B2(n9330), .C1(n9497), .C2(n9329), .ZN(n9425) );
  INV_X1 U10601 ( .A(n9427), .ZN(n9336) );
  AOI211_X1 U10602 ( .C1(n9427), .C2(n9352), .A(n9762), .B(n9332), .ZN(n9426)
         );
  NAND2_X1 U10603 ( .A1(n9426), .A2(n9515), .ZN(n9335) );
  AOI22_X1 U10604 ( .A1(n9519), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9508), .B2(
        n9333), .ZN(n9334) );
  OAI211_X1 U10605 ( .C1(n9336), .C2(n9357), .A(n9335), .B(n9334), .ZN(n9337)
         );
  AOI21_X1 U10606 ( .B1(n9425), .B2(n9338), .A(n9337), .ZN(n9339) );
  OAI21_X1 U10607 ( .B1(n9429), .B2(n9340), .A(n9339), .ZN(P1_U3275) );
  XNOR2_X1 U10608 ( .A(n9342), .B(n9341), .ZN(n9350) );
  OAI22_X1 U10609 ( .A1(n9344), .A2(n9502), .B1(n9501), .B2(n9343), .ZN(n9349)
         );
  XNOR2_X1 U10610 ( .A(n9346), .B(n9345), .ZN(n9434) );
  NOR2_X1 U10611 ( .A1(n9434), .A2(n9347), .ZN(n9348) );
  AOI211_X1 U10612 ( .C1(n9351), .C2(n9350), .A(n9349), .B(n9348), .ZN(n9433)
         );
  INV_X1 U10613 ( .A(n9352), .ZN(n9353) );
  AOI21_X1 U10614 ( .B1(n9430), .B2(n9354), .A(n9353), .ZN(n9431) );
  AOI22_X1 U10615 ( .A1(n9312), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9508), .B2(
        n9355), .ZN(n9356) );
  OAI21_X1 U10616 ( .B1(n5329), .B2(n9357), .A(n9356), .ZN(n9360) );
  NOR2_X1 U10617 ( .A1(n9434), .A2(n9358), .ZN(n9359) );
  AOI211_X1 U10618 ( .C1(n9431), .C2(n9361), .A(n9360), .B(n9359), .ZN(n9362)
         );
  OAI21_X1 U10619 ( .B1(n9433), .B2(n9519), .A(n9362), .ZN(P1_U3276) );
  NAND2_X1 U10620 ( .A1(n8876), .A2(n9750), .ZN(n9363) );
  OAI211_X1 U10621 ( .C1(n9364), .C2(n9762), .A(n9529), .B(n9363), .ZN(n9435)
         );
  MUX2_X1 U10622 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9435), .S(n9781), .Z(
        P1_U3554) );
  MUX2_X1 U10623 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9436), .S(n9781), .Z(
        P1_U3552) );
  MUX2_X1 U10624 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9369), .S(n9781), .Z(
        P1_U3551) );
  AOI22_X1 U10625 ( .A1(n9371), .A2(n9751), .B1(n9750), .B2(n9370), .ZN(n9372)
         );
  OAI211_X1 U10626 ( .C1(n9374), .C2(n9534), .A(n9373), .B(n9372), .ZN(n9437)
         );
  MUX2_X1 U10627 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9437), .S(n9781), .Z(
        P1_U3550) );
  AOI22_X1 U10628 ( .A1(n9376), .A2(n9751), .B1(n9750), .B2(n9375), .ZN(n9377)
         );
  OAI211_X1 U10629 ( .C1(n9379), .C2(n9534), .A(n9378), .B(n9377), .ZN(n9438)
         );
  MUX2_X1 U10630 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9438), .S(n9781), .Z(
        P1_U3549) );
  AOI211_X1 U10631 ( .C1(n9750), .C2(n9382), .A(n9381), .B(n9380), .ZN(n9383)
         );
  OAI21_X1 U10632 ( .B1(n9384), .B2(n9534), .A(n9383), .ZN(n9439) );
  MUX2_X1 U10633 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9439), .S(n9781), .Z(
        P1_U3548) );
  AOI211_X1 U10634 ( .C1(n9750), .C2(n9387), .A(n9386), .B(n9385), .ZN(n9388)
         );
  OAI21_X1 U10635 ( .B1(n9389), .B2(n9534), .A(n9388), .ZN(n9440) );
  MUX2_X1 U10636 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9440), .S(n9781), .Z(
        P1_U3547) );
  AOI22_X1 U10637 ( .A1(n9391), .A2(n9751), .B1(n9750), .B2(n9390), .ZN(n9392)
         );
  OAI211_X1 U10638 ( .C1(n9394), .C2(n9534), .A(n9393), .B(n9392), .ZN(n9441)
         );
  MUX2_X1 U10639 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9441), .S(n9781), .Z(
        P1_U3546) );
  AOI22_X1 U10640 ( .A1(n9396), .A2(n9751), .B1(n9750), .B2(n9395), .ZN(n9397)
         );
  OAI211_X1 U10641 ( .C1(n9399), .C2(n9534), .A(n9398), .B(n9397), .ZN(n9442)
         );
  MUX2_X1 U10642 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9442), .S(n9781), .Z(
        P1_U3545) );
  AOI211_X1 U10643 ( .C1(n9750), .C2(n9402), .A(n9401), .B(n9400), .ZN(n9403)
         );
  OAI21_X1 U10644 ( .B1(n9404), .B2(n9534), .A(n9403), .ZN(n9443) );
  MUX2_X1 U10645 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9443), .S(n9781), .Z(
        P1_U3544) );
  AOI22_X1 U10646 ( .A1(n9406), .A2(n9751), .B1(n9750), .B2(n9405), .ZN(n9407)
         );
  OAI211_X1 U10647 ( .C1(n9409), .C2(n9534), .A(n9408), .B(n9407), .ZN(n9444)
         );
  MUX2_X1 U10648 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9444), .S(n9781), .Z(
        P1_U3543) );
  AOI22_X1 U10649 ( .A1(n9411), .A2(n9751), .B1(n9750), .B2(n9410), .ZN(n9412)
         );
  OAI211_X1 U10650 ( .C1(n9414), .C2(n9534), .A(n9413), .B(n9412), .ZN(n9445)
         );
  MUX2_X1 U10651 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9445), .S(n9781), .Z(
        P1_U3542) );
  AOI211_X1 U10652 ( .C1(n9750), .C2(n9417), .A(n9416), .B(n9415), .ZN(n9418)
         );
  OAI21_X1 U10653 ( .B1(n9419), .B2(n9534), .A(n9418), .ZN(n9446) );
  MUX2_X1 U10654 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9446), .S(n9781), .Z(
        P1_U3541) );
  AOI22_X1 U10655 ( .A1(n9421), .A2(n9751), .B1(n9750), .B2(n9420), .ZN(n9422)
         );
  OAI211_X1 U10656 ( .C1(n9424), .C2(n9534), .A(n9423), .B(n9422), .ZN(n9447)
         );
  MUX2_X1 U10657 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9447), .S(n9781), .Z(
        P1_U3540) );
  AOI211_X1 U10658 ( .C1(n9750), .C2(n9427), .A(n9426), .B(n9425), .ZN(n9428)
         );
  OAI21_X1 U10659 ( .B1(n9429), .B2(n9534), .A(n9428), .ZN(n9448) );
  MUX2_X1 U10660 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9448), .S(n9781), .Z(
        P1_U3539) );
  AOI22_X1 U10661 ( .A1(n9431), .A2(n9751), .B1(n9750), .B2(n9430), .ZN(n9432)
         );
  OAI211_X1 U10662 ( .C1(n9756), .C2(n9434), .A(n9433), .B(n9432), .ZN(n9449)
         );
  MUX2_X1 U10663 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9449), .S(n9781), .Z(
        P1_U3538) );
  MUX2_X1 U10664 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9435), .S(n9759), .Z(
        P1_U3522) );
  MUX2_X1 U10665 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9436), .S(n9759), .Z(
        P1_U3520) );
  MUX2_X1 U10666 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9437), .S(n9759), .Z(
        P1_U3518) );
  MUX2_X1 U10667 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9438), .S(n9759), .Z(
        P1_U3517) );
  MUX2_X1 U10668 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9439), .S(n9759), .Z(
        P1_U3516) );
  MUX2_X1 U10669 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9440), .S(n9759), .Z(
        P1_U3515) );
  MUX2_X1 U10670 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9441), .S(n9759), .Z(
        P1_U3514) );
  MUX2_X1 U10671 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9442), .S(n9759), .Z(
        P1_U3513) );
  MUX2_X1 U10672 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9443), .S(n9759), .Z(
        P1_U3512) );
  MUX2_X1 U10673 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9444), .S(n9759), .Z(
        P1_U3511) );
  MUX2_X1 U10674 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9445), .S(n9759), .Z(
        P1_U3510) );
  MUX2_X1 U10675 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9446), .S(n9759), .Z(
        P1_U3508) );
  MUX2_X1 U10676 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9447), .S(n9759), .Z(
        P1_U3505) );
  MUX2_X1 U10677 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9448), .S(n9759), .Z(
        P1_U3502) );
  MUX2_X1 U10678 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9449), .S(n9759), .Z(
        P1_U3499) );
  MUX2_X1 U10679 ( .A(P1_D_REG_0__SCAN_IN), .B(n9450), .S(n9722), .Z(P1_U3440)
         );
  NOR4_X1 U10680 ( .A1(n9452), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n9451), .ZN(n9453) );
  AOI21_X1 U10681 ( .B1(n9463), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9453), .ZN(
        n9454) );
  OAI21_X1 U10682 ( .B1(n9455), .B2(n9460), .A(n9454), .ZN(P1_U3322) );
  AOI22_X1 U10683 ( .A1(n5395), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9463), .ZN(n9456) );
  OAI21_X1 U10684 ( .B1(n9457), .B2(n9460), .A(n9456), .ZN(P1_U3323) );
  AOI22_X1 U10685 ( .A1(n9458), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n9463), .ZN(n9459) );
  OAI21_X1 U10686 ( .B1(n9461), .B2(n9460), .A(n9459), .ZN(P1_U3324) );
  INV_X1 U10687 ( .A(n9462), .ZN(n9465) );
  AOI22_X1 U10688 ( .A1(n9572), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n9463), .ZN(n9464) );
  OAI21_X1 U10689 ( .B1(n9465), .B2(n9460), .A(n9464), .ZN(P1_U3325) );
  MUX2_X1 U10690 ( .A(n9466), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI22_X1 U10691 ( .A1(n9788), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n9477) );
  NAND2_X1 U10692 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9469) );
  AOI211_X1 U10693 ( .C1(n9469), .C2(n9468), .A(n9467), .B(n9786), .ZN(n9470)
         );
  AOI21_X1 U10694 ( .B1(n9483), .B2(n4461), .A(n9470), .ZN(n9476) );
  INV_X1 U10695 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10272) );
  NOR2_X1 U10696 ( .A1(n9791), .A2(n10272), .ZN(n9474) );
  OAI211_X1 U10697 ( .C1(n9474), .C2(n9473), .A(n9783), .B(n9472), .ZN(n9475)
         );
  NAND3_X1 U10698 ( .A1(n9477), .A2(n9476), .A3(n9475), .ZN(P2_U3246) );
  AOI22_X1 U10699 ( .A1(n9788), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9489) );
  AOI211_X1 U10700 ( .C1(n9480), .C2(n9479), .A(n9478), .B(n9786), .ZN(n9481)
         );
  AOI21_X1 U10701 ( .B1(n9483), .B2(n9482), .A(n9481), .ZN(n9488) );
  OAI211_X1 U10702 ( .C1(n9486), .C2(n9485), .A(n9783), .B(n9484), .ZN(n9487)
         );
  NAND3_X1 U10703 ( .A1(n9489), .A2(n9488), .A3(n9487), .ZN(P2_U3247) );
  XNOR2_X1 U10704 ( .A(n9490), .B(n9492), .ZN(n9525) );
  INV_X1 U10705 ( .A(n9491), .ZN(n9499) );
  INV_X1 U10706 ( .A(n9492), .ZN(n9493) );
  AOI21_X1 U10707 ( .B1(n9495), .B2(n9494), .A(n9493), .ZN(n9496) );
  AOI211_X1 U10708 ( .C1(n9499), .C2(n9498), .A(n9497), .B(n9496), .ZN(n9505)
         );
  OAI22_X1 U10709 ( .A1(n9503), .A2(n9502), .B1(n9501), .B2(n9500), .ZN(n9504)
         );
  AOI211_X1 U10710 ( .C1(n9525), .C2(n9506), .A(n9505), .B(n9504), .ZN(n9522)
         );
  AOI222_X1 U10711 ( .A1(n9510), .A2(n9509), .B1(P1_REG2_REG_10__SCAN_IN), 
        .B2(n9519), .C1(n9508), .C2(n9507), .ZN(n9518) );
  INV_X1 U10712 ( .A(n9511), .ZN(n9513) );
  OAI211_X1 U10713 ( .C1(n9513), .C2(n9521), .A(n9751), .B(n9512), .ZN(n9520)
         );
  INV_X1 U10714 ( .A(n9520), .ZN(n9514) );
  AOI22_X1 U10715 ( .A1(n9525), .A2(n9516), .B1(n9515), .B2(n9514), .ZN(n9517)
         );
  OAI211_X1 U10716 ( .C1(n9519), .C2(n9522), .A(n9518), .B(n9517), .ZN(
        P1_U3281) );
  OAI21_X1 U10717 ( .B1(n9521), .B2(n9760), .A(n9520), .ZN(n9524) );
  INV_X1 U10718 ( .A(n9522), .ZN(n9523) );
  AOI211_X1 U10719 ( .C1(n9767), .C2(n9525), .A(n9524), .B(n9523), .ZN(n9528)
         );
  INV_X1 U10720 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9526) );
  AOI22_X1 U10721 ( .A1(n9759), .A2(n9528), .B1(n9526), .B2(n9768), .ZN(
        P1_U3484) );
  AOI22_X1 U10722 ( .A1(n9781), .A2(n9528), .B1(n9527), .B2(n9779), .ZN(
        P1_U3533) );
  OAI21_X1 U10723 ( .B1(n9530), .B2(n9760), .A(n9529), .ZN(n9531) );
  AOI21_X1 U10724 ( .B1(n9532), .B2(n9751), .A(n9531), .ZN(n9563) );
  INV_X1 U10725 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9533) );
  AOI22_X1 U10726 ( .A1(n9781), .A2(n9563), .B1(n9533), .B2(n9779), .ZN(
        P1_U3553) );
  OAI211_X1 U10727 ( .C1(n9537), .C2(n9760), .A(n9536), .B(n9535), .ZN(n9538)
         );
  AOI21_X1 U10728 ( .B1(n9539), .B2(n5675), .A(n9538), .ZN(n9565) );
  AOI22_X1 U10729 ( .A1(n9781), .A2(n9565), .B1(n9540), .B2(n9779), .ZN(
        P1_U3537) );
  OAI22_X1 U10730 ( .A1(n9542), .A2(n9762), .B1(n9541), .B2(n9760), .ZN(n9543)
         );
  AOI21_X1 U10731 ( .B1(n9544), .B2(n9767), .A(n9543), .ZN(n9545) );
  AOI22_X1 U10732 ( .A1(n9781), .A2(n9567), .B1(n9547), .B2(n9779), .ZN(
        P1_U3536) );
  OAI21_X1 U10733 ( .B1(n9549), .B2(n9760), .A(n9548), .ZN(n9550) );
  AOI21_X1 U10734 ( .B1(n9551), .B2(n9767), .A(n9550), .ZN(n9552) );
  AND2_X1 U10735 ( .A1(n9553), .A2(n9552), .ZN(n9569) );
  AOI22_X1 U10736 ( .A1(n9781), .A2(n9569), .B1(n9554), .B2(n9779), .ZN(
        P1_U3535) );
  INV_X1 U10737 ( .A(n9555), .ZN(n9556) );
  OAI22_X1 U10738 ( .A1(n9557), .A2(n9762), .B1(n9556), .B2(n9760), .ZN(n9558)
         );
  AOI21_X1 U10739 ( .B1(n9559), .B2(n9767), .A(n9558), .ZN(n9560) );
  AND2_X1 U10740 ( .A1(n9561), .A2(n9560), .ZN(n9571) );
  AOI22_X1 U10741 ( .A1(n9781), .A2(n9571), .B1(n6503), .B2(n9779), .ZN(
        P1_U3534) );
  INV_X1 U10742 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9562) );
  AOI22_X1 U10743 ( .A1(n9759), .A2(n9563), .B1(n9562), .B2(n9768), .ZN(
        P1_U3521) );
  INV_X1 U10744 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9564) );
  AOI22_X1 U10745 ( .A1(n9759), .A2(n9565), .B1(n9564), .B2(n9768), .ZN(
        P1_U3496) );
  INV_X1 U10746 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9566) );
  AOI22_X1 U10747 ( .A1(n9759), .A2(n9567), .B1(n9566), .B2(n9768), .ZN(
        P1_U3493) );
  INV_X1 U10748 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9568) );
  AOI22_X1 U10749 ( .A1(n9759), .A2(n9569), .B1(n9568), .B2(n9768), .ZN(
        P1_U3490) );
  INV_X1 U10750 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9570) );
  AOI22_X1 U10751 ( .A1(n9759), .A2(n9571), .B1(n9570), .B2(n9768), .ZN(
        P1_U3487) );
  XNOR2_X1 U10752 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X1 U10753 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10143) );
  AOI211_X1 U10754 ( .C1(n9572), .C2(P1_REG2_REG_0__SCAN_IN), .A(
        P1_IR_REG_0__SCAN_IN), .B(n9589), .ZN(n9590) );
  INV_X1 U10755 ( .A(n9591), .ZN(n9575) );
  OAI21_X1 U10756 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n9578), .A(n9572), .ZN(
        n9573) );
  AOI21_X1 U10757 ( .B1(n9575), .B2(n9574), .A(n9573), .ZN(n9576) );
  OAI21_X1 U10758 ( .B1(n9590), .B2(n9576), .A(P1_STATE_REG_SCAN_IN), .ZN(
        n9577) );
  OAI211_X1 U10759 ( .C1(P1_STATE_REG_SCAN_IN), .C2(P1_REG3_REG_0__SCAN_IN), 
        .A(n9577), .B(P1_U3083), .ZN(n9580) );
  NAND3_X1 U10760 ( .A1(n9693), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9578), .ZN(
        n9579) );
  OAI211_X1 U10761 ( .C1(n10143), .C2(n9716), .A(n9580), .B(n9579), .ZN(
        P1_U3241) );
  XNOR2_X1 U10762 ( .A(n9582), .B(n9581), .ZN(n9598) );
  NAND2_X1 U10763 ( .A1(P1_U3084), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9587) );
  OAI211_X1 U10764 ( .C1(n9585), .C2(n9584), .A(n9693), .B(n9583), .ZN(n9586)
         );
  OAI211_X1 U10765 ( .C1(n9691), .C2(n9588), .A(n9587), .B(n9586), .ZN(n9597)
         );
  INV_X1 U10766 ( .A(n9589), .ZN(n9594) );
  AOI211_X1 U10767 ( .C1(n9592), .C2(n9591), .A(n9100), .B(n9590), .ZN(n9593)
         );
  OAI21_X1 U10768 ( .B1(n9595), .B2(n9594), .A(n9593), .ZN(n9615) );
  INV_X1 U10769 ( .A(n9615), .ZN(n9596) );
  AOI211_X1 U10770 ( .C1(n9687), .C2(n9598), .A(n9597), .B(n9596), .ZN(n9599)
         );
  OAI21_X1 U10771 ( .B1(n9716), .B2(n9600), .A(n9599), .ZN(P1_U3243) );
  AOI21_X1 U10772 ( .B1(n9603), .B2(n9602), .A(n9601), .ZN(n9604) );
  INV_X1 U10773 ( .A(n9604), .ZN(n9605) );
  NAND2_X1 U10774 ( .A1(n9687), .A2(n9605), .ZN(n9612) );
  OAI21_X1 U10775 ( .B1(n9608), .B2(n9607), .A(n9606), .ZN(n9610) );
  AOI21_X1 U10776 ( .B1(n9693), .B2(n9610), .A(n9609), .ZN(n9611) );
  OAI211_X1 U10777 ( .C1(n9691), .C2(n9613), .A(n9612), .B(n9611), .ZN(n9614)
         );
  INV_X1 U10778 ( .A(n9614), .ZN(n9616) );
  OAI211_X1 U10779 ( .C1(n9617), .C2(n9716), .A(n9616), .B(n9615), .ZN(
        P1_U3245) );
  INV_X1 U10780 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9631) );
  OAI211_X1 U10781 ( .C1(n9620), .C2(n9619), .A(n9687), .B(n9618), .ZN(n9621)
         );
  INV_X1 U10782 ( .A(n9621), .ZN(n9622) );
  AOI211_X1 U10783 ( .C1(n9707), .C2(n9624), .A(n9623), .B(n9622), .ZN(n9630)
         );
  AOI21_X1 U10784 ( .B1(n9627), .B2(n9626), .A(n9625), .ZN(n9628) );
  OR2_X1 U10785 ( .A1(n9712), .A2(n9628), .ZN(n9629) );
  OAI211_X1 U10786 ( .C1(n9631), .C2(n9716), .A(n9630), .B(n9629), .ZN(
        P1_U3253) );
  INV_X1 U10787 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9645) );
  NOR2_X1 U10788 ( .A1(n9633), .A2(n9632), .ZN(n9634) );
  NOR3_X1 U10789 ( .A1(n9701), .A2(n9635), .A3(n9634), .ZN(n9636) );
  AOI211_X1 U10790 ( .C1(n9707), .C2(n9638), .A(n9637), .B(n9636), .ZN(n9644)
         );
  AOI21_X1 U10791 ( .B1(n9641), .B2(n9640), .A(n9639), .ZN(n9642) );
  OR2_X1 U10792 ( .A1(n9642), .A2(n9712), .ZN(n9643) );
  OAI211_X1 U10793 ( .C1(n9645), .C2(n9716), .A(n9644), .B(n9643), .ZN(
        P1_U3254) );
  INV_X1 U10794 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9661) );
  AOI21_X1 U10795 ( .B1(n9648), .B2(n9647), .A(n9646), .ZN(n9649) );
  NAND2_X1 U10796 ( .A1(n9687), .A2(n9649), .ZN(n9652) );
  INV_X1 U10797 ( .A(n9650), .ZN(n9651) );
  OAI211_X1 U10798 ( .C1(n9691), .C2(n9653), .A(n9652), .B(n9651), .ZN(n9654)
         );
  INV_X1 U10799 ( .A(n9654), .ZN(n9660) );
  AOI21_X1 U10800 ( .B1(n9657), .B2(n9656), .A(n9655), .ZN(n9658) );
  OR2_X1 U10801 ( .A1(n9658), .A2(n9712), .ZN(n9659) );
  OAI211_X1 U10802 ( .C1(n9661), .C2(n9716), .A(n9660), .B(n9659), .ZN(
        P1_U3255) );
  INV_X1 U10803 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10255) );
  AOI211_X1 U10804 ( .C1(n9664), .C2(n9663), .A(n9662), .B(n9701), .ZN(n9665)
         );
  AOI211_X1 U10805 ( .C1(n9707), .C2(n9667), .A(n9666), .B(n9665), .ZN(n9671)
         );
  OAI211_X1 U10806 ( .C1(n9669), .C2(P1_REG1_REG_15__SCAN_IN), .A(n9693), .B(
        n9668), .ZN(n9670) );
  OAI211_X1 U10807 ( .C1(n10255), .C2(n9716), .A(n9671), .B(n9670), .ZN(
        P1_U3256) );
  INV_X1 U10808 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9682) );
  AOI211_X1 U10809 ( .C1(n4551), .C2(n9673), .A(n9672), .B(n9701), .ZN(n9674)
         );
  AOI211_X1 U10810 ( .C1(n9707), .C2(n9676), .A(n9675), .B(n9674), .ZN(n9681)
         );
  OAI211_X1 U10811 ( .C1(n9679), .C2(n9678), .A(n9693), .B(n9677), .ZN(n9680)
         );
  OAI211_X1 U10812 ( .C1(n9682), .C2(n9716), .A(n9681), .B(n9680), .ZN(
        P1_U3257) );
  INV_X1 U10813 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9699) );
  AOI21_X1 U10814 ( .B1(n9685), .B2(n9684), .A(n9683), .ZN(n9686) );
  NAND2_X1 U10815 ( .A1(n9687), .A2(n9686), .ZN(n9689) );
  OAI211_X1 U10816 ( .C1(n9691), .C2(n9690), .A(n9689), .B(n9688), .ZN(n9692)
         );
  INV_X1 U10817 ( .A(n9692), .ZN(n9698) );
  OAI211_X1 U10818 ( .C1(n9696), .C2(n9695), .A(n9694), .B(n9693), .ZN(n9697)
         );
  OAI211_X1 U10819 ( .C1(n9699), .C2(n9716), .A(n9698), .B(n9697), .ZN(
        P1_U3258) );
  INV_X1 U10820 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10338) );
  INV_X1 U10821 ( .A(n9700), .ZN(n9706) );
  AOI211_X1 U10822 ( .C1(n9704), .C2(n9703), .A(n9702), .B(n9701), .ZN(n9705)
         );
  AOI211_X1 U10823 ( .C1(n9708), .C2(n9707), .A(n9706), .B(n9705), .ZN(n9715)
         );
  AOI21_X1 U10824 ( .B1(n9711), .B2(n9710), .A(n9709), .ZN(n9713) );
  OR2_X1 U10825 ( .A1(n9713), .A2(n9712), .ZN(n9714) );
  OAI211_X1 U10826 ( .C1(n10338), .C2(n9716), .A(n9715), .B(n9714), .ZN(
        P1_U3259) );
  AND2_X1 U10827 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9719), .ZN(P1_U3292) );
  AND2_X1 U10828 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9719), .ZN(P1_U3293) );
  AND2_X1 U10829 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9719), .ZN(P1_U3294) );
  AND2_X1 U10830 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9719), .ZN(P1_U3295) );
  AND2_X1 U10831 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9719), .ZN(P1_U3296) );
  AND2_X1 U10832 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9719), .ZN(P1_U3297) );
  AND2_X1 U10833 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9719), .ZN(P1_U3298) );
  AND2_X1 U10834 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9719), .ZN(P1_U3299) );
  AND2_X1 U10835 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9719), .ZN(P1_U3300) );
  AND2_X1 U10836 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9719), .ZN(P1_U3301) );
  INV_X1 U10837 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10182) );
  NOR2_X1 U10838 ( .A1(n9718), .A2(n10182), .ZN(P1_U3302) );
  AND2_X1 U10839 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9719), .ZN(P1_U3303) );
  AND2_X1 U10840 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9719), .ZN(P1_U3304) );
  AND2_X1 U10841 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9719), .ZN(P1_U3305) );
  AND2_X1 U10842 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9719), .ZN(P1_U3306) );
  AND2_X1 U10843 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9719), .ZN(P1_U3307) );
  AND2_X1 U10844 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9719), .ZN(P1_U3308) );
  AND2_X1 U10845 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9719), .ZN(P1_U3309) );
  AND2_X1 U10846 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9719), .ZN(P1_U3310) );
  AND2_X1 U10847 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9719), .ZN(P1_U3311) );
  AND2_X1 U10848 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9719), .ZN(P1_U3312) );
  AND2_X1 U10849 ( .A1(n9719), .A2(P1_D_REG_10__SCAN_IN), .ZN(P1_U3313) );
  AND2_X1 U10850 ( .A1(n9719), .A2(P1_D_REG_9__SCAN_IN), .ZN(P1_U3314) );
  INV_X1 U10851 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10192) );
  NOR2_X1 U10852 ( .A1(n9718), .A2(n10192), .ZN(P1_U3315) );
  AND2_X1 U10853 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9719), .ZN(P1_U3316) );
  AND2_X1 U10854 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9719), .ZN(P1_U3317) );
  AND2_X1 U10855 ( .A1(n9719), .A2(P1_D_REG_5__SCAN_IN), .ZN(P1_U3318) );
  AND2_X1 U10856 ( .A1(n9719), .A2(P1_D_REG_4__SCAN_IN), .ZN(P1_U3319) );
  INV_X1 U10857 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10268) );
  NOR2_X1 U10858 ( .A1(n9718), .A2(n10268), .ZN(P1_U3320) );
  AND2_X1 U10859 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9719), .ZN(P1_U3321) );
  INV_X1 U10860 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9721) );
  OAI21_X1 U10861 ( .B1(n9722), .B2(n9721), .A(n9720), .ZN(P1_U3441) );
  INV_X1 U10862 ( .A(n9723), .ZN(n9728) );
  OAI21_X1 U10863 ( .B1(n9725), .B2(n9760), .A(n9724), .ZN(n9727) );
  AOI211_X1 U10864 ( .C1(n9767), .C2(n9728), .A(n9727), .B(n9726), .ZN(n9771)
         );
  AOI22_X1 U10865 ( .A1(n9759), .A2(n9771), .B1(n5398), .B2(n9768), .ZN(
        P1_U3457) );
  NAND3_X1 U10866 ( .A1(n9730), .A2(n9751), .A3(n9729), .ZN(n9731) );
  OAI21_X1 U10867 ( .B1(n9732), .B2(n9760), .A(n9731), .ZN(n9734) );
  AOI211_X1 U10868 ( .C1(n9767), .C2(n9735), .A(n9734), .B(n9733), .ZN(n9773)
         );
  AOI22_X1 U10869 ( .A1(n9759), .A2(n9773), .B1(n5408), .B2(n9768), .ZN(
        P1_U3460) );
  OAI22_X1 U10870 ( .A1(n9737), .A2(n9762), .B1(n9736), .B2(n9760), .ZN(n9739)
         );
  AOI211_X1 U10871 ( .C1(n9767), .C2(n9740), .A(n9739), .B(n9738), .ZN(n9775)
         );
  INV_X1 U10872 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9741) );
  AOI22_X1 U10873 ( .A1(n9759), .A2(n9775), .B1(n9741), .B2(n9768), .ZN(
        P1_U3466) );
  AOI22_X1 U10874 ( .A1(n9743), .A2(n9751), .B1(n9750), .B2(n9742), .ZN(n9744)
         );
  OAI211_X1 U10875 ( .C1(n9746), .C2(n9756), .A(n9745), .B(n9744), .ZN(n9747)
         );
  INV_X1 U10876 ( .A(n9747), .ZN(n9776) );
  INV_X1 U10877 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9748) );
  AOI22_X1 U10878 ( .A1(n9759), .A2(n9776), .B1(n9748), .B2(n9768), .ZN(
        P1_U3472) );
  AOI22_X1 U10879 ( .A1(n9752), .A2(n9751), .B1(n9750), .B2(n9749), .ZN(n9753)
         );
  OAI211_X1 U10880 ( .C1(n9756), .C2(n9755), .A(n9754), .B(n9753), .ZN(n9757)
         );
  INV_X1 U10881 ( .A(n9757), .ZN(n9778) );
  INV_X1 U10882 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9758) );
  AOI22_X1 U10883 ( .A1(n9759), .A2(n9778), .B1(n9758), .B2(n9768), .ZN(
        P1_U3478) );
  OAI22_X1 U10884 ( .A1(n9763), .A2(n9762), .B1(n9761), .B2(n9760), .ZN(n9765)
         );
  AOI211_X1 U10885 ( .C1(n9767), .C2(n9766), .A(n9765), .B(n9764), .ZN(n9780)
         );
  INV_X1 U10886 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9769) );
  AOI22_X1 U10887 ( .A1(n9759), .A2(n9780), .B1(n9769), .B2(n9768), .ZN(
        P1_U3481) );
  AOI22_X1 U10888 ( .A1(n9781), .A2(n9771), .B1(n9770), .B2(n9779), .ZN(
        P1_U3524) );
  INV_X1 U10889 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9772) );
  AOI22_X1 U10890 ( .A1(n9781), .A2(n9773), .B1(n9772), .B2(n9779), .ZN(
        P1_U3525) );
  INV_X1 U10891 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9774) );
  AOI22_X1 U10892 ( .A1(n9781), .A2(n9775), .B1(n9774), .B2(n9779), .ZN(
        P1_U3527) );
  AOI22_X1 U10893 ( .A1(n9781), .A2(n9776), .B1(n6288), .B2(n9779), .ZN(
        P1_U3529) );
  AOI22_X1 U10894 ( .A1(n9781), .A2(n9778), .B1(n9777), .B2(n9779), .ZN(
        P1_U3531) );
  AOI22_X1 U10895 ( .A1(n9781), .A2(n9780), .B1(n10207), .B2(n9779), .ZN(
        P1_U3532) );
  AOI22_X1 U10896 ( .A1(n9782), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9783), .ZN(n9792) );
  NAND2_X1 U10897 ( .A1(n9783), .A2(n10272), .ZN(n9784) );
  OAI211_X1 U10898 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n9786), .A(n9785), .B(
        n9784), .ZN(n9787) );
  INV_X1 U10899 ( .A(n9787), .ZN(n9790) );
  AOI22_X1 U10900 ( .A1(n9788), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9789) );
  OAI221_X1 U10901 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9792), .C1(n9791), .C2(
        n9790), .A(n9789), .ZN(P2_U3245) );
  AND2_X1 U10902 ( .A1(n9794), .A2(n9793), .ZN(n9795) );
  OR2_X1 U10903 ( .A1(n9796), .A2(n9795), .ZN(n9809) );
  NAND2_X1 U10904 ( .A1(n9798), .A2(n9797), .ZN(n9799) );
  NAND2_X1 U10905 ( .A1(n9800), .A2(n9799), .ZN(n9880) );
  OAI22_X1 U10906 ( .A1(n9809), .A2(n9801), .B1(n9836), .B2(n9880), .ZN(n9802)
         );
  INV_X1 U10907 ( .A(n9802), .ZN(n9819) );
  AOI21_X1 U10908 ( .B1(n9804), .B2(n9803), .A(n4562), .ZN(n9814) );
  AOI22_X1 U10909 ( .A1(n9808), .A2(n9807), .B1(n9806), .B2(n9805), .ZN(n9812)
         );
  INV_X1 U10910 ( .A(n9809), .ZN(n9883) );
  NAND2_X1 U10911 ( .A1(n9883), .A2(n9810), .ZN(n9811) );
  OAI211_X1 U10912 ( .C1(n9814), .C2(n9813), .A(n9812), .B(n9811), .ZN(n9881)
         );
  AOI22_X1 U10913 ( .A1(n9842), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n9815), .B2(
        n9838), .ZN(n9816) );
  OAI21_X1 U10914 ( .B1(n9879), .B2(n9835), .A(n9816), .ZN(n9817) );
  AOI21_X1 U10915 ( .B1(n9881), .B2(n9840), .A(n9817), .ZN(n9818) );
  NAND2_X1 U10916 ( .A1(n9819), .A2(n9818), .ZN(P2_U3288) );
  AOI22_X1 U10917 ( .A1(n9838), .A2(n10240), .B1(P2_REG2_REG_3__SCAN_IN), .B2(
        n9842), .ZN(n9829) );
  NAND2_X1 U10918 ( .A1(n9821), .A2(n9820), .ZN(n9825) );
  NAND2_X1 U10919 ( .A1(n9823), .A2(n9822), .ZN(n9824) );
  OAI211_X1 U10920 ( .C1(n9826), .C2(n9835), .A(n9825), .B(n9824), .ZN(n9827)
         );
  INV_X1 U10921 ( .A(n9827), .ZN(n9828) );
  OAI211_X1 U10922 ( .C1(n9842), .C2(n9830), .A(n9829), .B(n9828), .ZN(
        P2_U3293) );
  NOR2_X1 U10923 ( .A1(n9832), .A2(n9831), .ZN(n9854) );
  INV_X1 U10924 ( .A(n9854), .ZN(n9856) );
  OR2_X1 U10925 ( .A1(n9833), .A2(n9857), .ZN(n9834) );
  AOI21_X1 U10926 ( .B1(n9856), .B2(n9834), .A(n9851), .ZN(n9841) );
  AOI21_X1 U10927 ( .B1(n9836), .B2(n9835), .A(n4690), .ZN(n9837) );
  AOI21_X1 U10928 ( .B1(n9838), .B2(P2_REG3_REG_0__SCAN_IN), .A(n9837), .ZN(
        n9839) );
  OAI221_X1 U10929 ( .B1(n9842), .B2(n9841), .C1(n9840), .C2(n10075), .A(n9839), .ZN(P2_U3296) );
  AND2_X1 U10930 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9848), .ZN(P2_U3297) );
  AND2_X1 U10931 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9848), .ZN(P2_U3298) );
  AND2_X1 U10932 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9848), .ZN(P2_U3299) );
  AND2_X1 U10933 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9848), .ZN(P2_U3300) );
  AND2_X1 U10934 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9848), .ZN(P2_U3301) );
  AND2_X1 U10935 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9848), .ZN(P2_U3302) );
  AND2_X1 U10936 ( .A1(n9848), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3303) );
  AND2_X1 U10937 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9848), .ZN(P2_U3304) );
  AND2_X1 U10938 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9848), .ZN(P2_U3305) );
  AND2_X1 U10939 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9848), .ZN(P2_U3306) );
  AND2_X1 U10940 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9848), .ZN(P2_U3307) );
  AND2_X1 U10941 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9848), .ZN(P2_U3308) );
  AND2_X1 U10942 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9848), .ZN(P2_U3309) );
  AND2_X1 U10943 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9848), .ZN(P2_U3310) );
  AND2_X1 U10944 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9848), .ZN(P2_U3311) );
  INV_X1 U10945 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n10084) );
  NOR2_X1 U10946 ( .A1(n9845), .A2(n10084), .ZN(P2_U3312) );
  AND2_X1 U10947 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9848), .ZN(P2_U3313) );
  AND2_X1 U10948 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9848), .ZN(P2_U3314) );
  AND2_X1 U10949 ( .A1(n9848), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3315) );
  AND2_X1 U10950 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9848), .ZN(P2_U3316) );
  AND2_X1 U10951 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9848), .ZN(P2_U3317) );
  AND2_X1 U10952 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9848), .ZN(P2_U3318) );
  AND2_X1 U10953 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9848), .ZN(P2_U3319) );
  INV_X1 U10954 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n10142) );
  NOR2_X1 U10955 ( .A1(n9845), .A2(n10142), .ZN(P2_U3320) );
  AND2_X1 U10956 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9848), .ZN(P2_U3321) );
  INV_X1 U10957 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n10244) );
  NOR2_X1 U10958 ( .A1(n9845), .A2(n10244), .ZN(P2_U3322) );
  AND2_X1 U10959 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9848), .ZN(P2_U3323) );
  AND2_X1 U10960 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9848), .ZN(P2_U3324) );
  AND2_X1 U10961 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9848), .ZN(P2_U3325) );
  AND2_X1 U10962 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9848), .ZN(P2_U3326) );
  AOI22_X1 U10963 ( .A1(n9850), .A2(n9847), .B1(n9846), .B2(n9848), .ZN(
        P2_U3437) );
  AOI22_X1 U10964 ( .A1(n9850), .A2(n9849), .B1(n10076), .B2(n9848), .ZN(
        P2_U3438) );
  AOI21_X1 U10965 ( .B1(n9852), .B2(n6231), .A(n9851), .ZN(n9853) );
  OAI21_X1 U10966 ( .B1(n9854), .B2(n9864), .A(n9853), .ZN(n9855) );
  AOI21_X1 U10967 ( .B1(n9857), .B2(n9856), .A(n9855), .ZN(n9916) );
  INV_X1 U10968 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10186) );
  AOI22_X1 U10969 ( .A1(n9915), .A2(n9916), .B1(n10186), .B2(n9913), .ZN(
        P2_U3451) );
  OAI211_X1 U10970 ( .C1(n9860), .C2(n9905), .A(n9859), .B(n9858), .ZN(n9861)
         );
  AOI21_X1 U10971 ( .B1(n9912), .B2(n9862), .A(n9861), .ZN(n9917) );
  INV_X1 U10972 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9863) );
  AOI22_X1 U10973 ( .A1(n9915), .A2(n9917), .B1(n9863), .B2(n9913), .ZN(
        P2_U3466) );
  NOR2_X1 U10974 ( .A1(n9865), .A2(n9864), .ZN(n9870) );
  OAI22_X1 U10975 ( .A1(n9867), .A2(n9907), .B1(n9866), .B2(n9905), .ZN(n9869)
         );
  AOI211_X1 U10976 ( .C1(n9870), .C2(n7328), .A(n9869), .B(n9868), .ZN(n9918)
         );
  INV_X1 U10977 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9871) );
  AOI22_X1 U10978 ( .A1(n9915), .A2(n9918), .B1(n9871), .B2(n9913), .ZN(
        P2_U3469) );
  OAI22_X1 U10979 ( .A1(n9873), .A2(n9907), .B1(n9872), .B2(n9905), .ZN(n9875)
         );
  AOI211_X1 U10980 ( .C1(n9912), .C2(n9876), .A(n9875), .B(n9874), .ZN(n9919)
         );
  INV_X1 U10981 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9877) );
  AOI22_X1 U10982 ( .A1(n9915), .A2(n9919), .B1(n9877), .B2(n9913), .ZN(
        P2_U3472) );
  INV_X1 U10983 ( .A(n9878), .ZN(n9896) );
  OAI22_X1 U10984 ( .A1(n9880), .A2(n9907), .B1(n9879), .B2(n9905), .ZN(n9882)
         );
  AOI211_X1 U10985 ( .C1(n9896), .C2(n9883), .A(n9882), .B(n9881), .ZN(n9920)
         );
  INV_X1 U10986 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9884) );
  AOI22_X1 U10987 ( .A1(n9915), .A2(n9920), .B1(n9884), .B2(n9913), .ZN(
        P2_U3475) );
  OAI22_X1 U10988 ( .A1(n9885), .A2(n9907), .B1(n7385), .B2(n9905), .ZN(n9887)
         );
  AOI211_X1 U10989 ( .C1(n9896), .C2(n9888), .A(n9887), .B(n9886), .ZN(n9921)
         );
  INV_X1 U10990 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9889) );
  AOI22_X1 U10991 ( .A1(n9915), .A2(n9921), .B1(n9889), .B2(n9913), .ZN(
        P2_U3478) );
  INV_X1 U10992 ( .A(n9890), .ZN(n9895) );
  OAI22_X1 U10993 ( .A1(n9892), .A2(n9907), .B1(n9891), .B2(n9905), .ZN(n9894)
         );
  AOI211_X1 U10994 ( .C1(n9896), .C2(n9895), .A(n9894), .B(n9893), .ZN(n9922)
         );
  INV_X1 U10995 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9897) );
  AOI22_X1 U10996 ( .A1(n9915), .A2(n9922), .B1(n9897), .B2(n9913), .ZN(
        P2_U3481) );
  INV_X1 U10997 ( .A(n9898), .ZN(n9903) );
  OAI22_X1 U10998 ( .A1(n9900), .A2(n9907), .B1(n9899), .B2(n9905), .ZN(n9902)
         );
  AOI211_X1 U10999 ( .C1(n9903), .C2(n9912), .A(n9902), .B(n9901), .ZN(n9923)
         );
  INV_X1 U11000 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10130) );
  AOI22_X1 U11001 ( .A1(n9915), .A2(n9923), .B1(n10130), .B2(n9913), .ZN(
        P2_U3484) );
  INV_X1 U11002 ( .A(n9904), .ZN(n9911) );
  OAI22_X1 U11003 ( .A1(n9908), .A2(n9907), .B1(n9906), .B2(n9905), .ZN(n9910)
         );
  AOI211_X1 U11004 ( .C1(n9912), .C2(n9911), .A(n9910), .B(n9909), .ZN(n9926)
         );
  INV_X1 U11005 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9914) );
  AOI22_X1 U11006 ( .A1(n9915), .A2(n9926), .B1(n9914), .B2(n9913), .ZN(
        P2_U3487) );
  AOI22_X1 U11007 ( .A1(n9927), .A2(n9916), .B1(n10272), .B2(n9924), .ZN(
        P2_U3520) );
  AOI22_X1 U11008 ( .A1(n9927), .A2(n9917), .B1(n6954), .B2(n9924), .ZN(
        P2_U3525) );
  AOI22_X1 U11009 ( .A1(n9927), .A2(n9918), .B1(n6953), .B2(n9924), .ZN(
        P2_U3526) );
  AOI22_X1 U11010 ( .A1(n9927), .A2(n9919), .B1(n6952), .B2(n9924), .ZN(
        P2_U3527) );
  AOI22_X1 U11011 ( .A1(n9927), .A2(n9920), .B1(n6951), .B2(n9924), .ZN(
        P2_U3528) );
  AOI22_X1 U11012 ( .A1(n9927), .A2(n9921), .B1(n6950), .B2(n9924), .ZN(
        P2_U3529) );
  AOI22_X1 U11013 ( .A1(n9927), .A2(n9922), .B1(n6949), .B2(n9924), .ZN(
        P2_U3530) );
  AOI22_X1 U11014 ( .A1(n9927), .A2(n9923), .B1(n6967), .B2(n9924), .ZN(
        P2_U3531) );
  AOI22_X1 U11015 ( .A1(n9927), .A2(n9926), .B1(n9925), .B2(n9924), .ZN(
        P2_U3532) );
  INV_X1 U11016 ( .A(n9928), .ZN(n9929) );
  NAND2_X1 U11017 ( .A1(n9930), .A2(n9929), .ZN(n9931) );
  XOR2_X1 U11018 ( .A(n9932), .B(n9931), .Z(ADD_1071_U5) );
  INV_X1 U11019 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n9933) );
  AOI22_X1 U11020 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .B1(n9933), .B2(n10143), .ZN(ADD_1071_U46) );
  OAI21_X1 U11021 ( .B1(n9936), .B2(n9935), .A(n9934), .ZN(ADD_1071_U56) );
  OAI21_X1 U11022 ( .B1(n9939), .B2(n9938), .A(n9937), .ZN(ADD_1071_U57) );
  OAI21_X1 U11023 ( .B1(n9942), .B2(n9941), .A(n9940), .ZN(ADD_1071_U58) );
  OAI21_X1 U11024 ( .B1(n9945), .B2(n9944), .A(n9943), .ZN(ADD_1071_U59) );
  OAI21_X1 U11025 ( .B1(n9948), .B2(n9947), .A(n9946), .ZN(ADD_1071_U60) );
  OAI21_X1 U11026 ( .B1(n9951), .B2(n9950), .A(n9949), .ZN(ADD_1071_U61) );
  AOI21_X1 U11027 ( .B1(n9954), .B2(n9953), .A(n9952), .ZN(ADD_1071_U62) );
  AOI21_X1 U11028 ( .B1(n9957), .B2(n9956), .A(n9955), .ZN(ADD_1071_U63) );
  OAI22_X1 U11029 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(keyinput42), .B1(
        keyinput66), .B2(P2_REG0_REG_24__SCAN_IN), .ZN(n9958) );
  AOI221_X1 U11030 ( .B1(P1_REG3_REG_13__SCAN_IN), .B2(keyinput42), .C1(
        P2_REG0_REG_24__SCAN_IN), .C2(keyinput66), .A(n9958), .ZN(n9965) );
  OAI22_X1 U11031 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(keyinput68), .B1(
        keyinput85), .B2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9959) );
  AOI221_X1 U11032 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(keyinput68), .C1(
        P2_ADDR_REG_6__SCAN_IN), .C2(keyinput85), .A(n9959), .ZN(n9964) );
  OAI22_X1 U11033 ( .A1(P1_REG0_REG_16__SCAN_IN), .A2(keyinput0), .B1(
        P2_REG1_REG_20__SCAN_IN), .B2(keyinput112), .ZN(n9960) );
  AOI221_X1 U11034 ( .B1(P1_REG0_REG_16__SCAN_IN), .B2(keyinput0), .C1(
        keyinput112), .C2(P2_REG1_REG_20__SCAN_IN), .A(n9960), .ZN(n9963) );
  OAI22_X1 U11035 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(keyinput111), .B1(
        P1_REG2_REG_17__SCAN_IN), .B2(keyinput106), .ZN(n9961) );
  AOI221_X1 U11036 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(keyinput111), .C1(
        keyinput106), .C2(P1_REG2_REG_17__SCAN_IN), .A(n9961), .ZN(n9962) );
  NAND4_X1 U11037 ( .A1(n9965), .A2(n9964), .A3(n9963), .A4(n9962), .ZN(n9993)
         );
  OAI22_X1 U11038 ( .A1(P1_REG2_REG_19__SCAN_IN), .A2(keyinput49), .B1(
        P2_D_REG_1__SCAN_IN), .B2(keyinput2), .ZN(n9966) );
  AOI221_X1 U11039 ( .B1(P1_REG2_REG_19__SCAN_IN), .B2(keyinput49), .C1(
        keyinput2), .C2(P2_D_REG_1__SCAN_IN), .A(n9966), .ZN(n9973) );
  OAI22_X1 U11040 ( .A1(P1_REG0_REG_21__SCAN_IN), .A2(keyinput121), .B1(
        P2_WR_REG_SCAN_IN), .B2(keyinput36), .ZN(n9967) );
  AOI221_X1 U11041 ( .B1(P1_REG0_REG_21__SCAN_IN), .B2(keyinput121), .C1(
        keyinput36), .C2(P2_WR_REG_SCAN_IN), .A(n9967), .ZN(n9972) );
  OAI22_X1 U11042 ( .A1(SI_20_), .A2(keyinput87), .B1(P2_REG1_REG_8__SCAN_IN), 
        .B2(keyinput13), .ZN(n9968) );
  AOI221_X1 U11043 ( .B1(SI_20_), .B2(keyinput87), .C1(keyinput13), .C2(
        P2_REG1_REG_8__SCAN_IN), .A(n9968), .ZN(n9971) );
  OAI22_X1 U11044 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(keyinput46), .B1(
        keyinput40), .B2(P2_REG3_REG_12__SCAN_IN), .ZN(n9969) );
  AOI221_X1 U11045 ( .B1(P2_IR_REG_10__SCAN_IN), .B2(keyinput46), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput40), .A(n9969), .ZN(n9970) );
  NAND4_X1 U11046 ( .A1(n9973), .A2(n9972), .A3(n9971), .A4(n9970), .ZN(n9992)
         );
  OAI22_X1 U11047 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(keyinput94), .B1(
        keyinput71), .B2(P2_ADDR_REG_0__SCAN_IN), .ZN(n9974) );
  AOI221_X1 U11048 ( .B1(P2_IR_REG_25__SCAN_IN), .B2(keyinput94), .C1(
        P2_ADDR_REG_0__SCAN_IN), .C2(keyinput71), .A(n9974), .ZN(n9981) );
  OAI22_X1 U11049 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(keyinput95), .B1(
        keyinput58), .B2(P1_REG0_REG_9__SCAN_IN), .ZN(n9975) );
  AOI221_X1 U11050 ( .B1(P2_DATAO_REG_0__SCAN_IN), .B2(keyinput95), .C1(
        P1_REG0_REG_9__SCAN_IN), .C2(keyinput58), .A(n9975), .ZN(n9980) );
  OAI22_X1 U11051 ( .A1(P1_REG0_REG_22__SCAN_IN), .A2(keyinput48), .B1(
        keyinput113), .B2(P2_REG0_REG_7__SCAN_IN), .ZN(n9976) );
  AOI221_X1 U11052 ( .B1(P1_REG0_REG_22__SCAN_IN), .B2(keyinput48), .C1(
        P2_REG0_REG_7__SCAN_IN), .C2(keyinput113), .A(n9976), .ZN(n9979) );
  OAI22_X1 U11053 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(keyinput77), .B1(
        keyinput25), .B2(SI_6_), .ZN(n9977) );
  AOI221_X1 U11054 ( .B1(P1_DATAO_REG_25__SCAN_IN), .B2(keyinput77), .C1(SI_6_), .C2(keyinput25), .A(n9977), .ZN(n9978) );
  NAND4_X1 U11055 ( .A1(n9981), .A2(n9980), .A3(n9979), .A4(n9978), .ZN(n9991)
         );
  OAI22_X1 U11056 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(keyinput119), .B1(
        keyinput107), .B2(P1_REG2_REG_2__SCAN_IN), .ZN(n9982) );
  AOI221_X1 U11057 ( .B1(P1_DATAO_REG_14__SCAN_IN), .B2(keyinput119), .C1(
        P1_REG2_REG_2__SCAN_IN), .C2(keyinput107), .A(n9982), .ZN(n9989) );
  OAI22_X1 U11058 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(keyinput110), .B1(
        keyinput117), .B2(SI_30_), .ZN(n9983) );
  AOI221_X1 U11059 ( .B1(P1_DATAO_REG_24__SCAN_IN), .B2(keyinput110), .C1(
        SI_30_), .C2(keyinput117), .A(n9983), .ZN(n9988) );
  OAI22_X1 U11060 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(keyinput34), .B1(
        P2_REG0_REG_11__SCAN_IN), .B2(keyinput78), .ZN(n9984) );
  AOI221_X1 U11061 ( .B1(P1_IR_REG_30__SCAN_IN), .B2(keyinput34), .C1(
        keyinput78), .C2(P2_REG0_REG_11__SCAN_IN), .A(n9984), .ZN(n9987) );
  OAI22_X1 U11062 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(keyinput23), .B1(
        keyinput76), .B2(P2_REG1_REG_31__SCAN_IN), .ZN(n9985) );
  AOI221_X1 U11063 ( .B1(P1_DATAO_REG_0__SCAN_IN), .B2(keyinput23), .C1(
        P2_REG1_REG_31__SCAN_IN), .C2(keyinput76), .A(n9985), .ZN(n9986) );
  NAND4_X1 U11064 ( .A1(n9989), .A2(n9988), .A3(n9987), .A4(n9986), .ZN(n9990)
         );
  NOR4_X1 U11065 ( .A1(n9993), .A2(n9992), .A3(n9991), .A4(n9990), .ZN(n10325)
         );
  AOI22_X1 U11066 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(keyinput200), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput210), .ZN(n9994) );
  OAI221_X1 U11067 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(keyinput200), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput210), .A(n9994), .ZN(n10001) );
  AOI22_X1 U11068 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(keyinput254), .B1(
        P2_D_REG_25__SCAN_IN), .B2(keyinput202), .ZN(n9995) );
  OAI221_X1 U11069 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(keyinput254), .C1(
        P2_D_REG_25__SCAN_IN), .C2(keyinput202), .A(n9995), .ZN(n10000) );
  AOI22_X1 U11070 ( .A1(P2_D_REG_13__SCAN_IN), .A2(keyinput146), .B1(
        P1_REG0_REG_0__SCAN_IN), .B2(keyinput230), .ZN(n9996) );
  OAI221_X1 U11071 ( .B1(P2_D_REG_13__SCAN_IN), .B2(keyinput146), .C1(
        P1_REG0_REG_0__SCAN_IN), .C2(keyinput230), .A(n9996), .ZN(n9999) );
  AOI22_X1 U11072 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(keyinput150), .B1(
        P1_IR_REG_3__SCAN_IN), .B2(keyinput216), .ZN(n9997) );
  OAI221_X1 U11073 ( .B1(P1_DATAO_REG_30__SCAN_IN), .B2(keyinput150), .C1(
        P1_IR_REG_3__SCAN_IN), .C2(keyinput216), .A(n9997), .ZN(n9998) );
  NOR4_X1 U11074 ( .A1(n10001), .A2(n10000), .A3(n9999), .A4(n9998), .ZN(
        n10029) );
  AOI22_X1 U11075 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(keyinput228), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(keyinput149), .ZN(n10002) );
  OAI221_X1 U11076 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(keyinput228), .C1(
        P2_DATAO_REG_24__SCAN_IN), .C2(keyinput149), .A(n10002), .ZN(n10009)
         );
  AOI22_X1 U11077 ( .A1(P1_D_REG_10__SCAN_IN), .A2(keyinput135), .B1(
        P1_IR_REG_0__SCAN_IN), .B2(keyinput239), .ZN(n10003) );
  OAI221_X1 U11078 ( .B1(P1_D_REG_10__SCAN_IN), .B2(keyinput135), .C1(
        P1_IR_REG_0__SCAN_IN), .C2(keyinput239), .A(n10003), .ZN(n10008) );
  AOI22_X1 U11079 ( .A1(P2_REG0_REG_18__SCAN_IN), .A2(keyinput195), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(keyinput154), .ZN(n10004) );
  OAI221_X1 U11080 ( .B1(P2_REG0_REG_18__SCAN_IN), .B2(keyinput195), .C1(
        P2_DATAO_REG_10__SCAN_IN), .C2(keyinput154), .A(n10004), .ZN(n10007)
         );
  AOI22_X1 U11081 ( .A1(P1_D_REG_3__SCAN_IN), .A2(keyinput193), .B1(
        P1_D_REG_4__SCAN_IN), .B2(keyinput180), .ZN(n10005) );
  OAI221_X1 U11082 ( .B1(P1_D_REG_3__SCAN_IN), .B2(keyinput193), .C1(
        P1_D_REG_4__SCAN_IN), .C2(keyinput180), .A(n10005), .ZN(n10006) );
  NOR4_X1 U11083 ( .A1(n10009), .A2(n10008), .A3(n10007), .A4(n10006), .ZN(
        n10028) );
  AOI22_X1 U11084 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(keyinput141), .B1(
        P2_REG1_REG_26__SCAN_IN), .B2(keyinput157), .ZN(n10010) );
  OAI221_X1 U11085 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(keyinput141), .C1(
        P2_REG1_REG_26__SCAN_IN), .C2(keyinput157), .A(n10010), .ZN(n10017) );
  AOI22_X1 U11086 ( .A1(P2_REG1_REG_31__SCAN_IN), .A2(keyinput204), .B1(
        P1_REG3_REG_13__SCAN_IN), .B2(keyinput170), .ZN(n10011) );
  OAI221_X1 U11087 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(keyinput204), .C1(
        P1_REG3_REG_13__SCAN_IN), .C2(keyinput170), .A(n10011), .ZN(n10016) );
  AOI22_X1 U11088 ( .A1(P2_REG0_REG_24__SCAN_IN), .A2(keyinput194), .B1(
        P1_IR_REG_17__SCAN_IN), .B2(keyinput242), .ZN(n10012) );
  OAI221_X1 U11089 ( .B1(P2_REG0_REG_24__SCAN_IN), .B2(keyinput194), .C1(
        P1_IR_REG_17__SCAN_IN), .C2(keyinput242), .A(n10012), .ZN(n10015) );
  AOI22_X1 U11090 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput248), .B1(
        P2_IR_REG_4__SCAN_IN), .B2(keyinput246), .ZN(n10013) );
  OAI221_X1 U11091 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput248), .C1(
        P2_IR_REG_4__SCAN_IN), .C2(keyinput246), .A(n10013), .ZN(n10014) );
  NOR4_X1 U11092 ( .A1(n10017), .A2(n10016), .A3(n10015), .A4(n10014), .ZN(
        n10027) );
  AOI22_X1 U11093 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(keyinput213), .B1(
        P1_REG1_REG_26__SCAN_IN), .B2(keyinput209), .ZN(n10018) );
  OAI221_X1 U11094 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(keyinput213), .C1(
        P1_REG1_REG_26__SCAN_IN), .C2(keyinput209), .A(n10018), .ZN(n10025) );
  AOI22_X1 U11095 ( .A1(P2_REG0_REG_26__SCAN_IN), .A2(keyinput198), .B1(
        P2_ADDR_REG_19__SCAN_IN), .B2(keyinput237), .ZN(n10019) );
  OAI221_X1 U11096 ( .B1(P2_REG0_REG_26__SCAN_IN), .B2(keyinput198), .C1(
        P2_ADDR_REG_19__SCAN_IN), .C2(keyinput237), .A(n10019), .ZN(n10024) );
  AOI22_X1 U11097 ( .A1(P1_REG0_REG_17__SCAN_IN), .A2(keyinput212), .B1(SI_3_), 
        .B2(keyinput225), .ZN(n10020) );
  OAI221_X1 U11098 ( .B1(P1_REG0_REG_17__SCAN_IN), .B2(keyinput212), .C1(SI_3_), .C2(keyinput225), .A(n10020), .ZN(n10023) );
  AOI22_X1 U11099 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput164), .B1(
        P1_B_REG_SCAN_IN), .B2(keyinput252), .ZN(n10021) );
  OAI221_X1 U11100 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput164), .C1(
        P1_B_REG_SCAN_IN), .C2(keyinput252), .A(n10021), .ZN(n10022) );
  NOR4_X1 U11101 ( .A1(n10025), .A2(n10024), .A3(n10023), .A4(n10022), .ZN(
        n10026) );
  NAND4_X1 U11102 ( .A1(n10029), .A2(n10028), .A3(n10027), .A4(n10026), .ZN(
        n10170) );
  AOI22_X1 U11103 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(keyinput158), .B1(
        P1_REG2_REG_12__SCAN_IN), .B2(keyinput165), .ZN(n10030) );
  OAI221_X1 U11104 ( .B1(P2_IR_REG_13__SCAN_IN), .B2(keyinput158), .C1(
        P1_REG2_REG_12__SCAN_IN), .C2(keyinput165), .A(n10030), .ZN(n10037) );
  AOI22_X1 U11105 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(keyinput201), .B1(
        P1_REG1_REG_22__SCAN_IN), .B2(keyinput152), .ZN(n10031) );
  OAI221_X1 U11106 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(keyinput201), .C1(
        P1_REG1_REG_22__SCAN_IN), .C2(keyinput152), .A(n10031), .ZN(n10036) );
  AOI22_X1 U11107 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(keyinput222), .B1(
        P2_IR_REG_31__SCAN_IN), .B2(keyinput132), .ZN(n10032) );
  OAI221_X1 U11108 ( .B1(P2_IR_REG_25__SCAN_IN), .B2(keyinput222), .C1(
        P2_IR_REG_31__SCAN_IN), .C2(keyinput132), .A(n10032), .ZN(n10035) );
  AOI22_X1 U11109 ( .A1(P2_REG2_REG_1__SCAN_IN), .A2(keyinput188), .B1(
        P1_REG1_REG_9__SCAN_IN), .B2(keyinput172), .ZN(n10033) );
  OAI221_X1 U11110 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(keyinput188), .C1(
        P1_REG1_REG_9__SCAN_IN), .C2(keyinput172), .A(n10033), .ZN(n10034) );
  NOR4_X1 U11111 ( .A1(n10037), .A2(n10036), .A3(n10035), .A4(n10034), .ZN(
        n10065) );
  AOI22_X1 U11112 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(keyinput129), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput136), .ZN(n10038) );
  OAI221_X1 U11113 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(keyinput129), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput136), .A(n10038), .ZN(n10045) );
  AOI22_X1 U11114 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(keyinput224), .B1(
        P1_IR_REG_23__SCAN_IN), .B2(keyinput137), .ZN(n10039) );
  OAI221_X1 U11115 ( .B1(P2_DATAO_REG_30__SCAN_IN), .B2(keyinput224), .C1(
        P1_IR_REG_23__SCAN_IN), .C2(keyinput137), .A(n10039), .ZN(n10044) );
  AOI22_X1 U11116 ( .A1(P2_REG0_REG_2__SCAN_IN), .A2(keyinput187), .B1(
        P1_REG0_REG_25__SCAN_IN), .B2(keyinput133), .ZN(n10040) );
  OAI221_X1 U11117 ( .B1(P2_REG0_REG_2__SCAN_IN), .B2(keyinput187), .C1(
        P1_REG0_REG_25__SCAN_IN), .C2(keyinput133), .A(n10040), .ZN(n10043) );
  AOI22_X1 U11118 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(keyinput156), .B1(
        P1_IR_REG_7__SCAN_IN), .B2(keyinput139), .ZN(n10041) );
  OAI221_X1 U11119 ( .B1(P1_IR_REG_26__SCAN_IN), .B2(keyinput156), .C1(
        P1_IR_REG_7__SCAN_IN), .C2(keyinput139), .A(n10041), .ZN(n10042) );
  NOR4_X1 U11120 ( .A1(n10045), .A2(n10044), .A3(n10043), .A4(n10042), .ZN(
        n10064) );
  AOI22_X1 U11121 ( .A1(P1_REG0_REG_9__SCAN_IN), .A2(keyinput186), .B1(
        P1_IR_REG_31__SCAN_IN), .B2(keyinput163), .ZN(n10046) );
  OAI221_X1 U11122 ( .B1(P1_REG0_REG_9__SCAN_IN), .B2(keyinput186), .C1(
        P1_IR_REG_31__SCAN_IN), .C2(keyinput163), .A(n10046), .ZN(n10053) );
  AOI22_X1 U11123 ( .A1(P1_REG1_REG_31__SCAN_IN), .A2(keyinput171), .B1(
        P1_REG1_REG_24__SCAN_IN), .B2(keyinput203), .ZN(n10047) );
  OAI221_X1 U11124 ( .B1(P1_REG1_REG_31__SCAN_IN), .B2(keyinput171), .C1(
        P1_REG1_REG_24__SCAN_IN), .C2(keyinput203), .A(n10047), .ZN(n10052) );
  AOI22_X1 U11125 ( .A1(P2_REG0_REG_7__SCAN_IN), .A2(keyinput241), .B1(
        P2_IR_REG_12__SCAN_IN), .B2(keyinput143), .ZN(n10048) );
  OAI221_X1 U11126 ( .B1(P2_REG0_REG_7__SCAN_IN), .B2(keyinput241), .C1(
        P2_IR_REG_12__SCAN_IN), .C2(keyinput143), .A(n10048), .ZN(n10051) );
  AOI22_X1 U11127 ( .A1(P2_REG1_REG_20__SCAN_IN), .A2(keyinput240), .B1(
        P1_RD_REG_SCAN_IN), .B2(keyinput226), .ZN(n10049) );
  OAI221_X1 U11128 ( .B1(P2_REG1_REG_20__SCAN_IN), .B2(keyinput240), .C1(
        P1_RD_REG_SCAN_IN), .C2(keyinput226), .A(n10049), .ZN(n10050) );
  NOR4_X1 U11129 ( .A1(n10053), .A2(n10052), .A3(n10051), .A4(n10050), .ZN(
        n10063) );
  AOI22_X1 U11130 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput147), .B1(
        P1_REG3_REG_15__SCAN_IN), .B2(keyinput140), .ZN(n10054) );
  OAI221_X1 U11131 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput147), .C1(
        P1_REG3_REG_15__SCAN_IN), .C2(keyinput140), .A(n10054), .ZN(n10061) );
  AOI22_X1 U11132 ( .A1(P2_D_REG_6__SCAN_IN), .A2(keyinput255), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(keyinput151), .ZN(n10055) );
  OAI221_X1 U11133 ( .B1(P2_D_REG_6__SCAN_IN), .B2(keyinput255), .C1(
        P1_DATAO_REG_0__SCAN_IN), .C2(keyinput151), .A(n10055), .ZN(n10060) );
  AOI22_X1 U11134 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(keyinput182), .B1(
        P1_REG2_REG_1__SCAN_IN), .B2(keyinput192), .ZN(n10056) );
  OAI221_X1 U11135 ( .B1(P2_IR_REG_2__SCAN_IN), .B2(keyinput182), .C1(
        P1_REG2_REG_1__SCAN_IN), .C2(keyinput192), .A(n10056), .ZN(n10059) );
  AOI22_X1 U11136 ( .A1(P2_RD_REG_SCAN_IN), .A2(keyinput161), .B1(
        P1_D_REG_9__SCAN_IN), .B2(keyinput251), .ZN(n10057) );
  OAI221_X1 U11137 ( .B1(P2_RD_REG_SCAN_IN), .B2(keyinput161), .C1(
        P1_D_REG_9__SCAN_IN), .C2(keyinput251), .A(n10057), .ZN(n10058) );
  NOR4_X1 U11138 ( .A1(n10061), .A2(n10060), .A3(n10059), .A4(n10058), .ZN(
        n10062) );
  NAND4_X1 U11139 ( .A1(n10065), .A2(n10064), .A3(n10063), .A4(n10062), .ZN(
        n10169) );
  AOI22_X1 U11140 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput173), .B1(SI_20_), 
        .B2(keyinput215), .ZN(n10066) );
  OAI221_X1 U11141 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput173), .C1(SI_20_), .C2(keyinput215), .A(n10066), .ZN(n10073) );
  AOI22_X1 U11142 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(keyinput190), .B1(
        P1_REG2_REG_2__SCAN_IN), .B2(keyinput235), .ZN(n10067) );
  OAI221_X1 U11143 ( .B1(P2_IR_REG_18__SCAN_IN), .B2(keyinput190), .C1(
        P1_REG2_REG_2__SCAN_IN), .C2(keyinput235), .A(n10067), .ZN(n10072) );
  AOI22_X1 U11144 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput134), .B1(
        P1_D_REG_5__SCAN_IN), .B2(keyinput221), .ZN(n10068) );
  OAI221_X1 U11145 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput134), .C1(
        P1_D_REG_5__SCAN_IN), .C2(keyinput221), .A(n10068), .ZN(n10071) );
  AOI22_X1 U11146 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(keyinput199), .B1(n6288), 
        .B2(keyinput131), .ZN(n10069) );
  OAI221_X1 U11147 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(keyinput199), .C1(n6288), 
        .C2(keyinput131), .A(n10069), .ZN(n10070) );
  NOR4_X1 U11148 ( .A1(n10073), .A2(n10072), .A3(n10071), .A4(n10070), .ZN(
        n10114) );
  AOI22_X1 U11149 ( .A1(n10075), .A2(keyinput253), .B1(n10246), .B2(
        keyinput227), .ZN(n10074) );
  OAI221_X1 U11150 ( .B1(n10075), .B2(keyinput253), .C1(n10246), .C2(
        keyinput227), .A(n10074), .ZN(n10080) );
  XNOR2_X1 U11151 ( .A(n10076), .B(keyinput130), .ZN(n10079) );
  XNOR2_X1 U11152 ( .A(n10077), .B(keyinput208), .ZN(n10078) );
  OR3_X1 U11153 ( .A1(n10080), .A2(n10079), .A3(n10078), .ZN(n10087) );
  AOI22_X1 U11154 ( .A1(n10082), .A2(keyinput159), .B1(keyinput211), .B2(n5398), .ZN(n10081) );
  OAI221_X1 U11155 ( .B1(n10082), .B2(keyinput159), .C1(n5398), .C2(
        keyinput211), .A(n10081), .ZN(n10086) );
  INV_X1 U11156 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10194) );
  AOI22_X1 U11157 ( .A1(n10194), .A2(keyinput244), .B1(n10084), .B2(
        keyinput218), .ZN(n10083) );
  OAI221_X1 U11158 ( .B1(n10194), .B2(keyinput244), .C1(n10084), .C2(
        keyinput218), .A(n10083), .ZN(n10085) );
  NOR3_X1 U11159 ( .A1(n10087), .A2(n10086), .A3(n10085), .ZN(n10113) );
  INV_X1 U11160 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n10089) );
  AOI22_X1 U11161 ( .A1(n10089), .A2(keyinput145), .B1(keyinput207), .B2(n5967), .ZN(n10088) );
  OAI221_X1 U11162 ( .B1(n10089), .B2(keyinput145), .C1(n5967), .C2(
        keyinput207), .A(n10088), .ZN(n10099) );
  AOI22_X1 U11163 ( .A1(n10091), .A2(keyinput233), .B1(keyinput231), .B2(n8213), .ZN(n10090) );
  OAI221_X1 U11164 ( .B1(n10091), .B2(keyinput233), .C1(n8213), .C2(
        keyinput231), .A(n10090), .ZN(n10098) );
  INV_X1 U11165 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10093) );
  AOI22_X1 U11166 ( .A1(n10093), .A2(keyinput234), .B1(keyinput167), .B2(n6278), .ZN(n10092) );
  OAI221_X1 U11167 ( .B1(n10093), .B2(keyinput234), .C1(n6278), .C2(
        keyinput167), .A(n10092), .ZN(n10097) );
  AOI22_X1 U11168 ( .A1(n10095), .A2(keyinput247), .B1(keyinput177), .B2(n5544), .ZN(n10094) );
  OAI221_X1 U11169 ( .B1(n10095), .B2(keyinput247), .C1(n5544), .C2(
        keyinput177), .A(n10094), .ZN(n10096) );
  NOR4_X1 U11170 ( .A1(n10099), .A2(n10098), .A3(n10097), .A4(n10096), .ZN(
        n10112) );
  AOI22_X1 U11171 ( .A1(n10229), .A2(keyinput160), .B1(n10222), .B2(
        keyinput243), .ZN(n10100) );
  OAI221_X1 U11172 ( .B1(n10229), .B2(keyinput160), .C1(n10222), .C2(
        keyinput243), .A(n10100), .ZN(n10110) );
  AOI22_X1 U11173 ( .A1(n10271), .A2(keyinput232), .B1(n10102), .B2(
        keyinput191), .ZN(n10101) );
  OAI221_X1 U11174 ( .B1(n10271), .B2(keyinput232), .C1(n10102), .C2(
        keyinput191), .A(n10101), .ZN(n10109) );
  AOI22_X1 U11175 ( .A1(n10104), .A2(keyinput205), .B1(n10192), .B2(
        keyinput214), .ZN(n10103) );
  OAI221_X1 U11176 ( .B1(n10104), .B2(keyinput205), .C1(n10192), .C2(
        keyinput214), .A(n10103), .ZN(n10108) );
  AOI22_X1 U11177 ( .A1(n10106), .A2(keyinput223), .B1(keyinput220), .B2(n6487), .ZN(n10105) );
  OAI221_X1 U11178 ( .B1(n10106), .B2(keyinput223), .C1(n6487), .C2(
        keyinput220), .A(n10105), .ZN(n10107) );
  NOR4_X1 U11179 ( .A1(n10110), .A2(n10109), .A3(n10108), .A4(n10107), .ZN(
        n10111) );
  NAND4_X1 U11180 ( .A1(n10114), .A2(n10113), .A3(n10112), .A4(n10111), .ZN(
        n10168) );
  AOI22_X1 U11181 ( .A1(n10209), .A2(keyinput178), .B1(n10116), .B2(
        keyinput175), .ZN(n10115) );
  OAI221_X1 U11182 ( .B1(n10209), .B2(keyinput178), .C1(n10116), .C2(
        keyinput175), .A(n10115), .ZN(n10126) );
  AOI22_X1 U11183 ( .A1(n10118), .A2(keyinput181), .B1(keyinput148), .B2(n6949), .ZN(n10117) );
  OAI221_X1 U11184 ( .B1(n10118), .B2(keyinput181), .C1(n6949), .C2(
        keyinput148), .A(n10117), .ZN(n10125) );
  AOI22_X1 U11185 ( .A1(n10185), .A2(keyinput138), .B1(n10120), .B2(
        keyinput238), .ZN(n10119) );
  OAI221_X1 U11186 ( .B1(n10185), .B2(keyinput138), .C1(n10120), .C2(
        keyinput238), .A(n10119), .ZN(n10124) );
  INV_X1 U11187 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n10247) );
  AOI22_X1 U11188 ( .A1(n10122), .A2(keyinput249), .B1(keyinput179), .B2(
        n10247), .ZN(n10121) );
  OAI221_X1 U11189 ( .B1(n10122), .B2(keyinput249), .C1(n10247), .C2(
        keyinput179), .A(n10121), .ZN(n10123) );
  NOR4_X1 U11190 ( .A1(n10126), .A2(n10125), .A3(n10124), .A4(n10123), .ZN(
        n10166) );
  AOI22_X1 U11191 ( .A1(n10204), .A2(keyinput185), .B1(n10128), .B2(
        keyinput144), .ZN(n10127) );
  OAI221_X1 U11192 ( .B1(n10204), .B2(keyinput185), .C1(n10128), .C2(
        keyinput144), .A(n10127), .ZN(n10138) );
  INV_X1 U11193 ( .A(SI_18_), .ZN(n10183) );
  AOI22_X1 U11194 ( .A1(n10183), .A2(keyinput219), .B1(keyinput206), .B2(
        n10130), .ZN(n10129) );
  OAI221_X1 U11195 ( .B1(n10183), .B2(keyinput219), .C1(n10130), .C2(
        keyinput206), .A(n10129), .ZN(n10137) );
  AOI22_X1 U11196 ( .A1(n10182), .A2(keyinput169), .B1(keyinput168), .B2(
        n10132), .ZN(n10131) );
  OAI221_X1 U11197 ( .B1(n10182), .B2(keyinput169), .C1(n10132), .C2(
        keyinput168), .A(n10131), .ZN(n10136) );
  AOI22_X1 U11198 ( .A1(n10134), .A2(keyinput176), .B1(n10226), .B2(
        keyinput189), .ZN(n10133) );
  OAI221_X1 U11199 ( .B1(n10134), .B2(keyinput176), .C1(n10226), .C2(
        keyinput189), .A(n10133), .ZN(n10135) );
  NOR4_X1 U11200 ( .A1(n10138), .A2(n10137), .A3(n10136), .A4(n10135), .ZN(
        n10165) );
  AOI22_X1 U11201 ( .A1(n10266), .A2(keyinput184), .B1(keyinput166), .B2(
        n10186), .ZN(n10139) );
  OAI221_X1 U11202 ( .B1(n10266), .B2(keyinput184), .C1(n10186), .C2(
        keyinput166), .A(n10139), .ZN(n10150) );
  INV_X1 U11203 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10141) );
  AOI22_X1 U11204 ( .A1(n10142), .A2(keyinput183), .B1(n10141), .B2(
        keyinput128), .ZN(n10140) );
  OAI221_X1 U11205 ( .B1(n10142), .B2(keyinput183), .C1(n10141), .C2(
        keyinput128), .A(n10140), .ZN(n10146) );
  XNOR2_X1 U11206 ( .A(n10143), .B(keyinput196), .ZN(n10145) );
  XOR2_X1 U11207 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput162), .Z(n10144) );
  OR3_X1 U11208 ( .A1(n10146), .A2(n10145), .A3(n10144), .ZN(n10149) );
  AOI22_X1 U11209 ( .A1(n7778), .A2(keyinput155), .B1(keyinput217), .B2(n6990), 
        .ZN(n10147) );
  OAI221_X1 U11210 ( .B1(n7778), .B2(keyinput155), .C1(n6990), .C2(keyinput217), .A(n10147), .ZN(n10148) );
  NOR3_X1 U11211 ( .A1(n10150), .A2(n10149), .A3(n10148), .ZN(n10164) );
  INV_X1 U11212 ( .A(SI_30_), .ZN(n10152) );
  AOI22_X1 U11213 ( .A1(n6533), .A2(keyinput236), .B1(keyinput245), .B2(n10152), .ZN(n10151) );
  OAI221_X1 U11214 ( .B1(n6533), .B2(keyinput236), .C1(n10152), .C2(
        keyinput245), .A(n10151), .ZN(n10162) );
  INV_X1 U11215 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n10155) );
  AOI22_X1 U11216 ( .A1(n10155), .A2(keyinput250), .B1(n10154), .B2(
        keyinput153), .ZN(n10153) );
  OAI221_X1 U11217 ( .B1(n10155), .B2(keyinput250), .C1(n10154), .C2(
        keyinput153), .A(n10153), .ZN(n10161) );
  XNOR2_X1 U11218 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput174), .ZN(n10159) );
  XNOR2_X1 U11219 ( .A(P2_REG1_REG_2__SCAN_IN), .B(keyinput229), .ZN(n10158)
         );
  XNOR2_X1 U11220 ( .A(P1_REG1_REG_27__SCAN_IN), .B(keyinput142), .ZN(n10157)
         );
  XNOR2_X1 U11221 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput197), .ZN(n10156) );
  NAND4_X1 U11222 ( .A1(n10159), .A2(n10158), .A3(n10157), .A4(n10156), .ZN(
        n10160) );
  NOR3_X1 U11223 ( .A1(n10162), .A2(n10161), .A3(n10160), .ZN(n10163) );
  NAND4_X1 U11224 ( .A1(n10166), .A2(n10165), .A3(n10164), .A4(n10163), .ZN(
        n10167) );
  NOR4_X1 U11225 ( .A1(n10170), .A2(n10169), .A3(n10168), .A4(n10167), .ZN(
        n10286) );
  AOI22_X1 U11226 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(keyinput72), .B1(
        P1_REG1_REG_22__SCAN_IN), .B2(keyinput24), .ZN(n10171) );
  OAI221_X1 U11227 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(keyinput72), .C1(
        P1_REG1_REG_22__SCAN_IN), .C2(keyinput24), .A(n10171), .ZN(n10178) );
  AOI22_X1 U11228 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(keyinput100), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(keyinput63), .ZN(n10172) );
  OAI221_X1 U11229 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(keyinput100), .C1(
        P2_DATAO_REG_14__SCAN_IN), .C2(keyinput63), .A(n10172), .ZN(n10177) );
  AOI22_X1 U11230 ( .A1(P2_D_REG_25__SCAN_IN), .A2(keyinput74), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(keyinput53), .ZN(n10173) );
  OAI221_X1 U11231 ( .B1(P2_D_REG_25__SCAN_IN), .B2(keyinput74), .C1(
        P1_DATAO_REG_28__SCAN_IN), .C2(keyinput53), .A(n10173), .ZN(n10176) );
  AOI22_X1 U11232 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput45), .B1(
        P2_D_REG_16__SCAN_IN), .B2(keyinput90), .ZN(n10174) );
  OAI221_X1 U11233 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput45), .C1(
        P2_D_REG_16__SCAN_IN), .C2(keyinput90), .A(n10174), .ZN(n10175) );
  NOR4_X1 U11234 ( .A1(n10178), .A2(n10177), .A3(n10176), .A4(n10175), .ZN(
        n10220) );
  AOI22_X1 U11235 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput6), .B1(
        P1_REG3_REG_23__SCAN_IN), .B2(keyinput47), .ZN(n10179) );
  OAI221_X1 U11236 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput6), .C1(
        P1_REG3_REG_23__SCAN_IN), .C2(keyinput47), .A(n10179), .ZN(n10190) );
  AOI22_X1 U11237 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(keyinput1), .B1(
        P1_RD_REG_SCAN_IN), .B2(keyinput98), .ZN(n10180) );
  OAI221_X1 U11238 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(keyinput1), .C1(
        P1_RD_REG_SCAN_IN), .C2(keyinput98), .A(n10180), .ZN(n10189) );
  AOI22_X1 U11239 ( .A1(n10183), .A2(keyinput91), .B1(n10182), .B2(keyinput41), 
        .ZN(n10181) );
  OAI221_X1 U11240 ( .B1(n10183), .B2(keyinput91), .C1(n10182), .C2(keyinput41), .A(n10181), .ZN(n10188) );
  AOI22_X1 U11241 ( .A1(n10186), .A2(keyinput38), .B1(n10185), .B2(keyinput10), 
        .ZN(n10184) );
  OAI221_X1 U11242 ( .B1(n10186), .B2(keyinput38), .C1(n10185), .C2(keyinput10), .A(n10184), .ZN(n10187) );
  NOR4_X1 U11243 ( .A1(n10190), .A2(n10189), .A3(n10188), .A4(n10187), .ZN(
        n10219) );
  AOI22_X1 U11244 ( .A1(n10193), .A2(keyinput97), .B1(n10192), .B2(keyinput86), 
        .ZN(n10191) );
  OAI221_X1 U11245 ( .B1(n10193), .B2(keyinput97), .C1(n10192), .C2(keyinput86), .A(n10191), .ZN(n10202) );
  XOR2_X1 U11246 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput88), .Z(n10201) );
  XNOR2_X1 U11247 ( .A(keyinput116), .B(n10194), .ZN(n10200) );
  XNOR2_X1 U11248 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput118), .ZN(n10198) );
  XNOR2_X1 U11249 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput11), .ZN(n10197) );
  XNOR2_X1 U11250 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput8), .ZN(n10196) );
  XNOR2_X1 U11251 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput9), .ZN(n10195) );
  NAND4_X1 U11252 ( .A1(n10198), .A2(n10197), .A3(n10196), .A4(n10195), .ZN(
        n10199) );
  NOR4_X1 U11253 ( .A1(n10202), .A2(n10201), .A3(n10200), .A4(n10199), .ZN(
        n10218) );
  AOI22_X1 U11254 ( .A1(n10204), .A2(keyinput57), .B1(n6533), .B2(keyinput108), 
        .ZN(n10203) );
  OAI221_X1 U11255 ( .B1(n10204), .B2(keyinput57), .C1(n6533), .C2(keyinput108), .A(n10203), .ZN(n10216) );
  AOI22_X1 U11256 ( .A1(n10207), .A2(keyinput44), .B1(keyinput30), .B2(n10206), 
        .ZN(n10205) );
  OAI221_X1 U11257 ( .B1(n10207), .B2(keyinput44), .C1(n10206), .C2(keyinput30), .A(n10205), .ZN(n10215) );
  AOI22_X1 U11258 ( .A1(n10210), .A2(keyinput60), .B1(n10209), .B2(keyinput50), 
        .ZN(n10208) );
  OAI221_X1 U11259 ( .B1(n10210), .B2(keyinput60), .C1(n10209), .C2(keyinput50), .A(n10208), .ZN(n10214) );
  XNOR2_X1 U11260 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput4), .ZN(n10212) );
  XNOR2_X1 U11261 ( .A(keyinput20), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n10211)
         );
  NAND2_X1 U11262 ( .A1(n10212), .A2(n10211), .ZN(n10213) );
  NOR4_X1 U11263 ( .A1(n10216), .A2(n10215), .A3(n10214), .A4(n10213), .ZN(
        n10217) );
  NAND4_X1 U11264 ( .A1(n10220), .A2(n10219), .A3(n10218), .A4(n10217), .ZN(
        n10285) );
  AOI22_X1 U11265 ( .A1(n10223), .A2(keyinput21), .B1(keyinput115), .B2(n10222), .ZN(n10221) );
  OAI221_X1 U11266 ( .B1(n10223), .B2(keyinput21), .C1(n10222), .C2(
        keyinput115), .A(n10221), .ZN(n10235) );
  INV_X1 U11267 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n10225) );
  AOI22_X1 U11268 ( .A1(n10226), .A2(keyinput61), .B1(keyinput29), .B2(n10225), 
        .ZN(n10224) );
  OAI221_X1 U11269 ( .B1(n10226), .B2(keyinput61), .C1(n10225), .C2(keyinput29), .A(n10224), .ZN(n10234) );
  AOI22_X1 U11270 ( .A1(n10229), .A2(keyinput32), .B1(keyinput14), .B2(n10228), 
        .ZN(n10227) );
  OAI221_X1 U11271 ( .B1(n10229), .B2(keyinput32), .C1(n10228), .C2(keyinput14), .A(n10227), .ZN(n10233) );
  XNOR2_X1 U11272 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput28), .ZN(n10231) );
  XNOR2_X1 U11273 ( .A(keyinput89), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n10230) );
  NAND2_X1 U11274 ( .A1(n10231), .A2(n10230), .ZN(n10232) );
  NOR4_X1 U11275 ( .A1(n10235), .A2(n10234), .A3(n10233), .A4(n10232), .ZN(
        n10283) );
  INV_X1 U11276 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10238) );
  AOI22_X1 U11277 ( .A1(n10238), .A2(keyinput101), .B1(n10237), .B2(keyinput54), .ZN(n10236) );
  OAI221_X1 U11278 ( .B1(n10238), .B2(keyinput101), .C1(n10237), .C2(
        keyinput54), .A(n10236), .ZN(n10251) );
  AOI22_X1 U11279 ( .A1(n10241), .A2(keyinput114), .B1(keyinput19), .B2(n10240), .ZN(n10239) );
  OAI221_X1 U11280 ( .B1(n10241), .B2(keyinput114), .C1(n10240), .C2(
        keyinput19), .A(n10239), .ZN(n10250) );
  INV_X1 U11281 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10243) );
  AOI22_X1 U11282 ( .A1(n10244), .A2(keyinput127), .B1(keyinput120), .B2(
        n10243), .ZN(n10242) );
  OAI221_X1 U11283 ( .B1(n10244), .B2(keyinput127), .C1(n10243), .C2(
        keyinput120), .A(n10242), .ZN(n10249) );
  AOI22_X1 U11284 ( .A1(n10247), .A2(keyinput51), .B1(n10246), .B2(keyinput99), 
        .ZN(n10245) );
  OAI221_X1 U11285 ( .B1(n10247), .B2(keyinput51), .C1(n10246), .C2(keyinput99), .A(n10245), .ZN(n10248) );
  NOR4_X1 U11286 ( .A1(n10251), .A2(n10250), .A3(n10249), .A4(n10248), .ZN(
        n10282) );
  INV_X1 U11287 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n10253) );
  AOI22_X1 U11288 ( .A1(n6278), .A2(keyinput39), .B1(n10253), .B2(keyinput84), 
        .ZN(n10252) );
  OAI221_X1 U11289 ( .B1(n6278), .B2(keyinput39), .C1(n10253), .C2(keyinput84), 
        .A(n10252), .ZN(n10264) );
  INV_X1 U11290 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10256) );
  AOI22_X1 U11291 ( .A1(n10256), .A2(keyinput37), .B1(keyinput126), .B2(n10255), .ZN(n10254) );
  OAI221_X1 U11292 ( .B1(n10256), .B2(keyinput37), .C1(n10255), .C2(
        keyinput126), .A(n10254), .ZN(n10263) );
  INV_X1 U11293 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n10258) );
  AOI22_X1 U11294 ( .A1(n6487), .A2(keyinput92), .B1(n10258), .B2(keyinput70), 
        .ZN(n10257) );
  OAI221_X1 U11295 ( .B1(n6487), .B2(keyinput92), .C1(n10258), .C2(keyinput70), 
        .A(n10257), .ZN(n10262) );
  XNOR2_X1 U11296 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput35), .ZN(n10260) );
  XNOR2_X1 U11297 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput69), .ZN(n10259) );
  NAND2_X1 U11298 ( .A1(n10260), .A2(n10259), .ZN(n10261) );
  NOR4_X1 U11299 ( .A1(n10264), .A2(n10263), .A3(n10262), .A4(n10261), .ZN(
        n10281) );
  AOI22_X1 U11300 ( .A1(n10266), .A2(keyinput56), .B1(keyinput27), .B2(n7778), 
        .ZN(n10265) );
  OAI221_X1 U11301 ( .B1(n10266), .B2(keyinput56), .C1(n7778), .C2(keyinput27), 
        .A(n10265), .ZN(n10279) );
  INV_X1 U11302 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10269) );
  AOI22_X1 U11303 ( .A1(n10269), .A2(keyinput43), .B1(n10268), .B2(keyinput65), 
        .ZN(n10267) );
  OAI221_X1 U11304 ( .B1(n10269), .B2(keyinput43), .C1(n10268), .C2(keyinput65), .A(n10267), .ZN(n10278) );
  AOI22_X1 U11305 ( .A1(n10272), .A2(keyinput73), .B1(keyinput104), .B2(n10271), .ZN(n10270) );
  OAI221_X1 U11306 ( .B1(n10272), .B2(keyinput73), .C1(n10271), .C2(
        keyinput104), .A(n10270), .ZN(n10277) );
  XOR2_X1 U11307 ( .A(n10273), .B(keyinput59), .Z(n10275) );
  XNOR2_X1 U11308 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput33), .ZN(n10274) );
  NAND2_X1 U11309 ( .A1(n10275), .A2(n10274), .ZN(n10276) );
  NOR4_X1 U11310 ( .A1(n10279), .A2(n10278), .A3(n10277), .A4(n10276), .ZN(
        n10280) );
  NAND4_X1 U11311 ( .A1(n10283), .A2(n10282), .A3(n10281), .A4(n10280), .ZN(
        n10284) );
  NOR3_X1 U11312 ( .A1(n10286), .A2(n10285), .A3(n10284), .ZN(n10324) );
  OAI22_X1 U11313 ( .A1(P1_D_REG_10__SCAN_IN), .A2(keyinput7), .B1(
        P2_REG2_REG_0__SCAN_IN), .B2(keyinput125), .ZN(n10287) );
  AOI221_X1 U11314 ( .B1(P1_D_REG_10__SCAN_IN), .B2(keyinput7), .C1(
        keyinput125), .C2(P2_REG2_REG_0__SCAN_IN), .A(n10287), .ZN(n10294) );
  OAI22_X1 U11315 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(keyinput16), .B1(
        P2_D_REG_13__SCAN_IN), .B2(keyinput18), .ZN(n10288) );
  AOI221_X1 U11316 ( .B1(P1_DATAO_REG_22__SCAN_IN), .B2(keyinput16), .C1(
        keyinput18), .C2(P2_D_REG_13__SCAN_IN), .A(n10288), .ZN(n10293) );
  OAI22_X1 U11317 ( .A1(P1_REG2_REG_1__SCAN_IN), .A2(keyinput64), .B1(
        keyinput122), .B2(P2_REG0_REG_29__SCAN_IN), .ZN(n10289) );
  AOI221_X1 U11318 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(keyinput64), .C1(
        P2_REG0_REG_29__SCAN_IN), .C2(keyinput122), .A(n10289), .ZN(n10292) );
  OAI22_X1 U11319 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(keyinput105), .B1(
        P2_IR_REG_18__SCAN_IN), .B2(keyinput62), .ZN(n10290) );
  AOI221_X1 U11320 ( .B1(P1_DATAO_REG_1__SCAN_IN), .B2(keyinput105), .C1(
        keyinput62), .C2(P2_IR_REG_18__SCAN_IN), .A(n10290), .ZN(n10291) );
  NAND4_X1 U11321 ( .A1(n10294), .A2(n10293), .A3(n10292), .A4(n10291), .ZN(
        n10322) );
  OAI22_X1 U11322 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(keyinput109), .B1(
        keyinput82), .B2(P2_REG3_REG_26__SCAN_IN), .ZN(n10295) );
  AOI221_X1 U11323 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(keyinput109), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput82), .A(n10295), .ZN(n10302) );
  OAI22_X1 U11324 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(keyinput80), .B1(
        keyinput96), .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n10296) );
  AOI221_X1 U11325 ( .B1(P2_IR_REG_27__SCAN_IN), .B2(keyinput80), .C1(
        P2_DATAO_REG_30__SCAN_IN), .C2(keyinput96), .A(n10296), .ZN(n10301) );
  OAI22_X1 U11326 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(keyinput26), .B1(
        keyinput15), .B2(P2_IR_REG_12__SCAN_IN), .ZN(n10297) );
  AOI221_X1 U11327 ( .B1(P2_DATAO_REG_10__SCAN_IN), .B2(keyinput26), .C1(
        P2_IR_REG_12__SCAN_IN), .C2(keyinput15), .A(n10297), .ZN(n10300) );
  OAI22_X1 U11328 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(keyinput12), .B1(
        P1_REG1_REG_26__SCAN_IN), .B2(keyinput81), .ZN(n10298) );
  AOI221_X1 U11329 ( .B1(P1_REG3_REG_15__SCAN_IN), .B2(keyinput12), .C1(
        keyinput81), .C2(P1_REG1_REG_26__SCAN_IN), .A(n10298), .ZN(n10299) );
  NAND4_X1 U11330 ( .A1(n10302), .A2(n10301), .A3(n10300), .A4(n10299), .ZN(
        n10321) );
  OAI22_X1 U11331 ( .A1(P1_REG1_REG_6__SCAN_IN), .A2(keyinput3), .B1(
        keyinput22), .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n10303) );
  AOI221_X1 U11332 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(keyinput3), .C1(
        P1_DATAO_REG_30__SCAN_IN), .C2(keyinput22), .A(n10303), .ZN(n10310) );
  OAI22_X1 U11333 ( .A1(P1_REG1_REG_24__SCAN_IN), .A2(keyinput75), .B1(
        P2_D_REG_8__SCAN_IN), .B2(keyinput55), .ZN(n10304) );
  AOI221_X1 U11334 ( .B1(P1_REG1_REG_24__SCAN_IN), .B2(keyinput75), .C1(
        keyinput55), .C2(P2_D_REG_8__SCAN_IN), .A(n10304), .ZN(n10309) );
  OAI22_X1 U11335 ( .A1(P1_D_REG_9__SCAN_IN), .A2(keyinput123), .B1(
        keyinput103), .B2(P2_ADDR_REG_16__SCAN_IN), .ZN(n10305) );
  AOI221_X1 U11336 ( .B1(P1_D_REG_9__SCAN_IN), .B2(keyinput123), .C1(
        P2_ADDR_REG_16__SCAN_IN), .C2(keyinput103), .A(n10305), .ZN(n10308) );
  OAI22_X1 U11337 ( .A1(P1_D_REG_4__SCAN_IN), .A2(keyinput52), .B1(keyinput79), 
        .B2(P2_REG3_REG_13__SCAN_IN), .ZN(n10306) );
  AOI221_X1 U11338 ( .B1(P1_D_REG_4__SCAN_IN), .B2(keyinput52), .C1(
        P2_REG3_REG_13__SCAN_IN), .C2(keyinput79), .A(n10306), .ZN(n10307) );
  NAND4_X1 U11339 ( .A1(n10310), .A2(n10309), .A3(n10308), .A4(n10307), .ZN(
        n10320) );
  OAI22_X1 U11340 ( .A1(P1_REG2_REG_20__SCAN_IN), .A2(keyinput17), .B1(
        P1_REG0_REG_1__SCAN_IN), .B2(keyinput83), .ZN(n10311) );
  AOI221_X1 U11341 ( .B1(P1_REG2_REG_20__SCAN_IN), .B2(keyinput17), .C1(
        keyinput83), .C2(P1_REG0_REG_1__SCAN_IN), .A(n10311), .ZN(n10318) );
  OAI22_X1 U11342 ( .A1(P1_B_REG_SCAN_IN), .A2(keyinput124), .B1(
        P1_REG0_REG_0__SCAN_IN), .B2(keyinput102), .ZN(n10312) );
  AOI221_X1 U11343 ( .B1(P1_B_REG_SCAN_IN), .B2(keyinput124), .C1(keyinput102), 
        .C2(P1_REG0_REG_0__SCAN_IN), .A(n10312), .ZN(n10317) );
  OAI22_X1 U11344 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(keyinput31), .B1(
        keyinput67), .B2(P2_REG0_REG_18__SCAN_IN), .ZN(n10313) );
  AOI221_X1 U11345 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(keyinput31), .C1(
        P2_REG0_REG_18__SCAN_IN), .C2(keyinput67), .A(n10313), .ZN(n10316) );
  OAI22_X1 U11346 ( .A1(P1_D_REG_5__SCAN_IN), .A2(keyinput93), .B1(
        P1_REG0_REG_25__SCAN_IN), .B2(keyinput5), .ZN(n10314) );
  AOI221_X1 U11347 ( .B1(P1_D_REG_5__SCAN_IN), .B2(keyinput93), .C1(keyinput5), 
        .C2(P1_REG0_REG_25__SCAN_IN), .A(n10314), .ZN(n10315) );
  NAND4_X1 U11348 ( .A1(n10318), .A2(n10317), .A3(n10316), .A4(n10315), .ZN(
        n10319) );
  NOR4_X1 U11349 ( .A1(n10322), .A2(n10321), .A3(n10320), .A4(n10319), .ZN(
        n10323) );
  NAND3_X1 U11350 ( .A1(n10325), .A2(n10324), .A3(n10323), .ZN(n10328) );
  MUX2_X1 U11351 ( .A(n10326), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9100), .Z(
        n10327) );
  XNOR2_X1 U11352 ( .A(n10328), .B(n10327), .ZN(P1_U3573) );
  XOR2_X1 U11353 ( .A(n10329), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  XOR2_X1 U11354 ( .A(n10331), .B(n10330), .Z(ADD_1071_U54) );
  NOR2_X1 U11355 ( .A1(n10333), .A2(n10332), .ZN(n10334) );
  XOR2_X1 U11356 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10334), .Z(ADD_1071_U51) );
  OAI21_X1 U11357 ( .B1(n10337), .B2(n10336), .A(n10335), .ZN(n10339) );
  XOR2_X1 U11358 ( .A(n10339), .B(n10338), .Z(ADD_1071_U55) );
  AOI21_X1 U11359 ( .B1(n10342), .B2(n10341), .A(n10340), .ZN(ADD_1071_U47) );
  XOR2_X1 U11360 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10343), .Z(ADD_1071_U48) );
  XOR2_X1 U11361 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10344), .Z(ADD_1071_U49) );
  XOR2_X1 U11362 ( .A(n10346), .B(n10345), .Z(ADD_1071_U53) );
  XNOR2_X1 U11363 ( .A(n10348), .B(n10347), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4978 ( .A(n5905), .Z(n7752) );
endmodule

