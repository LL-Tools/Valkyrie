

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212;

  NOR2_X2 U4888 ( .A1(n7417), .A2(n7769), .ZN(n7732) );
  NAND2_X1 U4889 ( .A1(n6161), .A2(n6238), .ZN(n9771) );
  NAND2_X1 U4890 ( .A1(n5632), .A2(n6243), .ZN(n6978) );
  INV_X1 U4891 ( .A(n9688), .ZN(n7186) );
  INV_X4 U4892 ( .A(n6056), .ZN(n5789) );
  INV_X1 U4894 ( .A(n9350), .ZN(n4486) );
  CLKBUF_X2 U4895 ( .A(n5964), .Z(n4387) );
  CLKBUF_X3 U4896 ( .A(n5197), .Z(n5602) );
  INV_X1 U4897 ( .A(n4980), .ZN(n4749) );
  INV_X1 U4898 ( .A(n5349), .ZN(n6191) );
  INV_X2 U4900 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8011) );
  NAND2_X1 U4901 ( .A1(n6773), .A2(n6692), .ZN(n6851) );
  INV_X1 U4902 ( .A(n6058), .ZN(n6041) );
  INV_X1 U4903 ( .A(n5221), .ZN(n6188) );
  OAI22_X1 U4904 ( .A1(n8796), .A2(n4773), .B1(n4774), .B2(n8437), .ZN(n8768)
         );
  OAI211_X1 U4905 ( .C1(n6562), .C2(n6473), .A(n5223), .B(n5222), .ZN(n7102)
         );
  NOR2_X1 U4906 ( .A1(n9380), .A2(n9202), .ZN(n9193) );
  AOI21_X1 U4907 ( .B1(n9216), .B2(n9635), .A(n9215), .ZN(n9386) );
  AND4_X1 U4908 ( .A1(n5050), .A2(n5049), .A3(n5048), .A4(n5047), .ZN(n4383)
         );
  XOR2_X1 U4909 ( .A(n6064), .B(n6063), .Z(n4384) );
  OR2_X2 U4910 ( .A1(n6112), .A2(n8253), .ZN(n4443) );
  OAI211_X2 U4911 ( .C1(n4781), .C2(n5194), .A(n5219), .B(n4779), .ZN(n5236)
         );
  XNOR2_X2 U4912 ( .A(n4970), .B(n4969), .ZN(n5194) );
  AOI21_X2 U4913 ( .B1(n9771), .B2(n9781), .A(n6266), .ZN(n7328) );
  AND2_X2 U4914 ( .A1(n9510), .A2(n4725), .ZN(n4724) );
  NAND2_X4 U4915 ( .A1(n5684), .A2(n7677), .ZN(n6562) );
  OR2_X2 U4916 ( .A1(n7312), .A2(n6147), .ZN(n6691) );
  NOR2_X2 U4918 ( .A1(n9293), .A2(n9408), .ZN(n9279) );
  NAND2_X2 U4919 ( .A1(n5510), .A2(n5509), .ZN(n8932) );
  OR2_X1 U4920 ( .A1(n9249), .A2(n4801), .ZN(n4798) );
  NAND2_X1 U4921 ( .A1(n4560), .A2(n4852), .ZN(n5511) );
  INV_X2 U4922 ( .A(n8870), .ZN(n4388) );
  INV_X2 U4923 ( .A(n9665), .ZN(n4389) );
  NAND2_X2 U4924 ( .A1(n6244), .A2(n6252), .ZN(n7094) );
  INV_X4 U4925 ( .A(n6738), .ZN(n8062) );
  INV_X1 U4926 ( .A(n7166), .ZN(n9683) );
  NOR2_X1 U4927 ( .A1(n6646), .A2(n6645), .ZN(n6644) );
  INV_X2 U4929 ( .A(n5784), .ZN(n5790) );
  NAND2_X2 U4930 ( .A1(n8412), .A2(n6068), .ZN(n5778) );
  XNOR2_X1 U4931 ( .A(n5746), .B(n5745), .ZN(n8412) );
  OAI21_X1 U4932 ( .B1(n5744), .B2(n4951), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4747) );
  AND2_X1 U4933 ( .A1(n5727), .A2(n4415), .ZN(n6073) );
  NOR2_X1 U4934 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n7652) );
  BUF_X2 U4935 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n9765) );
  INV_X2 U4936 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X2 U4937 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  OAI21_X1 U4938 ( .B1(n4613), .B2(n8362), .A(n4612), .ZN(n4611) );
  XNOR2_X1 U4939 ( .A(n4764), .B(n8448), .ZN(n8901) );
  NAND2_X1 U4940 ( .A1(n4720), .A2(n4721), .ZN(n4584) );
  INV_X1 U4941 ( .A(n6156), .ZN(n4582) );
  NAND2_X1 U4942 ( .A1(n8661), .A2(n8443), .ZN(n4764) );
  OAI21_X1 U4943 ( .B1(n4669), .B2(n4474), .A(n4670), .ZN(n4666) );
  AOI21_X1 U4944 ( .B1(n8453), .B2(n9777), .A(n8452), .ZN(n8900) );
  NAND2_X1 U4945 ( .A1(n9077), .A2(n4917), .ZN(n4915) );
  AOI211_X1 U4946 ( .C1(n9774), .C2(n8695), .A(n8694), .B(n8693), .ZN(n8910)
         );
  AND2_X1 U4947 ( .A1(n4890), .A2(n6357), .ZN(n8449) );
  AOI21_X1 U4948 ( .B1(n8676), .B2(n9777), .A(n8675), .ZN(n8905) );
  OR2_X1 U4949 ( .A1(n8735), .A2(n8742), .ZN(n4755) );
  AND2_X1 U4950 ( .A1(n4843), .A2(n4841), .ZN(n8461) );
  OAI21_X1 U4951 ( .B1(n9242), .B2(n8397), .A(n8246), .ZN(n9226) );
  OAI21_X1 U4952 ( .B1(n4411), .B2(n8343), .A(n4585), .ZN(n9242) );
  AOI21_X1 U4953 ( .B1(n4533), .B2(n4537), .A(n4466), .ZN(n4531) );
  NAND2_X1 U4954 ( .A1(n8812), .A2(n4427), .ZN(n8796) );
  NOR2_X1 U4955 ( .A1(n8209), .A2(n4402), .ZN(n4585) );
  NOR2_X1 U4956 ( .A1(n6371), .A2(n6226), .ZN(n6367) );
  XNOR2_X1 U4957 ( .A(n5511), .B(n5530), .ZN(n8034) );
  NAND2_X1 U4958 ( .A1(n8813), .A2(n8820), .ZN(n8812) );
  AOI21_X1 U4959 ( .B1(n4753), .B2(n4757), .A(n4751), .ZN(n4750) );
  OAI21_X1 U4960 ( .B1(n8138), .B2(n8137), .A(n8136), .ZN(n9375) );
  AND2_X1 U4961 ( .A1(n4526), .A2(n4450), .ZN(n8813) );
  XNOR2_X1 U4962 ( .A(n4478), .B(n6202), .ZN(n8138) );
  NAND2_X1 U4963 ( .A1(n4804), .A2(n4807), .ZN(n9322) );
  AND2_X1 U4964 ( .A1(n9358), .A2(n8333), .ZN(n9345) );
  INV_X1 U4965 ( .A(n4711), .ZN(n4710) );
  NAND2_X1 U4966 ( .A1(n4880), .A2(n6338), .ZN(n4878) );
  OR2_X1 U4967 ( .A1(n4714), .A2(n8200), .ZN(n4713) );
  AND2_X1 U4968 ( .A1(n6344), .A2(n6343), .ZN(n8742) );
  OR2_X1 U4969 ( .A1(n8922), .A2(n8505), .ZN(n6344) );
  NAND2_X1 U4970 ( .A1(n6011), .A2(n6010), .ZN(n9398) );
  NAND2_X1 U4971 ( .A1(n6338), .A2(n6337), .ZN(n8775) );
  AOI21_X1 U4972 ( .B1(n7843), .B2(n6169), .A(n4959), .ZN(n7922) );
  NAND2_X1 U4973 ( .A1(n5994), .A2(n5993), .ZN(n9408) );
  XNOR2_X1 U4974 ( .A(n5541), .B(n5555), .ZN(n7458) );
  NAND2_X1 U4975 ( .A1(n7683), .A2(n7684), .ZN(n7682) );
  NAND2_X1 U4976 ( .A1(n5983), .A2(n5982), .ZN(n9413) );
  NAND2_X1 U4977 ( .A1(n5540), .A2(n5556), .ZN(n5541) );
  NOR2_X1 U4978 ( .A1(n8855), .A2(n4874), .ZN(n4873) );
  NAND2_X1 U4979 ( .A1(n5966), .A2(n5965), .ZN(n9423) );
  AND2_X1 U4980 ( .A1(n8183), .A2(n5932), .ZN(n8188) );
  NAND2_X1 U4981 ( .A1(n6313), .A2(n6314), .ZN(n8855) );
  OR2_X1 U4982 ( .A1(n7780), .A2(n7781), .ZN(n4790) );
  NAND2_X1 U4983 ( .A1(n5421), .A2(n5420), .ZN(n8953) );
  OR2_X1 U4984 ( .A1(n8960), .A2(n8830), .ZN(n6313) );
  NAND2_X1 U4985 ( .A1(n5103), .A2(n5102), .ZN(n8522) );
  OR2_X1 U4986 ( .A1(n8964), .A2(n8883), .ZN(n6309) );
  AND2_X1 U4987 ( .A1(n7920), .A2(n6305), .ZN(n8863) );
  NAND2_X1 U4988 ( .A1(n5064), .A2(n5063), .ZN(n8960) );
  AND2_X1 U4989 ( .A1(n6300), .A2(n7846), .ZN(n7834) );
  OR2_X1 U4990 ( .A1(n9491), .A2(n7999), .ZN(n7920) );
  NAND2_X1 U4991 ( .A1(n5116), .A2(n5115), .ZN(n8964) );
  OAI21_X1 U4992 ( .B1(n5414), .B2(n4586), .A(n5418), .ZN(n5438) );
  NAND2_X1 U4993 ( .A1(n5140), .A2(n5139), .ZN(n9491) );
  OAI21_X1 U4994 ( .B1(n5110), .B2(n5043), .A(n5042), .ZN(n5414) );
  NAND2_X1 U4995 ( .A1(n5880), .A2(n5879), .ZN(n9532) );
  NAND2_X1 U4996 ( .A1(n6280), .A2(n6281), .ZN(n7492) );
  OAI21_X1 U4997 ( .B1(n5134), .B2(n5030), .A(n5029), .ZN(n5110) );
  NAND2_X1 U4998 ( .A1(n4597), .A2(n4596), .ZN(n9634) );
  OR2_X1 U4999 ( .A1(n7687), .A2(n7779), .ZN(n6287) );
  INV_X1 U5000 ( .A(n6163), .ZN(n7714) );
  OAI21_X1 U5001 ( .B1(n5386), .B2(n5014), .A(n5013), .ZN(n5169) );
  OAI21_X1 U5002 ( .B1(n5010), .B2(n4829), .A(n4433), .ZN(n5154) );
  XNOR2_X1 U5003 ( .A(n5359), .B(n5358), .ZN(n6494) );
  NOR2_X1 U5004 ( .A1(n6113), .A2(n8315), .ZN(n9656) );
  NAND2_X2 U5005 ( .A1(n7039), .A2(n9629), .ZN(n9665) );
  OR2_X1 U5006 ( .A1(n9648), .A2(n9651), .ZN(n9649) );
  NAND2_X2 U5007 ( .A1(n6990), .A2(n9778), .ZN(n8870) );
  NAND2_X1 U5008 ( .A1(n5321), .A2(n5320), .ZN(n4995) );
  NAND2_X1 U5009 ( .A1(n4475), .A2(n4990), .ZN(n5321) );
  NAND2_X1 U5010 ( .A1(n4413), .A2(n5258), .ZN(n8584) );
  NAND2_X1 U5011 ( .A1(n4476), .A2(n4987), .ZN(n5301) );
  AND4_X1 U5012 ( .A1(n5202), .A2(n5201), .A3(n5200), .A4(n5199), .ZN(n8422)
         );
  AND4_X1 U5013 ( .A1(n5280), .A2(n5279), .A3(n5278), .A4(n5277), .ZN(n8547)
         );
  NAND2_X1 U5014 ( .A1(n6978), .A2(n5077), .ZN(n5197) );
  NAND2_X1 U5015 ( .A1(n6159), .A2(n7102), .ZN(n6252) );
  NAND4_X1 U5016 ( .A1(n5234), .A2(n5233), .A3(n5232), .A4(n5231), .ZN(n8585)
         );
  AND3_X1 U5017 ( .A1(n5243), .A2(n5242), .A3(n5241), .ZN(n7117) );
  AND2_X1 U5018 ( .A1(n4639), .A2(n4638), .ZN(n6646) );
  AND2_X1 U5019 ( .A1(n5764), .A2(n4594), .ZN(n9676) );
  INV_X1 U5020 ( .A(n7098), .ZN(n7008) );
  NAND2_X1 U5021 ( .A1(n4815), .A2(n4674), .ZN(n7142) );
  OAI211_X1 U5022 ( .C1(n6562), .C2(n6579), .A(n5196), .B(n5195), .ZN(n7098)
         );
  NAND4_X1 U5023 ( .A1(n5760), .A2(n5759), .A3(n5758), .A4(n5757), .ZN(n9129)
         );
  NOR2_X1 U5024 ( .A1(n6147), .A2(n4486), .ZN(n6716) );
  XNOR2_X1 U5025 ( .A(n5076), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8714) );
  AND2_X1 U5026 ( .A1(n6086), .A2(n6087), .ZN(n6081) );
  NAND2_X2 U5027 ( .A1(n5736), .A2(n5735), .ZN(n5791) );
  INV_X1 U5028 ( .A(n5083), .ZN(n5091) );
  XNOR2_X1 U5029 ( .A(n5082), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5083) );
  NAND2_X1 U5030 ( .A1(n5778), .A2(n6051), .ZN(n8137) );
  MUX2_X1 U5031 ( .A(n6693), .B(n6459), .S(n5778), .Z(n7148) );
  NAND2_X1 U5032 ( .A1(n4522), .A2(n5703), .ZN(n5715) );
  NAND2_X1 U5033 ( .A1(n8005), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5732) );
  INV_X1 U5034 ( .A(n5933), .ZN(n4522) );
  NAND2_X1 U5035 ( .A1(n4826), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5743) );
  XNOR2_X1 U5036 ( .A(n5055), .B(n10177), .ZN(n7677) );
  NAND2_X1 U5037 ( .A1(n5054), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5055) );
  NOR2_X1 U5038 ( .A1(n4541), .A2(n4540), .ZN(n4539) );
  AND3_X1 U5039 ( .A1(n5298), .A2(n4397), .A3(n4452), .ZN(n5170) );
  INV_X2 U5040 ( .A(n7450), .ZN(n4390) );
  AND4_X1 U5041 ( .A1(n5697), .A2(n4511), .A3(n4510), .A4(n5696), .ZN(n5899)
         );
  NAND2_X1 U5042 ( .A1(n5192), .A2(n4430), .ZN(n6579) );
  INV_X1 U5043 ( .A(n4540), .ZN(n5298) );
  AND2_X1 U5044 ( .A1(n4905), .A2(n4904), .ZN(n4903) );
  AND2_X1 U5045 ( .A1(n4509), .A2(n5699), .ZN(n4511) );
  INV_X1 U5046 ( .A(n4980), .ZN(n4391) );
  AND4_X1 U5047 ( .A1(n5068), .A2(n5059), .A3(n5057), .A4(n5061), .ZN(n5049)
         );
  AND4_X1 U5048 ( .A1(n5046), .A2(n5112), .A3(n5387), .A4(n5368), .ZN(n5050)
         );
  AND2_X1 U5049 ( .A1(n5045), .A2(n4906), .ZN(n4905) );
  AND4_X1 U5050 ( .A1(n5695), .A2(n10118), .A3(n5807), .A4(n5694), .ZN(n5696)
         );
  AND3_X1 U5051 ( .A1(n5864), .A2(n5836), .A3(n5698), .ZN(n4509) );
  AND2_X1 U5052 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7651) );
  INV_X1 U5053 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5722) );
  NOR2_X1 U5054 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5761) );
  INV_X1 U5055 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5912) );
  NOR2_X1 U5056 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5693) );
  INV_X1 U5057 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5724) );
  NOR2_X2 U5058 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5191) );
  INV_X1 U5059 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5112) );
  NOR2_X1 U5060 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4907) );
  INV_X1 U5061 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5387) );
  INV_X1 U5062 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5368) );
  NOR2_X1 U5063 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5046) );
  XNOR2_X2 U5064 ( .A(n5708), .B(n5724), .ZN(n9350) );
  XNOR2_X2 U5065 ( .A(n5743), .B(n5742), .ZN(n6068) );
  AND2_X4 U5066 ( .A1(n6691), .A2(n6773), .ZN(n6707) );
  OAI21_X2 U5067 ( .B1(n8819), .B2(n6174), .A(n6331), .ZN(n8789) );
  NOR2_X2 U5068 ( .A1(n8821), .A2(n8820), .ZN(n8819) );
  INV_X1 U5069 ( .A(n8551), .ZN(n5244) );
  INV_X1 U5070 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6083) );
  NAND2_X1 U5071 ( .A1(n5438), .A2(n5437), .ZN(n5441) );
  NAND2_X1 U5073 ( .A1(n4796), .A2(n4795), .ZN(n9200) );
  AOI21_X1 U5074 ( .B1(n4797), .B2(n4801), .A(n4438), .ZN(n4795) );
  OR2_X1 U5075 ( .A1(n8279), .A2(n6068), .ZN(n9660) );
  AOI21_X1 U5076 ( .B1(n4661), .B2(n6350), .A(n4660), .ZN(n4659) );
  INV_X1 U5077 ( .A(n6355), .ZN(n4660) );
  INV_X1 U5078 ( .A(n6370), .ZN(n4891) );
  NAND2_X1 U5079 ( .A1(n5367), .A2(n5366), .ZN(n5010) );
  NAND2_X1 U5080 ( .A1(n4997), .A2(n4996), .ZN(n5000) );
  NAND2_X1 U5081 ( .A1(n8494), .A2(n4854), .ZN(n4853) );
  INV_X1 U5082 ( .A(n5602), .ZN(n5629) );
  NAND2_X1 U5083 ( .A1(n4861), .A2(n5407), .ZN(n7995) );
  INV_X1 U5084 ( .A(n7939), .ZN(n4861) );
  OR2_X1 U5085 ( .A1(n8919), .A2(n8747), .ZN(n8703) );
  OR2_X1 U5086 ( .A1(n8759), .A2(n8746), .ZN(n4955) );
  OAI21_X1 U5087 ( .B1(n8804), .B2(n4776), .A(n8438), .ZN(n4775) );
  OR2_X1 U5088 ( .A1(n8942), .A2(n8496), .ZN(n6331) );
  NAND2_X1 U5089 ( .A1(n4872), .A2(n6313), .ZN(n4871) );
  NAND2_X1 U5090 ( .A1(n4873), .A2(n6312), .ZN(n4872) );
  OR3_X1 U5091 ( .A1(n5395), .A2(n5174), .A3(n7243), .ZN(n5159) );
  INV_X1 U5092 ( .A(n7487), .ZN(n7488) );
  INV_X1 U5093 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n4906) );
  INV_X1 U5094 ( .A(n8088), .ZN(n4923) );
  NAND2_X1 U5095 ( .A1(n8407), .A2(n8144), .ZN(n8354) );
  INV_X1 U5096 ( .A(n7799), .ZN(n5735) );
  INV_X1 U5097 ( .A(n5737), .ZN(n5736) );
  NOR2_X1 U5098 ( .A1(n6921), .A2(n4472), .ZN(n6406) );
  AND2_X1 U5099 ( .A1(n6144), .A2(n4451), .ZN(n4802) );
  OAI21_X1 U5100 ( .B1(n6183), .B2(n6182), .A(n6186), .ZN(n6198) );
  OAI21_X1 U5101 ( .B1(n5577), .B2(n5576), .A(n5575), .ZN(n5594) );
  AND2_X1 U5102 ( .A1(n5574), .A2(n5573), .ZN(n5575) );
  INV_X1 U5103 ( .A(n5415), .ZN(n4586) );
  NAND2_X1 U5104 ( .A1(n4772), .A2(n4994), .ZN(n4771) );
  INV_X1 U5105 ( .A(n5340), .ZN(n4772) );
  NOR2_X1 U5106 ( .A1(n5511), .A2(n4559), .ZN(n8473) );
  INV_X1 U5107 ( .A(n5530), .ZN(n4559) );
  NAND2_X1 U5108 ( .A1(n8551), .A2(n5246), .ZN(n5247) );
  NAND2_X1 U5109 ( .A1(n5632), .A2(n8649), .ZN(n6383) );
  INV_X2 U5110 ( .A(n5213), .ZN(n6189) );
  AND4_X1 U5111 ( .A1(n5380), .A2(n5379), .A3(n5378), .A4(n5377), .ZN(n7687)
         );
  NAND2_X2 U5112 ( .A1(n5085), .A2(n5091), .ZN(n5349) );
  NOR2_X1 U5113 ( .A1(n9469), .A2(n9468), .ZN(n9467) );
  OR2_X1 U5114 ( .A1(n6615), .A2(n6614), .ZN(n4637) );
  AND2_X1 U5115 ( .A1(n6361), .A2(n6362), .ZN(n8448) );
  NAND2_X1 U5116 ( .A1(n8753), .A2(n4955), .ZN(n8735) );
  XNOR2_X1 U5117 ( .A(n8927), .B(n8746), .ZN(n8754) );
  NAND2_X1 U5118 ( .A1(n4881), .A2(n6333), .ZN(n4880) );
  NAND2_X1 U5119 ( .A1(n4785), .A2(n4783), .ZN(n8841) );
  NOR2_X1 U5120 ( .A1(n4784), .A2(n8433), .ZN(n4783) );
  INV_X1 U5121 ( .A(n6168), .ZN(n6167) );
  NAND2_X1 U5122 ( .A1(n7929), .A2(n4956), .ZN(n8864) );
  INV_X1 U5123 ( .A(n9772), .ZN(n8880) );
  NAND2_X1 U5124 ( .A1(n6178), .A2(n6177), .ZN(n8898) );
  AND2_X1 U5125 ( .A1(n5632), .A2(n6991), .ZN(n9819) );
  NAND2_X1 U5126 ( .A1(n5069), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5076) );
  NAND2_X1 U5127 ( .A1(n4492), .A2(n4491), .ZN(n7284) );
  NAND2_X1 U5128 ( .A1(n4495), .A2(n4498), .ZN(n4491) );
  NAND2_X1 U5129 ( .A1(n7214), .A2(n7213), .ZN(n7212) );
  AND2_X1 U5130 ( .A1(n8143), .A2(n8142), .ZN(n9194) );
  AND2_X1 U5131 ( .A1(n6054), .A2(n6053), .ZN(n8236) );
  INV_X1 U5132 ( .A(n4808), .ZN(n4807) );
  NAND2_X1 U5133 ( .A1(n6133), .A2(n4805), .ZN(n4804) );
  OAI21_X1 U5134 ( .B1(n4809), .B2(n4410), .A(n6136), .ZN(n4808) );
  INV_X1 U5135 ( .A(n8137), .ZN(n8139) );
  NAND2_X1 U5136 ( .A1(n9659), .A2(n9688), .ZN(n8256) );
  INV_X1 U5137 ( .A(n9127), .ZN(n9659) );
  XNOR2_X1 U5138 ( .A(n4793), .B(n8276), .ZN(n9379) );
  AND2_X1 U5139 ( .A1(n9383), .A2(n9117), .ZN(n6145) );
  INV_X1 U5140 ( .A(n9718), .ZN(n9689) );
  NAND2_X1 U5141 ( .A1(n6073), .A2(n4589), .ZN(n4826) );
  AND2_X1 U5142 ( .A1(n5730), .A2(n5745), .ZN(n4589) );
  NAND2_X1 U5143 ( .A1(n7651), .A2(n4857), .ZN(n4480) );
  NAND2_X1 U5144 ( .A1(n7652), .A2(n4966), .ZN(n4481) );
  INV_X1 U5145 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4857) );
  NAND2_X1 U5146 ( .A1(n4720), .A2(n4721), .ZN(n4678) );
  NAND2_X1 U5147 ( .A1(n4673), .A2(n4672), .ZN(n6263) );
  NAND2_X1 U5148 ( .A1(n6260), .A2(n6372), .ZN(n4673) );
  NAND2_X1 U5149 ( .A1(n6234), .A2(n6360), .ZN(n4672) );
  NOR2_X1 U5150 ( .A1(n5860), .A2(n8232), .ZN(n4609) );
  NAND2_X1 U5151 ( .A1(n8264), .A2(n4607), .ZN(n4606) );
  NAND2_X1 U5152 ( .A1(n8156), .A2(n4608), .ZN(n4607) );
  OR2_X1 U5153 ( .A1(n8163), .A2(n8164), .ZN(n4605) );
  OAI22_X1 U5154 ( .A1(n8330), .A2(n4608), .B1(n8193), .B2(n4619), .ZN(n4617)
         );
  NOR2_X1 U5155 ( .A1(n4622), .A2(n8232), .ZN(n4621) );
  NOR2_X1 U5156 ( .A1(n4624), .A2(n4625), .ZN(n4622) );
  AND2_X1 U5157 ( .A1(n8196), .A2(n8195), .ZN(n4625) );
  INV_X1 U5158 ( .A(n4624), .ZN(n4623) );
  NAND2_X1 U5159 ( .A1(n8329), .A2(n8232), .ZN(n4619) );
  INV_X1 U5160 ( .A(n4621), .ZN(n4620) );
  AND2_X1 U5161 ( .A1(n4653), .A2(n4651), .ZN(n4650) );
  NAND2_X1 U5162 ( .A1(n4420), .A2(n4784), .ZN(n4651) );
  INV_X1 U5163 ( .A(n6318), .ZN(n4653) );
  INV_X1 U5164 ( .A(n4646), .ZN(n4645) );
  AND2_X1 U5165 ( .A1(n4650), .A2(n6323), .ZN(n4646) );
  AOI21_X1 U5166 ( .B1(n8197), .B2(n8201), .A(n8248), .ZN(n4593) );
  NAND2_X1 U5167 ( .A1(n4592), .A2(n4590), .ZN(n8206) );
  OAI21_X1 U5168 ( .B1(n4591), .B2(n8248), .A(n8232), .ZN(n4590) );
  OAI21_X1 U5169 ( .B1(n4593), .B2(n8247), .A(n4608), .ZN(n4592) );
  AOI21_X1 U5170 ( .B1(n8199), .B2(n8331), .A(n4442), .ZN(n4591) );
  AOI21_X1 U5171 ( .B1(n4664), .B2(n4662), .A(n8681), .ZN(n4661) );
  INV_X1 U5172 ( .A(n6352), .ZN(n4662) );
  OR2_X1 U5173 ( .A1(n8099), .A2(n8098), .ZN(n8100) );
  NOR2_X1 U5174 ( .A1(n9054), .A2(n8093), .ZN(n4912) );
  AND2_X1 U5175 ( .A1(n8318), .A2(n4742), .ZN(n4598) );
  INV_X1 U5176 ( .A(n5358), .ZN(n4769) );
  NAND2_X1 U5177 ( .A1(n5002), .A2(n5001), .ZN(n5005) );
  NAND2_X1 U5178 ( .A1(n4859), .A2(n5180), .ZN(n5406) );
  XNOR2_X1 U5179 ( .A(n6166), .B(n5629), .ZN(n5167) );
  NOR2_X1 U5180 ( .A1(n4855), .A2(n4850), .ZN(n4849) );
  INV_X1 U5181 ( .A(n5463), .ZN(n4850) );
  NAND2_X1 U5182 ( .A1(n8494), .A2(n4856), .ZN(n4855) );
  INV_X1 U5183 ( .A(n8559), .ZN(n4856) );
  NOR2_X1 U5184 ( .A1(n4842), .A2(n6453), .ZN(n4841) );
  INV_X1 U5185 ( .A(n4844), .ZN(n4842) );
  NAND2_X1 U5186 ( .A1(n4656), .A2(n4658), .ZN(n4655) );
  INV_X1 U5187 ( .A(n6372), .ZN(n6360) );
  NOR2_X1 U5188 ( .A1(n4891), .A2(n4892), .ZN(n4889) );
  NAND2_X1 U5189 ( .A1(n6374), .A2(n4425), .ZN(n4886) );
  NOR2_X1 U5190 ( .A1(n4884), .A2(n4477), .ZN(n4883) );
  AND2_X1 U5191 ( .A1(n4887), .A2(n6367), .ZN(n4477) );
  AOI22_X1 U5192 ( .A1(n4891), .A2(n6180), .B1(n4892), .B2(n4888), .ZN(n4887)
         );
  OR2_X1 U5193 ( .A1(n8907), .A2(n8707), .ZN(n6353) );
  OR2_X1 U5194 ( .A1(n8914), .A2(n8687), .ZN(n6347) );
  OR2_X1 U5195 ( .A1(n5490), .A2(n10151), .ZN(n5523) );
  NAND2_X1 U5196 ( .A1(n4444), .A2(n8802), .ZN(n4695) );
  INV_X1 U5197 ( .A(n4869), .ZN(n4865) );
  INV_X1 U5198 ( .A(n6315), .ZN(n4874) );
  NOR2_X1 U5199 ( .A1(n9491), .A2(n6166), .ZN(n4708) );
  NAND2_X1 U5200 ( .A1(n5088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5395) );
  AND2_X1 U5201 ( .A1(n7584), .A2(n7583), .ZN(n7778) );
  INV_X1 U5202 ( .A(n7224), .ZN(n4524) );
  NAND2_X1 U5203 ( .A1(n9752), .A2(n8550), .ZN(n6236) );
  NAND2_X1 U5204 ( .A1(n5298), .A2(n4397), .ZN(n5360) );
  NOR2_X1 U5205 ( .A1(n4497), .A2(n4496), .ZN(n4495) );
  INV_X1 U5206 ( .A(n7064), .ZN(n4496) );
  NOR2_X1 U5207 ( .A1(n6938), .A2(n4498), .ZN(n4497) );
  AND2_X1 U5208 ( .A1(n4929), .A2(n4502), .ZN(n4501) );
  NAND2_X1 U5209 ( .A1(n4503), .A2(n7956), .ZN(n4502) );
  NOR2_X1 U5210 ( .A1(n4436), .A2(n4930), .ZN(n4929) );
  INV_X1 U5211 ( .A(n7902), .ZN(n4503) );
  INV_X1 U5212 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5698) );
  INV_X1 U5213 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5695) );
  OR2_X1 U5214 ( .A1(n9388), .A2(n9107), .ZN(n8346) );
  INV_X1 U5215 ( .A(n8345), .ZN(n8246) );
  NOR2_X1 U5216 ( .A1(n9405), .A2(n9398), .ZN(n4680) );
  INV_X1 U5217 ( .A(n9266), .ZN(n4736) );
  NOR2_X1 U5218 ( .A1(n6138), .A2(n4822), .ZN(n4820) );
  INV_X1 U5219 ( .A(n4824), .ZN(n4817) );
  NAND2_X1 U5220 ( .A1(n8388), .A2(n8341), .ZN(n5999) );
  NAND2_X1 U5221 ( .A1(n9342), .A2(n8249), .ZN(n4712) );
  OR2_X1 U5222 ( .A1(n9420), .A2(n9083), .ZN(n8331) );
  OR2_X1 U5223 ( .A1(n9423), .A2(n9318), .ZN(n8250) );
  AND2_X1 U5224 ( .A1(n8269), .A2(n8293), .ZN(n4728) );
  NAND2_X1 U5225 ( .A1(n7473), .A2(n4728), .ZN(n7725) );
  INV_X1 U5226 ( .A(n9634), .ZN(n8152) );
  INV_X1 U5227 ( .A(n8256), .ZN(n4745) );
  OR2_X1 U5228 ( .A1(n5784), .A2(n5765), .ZN(n5767) );
  INV_X1 U5229 ( .A(n9129), .ZN(n7160) );
  NAND2_X1 U5230 ( .A1(n4484), .A2(n6050), .ZN(n6183) );
  NAND2_X1 U5231 ( .A1(n6047), .A2(n6046), .ZN(n4484) );
  AND4_X1 U5232 ( .A1(n10117), .A2(n5729), .A3(n5728), .A4(n6083), .ZN(n5730)
         );
  AND2_X1 U5233 ( .A1(n5539), .A2(n5538), .ZN(n5556) );
  NAND2_X1 U5234 ( .A1(n4482), .A2(n4574), .ZN(n5502) );
  AOI21_X1 U5235 ( .B1(n4577), .B2(n4579), .A(n4575), .ZN(n4574) );
  NAND2_X1 U5236 ( .A1(n5441), .A2(n4577), .ZN(n4482) );
  INV_X1 U5237 ( .A(n5486), .ZN(n4575) );
  INV_X1 U5238 ( .A(n4832), .ZN(n4829) );
  NAND2_X1 U5239 ( .A1(n4832), .A2(n4828), .ZN(n4827) );
  INV_X1 U5240 ( .A(n5000), .ZN(n4770) );
  NAND2_X1 U5241 ( .A1(n5000), .A2(n4999), .ZN(n5340) );
  NAND2_X1 U5242 ( .A1(n4748), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4968) );
  INV_X1 U5243 ( .A(n5755), .ZN(n4748) );
  NOR2_X1 U5244 ( .A1(n4839), .A2(n4838), .ZN(n4837) );
  INV_X1 U5245 ( .A(n5592), .ZN(n4839) );
  NOR2_X1 U5246 ( .A1(n4840), .A2(n4845), .ZN(n4838) );
  INV_X1 U5247 ( .A(n4841), .ZN(n4840) );
  AND2_X1 U5248 ( .A1(n7938), .A2(n5183), .ZN(n7939) );
  NAND2_X1 U5249 ( .A1(n4848), .A2(n5435), .ZN(n4847) );
  INV_X1 U5250 ( .A(n7949), .ZN(n4848) );
  AND2_X1 U5251 ( .A1(n5328), .A2(n5309), .ZN(n4550) );
  NOR2_X1 U5252 ( .A1(n5483), .A2(n5482), .ZN(n4854) );
  AOI22_X1 U5253 ( .A1(n8031), .A2(n5533), .B1(n5532), .B2(n5531), .ZN(n5550)
         );
  NAND2_X1 U5254 ( .A1(n8543), .A2(n5268), .ZN(n8542) );
  NAND2_X1 U5255 ( .A1(n4547), .A2(n7544), .ZN(n4546) );
  INV_X1 U5256 ( .A(n7556), .ZN(n4547) );
  NOR2_X1 U5257 ( .A1(n7540), .A2(n4549), .ZN(n4548) );
  INV_X1 U5258 ( .A(n5348), .ZN(n4549) );
  AND4_X1 U5259 ( .A1(n5479), .A2(n5478), .A3(n5477), .A4(n5476), .ZN(n8496)
         );
  NOR2_X1 U5260 ( .A1(n9467), .A2(n4414), .ZN(n6635) );
  OR2_X1 U5261 ( .A1(n6635), .A2(n6634), .ZN(n4627) );
  NOR2_X1 U5262 ( .A1(n6667), .A2(n4435), .ZN(n6573) );
  OR2_X1 U5263 ( .A1(n6573), .A2(n6572), .ZN(n4639) );
  AND2_X1 U5264 ( .A1(n4637), .A2(n4636), .ZN(n6813) );
  NAND2_X1 U5265 ( .A1(n6810), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4636) );
  OR2_X1 U5266 ( .A1(n6813), .A2(n6812), .ZN(n4635) );
  NOR2_X1 U5267 ( .A1(n8629), .A2(n4630), .ZN(n8641) );
  AND2_X1 U5268 ( .A1(n8630), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4630) );
  OR2_X1 U5269 ( .A1(n8907), .A2(n8672), .ZN(n8441) );
  NAND2_X1 U5270 ( .A1(n8914), .A2(n8687), .ZN(n8689) );
  NAND2_X1 U5271 ( .A1(n6347), .A2(n8689), .ZN(n8704) );
  AOI21_X1 U5272 ( .B1(n4756), .B2(n4754), .A(n4446), .ZN(n4753) );
  INV_X1 U5273 ( .A(n4760), .ZN(n4754) );
  NAND2_X1 U5274 ( .A1(n8742), .A2(n4760), .ZN(n4758) );
  NOR2_X1 U5275 ( .A1(n4536), .A2(n4534), .ZN(n4533) );
  AND2_X1 U5276 ( .A1(n4753), .A2(n4535), .ZN(n4534) );
  INV_X1 U5277 ( .A(n4750), .ZN(n4536) );
  INV_X1 U5278 ( .A(n4955), .ZN(n4535) );
  INV_X1 U5279 ( .A(n4753), .ZN(n4537) );
  NAND2_X1 U5280 ( .A1(n8703), .A2(n6227), .ZN(n8720) );
  NAND2_X1 U5281 ( .A1(n4761), .A2(n8505), .ZN(n4760) );
  NAND2_X1 U5282 ( .A1(n8735), .A2(n4760), .ZN(n4752) );
  NOR2_X1 U5283 ( .A1(n8769), .A2(n8927), .ZN(n8756) );
  NOR2_X1 U5284 ( .A1(n8932), .A2(n8439), .ZN(n8440) );
  NOR2_X1 U5285 ( .A1(n8789), .A2(n8788), .ZN(n4882) );
  NAND2_X1 U5286 ( .A1(n8796), .A2(n8804), .ZN(n8795) );
  INV_X1 U5287 ( .A(n4871), .ZN(n4868) );
  NOR2_X1 U5288 ( .A1(n4871), .A2(n8827), .ZN(n4869) );
  NAND2_X1 U5289 ( .A1(n7980), .A2(n4873), .ZN(n4870) );
  AND2_X1 U5290 ( .A1(n8522), .A2(n8575), .ZN(n8433) );
  NOR2_X1 U5291 ( .A1(n7986), .A2(n4787), .ZN(n4786) );
  NOR2_X1 U5292 ( .A1(n7839), .A2(n7844), .ZN(n4528) );
  AND2_X1 U5293 ( .A1(n7867), .A2(n9852), .ZN(n7857) );
  NOR2_X1 U5294 ( .A1(n4897), .A2(n4895), .ZN(n4894) );
  INV_X1 U5295 ( .A(n6288), .ZN(n4895) );
  INV_X1 U5296 ( .A(n6298), .ZN(n4897) );
  NAND2_X1 U5297 ( .A1(n7580), .A2(n7579), .ZN(n7586) );
  NOR2_X1 U5298 ( .A1(n7586), .A2(n7585), .ZN(n7780) );
  OAI21_X1 U5299 ( .B1(n9782), .B2(n7327), .A(n7326), .ZN(n7486) );
  AND2_X1 U5300 ( .A1(n5688), .A2(n6561), .ZN(n9772) );
  OR2_X1 U5301 ( .A1(n6203), .A2(n6468), .ZN(n5195) );
  NAND2_X1 U5302 ( .A1(n5622), .A2(n5621), .ZN(n8902) );
  AND2_X1 U5303 ( .A1(n5632), .A2(n5633), .ZN(n9845) );
  NAND2_X1 U5304 ( .A1(n4903), .A2(n5051), .ZN(n4541) );
  NAND2_X1 U5305 ( .A1(n5067), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5419) );
  AND2_X1 U5306 ( .A1(n5298), .A2(n4905), .ZN(n5056) );
  NAND2_X1 U5307 ( .A1(n4632), .A2(n8011), .ZN(n4631) );
  INV_X1 U5308 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4632) );
  NAND2_X1 U5309 ( .A1(n6737), .A2(n6736), .ZN(n6739) );
  NAND2_X1 U5310 ( .A1(n9003), .A2(n8114), .ZN(n4942) );
  AND2_X1 U5311 ( .A1(n8093), .A2(n9080), .ZN(n4917) );
  AND2_X1 U5312 ( .A1(n8093), .A2(n4923), .ZN(n4916) );
  NAND2_X1 U5313 ( .A1(n4946), .A2(n4945), .ZN(n7342) );
  AND2_X1 U5314 ( .A1(n7286), .A2(n4947), .ZN(n4945) );
  INV_X1 U5315 ( .A(n9018), .ZN(n4928) );
  NAND2_X1 U5316 ( .A1(n4919), .A2(n4923), .ZN(n4922) );
  NAND2_X1 U5317 ( .A1(n7424), .A2(n7423), .ZN(n4508) );
  INV_X1 U5318 ( .A(n9244), .ZN(n9107) );
  AND4_X1 U5319 ( .A1(n6062), .A2(n6061), .A3(n6060), .A4(n6059), .ZN(n8230)
         );
  NOR2_X1 U5320 ( .A1(n6601), .A2(n6600), .ZN(n6599) );
  NAND2_X1 U5321 ( .A1(n7212), .A2(n6407), .ZN(n7604) );
  OR2_X1 U5322 ( .A1(n7609), .A2(n7608), .ZN(n4566) );
  AOI21_X1 U5323 ( .B1(n4800), .B2(n4802), .A(n4445), .ZN(n4799) );
  INV_X1 U5324 ( .A(n9257), .ZN(n4800) );
  INV_X1 U5325 ( .A(n4802), .ZN(n4801) );
  NAND2_X1 U5326 ( .A1(n9254), .A2(n9268), .ZN(n6144) );
  NAND2_X1 U5327 ( .A1(n8396), .A2(n8398), .ZN(n9257) );
  AOI21_X1 U5328 ( .B1(n4739), .B2(n8248), .A(n4738), .ZN(n4737) );
  INV_X1 U5329 ( .A(n8388), .ZN(n4738) );
  AND2_X1 U5330 ( .A1(n9408), .A2(n9905), .ZN(n6139) );
  NAND2_X1 U5331 ( .A1(n9283), .A2(n9269), .ZN(n6140) );
  INV_X1 U5332 ( .A(n5999), .ZN(n9284) );
  NOR2_X1 U5333 ( .A1(n9314), .A2(n5981), .ZN(n9300) );
  NOR2_X1 U5334 ( .A1(n9306), .A2(n4825), .ZN(n4824) );
  INV_X1 U5335 ( .A(n4961), .ZN(n4825) );
  OAI22_X1 U5336 ( .A1(n9306), .A2(n4823), .B1(n9309), .B2(n9083), .ZN(n4822)
         );
  INV_X1 U5337 ( .A(n4965), .ZN(n4823) );
  NOR2_X1 U5338 ( .A1(n9315), .A2(n9316), .ZN(n9314) );
  AND2_X1 U5339 ( .A1(n8331), .A2(n8201), .ZN(n9306) );
  NAND2_X1 U5340 ( .A1(n4715), .A2(n8326), .ZN(n4714) );
  NAND2_X1 U5341 ( .A1(n9339), .A2(n5963), .ZN(n4715) );
  NOR2_X1 U5342 ( .A1(n6134), .A2(n4813), .ZN(n4812) );
  INV_X1 U5343 ( .A(n4957), .ZN(n4813) );
  NAND2_X1 U5344 ( .A1(n4810), .A2(n4814), .ZN(n4809) );
  INV_X1 U5345 ( .A(n9360), .ZN(n4810) );
  OR2_X1 U5346 ( .A1(n7888), .A2(n9362), .ZN(n4957) );
  NAND2_X1 U5347 ( .A1(n7887), .A2(n6132), .ZN(n6133) );
  NAND2_X1 U5348 ( .A1(n9512), .A2(n8183), .ZN(n7887) );
  AND2_X1 U5349 ( .A1(n8297), .A2(n8295), .ZN(n8269) );
  NOR2_X1 U5350 ( .A1(n5860), .A2(n4733), .ZN(n4732) );
  INV_X1 U5351 ( .A(n8175), .ZN(n4733) );
  OR2_X1 U5352 ( .A1(n7297), .A2(n8154), .ZN(n4734) );
  AND2_X1 U5353 ( .A1(n8311), .A2(n8301), .ZN(n7031) );
  AND3_X1 U5354 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5802) );
  NAND2_X1 U5355 ( .A1(n7176), .A2(n8317), .ZN(n4746) );
  INV_X1 U5356 ( .A(n9125), .ZN(n9661) );
  OR2_X1 U5357 ( .A1(n8279), .A2(n6729), .ZN(n9662) );
  XNOR2_X1 U5358 ( .A(n6198), .B(n6197), .ZN(n6196) );
  NAND2_X1 U5359 ( .A1(n5742), .A2(n5745), .ZN(n4951) );
  NAND2_X1 U5360 ( .A1(n5596), .A2(n5595), .ZN(n5618) );
  XNOR2_X1 U5361 ( .A(n6080), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6090) );
  OAI21_X1 U5362 ( .B1(n6079), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6080) );
  AND2_X1 U5363 ( .A1(n5538), .A2(n5518), .ZN(n5534) );
  NAND2_X1 U5364 ( .A1(n4522), .A2(n4521), .ZN(n5716) );
  AND2_X1 U5365 ( .A1(n5703), .A2(n5724), .ZN(n4521) );
  NAND2_X1 U5366 ( .A1(n4576), .A2(n5464), .ZN(n5485) );
  NAND2_X1 U5367 ( .A1(n5441), .A2(n4580), .ZN(n4576) );
  NAND2_X1 U5368 ( .A1(n4862), .A2(n4984), .ZN(n5283) );
  XNOR2_X1 U5369 ( .A(n4985), .B(SI_5_), .ZN(n5282) );
  XNOR2_X1 U5370 ( .A(n4972), .B(SI_2_), .ZN(n5219) );
  AND2_X1 U5371 ( .A1(n5677), .A2(n5625), .ZN(n8666) );
  INV_X1 U5372 ( .A(n8787), .ZN(n8937) );
  INV_X1 U5373 ( .A(n8584), .ZN(n9752) );
  AND3_X1 U5374 ( .A1(n5529), .A2(n5528), .A3(n5527), .ZN(n8746) );
  AND4_X1 U5375 ( .A1(n5496), .A2(n5495), .A3(n5494), .A4(n5493), .ZN(n8562)
         );
  AND4_X1 U5376 ( .A1(n5455), .A2(n5454), .A3(n5453), .A4(n5452), .ZN(n8831)
         );
  OAI22_X1 U5377 ( .A1(n8138), .A2(n5221), .B1(n6204), .B2(n6203), .ZN(n8890)
         );
  INV_X1 U5378 ( .A(n8902), .ZN(n8668) );
  OAI211_X1 U5379 ( .C1(n8901), .C2(n9485), .A(n4426), .B(n4693), .ZN(n8982)
         );
  NAND2_X1 U5380 ( .A1(n8899), .A2(n9819), .ZN(n4693) );
  NAND2_X1 U5381 ( .A1(n8898), .A2(n9818), .ZN(n4692) );
  AND2_X1 U5382 ( .A1(n4935), .A2(n4461), .ZN(n4933) );
  AND2_X1 U5383 ( .A1(n4936), .A2(n9102), .ZN(n4935) );
  OAI21_X1 U5384 ( .B1(n8118), .B2(n4938), .A(n4937), .ZN(n4936) );
  NOR2_X1 U5385 ( .A1(n4943), .A2(n4939), .ZN(n4938) );
  NAND2_X1 U5386 ( .A1(n8118), .A2(n4942), .ZN(n4937) );
  NAND2_X1 U5387 ( .A1(n4941), .A2(n4942), .ZN(n4940) );
  INV_X1 U5388 ( .A(n8118), .ZN(n4941) );
  NAND2_X1 U5389 ( .A1(n6038), .A2(n6037), .ZN(n9383) );
  NAND2_X1 U5390 ( .A1(n9103), .A2(n8111), .ZN(n9001) );
  NAND2_X1 U5391 ( .A1(n8110), .A2(n8109), .ZN(n8111) );
  INV_X1 U5392 ( .A(n8107), .ZN(n8110) );
  NAND2_X1 U5393 ( .A1(n7665), .A2(n7664), .ZN(n7668) );
  INV_X1 U5394 ( .A(n9905), .ZN(n9269) );
  NAND2_X1 U5395 ( .A1(n5783), .A2(n5782), .ZN(n9688) );
  INV_X1 U5396 ( .A(n9333), .ZN(n9083) );
  INV_X1 U5397 ( .A(n9243), .ZN(n9268) );
  NAND2_X1 U5398 ( .A1(n4615), .A2(n4614), .ZN(n4613) );
  NAND2_X1 U5399 ( .A1(n8359), .A2(n4486), .ZN(n4615) );
  AOI21_X1 U5400 ( .B1(n8411), .B2(n4490), .A(n8417), .ZN(n4612) );
  NAND4_X1 U5401 ( .A1(n5788), .A2(n5787), .A3(n5786), .A4(n5785), .ZN(n9127)
         );
  OAI21_X1 U5402 ( .B1(n9182), .B2(n4572), .A(n4571), .ZN(n4570) );
  NAND2_X1 U5403 ( .A1(n6435), .A2(n6433), .ZN(n4572) );
  AOI21_X1 U5404 ( .B1(n9183), .B2(n9593), .A(n9585), .ZN(n4571) );
  NAND2_X1 U5405 ( .A1(n4569), .A2(n9185), .ZN(n4568) );
  OR2_X1 U5406 ( .A1(n9619), .A2(n9186), .ZN(n4569) );
  INV_X1 U5407 ( .A(n9194), .ZN(n9547) );
  AND2_X1 U5408 ( .A1(n4723), .A2(n4722), .ZN(n4721) );
  OR2_X1 U5409 ( .A1(n6071), .A2(n6072), .ZN(n4722) );
  OR2_X1 U5410 ( .A1(n9229), .A2(n9660), .ZN(n4723) );
  AOI21_X1 U5411 ( .B1(n9381), .B2(n9337), .A(n6154), .ZN(n6155) );
  OR2_X1 U5412 ( .A1(n5778), .A2(n6461), .ZN(n4815) );
  NAND2_X1 U5413 ( .A1(n4675), .A2(n5778), .ZN(n4674) );
  OAI21_X1 U5414 ( .B1(n9379), .B2(n9710), .A(n9382), .ZN(n4792) );
  NAND2_X1 U5415 ( .A1(n4384), .A2(n9635), .ZN(n4720) );
  INV_X1 U5416 ( .A(n4792), .ZN(n4962) );
  AND2_X1 U5417 ( .A1(n4721), .A2(n4469), .ZN(n4718) );
  NAND2_X1 U5418 ( .A1(n5713), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5707) );
  AOI21_X1 U5419 ( .B1(n4416), .B2(n8163), .A(n4606), .ZN(n4602) );
  NAND2_X1 U5420 ( .A1(n8249), .A2(n8326), .ZN(n4624) );
  AND2_X1 U5421 ( .A1(n4620), .A2(n4619), .ZN(n4618) );
  NAND2_X1 U5422 ( .A1(n4647), .A2(n4650), .ZN(n6325) );
  AOI21_X1 U5423 ( .B1(n4646), .B2(n4649), .A(n4406), .ZN(n4643) );
  INV_X1 U5424 ( .A(n8341), .ZN(n8147) );
  INV_X1 U5425 ( .A(n4659), .ZN(n4658) );
  AOI21_X1 U5426 ( .B1(n4659), .B2(n4657), .A(n8669), .ZN(n4656) );
  INV_X1 U5427 ( .A(n4661), .ZN(n4657) );
  NAND2_X1 U5428 ( .A1(n8897), .A2(n6362), .ZN(n4888) );
  INV_X1 U5429 ( .A(n7962), .ZN(n4930) );
  AND2_X1 U5430 ( .A1(n9393), .A2(n9228), .ZN(n8345) );
  NAND2_X1 U5431 ( .A1(n9408), .A2(n9269), .ZN(n8341) );
  AND2_X1 U5432 ( .A1(n9383), .A2(n9229), .ZN(n8225) );
  INV_X1 U5433 ( .A(n4578), .ZN(n4577) );
  OAI21_X1 U5434 ( .B1(n4580), .B2(n4579), .A(n5484), .ZN(n4578) );
  INV_X1 U5435 ( .A(n5464), .ZN(n4579) );
  NOR2_X1 U5436 ( .A1(n5168), .A2(n4833), .ZN(n4832) );
  INV_X1 U5437 ( .A(n5013), .ZN(n4833) );
  INV_X1 U5438 ( .A(n5009), .ZN(n4828) );
  AOI21_X1 U5439 ( .B1(n4832), .B2(n5014), .A(n4831), .ZN(n4830) );
  INV_X1 U5440 ( .A(n5020), .ZN(n4831) );
  OR2_X1 U5441 ( .A1(n8502), .A2(n8501), .ZN(n4845) );
  INV_X1 U5442 ( .A(n8704), .ZN(n4751) );
  OR2_X1 U5443 ( .A1(n5374), .A2(n5373), .ZN(n5393) );
  NOR2_X1 U5444 ( .A1(n7517), .A2(n4901), .ZN(n4900) );
  INV_X1 U5445 ( .A(n6271), .ZN(n4901) );
  NAND2_X1 U5446 ( .A1(n7230), .A2(n9746), .ZN(n7333) );
  AND2_X1 U5447 ( .A1(n5250), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5273) );
  AND2_X1 U5448 ( .A1(n7117), .A2(n9800), .ZN(n4698) );
  NAND2_X1 U5449 ( .A1(n8736), .A2(n4759), .ZN(n8727) );
  AND2_X1 U5450 ( .A1(n7407), .A2(n7252), .ZN(n6991) );
  NAND2_X1 U5451 ( .A1(n5170), .A2(n5058), .ZN(n5111) );
  INV_X1 U5452 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5045) );
  NOR2_X1 U5453 ( .A1(n7066), .A2(n4494), .ZN(n4493) );
  INV_X1 U5454 ( .A(n6938), .ZN(n4494) );
  AND2_X1 U5455 ( .A1(n6707), .A2(n6695), .ZN(n4512) );
  AND2_X1 U5456 ( .A1(n8100), .A2(n9080), .ZN(n4911) );
  NOR2_X1 U5457 ( .A1(n9054), .A2(n4519), .ZN(n4518) );
  INV_X1 U5458 ( .A(n9011), .ZN(n4519) );
  AND2_X1 U5459 ( .A1(n8100), .A2(n4923), .ZN(n4909) );
  INV_X1 U5460 ( .A(n8100), .ZN(n4908) );
  INV_X1 U5461 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5836) );
  INV_X1 U5462 ( .A(n8346), .ZN(n8351) );
  AND2_X1 U5463 ( .A1(n4799), .A2(n9227), .ZN(n4797) );
  NOR2_X1 U5464 ( .A1(n9393), .A2(n9228), .ZN(n8397) );
  OR2_X1 U5465 ( .A1(n6030), .A2(n9005), .ZN(n6039) );
  OR2_X1 U5466 ( .A1(n6021), .A2(n9109), .ZN(n6030) );
  OR2_X1 U5467 ( .A1(n9408), .A2(n9269), .ZN(n8388) );
  NOR2_X1 U5468 ( .A1(n4410), .A2(n4806), .ZN(n4805) );
  INV_X1 U5469 ( .A(n4812), .ZN(n4806) );
  NOR2_X1 U5470 ( .A1(n9549), .A2(n7908), .ZN(n4683) );
  NAND2_X1 U5471 ( .A1(n4732), .A2(n8154), .ZN(n4731) );
  NAND2_X1 U5472 ( .A1(n4688), .A2(n4403), .ZN(n7417) );
  NOR2_X1 U5473 ( .A1(n7430), .A2(n4686), .ZN(n4685) );
  NAND2_X1 U5474 ( .A1(n9563), .A2(n4687), .ZN(n4686) );
  AOI21_X1 U5475 ( .B1(n4599), .B2(n8318), .A(n6116), .ZN(n4596) );
  NAND2_X1 U5476 ( .A1(n5802), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5817) );
  AOI21_X1 U5477 ( .B1(n4744), .B2(n4743), .A(n6113), .ZN(n4742) );
  INV_X1 U5478 ( .A(n8317), .ZN(n4743) );
  NAND2_X1 U5479 ( .A1(n4744), .A2(n4601), .ZN(n4600) );
  INV_X1 U5480 ( .A(n7176), .ZN(n4601) );
  INV_X1 U5481 ( .A(n6691), .ZN(n6692) );
  AND2_X1 U5482 ( .A1(n9380), .A2(n8230), .ZN(n8363) );
  NAND2_X1 U5483 ( .A1(n7732), .A2(n4682), .ZN(n9365) );
  AND2_X1 U5484 ( .A1(n9371), .A2(n4400), .ZN(n4682) );
  AND2_X1 U5485 ( .A1(n5556), .A2(n5555), .ZN(n5557) );
  AND2_X1 U5486 ( .A1(n5440), .A2(n4581), .ZN(n4580) );
  INV_X1 U5487 ( .A(n5465), .ZN(n4581) );
  OR2_X1 U5488 ( .A1(n5109), .A2(n5039), .ZN(n5043) );
  INV_X1 U5489 ( .A(n5040), .ZN(n5041) );
  INV_X1 U5490 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n4510) );
  AND2_X1 U5491 ( .A1(n5025), .A2(n5024), .ZN(n5153) );
  INV_X1 U5492 ( .A(n5385), .ZN(n5014) );
  XNOR2_X1 U5493 ( .A(n5011), .B(SI_11_), .ZN(n5385) );
  NAND2_X1 U5494 ( .A1(n4448), .A2(n4485), .ZN(n5367) );
  NAND2_X1 U5495 ( .A1(n4995), .A2(n4768), .ZN(n4485) );
  NAND2_X1 U5496 ( .A1(n4768), .A2(n4770), .ZN(n4765) );
  AND2_X1 U5497 ( .A1(n5009), .A2(n5008), .ZN(n5366) );
  INV_X1 U5498 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5807) );
  INV_X1 U5499 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4966) );
  OR2_X1 U5500 ( .A1(n5182), .A2(n5181), .ZN(n7938) );
  OR2_X1 U5501 ( .A1(n5119), .A2(n9982), .ZN(n5426) );
  NAND2_X1 U5502 ( .A1(n5408), .A2(n4860), .ZN(n7879) );
  NAND2_X1 U5503 ( .A1(n5184), .A2(n7995), .ZN(n4860) );
  XNOR2_X1 U5504 ( .A(n5602), .B(n7117), .ZN(n8551) );
  INV_X1 U5505 ( .A(n5166), .ZN(n4858) );
  AND2_X1 U5506 ( .A1(n4853), .A2(n4456), .ZN(n4852) );
  NAND2_X1 U5507 ( .A1(n8486), .A2(n4849), .ZN(n4560) );
  AND2_X1 U5508 ( .A1(n6158), .A2(n6989), .ZN(n5224) );
  INV_X1 U5509 ( .A(n8024), .ZN(n5228) );
  NAND2_X1 U5510 ( .A1(n8502), .A2(n8501), .ZN(n4844) );
  AND2_X1 U5511 ( .A1(n7996), .A2(n7995), .ZN(n8516) );
  NAND2_X1 U5512 ( .A1(n4385), .A2(n6229), .ZN(n6372) );
  NOR2_X1 U5513 ( .A1(n8890), .A2(n6206), .ZN(n6371) );
  NAND2_X1 U5514 ( .A1(n4483), .A2(n6517), .ZN(n4669) );
  XNOR2_X1 U5515 ( .A(n6207), .B(n4385), .ZN(n4483) );
  NOR2_X1 U5516 ( .A1(n4889), .A2(n4886), .ZN(n4885) );
  AND4_X1 U5517 ( .A1(n5337), .A2(n5336), .A3(n5335), .A4(n5334), .ZN(n7330)
         );
  NAND2_X1 U5518 ( .A1(n6621), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4638) );
  NAND2_X1 U5519 ( .A1(n6883), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4634) );
  NOR2_X1 U5520 ( .A1(n6963), .A2(n4641), .ZN(n6965) );
  AND2_X1 U5521 ( .A1(n6964), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4641) );
  NOR2_X1 U5522 ( .A1(n6965), .A2(n6966), .ZN(n7077) );
  NOR2_X1 U5523 ( .A1(n7077), .A2(n4640), .ZN(n7081) );
  AND2_X1 U5524 ( .A1(n7078), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4640) );
  NAND2_X1 U5525 ( .A1(n7081), .A2(n7080), .ZN(n7239) );
  NOR2_X1 U5526 ( .A1(n8444), .A2(n8898), .ZN(n8656) );
  NAND2_X1 U5527 ( .A1(n8736), .A2(n4703), .ZN(n8444) );
  AND2_X1 U5528 ( .A1(n4401), .A2(n8668), .ZN(n4703) );
  AND2_X1 U5529 ( .A1(n5590), .A2(n5589), .ZN(n8687) );
  NAND2_X1 U5530 ( .A1(n8736), .A2(n4394), .ZN(n8711) );
  AND2_X1 U5531 ( .A1(n8736), .A2(n4401), .ZN(n8684) );
  INV_X1 U5532 ( .A(n4533), .ZN(n4532) );
  INV_X1 U5533 ( .A(n5545), .ZN(n5544) );
  INV_X1 U5534 ( .A(n8720), .ZN(n8724) );
  AND2_X1 U5535 ( .A1(n8756), .A2(n4761), .ZN(n8736) );
  NAND2_X1 U5536 ( .A1(n4877), .A2(n8761), .ZN(n4876) );
  NAND2_X1 U5537 ( .A1(n4878), .A2(n4412), .ZN(n4877) );
  NAND2_X1 U5538 ( .A1(n4958), .A2(n4777), .ZN(n4773) );
  INV_X1 U5539 ( .A(n4775), .ZN(n4774) );
  NOR3_X1 U5540 ( .A1(n8832), .A2(n8942), .A3(n8949), .ZN(n8797) );
  OR2_X1 U5541 ( .A1(n5450), .A2(n5449), .ZN(n5474) );
  OAI21_X1 U5542 ( .B1(n4867), .B2(n4866), .A(n4864), .ZN(n8821) );
  NAND2_X1 U5543 ( .A1(n6324), .A2(n4873), .ZN(n4866) );
  NAND2_X1 U5544 ( .A1(n4865), .A2(n6324), .ZN(n4864) );
  OR2_X1 U5545 ( .A1(n8844), .A2(n8953), .ZN(n8832) );
  NOR2_X1 U5546 ( .A1(n8832), .A2(n8949), .ZN(n8814) );
  NAND2_X1 U5547 ( .A1(n8826), .A2(n8436), .ZN(n4526) );
  AND2_X1 U5548 ( .A1(n7857), .A2(n4459), .ZN(n8843) );
  INV_X1 U5549 ( .A(n8522), .ZN(n4706) );
  OR2_X1 U5550 ( .A1(n8964), .A2(n8576), .ZN(n4788) );
  NAND2_X1 U5551 ( .A1(n7857), .A2(n4398), .ZN(n7987) );
  NAND2_X1 U5552 ( .A1(n7857), .A2(n4708), .ZN(n8867) );
  NAND2_X1 U5553 ( .A1(n7857), .A2(n7928), .ZN(n8865) );
  AND4_X1 U5554 ( .A1(n5178), .A2(n5177), .A3(n5176), .A4(n5175), .ZN(n7849)
         );
  NAND2_X1 U5555 ( .A1(n7591), .A2(n6287), .ZN(n4896) );
  AND2_X1 U5556 ( .A1(n7523), .A2(n4408), .ZN(n7867) );
  NAND2_X1 U5557 ( .A1(n7523), .A2(n4396), .ZN(n7868) );
  AND2_X1 U5558 ( .A1(n6562), .A2(n4749), .ZN(n5445) );
  INV_X1 U5559 ( .A(n6562), .ZN(n6518) );
  AND4_X1 U5560 ( .A1(n5357), .A2(n5356), .A3(n5355), .A4(n5354), .ZN(n7593)
         );
  AND2_X1 U5561 ( .A1(n7523), .A2(n9840), .ZN(n7525) );
  NAND2_X1 U5562 ( .A1(n7523), .A2(n4393), .ZN(n7596) );
  NAND2_X1 U5563 ( .A1(n6162), .A2(n6271), .ZN(n7516) );
  NOR2_X1 U5564 ( .A1(n4963), .A2(n7335), .ZN(n7523) );
  AND2_X1 U5565 ( .A1(n6270), .A2(n6271), .ZN(n7487) );
  AOI21_X1 U5566 ( .B1(n7324), .B2(n4524), .A(n4437), .ZN(n4523) );
  INV_X1 U5567 ( .A(n7324), .ZN(n4525) );
  OR2_X1 U5568 ( .A1(n7333), .A2(n7332), .ZN(n4963) );
  AND4_X1 U5569 ( .A1(n4698), .A2(n9811), .A3(n7008), .A4(n9830), .ZN(n7230)
         );
  AND2_X1 U5570 ( .A1(n7226), .A2(n6235), .ZN(n4899) );
  CLKBUF_X1 U5571 ( .A(n7001), .Z(n6980) );
  OR2_X1 U5572 ( .A1(n5349), .A2(n7097), .ZN(n5216) );
  NAND2_X1 U5573 ( .A1(n7676), .A2(n6188), .ZN(n5601) );
  INV_X1 U5574 ( .A(n7117), .ZN(n9817) );
  INV_X1 U5575 ( .A(n6991), .ZN(n9801) );
  AND2_X1 U5576 ( .A1(n5653), .A2(n5652), .ZN(n9791) );
  NAND3_X1 U5577 ( .A1(n5052), .A2(n4700), .A3(n10177), .ZN(n4902) );
  AND2_X1 U5578 ( .A1(n5298), .A2(n4903), .ZN(n4699) );
  NOR2_X1 U5579 ( .A1(n5060), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n4642) );
  INV_X1 U5580 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5044) );
  AND2_X1 U5581 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4967) );
  XNOR2_X1 U5582 ( .A(n6944), .B(n6738), .ZN(n7064) );
  INV_X1 U5584 ( .A(n4942), .ZN(n4939) );
  NAND2_X1 U5585 ( .A1(n4944), .A2(n9002), .ZN(n4943) );
  INV_X1 U5586 ( .A(n9003), .ZN(n4944) );
  XOR2_X1 U5587 ( .A(n8117), .B(n8116), .Z(n8118) );
  INV_X1 U5588 ( .A(n6764), .ZN(n6850) );
  NAND2_X1 U5589 ( .A1(n7282), .A2(n7283), .ZN(n4947) );
  OR2_X1 U5590 ( .A1(n7282), .A2(n7283), .ZN(n4948) );
  OR2_X1 U5591 ( .A1(n5853), .A2(n6598), .ZN(n5871) );
  NAND2_X1 U5592 ( .A1(n4500), .A2(n4499), .ZN(n8056) );
  AOI21_X1 U5593 ( .B1(n4501), .B2(n4504), .A(n4432), .ZN(n4499) );
  INV_X1 U5594 ( .A(n7956), .ZN(n4504) );
  INV_X1 U5595 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n10118) );
  NOR2_X1 U5596 ( .A1(n9595), .A2(n9594), .ZN(n9597) );
  NOR2_X1 U5597 ( .A1(n9597), .A2(n4564), .ZN(n9143) );
  AND2_X1 U5598 ( .A1(n6479), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4564) );
  NAND2_X1 U5599 ( .A1(n9143), .A2(n9144), .ZN(n9142) );
  NAND2_X1 U5600 ( .A1(n9142), .A2(n4563), .ZN(n9606) );
  OR2_X1 U5601 ( .A1(n9148), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4563) );
  NOR2_X1 U5602 ( .A1(n6599), .A2(n4463), .ZN(n6795) );
  NAND2_X1 U5603 ( .A1(n6795), .A2(n6794), .ZN(n6793) );
  NAND2_X1 U5604 ( .A1(n6793), .A2(n4561), .ZN(n6830) );
  OR2_X1 U5605 ( .A1(n6515), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4561) );
  XNOR2_X1 U5606 ( .A(n6406), .B(n6430), .ZN(n7214) );
  AND2_X1 U5607 ( .A1(n4566), .A2(n4565), .ZN(n7808) );
  NAND2_X1 U5608 ( .A1(n7805), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4565) );
  NOR2_X1 U5609 ( .A1(n7808), .A2(n7807), .ZN(n9162) );
  AND2_X1 U5610 ( .A1(n8281), .A2(n8349), .ZN(n9211) );
  AND2_X1 U5611 ( .A1(n9279), .A2(n4407), .ZN(n9221) );
  NAND2_X1 U5612 ( .A1(n9279), .A2(n4395), .ZN(n9235) );
  NAND2_X1 U5613 ( .A1(n9279), .A2(n6148), .ZN(n9270) );
  INV_X1 U5614 ( .A(n6002), .ZN(n6004) );
  AOI21_X1 U5615 ( .B1(n4820), .B2(n4817), .A(n4441), .ZN(n4816) );
  INV_X1 U5616 ( .A(n4820), .ZN(n4818) );
  NOR2_X1 U5617 ( .A1(n5967), .A2(n10029), .ZN(n5976) );
  OAI21_X1 U5618 ( .B1(n4714), .B2(n4712), .A(n8250), .ZN(n4711) );
  NOR2_X1 U5619 ( .A1(n9365), .A2(n9429), .ZN(n9349) );
  INV_X1 U5620 ( .A(n5957), .ZN(n5958) );
  NAND2_X1 U5621 ( .A1(n5958), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5967) );
  AND2_X1 U5622 ( .A1(n9510), .A2(n4728), .ZN(n4726) );
  NAND2_X1 U5623 ( .A1(n7732), .A2(n4683), .ZN(n9514) );
  AND2_X1 U5624 ( .A1(n9357), .A2(n8192), .ZN(n8270) );
  NOR2_X1 U5625 ( .A1(n5928), .A2(n10111), .ZN(n5936) );
  NAND2_X1 U5626 ( .A1(n7725), .A2(n8295), .ZN(n9501) );
  NAND2_X1 U5627 ( .A1(n4794), .A2(n8188), .ZN(n9512) );
  INV_X1 U5628 ( .A(n8188), .ZN(n9510) );
  NAND2_X1 U5629 ( .A1(n5902), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5918) );
  OR2_X1 U5630 ( .A1(n5918), .A2(n5917), .ZN(n5928) );
  NAND2_X1 U5631 ( .A1(n7732), .A2(n7918), .ZN(n9513) );
  NOR2_X1 U5632 ( .A1(n4727), .A2(n8171), .ZN(n7726) );
  INV_X1 U5633 ( .A(n7473), .ZN(n4727) );
  AND2_X1 U5634 ( .A1(n5892), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5902) );
  NAND2_X1 U5635 ( .A1(n4688), .A2(n4685), .ZN(n9536) );
  NOR2_X1 U5636 ( .A1(n5871), .A2(n5870), .ZN(n5881) );
  NOR3_X1 U5637 ( .A1(n7302), .A2(n7430), .A3(n9479), .ZN(n9537) );
  AND2_X1 U5638 ( .A1(n4734), .A2(n8303), .ZN(n7361) );
  NOR2_X1 U5639 ( .A1(n7302), .A2(n9479), .ZN(n7366) );
  AOI21_X1 U5640 ( .B1(n7124), .B2(n6120), .A(n4960), .ZN(n7301) );
  OR2_X1 U5641 ( .A1(n5851), .A2(n5850), .ZN(n5853) );
  AND2_X1 U5642 ( .A1(n7052), .A2(n7037), .ZN(n9627) );
  NAND2_X1 U5643 ( .A1(n4746), .A2(n4744), .ZN(n7023) );
  NOR2_X1 U5644 ( .A1(n9649), .A2(n7059), .ZN(n7052) );
  NAND2_X1 U5645 ( .A1(n4600), .A2(n4742), .ZN(n7047) );
  NAND2_X1 U5646 ( .A1(n7047), .A2(n7046), .ZN(n7045) );
  NAND2_X1 U5647 ( .A1(n9644), .A2(n6114), .ZN(n9646) );
  NOR2_X1 U5648 ( .A1(n7202), .A2(n7166), .ZN(n7183) );
  INV_X1 U5649 ( .A(n7159), .ZN(n8253) );
  AND2_X1 U5650 ( .A1(n5772), .A2(n5771), .ZN(n9066) );
  NOR2_X1 U5651 ( .A1(n5770), .A2(n5769), .ZN(n5771) );
  NOR2_X1 U5652 ( .A1(n6056), .A2(n5768), .ZN(n5769) );
  NOR2_X1 U5653 ( .A1(n6695), .A2(n7148), .ZN(n7144) );
  NAND2_X1 U5654 ( .A1(n6149), .A2(n6716), .ZN(n7126) );
  INV_X1 U5655 ( .A(n8236), .ZN(n9380) );
  NOR2_X1 U5656 ( .A1(n8280), .A2(n8363), .ZN(n8276) );
  INV_X1 U5657 ( .A(n7142), .ZN(n9671) );
  OR2_X1 U5658 ( .A1(n6717), .A2(n6716), .ZN(n9718) );
  INV_X1 U5659 ( .A(SI_30_), .ZN(n4479) );
  XNOR2_X1 U5660 ( .A(n6196), .B(SI_30_), .ZN(n8140) );
  XNOR2_X1 U5661 ( .A(n6183), .B(n6052), .ZN(n7797) );
  NAND2_X1 U5662 ( .A1(n5620), .A2(n5619), .ZN(n6047) );
  NAND2_X1 U5663 ( .A1(n5618), .A2(n5617), .ZN(n5620) );
  XNOR2_X1 U5664 ( .A(n5594), .B(n5593), .ZN(n7532) );
  XNOR2_X1 U5665 ( .A(n5563), .B(n5572), .ZN(n7535) );
  AND2_X1 U5666 ( .A1(n5559), .A2(n5571), .ZN(n5563) );
  OR2_X1 U5667 ( .A1(n5577), .A2(n5570), .ZN(n5559) );
  OR2_X1 U5668 ( .A1(n5577), .A2(n5554), .ZN(n5540) );
  NAND2_X1 U5669 ( .A1(n5441), .A2(n5440), .ZN(n5466) );
  XNOR2_X1 U5670 ( .A(n5100), .B(n5099), .ZN(n6841) );
  XNOR2_X1 U5671 ( .A(n5154), .B(n5153), .ZN(n6787) );
  INV_X1 U5672 ( .A(n4766), .ZN(n5359) );
  INV_X1 U5673 ( .A(n4771), .ZN(n4767) );
  NAND2_X1 U5674 ( .A1(n4995), .A2(n4994), .ZN(n5341) );
  XNOR2_X1 U5675 ( .A(n4988), .B(SI_6_), .ZN(n5300) );
  XNOR2_X1 U5676 ( .A(n4982), .B(SI_4_), .ZN(n5263) );
  NAND2_X1 U5677 ( .A1(n8135), .A2(n5309), .ZN(n7445) );
  NAND2_X1 U5678 ( .A1(n4836), .A2(n4834), .ZN(n8470) );
  AOI21_X1 U5679 ( .B1(n4837), .B2(n4840), .A(n4835), .ZN(n4834) );
  INV_X1 U5680 ( .A(n8460), .ZN(n4835) );
  AND4_X1 U5681 ( .A1(n5124), .A2(n5123), .A3(n5122), .A4(n5121), .ZN(n8883)
         );
  NAND2_X1 U5682 ( .A1(n5520), .A2(n5519), .ZN(n8927) );
  AND4_X1 U5683 ( .A1(n5400), .A2(n5399), .A3(n5398), .A4(n5397), .ZN(n7788)
         );
  NAND2_X1 U5684 ( .A1(n4543), .A2(n7544), .ZN(n7557) );
  NAND2_X1 U5685 ( .A1(n7377), .A2(n4548), .ZN(n4543) );
  INV_X1 U5686 ( .A(n5462), .ZN(n8489) );
  AND4_X1 U5687 ( .A1(n5317), .A2(n5316), .A3(n5315), .A4(n5314), .ZN(n8129)
         );
  OAI21_X1 U5688 ( .B1(n8560), .B2(n8559), .A(n4851), .ZN(n8495) );
  INV_X1 U5689 ( .A(n4854), .ZN(n4851) );
  AND2_X1 U5690 ( .A1(n5290), .A2(n5272), .ZN(n4558) );
  NAND2_X1 U5691 ( .A1(n8542), .A2(n5272), .ZN(n9745) );
  NAND2_X1 U5692 ( .A1(n7377), .A2(n5348), .ZN(n7545) );
  NAND2_X1 U5693 ( .A1(n8486), .A2(n5463), .ZN(n8560) );
  AND4_X1 U5694 ( .A1(n5147), .A2(n5146), .A3(n5145), .A4(n5144), .ZN(n7999)
         );
  INV_X1 U5695 ( .A(n4859), .ZN(n7828) );
  INV_X1 U5696 ( .A(n4545), .ZN(n4544) );
  OAI22_X1 U5697 ( .A1(n4546), .A2(n4548), .B1(n5383), .B2(n5384), .ZN(n4545)
         );
  INV_X1 U5698 ( .A(n6456), .ZN(n4554) );
  INV_X1 U5699 ( .A(n6455), .ZN(n4553) );
  NOR2_X1 U5700 ( .A1(n8461), .A2(n9743), .ZN(n4557) );
  NAND2_X1 U5701 ( .A1(n6452), .A2(n6453), .ZN(n4556) );
  NAND2_X1 U5702 ( .A1(n4843), .A2(n4844), .ZN(n6452) );
  NAND2_X1 U5703 ( .A1(n4669), .A2(n7451), .ZN(n4668) );
  AND4_X1 U5704 ( .A1(n5164), .A2(n5163), .A3(n5162), .A4(n5161), .ZN(n8881)
         );
  INV_X1 U5705 ( .A(n7593), .ZN(n8582) );
  INV_X1 U5706 ( .A(n8422), .ZN(n6209) );
  INV_X1 U5707 ( .A(n4627), .ZN(n6633) );
  NAND2_X1 U5708 ( .A1(n6568), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4626) );
  INV_X1 U5709 ( .A(n4639), .ZN(n6611) );
  INV_X1 U5710 ( .A(n4637), .ZN(n6809) );
  INV_X1 U5711 ( .A(n4635), .ZN(n6878) );
  XNOR2_X1 U5712 ( .A(n4628), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8647) );
  NAND2_X1 U5713 ( .A1(n4629), .A2(n8644), .ZN(n4628) );
  NAND2_X1 U5714 ( .A1(n8641), .A2(n8642), .ZN(n4629) );
  XNOR2_X1 U5715 ( .A(n8890), .B(n8893), .ZN(n8892) );
  INV_X1 U5716 ( .A(n8451), .ZN(n8452) );
  AOI22_X1 U5717 ( .A1(n8695), .A2(n9772), .B1(n8450), .B2(n8568), .ZN(n8451)
         );
  AOI21_X1 U5718 ( .B1(n8672), .B2(n9774), .A(n8708), .ZN(n8709) );
  OAI21_X1 U5719 ( .B1(n8753), .B2(n4537), .A(n4533), .ZN(n8699) );
  OAI21_X1 U5720 ( .B1(n8735), .B2(n4757), .A(n4753), .ZN(n8700) );
  NAND2_X1 U5721 ( .A1(n4752), .A2(n4756), .ZN(n8719) );
  NAND2_X1 U5722 ( .A1(n4755), .A2(n4760), .ZN(n8721) );
  NOR2_X1 U5723 ( .A1(n4882), .A2(n4880), .ZN(n8773) );
  NAND2_X1 U5724 ( .A1(n4879), .A2(n6333), .ZN(n8774) );
  AND2_X1 U5725 ( .A1(n5488), .A2(n5487), .ZN(n8787) );
  NAND2_X1 U5726 ( .A1(n8795), .A2(n4958), .ZN(n8781) );
  NAND2_X1 U5727 ( .A1(n4870), .A2(n4868), .ZN(n8828) );
  OAI21_X1 U5728 ( .B1(n7980), .B2(n6312), .A(n6315), .ZN(n8856) );
  INV_X1 U5729 ( .A(n8433), .ZN(n4782) );
  AND2_X1 U5730 ( .A1(n4529), .A2(n7838), .ZN(n7841) );
  INV_X1 U5731 ( .A(n4790), .ZN(n7864) );
  NAND2_X1 U5732 ( .A1(n7225), .A2(n7224), .ZN(n7325) );
  OR2_X1 U5733 ( .A1(n6203), .A2(n10132), .ZN(n5222) );
  INV_X1 U5734 ( .A(n8851), .ZN(n8872) );
  NAND2_X1 U5735 ( .A1(n9845), .A2(n5650), .ZN(n9778) );
  INV_X1 U5736 ( .A(n9792), .ZN(n9795) );
  NAND2_X1 U5737 ( .A1(n5071), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5073) );
  INV_X1 U5738 ( .A(n8714), .ZN(n8649) );
  INV_X1 U5739 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6493) );
  INV_X1 U5740 ( .A(n5056), .ZN(n5338) );
  INV_X1 U5741 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6488) );
  INV_X1 U5742 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6478) );
  INV_X1 U5743 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6470) );
  INV_X1 U5744 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6472) );
  NAND2_X1 U5745 ( .A1(n4449), .A2(n9765), .ZN(n4633) );
  INV_X1 U5746 ( .A(n9259), .ZN(n9228) );
  NAND2_X1 U5747 ( .A1(n7676), .A2(n8139), .ZN(n6029) );
  AND2_X1 U5748 ( .A1(n4915), .A2(n4914), .ZN(n9010) );
  NOR2_X1 U5749 ( .A1(n4399), .A2(n4424), .ZN(n4925) );
  NAND2_X1 U5750 ( .A1(n5975), .A2(n5974), .ZN(n9420) );
  NAND2_X1 U5751 ( .A1(n7957), .A2(n7956), .ZN(n4931) );
  CLKBUF_X1 U5752 ( .A(n6860), .Z(n6859) );
  AND2_X1 U5753 ( .A1(n4920), .A2(n4913), .ZN(n9053) );
  NAND2_X1 U5754 ( .A1(n4431), .A2(n9091), .ZN(n4926) );
  NOR2_X1 U5755 ( .A1(n7432), .A2(n4507), .ZN(n4506) );
  INV_X1 U5756 ( .A(n7425), .ZN(n4507) );
  OR2_X1 U5757 ( .A1(n6730), .A2(n6068), .ZN(n9110) );
  AOI21_X1 U5758 ( .B1(n9031), .B2(n9032), .A(n4464), .ZN(n9105) );
  AND2_X1 U5759 ( .A1(n6780), .A2(n6779), .ZN(n9108) );
  OR2_X1 U5760 ( .A1(n6730), .A2(n6729), .ZN(n9106) );
  NAND4_X1 U5761 ( .A1(n5796), .A2(n5795), .A3(n5794), .A4(n5793), .ZN(n9126)
         );
  INV_X1 U5762 ( .A(n9066), .ZN(n9128) );
  OR2_X1 U5763 ( .A1(n5784), .A2(n9729), .ZN(n5760) );
  OR2_X1 U5764 ( .A1(n6058), .A2(n7199), .ZN(n5757) );
  OR2_X1 U5765 ( .A1(n5791), .A2(n7150), .ZN(n5739) );
  NAND2_X1 U5766 ( .A1(n5789), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5738) );
  OR2_X1 U5767 ( .A1(n6058), .A2(n5734), .ZN(n5741) );
  NAND2_X1 U5768 ( .A1(n4588), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5889) );
  NOR2_X1 U5769 ( .A1(n7605), .A2(n7606), .ZN(n7609) );
  INV_X1 U5770 ( .A(n4566), .ZN(n7804) );
  NAND2_X1 U5771 ( .A1(n4798), .A2(n4799), .ZN(n9220) );
  NAND2_X1 U5772 ( .A1(n9249), .A2(n9257), .ZN(n4803) );
  NAND2_X1 U5773 ( .A1(n4735), .A2(n4737), .ZN(n9265) );
  NAND2_X1 U5774 ( .A1(n4740), .A2(n8203), .ZN(n9285) );
  OR2_X1 U5775 ( .A1(n9300), .A2(n8248), .ZN(n4740) );
  NAND2_X1 U5776 ( .A1(n4821), .A2(n4819), .ZN(n9292) );
  INV_X1 U5777 ( .A(n4822), .ZN(n4819) );
  NAND2_X1 U5778 ( .A1(n6137), .A2(n4824), .ZN(n4821) );
  AOI21_X1 U5779 ( .B1(n6137), .B2(n4961), .A(n4965), .ZN(n9307) );
  INV_X1 U5780 ( .A(n4709), .ZN(n9330) );
  AOI21_X1 U5781 ( .B1(n9345), .B2(n9339), .A(n4714), .ZN(n4709) );
  OAI21_X1 U5782 ( .B1(n9345), .B2(n5963), .A(n9339), .ZN(n9343) );
  NAND2_X1 U5783 ( .A1(n4811), .A2(n4809), .ZN(n9340) );
  NAND2_X1 U5784 ( .A1(n6133), .A2(n4812), .ZN(n4811) );
  NAND2_X1 U5785 ( .A1(n6133), .A2(n4957), .ZN(n9356) );
  NAND2_X1 U5786 ( .A1(n5901), .A2(n5900), .ZN(n7769) );
  NAND2_X1 U5787 ( .A1(n4734), .A2(n4732), .ZN(n9521) );
  NAND2_X1 U5788 ( .A1(n6118), .A2(n6117), .ZN(n9623) );
  NAND2_X1 U5789 ( .A1(n5801), .A2(n5800), .ZN(n9651) );
  NAND2_X1 U5790 ( .A1(n4746), .A2(n8256), .ZN(n9655) );
  INV_X1 U5791 ( .A(n9676), .ZN(n7205) );
  OR2_X1 U5792 ( .A1(n9705), .A2(n6104), .ZN(n9629) );
  AOI211_X1 U5793 ( .C1(n9689), .C2(n9547), .A(n9546), .B(n9545), .ZN(n9567)
         );
  OAI21_X1 U5794 ( .B1(n6196), .B2(n4479), .A(n6199), .ZN(n4478) );
  NOR2_X1 U5795 ( .A1(n4951), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n4949) );
  XNOR2_X1 U5796 ( .A(n6047), .B(n6046), .ZN(n8457) );
  XNOR2_X1 U5797 ( .A(n5618), .B(n5617), .ZN(n7676) );
  XNOR2_X1 U5798 ( .A(n4587), .B(n5534), .ZN(n7454) );
  OAI21_X1 U5799 ( .B1(n5577), .B2(n5535), .A(n5536), .ZN(n4587) );
  INV_X1 U5800 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6491) );
  INV_X1 U5801 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9973) );
  AND2_X1 U5802 ( .A1(n5781), .A2(n5798), .ZN(n9584) );
  INV_X1 U5803 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6466) );
  XNOR2_X1 U5804 ( .A(n5747), .B(n4562), .ZN(n6461) );
  NAND2_X1 U5805 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4562) );
  NOR2_X1 U5806 ( .A1(n7644), .A2(n10203), .ZN(n9903) );
  NAND2_X1 U5807 ( .A1(n4555), .A2(n4551), .ZN(P2_U3242) );
  NOR2_X1 U5808 ( .A1(n6457), .A2(n4552), .ZN(n4551) );
  NAND2_X1 U5809 ( .A1(n4557), .A2(n4556), .ZN(n4555) );
  NAND2_X1 U5810 ( .A1(n4554), .A2(n4553), .ZN(n4552) );
  NOR2_X1 U5811 ( .A1(n8905), .A2(n4388), .ZN(n8677) );
  NAND2_X1 U5812 ( .A1(n4691), .A2(n4690), .ZN(P2_U3549) );
  NAND2_X1 U5813 ( .A1(n9873), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n4690) );
  NAND2_X1 U5814 ( .A1(n8982), .A2(n9875), .ZN(n4691) );
  NAND2_X1 U5815 ( .A1(n4763), .A2(n4762), .ZN(P2_U3517) );
  NAND2_X1 U5816 ( .A1(n9859), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n4762) );
  NAND2_X1 U5817 ( .A1(n8982), .A2(n9861), .ZN(n4763) );
  NAND2_X1 U5818 ( .A1(n4935), .A2(n4940), .ZN(n4934) );
  NAND2_X1 U5819 ( .A1(n6743), .A2(n6742), .ZN(n6746) );
  NAND2_X1 U5820 ( .A1(n4611), .A2(n4610), .ZN(P1_U3240) );
  OR2_X1 U5821 ( .A1(n8416), .A2(n8415), .ZN(n4610) );
  NAND2_X1 U5822 ( .A1(n4573), .A2(n4567), .ZN(P1_U3260) );
  OR2_X1 U5823 ( .A1(n9184), .A2(n4486), .ZN(n4573) );
  AOI21_X1 U5824 ( .B1(n4570), .B2(n4486), .A(n4568), .ZN(n4567) );
  NAND2_X1 U5825 ( .A1(n4677), .A2(n4471), .ZN(P1_U3552) );
  OAI21_X1 U5826 ( .B1(n4678), .B2(n4792), .A(n9742), .ZN(n4677) );
  INV_X1 U5827 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n4676) );
  NAND2_X1 U5828 ( .A1(n4717), .A2(n4716), .ZN(n4719) );
  NAND2_X1 U5829 ( .A1(n4469), .A2(n9724), .ZN(n4716) );
  NAND2_X1 U5830 ( .A1(n4962), .A2(n4718), .ZN(n4717) );
  OAI21_X1 U5831 ( .B1(n7154), .B2(n8419), .A(n4488), .ZN(P1_U3333) );
  AND2_X1 U5832 ( .A1(n4735), .A2(n4411), .ZN(n4392) );
  AND2_X1 U5833 ( .A1(n9840), .A2(n7714), .ZN(n4393) );
  AND2_X1 U5834 ( .A1(n4759), .A2(n4705), .ZN(n4394) );
  AND2_X1 U5835 ( .A1(n4680), .A2(n9240), .ZN(n4395) );
  AND2_X1 U5836 ( .A1(n4393), .A2(n4702), .ZN(n4396) );
  AND3_X1 U5837 ( .A1(n5549), .A2(n5548), .A3(n5547), .ZN(n8505) );
  AND2_X1 U5838 ( .A1(n4905), .A2(n4671), .ZN(n4397) );
  AND2_X1 U5839 ( .A1(n4708), .A2(n4707), .ZN(n4398) );
  AND2_X1 U5840 ( .A1(n9072), .A2(n4927), .ZN(n4399) );
  INV_X1 U5841 ( .A(n8855), .ZN(n4784) );
  AND2_X1 U5842 ( .A1(n4683), .A2(n7888), .ZN(n4400) );
  AND2_X1 U5843 ( .A1(n4394), .A2(n4704), .ZN(n4401) );
  AND2_X1 U5844 ( .A1(n9300), .A2(n4447), .ZN(n4402) );
  AND2_X1 U5845 ( .A1(n4685), .A2(n4689), .ZN(n4403) );
  AND3_X1 U5846 ( .A1(n4462), .A2(n5051), .A3(n4903), .ZN(n4404) );
  OR2_X1 U5847 ( .A1(n6110), .A2(n7177), .ZN(n4405) );
  OR2_X1 U5848 ( .A1(n4652), .A2(n6172), .ZN(n4406) );
  AND2_X1 U5849 ( .A1(n4395), .A2(n4679), .ZN(n4407) );
  AND2_X1 U5850 ( .A1(n4396), .A2(n4701), .ZN(n4408) );
  NAND2_X1 U5851 ( .A1(n5565), .A2(n5564), .ZN(n8919) );
  INV_X1 U5852 ( .A(n8919), .ZN(n4759) );
  NAND2_X1 U5853 ( .A1(n4980), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4409) );
  XNOR2_X1 U5854 ( .A(n5707), .B(n5722), .ZN(n6149) );
  NOR2_X1 U5855 ( .A1(n6382), .A2(P2_U3152), .ZN(n6517) );
  NAND2_X2 U5856 ( .A1(n7125), .A2(n6691), .ZN(n6738) );
  NAND2_X2 U5857 ( .A1(n5736), .A2(n7799), .ZN(n6058) );
  NAND4_X1 U5858 ( .A1(n5753), .A2(n5752), .A3(n5751), .A4(n5750), .ZN(n6695)
         );
  NAND2_X2 U5859 ( .A1(n6562), .A2(n4980), .ZN(n5221) );
  NAND2_X1 U5860 ( .A1(n5737), .A2(n7799), .ZN(n6056) );
  INV_X1 U5861 ( .A(n4757), .ZN(n4756) );
  NAND2_X1 U5862 ( .A1(n4758), .A2(n8720), .ZN(n4757) );
  INV_X1 U5863 ( .A(n8942), .ZN(n8802) );
  NAND2_X1 U5864 ( .A1(n5471), .A2(n5470), .ZN(n8942) );
  NOR2_X1 U5865 ( .A1(n6135), .A2(n9363), .ZN(n4410) );
  AND2_X1 U5866 ( .A1(n4737), .A2(n4736), .ZN(n4411) );
  INV_X1 U5867 ( .A(n6374), .ZN(n4884) );
  INV_X1 U5868 ( .A(n7066), .ZN(n4498) );
  OR2_X1 U5869 ( .A1(n6175), .A2(n8788), .ZN(n4412) );
  AND3_X1 U5870 ( .A1(n5257), .A2(n5256), .A3(n5255), .ZN(n4413) );
  NAND2_X1 U5871 ( .A1(n6081), .A2(n6090), .ZN(n6773) );
  AND2_X1 U5872 ( .A1(n9471), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4414) );
  OR2_X1 U5873 ( .A1(n8902), .A2(n8442), .ZN(n6357) );
  NAND2_X1 U5874 ( .A1(n6309), .A2(n6308), .ZN(n6170) );
  NAND2_X1 U5875 ( .A1(n4926), .A2(n8067), .ZN(n9071) );
  NAND4_X1 U5876 ( .A1(n5190), .A2(n5189), .A3(n5188), .A4(n4538), .ZN(n6157)
         );
  NAND2_X1 U5877 ( .A1(n5447), .A2(n5446), .ZN(n8949) );
  INV_X1 U5878 ( .A(n8949), .ZN(n4696) );
  AND3_X1 U5879 ( .A1(n4511), .A2(n5697), .A3(n5696), .ZN(n4415) );
  AND2_X1 U5880 ( .A1(n4605), .A2(n8232), .ZN(n4416) );
  NAND2_X1 U5881 ( .A1(n5362), .A2(n5361), .ZN(n6163) );
  AND2_X1 U5882 ( .A1(n4803), .A2(n6144), .ZN(n4417) );
  NOR2_X1 U5883 ( .A1(n7706), .A2(n9525), .ZN(n4418) );
  NAND2_X1 U5884 ( .A1(n5935), .A2(n5934), .ZN(n9440) );
  INV_X1 U5885 ( .A(n8295), .ZN(n4725) );
  NAND2_X1 U5886 ( .A1(n5916), .A2(n5915), .ZN(n7908) );
  OR3_X1 U5887 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        n9765), .ZN(n4419) );
  AND2_X1 U5888 ( .A1(n6312), .A2(n6372), .ZN(n4420) );
  AND2_X1 U5889 ( .A1(n4635), .A2(n4634), .ZN(n4421) );
  INV_X1 U5890 ( .A(n8209), .ZN(n8396) );
  INV_X1 U5891 ( .A(n8093), .ZN(n4918) );
  NAND2_X1 U5892 ( .A1(n6001), .A2(n6000), .ZN(n9405) );
  INV_X1 U5893 ( .A(n8336), .ZN(n8248) );
  AND2_X1 U5894 ( .A1(n4627), .A2(n4626), .ZN(n4422) );
  NAND2_X1 U5895 ( .A1(n5056), .A2(n4383), .ZN(n5074) );
  NAND2_X1 U5896 ( .A1(n4907), .A2(n5191), .ZN(n5259) );
  NAND2_X1 U5897 ( .A1(n5298), .A2(n5045), .ZN(n5318) );
  AND2_X1 U5898 ( .A1(n8448), .A2(n6359), .ZN(n4423) );
  NAND2_X1 U5899 ( .A1(n6020), .A2(n6019), .ZN(n9393) );
  AND2_X1 U5900 ( .A1(n8074), .A2(n8073), .ZN(n4424) );
  AOI21_X1 U5901 ( .B1(n4771), .B2(n5000), .A(n4769), .ZN(n4768) );
  AND2_X1 U5902 ( .A1(n8448), .A2(n6357), .ZN(n4425) );
  INV_X1 U5903 ( .A(n4649), .ZN(n4648) );
  AND2_X1 U5904 ( .A1(n8900), .A2(n4692), .ZN(n4426) );
  NAND2_X1 U5905 ( .A1(n9279), .A2(n4680), .ZN(n4681) );
  INV_X1 U5906 ( .A(n6350), .ZN(n4664) );
  OR2_X1 U5907 ( .A1(n4696), .A2(n8831), .ZN(n4427) );
  OR2_X1 U5908 ( .A1(n5778), .A2(n6463), .ZN(n4428) );
  OR2_X1 U5909 ( .A1(n8932), .A2(n8572), .ZN(n6338) );
  NAND2_X1 U5910 ( .A1(n4623), .A2(n8193), .ZN(n4429) );
  AND2_X1 U5911 ( .A1(n4633), .A2(n4631), .ZN(n4430) );
  AND4_X1 U5912 ( .A1(n5217), .A2(n5216), .A3(n5215), .A4(n5214), .ZN(n6159)
         );
  AND2_X1 U5913 ( .A1(n9096), .A2(n4928), .ZN(n4431) );
  NOR2_X1 U5914 ( .A1(n8050), .A2(n8049), .ZN(n4432) );
  AND2_X1 U5915 ( .A1(n4830), .A2(n4827), .ZN(n4433) );
  NAND2_X1 U5916 ( .A1(n9698), .A2(n9126), .ZN(n8316) );
  AND2_X1 U5917 ( .A1(n7496), .A2(n6274), .ZN(n7575) );
  INV_X1 U5918 ( .A(n8343), .ZN(n4741) );
  AOI21_X1 U5919 ( .B1(n8140), .B2(n6188), .A(n6187), .ZN(n8897) );
  INV_X1 U5920 ( .A(n8897), .ZN(n4893) );
  NOR2_X1 U5921 ( .A1(n4912), .A2(n4908), .ZN(n4434) );
  AND2_X1 U5922 ( .A1(n6569), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4435) );
  INV_X1 U5923 ( .A(n6134), .ZN(n4814) );
  AND2_X1 U5924 ( .A1(n9435), .A2(n9346), .ZN(n6134) );
  OR2_X1 U5925 ( .A1(n9040), .A2(n8050), .ZN(n4436) );
  AND2_X1 U5926 ( .A1(n8547), .A2(n9746), .ZN(n4437) );
  NOR2_X1 U5927 ( .A1(n9388), .A2(n9244), .ZN(n4438) );
  AND2_X1 U5928 ( .A1(n8937), .A2(n8807), .ZN(n8437) );
  AND2_X1 U5929 ( .A1(n9072), .A2(n4928), .ZN(n4439) );
  NAND2_X1 U5930 ( .A1(n4699), .A2(n4383), .ZN(n4440) );
  NOR2_X1 U5931 ( .A1(n9413), .A2(n9287), .ZN(n4441) );
  NAND2_X1 U5932 ( .A1(n8204), .A2(n8203), .ZN(n4442) );
  NAND2_X1 U5933 ( .A1(n6357), .A2(n6358), .ZN(n8669) );
  AND2_X1 U5934 ( .A1(n8787), .A2(n4696), .ZN(n4444) );
  INV_X1 U5935 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4700) );
  NAND2_X1 U5936 ( .A1(n6353), .A2(n6354), .ZN(n8681) );
  INV_X1 U5937 ( .A(n8681), .ZN(n4663) );
  INV_X1 U5938 ( .A(n4958), .ZN(n4776) );
  NOR2_X1 U5939 ( .A1(n9240), .A2(n9228), .ZN(n4445) );
  AND2_X1 U5940 ( .A1(n4759), .A2(n8747), .ZN(n4446) );
  AND2_X1 U5941 ( .A1(n4739), .A2(n4741), .ZN(n4447) );
  AND2_X1 U5942 ( .A1(n4765), .A2(n5005), .ZN(n4448) );
  AND2_X1 U5943 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4449) );
  OR2_X1 U5944 ( .A1(n8953), .A2(n8573), .ZN(n4450) );
  OR2_X1 U5945 ( .A1(n9393), .A2(n9259), .ZN(n4451) );
  AND3_X1 U5946 ( .A1(n5387), .A2(n5368), .A3(n5057), .ZN(n4452) );
  AND2_X1 U5947 ( .A1(n4642), .A2(n5061), .ZN(n4453) );
  NAND2_X1 U5948 ( .A1(n8346), .A2(n8348), .ZN(n9227) );
  AND2_X1 U5949 ( .A1(n8259), .A2(n6117), .ZN(n4454) );
  AND2_X1 U5950 ( .A1(n5435), .A2(n5412), .ZN(n4455) );
  NOR2_X1 U5951 ( .A1(n8315), .A2(n4745), .ZN(n4744) );
  NAND2_X1 U5952 ( .A1(n5499), .A2(n5498), .ZN(n4456) );
  OR2_X1 U5953 ( .A1(n4495), .A2(n4493), .ZN(n4457) );
  AND2_X1 U5954 ( .A1(n7666), .A2(n7664), .ZN(n4458) );
  AND2_X1 U5955 ( .A1(n4398), .A2(n4706), .ZN(n4459) );
  AND2_X1 U5956 ( .A1(n4655), .A2(n4423), .ZN(n4460) );
  NAND2_X1 U5957 ( .A1(n5945), .A2(n5944), .ZN(n9435) );
  NAND2_X1 U5958 ( .A1(n8118), .A2(n4943), .ZN(n4461) );
  AND2_X1 U5959 ( .A1(n5052), .A2(n4700), .ZN(n4462) );
  XNOR2_X1 U5960 ( .A(n5073), .B(n5072), .ZN(n5632) );
  NAND2_X1 U5961 ( .A1(n5543), .A2(n5542), .ZN(n8922) );
  INV_X1 U5962 ( .A(n8922), .ZN(n4761) );
  NAND2_X1 U5963 ( .A1(n5778), .A2(n4980), .ZN(n5964) );
  NAND2_X1 U5964 ( .A1(n4931), .A2(n7962), .ZN(n8039) );
  NAND2_X1 U5965 ( .A1(n5697), .A2(n5696), .ZN(n5824) );
  NAND2_X1 U5966 ( .A1(n6123), .A2(n7360), .ZN(n7409) );
  INV_X1 U5967 ( .A(n6989), .ZN(n6894) );
  OR2_X1 U5968 ( .A1(n6383), .A2(n9801), .ZN(n6989) );
  AND2_X1 U5969 ( .A1(n6603), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4463) );
  OAI21_X1 U5970 ( .B1(n7409), .B2(n6124), .A(n6127), .ZN(n7475) );
  NAND2_X1 U5971 ( .A1(n4896), .A2(n6288), .ZN(n7872) );
  INV_X1 U5972 ( .A(n8803), .ZN(n4652) );
  NAND2_X1 U5973 ( .A1(n7903), .A2(n7902), .ZN(n7957) );
  INV_X1 U5974 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4904) );
  INV_X1 U5975 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n4671) );
  NAND2_X1 U5976 ( .A1(n5582), .A2(n5581), .ZN(n8914) );
  INV_X1 U5977 ( .A(n8914), .ZN(n4705) );
  NAND2_X1 U5978 ( .A1(n4508), .A2(n4506), .ZN(n7665) );
  NAND2_X1 U5979 ( .A1(n4508), .A2(n7425), .ZN(n7431) );
  NAND2_X1 U5980 ( .A1(n6029), .A2(n6028), .ZN(n9388) );
  INV_X1 U5981 ( .A(n9388), .ZN(n4679) );
  NOR3_X1 U5982 ( .A1(n8832), .A2(n8932), .A3(n4695), .ZN(n4697) );
  NAND2_X1 U5983 ( .A1(n5899), .A2(n5700), .ZN(n5924) );
  AND2_X1 U5984 ( .A1(n8105), .A2(n8104), .ZN(n4464) );
  NAND2_X1 U5985 ( .A1(n5601), .A2(n5600), .ZN(n8907) );
  INV_X1 U5986 ( .A(n8907), .ZN(n4704) );
  NAND2_X1 U5987 ( .A1(n7732), .A2(n4400), .ZN(n4684) );
  AND2_X1 U5988 ( .A1(n4870), .A2(n4869), .ZN(n4465) );
  NOR2_X1 U5989 ( .A1(n8914), .A2(n8569), .ZN(n4466) );
  INV_X1 U5990 ( .A(n4694), .ZN(n8782) );
  NOR2_X1 U5991 ( .A1(n8832), .A2(n4695), .ZN(n4694) );
  INV_X1 U5992 ( .A(n6149), .ZN(n6146) );
  AND2_X1 U5993 ( .A1(n5170), .A2(n4642), .ZN(n4467) );
  AND2_X1 U5994 ( .A1(n4785), .A2(n4782), .ZN(n4468) );
  INV_X1 U5995 ( .A(n8232), .ZN(n4608) );
  NAND2_X1 U5996 ( .A1(n5372), .A2(n5371), .ZN(n7779) );
  INV_X1 U5997 ( .A(n7779), .ZN(n4702) );
  OR2_X1 U5998 ( .A1(n9726), .A2(n6055), .ZN(n4469) );
  OR2_X1 U5999 ( .A1(n5641), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4470) );
  XNOR2_X1 U6000 ( .A(n5053), .B(n5078), .ZN(n5684) );
  OR2_X1 U6001 ( .A1(n9742), .A2(n4676), .ZN(n4471) );
  AND2_X1 U6002 ( .A1(n6925), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4472) );
  NAND2_X1 U6003 ( .A1(n5891), .A2(n5890), .ZN(n7706) );
  INV_X1 U6004 ( .A(n7706), .ZN(n4689) );
  NAND2_X1 U6005 ( .A1(n9646), .A2(n6115), .ZN(n7044) );
  NAND2_X1 U6006 ( .A1(n6939), .A2(n6938), .ZN(n7065) );
  INV_X1 U6007 ( .A(n8964), .ZN(n4707) );
  NAND2_X1 U6008 ( .A1(n4946), .A2(n4947), .ZN(n7285) );
  OR2_X1 U6009 ( .A1(n9626), .A2(n7315), .ZN(n7302) );
  INV_X1 U6010 ( .A(n7302), .ZN(n4688) );
  NAND2_X1 U6011 ( .A1(n4539), .A2(n4383), .ZN(n5641) );
  INV_X1 U6012 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8006) );
  AND2_X1 U6013 ( .A1(n4791), .A2(n4789), .ZN(n4473) );
  INV_X1 U6014 ( .A(n4487), .ZN(n6721) );
  NOR2_X1 U6015 ( .A1(n6717), .A2(n4490), .ZN(n4487) );
  NAND2_X1 U6016 ( .A1(n5839), .A2(n5838), .ZN(n9479) );
  INV_X1 U6017 ( .A(n9479), .ZN(n4687) );
  NAND2_X1 U6018 ( .A1(n5392), .A2(n5391), .ZN(n8975) );
  INV_X1 U6019 ( .A(n8975), .ZN(n4701) );
  OAI21_X1 U6020 ( .B1(n6845), .B2(n6844), .A(n6843), .ZN(n9060) );
  AND2_X1 U6021 ( .A1(n6989), .A2(n6983), .ZN(n4474) );
  NAND2_X1 U6022 ( .A1(n5714), .A2(n5713), .ZN(n7312) );
  INV_X1 U6023 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n10119) );
  NOR2_X1 U6024 ( .A1(n5081), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n8010) );
  INV_X1 U6025 ( .A(n5085), .ZN(n8430) );
  NOR2_X1 U6026 ( .A1(n8421), .A2(n7123), .ZN(n4489) );
  INV_X2 U6027 ( .A(n8008), .ZN(n8421) );
  NAND2_X1 U6028 ( .A1(n5301), .A2(n5300), .ZN(n4475) );
  NAND2_X1 U6029 ( .A1(n5283), .A2(n5282), .ZN(n4476) );
  INV_X2 U6030 ( .A(n4980), .ZN(n6051) );
  MUX2_X1 U6031 ( .A(n6466), .B(n6472), .S(n4980), .Z(n4976) );
  AND2_X4 U6032 ( .A1(n4481), .A2(n4480), .ZN(n4980) );
  OAI21_X2 U6033 ( .B1(n5502), .B2(n5501), .A(n5504), .ZN(n5577) );
  NAND2_X1 U6034 ( .A1(n6147), .A2(n8367), .ZN(n5718) );
  AOI21_X1 U6035 ( .B1(n6147), .B2(P1_STATE_REG_SCAN_IN), .A(n4489), .ZN(n4488) );
  AOI21_X1 U6036 ( .B1(n8358), .B2(n9350), .A(n4490), .ZN(n4614) );
  INV_X1 U6037 ( .A(n6147), .ZN(n4490) );
  NAND2_X1 U6038 ( .A1(n6939), .A2(n4457), .ZN(n4492) );
  NAND2_X1 U6039 ( .A1(n7903), .A2(n4501), .ZN(n4500) );
  NAND3_X1 U6040 ( .A1(n6743), .A2(n4505), .A3(n6742), .ZN(n6760) );
  INV_X1 U6041 ( .A(n6744), .ZN(n4505) );
  XNOR2_X1 U6042 ( .A(n6755), .B(n6756), .ZN(n6744) );
  NAND2_X1 U6043 ( .A1(n6760), .A2(n6759), .ZN(n6845) );
  NAND2_X1 U6044 ( .A1(n6700), .A2(n6699), .ZN(n6705) );
  NAND2_X1 U6045 ( .A1(n7126), .A2(n4512), .ZN(n4513) );
  INV_X1 U6046 ( .A(n6694), .ZN(n4514) );
  NAND2_X1 U6047 ( .A1(n6705), .A2(n6706), .ZN(n4515) );
  AND2_X1 U6048 ( .A1(n4514), .A2(n4513), .ZN(n6706) );
  AND2_X2 U6049 ( .A1(n7126), .A2(n6707), .ZN(n6764) );
  OAI21_X1 U6050 ( .B1(n8062), .B2(n6705), .A(n4515), .ZN(n6711) );
  NAND2_X1 U6051 ( .A1(n4517), .A2(n4516), .ZN(n9031) );
  NAND3_X1 U6052 ( .A1(n4915), .A2(n4518), .A3(n4914), .ZN(n4516) );
  NAND2_X1 U6053 ( .A1(n4520), .A2(n4910), .ZN(n4517) );
  NAND2_X1 U6054 ( .A1(n4919), .A2(n4916), .ZN(n4914) );
  NAND3_X1 U6055 ( .A1(n4915), .A2(n4914), .A3(n9011), .ZN(n4913) );
  AOI21_X1 U6056 ( .B1(n4919), .B2(n4909), .A(n4434), .ZN(n4520) );
  OAI21_X1 U6057 ( .B1(n7225), .B2(n4525), .A(n4523), .ZN(n9782) );
  NAND2_X1 U6058 ( .A1(n4527), .A2(n4791), .ZN(n4529) );
  AND2_X1 U6059 ( .A1(n4789), .A2(n7840), .ZN(n4527) );
  NAND2_X1 U6060 ( .A1(n4529), .A2(n4528), .ZN(n7929) );
  INV_X1 U6061 ( .A(n8753), .ZN(n4530) );
  OAI21_X1 U6062 ( .B1(n4530), .B2(n4532), .A(n4531), .ZN(n8682) );
  OR2_X1 U6063 ( .A1(n5349), .A2(n6987), .ZN(n4538) );
  INV_X1 U6064 ( .A(n6157), .ZN(n7002) );
  NAND2_X1 U6065 ( .A1(n7008), .A2(n6157), .ZN(n6245) );
  NOR2_X2 U6066 ( .A1(n5641), .A2(n4902), .ZN(n5079) );
  OR2_X2 U6067 ( .A1(n5261), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n4540) );
  NAND3_X1 U6068 ( .A1(n5191), .A2(n4907), .A3(n5044), .ZN(n5261) );
  XNOR2_X2 U6069 ( .A(n4542), .B(n5080), .ZN(n5085) );
  NOR2_X1 U6070 ( .A1(n8010), .A2(n8011), .ZN(n4542) );
  OAI21_X2 U6071 ( .B1(n7377), .B2(n4546), .A(n4544), .ZN(n7683) );
  NAND2_X1 U6072 ( .A1(n8135), .A2(n4550), .ZN(n7442) );
  NAND2_X1 U6073 ( .A1(n7442), .A2(n5329), .ZN(n5344) );
  NAND2_X1 U6074 ( .A1(n8542), .A2(n4558), .ZN(n9755) );
  NAND2_X1 U6075 ( .A1(n5170), .A2(n4453), .ZN(n5065) );
  NAND2_X1 U6076 ( .A1(n4583), .A2(n4582), .ZN(P1_U3355) );
  NAND2_X1 U6077 ( .A1(n4584), .A2(n9665), .ZN(n4583) );
  MUX2_X1 U6078 ( .A(n4981), .B(n6470), .S(n4980), .Z(n4982) );
  INV_X1 U6079 ( .A(n4415), .ZN(n4588) );
  NAND3_X1 U6080 ( .A1(n5727), .A2(n4415), .A3(n5730), .ZN(n5744) );
  NAND2_X1 U6081 ( .A1(n9129), .A2(n9676), .ZN(n8371) );
  AND2_X1 U6082 ( .A1(n4595), .A2(n4428), .ZN(n4594) );
  OR2_X1 U6083 ( .A1(n8137), .A2(n6474), .ZN(n4595) );
  INV_X1 U6084 ( .A(n7046), .ZN(n4599) );
  NAND2_X1 U6085 ( .A1(n4598), .A2(n4600), .ZN(n4597) );
  NAND2_X1 U6086 ( .A1(n8157), .A2(n4609), .ZN(n4603) );
  NAND2_X1 U6087 ( .A1(n8165), .A2(n4416), .ZN(n4604) );
  NAND3_X1 U6088 ( .A1(n4604), .A2(n4603), .A3(n4602), .ZN(n8179) );
  NAND2_X1 U6089 ( .A1(n8179), .A2(n8287), .ZN(n8172) );
  OAI21_X1 U6090 ( .B1(n8194), .B2(n4618), .A(n4616), .ZN(n8198) );
  AOI21_X1 U6091 ( .B1(n4621), .B2(n4429), .A(n4617), .ZN(n4616) );
  MUX2_X1 U6092 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6565), .S(n6579), .Z(n9457)
         );
  INV_X1 U6093 ( .A(n5065), .ZN(n5066) );
  NAND2_X1 U6094 ( .A1(n6311), .A2(n4648), .ZN(n4647) );
  OR2_X1 U6095 ( .A1(n6311), .A2(n4645), .ZN(n4644) );
  NAND2_X1 U6096 ( .A1(n4644), .A2(n4643), .ZN(n6327) );
  NAND3_X1 U6097 ( .A1(n7986), .A2(n4784), .A3(n6310), .ZN(n4649) );
  NAND2_X1 U6098 ( .A1(n4654), .A2(n4460), .ZN(n6364) );
  NAND2_X1 U6099 ( .A1(n6351), .A2(n4656), .ZN(n4654) );
  NAND2_X1 U6100 ( .A1(n4667), .A2(n4665), .ZN(P2_U3244) );
  INV_X1 U6101 ( .A(n4666), .ZN(n4665) );
  NAND2_X1 U6102 ( .A1(n6381), .A2(n4668), .ZN(n4667) );
  INV_X1 U6103 ( .A(n6385), .ZN(n4670) );
  OAI21_X1 U6104 ( .B1(n6467), .B2(n4980), .A(n4409), .ZN(n4675) );
  INV_X1 U6105 ( .A(n4681), .ZN(n9250) );
  INV_X1 U6106 ( .A(n4684), .ZN(n9364) );
  INV_X1 U6107 ( .A(n4697), .ZN(n8769) );
  NAND3_X1 U6108 ( .A1(n4698), .A2(n9811), .A3(n7008), .ZN(n7111) );
  NAND3_X1 U6109 ( .A1(n7008), .A2(n9811), .A3(n9800), .ZN(n7100) );
  NAND3_X1 U6110 ( .A1(n4383), .A2(n4404), .A3(n5298), .ZN(n5054) );
  OAI21_X2 U6111 ( .B1(n9345), .B2(n4713), .A(n4710), .ZN(n9315) );
  OAI21_X1 U6112 ( .B1(n4720), .B2(n9724), .A(n4719), .ZN(P1_U3520) );
  AOI211_X2 U6113 ( .C1(n7473), .C2(n4726), .A(n4724), .B(n8284), .ZN(n7892)
         );
  NAND2_X1 U6114 ( .A1(n7297), .A2(n4732), .ZN(n4730) );
  NAND2_X1 U6115 ( .A1(n4730), .A2(n4729), .ZN(n5888) );
  AND2_X1 U6116 ( .A1(n4731), .A2(n5887), .ZN(n4729) );
  NOR2_X1 U6117 ( .A1(n5999), .A2(n8247), .ZN(n4739) );
  NAND2_X1 U6118 ( .A1(n9300), .A2(n4739), .ZN(n4735) );
  XNOR2_X2 U6119 ( .A(n4747), .B(n5733), .ZN(n7799) );
  NAND2_X1 U6120 ( .A1(n4391), .A2(SI_0_), .ZN(n5755) );
  AOI21_X1 U6121 ( .B1(n4995), .B2(n4767), .A(n4770), .ZN(n4766) );
  AOI21_X1 U6122 ( .B1(n8768), .B2(n8775), .A(n8440), .ZN(n8755) );
  INV_X1 U6123 ( .A(n8437), .ZN(n4777) );
  INV_X1 U6124 ( .A(n5193), .ZN(n4778) );
  NAND2_X1 U6125 ( .A1(n4778), .A2(n4971), .ZN(n4779) );
  NAND2_X1 U6126 ( .A1(n4780), .A2(n4971), .ZN(n5220) );
  NAND2_X1 U6127 ( .A1(n5194), .A2(n5193), .ZN(n4780) );
  INV_X1 U6128 ( .A(n4971), .ZN(n4781) );
  NAND2_X1 U6129 ( .A1(n7984), .A2(n4786), .ZN(n4785) );
  NAND2_X1 U6130 ( .A1(n7984), .A2(n4788), .ZN(n7985) );
  INV_X1 U6131 ( .A(n4785), .ZN(n8434) );
  INV_X1 U6132 ( .A(n4788), .ZN(n4787) );
  NAND2_X1 U6133 ( .A1(n4790), .A2(n7873), .ZN(n4789) );
  NAND3_X1 U6134 ( .A1(n7782), .A2(n7778), .A3(n7873), .ZN(n4791) );
  NOR2_X2 U6135 ( .A1(n9199), .A2(n6145), .ZN(n4793) );
  INV_X1 U6136 ( .A(n9509), .ZN(n4794) );
  NAND2_X1 U6137 ( .A1(n6131), .A2(n6130), .ZN(n9509) );
  NAND2_X1 U6138 ( .A1(n9249), .A2(n4797), .ZN(n4796) );
  OAI21_X2 U6139 ( .B1(n6137), .B2(n4818), .A(n4816), .ZN(n9278) );
  INV_X1 U6140 ( .A(n9278), .ZN(n6141) );
  NAND2_X1 U6141 ( .A1(n6118), .A2(n4454), .ZN(n9625) );
  NAND2_X1 U6142 ( .A1(n9625), .A2(n6119), .ZN(n7124) );
  OAI22_X2 U6143 ( .A1(n7475), .A2(n6128), .B1(n7769), .B2(n9119), .ZN(n7724)
         );
  NAND3_X1 U6144 ( .A1(n4443), .A2(n4405), .A3(n6111), .ZN(n9644) );
  NAND2_X1 U6145 ( .A1(n5010), .A2(n5009), .ZN(n5386) );
  NAND2_X1 U6146 ( .A1(n8504), .A2(n4837), .ZN(n4836) );
  NAND2_X1 U6147 ( .A1(n8504), .A2(n4845), .ZN(n4843) );
  NAND3_X1 U6148 ( .A1(n5413), .A2(n5411), .A3(n4455), .ZN(n4846) );
  NAND2_X1 U6149 ( .A1(n4846), .A2(n4847), .ZN(n5462) );
  NAND3_X1 U6150 ( .A1(n5413), .A2(n5411), .A3(n5412), .ZN(n7950) );
  XNOR2_X1 U6151 ( .A(n5167), .B(n4858), .ZN(n4859) );
  INV_X1 U6152 ( .A(n5406), .ZN(n5182) );
  NAND2_X1 U6153 ( .A1(n5236), .A2(n4975), .ZN(n4863) );
  NAND3_X1 U6154 ( .A1(n5263), .A2(n4863), .A3(n4979), .ZN(n4862) );
  AND2_X1 U6155 ( .A1(n4863), .A2(n4979), .ZN(n5264) );
  INV_X1 U6156 ( .A(n7980), .ZN(n4867) );
  OAI21_X1 U6157 ( .B1(n8789), .B2(n4412), .A(n4878), .ZN(n8762) );
  INV_X1 U6158 ( .A(n4875), .ZN(n8760) );
  AOI21_X1 U6159 ( .B1(n8789), .B2(n4878), .A(n4876), .ZN(n4875) );
  INV_X1 U6160 ( .A(n4882), .ZN(n4879) );
  INV_X1 U6161 ( .A(n8775), .ZN(n4881) );
  NAND2_X1 U6162 ( .A1(n8670), .A2(n6356), .ZN(n4890) );
  AOI21_X1 U6163 ( .B1(n4890), .B2(n4885), .A(n4883), .ZN(n6207) );
  NOR2_X1 U6164 ( .A1(n8019), .A2(n7252), .ZN(n4892) );
  NAND2_X1 U6165 ( .A1(n4896), .A2(n4894), .ZN(n7784) );
  NAND2_X1 U6166 ( .A1(n7105), .A2(n6260), .ZN(n6161) );
  NAND2_X1 U6167 ( .A1(n6160), .A2(n4898), .ZN(n7105) );
  AND2_X1 U6168 ( .A1(n4899), .A2(n6236), .ZN(n4898) );
  NAND2_X1 U6169 ( .A1(n6236), .A2(n7226), .ZN(n7222) );
  NAND2_X1 U6170 ( .A1(n6160), .A2(n6235), .ZN(n7106) );
  NAND2_X1 U6171 ( .A1(n6162), .A2(n4900), .ZN(n7495) );
  NAND2_X1 U6172 ( .A1(n7495), .A2(n7496), .ZN(n6165) );
  NAND2_X1 U6173 ( .A1(n5079), .A2(n5078), .ZN(n5081) );
  NAND2_X1 U6174 ( .A1(n9077), .A2(n9080), .ZN(n4921) );
  NAND2_X1 U6175 ( .A1(n9077), .A2(n4911), .ZN(n4910) );
  NAND3_X1 U6176 ( .A1(n4921), .A2(n4922), .A3(n4918), .ZN(n4920) );
  INV_X1 U6177 ( .A(n8089), .ZN(n4919) );
  INV_X1 U6178 ( .A(n4922), .ZN(n9081) );
  NAND2_X1 U6179 ( .A1(n4924), .A2(n4925), .ZN(n9024) );
  NAND3_X1 U6180 ( .A1(n9091), .A2(n9096), .A3(n4439), .ZN(n4924) );
  NAND2_X1 U6181 ( .A1(n9091), .A2(n9096), .ZN(n9019) );
  INV_X1 U6182 ( .A(n8067), .ZN(n4927) );
  NAND2_X1 U6183 ( .A1(n9001), .A2(n4933), .ZN(n4932) );
  OAI211_X1 U6184 ( .C1(n9001), .C2(n4934), .A(n4932), .B(n8122), .ZN(P1_U3218) );
  NAND2_X1 U6185 ( .A1(n7665), .A2(n4458), .ZN(n7696) );
  NAND2_X1 U6186 ( .A1(n7284), .A2(n4948), .ZN(n4946) );
  NAND2_X1 U6187 ( .A1(n4950), .A2(n4949), .ZN(n8005) );
  INV_X1 U6188 ( .A(n5744), .ZN(n4950) );
  NAND2_X1 U6189 ( .A1(n9066), .A2(n7166), .ZN(n8319) );
  AOI211_X2 U6190 ( .C1(n8899), .C2(n8834), .A(n8455), .B(n8454), .ZN(n8456)
         );
  AND2_X1 U6191 ( .A1(n8423), .A2(n5207), .ZN(n6870) );
  NAND2_X1 U6192 ( .A1(n8706), .A2(n9777), .ZN(n8710) );
  XNOR2_X1 U6193 ( .A(n8705), .B(n8704), .ZN(n8706) );
  NAND2_X1 U6194 ( .A1(n8710), .A2(n8709), .ZN(n8912) );
  NAND2_X1 U6195 ( .A1(n5229), .A2(n5228), .ZN(n8022) );
  OAI21_X1 U6196 ( .B1(n5715), .B2(n5705), .A(n5704), .ZN(n5706) );
  NAND2_X2 U6197 ( .A1(n5085), .A2(n5083), .ZN(n5352) );
  CLKBUF_X1 U6198 ( .A(n9061), .Z(n9062) );
  OR2_X1 U6199 ( .A1(n5079), .A2(n8011), .ZN(n5053) );
  NAND2_X1 U6200 ( .A1(n5081), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5082) );
  XNOR2_X1 U6201 ( .A(n8449), .B(n8448), .ZN(n8453) );
  AND2_X1 U6202 ( .A1(n6109), .A2(n7173), .ZN(n4952) );
  AND2_X1 U6203 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n4953) );
  NAND2_X1 U6204 ( .A1(n6158), .A2(n9811), .ZN(n6244) );
  NOR2_X1 U6205 ( .A1(n5039), .A2(n5097), .ZN(n4954) );
  OR2_X1 U6206 ( .A1(n7928), .A2(n8881), .ZN(n4956) );
  OR2_X1 U6207 ( .A1(n8802), .A2(n8496), .ZN(n4958) );
  NOR2_X1 U6208 ( .A1(n6168), .A2(n7844), .ZN(n4959) );
  AND4_X1 U6209 ( .A1(n5096), .A2(n5095), .A3(n5094), .A4(n5093), .ZN(n8830)
         );
  INV_X1 U6210 ( .A(n9117), .ZN(n9229) );
  INV_X1 U6211 ( .A(n9774), .ZN(n8882) );
  CLKBUF_X3 U6212 ( .A(n6846), .Z(n8113) );
  AND2_X1 U6213 ( .A1(n5513), .A2(n5512), .ZN(n8572) );
  INV_X1 U6214 ( .A(n8572), .ZN(n8439) );
  AND2_X1 U6215 ( .A1(n7315), .A2(n9122), .ZN(n4960) );
  OR2_X1 U6216 ( .A1(n9423), .A2(n9347), .ZN(n4961) );
  OR2_X1 U6217 ( .A1(n7269), .A2(n7268), .ZN(n9873) );
  OR2_X1 U6218 ( .A1(n7269), .A2(n7261), .ZN(n9859) );
  AND2_X1 U6219 ( .A1(n8742), .A2(n8743), .ZN(n4964) );
  INV_X1 U6220 ( .A(n8261), .ZN(n6121) );
  AND2_X1 U6221 ( .A1(n9423), .A2(n9347), .ZN(n4965) );
  NAND2_X1 U6222 ( .A1(n7919), .A2(n7924), .ZN(n6168) );
  INV_X1 U6223 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5694) );
  AND2_X1 U6224 ( .A1(n4663), .A2(n8689), .ZN(n6176) );
  OAI21_X1 U6225 ( .B1(n6735), .B2(n7148), .A(n6697), .ZN(n6698) );
  INV_X1 U6226 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5701) );
  INV_X1 U6227 ( .A(n5393), .ZN(n5088) );
  OR2_X1 U6228 ( .A1(n5523), .A2(n5521), .ZN(n5545) );
  NAND2_X1 U6229 ( .A1(n8582), .A2(n7714), .ZN(n6280) );
  INV_X1 U6230 ( .A(n6773), .ZN(n6696) );
  INV_X1 U6231 ( .A(n5986), .ZN(n5985) );
  INV_X1 U6232 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5816) );
  INV_X1 U6233 ( .A(n8276), .ZN(n6063) );
  NAND2_X1 U6234 ( .A1(n9128), .A2(n9683), .ZN(n8313) );
  OR2_X1 U6235 ( .A1(n5572), .A2(n5571), .ZN(n5574) );
  INV_X1 U6236 ( .A(n5099), .ZN(n5039) );
  INV_X1 U6237 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5864) );
  INV_X1 U6238 ( .A(n7444), .ZN(n5328) );
  AND2_X1 U6239 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5250) );
  INV_X1 U6240 ( .A(n8488), .ZN(n5461) );
  INV_X1 U6241 ( .A(n6190), .ZN(n5249) );
  OR2_X1 U6242 ( .A1(n5349), .A2(n5198), .ZN(n5200) );
  INV_X1 U6243 ( .A(n7578), .ZN(n7579) );
  OR2_X1 U6244 ( .A1(n5331), .A2(n5330), .ZN(n5350) );
  NAND2_X1 U6245 ( .A1(n7002), .A2(n7098), .ZN(n6251) );
  NAND2_X1 U6246 ( .A1(n8671), .A2(n9774), .ZN(n8674) );
  INV_X1 U6247 ( .A(n8754), .ZN(n8761) );
  NAND2_X1 U6248 ( .A1(n8056), .A2(n8057), .ZN(n9092) );
  NAND2_X1 U6249 ( .A1(n5985), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6002) );
  OR2_X1 U6250 ( .A1(n6039), .A2(n8119), .ZN(n6151) );
  NAND2_X1 U6251 ( .A1(n5946), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5957) );
  NOR2_X1 U6252 ( .A1(n5817), .A2(n5816), .ZN(n5829) );
  OR2_X1 U6253 ( .A1(n9590), .A2(n9589), .ZN(n6426) );
  INV_X1 U6254 ( .A(n8225), .ZN(n8349) );
  NAND2_X1 U6255 ( .A1(n6004), .A2(n6003), .ZN(n6013) );
  NAND2_X1 U6256 ( .A1(P1_REG3_REG_21__SCAN_IN), .A2(n5976), .ZN(n5986) );
  OR2_X1 U6257 ( .A1(n9440), .A2(n9504), .ZN(n6132) );
  AND2_X1 U6258 ( .A1(n5881), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U6259 ( .A1(n7186), .A2(n9127), .ZN(n8317) );
  OR2_X1 U6260 ( .A1(n5558), .A2(n5557), .ZN(n5571) );
  NAND2_X1 U6261 ( .A1(n5716), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5717) );
  NOR2_X1 U6262 ( .A1(n4954), .A2(n5041), .ZN(n5042) );
  AND2_X1 U6263 ( .A1(n5616), .A2(n5615), .ZN(n8460) );
  OR2_X1 U6264 ( .A1(n5671), .A2(n5670), .ZN(n5672) );
  NAND2_X1 U6265 ( .A1(n5544), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U6266 ( .A1(n5157), .A2(n5156), .ZN(n6166) );
  INV_X1 U6267 ( .A(n9744), .ZN(n5290) );
  OR3_X1 U6268 ( .A1(n5583), .A2(n8507), .A3(n6454), .ZN(n5604) );
  OR2_X1 U6269 ( .A1(n6571), .A2(n8017), .ZN(n9761) );
  OAI22_X1 U6270 ( .A1(n8864), .A2(n8863), .B1(n9491), .B2(n8577), .ZN(n7930)
         );
  AND2_X1 U6271 ( .A1(n6976), .A2(n6243), .ZN(n6561) );
  NAND2_X1 U6272 ( .A1(n6245), .A2(n6251), .ZN(n7001) );
  NAND2_X1 U6273 ( .A1(n8674), .A2(n8673), .ZN(n8675) );
  AND2_X1 U6274 ( .A1(n6208), .A2(n6315), .ZN(n7986) );
  OR2_X1 U6275 ( .A1(n7576), .A2(n7575), .ZN(n7514) );
  AND2_X1 U6276 ( .A1(n5936), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5946) );
  OR2_X1 U6277 ( .A1(n6058), .A2(n5748), .ZN(n5753) );
  NAND2_X1 U6278 ( .A1(n6148), .A2(n9034), .ZN(n6142) );
  OR2_X1 U6279 ( .A1(n9429), .A2(n9332), .ZN(n6136) );
  INV_X1 U6280 ( .A(n8267), .ZN(n5908) );
  NAND2_X1 U6281 ( .A1(n9214), .A2(n9213), .ZN(n9215) );
  AND2_X1 U6282 ( .A1(n7022), .A2(n8322), .ZN(n7046) );
  AND2_X1 U6283 ( .A1(n6774), .A2(n6722), .ZN(n6726) );
  AND2_X1 U6284 ( .A1(n5040), .A2(n5038), .ZN(n5099) );
  AND2_X1 U6285 ( .A1(n5005), .A2(n5004), .ZN(n5358) );
  NAND2_X1 U6286 ( .A1(n4978), .A2(n4977), .ZN(n4979) );
  INV_X1 U6287 ( .A(n8554), .ZN(n9751) );
  INV_X1 U6288 ( .A(n9747), .ZN(n8565) );
  AND2_X1 U6289 ( .A1(n5610), .A2(n5609), .ZN(n8707) );
  AND4_X1 U6290 ( .A1(n5108), .A2(n5107), .A3(n5106), .A4(n5105), .ZN(n8858)
         );
  AND2_X1 U6291 ( .A1(n6577), .A2(n6576), .ZN(n9764) );
  NOR2_X1 U6292 ( .A1(n8900), .A2(n4388), .ZN(n8454) );
  INV_X1 U6293 ( .A(n8874), .ZN(n8834) );
  INV_X1 U6294 ( .A(n9819), .ZN(n9853) );
  AND2_X1 U6295 ( .A1(n7842), .A2(n9824), .ZN(n9485) );
  AND2_X1 U6296 ( .A1(n7514), .A2(n7513), .ZN(n9844) );
  OR3_X1 U6297 ( .A1(n7260), .A2(n7259), .A3(n7258), .ZN(n7269) );
  OAI21_X1 U6298 ( .B1(n7758), .B2(n7757), .A(n7756), .ZN(n7898) );
  AND2_X1 U6299 ( .A1(n6947), .A2(n9689), .ZN(n9100) );
  AND4_X1 U6300 ( .A1(n5992), .A2(n5991), .A3(n5990), .A4(n5989), .ZN(n9319)
         );
  INV_X1 U6301 ( .A(n9370), .ZN(n9531) );
  OR2_X1 U6302 ( .A1(n6717), .A2(n6147), .ZN(n9705) );
  AND2_X1 U6303 ( .A1(n9378), .A2(n9694), .ZN(n9710) );
  XNOR2_X1 U6304 ( .A(n4992), .B(SI_7_), .ZN(n5320) );
  XNOR2_X1 U6305 ( .A(n4976), .B(SI_3_), .ZN(n5237) );
  INV_X1 U6306 ( .A(n8655), .ZN(n9766) );
  INV_X1 U6307 ( .A(n8465), .ZN(n9750) );
  INV_X1 U6308 ( .A(n7330), .ZN(n8583) );
  INV_X1 U6309 ( .A(P2_U3966), .ZN(n8586) );
  AND2_X1 U6310 ( .A1(n6522), .A2(n6521), .ZN(n8655) );
  AND2_X1 U6311 ( .A1(n6382), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9798) );
  INV_X1 U6312 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10175) );
  INV_X1 U6313 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6477) );
  INV_X1 U6314 ( .A(n9393), .ZN(n9240) );
  OAI21_X1 U6315 ( .B1(n9379), .B2(n9374), .A(n6155), .ZN(n6156) );
  OR2_X1 U6316 ( .A1(n6543), .A2(n6718), .ZN(n9739) );
  OR2_X1 U6317 ( .A1(n6543), .A2(n6542), .ZN(n9724) );
  INV_X1 U6318 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10129) );
  INV_X1 U6319 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6481) );
  NOR2_X1 U6320 ( .A1(n9903), .A2(n9902), .ZN(n9901) );
  INV_X1 U6321 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6464) );
  INV_X1 U6322 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10132) );
  MUX2_X1 U6323 ( .A(n6464), .B(n10132), .S(n4980), .Z(n4972) );
  INV_X1 U6324 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5754) );
  NAND2_X1 U6325 ( .A1(n4980), .A2(n4967), .ZN(n5206) );
  NAND2_X1 U6326 ( .A1(n4968), .A2(n5206), .ZN(n4970) );
  INV_X1 U6327 ( .A(SI_1_), .ZN(n4969) );
  MUX2_X1 U6328 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4391), .Z(n5193) );
  NAND2_X1 U6329 ( .A1(n4970), .A2(SI_1_), .ZN(n4971) );
  INV_X1 U6330 ( .A(n4972), .ZN(n4973) );
  NAND2_X1 U6331 ( .A1(n4973), .A2(SI_2_), .ZN(n5235) );
  INV_X1 U6332 ( .A(n4976), .ZN(n4974) );
  NAND2_X1 U6333 ( .A1(n4974), .A2(SI_3_), .ZN(n4978) );
  AND2_X1 U6334 ( .A1(n5235), .A2(n4978), .ZN(n4975) );
  INV_X1 U6335 ( .A(n5237), .ZN(n4977) );
  INV_X1 U6336 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n4981) );
  INV_X1 U6337 ( .A(n4982), .ZN(n4983) );
  NAND2_X1 U6338 ( .A1(n4983), .A2(SI_4_), .ZN(n4984) );
  MUX2_X1 U6339 ( .A(n6477), .B(n9973), .S(n6051), .Z(n4985) );
  INV_X1 U6340 ( .A(n4985), .ZN(n4986) );
  NAND2_X1 U6341 ( .A1(n4986), .A2(SI_5_), .ZN(n4987) );
  MUX2_X1 U6342 ( .A(n6478), .B(n6481), .S(n6051), .Z(n4988) );
  INV_X1 U6343 ( .A(n4988), .ZN(n4989) );
  NAND2_X1 U6344 ( .A1(n4989), .A2(SI_6_), .ZN(n4990) );
  INV_X1 U6345 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n4991) );
  MUX2_X1 U6346 ( .A(n6488), .B(n4991), .S(n4749), .Z(n4992) );
  INV_X1 U6347 ( .A(n4992), .ZN(n4993) );
  NAND2_X1 U6348 ( .A1(n4993), .A2(SI_7_), .ZN(n4994) );
  MUX2_X1 U6349 ( .A(n6493), .B(n6491), .S(n6051), .Z(n4997) );
  INV_X1 U6350 ( .A(SI_8_), .ZN(n4996) );
  INV_X1 U6351 ( .A(n4997), .ZN(n4998) );
  NAND2_X1 U6352 ( .A1(n4998), .A2(SI_8_), .ZN(n4999) );
  INV_X1 U6353 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6495) );
  MUX2_X1 U6354 ( .A(n10175), .B(n6495), .S(n4749), .Z(n5002) );
  INV_X1 U6355 ( .A(SI_9_), .ZN(n5001) );
  INV_X1 U6356 ( .A(n5002), .ZN(n5003) );
  NAND2_X1 U6357 ( .A1(n5003), .A2(SI_9_), .ZN(n5004) );
  INV_X1 U6358 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6512) );
  INV_X1 U6359 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6509) );
  MUX2_X1 U6360 ( .A(n6512), .B(n6509), .S(n4749), .Z(n5006) );
  INV_X1 U6361 ( .A(SI_10_), .ZN(n9968) );
  NAND2_X1 U6362 ( .A1(n5006), .A2(n9968), .ZN(n5009) );
  INV_X1 U6363 ( .A(n5006), .ZN(n5007) );
  NAND2_X1 U6364 ( .A1(n5007), .A2(SI_10_), .ZN(n5008) );
  INV_X1 U6365 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6514) );
  MUX2_X1 U6366 ( .A(n6514), .B(n10129), .S(n4749), .Z(n5011) );
  INV_X1 U6367 ( .A(n5011), .ZN(n5012) );
  NAND2_X1 U6368 ( .A1(n5012), .A2(SI_11_), .ZN(n5013) );
  INV_X1 U6369 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5016) );
  INV_X1 U6370 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5015) );
  MUX2_X1 U6371 ( .A(n5016), .B(n5015), .S(n6051), .Z(n5017) );
  INV_X1 U6372 ( .A(SI_12_), .ZN(n9908) );
  NAND2_X1 U6373 ( .A1(n5017), .A2(n9908), .ZN(n5020) );
  INV_X1 U6374 ( .A(n5017), .ZN(n5018) );
  NAND2_X1 U6375 ( .A1(n5018), .A2(SI_12_), .ZN(n5019) );
  NAND2_X1 U6376 ( .A1(n5020), .A2(n5019), .ZN(n5168) );
  INV_X1 U6377 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6803) );
  INV_X1 U6378 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10178) );
  MUX2_X1 U6379 ( .A(n6803), .B(n10178), .S(n6051), .Z(n5022) );
  INV_X1 U6380 ( .A(SI_13_), .ZN(n5021) );
  NAND2_X1 U6381 ( .A1(n5022), .A2(n5021), .ZN(n5025) );
  INV_X1 U6382 ( .A(n5022), .ZN(n5023) );
  NAND2_X1 U6383 ( .A1(n5023), .A2(SI_13_), .ZN(n5024) );
  NAND2_X1 U6384 ( .A1(n5154), .A2(n5153), .ZN(n5026) );
  NAND2_X1 U6385 ( .A1(n5026), .A2(n5025), .ZN(n5134) );
  INV_X1 U6386 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6806) );
  INV_X1 U6387 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10160) );
  MUX2_X1 U6388 ( .A(n6806), .B(n10160), .S(n4749), .Z(n5027) );
  XNOR2_X1 U6389 ( .A(n5027), .B(SI_14_), .ZN(n5133) );
  INV_X1 U6390 ( .A(n5133), .ZN(n5030) );
  INV_X1 U6391 ( .A(n5027), .ZN(n5028) );
  NAND2_X1 U6392 ( .A1(n5028), .A2(SI_14_), .ZN(n5029) );
  INV_X1 U6393 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6838) );
  INV_X1 U6394 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6840) );
  MUX2_X1 U6395 ( .A(n6838), .B(n6840), .S(n6051), .Z(n5031) );
  INV_X1 U6396 ( .A(SI_15_), .ZN(n10137) );
  NAND2_X1 U6397 ( .A1(n5031), .A2(n10137), .ZN(n5097) );
  INV_X1 U6398 ( .A(n5031), .ZN(n5032) );
  NAND2_X1 U6399 ( .A1(n5032), .A2(SI_15_), .ZN(n5033) );
  NAND2_X1 U6400 ( .A1(n5097), .A2(n5033), .ZN(n5109) );
  INV_X1 U6401 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5034) );
  INV_X1 U6402 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6876) );
  MUX2_X1 U6403 ( .A(n5034), .B(n6876), .S(n6051), .Z(n5036) );
  INV_X1 U6404 ( .A(SI_16_), .ZN(n5035) );
  NAND2_X1 U6405 ( .A1(n5036), .A2(n5035), .ZN(n5040) );
  INV_X1 U6406 ( .A(n5036), .ZN(n5037) );
  NAND2_X1 U6407 ( .A1(n5037), .A2(SI_16_), .ZN(n5038) );
  INV_X1 U6408 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6930) );
  INV_X1 U6409 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10161) );
  MUX2_X1 U6410 ( .A(n6930), .B(n10161), .S(n6051), .Z(n5416) );
  XNOR2_X1 U6411 ( .A(n5416), .B(SI_17_), .ZN(n5415) );
  XNOR2_X1 U6412 ( .A(n5414), .B(n5415), .ZN(n6902) );
  INV_X1 U6413 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5068) );
  INV_X1 U6414 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5059) );
  INV_X1 U6415 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5057) );
  INV_X1 U6416 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5061) );
  NOR2_X1 U6417 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5048) );
  NOR2_X1 U6418 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5047) );
  NOR3_X1 U6419 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n5051) );
  INV_X1 U6420 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5052) );
  INV_X1 U6421 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5078) );
  INV_X1 U6422 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n10177) );
  NAND2_X1 U6423 ( .A1(n6902), .A2(n6188), .ZN(n5064) );
  INV_X1 U6424 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5058) );
  INV_X1 U6425 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5135) );
  NAND3_X1 U6426 ( .A1(n5112), .A2(n5135), .A3(n5059), .ZN(n5060) );
  NAND2_X1 U6427 ( .A1(n5065), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5062) );
  XNOR2_X1 U6428 ( .A(n5062), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8630) );
  AOI22_X1 U6429 ( .A1(n5445), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6518), .B2(
        n8630), .ZN(n5063) );
  INV_X1 U6430 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n10139) );
  NAND2_X1 U6431 ( .A1(n5066), .A2(n10139), .ZN(n5067) );
  NAND2_X1 U6432 ( .A1(n5419), .A2(n5068), .ZN(n5069) );
  INV_X1 U6433 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5070) );
  NAND2_X1 U6434 ( .A1(n5076), .A2(n5070), .ZN(n5071) );
  INV_X1 U6435 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5072) );
  NAND2_X1 U6436 ( .A1(n5074), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5075) );
  XNOR2_X1 U6437 ( .A(n5075), .B(n4904), .ZN(n7252) );
  INV_X1 U6438 ( .A(n7252), .ZN(n6243) );
  NAND2_X1 U6439 ( .A1(n4440), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5635) );
  INV_X1 U6440 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5634) );
  XNOR2_X1 U6441 ( .A(n5635), .B(n5634), .ZN(n7407) );
  INV_X1 U6442 ( .A(n7407), .ZN(n6976) );
  NAND2_X1 U6443 ( .A1(n4385), .A2(n6976), .ZN(n6982) );
  NAND3_X1 U6444 ( .A1(n6982), .A2(n7252), .A3(n9801), .ZN(n5077) );
  XNOR2_X1 U6445 ( .A(n8960), .B(n5602), .ZN(n5186) );
  INV_X1 U6446 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5080) );
  NAND2_X1 U6447 ( .A1(n6191), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5096) );
  AND2_X4 U6448 ( .A1(n8430), .A2(n5083), .ZN(n6190) );
  INV_X1 U6449 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n5084) );
  OR2_X1 U6450 ( .A1(n5249), .A2(n5084), .ZN(n5095) );
  NAND2_X1 U6451 ( .A1(n5273), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5311) );
  INV_X1 U6452 ( .A(n5311), .ZN(n5086) );
  NAND2_X1 U6453 ( .A1(n5086), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5331) );
  INV_X1 U6454 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5330) );
  INV_X1 U6455 ( .A(n5350), .ZN(n5087) );
  NAND2_X1 U6456 ( .A1(n5087), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5374) );
  INV_X1 U6457 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5373) );
  INV_X1 U6458 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5174) );
  INV_X1 U6459 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7243) );
  INV_X1 U6460 ( .A(n5159), .ZN(n5089) );
  NAND2_X1 U6461 ( .A1(n5089), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5143) );
  INV_X1 U6462 ( .A(n5143), .ZN(n5090) );
  NAND2_X1 U6463 ( .A1(n5090), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5119) );
  INV_X1 U6464 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9982) );
  INV_X1 U6465 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5425) );
  XNOR2_X1 U6466 ( .A(n5426), .B(n5425), .ZN(n8847) );
  OR2_X1 U6467 ( .A1(n5352), .A2(n8847), .ZN(n5094) );
  NAND2_X1 U6468 ( .A1(n8430), .A2(n5091), .ZN(n5213) );
  INV_X1 U6469 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n5092) );
  OR2_X1 U6470 ( .A1(n6195), .A2(n5092), .ZN(n5093) );
  NOR2_X1 U6471 ( .A1(n8830), .A2(n6894), .ZN(n5185) );
  XNOR2_X1 U6472 ( .A(n5186), .B(n5185), .ZN(n7881) );
  OR2_X1 U6473 ( .A1(n5110), .A2(n5109), .ZN(n5098) );
  NAND2_X1 U6474 ( .A1(n5098), .A2(n5097), .ZN(n5100) );
  NAND2_X1 U6475 ( .A1(n6841), .A2(n6188), .ZN(n5103) );
  OR2_X1 U6476 ( .A1(n4467), .A2(n8011), .ZN(n5101) );
  XNOR2_X1 U6477 ( .A(n5101), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8613) );
  AOI22_X1 U6478 ( .A1(n5445), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6518), .B2(
        n8613), .ZN(n5102) );
  XNOR2_X1 U6479 ( .A(n8522), .B(n5197), .ZN(n5125) );
  NAND2_X1 U6480 ( .A1(n6189), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5108) );
  INV_X1 U6481 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7989) );
  OR2_X1 U6482 ( .A1(n5349), .A2(n7989), .ZN(n5107) );
  INV_X1 U6483 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8591) );
  OR2_X1 U6484 ( .A1(n5249), .A2(n8591), .ZN(n5106) );
  NAND2_X1 U6485 ( .A1(n5119), .A2(n9982), .ZN(n5104) );
  NAND2_X1 U6486 ( .A1(n5426), .A2(n5104), .ZN(n8527) );
  OR2_X1 U6487 ( .A1(n5352), .A2(n8527), .ZN(n5105) );
  NOR2_X1 U6488 ( .A1(n8858), .A2(n6894), .ZN(n5126) );
  NAND2_X1 U6489 ( .A1(n5125), .A2(n5126), .ZN(n8515) );
  XNOR2_X1 U6490 ( .A(n5110), .B(n5109), .ZN(n6837) );
  NAND2_X1 U6491 ( .A1(n6837), .A2(n6188), .ZN(n5116) );
  NAND2_X1 U6492 ( .A1(n5111), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5155) );
  NAND2_X1 U6493 ( .A1(n5155), .A2(n5112), .ZN(n5113) );
  NAND2_X1 U6494 ( .A1(n5113), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5136) );
  NAND2_X1 U6495 ( .A1(n5136), .A2(n5135), .ZN(n5138) );
  NAND2_X1 U6496 ( .A1(n5138), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5114) );
  XNOR2_X1 U6497 ( .A(n5114), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8597) );
  AOI22_X1 U6498 ( .A1(n5445), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6518), .B2(
        n8597), .ZN(n5115) );
  XNOR2_X1 U6499 ( .A(n8964), .B(n5602), .ZN(n5131) );
  INV_X1 U6500 ( .A(n5131), .ZN(n8517) );
  NAND2_X1 U6501 ( .A1(n6190), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5124) );
  INV_X1 U6502 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5117) );
  NAND2_X1 U6503 ( .A1(n5143), .A2(n5117), .ZN(n5118) );
  NAND2_X1 U6504 ( .A1(n5119), .A2(n5118), .ZN(n8000) );
  OR2_X1 U6505 ( .A1(n5352), .A2(n8000), .ZN(n5123) );
  INV_X1 U6506 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n5120) );
  OR2_X1 U6507 ( .A1(n6195), .A2(n5120), .ZN(n5122) );
  INV_X1 U6508 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7932) );
  OR2_X1 U6509 ( .A1(n5349), .A2(n7932), .ZN(n5121) );
  NOR2_X1 U6510 ( .A1(n8883), .A2(n6894), .ZN(n5130) );
  INV_X1 U6511 ( .A(n5130), .ZN(n8518) );
  NAND3_X1 U6512 ( .A1(n8515), .A2(n8517), .A3(n8518), .ZN(n5129) );
  INV_X1 U6513 ( .A(n5125), .ZN(n5128) );
  INV_X1 U6514 ( .A(n5126), .ZN(n5127) );
  NAND2_X1 U6515 ( .A1(n5128), .A2(n5127), .ZN(n8514) );
  AND2_X1 U6516 ( .A1(n5129), .A2(n8514), .ZN(n5408) );
  NAND2_X1 U6517 ( .A1(n5131), .A2(n5130), .ZN(n5132) );
  AND2_X1 U6518 ( .A1(n8515), .A2(n5132), .ZN(n5184) );
  XNOR2_X1 U6519 ( .A(n5134), .B(n5133), .ZN(n6804) );
  NAND2_X1 U6520 ( .A1(n6804), .A2(n6188), .ZN(n5140) );
  OR2_X1 U6521 ( .A1(n5136), .A2(n5135), .ZN(n5137) );
  AND2_X1 U6522 ( .A1(n5138), .A2(n5137), .ZN(n7743) );
  AOI22_X1 U6523 ( .A1(n5445), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6518), .B2(
        n7743), .ZN(n5139) );
  XNOR2_X1 U6524 ( .A(n9491), .B(n5629), .ZN(n5148) );
  NAND2_X1 U6525 ( .A1(n6189), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5147) );
  INV_X1 U6526 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n5141) );
  OR2_X1 U6527 ( .A1(n5249), .A2(n5141), .ZN(n5146) );
  INV_X1 U6528 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9939) );
  NAND2_X1 U6529 ( .A1(n5159), .A2(n9939), .ZN(n5142) );
  NAND2_X1 U6530 ( .A1(n5143), .A2(n5142), .ZN(n8868) );
  OR2_X1 U6531 ( .A1(n5352), .A2(n8868), .ZN(n5145) );
  INV_X1 U6532 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8869) );
  OR2_X1 U6533 ( .A1(n5349), .A2(n8869), .ZN(n5144) );
  INV_X1 U6534 ( .A(n7999), .ZN(n8577) );
  NAND2_X1 U6535 ( .A1(n8577), .A2(n6989), .ZN(n5149) );
  NAND2_X1 U6536 ( .A1(n5148), .A2(n5149), .ZN(n5407) );
  INV_X1 U6537 ( .A(n5148), .ZN(n5151) );
  INV_X1 U6538 ( .A(n5149), .ZN(n5150) );
  NAND2_X1 U6539 ( .A1(n5151), .A2(n5150), .ZN(n5152) );
  NAND2_X1 U6540 ( .A1(n5407), .A2(n5152), .ZN(n7943) );
  INV_X1 U6541 ( .A(n7943), .ZN(n5183) );
  NAND2_X1 U6542 ( .A1(n6787), .A2(n6188), .ZN(n5157) );
  XNOR2_X1 U6543 ( .A(n5155), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7389) );
  AOI22_X1 U6544 ( .A1(n5445), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6518), .B2(
        n7389), .ZN(n5156) );
  INV_X1 U6545 ( .A(n5167), .ZN(n5165) );
  NAND2_X1 U6546 ( .A1(n6189), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5164) );
  INV_X1 U6547 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5158) );
  OR2_X1 U6548 ( .A1(n5249), .A2(n5158), .ZN(n5163) );
  OAI21_X1 U6549 ( .B1(n5395), .B2(n5174), .A(n7243), .ZN(n5160) );
  NAND2_X1 U6550 ( .A1(n5160), .A2(n5159), .ZN(n7854) );
  OR2_X1 U6551 ( .A1(n5352), .A2(n7854), .ZN(n5162) );
  INV_X1 U6552 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7855) );
  OR2_X1 U6553 ( .A1(n5349), .A2(n7855), .ZN(n5161) );
  NOR2_X1 U6554 ( .A1(n8881), .A2(n6894), .ZN(n5166) );
  NAND2_X1 U6555 ( .A1(n5165), .A2(n5166), .ZN(n5180) );
  XNOR2_X1 U6556 ( .A(n5169), .B(n5168), .ZN(n6528) );
  NAND2_X1 U6557 ( .A1(n6528), .A2(n6188), .ZN(n5173) );
  OR2_X1 U6558 ( .A1(n5170), .A2(n8011), .ZN(n5171) );
  XNOR2_X1 U6559 ( .A(n5171), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7240) );
  AOI22_X1 U6560 ( .A1(n5445), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6518), .B2(
        n7240), .ZN(n5172) );
  NAND2_X1 U6561 ( .A1(n5173), .A2(n5172), .ZN(n7837) );
  XNOR2_X1 U6562 ( .A(n7837), .B(n5197), .ZN(n5405) );
  NAND2_X1 U6563 ( .A1(n6189), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5178) );
  INV_X1 U6564 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7079) );
  OR2_X1 U6565 ( .A1(n5249), .A2(n7079), .ZN(n5177) );
  XNOR2_X1 U6566 ( .A(n5395), .B(n5174), .ZN(n7790) );
  OR2_X1 U6567 ( .A1(n5352), .A2(n7790), .ZN(n5176) );
  INV_X1 U6568 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7791) );
  OR2_X1 U6569 ( .A1(n5349), .A2(n7791), .ZN(n5175) );
  INV_X1 U6570 ( .A(n7849), .ZN(n8579) );
  NAND2_X1 U6571 ( .A1(n8579), .A2(n6989), .ZN(n5404) );
  INV_X1 U6572 ( .A(n5404), .ZN(n5179) );
  NAND2_X1 U6573 ( .A1(n5405), .A2(n5179), .ZN(n7826) );
  AND2_X1 U6574 ( .A1(n7826), .A2(n5180), .ZN(n5181) );
  OR2_X1 U6575 ( .A1(n7881), .A2(n7879), .ZN(n5413) );
  NAND2_X1 U6576 ( .A1(n5186), .A2(n5185), .ZN(n5412) );
  NAND2_X1 U6577 ( .A1(n6190), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5190) );
  INV_X1 U6578 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5187) );
  OR2_X1 U6579 ( .A1(n5213), .A2(n5187), .ZN(n5189) );
  INV_X1 U6580 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6871) );
  OR2_X1 U6581 ( .A1(n5352), .A2(n6871), .ZN(n5188) );
  INV_X1 U6582 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6987) );
  NAND2_X1 U6583 ( .A1(n6157), .A2(n6989), .ZN(n5210) );
  INV_X1 U6584 ( .A(n5191), .ZN(n5192) );
  XNOR2_X1 U6585 ( .A(n5194), .B(n5193), .ZN(n6467) );
  OR2_X1 U6586 ( .A1(n5221), .A2(n6467), .ZN(n5196) );
  NAND2_X4 U6587 ( .A1(n6562), .A2(n4749), .ZN(n6203) );
  INV_X1 U6588 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6468) );
  XNOR2_X1 U6589 ( .A(n5197), .B(n7098), .ZN(n5208) );
  XNOR2_X1 U6590 ( .A(n5210), .B(n5208), .ZN(n6869) );
  INV_X1 U6591 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7018) );
  OR2_X1 U6592 ( .A1(n5352), .A2(n7018), .ZN(n5202) );
  NAND2_X1 U6593 ( .A1(n6190), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5201) );
  INV_X1 U6594 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U6595 ( .A1(n6189), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5199) );
  INV_X1 U6596 ( .A(SI_0_), .ZN(n5204) );
  INV_X1 U6597 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5203) );
  OAI21_X1 U6598 ( .B1(n6051), .B2(n5204), .A(n5203), .ZN(n5205) );
  AND2_X1 U6599 ( .A1(n5206), .A2(n5205), .ZN(n9000) );
  MUX2_X1 U6600 ( .A(n9765), .B(n9000), .S(n6562), .Z(n8426) );
  NAND2_X1 U6601 ( .A1(n6209), .A2(n8426), .ZN(n7000) );
  INV_X1 U6602 ( .A(n7000), .ZN(n6974) );
  NAND2_X1 U6603 ( .A1(n6974), .A2(n6989), .ZN(n8423) );
  OR2_X1 U6604 ( .A1(n5197), .A2(n8426), .ZN(n5207) );
  NAND2_X1 U6605 ( .A1(n6869), .A2(n6870), .ZN(n6868) );
  INV_X1 U6606 ( .A(n5208), .ZN(n5209) );
  NAND2_X1 U6607 ( .A1(n5210), .A2(n5209), .ZN(n5211) );
  NAND2_X1 U6608 ( .A1(n6868), .A2(n5211), .ZN(n8025) );
  INV_X1 U6609 ( .A(n8025), .ZN(n5229) );
  NAND2_X1 U6610 ( .A1(n6190), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5217) );
  INV_X1 U6611 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7097) );
  INV_X1 U6612 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5212) );
  OR2_X1 U6613 ( .A1(n5213), .A2(n5212), .ZN(n5215) );
  INV_X1 U6614 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n8026) );
  OR2_X1 U6615 ( .A1(n5352), .A2(n8026), .ZN(n5214) );
  OR2_X1 U6616 ( .A1(n5191), .A2(n8011), .ZN(n5218) );
  XNOR2_X1 U6617 ( .A(n5218), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9471) );
  INV_X1 U6618 ( .A(n9471), .ZN(n6473) );
  XNOR2_X1 U6619 ( .A(n5220), .B(n5219), .ZN(n6474) );
  OR2_X1 U6620 ( .A1(n5221), .A2(n6474), .ZN(n5223) );
  XNOR2_X1 U6621 ( .A(n7102), .B(n5197), .ZN(n5225) );
  NAND2_X1 U6622 ( .A1(n5224), .A2(n5225), .ZN(n5230) );
  INV_X1 U6623 ( .A(n5224), .ZN(n5226) );
  INV_X1 U6624 ( .A(n5225), .ZN(n6895) );
  NAND2_X1 U6625 ( .A1(n5226), .A2(n6895), .ZN(n5227) );
  NAND2_X1 U6626 ( .A1(n5230), .A2(n5227), .ZN(n8024) );
  NAND2_X1 U6627 ( .A1(n8022), .A2(n5230), .ZN(n5248) );
  OR2_X1 U6628 ( .A1(n5352), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5234) );
  NAND2_X1 U6629 ( .A1(n6190), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5233) );
  INV_X1 U6630 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6999) );
  OR2_X1 U6631 ( .A1(n5349), .A2(n6999), .ZN(n5232) );
  NAND2_X1 U6632 ( .A1(n6189), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5231) );
  AND2_X1 U6633 ( .A1(n8585), .A2(n6989), .ZN(n5245) );
  NAND2_X1 U6634 ( .A1(n5236), .A2(n5235), .ZN(n5238) );
  XNOR2_X1 U6635 ( .A(n5238), .B(n5237), .ZN(n6471) );
  OR2_X1 U6636 ( .A1(n5221), .A2(n6471), .ZN(n5243) );
  OR2_X1 U6637 ( .A1(n6203), .A2(n6472), .ZN(n5242) );
  INV_X1 U6638 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5240) );
  NAND2_X1 U6639 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4419), .ZN(n5239) );
  XNOR2_X1 U6640 ( .A(n5240), .B(n5239), .ZN(n6643) );
  OR2_X1 U6641 ( .A1(n6562), .A2(n6643), .ZN(n5241) );
  NAND2_X1 U6642 ( .A1(n5245), .A2(n5244), .ZN(n5267) );
  INV_X1 U6643 ( .A(n5245), .ZN(n5246) );
  AND2_X1 U6644 ( .A1(n5267), .A2(n5247), .ZN(n6892) );
  NAND2_X1 U6645 ( .A1(n5248), .A2(n6892), .ZN(n8543) );
  INV_X1 U6646 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6564) );
  OR2_X1 U6647 ( .A1(n5249), .A2(n6564), .ZN(n5257) );
  INV_X1 U6648 ( .A(n5250), .ZN(n5274) );
  INV_X1 U6649 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5252) );
  INV_X1 U6650 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5251) );
  NAND2_X1 U6651 ( .A1(n5252), .A2(n5251), .ZN(n5253) );
  NAND2_X1 U6652 ( .A1(n5274), .A2(n5253), .ZN(n8546) );
  OR2_X1 U6653 ( .A1(n5352), .A2(n8546), .ZN(n5256) );
  INV_X1 U6654 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5254) );
  OR2_X1 U6655 ( .A1(n5213), .A2(n5254), .ZN(n5255) );
  NAND2_X1 U6656 ( .A1(n6191), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5258) );
  NAND2_X1 U6657 ( .A1(n8584), .A2(n6989), .ZN(n5271) );
  NAND2_X1 U6658 ( .A1(n5259), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5260) );
  MUX2_X1 U6659 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5260), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5262) );
  NAND2_X1 U6660 ( .A1(n5262), .A2(n5261), .ZN(n6676) );
  XNOR2_X1 U6661 ( .A(n5264), .B(n5263), .ZN(n6469) );
  OR2_X1 U6662 ( .A1(n5221), .A2(n6469), .ZN(n5266) );
  OR2_X1 U6663 ( .A1(n6203), .A2(n6470), .ZN(n5265) );
  OAI211_X1 U6664 ( .C1(n6562), .C2(n6676), .A(n5266), .B(n5265), .ZN(n8550)
         );
  XNOR2_X1 U6665 ( .A(n5602), .B(n8550), .ZN(n5269) );
  XNOR2_X1 U6666 ( .A(n5271), .B(n5269), .ZN(n8553) );
  AND2_X1 U6667 ( .A1(n8553), .A2(n5267), .ZN(n5268) );
  INV_X1 U6668 ( .A(n5269), .ZN(n5270) );
  NAND2_X1 U6669 ( .A1(n5271), .A2(n5270), .ZN(n5272) );
  NAND2_X1 U6670 ( .A1(n6190), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5280) );
  INV_X1 U6671 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7229) );
  OR2_X1 U6672 ( .A1(n5349), .A2(n7229), .ZN(n5279) );
  INV_X1 U6673 ( .A(n5273), .ZN(n5292) );
  INV_X1 U6674 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10169) );
  NAND2_X1 U6675 ( .A1(n5274), .A2(n10169), .ZN(n5275) );
  NAND2_X1 U6676 ( .A1(n5292), .A2(n5275), .ZN(n9758) );
  OR2_X1 U6677 ( .A1(n5352), .A2(n9758), .ZN(n5278) );
  INV_X1 U6678 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5276) );
  OR2_X1 U6679 ( .A1(n6195), .A2(n5276), .ZN(n5277) );
  NOR2_X1 U6680 ( .A1(n8547), .A2(n6894), .ZN(n5286) );
  NAND2_X1 U6681 ( .A1(n5261), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5281) );
  XNOR2_X1 U6682 ( .A(n5281), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6621) );
  INV_X1 U6683 ( .A(n6621), .ZN(n6585) );
  XNOR2_X1 U6684 ( .A(n5283), .B(n5282), .ZN(n6476) );
  OR2_X1 U6685 ( .A1(n5221), .A2(n6476), .ZN(n5285) );
  OR2_X1 U6686 ( .A1(n6203), .A2(n6477), .ZN(n5284) );
  OAI211_X1 U6687 ( .C1(n6562), .C2(n6585), .A(n5285), .B(n5284), .ZN(n7263)
         );
  XNOR2_X1 U6688 ( .A(n5602), .B(n7263), .ZN(n8123) );
  NAND2_X1 U6689 ( .A1(n5286), .A2(n8123), .ZN(n5304) );
  INV_X1 U6690 ( .A(n5286), .ZN(n5288) );
  INV_X1 U6691 ( .A(n8123), .ZN(n5287) );
  NAND2_X1 U6692 ( .A1(n5288), .A2(n5287), .ZN(n5289) );
  NAND2_X1 U6693 ( .A1(n5304), .A2(n5289), .ZN(n9744) );
  INV_X1 U6694 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U6695 ( .A1(n5292), .A2(n5291), .ZN(n5293) );
  NAND2_X1 U6696 ( .A1(n5311), .A2(n5293), .ZN(n9779) );
  OR2_X1 U6697 ( .A1(n5352), .A2(n9779), .ZN(n5297) );
  NAND2_X1 U6698 ( .A1(n6190), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5296) );
  INV_X1 U6699 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6620) );
  OR2_X1 U6700 ( .A1(n5349), .A2(n6620), .ZN(n5295) );
  NAND2_X1 U6701 ( .A1(n6189), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5294) );
  NAND4_X1 U6702 ( .A1(n5297), .A2(n5296), .A3(n5295), .A4(n5294), .ZN(n9748)
         );
  NAND2_X1 U6703 ( .A1(n9748), .A2(n6989), .ZN(n5307) );
  OR2_X1 U6704 ( .A1(n5298), .A2(n8011), .ZN(n5299) );
  XNOR2_X1 U6705 ( .A(n5299), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6619) );
  INV_X1 U6706 ( .A(n6619), .ZN(n6654) );
  XNOR2_X1 U6707 ( .A(n5301), .B(n5300), .ZN(n6480) );
  OR2_X1 U6708 ( .A1(n5221), .A2(n6480), .ZN(n5303) );
  OR2_X1 U6709 ( .A1(n6203), .A2(n6478), .ZN(n5302) );
  OAI211_X1 U6710 ( .C1(n6562), .C2(n6654), .A(n5303), .B(n5302), .ZN(n7332)
         );
  XNOR2_X1 U6711 ( .A(n5197), .B(n7332), .ZN(n5306) );
  XNOR2_X1 U6712 ( .A(n5307), .B(n5306), .ZN(n8125) );
  AND2_X1 U6713 ( .A1(n5304), .A2(n8125), .ZN(n5305) );
  NAND2_X1 U6714 ( .A1(n9755), .A2(n5305), .ZN(n8135) );
  INV_X1 U6715 ( .A(n5306), .ZN(n5308) );
  NAND2_X1 U6716 ( .A1(n5308), .A2(n5307), .ZN(n5309) );
  NAND2_X1 U6717 ( .A1(n6190), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5317) );
  INV_X1 U6718 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5310) );
  OR2_X1 U6719 ( .A1(n5349), .A2(n5310), .ZN(n5316) );
  INV_X1 U6720 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6655) );
  NAND2_X1 U6721 ( .A1(n5311), .A2(n6655), .ZN(n5312) );
  NAND2_X1 U6722 ( .A1(n5331), .A2(n5312), .ZN(n7398) );
  OR2_X1 U6723 ( .A1(n5352), .A2(n7398), .ZN(n5315) );
  INV_X1 U6724 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5313) );
  OR2_X1 U6725 ( .A1(n6195), .A2(n5313), .ZN(n5314) );
  NOR2_X1 U6726 ( .A1(n8129), .A2(n6894), .ZN(n5324) );
  NAND2_X1 U6727 ( .A1(n5318), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5319) );
  XNOR2_X1 U6728 ( .A(n5319), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6617) );
  INV_X1 U6729 ( .A(n6617), .ZN(n6666) );
  XNOR2_X1 U6730 ( .A(n5321), .B(n5320), .ZN(n6487) );
  OR2_X1 U6731 ( .A1(n5221), .A2(n6487), .ZN(n5323) );
  OR2_X1 U6732 ( .A1(n6203), .A2(n6488), .ZN(n5322) );
  OAI211_X1 U6733 ( .C1(n6562), .C2(n6666), .A(n5323), .B(n5322), .ZN(n7335)
         );
  XNOR2_X1 U6734 ( .A(n5602), .B(n7335), .ZN(n5325) );
  NAND2_X1 U6735 ( .A1(n5324), .A2(n5325), .ZN(n5329) );
  INV_X1 U6736 ( .A(n5324), .ZN(n5326) );
  INV_X1 U6737 ( .A(n5325), .ZN(n7376) );
  NAND2_X1 U6738 ( .A1(n5326), .A2(n7376), .ZN(n5327) );
  NAND2_X1 U6739 ( .A1(n5329), .A2(n5327), .ZN(n7444) );
  NAND2_X1 U6740 ( .A1(n6190), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5337) );
  INV_X1 U6741 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7522) );
  OR2_X1 U6742 ( .A1(n5349), .A2(n7522), .ZN(n5336) );
  NAND2_X1 U6743 ( .A1(n5331), .A2(n5330), .ZN(n5332) );
  NAND2_X1 U6744 ( .A1(n5350), .A2(n5332), .ZN(n7521) );
  OR2_X1 U6745 ( .A1(n5352), .A2(n7521), .ZN(n5335) );
  INV_X1 U6746 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5333) );
  OR2_X1 U6747 ( .A1(n5213), .A2(n5333), .ZN(n5334) );
  NAND2_X1 U6748 ( .A1(n8583), .A2(n6989), .ZN(n5345) );
  NAND2_X1 U6749 ( .A1(n5338), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5339) );
  XNOR2_X1 U6750 ( .A(n5339), .B(n4671), .ZN(n6817) );
  XNOR2_X1 U6751 ( .A(n5341), .B(n5340), .ZN(n6489) );
  NAND2_X1 U6752 ( .A1(n6489), .A2(n6188), .ZN(n5343) );
  OR2_X1 U6753 ( .A1(n6203), .A2(n6493), .ZN(n5342) );
  OAI211_X1 U6754 ( .C1(n6562), .C2(n6817), .A(n5343), .B(n5342), .ZN(n7528)
         );
  XNOR2_X1 U6755 ( .A(n7528), .B(n5197), .ZN(n5346) );
  XNOR2_X1 U6756 ( .A(n5345), .B(n5346), .ZN(n7374) );
  NAND2_X1 U6757 ( .A1(n5344), .A2(n7374), .ZN(n7377) );
  INV_X1 U6758 ( .A(n5345), .ZN(n5347) );
  NAND2_X1 U6759 ( .A1(n5347), .A2(n5346), .ZN(n5348) );
  NAND2_X1 U6760 ( .A1(n6190), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5357) );
  INV_X1 U6761 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7507) );
  OR2_X1 U6762 ( .A1(n5349), .A2(n7507), .ZN(n5356) );
  INV_X1 U6763 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7550) );
  NAND2_X1 U6764 ( .A1(n5350), .A2(n7550), .ZN(n5351) );
  NAND2_X1 U6765 ( .A1(n5374), .A2(n5351), .ZN(n7549) );
  OR2_X1 U6766 ( .A1(n5352), .A2(n7549), .ZN(n5355) );
  INV_X1 U6767 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5353) );
  OR2_X1 U6768 ( .A1(n5213), .A2(n5353), .ZN(n5354) );
  NOR2_X1 U6769 ( .A1(n7593), .A2(n6894), .ZN(n5363) );
  NAND2_X1 U6770 ( .A1(n6494), .A2(n6188), .ZN(n5362) );
  NAND2_X1 U6771 ( .A1(n5360), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5369) );
  XNOR2_X1 U6772 ( .A(n5369), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6883) );
  AOI22_X1 U6773 ( .A1(n5445), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6518), .B2(
        n6883), .ZN(n5361) );
  XNOR2_X1 U6774 ( .A(n6163), .B(n5197), .ZN(n7542) );
  AND2_X1 U6775 ( .A1(n5363), .A2(n7542), .ZN(n7540) );
  INV_X1 U6776 ( .A(n5363), .ZN(n5365) );
  INV_X1 U6777 ( .A(n7542), .ZN(n5364) );
  NAND2_X1 U6778 ( .A1(n5365), .A2(n5364), .ZN(n7544) );
  XNOR2_X1 U6779 ( .A(n5367), .B(n5366), .ZN(n6508) );
  NAND2_X1 U6780 ( .A1(n6508), .A2(n6188), .ZN(n5372) );
  NAND2_X1 U6781 ( .A1(n5369), .A2(n5368), .ZN(n5370) );
  NAND2_X1 U6782 ( .A1(n5370), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5388) );
  XNOR2_X1 U6783 ( .A(n5388), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6964) );
  AOI22_X1 U6784 ( .A1(n5445), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6518), .B2(
        n6964), .ZN(n5371) );
  XNOR2_X1 U6785 ( .A(n7779), .B(n5602), .ZN(n5381) );
  NAND2_X1 U6786 ( .A1(n6190), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5380) );
  INV_X1 U6787 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7595) );
  OR2_X1 U6788 ( .A1(n5349), .A2(n7595), .ZN(n5379) );
  NAND2_X1 U6789 ( .A1(n5374), .A2(n5373), .ZN(n5375) );
  NAND2_X1 U6790 ( .A1(n5393), .A2(n5375), .ZN(n7594) );
  OR2_X1 U6791 ( .A1(n5352), .A2(n7594), .ZN(n5378) );
  INV_X1 U6792 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5376) );
  OR2_X1 U6793 ( .A1(n5213), .A2(n5376), .ZN(n5377) );
  NOR2_X1 U6794 ( .A1(n7687), .A2(n6894), .ZN(n5382) );
  XNOR2_X1 U6795 ( .A(n5381), .B(n5382), .ZN(n7556) );
  INV_X1 U6796 ( .A(n5381), .ZN(n5384) );
  INV_X1 U6797 ( .A(n5382), .ZN(n5383) );
  XNOR2_X1 U6798 ( .A(n5386), .B(n5385), .ZN(n6513) );
  NAND2_X1 U6799 ( .A1(n6513), .A2(n6188), .ZN(n5392) );
  NAND2_X1 U6800 ( .A1(n5388), .A2(n5387), .ZN(n5389) );
  NAND2_X1 U6801 ( .A1(n5389), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5390) );
  XNOR2_X1 U6802 ( .A(n5390), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7078) );
  AOI22_X1 U6803 ( .A1(n5445), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6518), .B2(
        n7078), .ZN(n5391) );
  XNOR2_X1 U6804 ( .A(n8975), .B(n5629), .ZN(n7680) );
  NAND2_X1 U6805 ( .A1(n6190), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5400) );
  INV_X1 U6806 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6959) );
  OR2_X1 U6807 ( .A1(n5349), .A2(n6959), .ZN(n5399) );
  INV_X1 U6808 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7686) );
  NAND2_X1 U6809 ( .A1(n5393), .A2(n7686), .ZN(n5394) );
  NAND2_X1 U6810 ( .A1(n5395), .A2(n5394), .ZN(n7869) );
  OR2_X1 U6811 ( .A1(n5352), .A2(n7869), .ZN(n5398) );
  INV_X1 U6812 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5396) );
  OR2_X1 U6813 ( .A1(n5213), .A2(n5396), .ZN(n5397) );
  INV_X1 U6814 ( .A(n7788), .ZN(n8580) );
  NAND2_X1 U6815 ( .A1(n8580), .A2(n6989), .ZN(n5401) );
  NAND2_X1 U6816 ( .A1(n7680), .A2(n5401), .ZN(n7684) );
  INV_X1 U6817 ( .A(n7680), .ZN(n5403) );
  INV_X1 U6818 ( .A(n5401), .ZN(n5402) );
  NAND2_X1 U6819 ( .A1(n5403), .A2(n5402), .ZN(n7685) );
  NAND2_X1 U6820 ( .A1(n7682), .A2(n7685), .ZN(n7772) );
  XNOR2_X1 U6821 ( .A(n5405), .B(n5404), .ZN(n7825) );
  AND2_X1 U6822 ( .A1(n7825), .A2(n5406), .ZN(n7937) );
  AND2_X1 U6823 ( .A1(n7937), .A2(n5407), .ZN(n7994) );
  AND2_X1 U6824 ( .A1(n7994), .A2(n5408), .ZN(n7878) );
  INV_X1 U6825 ( .A(n7881), .ZN(n5409) );
  AND2_X1 U6826 ( .A1(n7878), .A2(n5409), .ZN(n5410) );
  NAND2_X1 U6827 ( .A1(n7772), .A2(n5410), .ZN(n5411) );
  INV_X1 U6828 ( .A(n5416), .ZN(n5417) );
  NAND2_X1 U6829 ( .A1(n5417), .A2(SI_17_), .ZN(n5418) );
  MUX2_X1 U6830 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4749), .Z(n5439) );
  XNOR2_X1 U6831 ( .A(n5439), .B(SI_18_), .ZN(n5436) );
  XNOR2_X1 U6832 ( .A(n5438), .B(n5436), .ZN(n6931) );
  NAND2_X1 U6833 ( .A1(n6931), .A2(n6188), .ZN(n5421) );
  XNOR2_X1 U6834 ( .A(n5419), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8643) );
  AOI22_X1 U6835 ( .A1(n5445), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6518), .B2(
        n8643), .ZN(n5420) );
  XNOR2_X1 U6836 ( .A(n8953), .B(n5602), .ZN(n5434) );
  INV_X1 U6837 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8631) );
  OR2_X1 U6838 ( .A1(n5249), .A2(n8631), .ZN(n5431) );
  NAND2_X1 U6839 ( .A1(n6189), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5430) );
  INV_X1 U6840 ( .A(n5426), .ZN(n5423) );
  AND2_X1 U6841 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n5422) );
  NAND2_X1 U6842 ( .A1(n5423), .A2(n5422), .ZN(n5450) );
  INV_X1 U6843 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5424) );
  OAI21_X1 U6844 ( .B1(n5426), .B2(n5425), .A(n5424), .ZN(n5427) );
  NAND2_X1 U6845 ( .A1(n5450), .A2(n5427), .ZN(n7951) );
  OR2_X1 U6846 ( .A1(n5352), .A2(n7951), .ZN(n5429) );
  NAND2_X1 U6847 ( .A1(n6191), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5428) );
  NAND4_X1 U6848 ( .A1(n5431), .A2(n5430), .A3(n5429), .A4(n5428), .ZN(n8573)
         );
  NAND2_X1 U6849 ( .A1(n8573), .A2(n6989), .ZN(n5432) );
  XNOR2_X1 U6850 ( .A(n5434), .B(n5432), .ZN(n7949) );
  INV_X1 U6851 ( .A(n5432), .ZN(n5433) );
  NAND2_X1 U6852 ( .A1(n5434), .A2(n5433), .ZN(n5435) );
  INV_X1 U6853 ( .A(n5436), .ZN(n5437) );
  NAND2_X1 U6854 ( .A1(n5439), .A2(SI_18_), .ZN(n5440) );
  INV_X1 U6855 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7015) );
  INV_X1 U6856 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7017) );
  MUX2_X1 U6857 ( .A(n7015), .B(n7017), .S(n4749), .Z(n5442) );
  INV_X1 U6858 ( .A(SI_19_), .ZN(n10064) );
  NAND2_X1 U6859 ( .A1(n5442), .A2(n10064), .ZN(n5464) );
  INV_X1 U6860 ( .A(n5442), .ZN(n5443) );
  NAND2_X1 U6861 ( .A1(n5443), .A2(SI_19_), .ZN(n5444) );
  NAND2_X1 U6862 ( .A1(n5464), .A2(n5444), .ZN(n5465) );
  XNOR2_X1 U6863 ( .A(n5466), .B(n5465), .ZN(n7014) );
  NAND2_X1 U6864 ( .A1(n7014), .A2(n6188), .ZN(n5447) );
  AOI22_X1 U6865 ( .A1(n5445), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n4385), .B2(
        n6518), .ZN(n5446) );
  XNOR2_X1 U6866 ( .A(n8949), .B(n5629), .ZN(n5456) );
  NAND2_X1 U6867 ( .A1(n6189), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5455) );
  INV_X1 U6868 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n5448) );
  OR2_X1 U6869 ( .A1(n5249), .A2(n5448), .ZN(n5454) );
  INV_X1 U6870 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8816) );
  OR2_X1 U6871 ( .A1(n5349), .A2(n8816), .ZN(n5453) );
  INV_X1 U6872 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5449) );
  NAND2_X1 U6873 ( .A1(n5450), .A2(n5449), .ZN(n5451) );
  NAND2_X1 U6874 ( .A1(n5474), .A2(n5451), .ZN(n8815) );
  OR2_X1 U6875 ( .A1(n5352), .A2(n8815), .ZN(n5452) );
  INV_X1 U6876 ( .A(n8831), .ZN(n8806) );
  NAND2_X1 U6877 ( .A1(n8806), .A2(n6989), .ZN(n5457) );
  NAND2_X1 U6878 ( .A1(n5456), .A2(n5457), .ZN(n5463) );
  INV_X1 U6879 ( .A(n5456), .ZN(n5459) );
  INV_X1 U6880 ( .A(n5457), .ZN(n5458) );
  NAND2_X1 U6881 ( .A1(n5459), .A2(n5458), .ZN(n5460) );
  NAND2_X1 U6882 ( .A1(n5463), .A2(n5460), .ZN(n8488) );
  NAND2_X1 U6883 ( .A1(n5462), .A2(n5461), .ZN(n8486) );
  INV_X1 U6884 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n9957) );
  INV_X1 U6885 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7123) );
  MUX2_X1 U6886 ( .A(n9957), .B(n7123), .S(n6051), .Z(n5467) );
  INV_X1 U6887 ( .A(SI_20_), .ZN(n10144) );
  NAND2_X1 U6888 ( .A1(n5467), .A2(n10144), .ZN(n5486) );
  INV_X1 U6889 ( .A(n5467), .ZN(n5468) );
  NAND2_X1 U6890 ( .A1(n5468), .A2(SI_20_), .ZN(n5469) );
  AND2_X1 U6891 ( .A1(n5486), .A2(n5469), .ZN(n5484) );
  XNOR2_X1 U6892 ( .A(n5485), .B(n5484), .ZN(n7122) );
  NAND2_X1 U6893 ( .A1(n7122), .A2(n6188), .ZN(n5471) );
  OR2_X1 U6894 ( .A1(n6203), .A2(n9957), .ZN(n5470) );
  XNOR2_X1 U6895 ( .A(n8942), .B(n5602), .ZN(n5480) );
  NAND2_X1 U6896 ( .A1(n6190), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5479) );
  INV_X1 U6897 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n5472) );
  OR2_X1 U6898 ( .A1(n5349), .A2(n5472), .ZN(n5478) );
  INV_X1 U6899 ( .A(n5474), .ZN(n5473) );
  NAND2_X1 U6900 ( .A1(n5473), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5490) );
  INV_X1 U6901 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8561) );
  NAND2_X1 U6902 ( .A1(n5474), .A2(n8561), .ZN(n5475) );
  NAND2_X1 U6903 ( .A1(n5490), .A2(n5475), .ZN(n8799) );
  OR2_X1 U6904 ( .A1(n5352), .A2(n8799), .ZN(n5477) );
  INV_X1 U6905 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n10173) );
  OR2_X1 U6906 ( .A1(n6195), .A2(n10173), .ZN(n5476) );
  NOR2_X1 U6907 ( .A1(n8496), .A2(n6894), .ZN(n5481) );
  XNOR2_X1 U6908 ( .A(n5480), .B(n5481), .ZN(n8559) );
  INV_X1 U6909 ( .A(n5480), .ZN(n5483) );
  INV_X1 U6910 ( .A(n5481), .ZN(n5482) );
  MUX2_X1 U6911 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n6051), .Z(n5503) );
  INV_X1 U6912 ( .A(SI_21_), .ZN(n9970) );
  XNOR2_X1 U6913 ( .A(n5503), .B(n9970), .ZN(n5500) );
  XNOR2_X1 U6914 ( .A(n5502), .B(n5500), .ZN(n7251) );
  NAND2_X1 U6915 ( .A1(n7251), .A2(n6188), .ZN(n5488) );
  INV_X1 U6916 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7253) );
  OR2_X1 U6917 ( .A1(n6203), .A2(n7253), .ZN(n5487) );
  XNOR2_X1 U6918 ( .A(n8787), .B(n5602), .ZN(n5497) );
  NAND2_X1 U6919 ( .A1(n6190), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5496) );
  INV_X1 U6920 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n5489) );
  OR2_X1 U6921 ( .A1(n5349), .A2(n5489), .ZN(n5495) );
  INV_X1 U6922 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10151) );
  NAND2_X1 U6923 ( .A1(n5490), .A2(n10151), .ZN(n5491) );
  NAND2_X1 U6924 ( .A1(n5523), .A2(n5491), .ZN(n8784) );
  OR2_X1 U6925 ( .A1(n5352), .A2(n8784), .ZN(n5494) );
  INV_X1 U6926 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n5492) );
  OR2_X1 U6927 ( .A1(n6195), .A2(n5492), .ZN(n5493) );
  NOR2_X1 U6928 ( .A1(n8562), .A2(n6894), .ZN(n5498) );
  XNOR2_X1 U6929 ( .A(n5497), .B(n5498), .ZN(n8494) );
  INV_X1 U6930 ( .A(n5497), .ZN(n5499) );
  INV_X1 U6931 ( .A(n5500), .ZN(n5501) );
  NAND2_X1 U6932 ( .A1(n5503), .A2(SI_21_), .ZN(n5504) );
  INV_X1 U6933 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7408) );
  INV_X1 U6934 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8420) );
  MUX2_X1 U6935 ( .A(n7408), .B(n8420), .S(n4749), .Z(n5506) );
  INV_X1 U6936 ( .A(SI_22_), .ZN(n5505) );
  NAND2_X1 U6937 ( .A1(n5506), .A2(n5505), .ZN(n5536) );
  INV_X1 U6938 ( .A(n5506), .ZN(n5507) );
  NAND2_X1 U6939 ( .A1(n5507), .A2(SI_22_), .ZN(n5508) );
  NAND2_X1 U6940 ( .A1(n5536), .A2(n5508), .ZN(n5535) );
  XNOR2_X1 U6941 ( .A(n5577), .B(n5535), .ZN(n7406) );
  NAND2_X1 U6942 ( .A1(n7406), .A2(n6188), .ZN(n5510) );
  OR2_X1 U6943 ( .A1(n6203), .A2(n7408), .ZN(n5509) );
  XNOR2_X1 U6944 ( .A(n8932), .B(n5629), .ZN(n5530) );
  XNOR2_X1 U6945 ( .A(n5523), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n8770) );
  INV_X1 U6946 ( .A(n5352), .ZN(n5682) );
  AOI22_X1 U6947 ( .A1(n8770), .A2(n5682), .B1(n6189), .B2(
        P2_REG0_REG_22__SCAN_IN), .ZN(n5513) );
  AOI22_X1 U6948 ( .A1(n6190), .A2(P2_REG1_REG_22__SCAN_IN), .B1(n6191), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n5512) );
  OR2_X1 U6949 ( .A1(n8572), .A2(n6894), .ZN(n5514) );
  NAND2_X1 U6950 ( .A1(n8034), .A2(n5514), .ZN(n8031) );
  INV_X1 U6951 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7453) );
  INV_X1 U6952 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7457) );
  MUX2_X1 U6953 ( .A(n7453), .B(n7457), .S(n6051), .Z(n5516) );
  INV_X1 U6954 ( .A(SI_23_), .ZN(n5515) );
  NAND2_X1 U6955 ( .A1(n5516), .A2(n5515), .ZN(n5538) );
  INV_X1 U6956 ( .A(n5516), .ZN(n5517) );
  NAND2_X1 U6957 ( .A1(n5517), .A2(SI_23_), .ZN(n5518) );
  NAND2_X1 U6958 ( .A1(n7454), .A2(n6188), .ZN(n5520) );
  OR2_X1 U6959 ( .A1(n6203), .A2(n7453), .ZN(n5519) );
  XNOR2_X1 U6960 ( .A(n8927), .B(n5629), .ZN(n8475) );
  NAND2_X1 U6961 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n5521) );
  INV_X1 U6962 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n5522) );
  INV_X1 U6963 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9984) );
  OAI21_X1 U6964 ( .B1(n5523), .B2(n5522), .A(n9984), .ZN(n5524) );
  AND2_X1 U6965 ( .A1(n5545), .A2(n5524), .ZN(n8757) );
  NAND2_X1 U6966 ( .A1(n8757), .A2(n5682), .ZN(n5529) );
  NAND2_X1 U6967 ( .A1(n6190), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U6968 ( .A1(n6189), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5525) );
  AND2_X1 U6969 ( .A1(n5526), .A2(n5525), .ZN(n5528) );
  NAND2_X1 U6970 ( .A1(n6191), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5527) );
  INV_X1 U6971 ( .A(n8746), .ZN(n8571) );
  NAND2_X1 U6972 ( .A1(n8571), .A2(n6989), .ZN(n8478) );
  AOI21_X1 U6973 ( .B1(n8475), .B2(n8478), .A(n8473), .ZN(n5533) );
  INV_X1 U6974 ( .A(n8478), .ZN(n5532) );
  INV_X1 U6975 ( .A(n8475), .ZN(n5531) );
  INV_X1 U6976 ( .A(n5534), .ZN(n5537) );
  OR2_X1 U6977 ( .A1(n5535), .A2(n5537), .ZN(n5554) );
  OR2_X1 U6978 ( .A1(n5537), .A2(n5536), .ZN(n5539) );
  MUX2_X1 U6979 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n4749), .Z(n5553) );
  XNOR2_X1 U6980 ( .A(n5553), .B(n10027), .ZN(n5555) );
  NAND2_X1 U6981 ( .A1(n7458), .A2(n6188), .ZN(n5543) );
  INV_X1 U6982 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7483) );
  OR2_X1 U6983 ( .A1(n6203), .A2(n7483), .ZN(n5542) );
  XNOR2_X1 U6984 ( .A(n8922), .B(n5602), .ZN(n5551) );
  XNOR2_X1 U6985 ( .A(n5550), .B(n5551), .ZN(n8535) );
  INV_X1 U6986 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10109) );
  NAND2_X1 U6987 ( .A1(n5545), .A2(n10109), .ZN(n5546) );
  NAND2_X1 U6988 ( .A1(n5583), .A2(n5546), .ZN(n8738) );
  OR2_X1 U6989 ( .A1(n8738), .A2(n5352), .ZN(n5549) );
  AOI22_X1 U6990 ( .A1(n6190), .A2(P2_REG1_REG_24__SCAN_IN), .B1(n6191), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U6991 ( .A1(n6189), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5547) );
  NOR2_X1 U6992 ( .A1(n8505), .A2(n6894), .ZN(n8534) );
  INV_X1 U6993 ( .A(n5550), .ZN(n5552) );
  AOI22_X2 U6994 ( .A1(n8535), .A2(n8534), .B1(n5552), .B2(n5551), .ZN(n8504)
         );
  AND2_X1 U6995 ( .A1(n5553), .A2(SI_24_), .ZN(n5558) );
  OR2_X1 U6996 ( .A1(n5554), .A2(n5558), .ZN(n5570) );
  INV_X1 U6997 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7537) );
  INV_X1 U6998 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9958) );
  MUX2_X1 U6999 ( .A(n7537), .B(n9958), .S(n4749), .Z(n5560) );
  INV_X1 U7000 ( .A(SI_25_), .ZN(n10009) );
  NAND2_X1 U7001 ( .A1(n5560), .A2(n10009), .ZN(n5573) );
  INV_X1 U7002 ( .A(n5560), .ZN(n5561) );
  NAND2_X1 U7003 ( .A1(n5561), .A2(SI_25_), .ZN(n5562) );
  NAND2_X1 U7004 ( .A1(n5573), .A2(n5562), .ZN(n5572) );
  NAND2_X1 U7005 ( .A1(n7535), .A2(n6188), .ZN(n5565) );
  OR2_X1 U7006 ( .A1(n6203), .A2(n7537), .ZN(n5564) );
  XNOR2_X1 U7007 ( .A(n4759), .B(n5602), .ZN(n8502) );
  XNOR2_X1 U7008 ( .A(n5583), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n8730) );
  INV_X1 U7009 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U7010 ( .A1(n6189), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5567) );
  NAND2_X1 U7011 ( .A1(n6190), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5566) );
  OAI211_X1 U7012 ( .C1(n5349), .C2(n5568), .A(n5567), .B(n5566), .ZN(n5569)
         );
  AOI21_X1 U7013 ( .B1(n8730), .B2(n5682), .A(n5569), .ZN(n8747) );
  INV_X1 U7014 ( .A(n8747), .ZN(n8570) );
  NAND2_X1 U7015 ( .A1(n8570), .A2(n6989), .ZN(n8501) );
  OR2_X1 U7016 ( .A1(n5570), .A2(n5572), .ZN(n5576) );
  INV_X1 U7017 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7563) );
  INV_X1 U7018 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7533) );
  MUX2_X1 U7019 ( .A(n7563), .B(n7533), .S(n6051), .Z(n5578) );
  INV_X1 U7020 ( .A(SI_26_), .ZN(n10155) );
  NAND2_X1 U7021 ( .A1(n5578), .A2(n10155), .ZN(n5595) );
  INV_X1 U7022 ( .A(n5578), .ZN(n5579) );
  NAND2_X1 U7023 ( .A1(n5579), .A2(SI_26_), .ZN(n5580) );
  AND2_X1 U7024 ( .A1(n5595), .A2(n5580), .ZN(n5593) );
  NAND2_X1 U7025 ( .A1(n7532), .A2(n6188), .ZN(n5582) );
  OR2_X1 U7026 ( .A1(n6203), .A2(n7563), .ZN(n5581) );
  XNOR2_X1 U7027 ( .A(n8914), .B(n5602), .ZN(n8462) );
  INV_X1 U7028 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8507) );
  INV_X1 U7029 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6454) );
  OAI21_X1 U7030 ( .B1(n5583), .B2(n8507), .A(n6454), .ZN(n5584) );
  NAND2_X1 U7031 ( .A1(n5584), .A2(n5604), .ZN(n8713) );
  OR2_X1 U7032 ( .A1(n8713), .A2(n5352), .ZN(n5590) );
  INV_X1 U7033 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U7034 ( .A1(n6191), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5586) );
  NAND2_X1 U7035 ( .A1(n6190), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5585) );
  OAI211_X1 U7036 ( .C1(n5587), .C2(n6195), .A(n5586), .B(n5585), .ZN(n5588)
         );
  INV_X1 U7037 ( .A(n5588), .ZN(n5589) );
  NOR2_X1 U7038 ( .A1(n8687), .A2(n6894), .ZN(n5591) );
  NAND2_X1 U7039 ( .A1(n8462), .A2(n5591), .ZN(n5592) );
  OAI21_X1 U7040 ( .B1(n8462), .B2(n5591), .A(n5592), .ZN(n6453) );
  NAND2_X1 U7041 ( .A1(n5594), .A2(n5593), .ZN(n5596) );
  INV_X1 U7042 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7679) );
  INV_X1 U7043 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7603) );
  MUX2_X1 U7044 ( .A(n7679), .B(n7603), .S(n4749), .Z(n5597) );
  INV_X1 U7045 ( .A(SI_27_), .ZN(n10150) );
  NAND2_X1 U7046 ( .A1(n5597), .A2(n10150), .ZN(n5619) );
  INV_X1 U7047 ( .A(n5597), .ZN(n5598) );
  NAND2_X1 U7048 ( .A1(n5598), .A2(SI_27_), .ZN(n5599) );
  AND2_X1 U7049 ( .A1(n5619), .A2(n5599), .ZN(n5617) );
  OR2_X1 U7050 ( .A1(n6203), .A2(n7679), .ZN(n5600) );
  XNOR2_X1 U7051 ( .A(n8907), .B(n5602), .ZN(n5611) );
  INV_X1 U7052 ( .A(n5604), .ZN(n5603) );
  NAND2_X1 U7053 ( .A1(n5603), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5624) );
  INV_X1 U7054 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10176) );
  NAND2_X1 U7055 ( .A1(n5604), .A2(n10176), .ZN(n5605) );
  NAND2_X1 U7056 ( .A1(n5624), .A2(n5605), .ZN(n8466) );
  OR2_X1 U7057 ( .A1(n8466), .A2(n5352), .ZN(n5610) );
  INV_X1 U7058 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n10039) );
  NAND2_X1 U7059 ( .A1(n6190), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5607) );
  NAND2_X1 U7060 ( .A1(n6191), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5606) );
  OAI211_X1 U7061 ( .C1(n10039), .C2(n6195), .A(n5607), .B(n5606), .ZN(n5608)
         );
  INV_X1 U7062 ( .A(n5608), .ZN(n5609) );
  NOR2_X1 U7063 ( .A1(n8707), .A2(n6894), .ZN(n5612) );
  NAND2_X1 U7064 ( .A1(n5611), .A2(n5612), .ZN(n5616) );
  INV_X1 U7065 ( .A(n5611), .ZN(n5614) );
  INV_X1 U7066 ( .A(n5612), .ZN(n5613) );
  NAND2_X1 U7067 ( .A1(n5614), .A2(n5613), .ZN(n5615) );
  NAND2_X1 U7068 ( .A1(n8470), .A2(n5616), .ZN(n5676) );
  INV_X1 U7069 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n10145) );
  INV_X1 U7070 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7713) );
  MUX2_X1 U7071 ( .A(n10145), .B(n7713), .S(n6051), .Z(n6049) );
  XNOR2_X1 U7072 ( .A(n6049), .B(SI_28_), .ZN(n6046) );
  NAND2_X1 U7073 ( .A1(n8457), .A2(n6188), .ZN(n5622) );
  OR2_X1 U7074 ( .A1(n6203), .A2(n10145), .ZN(n5621) );
  INV_X1 U7075 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5623) );
  OR2_X1 U7076 ( .A1(n5624), .A2(n5623), .ZN(n5677) );
  NAND2_X1 U7077 ( .A1(n5624), .A2(n5623), .ZN(n5625) );
  INV_X1 U7078 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9985) );
  NAND2_X1 U7079 ( .A1(n6191), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U7080 ( .A1(n6189), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5626) );
  OAI211_X1 U7081 ( .C1(n5249), .C2(n9985), .A(n5627), .B(n5626), .ZN(n5628)
         );
  AOI21_X1 U7082 ( .B1(n8666), .B2(n5682), .A(n5628), .ZN(n8442) );
  OR2_X1 U7083 ( .A1(n8442), .A2(n6894), .ZN(n5630) );
  XNOR2_X1 U7084 ( .A(n5630), .B(n5629), .ZN(n5668) );
  INV_X1 U7085 ( .A(n5668), .ZN(n5669) );
  AND2_X2 U7086 ( .A1(n6383), .A2(n6991), .ZN(n9818) );
  NOR3_X1 U7087 ( .A1(n8668), .A2(n9818), .A3(n5669), .ZN(n5631) );
  AOI21_X1 U7088 ( .B1(n8668), .B2(n5669), .A(n5631), .ZN(n5675) );
  AND2_X1 U7089 ( .A1(n4385), .A2(n7407), .ZN(n5633) );
  NAND2_X1 U7090 ( .A1(n5635), .A2(n5634), .ZN(n5636) );
  NAND2_X1 U7091 ( .A1(n5636), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5647) );
  INV_X1 U7092 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5646) );
  NAND2_X1 U7093 ( .A1(n5647), .A2(n5646), .ZN(n5649) );
  NAND2_X1 U7094 ( .A1(n5649), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5638) );
  INV_X1 U7095 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5637) );
  XNOR2_X1 U7096 ( .A(n5638), .B(n5637), .ZN(n7485) );
  INV_X1 U7097 ( .A(n7485), .ZN(n5645) );
  NAND2_X1 U7098 ( .A1(n4470), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5639) );
  MUX2_X1 U7099 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5639), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5640) );
  NAND2_X1 U7100 ( .A1(n5640), .A2(n5054), .ZN(n7565) );
  NAND2_X1 U7101 ( .A1(n5641), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5642) );
  MUX2_X1 U7102 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5642), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5643) );
  NAND2_X1 U7103 ( .A1(n5643), .A2(n4470), .ZN(n7536) );
  NOR2_X1 U7104 ( .A1(n7565), .A2(n7536), .ZN(n5644) );
  NAND2_X1 U7105 ( .A1(n5645), .A2(n5644), .ZN(n6558) );
  OR2_X1 U7106 ( .A1(n5647), .A2(n5646), .ZN(n5648) );
  NAND2_X1 U7107 ( .A1(n5649), .A2(n5648), .ZN(n6382) );
  NAND2_X1 U7108 ( .A1(n6558), .A2(n9798), .ZN(n9790) );
  NOR2_X1 U7109 ( .A1(n9790), .A2(n6243), .ZN(n5650) );
  XNOR2_X1 U7110 ( .A(n7485), .B(P2_B_REG_SCAN_IN), .ZN(n5651) );
  NAND2_X1 U7111 ( .A1(n5651), .A2(n7536), .ZN(n5653) );
  INV_X1 U7112 ( .A(n7565), .ZN(n5652) );
  INV_X1 U7113 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9796) );
  AND2_X1 U7114 ( .A1(n7565), .A2(n7536), .ZN(n9797) );
  AOI21_X1 U7115 ( .B1(n9791), .B2(n9796), .A(n9797), .ZN(n7259) );
  NOR2_X1 U7116 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .ZN(
        n5657) );
  NOR4_X1 U7117 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n5656) );
  NOR4_X1 U7118 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n5655) );
  NOR4_X1 U7119 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5654) );
  NAND4_X1 U7120 ( .A1(n5657), .A2(n5656), .A3(n5655), .A4(n5654), .ZN(n5663)
         );
  NOR4_X1 U7121 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n5661) );
  NOR4_X1 U7122 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n5660) );
  NOR4_X1 U7123 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n5659) );
  NOR4_X1 U7124 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n5658) );
  NAND4_X1 U7125 ( .A1(n5661), .A2(n5660), .A3(n5659), .A4(n5658), .ZN(n5662)
         );
  OAI21_X1 U7126 ( .B1(n5663), .B2(n5662), .A(n9791), .ZN(n7256) );
  NAND2_X1 U7127 ( .A1(n7259), .A2(n7256), .ZN(n5685) );
  NOR2_X1 U7128 ( .A1(n9790), .A2(n5685), .ZN(n6975) );
  INV_X1 U7129 ( .A(n6975), .ZN(n5666) );
  INV_X1 U7130 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9794) );
  NAND2_X1 U7131 ( .A1(n9791), .A2(n9794), .ZN(n5665) );
  AND2_X1 U7132 ( .A1(n7565), .A2(n7485), .ZN(n9793) );
  INV_X1 U7133 ( .A(n9793), .ZN(n5664) );
  NAND2_X1 U7134 ( .A1(n5665), .A2(n5664), .ZN(n7268) );
  OR2_X1 U7135 ( .A1(n5666), .A2(n7268), .ZN(n5683) );
  NAND2_X1 U7136 ( .A1(n9778), .A2(n5683), .ZN(n8529) );
  NAND2_X1 U7137 ( .A1(n8529), .A2(n9818), .ZN(n9747) );
  OR2_X1 U7138 ( .A1(n9818), .A2(n6561), .ZN(n5667) );
  OR2_X2 U7139 ( .A1(n5667), .A2(n5683), .ZN(n9743) );
  OAI21_X1 U7140 ( .B1(n8668), .B2(n9747), .A(n9743), .ZN(n5674) );
  NOR3_X1 U7141 ( .A1(n8668), .A2(n9818), .A3(n5668), .ZN(n5671) );
  NOR2_X1 U7142 ( .A1(n8902), .A2(n5669), .ZN(n5670) );
  NAND2_X1 U7143 ( .A1(n5676), .A2(n5672), .ZN(n5673) );
  OAI211_X1 U7144 ( .C1(n5676), .C2(n5675), .A(n5674), .B(n5673), .ZN(n5692)
         );
  INV_X1 U7145 ( .A(n5677), .ZN(n8445) );
  INV_X1 U7146 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5680) );
  NAND2_X1 U7147 ( .A1(n6190), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U7148 ( .A1(n6191), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5678) );
  OAI211_X1 U7149 ( .C1(n5680), .C2(n6195), .A(n5679), .B(n5678), .ZN(n5681)
         );
  AOI21_X1 U7150 ( .B1(n8445), .B2(n5682), .A(n5681), .ZN(n6179) );
  INV_X1 U7151 ( .A(n6179), .ZN(n8671) );
  OR2_X1 U7152 ( .A1(n5683), .A2(n6383), .ZN(n8508) );
  AND2_X1 U7153 ( .A1(n5684), .A2(n6561), .ZN(n9774) );
  NOR2_X1 U7154 ( .A1(n8508), .A2(n8882), .ZN(n8465) );
  NAND2_X1 U7155 ( .A1(n9845), .A2(n7252), .ZN(n7255) );
  OAI21_X1 U7156 ( .B1(n5685), .B2(n7268), .A(n7255), .ZN(n5686) );
  NAND2_X1 U7157 ( .A1(n6383), .A2(n6561), .ZN(n7257) );
  NAND4_X1 U7158 ( .A1(n5686), .A2(n6558), .A3(n6382), .A4(n7257), .ZN(n5687)
         );
  NAND2_X1 U7159 ( .A1(n5687), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9759) );
  INV_X1 U7160 ( .A(n9759), .ZN(n8511) );
  AOI22_X1 U7161 ( .A1(n8671), .A2(n8465), .B1(n8666), .B2(n8511), .ZN(n5690)
         );
  INV_X1 U7162 ( .A(n8707), .ZN(n8672) );
  INV_X1 U7163 ( .A(n5684), .ZN(n5688) );
  NOR2_X1 U7164 ( .A1(n8508), .A2(n8880), .ZN(n8554) );
  AOI22_X1 U7165 ( .A1(n8672), .A2(n8554), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n5689) );
  AND2_X1 U7166 ( .A1(n5690), .A2(n5689), .ZN(n5691) );
  NAND2_X1 U7167 ( .A1(n5692), .A2(n5691), .ZN(P2_U3222) );
  NAND2_X1 U7168 ( .A1(n5761), .A2(n5693), .ZN(n5779) );
  INV_X1 U7169 ( .A(n5779), .ZN(n5697) );
  NOR2_X1 U7170 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5699) );
  NOR2_X1 U7171 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5700) );
  INV_X1 U7172 ( .A(n5924), .ZN(n5702) );
  NAND2_X1 U7173 ( .A1(n5702), .A2(n5701), .ZN(n5933) );
  NOR2_X1 U7174 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5703) );
  OR2_X1 U7175 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5709) );
  OR2_X1 U7176 ( .A1(n5709), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n5705) );
  OR2_X1 U7177 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n5704) );
  INV_X1 U7178 ( .A(n5706), .ZN(n5713) );
  NAND2_X1 U7179 ( .A1(n5715), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5708) );
  OR2_X1 U7180 ( .A1(n6149), .A2(n9350), .ZN(n5719) );
  INV_X1 U7181 ( .A(n5715), .ZN(n5711) );
  INV_X1 U7182 ( .A(n5709), .ZN(n5710) );
  NAND2_X1 U7183 ( .A1(n5711), .A2(n5710), .ZN(n5712) );
  NAND2_X1 U7184 ( .A1(n5712), .A2(n4953), .ZN(n5714) );
  XNOR2_X1 U7185 ( .A(n5717), .B(P1_IR_REG_20__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7186 ( .A1(n5719), .A2(n5718), .ZN(n9635) );
  NOR2_X1 U7187 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5721) );
  NOR2_X1 U7188 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5720) );
  NAND4_X1 U7189 ( .A1(n5721), .A2(n5720), .A3(n5701), .A4(n10119), .ZN(n5726)
         );
  INV_X1 U7190 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5723) );
  NAND4_X1 U7191 ( .A1(n5724), .A2(n5912), .A3(n5723), .A4(n5722), .ZN(n5725)
         );
  NOR2_X1 U7192 ( .A1(n5726), .A2(n5725), .ZN(n5727) );
  INV_X1 U7193 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n10117) );
  INV_X1 U7194 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5729) );
  INV_X1 U7195 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5728) );
  INV_X1 U7196 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5742) );
  INV_X1 U7197 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5731) );
  XNOR2_X2 U7198 ( .A(n5732), .B(n5731), .ZN(n5737) );
  INV_X1 U7199 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5733) );
  INV_X1 U7200 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5734) );
  NAND2_X2 U7201 ( .A1(n5737), .A2(n5735), .ZN(n5784) );
  NAND2_X1 U7202 ( .A1(n5790), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5740) );
  INV_X1 U7203 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7150) );
  NAND4_X2 U7204 ( .A1(n5741), .A2(n5740), .A3(n5739), .A4(n5738), .ZN(n9130)
         );
  NAND2_X1 U7205 ( .A1(n5744), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5746) );
  INV_X1 U7206 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5745) );
  INV_X1 U7207 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5747) );
  INV_X1 U7208 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6462) );
  XNOR2_X2 U7209 ( .A(n9130), .B(n7142), .ZN(n8255) );
  INV_X1 U7210 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5748) );
  NAND2_X1 U7211 ( .A1(n5790), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5752) );
  INV_X1 U7212 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5749) );
  OR2_X1 U7213 ( .A1(n5791), .A2(n5749), .ZN(n5751) );
  NAND2_X1 U7214 ( .A1(n5789), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5750) );
  INV_X1 U7215 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6693) );
  XNOR2_X1 U7216 ( .A(n5755), .B(n5754), .ZN(n6459) );
  NAND2_X1 U7217 ( .A1(n8255), .A2(n7144), .ZN(n7143) );
  INV_X1 U7218 ( .A(n9130), .ZN(n7194) );
  NAND2_X1 U7219 ( .A1(n7194), .A2(n7142), .ZN(n5756) );
  NAND2_X1 U7220 ( .A1(n7143), .A2(n5756), .ZN(n8373) );
  INV_X1 U7221 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9729) );
  INV_X1 U7222 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7198) );
  OR2_X1 U7223 ( .A1(n5791), .A2(n7198), .ZN(n5759) );
  NAND2_X1 U7224 ( .A1(n5789), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5758) );
  INV_X1 U7225 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7199) );
  OR2_X1 U7226 ( .A1(n5761), .A2(n8006), .ZN(n5763) );
  INV_X1 U7227 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5762) );
  NAND2_X1 U7228 ( .A1(n5763), .A2(n5762), .ZN(n5773) );
  OAI21_X1 U7229 ( .B1(n5763), .B2(n5762), .A(n5773), .ZN(n6463) );
  OR2_X1 U7230 ( .A1(n4387), .A2(n6464), .ZN(n5764) );
  NAND2_X1 U7231 ( .A1(n7160), .A2(n7205), .ZN(n8370) );
  AND2_X1 U7232 ( .A1(n8370), .A2(n8371), .ZN(n7193) );
  NAND2_X1 U7233 ( .A1(n8373), .A2(n7193), .ZN(n7192) );
  NAND2_X1 U7234 ( .A1(n7192), .A2(n8370), .ZN(n7157) );
  NAND2_X1 U7235 ( .A1(n6041), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5772) );
  INV_X1 U7236 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5765) );
  OR2_X1 U7237 ( .A1(n5791), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5766) );
  NAND2_X1 U7238 ( .A1(n5767), .A2(n5766), .ZN(n5770) );
  INV_X1 U7239 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5768) );
  NAND2_X1 U7240 ( .A1(n5773), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5775) );
  INV_X1 U7241 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5774) );
  XNOR2_X1 U7242 ( .A(n5775), .B(n5774), .ZN(n6465) );
  OR2_X1 U7243 ( .A1(n4386), .A2(n6466), .ZN(n5777) );
  OR2_X1 U7244 ( .A1(n8137), .A2(n6471), .ZN(n5776) );
  OAI211_X1 U7245 ( .C1(n5778), .C2(n6465), .A(n5777), .B(n5776), .ZN(n7166)
         );
  AND2_X1 U7246 ( .A1(n8319), .A2(n8313), .ZN(n7159) );
  NAND2_X1 U7247 ( .A1(n7157), .A2(n7159), .ZN(n7158) );
  NAND2_X1 U7248 ( .A1(n7158), .A2(n8319), .ZN(n7176) );
  INV_X2 U7249 ( .A(n5778), .ZN(n6387) );
  NAND2_X1 U7250 ( .A1(n5779), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5780) );
  MUX2_X1 U7251 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5780), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5781) );
  NOR2_X1 U7252 ( .A1(n5779), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5808) );
  INV_X1 U7253 ( .A(n5808), .ZN(n5798) );
  AOI22_X1 U7254 ( .A1(n5797), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n6387), .B2(
        n9584), .ZN(n5783) );
  OR2_X1 U7255 ( .A1(n6469), .A2(n8137), .ZN(n5782) );
  OR2_X1 U7256 ( .A1(n5784), .A2(n9732), .ZN(n5788) );
  XNOR2_X1 U7257 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n9064) );
  OR2_X1 U7258 ( .A1(n5791), .A2(n9064), .ZN(n5787) );
  INV_X1 U7259 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7182) );
  OR2_X1 U7260 ( .A1(n6058), .A2(n7182), .ZN(n5786) );
  NAND2_X1 U7261 ( .A1(n5789), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U7262 ( .A1(n5789), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5796) );
  INV_X1 U7263 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6398) );
  OR2_X1 U7264 ( .A1(n6058), .A2(n6398), .ZN(n5795) );
  NAND2_X1 U7265 ( .A1(n5790), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5794) );
  INV_X1 U7266 ( .A(n5791), .ZN(n5948) );
  AOI21_X1 U7267 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5792) );
  NOR2_X1 U7268 ( .A1(n5792), .A2(n5802), .ZN(n9652) );
  NAND2_X1 U7269 ( .A1(n5948), .A2(n9652), .ZN(n5793) );
  INV_X1 U7270 ( .A(n9126), .ZN(n7048) );
  OR2_X1 U7271 ( .A1(n6476), .A2(n8137), .ZN(n5801) );
  NAND2_X1 U7272 ( .A1(n5798), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5799) );
  XNOR2_X1 U7273 ( .A(n5799), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6590) );
  AOI22_X1 U7274 ( .A1(n5797), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6387), .B2(
        n6590), .ZN(n5800) );
  AND2_X1 U7275 ( .A1(n7048), .A2(n9651), .ZN(n8315) );
  INV_X1 U7276 ( .A(n9651), .ZN(n9698) );
  OAI21_X1 U7277 ( .B1(n5802), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5817), .ZN(
        n7056) );
  OR2_X1 U7278 ( .A1(n5791), .A2(n7056), .ZN(n5806) );
  INV_X1 U7279 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7057) );
  OR2_X1 U7280 ( .A1(n6058), .A2(n7057), .ZN(n5805) );
  NAND2_X1 U7281 ( .A1(n5790), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U7282 ( .A1(n5789), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5803) );
  NAND4_X1 U7283 ( .A1(n5806), .A2(n5805), .A3(n5804), .A4(n5803), .ZN(n9125)
         );
  OR2_X1 U7284 ( .A1(n6480), .A2(n8137), .ZN(n5811) );
  NAND2_X1 U7285 ( .A1(n5808), .A2(n5807), .ZN(n5812) );
  NAND2_X1 U7286 ( .A1(n5812), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5809) );
  XNOR2_X1 U7287 ( .A(n5809), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6479) );
  AOI22_X1 U7288 ( .A1(n5797), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6387), .B2(
        n6479), .ZN(n5810) );
  NAND2_X1 U7289 ( .A1(n5811), .A2(n5810), .ZN(n7059) );
  OR2_X1 U7290 ( .A1(n9661), .A2(n7059), .ZN(n7022) );
  NAND2_X1 U7291 ( .A1(n7059), .A2(n9661), .ZN(n8322) );
  OR2_X1 U7292 ( .A1(n6487), .A2(n8137), .ZN(n5815) );
  OAI21_X1 U7293 ( .B1(n5812), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5813) );
  XNOR2_X1 U7294 ( .A(n5813), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9148) );
  AOI22_X1 U7295 ( .A1(n5797), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6387), .B2(
        n9148), .ZN(n5814) );
  NAND2_X1 U7296 ( .A1(n5815), .A2(n5814), .ZN(n7036) );
  INV_X1 U7297 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7034) );
  OR2_X1 U7298 ( .A1(n6058), .A2(n7034), .ZN(n5823) );
  AND2_X1 U7299 ( .A1(n5817), .A2(n5816), .ZN(n5818) );
  OR2_X1 U7300 ( .A1(n5818), .A2(n5829), .ZN(n7033) );
  OR2_X1 U7301 ( .A1(n5791), .A2(n7033), .ZN(n5822) );
  INV_X1 U7302 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5819) );
  OR2_X1 U7303 ( .A1(n5784), .A2(n5819), .ZN(n5821) );
  NAND2_X1 U7304 ( .A1(n5789), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5820) );
  NAND4_X1 U7305 ( .A1(n5823), .A2(n5822), .A3(n5821), .A4(n5820), .ZN(n9124)
         );
  INV_X1 U7306 ( .A(n9124), .ZN(n9638) );
  OR2_X1 U7307 ( .A1(n7036), .A2(n9638), .ZN(n8311) );
  AND2_X1 U7308 ( .A1(n8311), .A2(n7022), .ZN(n8318) );
  AND2_X1 U7309 ( .A1(n7036), .A2(n9638), .ZN(n6116) );
  NAND2_X1 U7310 ( .A1(n6489), .A2(n8139), .ZN(n5827) );
  NAND2_X1 U7311 ( .A1(n5824), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5825) );
  XNOR2_X1 U7312 ( .A(n5825), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6490) );
  AOI22_X1 U7313 ( .A1(n5797), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6387), .B2(
        n6490), .ZN(n5826) );
  NAND2_X1 U7314 ( .A1(n5827), .A2(n5826), .ZN(n9631) );
  INV_X1 U7315 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5828) );
  OR2_X1 U7316 ( .A1(n6058), .A2(n5828), .ZN(n5834) );
  NAND2_X1 U7317 ( .A1(n5829), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5851) );
  OR2_X1 U7318 ( .A1(n5829), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5830) );
  NAND2_X1 U7319 ( .A1(n5851), .A2(n5830), .ZN(n9628) );
  OR2_X1 U7320 ( .A1(n5791), .A2(n9628), .ZN(n5833) );
  NAND2_X1 U7321 ( .A1(n5789), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5832) );
  NAND2_X1 U7322 ( .A1(n5790), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5831) );
  NAND4_X1 U7323 ( .A1(n5834), .A2(n5833), .A3(n5832), .A4(n5831), .ZN(n9123)
         );
  INV_X1 U7324 ( .A(n9123), .ZN(n7027) );
  NAND2_X1 U7325 ( .A1(n9631), .A2(n7027), .ZN(n8302) );
  NAND2_X1 U7326 ( .A1(n8152), .A2(n8302), .ZN(n5835) );
  OR2_X1 U7327 ( .A1(n9631), .A2(n7027), .ZN(n8158) );
  NAND2_X1 U7328 ( .A1(n5835), .A2(n8158), .ZN(n7297) );
  NAND2_X1 U7329 ( .A1(n6508), .A2(n8139), .ZN(n5839) );
  NOR2_X1 U7330 ( .A1(n5824), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5846) );
  AND2_X1 U7331 ( .A1(n5846), .A2(n5836), .ZN(n5862) );
  OR2_X1 U7332 ( .A1(n5862), .A2(n8006), .ZN(n5837) );
  XNOR2_X1 U7333 ( .A(n5837), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6603) );
  AOI22_X1 U7334 ( .A1(n5797), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6387), .B2(
        n6603), .ZN(n5838) );
  INV_X1 U7335 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5850) );
  INV_X1 U7336 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6598) );
  NAND2_X1 U7337 ( .A1(n5853), .A2(n6598), .ZN(n5840) );
  NAND2_X1 U7338 ( .A1(n5871), .A2(n5840), .ZN(n7353) );
  OR2_X1 U7339 ( .A1(n5791), .A2(n7353), .ZN(n5845) );
  INV_X1 U7340 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7305) );
  OR2_X1 U7341 ( .A1(n6058), .A2(n7305), .ZN(n5844) );
  INV_X1 U7342 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n5841) );
  OR2_X1 U7343 ( .A1(n5784), .A2(n5841), .ZN(n5843) );
  NAND2_X1 U7344 ( .A1(n5789), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5842) );
  NAND4_X1 U7345 ( .A1(n5845), .A2(n5844), .A3(n5843), .A4(n5842), .ZN(n9121)
         );
  INV_X1 U7346 ( .A(n9121), .ZN(n7434) );
  OR2_X1 U7347 ( .A1(n9479), .A2(n7434), .ZN(n5858) );
  NAND2_X1 U7348 ( .A1(n6494), .A2(n8139), .ZN(n5849) );
  OR2_X1 U7349 ( .A1(n5846), .A2(n8006), .ZN(n5847) );
  XNOR2_X1 U7350 ( .A(n5847), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6448) );
  AOI22_X1 U7351 ( .A1(n5797), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6387), .B2(
        n6448), .ZN(n5848) );
  NAND2_X1 U7352 ( .A1(n5849), .A2(n5848), .ZN(n7315) );
  INV_X1 U7353 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6427) );
  OR2_X1 U7354 ( .A1(n5784), .A2(n6427), .ZN(n5857) );
  NAND2_X1 U7355 ( .A1(n5851), .A2(n5850), .ZN(n5852) );
  NAND2_X1 U7356 ( .A1(n5853), .A2(n5852), .ZN(n7289) );
  OR2_X1 U7357 ( .A1(n5791), .A2(n7289), .ZN(n5856) );
  NAND2_X1 U7358 ( .A1(n5789), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5855) );
  NAND2_X1 U7359 ( .A1(n6041), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5854) );
  NAND4_X1 U7360 ( .A1(n5857), .A2(n5856), .A3(n5855), .A4(n5854), .ZN(n9122)
         );
  INV_X1 U7361 ( .A(n9122), .ZN(n9637) );
  OR2_X1 U7362 ( .A1(n7315), .A2(n9637), .ZN(n7295) );
  AND2_X1 U7363 ( .A1(n5858), .A2(n7295), .ZN(n8164) );
  INV_X1 U7364 ( .A(n8164), .ZN(n8154) );
  NAND2_X1 U7365 ( .A1(n9479), .A2(n7434), .ZN(n8162) );
  NAND2_X1 U7366 ( .A1(n7315), .A2(n9637), .ZN(n8160) );
  NAND2_X1 U7367 ( .A1(n8162), .A2(n8160), .ZN(n5859) );
  NAND2_X1 U7368 ( .A1(n5859), .A2(n5858), .ZN(n8303) );
  INV_X1 U7369 ( .A(n8303), .ZN(n5860) );
  NAND2_X1 U7370 ( .A1(n6513), .A2(n8139), .ZN(n5869) );
  INV_X1 U7371 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5861) );
  AND2_X1 U7372 ( .A1(n5862), .A2(n5861), .ZN(n5865) );
  NOR2_X1 U7373 ( .A1(n5865), .A2(n8006), .ZN(n5863) );
  MUX2_X1 U7374 ( .A(n8006), .B(n5863), .S(P1_IR_REG_11__SCAN_IN), .Z(n5867)
         );
  NAND2_X1 U7375 ( .A1(n5865), .A2(n5864), .ZN(n5877) );
  INV_X1 U7376 ( .A(n5877), .ZN(n5866) );
  NOR2_X1 U7377 ( .A1(n5867), .A2(n5866), .ZN(n6515) );
  AOI22_X1 U7378 ( .A1(n5797), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6387), .B2(
        n6515), .ZN(n5868) );
  NAND2_X1 U7379 ( .A1(n5869), .A2(n5868), .ZN(n7430) );
  INV_X1 U7380 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6428) );
  OR2_X1 U7381 ( .A1(n5784), .A2(n6428), .ZN(n5876) );
  INV_X1 U7382 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5870) );
  AND2_X1 U7383 ( .A1(n5871), .A2(n5870), .ZN(n5872) );
  OR2_X1 U7384 ( .A1(n5872), .A2(n5881), .ZN(n7435) );
  OR2_X1 U7385 ( .A1(n5791), .A2(n7435), .ZN(n5875) );
  INV_X1 U7386 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7368) );
  OR2_X1 U7387 ( .A1(n6058), .A2(n7368), .ZN(n5874) );
  NAND2_X1 U7388 ( .A1(n5789), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5873) );
  NAND4_X1 U7389 ( .A1(n5876), .A2(n5875), .A3(n5874), .A4(n5873), .ZN(n9527)
         );
  INV_X1 U7390 ( .A(n9527), .ZN(n7671) );
  NAND2_X1 U7391 ( .A1(n7430), .A2(n7671), .ZN(n8175) );
  NAND2_X1 U7392 ( .A1(n6528), .A2(n8139), .ZN(n5880) );
  NAND2_X1 U7393 ( .A1(n5877), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5878) );
  XNOR2_X1 U7394 ( .A(n5878), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6833) );
  AOI22_X1 U7395 ( .A1(n5797), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6387), .B2(
        n6833), .ZN(n5879) );
  INV_X1 U7396 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6429) );
  OR2_X1 U7397 ( .A1(n5784), .A2(n6429), .ZN(n5886) );
  NOR2_X1 U7398 ( .A1(n5881), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5882) );
  OR2_X1 U7399 ( .A1(n5892), .A2(n5882), .ZN(n9529) );
  OR2_X1 U7400 ( .A1(n5791), .A2(n9529), .ZN(n5885) );
  NAND2_X1 U7401 ( .A1(n5789), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5884) );
  NAND2_X1 U7402 ( .A1(n6041), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5883) );
  NAND4_X1 U7403 ( .A1(n5886), .A2(n5885), .A3(n5884), .A4(n5883), .ZN(n9120)
         );
  INV_X1 U7404 ( .A(n9120), .ZN(n7658) );
  NOR2_X1 U7405 ( .A1(n9532), .A2(n7658), .ZN(n8156) );
  INV_X1 U7406 ( .A(n8156), .ZN(n8177) );
  OR2_X1 U7407 ( .A1(n7430), .A2(n7671), .ZN(n9520) );
  NAND2_X1 U7408 ( .A1(n8177), .A2(n9520), .ZN(n8166) );
  INV_X1 U7409 ( .A(n8166), .ZN(n5887) );
  NAND2_X1 U7410 ( .A1(n9532), .A2(n7658), .ZN(n8176) );
  NAND2_X1 U7411 ( .A1(n5888), .A2(n8176), .ZN(n7413) );
  NAND2_X1 U7412 ( .A1(n6787), .A2(n8139), .ZN(n5891) );
  XNOR2_X1 U7413 ( .A(n5889), .B(P1_IR_REG_13__SCAN_IN), .ZN(n6925) );
  AOI22_X1 U7414 ( .A1(n5797), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6387), .B2(
        n6925), .ZN(n5890) );
  INV_X1 U7415 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6413) );
  OR2_X1 U7416 ( .A1(n5784), .A2(n6413), .ZN(n5897) );
  NOR2_X1 U7417 ( .A1(n5892), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5893) );
  OR2_X1 U7418 ( .A1(n5902), .A2(n5893), .ZN(n7703) );
  OR2_X1 U7419 ( .A1(n5791), .A2(n7703), .ZN(n5896) );
  INV_X1 U7420 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7418) );
  OR2_X1 U7421 ( .A1(n6058), .A2(n7418), .ZN(n5895) );
  NAND2_X1 U7422 ( .A1(n5789), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5894) );
  NAND4_X1 U7423 ( .A1(n5897), .A2(n5896), .A3(n5895), .A4(n5894), .ZN(n9525)
         );
  INV_X1 U7424 ( .A(n9525), .ZN(n7700) );
  OR2_X1 U7425 ( .A1(n7706), .A2(n7700), .ZN(n8168) );
  NAND2_X1 U7426 ( .A1(n7706), .A2(n7700), .ZN(n8169) );
  NAND2_X1 U7427 ( .A1(n8168), .A2(n8169), .ZN(n8266) );
  INV_X1 U7428 ( .A(n8266), .ZN(n7411) );
  NAND2_X1 U7429 ( .A1(n7413), .A2(n7411), .ZN(n5898) );
  NAND2_X1 U7430 ( .A1(n5898), .A2(n8169), .ZN(n7471) );
  INV_X1 U7431 ( .A(n7471), .ZN(n5909) );
  NAND2_X1 U7432 ( .A1(n6804), .A2(n8139), .ZN(n5901) );
  OR2_X1 U7433 ( .A1(n5899), .A2(n8006), .ZN(n5910) );
  XNOR2_X1 U7434 ( .A(n5910), .B(P1_IR_REG_14__SCAN_IN), .ZN(n6430) );
  AOI22_X1 U7435 ( .A1(n5797), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6387), .B2(
        n6430), .ZN(n5900) );
  INV_X1 U7436 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6412) );
  OR2_X1 U7437 ( .A1(n5784), .A2(n6412), .ZN(n5907) );
  NAND2_X1 U7438 ( .A1(n5789), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5906) );
  OR2_X1 U7439 ( .A1(n5902), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5903) );
  AND2_X1 U7440 ( .A1(n5903), .A2(n5918), .ZN(n7765) );
  NAND2_X1 U7441 ( .A1(n5948), .A2(n7765), .ZN(n5905) );
  NAND2_X1 U7442 ( .A1(n6041), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5904) );
  NAND4_X1 U7443 ( .A1(n5907), .A2(n5906), .A3(n5905), .A4(n5904), .ZN(n9119)
         );
  INV_X1 U7444 ( .A(n9119), .ZN(n7762) );
  NOR2_X1 U7445 ( .A1(n7769), .A2(n7762), .ZN(n8171) );
  INV_X1 U7446 ( .A(n8171), .ZN(n8293) );
  NAND2_X1 U7447 ( .A1(n7769), .A2(n7762), .ZN(n8170) );
  NAND2_X1 U7448 ( .A1(n8293), .A2(n8170), .ZN(n8267) );
  NAND2_X1 U7449 ( .A1(n5909), .A2(n5908), .ZN(n7473) );
  NAND2_X1 U7450 ( .A1(n6837), .A2(n8139), .ZN(n5916) );
  NAND2_X1 U7451 ( .A1(n5910), .A2(n10119), .ZN(n5911) );
  NAND2_X1 U7452 ( .A1(n5911), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5913) );
  XNOR2_X1 U7453 ( .A(n5913), .B(n5912), .ZN(n7611) );
  INV_X1 U7454 ( .A(n7611), .ZN(n5914) );
  AOI22_X1 U7455 ( .A1(n5797), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6387), .B2(
        n5914), .ZN(n5915) );
  NAND2_X1 U7456 ( .A1(n5790), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5923) );
  INV_X1 U7457 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5917) );
  NAND2_X1 U7458 ( .A1(n5918), .A2(n5917), .ZN(n5919) );
  AND2_X1 U7459 ( .A1(n5928), .A2(n5919), .ZN(n7911) );
  NAND2_X1 U7460 ( .A1(n5948), .A2(n7911), .ZN(n5922) );
  NAND2_X1 U7461 ( .A1(n5789), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5921) );
  NAND2_X1 U7462 ( .A1(n6041), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5920) );
  NAND4_X1 U7463 ( .A1(n5923), .A2(n5922), .A3(n5921), .A4(n5920), .ZN(n9503)
         );
  INV_X1 U7464 ( .A(n9503), .ZN(n7975) );
  OR2_X1 U7465 ( .A1(n7908), .A2(n7975), .ZN(n8297) );
  NAND2_X1 U7466 ( .A1(n7908), .A2(n7975), .ZN(n8295) );
  NAND2_X1 U7467 ( .A1(n6841), .A2(n8139), .ZN(n5927) );
  NAND2_X1 U7468 ( .A1(n5924), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5925) );
  XNOR2_X1 U7469 ( .A(n5925), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7805) );
  AOI22_X1 U7470 ( .A1(n5797), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6387), .B2(
        n7805), .ZN(n5926) );
  NAND2_X2 U7471 ( .A1(n5927), .A2(n5926), .ZN(n9549) );
  INV_X1 U7472 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n10111) );
  AND2_X1 U7473 ( .A1(n5928), .A2(n10111), .ZN(n5929) );
  OR2_X1 U7474 ( .A1(n5929), .A2(n5936), .ZN(n9507) );
  AOI22_X1 U7475 ( .A1(n5790), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n5789), .B2(
        P1_REG0_REG_16__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U7476 ( .A1(n6041), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5930) );
  OAI211_X1 U7477 ( .C1(n9507), .C2(n5791), .A(n5931), .B(n5930), .ZN(n9118)
         );
  NAND2_X1 U7478 ( .A1(n9549), .A2(n9118), .ZN(n8183) );
  OR2_X1 U7479 ( .A1(n9549), .A2(n9118), .ZN(n5932) );
  INV_X1 U7480 ( .A(n9118), .ZN(n9046) );
  AND2_X1 U7481 ( .A1(n9549), .A2(n9046), .ZN(n8284) );
  NAND2_X1 U7482 ( .A1(n6902), .A2(n8139), .ZN(n5935) );
  NAND2_X1 U7483 ( .A1(n5933), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5941) );
  XNOR2_X1 U7484 ( .A(n5941), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9163) );
  AOI22_X1 U7485 ( .A1(n5797), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6387), .B2(
        n9163), .ZN(n5934) );
  NOR2_X1 U7486 ( .A1(n5936), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5937) );
  OR2_X1 U7487 ( .A1(n5946), .A2(n5937), .ZN(n9048) );
  AOI22_X1 U7488 ( .A1(n5790), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n5789), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n5939) );
  NAND2_X1 U7489 ( .A1(n6041), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5938) );
  OAI211_X1 U7490 ( .C1(n9048), .C2(n5791), .A(n5939), .B(n5938), .ZN(n9504)
         );
  INV_X1 U7491 ( .A(n9504), .ZN(n9362) );
  NAND2_X1 U7492 ( .A1(n9440), .A2(n9362), .ZN(n8192) );
  NAND2_X1 U7493 ( .A1(n7892), .A2(n8192), .ZN(n9358) );
  NAND2_X1 U7494 ( .A1(n6931), .A2(n8139), .ZN(n5945) );
  INV_X1 U7495 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U7496 ( .A1(n5941), .A2(n5940), .ZN(n5942) );
  NAND2_X1 U7497 ( .A1(n5942), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5943) );
  XNOR2_X1 U7498 ( .A(n5943), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9175) );
  AOI22_X1 U7499 ( .A1(n5797), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9175), .B2(
        n6387), .ZN(n5944) );
  OR2_X1 U7500 ( .A1(n5946), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5947) );
  AND2_X1 U7501 ( .A1(n5947), .A2(n5957), .ZN(n9367) );
  NAND2_X1 U7502 ( .A1(n9367), .A2(n5948), .ZN(n5953) );
  INV_X1 U7503 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9156) );
  NAND2_X1 U7504 ( .A1(n5789), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5950) );
  INV_X1 U7505 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n10171) );
  OR2_X1 U7506 ( .A1(n6058), .A2(n10171), .ZN(n5949) );
  OAI211_X1 U7507 ( .C1(n9156), .C2(n5784), .A(n5950), .B(n5949), .ZN(n5951)
         );
  INV_X1 U7508 ( .A(n5951), .ZN(n5952) );
  NAND2_X1 U7509 ( .A1(n5953), .A2(n5952), .ZN(n9346) );
  INV_X1 U7510 ( .A(n9346), .ZN(n9047) );
  OR2_X1 U7511 ( .A1(n9435), .A2(n9047), .ZN(n8195) );
  OR2_X1 U7512 ( .A1(n9440), .A2(n9362), .ZN(n9357) );
  AND2_X1 U7513 ( .A1(n8195), .A2(n9357), .ZN(n8333) );
  NAND2_X1 U7514 ( .A1(n9435), .A2(n9047), .ZN(n9341) );
  INV_X1 U7515 ( .A(n9341), .ZN(n5963) );
  NAND2_X1 U7516 ( .A1(n7014), .A2(n8139), .ZN(n5956) );
  AOI22_X1 U7517 ( .A1(n5797), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n4486), .B2(
        n6387), .ZN(n5955) );
  NAND2_X2 U7518 ( .A1(n5956), .A2(n5955), .ZN(n9429) );
  INV_X1 U7519 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9176) );
  OR2_X1 U7520 ( .A1(n5784), .A2(n9176), .ZN(n5962) );
  OAI21_X1 U7521 ( .B1(P1_REG3_REG_19__SCAN_IN), .B2(n5958), .A(n5967), .ZN(
        n9352) );
  OR2_X1 U7522 ( .A1(n5791), .A2(n9352), .ZN(n5961) );
  INV_X1 U7523 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9173) );
  OR2_X1 U7524 ( .A1(n6058), .A2(n9173), .ZN(n5960) );
  NAND2_X1 U7525 ( .A1(n5789), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5959) );
  NAND4_X1 U7526 ( .A1(n5962), .A2(n5961), .A3(n5960), .A4(n5959), .ZN(n9332)
         );
  INV_X1 U7527 ( .A(n9332), .ZN(n9363) );
  OR2_X1 U7528 ( .A1(n9429), .A2(n9363), .ZN(n8196) );
  NAND2_X1 U7529 ( .A1(n9429), .A2(n9363), .ZN(n8326) );
  NAND2_X1 U7530 ( .A1(n8196), .A2(n8326), .ZN(n9342) );
  INV_X1 U7531 ( .A(n9342), .ZN(n9339) );
  NAND2_X1 U7532 ( .A1(n7122), .A2(n8139), .ZN(n5966) );
  OR2_X1 U7533 ( .A1(n4387), .A2(n7123), .ZN(n5965) );
  INV_X1 U7534 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10152) );
  OR2_X1 U7535 ( .A1(n5784), .A2(n10152), .ZN(n5973) );
  INV_X1 U7536 ( .A(n5967), .ZN(n5969) );
  INV_X1 U7537 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n10029) );
  INV_X1 U7538 ( .A(n5976), .ZN(n5968) );
  OAI21_X1 U7539 ( .B1(P1_REG3_REG_20__SCAN_IN), .B2(n5969), .A(n5968), .ZN(
        n9326) );
  OR2_X1 U7540 ( .A1(n5791), .A2(n9326), .ZN(n5972) );
  NAND2_X1 U7541 ( .A1(n5789), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5971) );
  NAND2_X1 U7542 ( .A1(n6041), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5970) );
  NAND4_X1 U7543 ( .A1(n5973), .A2(n5972), .A3(n5971), .A4(n5970), .ZN(n9347)
         );
  INV_X1 U7544 ( .A(n9347), .ZN(n9318) );
  NAND2_X1 U7545 ( .A1(n9423), .A2(n9318), .ZN(n8249) );
  INV_X1 U7546 ( .A(n8249), .ZN(n8200) );
  NAND2_X1 U7547 ( .A1(n7251), .A2(n8139), .ZN(n5975) );
  INV_X1 U7548 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7311) );
  OR2_X1 U7549 ( .A1(n4387), .A2(n7311), .ZN(n5974) );
  OAI21_X1 U7550 ( .B1(P1_REG3_REG_21__SCAN_IN), .B2(n5976), .A(n5986), .ZN(
        n9310) );
  OR2_X1 U7551 ( .A1(n5791), .A2(n9310), .ZN(n5980) );
  INV_X1 U7552 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9311) );
  OR2_X1 U7553 ( .A1(n6058), .A2(n9311), .ZN(n5979) );
  NAND2_X1 U7554 ( .A1(n5789), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5978) );
  NAND2_X1 U7555 ( .A1(n5790), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5977) );
  NAND4_X1 U7556 ( .A1(n5980), .A2(n5979), .A3(n5978), .A4(n5977), .ZN(n9333)
         );
  NAND2_X1 U7557 ( .A1(n9420), .A2(n9083), .ZN(n8201) );
  INV_X1 U7558 ( .A(n9306), .ZN(n9316) );
  INV_X1 U7559 ( .A(n8201), .ZN(n5981) );
  NAND2_X1 U7560 ( .A1(n7406), .A2(n8139), .ZN(n5983) );
  OR2_X1 U7561 ( .A1(n4387), .A2(n8420), .ZN(n5982) );
  NAND2_X1 U7562 ( .A1(n5790), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5992) );
  INV_X1 U7563 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n5984) );
  OR2_X1 U7564 ( .A1(n6056), .A2(n5984), .ZN(n5991) );
  INV_X1 U7565 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9955) );
  NAND2_X1 U7566 ( .A1(n9955), .A2(n5986), .ZN(n5987) );
  NAND2_X1 U7567 ( .A1(n6002), .A2(n5987), .ZN(n9296) );
  OR2_X1 U7568 ( .A1(n5791), .A2(n9296), .ZN(n5990) );
  INV_X1 U7569 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n5988) );
  OR2_X1 U7570 ( .A1(n6058), .A2(n5988), .ZN(n5989) );
  OR2_X1 U7571 ( .A1(n9413), .A2(n9319), .ZN(n8336) );
  AND2_X1 U7572 ( .A1(n9413), .A2(n9319), .ZN(n8247) );
  INV_X1 U7573 ( .A(n8247), .ZN(n8203) );
  NAND2_X1 U7574 ( .A1(n7454), .A2(n8139), .ZN(n5994) );
  OR2_X1 U7575 ( .A1(n4387), .A2(n7457), .ZN(n5993) );
  NAND2_X1 U7576 ( .A1(n5789), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5998) );
  INV_X1 U7577 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9013) );
  XNOR2_X1 U7578 ( .A(n6002), .B(n9013), .ZN(n9280) );
  OR2_X1 U7579 ( .A1(n5791), .A2(n9280), .ZN(n5997) );
  NAND2_X1 U7580 ( .A1(n6041), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5996) );
  NAND2_X1 U7581 ( .A1(n5790), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5995) );
  NAND4_X1 U7582 ( .A1(n5998), .A2(n5997), .A3(n5996), .A4(n5995), .ZN(n9905)
         );
  NAND2_X1 U7583 ( .A1(n7458), .A2(n8139), .ZN(n6001) );
  INV_X1 U7584 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7459) );
  OR2_X1 U7585 ( .A1(n4387), .A2(n7459), .ZN(n6000) );
  INV_X1 U7586 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9055) );
  OAI21_X1 U7587 ( .B1(n6002), .B2(n9013), .A(n9055), .ZN(n6005) );
  AND2_X1 U7588 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(P1_REG3_REG_24__SCAN_IN), 
        .ZN(n6003) );
  NAND2_X1 U7589 ( .A1(n6005), .A2(n6013), .ZN(n9273) );
  OR2_X1 U7590 ( .A1(n5791), .A2(n9273), .ZN(n6009) );
  INV_X1 U7591 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n10089) );
  OR2_X1 U7592 ( .A1(n6058), .A2(n10089), .ZN(n6008) );
  NAND2_X1 U7593 ( .A1(n5790), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7594 ( .A1(n5789), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6006) );
  NAND4_X1 U7595 ( .A1(n6009), .A2(n6008), .A3(n6007), .A4(n6006), .ZN(n9286)
         );
  INV_X1 U7596 ( .A(n9286), .ZN(n9034) );
  OR2_X1 U7597 ( .A1(n9405), .A2(n9034), .ZN(n8394) );
  NAND2_X1 U7598 ( .A1(n9405), .A2(n9034), .ZN(n9255) );
  NAND2_X1 U7599 ( .A1(n8394), .A2(n9255), .ZN(n9266) );
  NAND2_X1 U7600 ( .A1(n7535), .A2(n8139), .ZN(n6011) );
  OR2_X1 U7601 ( .A1(n4387), .A2(n9958), .ZN(n6010) );
  NAND2_X1 U7602 ( .A1(n5789), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6018) );
  INV_X1 U7603 ( .A(n6013), .ZN(n6012) );
  NAND2_X1 U7604 ( .A1(n6012), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6021) );
  INV_X1 U7605 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9035) );
  NAND2_X1 U7606 ( .A1(n6013), .A2(n9035), .ZN(n6014) );
  NAND2_X1 U7607 ( .A1(n6021), .A2(n6014), .ZN(n9251) );
  OR2_X1 U7608 ( .A1(n5791), .A2(n9251), .ZN(n6017) );
  NAND2_X1 U7609 ( .A1(n6041), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U7610 ( .A1(n5790), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6015) );
  NAND4_X1 U7611 ( .A1(n6018), .A2(n6017), .A3(n6016), .A4(n6015), .ZN(n9243)
         );
  NAND2_X1 U7612 ( .A1(n9398), .A2(n9268), .ZN(n8398) );
  NAND2_X1 U7613 ( .A1(n8398), .A2(n9255), .ZN(n8343) );
  NOR2_X1 U7614 ( .A1(n9398), .A2(n9268), .ZN(n8209) );
  NAND2_X1 U7615 ( .A1(n7532), .A2(n8139), .ZN(n6020) );
  OR2_X1 U7616 ( .A1(n4387), .A2(n7533), .ZN(n6019) );
  INV_X1 U7617 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9109) );
  NAND2_X1 U7618 ( .A1(n6021), .A2(n9109), .ZN(n6022) );
  NAND2_X1 U7619 ( .A1(n6030), .A2(n6022), .ZN(n9237) );
  OR2_X1 U7620 ( .A1(n5791), .A2(n9237), .ZN(n6027) );
  INV_X1 U7621 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n6023) );
  OR2_X1 U7622 ( .A1(n6058), .A2(n6023), .ZN(n6026) );
  NAND2_X1 U7623 ( .A1(n5790), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6025) );
  NAND2_X1 U7624 ( .A1(n5789), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6024) );
  NAND4_X1 U7625 ( .A1(n6027), .A2(n6026), .A3(n6025), .A4(n6024), .ZN(n9259)
         );
  OR2_X1 U7626 ( .A1(n4387), .A2(n7603), .ZN(n6028) );
  INV_X1 U7627 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10138) );
  OR2_X1 U7628 ( .A1(n5784), .A2(n10138), .ZN(n6036) );
  INV_X1 U7629 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9005) );
  NAND2_X1 U7630 ( .A1(n6030), .A2(n9005), .ZN(n6031) );
  NAND2_X1 U7631 ( .A1(n6039), .A2(n6031), .ZN(n9222) );
  OR2_X1 U7632 ( .A1(n5791), .A2(n9222), .ZN(n6035) );
  INV_X1 U7633 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6032) );
  OR2_X1 U7634 ( .A1(n6058), .A2(n6032), .ZN(n6034) );
  NAND2_X1 U7635 ( .A1(n5789), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6033) );
  NAND4_X1 U7636 ( .A1(n6036), .A2(n6035), .A3(n6034), .A4(n6033), .ZN(n9244)
         );
  NAND2_X1 U7637 ( .A1(n9388), .A2(n9107), .ZN(n8348) );
  NOR2_X2 U7638 ( .A1(n9226), .A2(n9227), .ZN(n9225) );
  NOR2_X1 U7639 ( .A1(n9225), .A2(n8351), .ZN(n9210) );
  NAND2_X1 U7640 ( .A1(n8457), .A2(n8139), .ZN(n6038) );
  OR2_X1 U7641 ( .A1(n4387), .A2(n7713), .ZN(n6037) );
  INV_X1 U7642 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n10154) );
  OR2_X1 U7643 ( .A1(n5784), .A2(n10154), .ZN(n6045) );
  INV_X1 U7644 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8119) );
  NAND2_X1 U7645 ( .A1(n6039), .A2(n8119), .ZN(n6040) );
  NAND2_X1 U7646 ( .A1(n6151), .A2(n6040), .ZN(n9205) );
  OR2_X1 U7647 ( .A1(n5791), .A2(n9205), .ZN(n6044) );
  NAND2_X1 U7648 ( .A1(n5789), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U7649 ( .A1(n6041), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6042) );
  NAND4_X1 U7650 ( .A1(n6045), .A2(n6044), .A3(n6043), .A4(n6042), .ZN(n9117)
         );
  NOR2_X1 U7651 ( .A1(n9383), .A2(n9229), .ZN(n8224) );
  INV_X1 U7652 ( .A(n8224), .ZN(n8281) );
  NAND2_X1 U7653 ( .A1(n9210), .A2(n9211), .ZN(n9209) );
  NAND2_X1 U7654 ( .A1(n9209), .A2(n8349), .ZN(n6064) );
  INV_X1 U7655 ( .A(SI_28_), .ZN(n6048) );
  NAND2_X1 U7656 ( .A1(n6049), .A2(n6048), .ZN(n6050) );
  INV_X1 U7657 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n10131) );
  INV_X1 U7658 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7798) );
  MUX2_X1 U7659 ( .A(n10131), .B(n7798), .S(n4749), .Z(n6184) );
  XNOR2_X1 U7660 ( .A(n6184), .B(SI_29_), .ZN(n6052) );
  NAND2_X1 U7661 ( .A1(n7797), .A2(n8139), .ZN(n6054) );
  OR2_X1 U7662 ( .A1(n4387), .A2(n7798), .ZN(n6053) );
  NAND2_X1 U7663 ( .A1(n5790), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6062) );
  INV_X1 U7664 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6055) );
  OR2_X1 U7665 ( .A1(n6056), .A2(n6055), .ZN(n6061) );
  OR2_X1 U7666 ( .A1(n5791), .A2(n6151), .ZN(n6060) );
  INV_X1 U7667 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n6057) );
  OR2_X1 U7668 ( .A1(n6058), .A2(n6057), .ZN(n6059) );
  NOR2_X1 U7669 ( .A1(n9380), .A2(n8230), .ZN(n8280) );
  INV_X1 U7670 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n6067) );
  NAND2_X1 U7671 ( .A1(n5789), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6066) );
  NAND2_X1 U7672 ( .A1(n5790), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6065) );
  OAI211_X1 U7673 ( .C1(n6058), .C2(n6067), .A(n6066), .B(n6065), .ZN(n9116)
         );
  INV_X1 U7674 ( .A(n9116), .ZN(n6072) );
  INV_X1 U7675 ( .A(n7312), .ZN(n8367) );
  NAND2_X1 U7676 ( .A1(n6146), .A2(n8367), .ZN(n8279) );
  INV_X1 U7677 ( .A(n6068), .ZN(n6729) );
  INV_X1 U7678 ( .A(P1_B_REG_SCAN_IN), .ZN(n6069) );
  NOR2_X1 U7679 ( .A1(n8412), .A2(n6069), .ZN(n6070) );
  NOR2_X1 U7680 ( .A1(n9662), .A2(n6070), .ZN(n9189) );
  INV_X1 U7681 ( .A(n9189), .ZN(n6071) );
  OR2_X1 U7682 ( .A1(n8279), .A2(n6716), .ZN(n6774) );
  NAND2_X1 U7683 ( .A1(n6073), .A2(n6083), .ZN(n6076) );
  INV_X1 U7684 ( .A(n6076), .ZN(n6074) );
  NAND2_X1 U7685 ( .A1(n6074), .A2(n5728), .ZN(n6079) );
  NAND2_X1 U7686 ( .A1(n6079), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6075) );
  XNOR2_X1 U7687 ( .A(n6075), .B(P1_IR_REG_25__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7688 ( .A1(n6076), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6077) );
  MUX2_X1 U7689 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6077), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n6078) );
  AND2_X1 U7690 ( .A1(n6078), .A2(n6079), .ZN(n6087) );
  INV_X1 U7691 ( .A(n6073), .ZN(n6082) );
  NAND2_X1 U7692 ( .A1(n6082), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6084) );
  XNOR2_X1 U7693 ( .A(n6084), .B(n6083), .ZN(n6772) );
  AND2_X1 U7694 ( .A1(n6772), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6085) );
  AND2_X1 U7695 ( .A1(n6773), .A2(n6085), .ZN(n6722) );
  INV_X1 U7696 ( .A(n6086), .ZN(n7538) );
  NAND2_X1 U7697 ( .A1(n7538), .A2(P1_B_REG_SCAN_IN), .ZN(n6088) );
  INV_X1 U7698 ( .A(n6087), .ZN(n7460) );
  MUX2_X1 U7699 ( .A(P1_B_REG_SCAN_IN), .B(n6088), .S(n7460), .Z(n6089) );
  NAND2_X1 U7700 ( .A1(n6089), .A2(n6090), .ZN(n6536) );
  INV_X1 U7701 ( .A(n6090), .ZN(n7534) );
  NAND2_X1 U7702 ( .A1(n7534), .A2(n7460), .ZN(n6534) );
  OAI21_X1 U7703 ( .B1(n6536), .B2(P1_D_REG_0__SCAN_IN), .A(n6534), .ZN(n6102)
         );
  INV_X1 U7704 ( .A(n6536), .ZN(n6100) );
  NOR4_X1 U7705 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n10126) );
  NOR2_X1 U7706 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .ZN(
        n6093) );
  NOR4_X1 U7707 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6092) );
  NOR4_X1 U7708 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n6091) );
  AND4_X1 U7709 ( .A1(n10126), .A2(n6093), .A3(n6092), .A4(n6091), .ZN(n6099)
         );
  NOR4_X1 U7710 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n6097) );
  NOR4_X1 U7711 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6096) );
  NOR4_X1 U7712 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6095) );
  NOR4_X1 U7713 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n6094) );
  AND4_X1 U7714 ( .A1(n6097), .A2(n6096), .A3(n6095), .A4(n6094), .ZN(n6098)
         );
  NAND2_X1 U7715 ( .A1(n6099), .A2(n6098), .ZN(n6533) );
  NAND2_X1 U7716 ( .A1(n6100), .A2(n6533), .ZN(n6101) );
  NAND2_X1 U7717 ( .A1(n6102), .A2(n6101), .ZN(n6542) );
  NAND2_X1 U7718 ( .A1(n7534), .A2(n7538), .ZN(n6482) );
  OAI21_X1 U7719 ( .B1(n6536), .B2(P1_D_REG_1__SCAN_IN), .A(n6482), .ZN(n6719)
         );
  NOR2_X1 U7720 ( .A1(n6542), .A2(n6719), .ZN(n6103) );
  NAND2_X1 U7721 ( .A1(n6726), .A2(n6103), .ZN(n7039) );
  NAND2_X1 U7722 ( .A1(n6149), .A2(n7312), .ZN(n6717) );
  NAND2_X1 U7723 ( .A1(n6722), .A2(n4486), .ZN(n6104) );
  INV_X1 U7724 ( .A(n9405), .ZN(n6148) );
  INV_X1 U7725 ( .A(n8255), .ZN(n6105) );
  INV_X1 U7726 ( .A(n7148), .ZN(n6951) );
  AND2_X1 U7727 ( .A1(n6695), .A2(n6951), .ZN(n7139) );
  NAND2_X1 U7728 ( .A1(n6105), .A2(n7139), .ZN(n7138) );
  NAND2_X1 U7729 ( .A1(n9130), .A2(n7142), .ZN(n6106) );
  NAND2_X1 U7730 ( .A1(n7138), .A2(n6106), .ZN(n7191) );
  INV_X1 U7731 ( .A(n7191), .ZN(n6107) );
  INV_X1 U7732 ( .A(n7193), .ZN(n8252) );
  NAND2_X1 U7733 ( .A1(n6107), .A2(n8252), .ZN(n7155) );
  NAND2_X1 U7734 ( .A1(n7160), .A2(n9676), .ZN(n7156) );
  NAND2_X1 U7735 ( .A1(n9659), .A2(n7186), .ZN(n6109) );
  NAND2_X1 U7736 ( .A1(n9066), .A2(n9683), .ZN(n7173) );
  AND2_X1 U7737 ( .A1(n7156), .A2(n4952), .ZN(n6108) );
  NAND2_X1 U7738 ( .A1(n7155), .A2(n6108), .ZN(n6111) );
  INV_X1 U7739 ( .A(n6109), .ZN(n6110) );
  NAND2_X1 U7740 ( .A1(n8256), .A2(n8317), .ZN(n7177) );
  INV_X1 U7741 ( .A(n4952), .ZN(n6112) );
  INV_X1 U7742 ( .A(n8316), .ZN(n6113) );
  INV_X1 U7743 ( .A(n9656), .ZN(n6114) );
  NAND2_X1 U7744 ( .A1(n9126), .A2(n9651), .ZN(n6115) );
  OAI22_X2 U7745 ( .A1(n7044), .A2(n7046), .B1(n9125), .B2(n7059), .ZN(n7032)
         );
  INV_X1 U7746 ( .A(n6116), .ZN(n8301) );
  INV_X1 U7747 ( .A(n7031), .ZN(n8258) );
  NAND2_X1 U7748 ( .A1(n7032), .A2(n8258), .ZN(n6118) );
  OR2_X1 U7749 ( .A1(n7036), .A2(n9124), .ZN(n6117) );
  NAND2_X1 U7750 ( .A1(n8158), .A2(n8302), .ZN(n8259) );
  INV_X1 U7751 ( .A(n8259), .ZN(n9633) );
  NAND2_X1 U7752 ( .A1(n9631), .A2(n9123), .ZN(n6119) );
  OR2_X1 U7753 ( .A1(n7315), .A2(n9122), .ZN(n6120) );
  XNOR2_X1 U7754 ( .A(n9479), .B(n9121), .ZN(n8261) );
  NAND2_X1 U7755 ( .A1(n7301), .A2(n6121), .ZN(n7300) );
  OR2_X1 U7756 ( .A1(n9479), .A2(n9121), .ZN(n6122) );
  NAND2_X1 U7757 ( .A1(n7300), .A2(n6122), .ZN(n7362) );
  NAND2_X1 U7758 ( .A1(n7430), .A2(n9527), .ZN(n7359) );
  NAND2_X1 U7759 ( .A1(n7362), .A2(n7359), .ZN(n6123) );
  OR2_X1 U7760 ( .A1(n7430), .A2(n9527), .ZN(n7360) );
  NAND2_X1 U7761 ( .A1(n8177), .A2(n8176), .ZN(n9522) );
  INV_X1 U7762 ( .A(n9522), .ZN(n9535) );
  OR2_X1 U7763 ( .A1(n9535), .A2(n4418), .ZN(n6124) );
  NAND2_X1 U7764 ( .A1(n9532), .A2(n9120), .ZN(n7410) );
  NAND2_X1 U7765 ( .A1(n7706), .A2(n9525), .ZN(n6125) );
  AND2_X1 U7766 ( .A1(n7410), .A2(n6125), .ZN(n6126) );
  OR2_X1 U7767 ( .A1(n4418), .A2(n6126), .ZN(n6127) );
  AND2_X1 U7768 ( .A1(n7769), .A2(n9119), .ZN(n6128) );
  NAND2_X1 U7769 ( .A1(n7908), .A2(n9503), .ZN(n6129) );
  NAND2_X1 U7770 ( .A1(n7724), .A2(n6129), .ZN(n6131) );
  OR2_X1 U7771 ( .A1(n7908), .A2(n9503), .ZN(n6130) );
  INV_X1 U7772 ( .A(n9440), .ZN(n7888) );
  NAND2_X1 U7773 ( .A1(n8195), .A2(n9341), .ZN(n9360) );
  INV_X1 U7774 ( .A(n9429), .ZN(n6135) );
  INV_X1 U7775 ( .A(n9322), .ZN(n6137) );
  INV_X1 U7776 ( .A(n9423), .ZN(n9329) );
  INV_X1 U7777 ( .A(n9420), .ZN(n9309) );
  INV_X1 U7778 ( .A(n9413), .ZN(n9299) );
  NOR2_X1 U7779 ( .A1(n9299), .A2(n9319), .ZN(n6138) );
  INV_X1 U7780 ( .A(n9319), .ZN(n9287) );
  INV_X1 U7781 ( .A(n9408), .ZN(n9283) );
  AOI21_X2 U7782 ( .B1(n6141), .B2(n6140), .A(n6139), .ZN(n9264) );
  OAI21_X1 U7783 ( .B1(n9034), .B2(n6148), .A(n9264), .ZN(n6143) );
  NAND2_X2 U7784 ( .A1(n6143), .A2(n6142), .ZN(n9249) );
  INV_X1 U7785 ( .A(n9398), .ZN(n9254) );
  INV_X1 U7786 ( .A(n9227), .ZN(n8275) );
  NOR2_X1 U7787 ( .A1(n9200), .A2(n9211), .ZN(n9199) );
  NAND2_X1 U7788 ( .A1(n6146), .A2(n9350), .ZN(n7125) );
  OR2_X1 U7789 ( .A1(n7125), .A2(n6691), .ZN(n8414) );
  AND2_X1 U7790 ( .A1(n8414), .A2(n6738), .ZN(n9664) );
  NAND2_X1 U7791 ( .A1(n9665), .A2(n9664), .ZN(n9374) );
  INV_X1 U7792 ( .A(n9383), .ZN(n9208) );
  INV_X1 U7793 ( .A(n9435), .ZN(n9371) );
  NAND2_X1 U7794 ( .A1(n9671), .A2(n7148), .ZN(n7200) );
  OR2_X1 U7795 ( .A1(n7200), .A2(n7205), .ZN(n7202) );
  NAND2_X1 U7796 ( .A1(n7183), .A2(n7186), .ZN(n9648) );
  INV_X1 U7797 ( .A(n7036), .ZN(n7037) );
  INV_X1 U7798 ( .A(n9631), .ZN(n9719) );
  NAND2_X1 U7799 ( .A1(n9627), .A2(n9719), .ZN(n9626) );
  INV_X1 U7800 ( .A(n7430), .ZN(n7461) );
  INV_X1 U7801 ( .A(n9532), .ZN(n9563) );
  INV_X1 U7802 ( .A(n7908), .ZN(n7918) );
  NAND2_X1 U7803 ( .A1(n9329), .A2(n9349), .ZN(n9323) );
  NOR2_X2 U7804 ( .A1(n9323), .A2(n9420), .ZN(n9308) );
  NAND2_X1 U7805 ( .A1(n9299), .A2(n9308), .ZN(n9293) );
  NAND2_X1 U7806 ( .A1(n9208), .A2(n9221), .ZN(n9202) );
  AOI21_X1 U7807 ( .B1(n9380), .B2(n9202), .A(n9193), .ZN(n9381) );
  NOR2_X1 U7808 ( .A1(n7126), .A2(n8367), .ZN(n6150) );
  AND2_X1 U7809 ( .A1(n9665), .A2(n6150), .ZN(n9337) );
  NAND2_X1 U7810 ( .A1(n9665), .A2(n4487), .ZN(n9370) );
  INV_X1 U7811 ( .A(n6151), .ZN(n6152) );
  INV_X1 U7812 ( .A(n9629), .ZN(n9653) );
  AOI22_X1 U7813 ( .A1(n4389), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n6152), .B2(
        n9653), .ZN(n6153) );
  OAI21_X1 U7814 ( .B1(n8236), .B2(n9370), .A(n6153), .ZN(n6154) );
  NAND2_X1 U7815 ( .A1(n8422), .A2(n8426), .ZN(n6981) );
  NAND2_X1 U7816 ( .A1(n6981), .A2(n6251), .ZN(n6247) );
  NAND2_X1 U7817 ( .A1(n6247), .A2(n6245), .ZN(n7095) );
  INV_X1 U7818 ( .A(n6159), .ZN(n6158) );
  INV_X2 U7819 ( .A(n7102), .ZN(n9811) );
  OAI21_X1 U7820 ( .B1(n7095), .B2(n7094), .A(n6252), .ZN(n6996) );
  XNOR2_X1 U7821 ( .A(n8585), .B(n7117), .ZN(n7115) );
  INV_X1 U7822 ( .A(n7115), .ZN(n7007) );
  NAND2_X1 U7823 ( .A1(n6996), .A2(n7007), .ZN(n6160) );
  INV_X1 U7824 ( .A(n8585), .ZN(n8027) );
  NAND2_X1 U7825 ( .A1(n8027), .A2(n9817), .ZN(n6235) );
  INV_X1 U7826 ( .A(n8550), .ZN(n9830) );
  NAND2_X1 U7827 ( .A1(n9830), .A2(n8584), .ZN(n7226) );
  INV_X1 U7828 ( .A(n8547), .ZN(n9773) );
  INV_X1 U7829 ( .A(n7263), .ZN(n9746) );
  NAND2_X1 U7830 ( .A1(n9773), .A2(n9746), .ZN(n6259) );
  AND2_X1 U7831 ( .A1(n6259), .A2(n7226), .ZN(n6260) );
  NAND2_X1 U7832 ( .A1(n8547), .A2(n7263), .ZN(n6238) );
  XNOR2_X1 U7833 ( .A(n9748), .B(n7332), .ZN(n9781) );
  INV_X1 U7834 ( .A(n7332), .ZN(n9785) );
  NOR2_X1 U7835 ( .A1(n9748), .A2(n9785), .ZN(n6266) );
  NAND2_X1 U7836 ( .A1(n8129), .A2(n7335), .ZN(n6270) );
  NAND2_X1 U7837 ( .A1(n7328), .A2(n6270), .ZN(n6162) );
  INV_X1 U7838 ( .A(n8129), .ZN(n9775) );
  INV_X1 U7839 ( .A(n7335), .ZN(n7490) );
  NAND2_X1 U7840 ( .A1(n9775), .A2(n7490), .ZN(n6271) );
  NAND2_X1 U7841 ( .A1(n7330), .A2(n7528), .ZN(n7496) );
  INV_X1 U7842 ( .A(n7528), .ZN(n9840) );
  NAND2_X1 U7843 ( .A1(n8583), .A2(n9840), .ZN(n6274) );
  INV_X1 U7844 ( .A(n7575), .ZN(n7517) );
  NAND2_X1 U7845 ( .A1(n7593), .A2(n6163), .ZN(n6281) );
  INV_X1 U7846 ( .A(n7492), .ZN(n6164) );
  NAND2_X1 U7847 ( .A1(n6165), .A2(n6164), .ZN(n7498) );
  NAND2_X1 U7848 ( .A1(n7498), .A2(n6281), .ZN(n7591) );
  NAND2_X1 U7849 ( .A1(n7779), .A2(n7687), .ZN(n6288) );
  NAND2_X1 U7850 ( .A1(n8975), .A2(n7788), .ZN(n6298) );
  OR2_X1 U7851 ( .A1(n7837), .A2(n7849), .ZN(n6300) );
  OR2_X1 U7852 ( .A1(n8975), .A2(n7788), .ZN(n7785) );
  AND2_X1 U7853 ( .A1(n6300), .A2(n7785), .ZN(n6294) );
  NAND2_X1 U7854 ( .A1(n7784), .A2(n6294), .ZN(n7843) );
  NAND2_X1 U7855 ( .A1(n7837), .A2(n7849), .ZN(n7846) );
  NAND2_X1 U7856 ( .A1(n9491), .A2(n7999), .ZN(n6305) );
  NAND2_X1 U7857 ( .A1(n6166), .A2(n8881), .ZN(n8875) );
  AND2_X1 U7858 ( .A1(n8863), .A2(n8875), .ZN(n7919) );
  NAND2_X1 U7859 ( .A1(n8964), .A2(n8883), .ZN(n6308) );
  INV_X1 U7860 ( .A(n6170), .ZN(n7924) );
  AND2_X1 U7861 ( .A1(n7846), .A2(n6167), .ZN(n6169) );
  OR2_X1 U7862 ( .A1(n6166), .A2(n8881), .ZN(n6296) );
  NAND2_X1 U7863 ( .A1(n6296), .A2(n8875), .ZN(n7847) );
  INV_X1 U7864 ( .A(n7847), .ZN(n7844) );
  OR2_X1 U7865 ( .A1(n6170), .A2(n7920), .ZN(n7921) );
  AND2_X1 U7866 ( .A1(n6309), .A2(n7921), .ZN(n6171) );
  NAND2_X1 U7867 ( .A1(n7922), .A2(n6171), .ZN(n7980) );
  OR2_X1 U7868 ( .A1(n8522), .A2(n8858), .ZN(n6208) );
  INV_X1 U7869 ( .A(n6208), .ZN(n6312) );
  NAND2_X1 U7870 ( .A1(n8522), .A2(n8858), .ZN(n6315) );
  NAND2_X1 U7871 ( .A1(n8960), .A2(n8830), .ZN(n6314) );
  INV_X1 U7872 ( .A(n8573), .ZN(n8859) );
  OR2_X1 U7873 ( .A1(n8953), .A2(n8859), .ZN(n6323) );
  NAND2_X1 U7874 ( .A1(n8953), .A2(n8859), .ZN(n6324) );
  NAND2_X1 U7875 ( .A1(n6323), .A2(n6324), .ZN(n8827) );
  INV_X1 U7876 ( .A(n6324), .ZN(n6172) );
  OR2_X1 U7877 ( .A1(n8949), .A2(n8831), .ZN(n6326) );
  NAND2_X1 U7878 ( .A1(n8949), .A2(n8831), .ZN(n8803) );
  NAND2_X1 U7879 ( .A1(n6326), .A2(n8803), .ZN(n8820) );
  NAND2_X1 U7880 ( .A1(n8942), .A2(n8496), .ZN(n6328) );
  NAND2_X1 U7881 ( .A1(n6331), .A2(n6328), .ZN(n8804) );
  INV_X1 U7882 ( .A(n8804), .ZN(n6173) );
  NAND2_X1 U7883 ( .A1(n6173), .A2(n8803), .ZN(n6174) );
  XNOR2_X1 U7884 ( .A(n8937), .B(n8562), .ZN(n8788) );
  NAND2_X1 U7885 ( .A1(n8937), .A2(n8562), .ZN(n6333) );
  NAND2_X1 U7886 ( .A1(n8932), .A2(n8572), .ZN(n6337) );
  INV_X1 U7887 ( .A(n6338), .ZN(n6175) );
  NAND2_X1 U7888 ( .A1(n8922), .A2(n8505), .ZN(n6343) );
  NAND2_X1 U7889 ( .A1(n8927), .A2(n8746), .ZN(n8743) );
  NAND2_X1 U7890 ( .A1(n8760), .A2(n4964), .ZN(n8741) );
  NAND2_X1 U7891 ( .A1(n8741), .A2(n6344), .ZN(n8723) );
  NAND2_X1 U7892 ( .A1(n8919), .A2(n8747), .ZN(n6227) );
  NAND2_X1 U7893 ( .A1(n8723), .A2(n8724), .ZN(n8702) );
  AND2_X1 U7894 ( .A1(n6347), .A2(n8703), .ZN(n6231) );
  NAND2_X1 U7895 ( .A1(n8702), .A2(n6231), .ZN(n8690) );
  NAND2_X1 U7896 ( .A1(n8907), .A2(n8707), .ZN(n6354) );
  NAND2_X1 U7897 ( .A1(n8690), .A2(n6176), .ZN(n8688) );
  NAND2_X1 U7898 ( .A1(n8688), .A2(n6353), .ZN(n8670) );
  NAND2_X1 U7899 ( .A1(n8902), .A2(n8442), .ZN(n6358) );
  INV_X1 U7900 ( .A(n8669), .ZN(n6356) );
  NAND2_X1 U7901 ( .A1(n7797), .A2(n6188), .ZN(n6178) );
  OR2_X1 U7902 ( .A1(n6203), .A2(n10131), .ZN(n6177) );
  OR2_X1 U7903 ( .A1(n8898), .A2(n6179), .ZN(n6361) );
  NAND2_X1 U7904 ( .A1(n8898), .A2(n6179), .ZN(n6362) );
  INV_X1 U7905 ( .A(n6362), .ZN(n6180) );
  INV_X1 U7906 ( .A(SI_29_), .ZN(n6181) );
  AND2_X1 U7907 ( .A1(n6184), .A2(n6181), .ZN(n6182) );
  INV_X1 U7908 ( .A(n6184), .ZN(n6185) );
  NAND2_X1 U7909 ( .A1(n6185), .A2(SI_29_), .ZN(n6186) );
  MUX2_X1 U7910 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n4980), .Z(n6197) );
  INV_X1 U7911 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8431) );
  NOR2_X1 U7912 ( .A1(n6203), .A2(n8431), .ZN(n6187) );
  AOI222_X1 U7913 ( .A1(n6189), .A2(P2_REG0_REG_31__SCAN_IN), .B1(n6191), .B2(
        P2_REG2_REG_31__SCAN_IN), .C1(n6190), .C2(P2_REG1_REG_31__SCAN_IN), 
        .ZN(n6206) );
  INV_X1 U7914 ( .A(n6206), .ZN(n8019) );
  INV_X1 U7915 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7916 ( .A1(n6190), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6193) );
  NAND2_X1 U7917 ( .A1(n6191), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6192) );
  OAI211_X1 U7918 ( .C1(n6195), .C2(n6194), .A(n6193), .B(n6192), .ZN(n8568)
         );
  AND2_X1 U7919 ( .A1(n8897), .A2(n8568), .ZN(n6370) );
  NAND2_X1 U7920 ( .A1(n6198), .A2(n6197), .ZN(n6199) );
  MUX2_X1 U7921 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n4980), .Z(n6201) );
  INV_X1 U7922 ( .A(SI_31_), .ZN(n6200) );
  XNOR2_X1 U7923 ( .A(n6201), .B(n6200), .ZN(n6202) );
  INV_X1 U7924 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6204) );
  INV_X1 U7925 ( .A(n8568), .ZN(n6205) );
  AND2_X1 U7926 ( .A1(n4893), .A2(n6205), .ZN(n6226) );
  NAND2_X1 U7927 ( .A1(n8890), .A2(n6206), .ZN(n6374) );
  INV_X1 U7928 ( .A(n5632), .ZN(n6375) );
  NAND2_X1 U7929 ( .A1(n6375), .A2(n6243), .ZN(n6983) );
  NOR2_X1 U7930 ( .A1(n4884), .A2(n6370), .ZN(n6366) );
  NAND2_X1 U7931 ( .A1(n6238), .A2(n6259), .ZN(n7324) );
  NOR2_X1 U7932 ( .A1(n7324), .A2(n6980), .ZN(n6212) );
  INV_X1 U7933 ( .A(n8426), .ZN(n9800) );
  NAND2_X1 U7934 ( .A1(n6209), .A2(n9800), .ZN(n6250) );
  NAND2_X1 U7935 ( .A1(n6981), .A2(n6250), .ZN(n9803) );
  NOR2_X1 U7936 ( .A1(n7094), .A2(n9803), .ZN(n6211) );
  NOR2_X1 U7937 ( .A1(n7222), .A2(n5632), .ZN(n6210) );
  AND4_X1 U7938 ( .A1(n6212), .A2(n6211), .A3(n6210), .A4(n7007), .ZN(n6213)
         );
  NAND4_X1 U7939 ( .A1(n6213), .A2(n7487), .A3(n7575), .A4(n9781), .ZN(n6214)
         );
  NAND2_X1 U7940 ( .A1(n7785), .A2(n6298), .ZN(n7873) );
  NAND2_X1 U7941 ( .A1(n6287), .A2(n6288), .ZN(n7590) );
  NOR4_X1 U7942 ( .A1(n6214), .A2(n7873), .A3(n7590), .A4(n7492), .ZN(n6215)
         );
  NAND4_X1 U7943 ( .A1(n8863), .A2(n7844), .A3(n7834), .A4(n6215), .ZN(n6216)
         );
  NOR2_X1 U7944 ( .A1(n6170), .A2(n6216), .ZN(n6217) );
  NAND3_X1 U7945 ( .A1(n4784), .A2(n7986), .A3(n6217), .ZN(n6218) );
  OR3_X1 U7946 ( .A1(n8820), .A2(n8827), .A3(n6218), .ZN(n6219) );
  NOR4_X1 U7947 ( .A1(n8775), .A2(n8788), .A3(n8804), .A4(n6219), .ZN(n6220)
         );
  NAND4_X1 U7948 ( .A1(n8724), .A2(n8742), .A3(n6220), .A4(n8761), .ZN(n6221)
         );
  NOR4_X1 U7949 ( .A1(n8669), .A2(n8681), .A3(n8704), .A4(n6221), .ZN(n6222)
         );
  NAND4_X1 U7950 ( .A1(n6366), .A2(n6367), .A3(n8448), .A4(n6222), .ZN(n6223)
         );
  XNOR2_X1 U7951 ( .A(n6223), .B(n4385), .ZN(n6225) );
  INV_X1 U7952 ( .A(n6982), .ZN(n6224) );
  AOI22_X1 U7953 ( .A1(n6225), .A2(n7252), .B1(n6224), .B2(n5632), .ZN(n6380)
         );
  INV_X1 U7954 ( .A(n6226), .ZN(n6365) );
  INV_X1 U7955 ( .A(n6227), .ZN(n6228) );
  NOR2_X1 U7956 ( .A1(n8704), .A2(n6228), .ZN(n6230) );
  AND2_X1 U7957 ( .A1(n7407), .A2(n6243), .ZN(n6229) );
  MUX2_X1 U7958 ( .A(n6231), .B(n6230), .S(n6372), .Z(n6352) );
  OAI21_X1 U7959 ( .B1(n8746), .B2(n8927), .A(n8742), .ZN(n6233) );
  NAND2_X1 U7960 ( .A1(n6343), .A2(n6372), .ZN(n6232) );
  NAND2_X1 U7961 ( .A1(n6233), .A2(n6232), .ZN(n6342) );
  AND2_X1 U7962 ( .A1(n6236), .A2(n6238), .ZN(n6234) );
  NAND2_X1 U7963 ( .A1(n6236), .A2(n6235), .ZN(n6237) );
  NAND2_X1 U7964 ( .A1(n6263), .A2(n6237), .ZN(n6241) );
  INV_X1 U7965 ( .A(n6238), .ZN(n6239) );
  NOR2_X1 U7966 ( .A1(n6239), .A2(n6266), .ZN(n6240) );
  NAND2_X1 U7967 ( .A1(n6241), .A2(n6240), .ZN(n6242) );
  NAND2_X1 U7968 ( .A1(n6242), .A2(n6372), .ZN(n6258) );
  AND2_X1 U7969 ( .A1(n6250), .A2(n6243), .ZN(n6246) );
  OAI211_X1 U7970 ( .C1(n6247), .C2(n6246), .A(n6244), .B(n6245), .ZN(n6248)
         );
  NAND3_X1 U7971 ( .A1(n6248), .A2(n6252), .A3(n6372), .ZN(n6249) );
  NAND3_X1 U7972 ( .A1(n6263), .A2(n7007), .A3(n6249), .ZN(n6257) );
  NAND2_X1 U7973 ( .A1(n6245), .A2(n6250), .ZN(n6253) );
  NAND3_X1 U7974 ( .A1(n6253), .A2(n6252), .A3(n6251), .ZN(n6254) );
  NAND3_X1 U7975 ( .A1(n6254), .A2(n6360), .A3(n6244), .ZN(n6255) );
  NAND2_X1 U7976 ( .A1(n9748), .A2(n9785), .ZN(n6264) );
  NAND2_X1 U7977 ( .A1(n6255), .A2(n6264), .ZN(n6256) );
  AOI21_X1 U7978 ( .B1(n6258), .B2(n6257), .A(n6256), .ZN(n6269) );
  INV_X1 U7979 ( .A(n6259), .ZN(n6262) );
  OAI21_X1 U7980 ( .B1(n8027), .B2(n9817), .A(n6260), .ZN(n6261) );
  OAI21_X1 U7981 ( .B1(n6263), .B2(n6262), .A(n6261), .ZN(n6265) );
  AOI21_X1 U7982 ( .B1(n6265), .B2(n6264), .A(n6372), .ZN(n6268) );
  NAND2_X1 U7983 ( .A1(n6266), .A2(n6360), .ZN(n6267) );
  OAI211_X1 U7984 ( .C1(n6269), .C2(n6268), .A(n7487), .B(n6267), .ZN(n6273)
         );
  MUX2_X1 U7985 ( .A(n6271), .B(n6270), .S(n6372), .Z(n6272) );
  NAND3_X1 U7986 ( .A1(n6273), .A2(n7575), .A3(n6272), .ZN(n6279) );
  NAND2_X1 U7987 ( .A1(n6280), .A2(n6274), .ZN(n6276) );
  INV_X1 U7988 ( .A(n7496), .ZN(n6275) );
  MUX2_X1 U7989 ( .A(n6276), .B(n6275), .S(n6360), .Z(n6277) );
  INV_X1 U7990 ( .A(n6277), .ZN(n6278) );
  NAND3_X1 U7991 ( .A1(n6279), .A2(n6281), .A3(n6278), .ZN(n6286) );
  NAND2_X1 U7992 ( .A1(n6287), .A2(n6280), .ZN(n6283) );
  INV_X1 U7993 ( .A(n6281), .ZN(n6282) );
  MUX2_X1 U7994 ( .A(n6283), .B(n6282), .S(n6372), .Z(n6284) );
  INV_X1 U7995 ( .A(n6284), .ZN(n6285) );
  NAND3_X1 U7996 ( .A1(n6286), .A2(n6288), .A3(n6285), .ZN(n6293) );
  NAND2_X1 U7997 ( .A1(n7785), .A2(n6287), .ZN(n6290) );
  NAND2_X1 U7998 ( .A1(n6298), .A2(n6288), .ZN(n6289) );
  MUX2_X1 U7999 ( .A(n6290), .B(n6289), .S(n6360), .Z(n6291) );
  INV_X1 U8000 ( .A(n6291), .ZN(n6292) );
  NAND2_X1 U8001 ( .A1(n6293), .A2(n6292), .ZN(n6299) );
  NAND2_X1 U8002 ( .A1(n6299), .A2(n6294), .ZN(n6295) );
  NAND3_X1 U8003 ( .A1(n6295), .A2(n7844), .A3(n7846), .ZN(n6297) );
  NAND2_X1 U8004 ( .A1(n6297), .A2(n6296), .ZN(n6304) );
  NAND3_X1 U8005 ( .A1(n6299), .A2(n7846), .A3(n6298), .ZN(n6301) );
  NAND3_X1 U8006 ( .A1(n6301), .A2(n7844), .A3(n6300), .ZN(n6302) );
  NAND2_X1 U8007 ( .A1(n6302), .A2(n8875), .ZN(n6303) );
  MUX2_X1 U8008 ( .A(n6304), .B(n6303), .S(n6372), .Z(n6307) );
  INV_X1 U8009 ( .A(n8863), .ZN(n8878) );
  MUX2_X1 U8010 ( .A(n6305), .B(n7920), .S(n6372), .Z(n6306) );
  OAI211_X1 U8011 ( .C1(n6307), .C2(n8878), .A(n7924), .B(n6306), .ZN(n6311)
         );
  MUX2_X1 U8012 ( .A(n6309), .B(n6308), .S(n6372), .Z(n6310) );
  INV_X1 U8013 ( .A(n6313), .ZN(n6317) );
  OAI211_X1 U8014 ( .C1(n8855), .C2(n6315), .A(n6324), .B(n6314), .ZN(n6316)
         );
  MUX2_X1 U8015 ( .A(n6317), .B(n6316), .S(n6360), .Z(n6318) );
  NAND2_X1 U8016 ( .A1(n6325), .A2(n6323), .ZN(n6319) );
  NAND2_X1 U8017 ( .A1(n6319), .A2(n8803), .ZN(n6320) );
  NAND3_X1 U8018 ( .A1(n6320), .A2(n6331), .A3(n6326), .ZN(n6321) );
  NAND3_X1 U8019 ( .A1(n6321), .A2(n6328), .A3(n6333), .ZN(n6322) );
  INV_X1 U8020 ( .A(n8562), .ZN(n8807) );
  NAND2_X1 U8021 ( .A1(n8787), .A2(n8807), .ZN(n6330) );
  NAND3_X1 U8022 ( .A1(n6322), .A2(n6338), .A3(n6330), .ZN(n6336) );
  NAND2_X1 U8023 ( .A1(n6327), .A2(n6326), .ZN(n6329) );
  NAND2_X1 U8024 ( .A1(n6329), .A2(n6328), .ZN(n6332) );
  NAND3_X1 U8025 ( .A1(n6332), .A2(n6331), .A3(n6330), .ZN(n6334) );
  NAND3_X1 U8026 ( .A1(n6334), .A2(n6337), .A3(n6333), .ZN(n6335) );
  MUX2_X1 U8027 ( .A(n6336), .B(n6335), .S(n6372), .Z(n6340) );
  MUX2_X1 U8028 ( .A(n6338), .B(n6337), .S(n6360), .Z(n6339) );
  NAND3_X1 U8029 ( .A1(n6340), .A2(n8761), .A3(n6339), .ZN(n6341) );
  OAI211_X1 U8030 ( .C1(n6360), .C2(n8743), .A(n6342), .B(n6341), .ZN(n6346)
         );
  MUX2_X1 U8031 ( .A(n6344), .B(n6343), .S(n6360), .Z(n6345) );
  NAND3_X1 U8032 ( .A1(n6346), .A2(n8724), .A3(n6345), .ZN(n6351) );
  INV_X1 U8033 ( .A(n8689), .ZN(n6349) );
  INV_X1 U8034 ( .A(n6347), .ZN(n6348) );
  MUX2_X1 U8035 ( .A(n6349), .B(n6348), .S(n6372), .Z(n6350) );
  MUX2_X1 U8036 ( .A(n6354), .B(n6353), .S(n6372), .Z(n6355) );
  MUX2_X1 U8037 ( .A(n6358), .B(n6357), .S(n6372), .Z(n6359) );
  MUX2_X1 U8038 ( .A(n6362), .B(n6361), .S(n6360), .Z(n6363) );
  NAND3_X1 U8039 ( .A1(n6365), .A2(n6364), .A3(n6363), .ZN(n6369) );
  MUX2_X1 U8040 ( .A(n6367), .B(n6366), .S(n6372), .Z(n6368) );
  OAI21_X1 U8041 ( .B1(n6370), .B2(n6369), .A(n6368), .ZN(n6377) );
  INV_X1 U8042 ( .A(n6371), .ZN(n6373) );
  MUX2_X1 U8043 ( .A(n6374), .B(n6373), .S(n6372), .Z(n6376) );
  AOI21_X1 U8044 ( .B1(n6377), .B2(n6376), .A(n6375), .ZN(n6379) );
  NAND3_X1 U8045 ( .A1(n6379), .A2(n6982), .A3(n9801), .ZN(n6378) );
  OAI21_X1 U8046 ( .B1(n6380), .B2(n6379), .A(n6378), .ZN(n6381) );
  INV_X1 U8047 ( .A(P2_B_REG_SCAN_IN), .ZN(n9994) );
  NOR4_X1 U8048 ( .A1(n6383), .A2(n8880), .A3(n7677), .A4(n9790), .ZN(n6384)
         );
  AOI211_X1 U8049 ( .C1(n6517), .C2(n7407), .A(n9994), .B(n6384), .ZN(n6385)
         );
  INV_X1 U8050 ( .A(n6772), .ZN(n7455) );
  OR2_X1 U8051 ( .A1(n8279), .A2(n7455), .ZN(n6386) );
  OR2_X1 U8052 ( .A1(n6773), .A2(n7455), .ZN(n6701) );
  NAND2_X1 U8053 ( .A1(n6386), .A2(n6701), .ZN(n9181) );
  OR2_X1 U8054 ( .A1(n9181), .A2(n6387), .ZN(n6388) );
  NAND2_X1 U8055 ( .A1(n6388), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U8056 ( .A(n9798), .ZN(n6389) );
  NOR2_X2 U8057 ( .A1(n6558), .A2(n6389), .ZN(P2_U3966) );
  NOR2_X2 U8058 ( .A1(n6701), .A2(P1_U3084), .ZN(P1_U4006) );
  MUX2_X1 U8059 ( .A(n7368), .B(P1_REG2_REG_11__SCAN_IN), .S(n6515), .Z(n6390)
         );
  INV_X1 U8060 ( .A(n6390), .ZN(n6794) );
  NOR2_X1 U8061 ( .A1(n6490), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6391) );
  AOI21_X1 U8062 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6490), .A(n6391), .ZN(
        n9607) );
  NOR2_X1 U8063 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n9148), .ZN(n6392) );
  AOI21_X1 U8064 ( .B1(n9148), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6392), .ZN(
        n9144) );
  MUX2_X1 U8065 ( .A(n5734), .B(P1_REG2_REG_1__SCAN_IN), .S(n6461), .Z(n9137)
         );
  AND2_X1 U8066 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9136) );
  NAND2_X1 U8067 ( .A1(n9137), .A2(n9136), .ZN(n9135) );
  INV_X1 U8068 ( .A(n6461), .ZN(n9131) );
  NAND2_X1 U8069 ( .A1(n9131), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6393) );
  NAND2_X1 U8070 ( .A1(n9135), .A2(n6393), .ZN(n6677) );
  XNOR2_X1 U8071 ( .A(n6463), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n6678) );
  AND2_X1 U8072 ( .A1(n6677), .A2(n6678), .ZN(n6679) );
  INV_X1 U8073 ( .A(n6679), .ZN(n6395) );
  INV_X1 U8074 ( .A(n6463), .ZN(n6684) );
  NAND2_X1 U8075 ( .A1(n6684), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6394) );
  NAND2_X1 U8076 ( .A1(n6395), .A2(n6394), .ZN(n6548) );
  INV_X1 U8077 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10074) );
  MUX2_X1 U8078 ( .A(n10074), .B(P1_REG2_REG_3__SCAN_IN), .S(n6465), .Z(n6549)
         );
  NAND2_X1 U8079 ( .A1(n6548), .A2(n6549), .ZN(n6547) );
  INV_X1 U8080 ( .A(n6465), .ZN(n6552) );
  NAND2_X1 U8081 ( .A1(n6552), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6396) );
  NAND2_X1 U8082 ( .A1(n6547), .A2(n6396), .ZN(n9577) );
  MUX2_X1 U8083 ( .A(n7182), .B(P1_REG2_REG_4__SCAN_IN), .S(n9584), .Z(n9578)
         );
  NOR2_X1 U8084 ( .A1(n9577), .A2(n9578), .ZN(n9576) );
  NOR2_X1 U8085 ( .A1(n9584), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6397) );
  OR2_X1 U8086 ( .A1(n9576), .A2(n6397), .ZN(n6592) );
  XNOR2_X1 U8087 ( .A(n6590), .B(n6398), .ZN(n6593) );
  NAND2_X1 U8088 ( .A1(n6592), .A2(n6593), .ZN(n6591) );
  OR2_X1 U8089 ( .A1(n6590), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6399) );
  NAND2_X1 U8090 ( .A1(n6591), .A2(n6399), .ZN(n9595) );
  OR2_X1 U8091 ( .A1(n6479), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6401) );
  NAND2_X1 U8092 ( .A1(n6479), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6400) );
  NAND2_X1 U8093 ( .A1(n6401), .A2(n6400), .ZN(n9594) );
  NAND2_X1 U8094 ( .A1(n9607), .A2(n9606), .ZN(n9605) );
  OAI21_X1 U8095 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6490), .A(n9605), .ZN(
        n6443) );
  NAND2_X1 U8096 ( .A1(n6448), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6402) );
  OAI21_X1 U8097 ( .B1(n6448), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6402), .ZN(
        n6442) );
  NOR2_X1 U8098 ( .A1(n6443), .A2(n6442), .ZN(n6441) );
  AOI21_X1 U8099 ( .B1(n6448), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6441), .ZN(
        n6601) );
  NAND2_X1 U8100 ( .A1(n6603), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6403) );
  OAI21_X1 U8101 ( .B1(n6603), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6403), .ZN(
        n6600) );
  NAND2_X1 U8102 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6833), .ZN(n6404) );
  OAI21_X1 U8103 ( .B1(n6833), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6404), .ZN(
        n6829) );
  NOR2_X1 U8104 ( .A1(n6830), .A2(n6829), .ZN(n6828) );
  AOI21_X1 U8105 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n6833), .A(n6828), .ZN(
        n6923) );
  NAND2_X1 U8106 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n6925), .ZN(n6405) );
  OAI21_X1 U8107 ( .B1(n6925), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6405), .ZN(
        n6922) );
  NOR2_X1 U8108 ( .A1(n6923), .A2(n6922), .ZN(n6921) );
  INV_X1 U8109 ( .A(n6430), .ZN(n7217) );
  NAND2_X1 U8110 ( .A1(n6406), .A2(n7217), .ZN(n6407) );
  INV_X1 U8111 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7213) );
  XNOR2_X1 U8112 ( .A(n7604), .B(n7611), .ZN(n6410) );
  INV_X1 U8113 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n6409) );
  NOR2_X1 U8114 ( .A1(n6409), .A2(n6410), .ZN(n7605) );
  OR2_X1 U8115 ( .A1(n6068), .A2(P1_U3084), .ZN(n7711) );
  OR2_X1 U8116 ( .A1(n9181), .A2(n7711), .ZN(n6431) );
  INV_X1 U8117 ( .A(n6431), .ZN(n6408) );
  INV_X1 U8118 ( .A(n8412), .ZN(n6498) );
  NAND2_X1 U8119 ( .A1(n6408), .A2(n6498), .ZN(n9598) );
  AOI211_X1 U8120 ( .C1(n6410), .C2(n6409), .A(n7605), .B(n9598), .ZN(n6440)
         );
  INV_X1 U8121 ( .A(P1_U3083), .ZN(n6503) );
  NAND2_X1 U8122 ( .A1(n6503), .A2(n6701), .ZN(n9619) );
  INV_X1 U8123 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n6411) );
  NOR2_X1 U8124 ( .A1(n9619), .A2(n6411), .ZN(n6439) );
  INV_X1 U8125 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7823) );
  MUX2_X1 U8126 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n6412), .S(n6430), .Z(n7211)
         );
  INV_X1 U8127 ( .A(n6925), .ZN(n6788) );
  NOR2_X1 U8128 ( .A1(n6788), .A2(n6413), .ZN(n6414) );
  AOI21_X1 U8129 ( .B1(n6413), .B2(n6788), .A(n6414), .ZN(n6918) );
  INV_X1 U8130 ( .A(n6603), .ZN(n6510) );
  AOI22_X1 U8131 ( .A1(n6603), .A2(P1_REG1_REG_10__SCAN_IN), .B1(n5841), .B2(
        n6510), .ZN(n6605) );
  NAND2_X1 U8132 ( .A1(n6490), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6415) );
  OAI21_X1 U8133 ( .B1(n6490), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6415), .ZN(
        n9610) );
  NOR2_X1 U8134 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n9148), .ZN(n6416) );
  AOI21_X1 U8135 ( .B1(n9148), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6416), .ZN(
        n9151) );
  INV_X1 U8136 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9727) );
  MUX2_X1 U8137 ( .A(n9727), .B(P1_REG1_REG_1__SCAN_IN), .S(n6461), .Z(n9134)
         );
  AND2_X1 U8138 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9133) );
  NAND2_X1 U8139 ( .A1(n9134), .A2(n9133), .ZN(n9132) );
  NAND2_X1 U8140 ( .A1(n9131), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6417) );
  NAND2_X1 U8141 ( .A1(n9132), .A2(n6417), .ZN(n6686) );
  XNOR2_X1 U8142 ( .A(n6463), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n6687) );
  NAND2_X1 U8143 ( .A1(n6686), .A2(n6687), .ZN(n6685) );
  NAND2_X1 U8144 ( .A1(n6684), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6418) );
  NAND2_X1 U8145 ( .A1(n6685), .A2(n6418), .ZN(n6554) );
  MUX2_X1 U8146 ( .A(n5765), .B(P1_REG1_REG_3__SCAN_IN), .S(n6465), .Z(n6555)
         );
  NAND2_X1 U8147 ( .A1(n6554), .A2(n6555), .ZN(n6553) );
  NAND2_X1 U8148 ( .A1(n6552), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6419) );
  NAND2_X1 U8149 ( .A1(n6553), .A2(n6419), .ZN(n9574) );
  INV_X1 U8150 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9732) );
  MUX2_X1 U8151 ( .A(n9732), .B(P1_REG1_REG_4__SCAN_IN), .S(n9584), .Z(n9575)
         );
  NOR2_X1 U8152 ( .A1(n9574), .A2(n9575), .ZN(n9573) );
  NOR2_X1 U8153 ( .A1(n9584), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6420) );
  OR2_X1 U8154 ( .A1(n9573), .A2(n6420), .ZN(n6588) );
  NAND2_X1 U8155 ( .A1(n6590), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6422) );
  OR2_X1 U8156 ( .A1(n6590), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6421) );
  NAND2_X1 U8157 ( .A1(n6422), .A2(n6421), .ZN(n6587) );
  NOR2_X1 U8158 ( .A1(n6588), .A2(n6587), .ZN(n6586) );
  INV_X1 U8159 ( .A(n6422), .ZN(n6423) );
  OR2_X1 U8160 ( .A1(n6586), .A2(n6423), .ZN(n9590) );
  NAND2_X1 U8161 ( .A1(n6479), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6425) );
  OR2_X1 U8162 ( .A1(n6479), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6424) );
  NAND2_X1 U8163 ( .A1(n6425), .A2(n6424), .ZN(n9589) );
  OAI21_X1 U8164 ( .B1(n6479), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6426), .ZN(
        n9150) );
  NAND2_X1 U8165 ( .A1(n9151), .A2(n9150), .ZN(n9149) );
  OAI21_X1 U8166 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n9148), .A(n9149), .ZN(
        n9611) );
  NOR2_X1 U8167 ( .A1(n9610), .A2(n9611), .ZN(n9609) );
  AOI21_X1 U8168 ( .B1(n6490), .B2(P1_REG1_REG_8__SCAN_IN), .A(n9609), .ZN(
        n6445) );
  MUX2_X1 U8169 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n6427), .S(n6448), .Z(n6446)
         );
  NAND2_X1 U8170 ( .A1(n6445), .A2(n6446), .ZN(n6444) );
  OAI21_X1 U8171 ( .B1(n6448), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6444), .ZN(
        n6606) );
  NAND2_X1 U8172 ( .A1(n6605), .A2(n6606), .ZN(n6604) );
  OAI21_X1 U8173 ( .B1(n6603), .B2(P1_REG1_REG_10__SCAN_IN), .A(n6604), .ZN(
        n6791) );
  MUX2_X1 U8174 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n6428), .S(n6515), .Z(n6790)
         );
  NAND2_X1 U8175 ( .A1(n6791), .A2(n6790), .ZN(n6789) );
  OAI21_X1 U8176 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n6515), .A(n6789), .ZN(
        n6825) );
  MUX2_X1 U8177 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6429), .S(n6833), .Z(n6826)
         );
  NAND2_X1 U8178 ( .A1(n6825), .A2(n6826), .ZN(n6824) );
  OAI21_X1 U8179 ( .B1(n6833), .B2(P1_REG1_REG_12__SCAN_IN), .A(n6824), .ZN(
        n6919) );
  NAND2_X1 U8180 ( .A1(n6918), .A2(n6919), .ZN(n6917) );
  OAI21_X1 U8181 ( .B1(n6925), .B2(P1_REG1_REG_13__SCAN_IN), .A(n6917), .ZN(
        n7210) );
  NAND2_X1 U8182 ( .A1(n7211), .A2(n7210), .ZN(n7209) );
  OAI21_X1 U8183 ( .B1(n6430), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7209), .ZN(
        n7610) );
  XNOR2_X1 U8184 ( .A(n7611), .B(n7610), .ZN(n6432) );
  NOR2_X1 U8185 ( .A1(n7823), .A2(n6432), .ZN(n7612) );
  NOR2_X2 U8186 ( .A1(n6431), .A2(n6498), .ZN(n9593) );
  INV_X1 U8187 ( .A(n9593), .ZN(n9608) );
  AOI211_X1 U8188 ( .C1(n7823), .C2(n6432), .A(n7612), .B(n9608), .ZN(n6438)
         );
  INV_X1 U8189 ( .A(n9181), .ZN(n6435) );
  OR2_X1 U8190 ( .A1(n8412), .A2(P1_U3084), .ZN(n9180) );
  INV_X1 U8191 ( .A(n9180), .ZN(n6433) );
  AND2_X1 U8192 ( .A1(n6433), .A2(n6068), .ZN(n6434) );
  AND2_X1 U8193 ( .A1(n6435), .A2(n6434), .ZN(n9585) );
  INV_X1 U8194 ( .A(n9585), .ZN(n9617) );
  NOR2_X1 U8195 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5917), .ZN(n7914) );
  INV_X1 U8196 ( .A(n7914), .ZN(n6436) );
  OAI21_X1 U8197 ( .B1(n9617), .B2(n7611), .A(n6436), .ZN(n6437) );
  OR4_X1 U8198 ( .A1(n6440), .A2(n6439), .A3(n6438), .A4(n6437), .ZN(P1_U3256)
         );
  NOR2_X1 U8199 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5850), .ZN(n7291) );
  AOI211_X1 U8200 ( .C1(n6443), .C2(n6442), .A(n6441), .B(n9598), .ZN(n6451)
         );
  OAI21_X1 U8201 ( .B1(n6446), .B2(n6445), .A(n6444), .ZN(n6447) );
  AND2_X1 U8202 ( .A1(n9593), .A2(n6447), .ZN(n6450) );
  INV_X1 U8203 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10205) );
  INV_X1 U8204 ( .A(n6448), .ZN(n6496) );
  OAI22_X1 U8205 ( .A1(n9619), .A2(n10205), .B1(n9617), .B2(n6496), .ZN(n6449)
         );
  OR4_X1 U8206 ( .A1(n7291), .A2(n6451), .A3(n6450), .A4(n6449), .ZN(P1_U3250)
         );
  NOR2_X1 U8207 ( .A1(n4705), .A2(n9747), .ZN(n6457) );
  OAI22_X1 U8208 ( .A1(n8707), .A2(n9750), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6454), .ZN(n6456) );
  OAI22_X1 U8209 ( .A1(n8747), .A2(n9751), .B1(n8713), .B2(n9759), .ZN(n6455)
         );
  XNOR2_X1 U8210 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AND2_X1 U8211 ( .A1(P1_STATE_REG_SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6499) );
  INV_X1 U8212 ( .A(n6499), .ZN(n6458) );
  OAI21_X1 U8213 ( .B1(n6459), .B2(P1_STATE_REG_SCAN_IN), .A(n6458), .ZN(
        P1_U3353) );
  AND2_X1 U8214 ( .A1(n6051), .A2(P1_U3084), .ZN(n7710) );
  INV_X2 U8215 ( .A(n7710), .ZN(n8419) );
  AND2_X1 U8216 ( .A1(n4980), .A2(P1_U3084), .ZN(n8008) );
  AOI22_X1 U8217 ( .A1(n9584), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n8008), .ZN(n6460) );
  OAI21_X1 U8218 ( .B1(n6469), .B2(n8419), .A(n6460), .ZN(P1_U3349) );
  OAI222_X1 U8219 ( .A1(n8421), .A2(n6462), .B1(n8419), .B2(n6467), .C1(
        P1_U3084), .C2(n6461), .ZN(P1_U3352) );
  OAI222_X1 U8220 ( .A1(n8421), .A2(n6464), .B1(n8419), .B2(n6474), .C1(
        P1_U3084), .C2(n6463), .ZN(P1_U3351) );
  OAI222_X1 U8221 ( .A1(n8421), .A2(n6466), .B1(n8419), .B2(n6471), .C1(
        P1_U3084), .C2(n6465), .ZN(P1_U3350) );
  NOR2_X1 U8222 ( .A1(n4980), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8014) );
  INV_X2 U8223 ( .A(n8014), .ZN(n8459) );
  AND2_X1 U8224 ( .A1(n4980), .A2(P2_U3152), .ZN(n7450) );
  OAI222_X1 U8225 ( .A1(n8459), .A2(n6468), .B1(n4390), .B2(n6467), .C1(
        P2_U3152), .C2(n6579), .ZN(P2_U3357) );
  OAI222_X1 U8226 ( .A1(n8459), .A2(n6470), .B1(n4390), .B2(n6469), .C1(
        P2_U3152), .C2(n6676), .ZN(P2_U3354) );
  OAI222_X1 U8227 ( .A1(n8459), .A2(n6472), .B1(n4390), .B2(n6471), .C1(
        P2_U3152), .C2(n6643), .ZN(P2_U3355) );
  OAI222_X1 U8228 ( .A1(n8459), .A2(n10132), .B1(n4390), .B2(n6474), .C1(
        P2_U3152), .C2(n6473), .ZN(P2_U3356) );
  INV_X1 U8229 ( .A(n6590), .ZN(n6475) );
  OAI222_X1 U8230 ( .A1(n8421), .A2(n9973), .B1(n8419), .B2(n6476), .C1(
        P1_U3084), .C2(n6475), .ZN(P1_U3348) );
  OAI222_X1 U8231 ( .A1(n8459), .A2(n6477), .B1(n4390), .B2(n6476), .C1(
        P2_U3152), .C2(n6585), .ZN(P2_U3353) );
  OAI222_X1 U8232 ( .A1(n8459), .A2(n6478), .B1(n4390), .B2(n6480), .C1(
        P2_U3152), .C2(n6654), .ZN(P2_U3352) );
  INV_X1 U8233 ( .A(n6479), .ZN(n9601) );
  OAI222_X1 U8234 ( .A1(n8421), .A2(n6481), .B1(n8419), .B2(n6480), .C1(
        P1_U3084), .C2(n9601), .ZN(P1_U3347) );
  NAND2_X1 U8235 ( .A1(n6722), .A2(n6536), .ZN(n9668) );
  INV_X1 U8236 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6484) );
  INV_X1 U8237 ( .A(n6482), .ZN(n6483) );
  AOI22_X1 U8238 ( .A1(n9668), .A2(n6484), .B1(n6722), .B2(n6483), .ZN(
        P1_U3441) );
  INV_X1 U8239 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6532) );
  INV_X1 U8240 ( .A(n6534), .ZN(n6485) );
  AOI22_X1 U8241 ( .A1(n9668), .A2(n6532), .B1(n6722), .B2(n6485), .ZN(
        P1_U3440) );
  AOI22_X1 U8242 ( .A1(n9148), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n8008), .ZN(n6486) );
  OAI21_X1 U8243 ( .B1(n6487), .B2(n8419), .A(n6486), .ZN(P1_U3346) );
  OAI222_X1 U8244 ( .A1(n8459), .A2(n6488), .B1(n4390), .B2(n6487), .C1(
        P2_U3152), .C2(n6666), .ZN(P2_U3351) );
  INV_X1 U8245 ( .A(n6489), .ZN(n6492) );
  INV_X1 U8246 ( .A(n6490), .ZN(n9616) );
  OAI222_X1 U8247 ( .A1(n8421), .A2(n6491), .B1(n8419), .B2(n6492), .C1(
        P1_U3084), .C2(n9616), .ZN(P1_U3345) );
  OAI222_X1 U8248 ( .A1(n8459), .A2(n6493), .B1(n4390), .B2(n6492), .C1(
        P2_U3152), .C2(n6817), .ZN(P2_U3350) );
  INV_X1 U8249 ( .A(n6494), .ZN(n6497) );
  OAI222_X1 U8250 ( .A1(n8419), .A2(n6497), .B1(n6496), .B2(P1_U3084), .C1(
        n6495), .C2(n8421), .ZN(P1_U3344) );
  INV_X1 U8251 ( .A(n6883), .ZN(n6823) );
  OAI222_X1 U8252 ( .A1(n8459), .A2(n10175), .B1(n4390), .B2(n6497), .C1(n6823), .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U8253 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6507) );
  AOI21_X1 U8254 ( .B1(n6498), .B2(n5748), .A(n7711), .ZN(n6500) );
  NOR2_X1 U8255 ( .A1(n6500), .A2(n6499), .ZN(n6702) );
  AOI21_X1 U8256 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(P1_REG2_REG_0__SCAN_IN), .A(
        n8412), .ZN(n6501) );
  AOI211_X1 U8257 ( .C1(n6693), .C2(P1_REG1_REG_0__SCAN_IN), .A(n6068), .B(
        n6501), .ZN(n6502) );
  NOR3_X1 U8258 ( .A1(n6503), .A2(n6702), .A3(n6502), .ZN(n6504) );
  AOI21_X1 U8259 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .A(n6504), .ZN(
        n6506) );
  INV_X1 U8260 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6541) );
  NAND3_X1 U8261 ( .A1(n9593), .A2(P1_IR_REG_0__SCAN_IN), .A3(n6541), .ZN(
        n6505) );
  OAI211_X1 U8262 ( .C1(n6507), .C2(n9619), .A(n6506), .B(n6505), .ZN(P1_U3241) );
  INV_X1 U8263 ( .A(n6508), .ZN(n6511) );
  OAI222_X1 U8264 ( .A1(n8419), .A2(n6511), .B1(n6510), .B2(P1_U3084), .C1(
        n6509), .C2(n8421), .ZN(P1_U3343) );
  INV_X1 U8265 ( .A(n6964), .ZN(n6891) );
  OAI222_X1 U8266 ( .A1(n8459), .A2(n6512), .B1(n4390), .B2(n6511), .C1(n6891), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U8267 ( .A(n7078), .ZN(n7087) );
  INV_X1 U8268 ( .A(n6513), .ZN(n6516) );
  OAI222_X1 U8269 ( .A1(P2_U3152), .A2(n7087), .B1(n4390), .B2(n6516), .C1(
        n6514), .C2(n8459), .ZN(P2_U3347) );
  INV_X1 U8270 ( .A(n6515), .ZN(n6796) );
  OAI222_X1 U8271 ( .A1(n8421), .A2(n10129), .B1(n6796), .B2(P1_U3084), .C1(
        n8419), .C2(n6516), .ZN(P1_U3342) );
  INV_X1 U8272 ( .A(n6517), .ZN(n7451) );
  NAND2_X1 U8273 ( .A1(n9790), .A2(n7451), .ZN(n6519) );
  NAND2_X1 U8274 ( .A1(n6519), .A2(n6518), .ZN(n6522) );
  INV_X1 U8275 ( .A(n6561), .ZN(n6520) );
  OR2_X1 U8276 ( .A1(n9790), .A2(n6520), .ZN(n6521) );
  NOR2_X1 U8277 ( .A1(n9766), .A2(P2_U3966), .ZN(P2_U3151) );
  CLKBUF_X1 U8278 ( .A(P1_U4006), .Z(n9904) );
  NAND2_X1 U8279 ( .A1(n5790), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6526) );
  NAND2_X1 U8280 ( .A1(n5789), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6525) );
  INV_X1 U8281 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9187) );
  OR2_X1 U8282 ( .A1(n6058), .A2(n9187), .ZN(n6524) );
  AND3_X1 U8283 ( .A1(n6526), .A2(n6525), .A3(n6524), .ZN(n8231) );
  INV_X1 U8284 ( .A(n8231), .ZN(n9188) );
  NAND2_X1 U8285 ( .A1(n9188), .A2(n9904), .ZN(n6527) );
  OAI21_X1 U8286 ( .B1(n9904), .B2(n6204), .A(n6527), .ZN(P1_U3586) );
  INV_X1 U8287 ( .A(n6528), .ZN(n6531) );
  AOI22_X1 U8288 ( .A1(n6833), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n8008), .ZN(n6529) );
  OAI21_X1 U8289 ( .B1(n6531), .B2(n8419), .A(n6529), .ZN(P1_U3341) );
  AOI22_X1 U8290 ( .A1(n7240), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n8014), .ZN(n6530) );
  OAI21_X1 U8291 ( .B1(n6531), .B2(n4390), .A(n6530), .ZN(P2_U3346) );
  OAI211_X1 U8292 ( .C1(n9350), .C2(n9705), .A(n6726), .B(n6719), .ZN(n6543)
         );
  NOR2_X1 U8293 ( .A1(n6533), .A2(n6532), .ZN(n6535) );
  OAI21_X1 U8294 ( .B1(n6536), .B2(n6535), .A(n6534), .ZN(n6718) );
  INV_X2 U8295 ( .A(n9739), .ZN(n9742) );
  INV_X1 U8296 ( .A(n7144), .ZN(n6537) );
  NAND2_X1 U8297 ( .A1(n6695), .A2(n7148), .ZN(n8368) );
  NAND2_X1 U8298 ( .A1(n6537), .A2(n8368), .ZN(n8251) );
  NAND3_X1 U8299 ( .A1(n8251), .A2(n8414), .A3(n6717), .ZN(n6538) );
  OAI21_X1 U8300 ( .B1(n7194), .B2(n9662), .A(n6538), .ZN(n6952) );
  INV_X1 U8301 ( .A(n6952), .ZN(n6539) );
  OAI21_X1 U8302 ( .B1(n7148), .B2(n6717), .A(n6539), .ZN(n6544) );
  NAND2_X1 U8303 ( .A1(n6544), .A2(n9742), .ZN(n6540) );
  OAI21_X1 U8304 ( .B1(n9742), .B2(n6541), .A(n6540), .ZN(P1_U3523) );
  INV_X2 U8305 ( .A(n9724), .ZN(n9726) );
  INV_X1 U8306 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U8307 ( .A1(n6544), .A2(n9726), .ZN(n6545) );
  OAI21_X1 U8308 ( .B1(n9726), .B2(n6546), .A(n6545), .ZN(P1_U3454) );
  INV_X1 U8309 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10051) );
  AND2_X1 U8310 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6783) );
  INV_X1 U8311 ( .A(n9598), .ZN(n9615) );
  OAI211_X1 U8312 ( .C1(n6549), .C2(n6548), .A(n9615), .B(n6547), .ZN(n6550)
         );
  INV_X1 U8313 ( .A(n6550), .ZN(n6551) );
  AOI211_X1 U8314 ( .C1(n9585), .C2(n6552), .A(n6783), .B(n6551), .ZN(n6557)
         );
  OAI211_X1 U8315 ( .C1(n6555), .C2(n6554), .A(n9593), .B(n6553), .ZN(n6556)
         );
  OAI211_X1 U8316 ( .C1(n10051), .C2(n9619), .A(n6557), .B(n6556), .ZN(
        P1_U3244) );
  INV_X1 U8317 ( .A(n6558), .ZN(n6559) );
  NAND2_X1 U8318 ( .A1(n6559), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6560) );
  OAI211_X1 U8319 ( .C1(n9790), .C2(n6561), .A(n7451), .B(n6560), .ZN(n6563)
         );
  NAND2_X1 U8320 ( .A1(n6563), .A2(n6562), .ZN(n6571) );
  NAND2_X1 U8321 ( .A1(n6571), .A2(n8586), .ZN(n6577) );
  NAND2_X1 U8322 ( .A1(n6577), .A2(n5684), .ZN(n9760) );
  NOR2_X1 U8323 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10169), .ZN(n6575) );
  INV_X1 U8324 ( .A(n6676), .ZN(n6569) );
  MUX2_X1 U8325 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6564), .S(n6676), .Z(n6668)
         );
  INV_X1 U8326 ( .A(n6643), .ZN(n6568) );
  INV_X1 U8327 ( .A(n6579), .ZN(n9460) );
  NAND2_X1 U8328 ( .A1(n9765), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9458) );
  INV_X1 U8329 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6565) );
  NOR2_X1 U8330 ( .A1(n9458), .A2(n9457), .ZN(n9456) );
  AOI21_X1 U8331 ( .B1(n9460), .B2(P2_REG1_REG_1__SCAN_IN), .A(n9456), .ZN(
        n9469) );
  NAND2_X1 U8332 ( .A1(n9471), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6566) );
  OAI21_X1 U8333 ( .B1(n9471), .B2(P2_REG1_REG_2__SCAN_IN), .A(n6566), .ZN(
        n9468) );
  INV_X1 U8334 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6567) );
  MUX2_X1 U8335 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6567), .S(n6643), .Z(n6634)
         );
  NOR2_X1 U8336 ( .A1(n6668), .A2(n4422), .ZN(n6667) );
  NAND2_X1 U8337 ( .A1(n6621), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6570) );
  OAI21_X1 U8338 ( .B1(n6621), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6570), .ZN(
        n6572) );
  INV_X1 U8339 ( .A(n7677), .ZN(n8017) );
  AOI211_X1 U8340 ( .C1(n6573), .C2(n6572), .A(n6611), .B(n9761), .ZN(n6574)
         );
  AOI211_X1 U8341 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n9766), .A(n6575), .B(
        n6574), .ZN(n6584) );
  NOR2_X1 U8342 ( .A1(n5684), .A2(n7677), .ZN(n6576) );
  INV_X1 U8343 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7110) );
  MUX2_X1 U8344 ( .A(n7110), .B(P2_REG2_REG_4__SCAN_IN), .S(n6676), .Z(n6581)
         );
  MUX2_X1 U8345 ( .A(n6999), .B(P2_REG2_REG_3__SCAN_IN), .S(n6643), .Z(n6639)
         );
  NAND2_X1 U8346 ( .A1(n9471), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6580) );
  MUX2_X1 U8347 ( .A(n7097), .B(P2_REG2_REG_2__SCAN_IN), .S(n9471), .Z(n6578)
         );
  INV_X1 U8348 ( .A(n6578), .ZN(n9474) );
  MUX2_X1 U8349 ( .A(n6987), .B(P2_REG2_REG_1__SCAN_IN), .S(n6579), .Z(n9462)
         );
  NAND3_X1 U8350 ( .A1(n9765), .A2(P2_REG2_REG_0__SCAN_IN), .A3(n9462), .ZN(
        n9461) );
  OAI21_X1 U8351 ( .B1(n6579), .B2(n6987), .A(n9461), .ZN(n9475) );
  NAND2_X1 U8352 ( .A1(n9474), .A2(n9475), .ZN(n9473) );
  NAND2_X1 U8353 ( .A1(n6580), .A2(n9473), .ZN(n6640) );
  NAND2_X1 U8354 ( .A1(n6639), .A2(n6640), .ZN(n6638) );
  OAI21_X1 U8355 ( .B1(n6643), .B2(n6999), .A(n6638), .ZN(n6672) );
  NAND2_X1 U8356 ( .A1(n6581), .A2(n6672), .ZN(n6671) );
  OAI21_X1 U8357 ( .B1(n7110), .B2(n6676), .A(n6671), .ZN(n6623) );
  MUX2_X1 U8358 ( .A(n7229), .B(P2_REG2_REG_5__SCAN_IN), .S(n6621), .Z(n6622)
         );
  XNOR2_X1 U8359 ( .A(n6623), .B(n6622), .ZN(n6582) );
  NAND2_X1 U8360 ( .A1(n9764), .A2(n6582), .ZN(n6583) );
  OAI211_X1 U8361 ( .C1(n9760), .C2(n6585), .A(n6584), .B(n6583), .ZN(P2_U3250) );
  INV_X1 U8362 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6597) );
  AND2_X1 U8363 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6862) );
  AOI211_X1 U8364 ( .C1(n6588), .C2(n6587), .A(n6586), .B(n9608), .ZN(n6589)
         );
  AOI211_X1 U8365 ( .C1(n9585), .C2(n6590), .A(n6862), .B(n6589), .ZN(n6596)
         );
  OAI21_X1 U8366 ( .B1(n6593), .B2(n6592), .A(n6591), .ZN(n6594) );
  NAND2_X1 U8367 ( .A1(n9615), .A2(n6594), .ZN(n6595) );
  OAI211_X1 U8368 ( .C1(n6597), .C2(n9619), .A(n6596), .B(n6595), .ZN(P1_U3246) );
  INV_X1 U8369 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6610) );
  NOR2_X1 U8370 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6598), .ZN(n7355) );
  AOI211_X1 U8371 ( .C1(n6601), .C2(n6600), .A(n6599), .B(n9598), .ZN(n6602)
         );
  AOI211_X1 U8372 ( .C1(n9585), .C2(n6603), .A(n7355), .B(n6602), .ZN(n6609)
         );
  OAI21_X1 U8373 ( .B1(n6606), .B2(n6605), .A(n6604), .ZN(n6607) );
  NAND2_X1 U8374 ( .A1(n6607), .A2(n9593), .ZN(n6608) );
  OAI211_X1 U8375 ( .C1(n9619), .C2(n6610), .A(n6609), .B(n6608), .ZN(P1_U3251) );
  AND2_X1 U8376 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n7381) );
  NAND2_X1 U8377 ( .A1(n6619), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6612) );
  OAI21_X1 U8378 ( .B1(n6619), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6612), .ZN(
        n6645) );
  AOI21_X1 U8379 ( .B1(n6619), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6644), .ZN(
        n6658) );
  NAND2_X1 U8380 ( .A1(n6617), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6613) );
  OAI21_X1 U8381 ( .B1(n6617), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6613), .ZN(
        n6657) );
  NOR2_X1 U8382 ( .A1(n6658), .A2(n6657), .ZN(n6656) );
  AOI21_X1 U8383 ( .B1(n6617), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6656), .ZN(
        n6615) );
  XOR2_X1 U8384 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6817), .Z(n6614) );
  AOI211_X1 U8385 ( .C1(n6615), .C2(n6614), .A(n6809), .B(n9761), .ZN(n6616)
         );
  AOI211_X1 U8386 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n9766), .A(n7381), .B(
        n6616), .ZN(n6632) );
  NAND2_X1 U8387 ( .A1(n6617), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6628) );
  MUX2_X1 U8388 ( .A(n5310), .B(P2_REG2_REG_7__SCAN_IN), .S(n6617), .Z(n6618)
         );
  INV_X1 U8389 ( .A(n6618), .ZN(n6662) );
  NAND2_X1 U8390 ( .A1(n6619), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6627) );
  MUX2_X1 U8391 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6620), .S(n6619), .Z(n6650)
         );
  NAND2_X1 U8392 ( .A1(n6621), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6626) );
  INV_X1 U8393 ( .A(n6622), .ZN(n6624) );
  NAND2_X1 U8394 ( .A1(n6624), .A2(n6623), .ZN(n6625) );
  NAND2_X1 U8395 ( .A1(n6626), .A2(n6625), .ZN(n6651) );
  NAND2_X1 U8396 ( .A1(n6650), .A2(n6651), .ZN(n6649) );
  NAND2_X1 U8397 ( .A1(n6627), .A2(n6649), .ZN(n6663) );
  NAND2_X1 U8398 ( .A1(n6662), .A2(n6663), .ZN(n6661) );
  NAND2_X1 U8399 ( .A1(n6628), .A2(n6661), .ZN(n6630) );
  MUX2_X1 U8400 ( .A(n7522), .B(P2_REG2_REG_8__SCAN_IN), .S(n6817), .Z(n6629)
         );
  NAND2_X1 U8401 ( .A1(n6630), .A2(n6629), .ZN(n6816) );
  OAI211_X1 U8402 ( .C1(n6630), .C2(n6629), .A(n9764), .B(n6816), .ZN(n6631)
         );
  OAI211_X1 U8403 ( .C1(n9760), .C2(n6817), .A(n6632), .B(n6631), .ZN(P2_U3253) );
  NOR2_X1 U8404 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5252), .ZN(n6637) );
  AOI211_X1 U8405 ( .C1(n6635), .C2(n6634), .A(n6633), .B(n9761), .ZN(n6636)
         );
  AOI211_X1 U8406 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n9766), .A(n6637), .B(
        n6636), .ZN(n6642) );
  OAI211_X1 U8407 ( .C1(n6640), .C2(n6639), .A(n9764), .B(n6638), .ZN(n6641)
         );
  OAI211_X1 U8408 ( .C1(n9760), .C2(n6643), .A(n6642), .B(n6641), .ZN(P2_U3248) );
  NAND2_X1 U8409 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8128) );
  INV_X1 U8410 ( .A(n8128), .ZN(n6648) );
  AOI211_X1 U8411 ( .C1(n6646), .C2(n6645), .A(n6644), .B(n9761), .ZN(n6647)
         );
  AOI211_X1 U8412 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n9766), .A(n6648), .B(
        n6647), .ZN(n6653) );
  OAI211_X1 U8413 ( .C1(n6651), .C2(n6650), .A(n9764), .B(n6649), .ZN(n6652)
         );
  OAI211_X1 U8414 ( .C1(n9760), .C2(n6654), .A(n6653), .B(n6652), .ZN(P2_U3251) );
  NOR2_X1 U8415 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6655), .ZN(n6660) );
  AOI211_X1 U8416 ( .C1(n6658), .C2(n6657), .A(n6656), .B(n9761), .ZN(n6659)
         );
  AOI211_X1 U8417 ( .C1(P2_ADDR_REG_7__SCAN_IN), .C2(n9766), .A(n6660), .B(
        n6659), .ZN(n6665) );
  OAI211_X1 U8418 ( .C1(n6663), .C2(n6662), .A(n9764), .B(n6661), .ZN(n6664)
         );
  OAI211_X1 U8419 ( .C1(n9760), .C2(n6666), .A(n6665), .B(n6664), .ZN(P2_U3252) );
  AND2_X1 U8420 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n8549) );
  AOI211_X1 U8421 ( .C1(n4422), .C2(n6668), .A(n6667), .B(n9761), .ZN(n6669)
         );
  AOI211_X1 U8422 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n9766), .A(n8549), .B(
        n6669), .ZN(n6675) );
  MUX2_X1 U8423 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7110), .S(n6676), .Z(n6670)
         );
  INV_X1 U8424 ( .A(n6670), .ZN(n6673) );
  OAI211_X1 U8425 ( .C1(n6673), .C2(n6672), .A(n9764), .B(n6671), .ZN(n6674)
         );
  OAI211_X1 U8426 ( .C1(n9760), .C2(n6676), .A(n6675), .B(n6674), .ZN(P2_U3249) );
  INV_X1 U8427 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6690) );
  NOR2_X1 U8428 ( .A1(n7198), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6683) );
  INV_X1 U8429 ( .A(n6677), .ZN(n6681) );
  INV_X1 U8430 ( .A(n6678), .ZN(n6680) );
  AOI211_X1 U8431 ( .C1(n6681), .C2(n6680), .A(n6679), .B(n9598), .ZN(n6682)
         );
  AOI211_X1 U8432 ( .C1(n9585), .C2(n6684), .A(n6683), .B(n6682), .ZN(n6689)
         );
  OAI211_X1 U8433 ( .C1(n6687), .C2(n6686), .A(n9593), .B(n6685), .ZN(n6688)
         );
  OAI211_X1 U8434 ( .C1(n6690), .C2(n9619), .A(n6689), .B(n6688), .ZN(n6704)
         );
  OAI22_X1 U8435 ( .A1(n6851), .A2(n7148), .B1(n6773), .B2(n6693), .ZN(n6694)
         );
  INV_X2 U8436 ( .A(n6851), .ZN(n6846) );
  NAND2_X1 U8437 ( .A1(n6695), .A2(n6846), .ZN(n6700) );
  INV_X1 U8438 ( .A(n6707), .ZN(n6735) );
  NAND2_X1 U8439 ( .A1(n6696), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6697) );
  INV_X1 U8440 ( .A(n6698), .ZN(n6699) );
  XOR2_X1 U8441 ( .A(n6706), .B(n6705), .Z(n6754) );
  MUX2_X1 U8442 ( .A(n9136), .B(n6754), .S(n8412), .Z(n6703) );
  AOI211_X1 U8443 ( .C1(n6703), .C2(n6729), .A(n6702), .B(n6701), .ZN(n9582)
         );
  OR2_X1 U8444 ( .A1(n6704), .A2(n9582), .ZN(P1_U3243) );
  OAI22_X1 U8445 ( .A1(n6850), .A2(n7194), .B1(n9671), .B2(n6851), .ZN(n6740)
         );
  NAND2_X1 U8446 ( .A1(n6846), .A2(n9130), .ZN(n6709) );
  NAND2_X1 U8447 ( .A1(n6707), .A2(n7142), .ZN(n6708) );
  NAND2_X1 U8448 ( .A1(n6709), .A2(n6708), .ZN(n6710) );
  XNOR2_X1 U8449 ( .A(n6710), .B(n8062), .ZN(n6712) );
  NAND2_X1 U8450 ( .A1(n6711), .A2(n6712), .ZN(n6741) );
  INV_X1 U8451 ( .A(n6711), .ZN(n6714) );
  INV_X1 U8452 ( .A(n6712), .ZN(n6713) );
  NAND2_X1 U8453 ( .A1(n6714), .A2(n6713), .ZN(n6742) );
  NAND2_X1 U8454 ( .A1(n6741), .A2(n6742), .ZN(n6715) );
  XOR2_X1 U8455 ( .A(n6740), .B(n6715), .Z(n6734) );
  NAND2_X1 U8456 ( .A1(n9718), .A2(n8279), .ZN(n6777) );
  INV_X1 U8457 ( .A(n6777), .ZN(n6720) );
  OR2_X1 U8458 ( .A1(n6719), .A2(n6718), .ZN(n6723) );
  INV_X1 U8459 ( .A(n6722), .ZN(n8413) );
  NOR2_X1 U8460 ( .A1(n6723), .A2(n8413), .ZN(n6727) );
  NAND2_X1 U8461 ( .A1(n6720), .A2(n6727), .ZN(n9095) );
  INV_X1 U8462 ( .A(n6723), .ZN(n6776) );
  NAND2_X1 U8463 ( .A1(n6721), .A2(n8414), .ZN(n6725) );
  AND2_X1 U8464 ( .A1(n6723), .A2(n6722), .ZN(n6724) );
  NAND2_X1 U8465 ( .A1(n6725), .A2(n6724), .ZN(n6779) );
  AND2_X1 U8466 ( .A1(n6779), .A2(n6726), .ZN(n6947) );
  AOI21_X1 U8467 ( .B1(n6726), .B2(n6776), .A(n9100), .ZN(n6752) );
  INV_X1 U8468 ( .A(n9100), .ZN(n9115) );
  INV_X1 U8469 ( .A(n8414), .ZN(n6728) );
  NAND2_X1 U8470 ( .A1(n6728), .A2(n6727), .ZN(n6730) );
  INV_X1 U8471 ( .A(n9110), .ZN(n7915) );
  INV_X1 U8472 ( .A(n9106), .ZN(n9088) );
  AOI22_X1 U8473 ( .A1(n7915), .A2(n6695), .B1(n9088), .B2(n9129), .ZN(n6731)
         );
  OAI21_X1 U8474 ( .B1(n9115), .B2(n9671), .A(n6731), .ZN(n6732) );
  AOI21_X1 U8475 ( .B1(n6752), .B2(P1_REG3_REG_1__SCAN_IN), .A(n6732), .ZN(
        n6733) );
  OAI21_X1 U8476 ( .B1(n6734), .B2(n9095), .A(n6733), .ZN(P1_U3220) );
  NAND2_X1 U8477 ( .A1(n6846), .A2(n9129), .ZN(n6737) );
  NAND2_X1 U8478 ( .A1(n6707), .A2(n7205), .ZN(n6736) );
  XNOR2_X1 U8479 ( .A(n6739), .B(n6738), .ZN(n6755) );
  OAI22_X1 U8480 ( .A1(n6850), .A2(n7160), .B1(n9676), .B2(n6851), .ZN(n6756)
         );
  NAND2_X1 U8481 ( .A1(n6741), .A2(n6740), .ZN(n6743) );
  INV_X1 U8482 ( .A(n6760), .ZN(n6745) );
  AOI21_X1 U8483 ( .B1(n6744), .B2(n6746), .A(n6745), .ZN(n6750) );
  AOI22_X1 U8484 ( .A1(n9088), .A2(n9128), .B1(n7915), .B2(n9130), .ZN(n6747)
         );
  OAI21_X1 U8485 ( .B1(n9115), .B2(n9676), .A(n6747), .ZN(n6748) );
  AOI21_X1 U8486 ( .B1(n6752), .B2(P1_REG3_REG_2__SCAN_IN), .A(n6748), .ZN(
        n6749) );
  OAI21_X1 U8487 ( .B1(n6750), .B2(n9095), .A(n6749), .ZN(P1_U3235) );
  OAI22_X1 U8488 ( .A1(n9115), .A2(n7148), .B1(n7194), .B2(n9106), .ZN(n6751)
         );
  AOI21_X1 U8489 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n6752), .A(n6751), .ZN(
        n6753) );
  OAI21_X1 U8490 ( .B1(n9095), .B2(n6754), .A(n6753), .ZN(P1_U3230) );
  INV_X1 U8491 ( .A(n6755), .ZN(n6758) );
  INV_X1 U8492 ( .A(n6756), .ZN(n6757) );
  NAND2_X1 U8493 ( .A1(n6758), .A2(n6757), .ZN(n6759) );
  NAND2_X1 U8494 ( .A1(n8113), .A2(n9128), .ZN(n6762) );
  NAND2_X1 U8495 ( .A1(n6707), .A2(n7166), .ZN(n6761) );
  NAND2_X1 U8496 ( .A1(n6762), .A2(n6761), .ZN(n6763) );
  XNOR2_X1 U8497 ( .A(n6763), .B(n8062), .ZN(n6766) );
  NOR2_X1 U8498 ( .A1(n6851), .A2(n9683), .ZN(n6765) );
  AOI21_X1 U8499 ( .B1(n6764), .B2(n9128), .A(n6765), .ZN(n6767) );
  AND2_X1 U8500 ( .A1(n6766), .A2(n6767), .ZN(n6844) );
  INV_X1 U8501 ( .A(n6844), .ZN(n6770) );
  INV_X1 U8502 ( .A(n6766), .ZN(n6769) );
  INV_X1 U8503 ( .A(n6767), .ZN(n6768) );
  NAND2_X1 U8504 ( .A1(n6769), .A2(n6768), .ZN(n6843) );
  NAND2_X1 U8505 ( .A1(n6770), .A2(n6843), .ZN(n6771) );
  XNOR2_X1 U8506 ( .A(n6845), .B(n6771), .ZN(n6786) );
  AND3_X1 U8507 ( .A1(n6774), .A2(n6773), .A3(n6772), .ZN(n6775) );
  OAI21_X1 U8508 ( .B1(n6777), .B2(n6776), .A(n6775), .ZN(n6778) );
  NAND2_X1 U8509 ( .A1(n6778), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6780) );
  INV_X1 U8510 ( .A(n9108), .ZN(n9089) );
  INV_X1 U8511 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6781) );
  AOI22_X1 U8512 ( .A1(n9089), .A2(n6781), .B1(n7915), .B2(n9129), .ZN(n6785)
         );
  NOR2_X1 U8513 ( .A1(n9106), .A2(n9659), .ZN(n6782) );
  AOI211_X1 U8514 ( .C1(n9100), .C2(n7166), .A(n6783), .B(n6782), .ZN(n6784)
         );
  OAI211_X1 U8515 ( .C1(n6786), .C2(n9095), .A(n6785), .B(n6784), .ZN(P1_U3216) );
  INV_X1 U8516 ( .A(n6787), .ZN(n6802) );
  OAI222_X1 U8517 ( .A1(n8419), .A2(n6802), .B1(n6788), .B2(P1_U3084), .C1(
        n10178), .C2(n8421), .ZN(P1_U3340) );
  INV_X1 U8518 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6801) );
  OAI21_X1 U8519 ( .B1(n6791), .B2(n6790), .A(n6789), .ZN(n6792) );
  NAND2_X1 U8520 ( .A1(n6792), .A2(n9593), .ZN(n6800) );
  OAI21_X1 U8521 ( .B1(n6795), .B2(n6794), .A(n6793), .ZN(n6798) );
  AND2_X1 U8522 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3084), .ZN(n7437) );
  NOR2_X1 U8523 ( .A1(n9617), .A2(n6796), .ZN(n6797) );
  AOI211_X1 U8524 ( .C1(n9615), .C2(n6798), .A(n7437), .B(n6797), .ZN(n6799)
         );
  OAI211_X1 U8525 ( .C1(n9619), .C2(n6801), .A(n6800), .B(n6799), .ZN(P1_U3252) );
  INV_X1 U8526 ( .A(n7389), .ZN(n7245) );
  OAI222_X1 U8527 ( .A1(n8459), .A2(n6803), .B1(n4390), .B2(n6802), .C1(n7245), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8528 ( .A(n6804), .ZN(n6805) );
  OAI222_X1 U8529 ( .A1(n8419), .A2(n6805), .B1(n7217), .B2(P1_U3084), .C1(
        n10160), .C2(n8421), .ZN(P1_U3339) );
  INV_X1 U8530 ( .A(n7743), .ZN(n7740) );
  OAI222_X1 U8531 ( .A1(n8459), .A2(n6806), .B1(n4390), .B2(n6805), .C1(n7740), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8532 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6808) );
  NAND2_X1 U8533 ( .A1(n8019), .A2(P2_U3966), .ZN(n6807) );
  OAI21_X1 U8534 ( .B1(P2_U3966), .B2(n6808), .A(n6807), .ZN(P2_U3583) );
  NOR2_X1 U8535 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7550), .ZN(n6815) );
  INV_X1 U8536 ( .A(n6817), .ZN(n6810) );
  INV_X1 U8537 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6811) );
  MUX2_X1 U8538 ( .A(n6811), .B(P2_REG1_REG_9__SCAN_IN), .S(n6883), .Z(n6812)
         );
  AOI211_X1 U8539 ( .C1(n6813), .C2(n6812), .A(n6878), .B(n9761), .ZN(n6814)
         );
  AOI211_X1 U8540 ( .C1(P2_ADDR_REG_9__SCAN_IN), .C2(n9766), .A(n6815), .B(
        n6814), .ZN(n6822) );
  OAI21_X1 U8541 ( .B1(n6817), .B2(n7522), .A(n6816), .ZN(n6820) );
  MUX2_X1 U8542 ( .A(n7507), .B(P2_REG2_REG_9__SCAN_IN), .S(n6883), .Z(n6818)
         );
  INV_X1 U8543 ( .A(n6818), .ZN(n6819) );
  NAND2_X1 U8544 ( .A1(n6819), .A2(n6820), .ZN(n6884) );
  OAI211_X1 U8545 ( .C1(n6820), .C2(n6819), .A(n9764), .B(n6884), .ZN(n6821)
         );
  OAI211_X1 U8546 ( .C1(n9760), .C2(n6823), .A(n6822), .B(n6821), .ZN(P2_U3254) );
  INV_X1 U8547 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n6836) );
  OAI21_X1 U8548 ( .B1(n6826), .B2(n6825), .A(n6824), .ZN(n6827) );
  NAND2_X1 U8549 ( .A1(n6827), .A2(n9593), .ZN(n6835) );
  NAND2_X1 U8550 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n7670) );
  INV_X1 U8551 ( .A(n7670), .ZN(n6832) );
  AOI211_X1 U8552 ( .C1(n6830), .C2(n6829), .A(n6828), .B(n9598), .ZN(n6831)
         );
  AOI211_X1 U8553 ( .C1(n9585), .C2(n6833), .A(n6832), .B(n6831), .ZN(n6834)
         );
  OAI211_X1 U8554 ( .C1(n9619), .C2(n6836), .A(n6835), .B(n6834), .ZN(P1_U3253) );
  INV_X1 U8555 ( .A(n6837), .ZN(n6839) );
  INV_X1 U8556 ( .A(n8597), .ZN(n8588) );
  OAI222_X1 U8557 ( .A1(n8459), .A2(n6838), .B1(n4390), .B2(n6839), .C1(
        P2_U3152), .C2(n8588), .ZN(P2_U3343) );
  OAI222_X1 U8558 ( .A1(n8421), .A2(n6840), .B1(n8419), .B2(n6839), .C1(
        P1_U3084), .C2(n7611), .ZN(P1_U3338) );
  INV_X1 U8559 ( .A(n6841), .ZN(n6877) );
  AOI22_X1 U8560 ( .A1(n8613), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n8014), .ZN(n6842) );
  OAI21_X1 U8561 ( .B1(n6877), .B2(n4390), .A(n6842), .ZN(P2_U3342) );
  NAND2_X1 U8562 ( .A1(n8113), .A2(n9127), .ZN(n6848) );
  NAND2_X1 U8563 ( .A1(n6707), .A2(n9688), .ZN(n6847) );
  NAND2_X1 U8564 ( .A1(n6848), .A2(n6847), .ZN(n6849) );
  XNOR2_X1 U8565 ( .A(n6849), .B(n8062), .ZN(n6852) );
  OAI22_X1 U8566 ( .A1(n8101), .A2(n9659), .B1(n7186), .B2(n6851), .ZN(n6853)
         );
  XNOR2_X1 U8567 ( .A(n6852), .B(n6853), .ZN(n9063) );
  NAND2_X1 U8568 ( .A1(n9060), .A2(n9063), .ZN(n9061) );
  INV_X1 U8569 ( .A(n6852), .ZN(n6854) );
  NAND2_X1 U8570 ( .A1(n6854), .A2(n6853), .ZN(n6855) );
  NAND2_X1 U8571 ( .A1(n9061), .A2(n6855), .ZN(n6905) );
  NAND2_X1 U8572 ( .A1(n8113), .A2(n9126), .ZN(n6857) );
  NAND2_X1 U8573 ( .A1(n6707), .A2(n9651), .ZN(n6856) );
  NAND2_X1 U8574 ( .A1(n6857), .A2(n6856), .ZN(n6858) );
  XNOR2_X1 U8575 ( .A(n6858), .B(n8062), .ZN(n6903) );
  XNOR2_X1 U8576 ( .A(n6905), .B(n6903), .ZN(n6860) );
  AOI22_X1 U8577 ( .A1(n6764), .A2(n9126), .B1(n8113), .B2(n9651), .ZN(n6861)
         );
  NAND2_X1 U8578 ( .A1(n6860), .A2(n6861), .ZN(n6907) );
  OAI21_X1 U8579 ( .B1(n6859), .B2(n6861), .A(n6907), .ZN(n6866) );
  INV_X1 U8580 ( .A(n9095), .ZN(n9102) );
  AOI22_X1 U8581 ( .A1(n9089), .A2(n9652), .B1(n7915), .B2(n9127), .ZN(n6864)
         );
  AOI21_X1 U8582 ( .B1(n9088), .B2(n9125), .A(n6862), .ZN(n6863) );
  OAI211_X1 U8583 ( .C1(n9698), .C2(n9115), .A(n6864), .B(n6863), .ZN(n6865)
         );
  AOI21_X1 U8584 ( .B1(n6866), .B2(n9102), .A(n6865), .ZN(n6867) );
  INV_X1 U8585 ( .A(n6867), .ZN(P1_U3225) );
  OAI21_X1 U8586 ( .B1(n6870), .B2(n6869), .A(n6868), .ZN(n6874) );
  INV_X1 U8587 ( .A(n9743), .ZN(n8544) );
  AND2_X1 U8588 ( .A1(n8529), .A2(n7257), .ZN(n8425) );
  OAI22_X1 U8589 ( .A1(n8425), .A2(n6871), .B1(n9747), .B2(n7008), .ZN(n6873)
         );
  OAI22_X1 U8590 ( .A1(n8422), .A2(n9751), .B1(n9750), .B2(n6159), .ZN(n6872)
         );
  AOI211_X1 U8591 ( .C1(n6874), .C2(n8544), .A(n6873), .B(n6872), .ZN(n6875)
         );
  INV_X1 U8592 ( .A(n6875), .ZN(P2_U3224) );
  INV_X1 U8593 ( .A(n7805), .ZN(n7618) );
  OAI222_X1 U8594 ( .A1(n8419), .A2(n6877), .B1(n7618), .B2(P1_U3084), .C1(
        n6876), .C2(n8421), .ZN(P1_U3337) );
  NAND2_X1 U8595 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n7558) );
  INV_X1 U8596 ( .A(n7558), .ZN(n6882) );
  INV_X1 U8597 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6879) );
  MUX2_X1 U8598 ( .A(n6879), .B(P2_REG1_REG_10__SCAN_IN), .S(n6964), .Z(n6880)
         );
  NOR2_X1 U8599 ( .A1(n4421), .A2(n6880), .ZN(n6963) );
  AOI211_X1 U8600 ( .C1(n4421), .C2(n6880), .A(n6963), .B(n9761), .ZN(n6881)
         );
  AOI211_X1 U8601 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n9766), .A(n6882), .B(
        n6881), .ZN(n6890) );
  NAND2_X1 U8602 ( .A1(n6883), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6885) );
  NAND2_X1 U8603 ( .A1(n6885), .A2(n6884), .ZN(n6888) );
  MUX2_X1 U8604 ( .A(n7595), .B(P2_REG2_REG_10__SCAN_IN), .S(n6964), .Z(n6886)
         );
  INV_X1 U8605 ( .A(n6886), .ZN(n6887) );
  NAND2_X1 U8606 ( .A1(n6887), .A2(n6888), .ZN(n6957) );
  OAI211_X1 U8607 ( .C1(n6888), .C2(n6887), .A(n9764), .B(n6957), .ZN(n6889)
         );
  OAI211_X1 U8608 ( .C1(n9760), .C2(n6891), .A(n6890), .B(n6889), .ZN(P2_U3255) );
  INV_X1 U8609 ( .A(n6892), .ZN(n6893) );
  AOI21_X1 U8610 ( .B1(n8022), .B2(n6893), .A(n9743), .ZN(n6897) );
  NOR2_X1 U8611 ( .A1(n9743), .A2(n6894), .ZN(n8533) );
  INV_X1 U8612 ( .A(n8533), .ZN(n8552) );
  NOR3_X1 U8613 ( .A1(n8552), .A2(n6895), .A3(n6159), .ZN(n6896) );
  OAI21_X1 U8614 ( .B1(n6897), .B2(n6896), .A(n8543), .ZN(n6901) );
  OAI22_X1 U8615 ( .A1(n6159), .A2(n8880), .B1(n9752), .B2(n8882), .ZN(n6997)
         );
  INV_X1 U8616 ( .A(n8508), .ZN(n8523) );
  AOI22_X1 U8617 ( .A1(n6997), .A2(n8523), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        P2_U3152), .ZN(n6898) );
  OAI21_X1 U8618 ( .B1(n7117), .B2(n9747), .A(n6898), .ZN(n6899) );
  AOI21_X1 U8619 ( .B1(n8511), .B2(n5252), .A(n6899), .ZN(n6900) );
  NAND2_X1 U8620 ( .A1(n6901), .A2(n6900), .ZN(P2_U3220) );
  INV_X1 U8621 ( .A(n6902), .ZN(n6929) );
  INV_X1 U8622 ( .A(n9163), .ZN(n7809) );
  OAI222_X1 U8623 ( .A1(n8419), .A2(n6929), .B1(n7809), .B2(P1_U3084), .C1(
        n10161), .C2(n8421), .ZN(P1_U3336) );
  INV_X1 U8624 ( .A(n6903), .ZN(n6904) );
  OR2_X1 U8625 ( .A1(n6905), .A2(n6904), .ZN(n6906) );
  NAND2_X1 U8626 ( .A1(n6907), .A2(n6906), .ZN(n6934) );
  NAND2_X1 U8627 ( .A1(n7059), .A2(n6707), .ZN(n6909) );
  NAND2_X1 U8628 ( .A1(n8113), .A2(n9125), .ZN(n6908) );
  NAND2_X1 U8629 ( .A1(n6909), .A2(n6908), .ZN(n6910) );
  XNOR2_X1 U8630 ( .A(n6910), .B(n8062), .ZN(n6935) );
  NAND2_X1 U8631 ( .A1(n7059), .A2(n8113), .ZN(n6911) );
  OAI21_X1 U8632 ( .B1(n8101), .B2(n9661), .A(n6911), .ZN(n6936) );
  XNOR2_X1 U8633 ( .A(n6935), .B(n6936), .ZN(n6933) );
  XOR2_X1 U8634 ( .A(n6934), .B(n6933), .Z(n6916) );
  INV_X1 U8635 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6912) );
  NOR2_X1 U8636 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6912), .ZN(n9591) );
  OAI22_X1 U8637 ( .A1(n9108), .A2(n7056), .B1(n9638), .B2(n9106), .ZN(n6913)
         );
  AOI211_X1 U8638 ( .C1(n7915), .C2(n9126), .A(n9591), .B(n6913), .ZN(n6915)
         );
  INV_X1 U8639 ( .A(n7059), .ZN(n7055) );
  NOR2_X1 U8640 ( .A1(n7055), .A2(n9718), .ZN(n9703) );
  NAND2_X1 U8641 ( .A1(n6947), .A2(n9703), .ZN(n6914) );
  OAI211_X1 U8642 ( .C1(n6916), .C2(n9095), .A(n6915), .B(n6914), .ZN(P1_U3237) );
  INV_X1 U8643 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6928) );
  OAI21_X1 U8644 ( .B1(n6919), .B2(n6918), .A(n6917), .ZN(n6920) );
  NAND2_X1 U8645 ( .A1(n6920), .A2(n9593), .ZN(n6927) );
  AND2_X1 U8646 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7705) );
  AOI211_X1 U8647 ( .C1(n6923), .C2(n6922), .A(n6921), .B(n9598), .ZN(n6924)
         );
  AOI211_X1 U8648 ( .C1(n9585), .C2(n6925), .A(n7705), .B(n6924), .ZN(n6926)
         );
  OAI211_X1 U8649 ( .C1(n9619), .C2(n6928), .A(n6927), .B(n6926), .ZN(P1_U3254) );
  INV_X1 U8650 ( .A(n8630), .ZN(n8612) );
  OAI222_X1 U8651 ( .A1(n8459), .A2(n6930), .B1(n4390), .B2(n6929), .C1(n8612), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U8652 ( .A(n6931), .ZN(n6956) );
  AOI22_X1 U8653 ( .A1(n9175), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n8008), .ZN(n6932) );
  OAI21_X1 U8654 ( .B1(n6956), .B2(n8419), .A(n6932), .ZN(P1_U3335) );
  NAND2_X1 U8655 ( .A1(n6934), .A2(n6933), .ZN(n6939) );
  INV_X1 U8656 ( .A(n6935), .ZN(n6937) );
  OR2_X1 U8657 ( .A1(n6937), .A2(n6936), .ZN(n6938) );
  NAND2_X1 U8658 ( .A1(n7036), .A2(n8113), .ZN(n6941) );
  NAND2_X1 U8659 ( .A1(n6764), .A2(n9124), .ZN(n6940) );
  AND2_X1 U8660 ( .A1(n6941), .A2(n6940), .ZN(n7066) );
  NAND2_X1 U8661 ( .A1(n7036), .A2(n6707), .ZN(n6943) );
  NAND2_X1 U8662 ( .A1(n8113), .A2(n9124), .ZN(n6942) );
  NAND2_X1 U8663 ( .A1(n6943), .A2(n6942), .ZN(n6944) );
  XOR2_X1 U8664 ( .A(n7066), .B(n7064), .Z(n6945) );
  XNOR2_X1 U8665 ( .A(n7065), .B(n6945), .ZN(n6950) );
  AND2_X1 U8666 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9147) );
  OAI22_X1 U8667 ( .A1(n9108), .A2(n7033), .B1(n7027), .B2(n9106), .ZN(n6946)
         );
  AOI211_X1 U8668 ( .C1(n7915), .C2(n9125), .A(n9147), .B(n6946), .ZN(n6949)
         );
  AND2_X1 U8669 ( .A1(n7036), .A2(n9689), .ZN(n9714) );
  NAND2_X1 U8670 ( .A1(n6947), .A2(n9714), .ZN(n6948) );
  OAI211_X1 U8671 ( .C1(n6950), .C2(n9095), .A(n6949), .B(n6948), .ZN(P1_U3211) );
  OAI21_X1 U8672 ( .B1(n9531), .B2(n9337), .A(n6951), .ZN(n6954) );
  AOI22_X1 U8673 ( .A1(n6952), .A2(n9665), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n9653), .ZN(n6953) );
  OAI211_X1 U8674 ( .C1(n5748), .C2(n9665), .A(n6954), .B(n6953), .ZN(P1_U3291) );
  INV_X1 U8675 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10153) );
  INV_X1 U8676 ( .A(n8643), .ZN(n6955) );
  OAI222_X1 U8677 ( .A1(n8459), .A2(n10153), .B1(n4390), .B2(n6956), .C1(
        P2_U3152), .C2(n6955), .ZN(P2_U3340) );
  NAND2_X1 U8678 ( .A1(n6964), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6958) );
  NAND2_X1 U8679 ( .A1(n6958), .A2(n6957), .ZN(n6961) );
  MUX2_X1 U8680 ( .A(n6959), .B(P2_REG2_REG_11__SCAN_IN), .S(n7078), .Z(n6960)
         );
  NOR2_X1 U8681 ( .A1(n6961), .A2(n6960), .ZN(n7086) );
  AOI21_X1 U8682 ( .B1(n6961), .B2(n6960), .A(n7086), .ZN(n6973) );
  INV_X1 U8683 ( .A(n9764), .ZN(n8633) );
  INV_X1 U8684 ( .A(n9761), .ZN(n9763) );
  INV_X1 U8685 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6962) );
  MUX2_X1 U8686 ( .A(n6962), .B(P2_REG1_REG_11__SCAN_IN), .S(n7078), .Z(n6966)
         );
  AOI21_X1 U8687 ( .B1(n6966), .B2(n6965), .A(n7077), .ZN(n6967) );
  NAND2_X1 U8688 ( .A1(n9763), .A2(n6967), .ZN(n6970) );
  NOR2_X1 U8689 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7686), .ZN(n6968) );
  AOI21_X1 U8690 ( .B1(n9766), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n6968), .ZN(
        n6969) );
  OAI211_X1 U8691 ( .C1(n9760), .C2(n7087), .A(n6970), .B(n6969), .ZN(n6971)
         );
  INV_X1 U8692 ( .A(n6971), .ZN(n6972) );
  OAI21_X1 U8693 ( .B1(n6973), .B2(n8633), .A(n6972), .ZN(P2_U3256) );
  XNOR2_X1 U8694 ( .A(n6980), .B(n6974), .ZN(n9805) );
  NAND3_X1 U8695 ( .A1(n7257), .A2(n6975), .A3(n7268), .ZN(n6990) );
  XNOR2_X1 U8696 ( .A(n6978), .B(n6976), .ZN(n6977) );
  NAND2_X1 U8697 ( .A1(n6977), .A2(n8649), .ZN(n7842) );
  OR2_X1 U8698 ( .A1(n6978), .A2(n8649), .ZN(n7504) );
  NAND2_X1 U8699 ( .A1(n7842), .A2(n7504), .ZN(n6979) );
  NAND2_X1 U8700 ( .A1(n8870), .A2(n6979), .ZN(n8862) );
  XNOR2_X1 U8701 ( .A(n6981), .B(n6980), .ZN(n6986) );
  NAND2_X1 U8702 ( .A1(n6983), .A2(n6982), .ZN(n9777) );
  NAND2_X1 U8703 ( .A1(n6209), .A2(n9772), .ZN(n6984) );
  OAI21_X1 U8704 ( .B1(n6159), .B2(n8882), .A(n6984), .ZN(n6985) );
  AOI21_X1 U8705 ( .B1(n6986), .B2(n9777), .A(n6985), .ZN(n9806) );
  MUX2_X1 U8706 ( .A(n6987), .B(n9806), .S(n8870), .Z(n6995) );
  NOR2_X1 U8707 ( .A1(n5632), .A2(n9801), .ZN(n6988) );
  NAND2_X1 U8708 ( .A1(n8870), .A2(n6988), .ZN(n8851) );
  OR2_X1 U8709 ( .A1(n6990), .A2(n6989), .ZN(n8874) );
  NAND2_X1 U8710 ( .A1(n8851), .A2(n8874), .ZN(n9786) );
  AND2_X1 U8711 ( .A1(n9819), .A2(n8426), .ZN(n6993) );
  INV_X1 U8712 ( .A(n9818), .ZN(n9851) );
  OAI21_X1 U8713 ( .B1(n8426), .B2(n9853), .A(n9851), .ZN(n6992) );
  MUX2_X1 U8714 ( .A(n6993), .B(n6992), .S(n7098), .Z(n9808) );
  INV_X1 U8715 ( .A(n9778), .ZN(n8848) );
  AOI22_X1 U8716 ( .A1(n9786), .A2(n9808), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8848), .ZN(n6994) );
  OAI211_X1 U8717 ( .C1(n9805), .C2(n8862), .A(n6995), .B(n6994), .ZN(P2_U3295) );
  XNOR2_X1 U8718 ( .A(n6996), .B(n7007), .ZN(n6998) );
  AOI21_X1 U8719 ( .B1(n6998), .B2(n9777), .A(n6997), .ZN(n9822) );
  MUX2_X1 U8720 ( .A(n9822), .B(n6999), .S(n4388), .Z(n7013) );
  NAND2_X1 U8721 ( .A1(n7001), .A2(n7000), .ZN(n7004) );
  NAND2_X1 U8722 ( .A1(n7002), .A2(n7008), .ZN(n7003) );
  NAND2_X1 U8723 ( .A1(n7004), .A2(n7003), .ZN(n7093) );
  NAND2_X1 U8724 ( .A1(n7093), .A2(n7094), .ZN(n7006) );
  NAND2_X1 U8725 ( .A1(n6159), .A2(n9811), .ZN(n7005) );
  NAND2_X1 U8726 ( .A1(n7006), .A2(n7005), .ZN(n7116) );
  XNOR2_X1 U8727 ( .A(n7116), .B(n7007), .ZN(n9823) );
  INV_X1 U8728 ( .A(n9823), .ZN(n9826) );
  INV_X1 U8729 ( .A(n8862), .ZN(n9787) );
  NAND2_X1 U8730 ( .A1(n7100), .A2(n9817), .ZN(n7009) );
  AND2_X1 U8731 ( .A1(n7111), .A2(n7009), .ZN(n9820) );
  AOI22_X1 U8732 ( .A1(n9820), .A2(n8834), .B1(n8848), .B2(n5252), .ZN(n7010)
         );
  OAI21_X1 U8733 ( .B1(n7117), .B2(n8851), .A(n7010), .ZN(n7011) );
  AOI21_X1 U8734 ( .B1(n9826), .B2(n9787), .A(n7011), .ZN(n7012) );
  NAND2_X1 U8735 ( .A1(n7013), .A2(n7012), .ZN(P2_U3293) );
  INV_X1 U8736 ( .A(n7014), .ZN(n7016) );
  OAI222_X1 U8737 ( .A1(n8459), .A2(n7015), .B1(n4390), .B2(n7016), .C1(
        P2_U3152), .C2(n8649), .ZN(P2_U3339) );
  OAI222_X1 U8738 ( .A1(n8421), .A2(n7017), .B1(n8419), .B2(n7016), .C1(n9350), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  AOI22_X1 U8739 ( .A1(n9803), .A2(n9777), .B1(n9774), .B2(n6157), .ZN(n9799)
         );
  OAI21_X1 U8740 ( .B1(n7018), .B2(n9778), .A(n9799), .ZN(n7019) );
  AOI22_X1 U8741 ( .A1(n7019), .A2(n8870), .B1(n8426), .B2(n9786), .ZN(n7021)
         );
  AOI22_X1 U8742 ( .A1(n9787), .A2(n9803), .B1(P2_REG2_REG_0__SCAN_IN), .B2(
        n4388), .ZN(n7020) );
  NAND2_X1 U8743 ( .A1(n7021), .A2(n7020), .ZN(P2_U3296) );
  AND2_X1 U8744 ( .A1(n7022), .A2(n8316), .ZN(n8309) );
  NAND2_X1 U8745 ( .A1(n7023), .A2(n8309), .ZN(n7024) );
  NAND2_X1 U8746 ( .A1(n7024), .A2(n8322), .ZN(n7025) );
  XNOR2_X1 U8747 ( .A(n7025), .B(n7031), .ZN(n7026) );
  NAND2_X1 U8748 ( .A1(n7026), .A2(n9635), .ZN(n7030) );
  OAI22_X1 U8749 ( .A1(n9661), .A2(n9660), .B1(n9662), .B2(n7027), .ZN(n7028)
         );
  INV_X1 U8750 ( .A(n7028), .ZN(n7029) );
  NAND2_X1 U8751 ( .A1(n7030), .A2(n7029), .ZN(n9712) );
  XNOR2_X1 U8752 ( .A(n7032), .B(n7031), .ZN(n9711) );
  OAI22_X1 U8753 ( .A1(n9665), .A2(n7034), .B1(n7033), .B2(n9629), .ZN(n7035)
         );
  AOI21_X1 U8754 ( .B1(n9531), .B2(n7036), .A(n7035), .ZN(n7041) );
  INV_X1 U8755 ( .A(n9705), .ZN(n9690) );
  OAI21_X1 U8756 ( .B1(n7052), .B2(n7037), .A(n9690), .ZN(n7038) );
  NOR2_X1 U8757 ( .A1(n7038), .A2(n9627), .ZN(n9713) );
  OR2_X1 U8758 ( .A1(n7039), .A2(n4486), .ZN(n9516) );
  INV_X1 U8759 ( .A(n9516), .ZN(n9539) );
  NAND2_X1 U8760 ( .A1(n9713), .A2(n9539), .ZN(n7040) );
  OAI211_X1 U8761 ( .C1(n9711), .C2(n9374), .A(n7041), .B(n7040), .ZN(n7042)
         );
  AOI21_X1 U8762 ( .B1(n9665), .B2(n9712), .A(n7042), .ZN(n7043) );
  INV_X1 U8763 ( .A(n7043), .ZN(P1_U3284) );
  XNOR2_X1 U8764 ( .A(n7044), .B(n7046), .ZN(n9709) );
  INV_X1 U8765 ( .A(n9709), .ZN(n7063) );
  OAI211_X1 U8766 ( .C1(n7047), .C2(n7046), .A(n7045), .B(n9635), .ZN(n7051)
         );
  OAI22_X1 U8767 ( .A1(n9638), .A2(n9662), .B1(n9660), .B2(n7048), .ZN(n7049)
         );
  INV_X1 U8768 ( .A(n7049), .ZN(n7050) );
  NAND2_X1 U8769 ( .A1(n7051), .A2(n7050), .ZN(n9707) );
  INV_X1 U8770 ( .A(n9649), .ZN(n7054) );
  INV_X1 U8771 ( .A(n7052), .ZN(n7053) );
  OAI21_X1 U8772 ( .B1(n7055), .B2(n7054), .A(n7053), .ZN(n9706) );
  INV_X1 U8773 ( .A(n9337), .ZN(n9198) );
  OAI22_X1 U8774 ( .A1(n9665), .A2(n7057), .B1(n7056), .B2(n9629), .ZN(n7058)
         );
  AOI21_X1 U8775 ( .B1(n9531), .B2(n7059), .A(n7058), .ZN(n7060) );
  OAI21_X1 U8776 ( .B1(n9706), .B2(n9198), .A(n7060), .ZN(n7061) );
  AOI21_X1 U8777 ( .B1(n9707), .B2(n9665), .A(n7061), .ZN(n7062) );
  OAI21_X1 U8778 ( .B1(n7063), .B2(n9374), .A(n7062), .ZN(P1_U3285) );
  NAND2_X1 U8779 ( .A1(n9631), .A2(n6707), .ZN(n7068) );
  NAND2_X1 U8780 ( .A1(n8113), .A2(n9123), .ZN(n7067) );
  NAND2_X1 U8781 ( .A1(n7068), .A2(n7067), .ZN(n7069) );
  XNOR2_X1 U8782 ( .A(n7069), .B(n6738), .ZN(n7282) );
  NAND2_X1 U8783 ( .A1(n9631), .A2(n8113), .ZN(n7071) );
  NAND2_X1 U8784 ( .A1(n6764), .A2(n9123), .ZN(n7070) );
  NAND2_X1 U8785 ( .A1(n7071), .A2(n7070), .ZN(n7283) );
  XNOR2_X1 U8786 ( .A(n7282), .B(n7283), .ZN(n7072) );
  XNOR2_X1 U8787 ( .A(n7284), .B(n7072), .ZN(n7073) );
  NAND2_X1 U8788 ( .A1(n7073), .A2(n9102), .ZN(n7076) );
  INV_X1 U8789 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10106) );
  NOR2_X1 U8790 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10106), .ZN(n9613) );
  OAI22_X1 U8791 ( .A1(n9108), .A2(n9628), .B1(n9637), .B2(n9106), .ZN(n7074)
         );
  AOI211_X1 U8792 ( .C1(n7915), .C2(n9124), .A(n9613), .B(n7074), .ZN(n7075)
         );
  OAI211_X1 U8793 ( .C1(n9719), .C2(n9115), .A(n7076), .B(n7075), .ZN(P1_U3219) );
  INV_X1 U8794 ( .A(n7240), .ZN(n7092) );
  MUX2_X1 U8795 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7079), .S(n7240), .Z(n7080)
         );
  OAI21_X1 U8796 ( .B1(n7081), .B2(n7080), .A(n7239), .ZN(n7085) );
  NAND2_X1 U8797 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7773) );
  INV_X1 U8798 ( .A(n7773), .ZN(n7084) );
  INV_X1 U8799 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7082) );
  NOR2_X1 U8800 ( .A1(n8655), .A2(n7082), .ZN(n7083) );
  AOI211_X1 U8801 ( .C1(n9763), .C2(n7085), .A(n7084), .B(n7083), .ZN(n7091)
         );
  AOI21_X1 U8802 ( .B1(n7087), .B2(n6959), .A(n7086), .ZN(n7089) );
  MUX2_X1 U8803 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n7791), .S(n7240), .Z(n7088)
         );
  NAND2_X1 U8804 ( .A1(n7240), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7236) );
  OAI211_X1 U8805 ( .C1(n7240), .C2(P2_REG2_REG_12__SCAN_IN), .A(n7089), .B(
        n7236), .ZN(n7235) );
  OAI211_X1 U8806 ( .C1(n7089), .C2(n7088), .A(n9764), .B(n7235), .ZN(n7090)
         );
  OAI211_X1 U8807 ( .C1(n9760), .C2(n7092), .A(n7091), .B(n7090), .ZN(P2_U3257) );
  XOR2_X1 U8808 ( .A(n7093), .B(n7094), .Z(n9810) );
  XNOR2_X1 U8809 ( .A(n7095), .B(n7094), .ZN(n7096) );
  AOI222_X1 U8810 ( .A1(n9777), .A2(n7096), .B1(n6157), .B2(n9772), .C1(n8585), 
        .C2(n9774), .ZN(n9813) );
  MUX2_X1 U8811 ( .A(n7097), .B(n9813), .S(n8870), .Z(n7104) );
  OAI21_X1 U8812 ( .B1(n7098), .B2(n8426), .A(n7102), .ZN(n7099) );
  NAND2_X1 U8813 ( .A1(n7100), .A2(n7099), .ZN(n9812) );
  OAI22_X1 U8814 ( .A1(n9812), .A2(n8874), .B1(n8026), .B2(n9778), .ZN(n7101)
         );
  AOI21_X1 U8815 ( .B1(n8872), .B2(n7102), .A(n7101), .ZN(n7103) );
  OAI211_X1 U8816 ( .C1(n9810), .C2(n8862), .A(n7104), .B(n7103), .ZN(P2_U3294) );
  NAND2_X1 U8817 ( .A1(n7106), .A2(n7222), .ZN(n7107) );
  NAND3_X1 U8818 ( .A1(n7105), .A2(n9777), .A3(n7107), .ZN(n7109) );
  AOI22_X1 U8819 ( .A1(n9773), .A2(n9774), .B1(n9772), .B2(n8585), .ZN(n7108)
         );
  AND2_X1 U8820 ( .A1(n7109), .A2(n7108), .ZN(n9834) );
  OAI22_X1 U8821 ( .A1(n8870), .A2(n7110), .B1(n8546), .B2(n9778), .ZN(n7114)
         );
  AND2_X1 U8822 ( .A1(n7111), .A2(n8550), .ZN(n7112) );
  OR2_X1 U8823 ( .A1(n7112), .A2(n7230), .ZN(n9831) );
  NOR2_X1 U8824 ( .A1(n9831), .A2(n8874), .ZN(n7113) );
  AOI211_X1 U8825 ( .C1(n8872), .C2(n8550), .A(n7114), .B(n7113), .ZN(n7121)
         );
  NAND2_X1 U8826 ( .A1(n7116), .A2(n7115), .ZN(n7119) );
  NAND2_X1 U8827 ( .A1(n8027), .A2(n7117), .ZN(n7118) );
  NAND2_X1 U8828 ( .A1(n7119), .A2(n7118), .ZN(n7223) );
  XNOR2_X1 U8829 ( .A(n7222), .B(n7223), .ZN(n9829) );
  NAND2_X1 U8830 ( .A1(n9829), .A2(n9787), .ZN(n7120) );
  OAI211_X1 U8831 ( .C1(n9834), .C2(n4388), .A(n7121), .B(n7120), .ZN(P2_U3292) );
  INV_X1 U8832 ( .A(n7122), .ZN(n7154) );
  AND2_X1 U8833 ( .A1(n7295), .A2(n8160), .ZN(n8263) );
  XNOR2_X1 U8834 ( .A(n7124), .B(n8263), .ZN(n7314) );
  OR2_X1 U8835 ( .A1(n7125), .A2(n6692), .ZN(n7128) );
  OR2_X1 U8836 ( .A1(n7126), .A2(n7312), .ZN(n7127) );
  AND2_X1 U8837 ( .A1(n7128), .A2(n7127), .ZN(n9378) );
  INV_X1 U8838 ( .A(n9378), .ZN(n7731) );
  XNOR2_X1 U8839 ( .A(n7297), .B(n8263), .ZN(n7130) );
  INV_X1 U8840 ( .A(n9635), .ZN(n9657) );
  INV_X1 U8841 ( .A(n9660), .ZN(n9526) );
  INV_X1 U8842 ( .A(n9662), .ZN(n9524) );
  AOI22_X1 U8843 ( .A1(n9526), .A2(n9123), .B1(n9524), .B2(n9121), .ZN(n7129)
         );
  OAI21_X1 U8844 ( .B1(n7130), .B2(n9657), .A(n7129), .ZN(n7131) );
  AOI21_X1 U8845 ( .B1(n7314), .B2(n7731), .A(n7131), .ZN(n7318) );
  AOI21_X1 U8846 ( .B1(n7315), .B2(n9626), .A(n4688), .ZN(n7316) );
  INV_X1 U8847 ( .A(n7315), .ZN(n7132) );
  NOR2_X1 U8848 ( .A1(n7132), .A2(n9370), .ZN(n7135) );
  INV_X1 U8849 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7133) );
  OAI22_X1 U8850 ( .A1(n9665), .A2(n7133), .B1(n7289), .B2(n9629), .ZN(n7134)
         );
  AOI211_X1 U8851 ( .C1(n7316), .C2(n9337), .A(n7135), .B(n7134), .ZN(n7137)
         );
  NOR3_X1 U8852 ( .A1(n4389), .A2(n9350), .A3(n6691), .ZN(n7737) );
  NAND2_X1 U8853 ( .A1(n7314), .A2(n7737), .ZN(n7136) );
  OAI211_X1 U8854 ( .C1(n7318), .C2(n4389), .A(n7137), .B(n7136), .ZN(P1_U3282) );
  INV_X1 U8855 ( .A(n7737), .ZN(n7208) );
  INV_X1 U8856 ( .A(n7139), .ZN(n7140) );
  NAND2_X1 U8857 ( .A1(n8255), .A2(n7140), .ZN(n7141) );
  NAND2_X1 U8858 ( .A1(n7138), .A2(n7141), .ZN(n9669) );
  AOI22_X1 U8859 ( .A1(n9531), .A2(n7142), .B1(n4389), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7153) );
  AOI22_X1 U8860 ( .A1(n9526), .A2(n6695), .B1(n9524), .B2(n9129), .ZN(n7147)
         );
  OAI21_X1 U8861 ( .B1(n7144), .B2(n8255), .A(n7143), .ZN(n7145) );
  NAND2_X1 U8862 ( .A1(n7145), .A2(n9635), .ZN(n7146) );
  OAI211_X1 U8863 ( .C1(n9669), .C2(n9378), .A(n7147), .B(n7146), .ZN(n9672)
         );
  OAI21_X1 U8864 ( .B1(n9671), .B2(n7148), .A(n7200), .ZN(n7149) );
  OR2_X1 U8865 ( .A1(n9705), .A2(n7149), .ZN(n9670) );
  OAI22_X1 U8866 ( .A1(n9629), .A2(n7150), .B1(n9670), .B2(n4486), .ZN(n7151)
         );
  OAI21_X1 U8867 ( .B1(n9672), .B2(n7151), .A(n9665), .ZN(n7152) );
  OAI211_X1 U8868 ( .C1(n7208), .C2(n9669), .A(n7153), .B(n7152), .ZN(P1_U3290) );
  OAI222_X1 U8869 ( .A1(n8459), .A2(n9957), .B1(n4390), .B2(n7154), .C1(n5632), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  NAND2_X1 U8870 ( .A1(n7155), .A2(n7156), .ZN(n7172) );
  XNOR2_X1 U8871 ( .A(n7172), .B(n8253), .ZN(n9686) );
  INV_X1 U8872 ( .A(n9686), .ZN(n7171) );
  NAND2_X1 U8873 ( .A1(n9686), .A2(n7731), .ZN(n7164) );
  OAI21_X1 U8874 ( .B1(n7159), .B2(n7157), .A(n7158), .ZN(n7162) );
  OAI22_X1 U8875 ( .A1(n9659), .A2(n9662), .B1(n9660), .B2(n7160), .ZN(n7161)
         );
  AOI21_X1 U8876 ( .B1(n7162), .B2(n9635), .A(n7161), .ZN(n7163) );
  NAND2_X1 U8877 ( .A1(n7164), .A2(n7163), .ZN(n9684) );
  MUX2_X1 U8878 ( .A(n9684), .B(P1_REG2_REG_3__SCAN_IN), .S(n4389), .Z(n7165)
         );
  INV_X1 U8879 ( .A(n7165), .ZN(n7170) );
  AND2_X1 U8880 ( .A1(n7202), .A2(n7166), .ZN(n7167) );
  NOR2_X1 U8881 ( .A1(n7183), .A2(n7167), .ZN(n9681) );
  OAI22_X1 U8882 ( .A1(n9370), .A2(n9683), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9629), .ZN(n7168) );
  AOI21_X1 U8883 ( .B1(n9337), .B2(n9681), .A(n7168), .ZN(n7169) );
  OAI211_X1 U8884 ( .C1(n7171), .C2(n7208), .A(n7170), .B(n7169), .ZN(P1_U3288) );
  NAND2_X1 U8885 ( .A1(n7172), .A2(n8253), .ZN(n7174) );
  NAND2_X1 U8886 ( .A1(n7174), .A2(n7173), .ZN(n7175) );
  XNOR2_X1 U8887 ( .A(n7177), .B(n7175), .ZN(n7181) );
  INV_X1 U8888 ( .A(n7181), .ZN(n9695) );
  XNOR2_X1 U8889 ( .A(n7177), .B(n7176), .ZN(n7179) );
  AOI22_X1 U8890 ( .A1(n9524), .A2(n9126), .B1(n9526), .B2(n9128), .ZN(n7178)
         );
  OAI21_X1 U8891 ( .B1(n7179), .B2(n9657), .A(n7178), .ZN(n7180) );
  AOI21_X1 U8892 ( .B1(n7731), .B2(n7181), .A(n7180), .ZN(n9693) );
  MUX2_X1 U8893 ( .A(n7182), .B(n9693), .S(n9665), .Z(n7189) );
  INV_X1 U8894 ( .A(n7183), .ZN(n7185) );
  INV_X1 U8895 ( .A(n9648), .ZN(n7184) );
  AOI21_X1 U8896 ( .B1(n9688), .B2(n7185), .A(n7184), .ZN(n9691) );
  OAI22_X1 U8897 ( .A1(n9370), .A2(n7186), .B1(n9064), .B2(n9629), .ZN(n7187)
         );
  AOI21_X1 U8898 ( .B1(n9337), .B2(n9691), .A(n7187), .ZN(n7188) );
  OAI211_X1 U8899 ( .C1(n9695), .C2(n7208), .A(n7189), .B(n7188), .ZN(P1_U3287) );
  INV_X1 U8900 ( .A(n7155), .ZN(n7190) );
  AOI21_X1 U8901 ( .B1(n7193), .B2(n7191), .A(n7190), .ZN(n9675) );
  OAI21_X1 U8902 ( .B1(n7193), .B2(n8373), .A(n7192), .ZN(n7196) );
  OAI22_X1 U8903 ( .A1(n9066), .A2(n9662), .B1(n9660), .B2(n7194), .ZN(n7195)
         );
  AOI21_X1 U8904 ( .B1(n7196), .B2(n9635), .A(n7195), .ZN(n7197) );
  OAI21_X1 U8905 ( .B1(n9675), .B2(n9378), .A(n7197), .ZN(n9678) );
  NAND2_X1 U8906 ( .A1(n9678), .A2(n9665), .ZN(n7207) );
  OAI22_X1 U8907 ( .A1(n9665), .A2(n7199), .B1(n7198), .B2(n9629), .ZN(n7204)
         );
  NAND2_X1 U8908 ( .A1(n7200), .A2(n7205), .ZN(n7201) );
  NAND2_X1 U8909 ( .A1(n7202), .A2(n7201), .ZN(n9677) );
  NOR2_X1 U8910 ( .A1(n9198), .A2(n9677), .ZN(n7203) );
  AOI211_X1 U8911 ( .C1(n9531), .C2(n7205), .A(n7204), .B(n7203), .ZN(n7206)
         );
  OAI211_X1 U8912 ( .C1(n9675), .C2(n7208), .A(n7207), .B(n7206), .ZN(P1_U3289) );
  INV_X1 U8913 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7221) );
  OAI21_X1 U8914 ( .B1(n7211), .B2(n7210), .A(n7209), .ZN(n7219) );
  OAI21_X1 U8915 ( .B1(n7214), .B2(n7213), .A(n7212), .ZN(n7215) );
  NAND2_X1 U8916 ( .A1(n9615), .A2(n7215), .ZN(n7216) );
  NAND2_X1 U8917 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3084), .ZN(n7766) );
  OAI211_X1 U8918 ( .C1(n9617), .C2(n7217), .A(n7216), .B(n7766), .ZN(n7218)
         );
  AOI21_X1 U8919 ( .B1(n9593), .B2(n7219), .A(n7218), .ZN(n7220) );
  OAI21_X1 U8920 ( .B1(n9619), .B2(n7221), .A(n7220), .ZN(P1_U3255) );
  NAND2_X1 U8921 ( .A1(n7223), .A2(n7222), .ZN(n7225) );
  NAND2_X1 U8922 ( .A1(n9752), .A2(n9830), .ZN(n7224) );
  XOR2_X1 U8923 ( .A(n7325), .B(n7324), .Z(n7266) );
  NAND2_X1 U8924 ( .A1(n7105), .A2(n7226), .ZN(n7227) );
  XNOR2_X1 U8925 ( .A(n7227), .B(n7324), .ZN(n7228) );
  AOI222_X1 U8926 ( .A1(n9777), .A2(n7228), .B1(n9748), .B2(n9774), .C1(n8584), 
        .C2(n9772), .ZN(n7265) );
  MUX2_X1 U8927 ( .A(n7229), .B(n7265), .S(n8870), .Z(n7234) );
  INV_X1 U8928 ( .A(n7230), .ZN(n7231) );
  INV_X1 U8929 ( .A(n7333), .ZN(n9783) );
  AOI211_X1 U8930 ( .C1(n7263), .C2(n7231), .A(n9853), .B(n9783), .ZN(n7262)
         );
  NOR2_X1 U8931 ( .A1(n4388), .A2(n4385), .ZN(n8854) );
  OAI22_X1 U8932 ( .A1(n8851), .A2(n9746), .B1(n9778), .B2(n9758), .ZN(n7232)
         );
  AOI21_X1 U8933 ( .B1(n7262), .B2(n8854), .A(n7232), .ZN(n7233) );
  OAI211_X1 U8934 ( .C1(n7266), .C2(n8862), .A(n7234), .B(n7233), .ZN(P2_U3291) );
  NAND2_X1 U8935 ( .A1(n7236), .A2(n7235), .ZN(n7238) );
  AOI22_X1 U8936 ( .A1(n7389), .A2(n7855), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7245), .ZN(n7237) );
  NOR2_X1 U8937 ( .A1(n7238), .A2(n7237), .ZN(n7384) );
  AOI21_X1 U8938 ( .B1(n7238), .B2(n7237), .A(n7384), .ZN(n7250) );
  OAI21_X1 U8939 ( .B1(n7240), .B2(P2_REG1_REG_12__SCAN_IN), .A(n7239), .ZN(
        n7242) );
  AOI22_X1 U8940 ( .A1(n7389), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n5158), .B2(
        n7245), .ZN(n7241) );
  NAND2_X1 U8941 ( .A1(n7241), .A2(n7242), .ZN(n7388) );
  OAI21_X1 U8942 ( .B1(n7242), .B2(n7241), .A(n7388), .ZN(n7248) );
  INV_X1 U8943 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7244) );
  OAI22_X1 U8944 ( .A1(n8655), .A2(n7244), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7243), .ZN(n7247) );
  NOR2_X1 U8945 ( .A1(n9760), .A2(n7245), .ZN(n7246) );
  AOI211_X1 U8946 ( .C1(n9763), .C2(n7248), .A(n7247), .B(n7246), .ZN(n7249)
         );
  OAI21_X1 U8947 ( .B1(n7250), .B2(n8633), .A(n7249), .ZN(P2_U3258) );
  INV_X1 U8948 ( .A(n7251), .ZN(n7313) );
  OAI222_X1 U8949 ( .A1(n8459), .A2(n7253), .B1(n4390), .B2(n7313), .C1(n7252), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  INV_X1 U8950 ( .A(n9790), .ZN(n7254) );
  NAND2_X1 U8951 ( .A1(n7255), .A2(n7254), .ZN(n7260) );
  NAND2_X1 U8952 ( .A1(n7257), .A2(n7256), .ZN(n7258) );
  INV_X1 U8953 ( .A(n7268), .ZN(n7261) );
  INV_X1 U8954 ( .A(n9845), .ZN(n9824) );
  AOI21_X1 U8955 ( .B1(n9818), .B2(n7263), .A(n7262), .ZN(n7264) );
  OAI211_X1 U8956 ( .C1(n9485), .C2(n7266), .A(n7265), .B(n7264), .ZN(n7270)
         );
  NAND2_X1 U8957 ( .A1(n7270), .A2(n9861), .ZN(n7267) );
  OAI21_X1 U8958 ( .B1(n9861), .B2(n5276), .A(n7267), .ZN(P2_U3466) );
  INV_X1 U8959 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7272) );
  NAND2_X1 U8960 ( .A1(n7270), .A2(n9875), .ZN(n7271) );
  OAI21_X1 U8961 ( .B1(n9875), .B2(n7272), .A(n7271), .ZN(P2_U3525) );
  NAND2_X1 U8962 ( .A1(n7315), .A2(n6707), .ZN(n7274) );
  NAND2_X1 U8963 ( .A1(n8113), .A2(n9122), .ZN(n7273) );
  NAND2_X1 U8964 ( .A1(n7274), .A2(n7273), .ZN(n7275) );
  XNOR2_X1 U8965 ( .A(n7275), .B(n8062), .ZN(n7277) );
  NOR2_X1 U8966 ( .A1(n8101), .A2(n9637), .ZN(n7276) );
  AOI21_X1 U8967 ( .B1(n7315), .B2(n8113), .A(n7276), .ZN(n7278) );
  NAND2_X1 U8968 ( .A1(n7277), .A2(n7278), .ZN(n7341) );
  INV_X1 U8969 ( .A(n7277), .ZN(n7280) );
  INV_X1 U8970 ( .A(n7278), .ZN(n7279) );
  NAND2_X1 U8971 ( .A1(n7280), .A2(n7279), .ZN(n7281) );
  NAND2_X1 U8972 ( .A1(n7341), .A2(n7281), .ZN(n7288) );
  INV_X1 U8973 ( .A(n7288), .ZN(n7286) );
  INV_X1 U8974 ( .A(n7342), .ZN(n7287) );
  AOI21_X1 U8975 ( .B1(n7288), .B2(n7285), .A(n7287), .ZN(n7294) );
  OAI22_X1 U8976 ( .A1(n9108), .A2(n7289), .B1(n7434), .B2(n9106), .ZN(n7290)
         );
  AOI211_X1 U8977 ( .C1(n7915), .C2(n9123), .A(n7291), .B(n7290), .ZN(n7293)
         );
  NAND2_X1 U8978 ( .A1(n7315), .A2(n9100), .ZN(n7292) );
  OAI211_X1 U8979 ( .C1(n7294), .C2(n9095), .A(n7293), .B(n7292), .ZN(P1_U3229) );
  INV_X1 U8980 ( .A(n7295), .ZN(n7296) );
  AOI21_X1 U8981 ( .B1(n7297), .B2(n8160), .A(n7296), .ZN(n7298) );
  XOR2_X1 U8982 ( .A(n8261), .B(n7298), .Z(n7299) );
  OAI222_X1 U8983 ( .A1(n9662), .A2(n7671), .B1(n9660), .B2(n9637), .C1(n7299), 
        .C2(n9657), .ZN(n9481) );
  INV_X1 U8984 ( .A(n9481), .ZN(n7310) );
  OAI21_X1 U8985 ( .B1(n7301), .B2(n6121), .A(n7300), .ZN(n9483) );
  INV_X1 U8986 ( .A(n9374), .ZN(n9540) );
  NAND2_X1 U8987 ( .A1(n7302), .A2(n9479), .ZN(n7303) );
  NAND2_X1 U8988 ( .A1(n7303), .A2(n9690), .ZN(n7304) );
  OR2_X1 U8989 ( .A1(n7366), .A2(n7304), .ZN(n9480) );
  OAI22_X1 U8990 ( .A1(n9665), .A2(n7305), .B1(n7353), .B2(n9629), .ZN(n7306)
         );
  AOI21_X1 U8991 ( .B1(n9479), .B2(n9531), .A(n7306), .ZN(n7307) );
  OAI21_X1 U8992 ( .B1(n9480), .B2(n9516), .A(n7307), .ZN(n7308) );
  AOI21_X1 U8993 ( .B1(n9483), .B2(n9540), .A(n7308), .ZN(n7309) );
  OAI21_X1 U8994 ( .B1(n7310), .B2(n4389), .A(n7309), .ZN(P1_U3281) );
  OAI222_X1 U8995 ( .A1(n8419), .A2(n7313), .B1(P1_U3084), .B2(n7312), .C1(
        n7311), .C2(n8421), .ZN(P1_U3332) );
  NAND2_X1 U8996 ( .A1(n6149), .A2(n4486), .ZN(n8232) );
  OR2_X1 U8997 ( .A1(n8232), .A2(n6147), .ZN(n9694) );
  INV_X1 U8998 ( .A(n7314), .ZN(n7319) );
  AOI22_X1 U8999 ( .A1(n7316), .A2(n9690), .B1(n9689), .B2(n7315), .ZN(n7317)
         );
  OAI211_X1 U9000 ( .C1(n9694), .C2(n7319), .A(n7318), .B(n7317), .ZN(n7321)
         );
  NAND2_X1 U9001 ( .A1(n7321), .A2(n9742), .ZN(n7320) );
  OAI21_X1 U9002 ( .B1(n9742), .B2(n6427), .A(n7320), .ZN(P1_U3532) );
  INV_X1 U9003 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7323) );
  NAND2_X1 U9004 ( .A1(n7321), .A2(n9726), .ZN(n7322) );
  OAI21_X1 U9005 ( .B1(n9726), .B2(n7323), .A(n7322), .ZN(P1_U3481) );
  INV_X1 U9006 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7338) );
  NOR2_X1 U9007 ( .A1(n9748), .A2(n7332), .ZN(n7327) );
  NAND2_X1 U9008 ( .A1(n9748), .A2(n7332), .ZN(n7326) );
  XOR2_X1 U9009 ( .A(n7486), .B(n7487), .Z(n7405) );
  XOR2_X1 U9010 ( .A(n7328), .B(n7487), .Z(n7331) );
  NAND2_X1 U9011 ( .A1(n9748), .A2(n9772), .ZN(n7329) );
  OAI21_X1 U9012 ( .B1(n7330), .B2(n8882), .A(n7329), .ZN(n7440) );
  AOI21_X1 U9013 ( .B1(n7331), .B2(n9777), .A(n7440), .ZN(n7400) );
  AND2_X1 U9014 ( .A1(n4963), .A2(n7335), .ZN(n7334) );
  NOR2_X1 U9015 ( .A1(n7523), .A2(n7334), .ZN(n7403) );
  AOI22_X1 U9016 ( .A1(n7403), .A2(n9819), .B1(n9818), .B2(n7335), .ZN(n7336)
         );
  OAI211_X1 U9017 ( .C1(n7405), .C2(n9485), .A(n7400), .B(n7336), .ZN(n7339)
         );
  NAND2_X1 U9018 ( .A1(n7339), .A2(n9875), .ZN(n7337) );
  OAI21_X1 U9019 ( .B1(n9875), .B2(n7338), .A(n7337), .ZN(P2_U3527) );
  NAND2_X1 U9020 ( .A1(n7339), .A2(n9861), .ZN(n7340) );
  OAI21_X1 U9021 ( .B1(n9861), .B2(n5313), .A(n7340), .ZN(P2_U3472) );
  NAND2_X1 U9022 ( .A1(n7342), .A2(n7341), .ZN(n7424) );
  NAND2_X1 U9023 ( .A1(n9479), .A2(n6707), .ZN(n7344) );
  NAND2_X1 U9024 ( .A1(n8113), .A2(n9121), .ZN(n7343) );
  NAND2_X1 U9025 ( .A1(n7344), .A2(n7343), .ZN(n7345) );
  XNOR2_X1 U9026 ( .A(n7345), .B(n6738), .ZN(n7348) );
  NAND2_X1 U9027 ( .A1(n9479), .A2(n8113), .ZN(n7347) );
  NAND2_X1 U9028 ( .A1(n6764), .A2(n9121), .ZN(n7346) );
  NAND2_X1 U9029 ( .A1(n7347), .A2(n7346), .ZN(n7349) );
  NAND2_X1 U9030 ( .A1(n7348), .A2(n7349), .ZN(n7423) );
  INV_X1 U9031 ( .A(n7348), .ZN(n7351) );
  INV_X1 U9032 ( .A(n7349), .ZN(n7350) );
  NAND2_X1 U9033 ( .A1(n7351), .A2(n7350), .ZN(n7425) );
  NAND2_X1 U9034 ( .A1(n7423), .A2(n7425), .ZN(n7352) );
  XNOR2_X1 U9035 ( .A(n7424), .B(n7352), .ZN(n7358) );
  OAI22_X1 U9036 ( .A1(n9108), .A2(n7353), .B1(n9637), .B2(n9110), .ZN(n7354)
         );
  AOI211_X1 U9037 ( .C1(n9088), .C2(n9527), .A(n7355), .B(n7354), .ZN(n7357)
         );
  NAND2_X1 U9038 ( .A1(n9479), .A2(n9100), .ZN(n7356) );
  OAI211_X1 U9039 ( .C1(n7358), .C2(n9095), .A(n7357), .B(n7356), .ZN(P1_U3215) );
  NAND2_X1 U9040 ( .A1(n7360), .A2(n7359), .ZN(n8264) );
  XOR2_X1 U9041 ( .A(n7361), .B(n8264), .Z(n7365) );
  OAI22_X1 U9042 ( .A1(n7434), .A2(n9660), .B1(n9662), .B2(n7658), .ZN(n7364)
         );
  XNOR2_X1 U9043 ( .A(n7362), .B(n8264), .ZN(n7466) );
  NOR2_X1 U9044 ( .A1(n7466), .A2(n9378), .ZN(n7363) );
  AOI211_X1 U9045 ( .C1(n9635), .C2(n7365), .A(n7364), .B(n7363), .ZN(n7465)
         );
  INV_X1 U9046 ( .A(n7466), .ZN(n7372) );
  NOR2_X1 U9047 ( .A1(n7366), .A2(n7461), .ZN(n7367) );
  OR2_X1 U9048 ( .A1(n9537), .A2(n7367), .ZN(n7462) );
  OAI22_X1 U9049 ( .A1(n9665), .A2(n7368), .B1(n7435), .B2(n9629), .ZN(n7369)
         );
  AOI21_X1 U9050 ( .B1(n7430), .B2(n9531), .A(n7369), .ZN(n7370) );
  OAI21_X1 U9051 ( .B1(n7462), .B2(n9198), .A(n7370), .ZN(n7371) );
  AOI21_X1 U9052 ( .B1(n7372), .B2(n7737), .A(n7371), .ZN(n7373) );
  OAI21_X1 U9053 ( .B1(n7465), .B2(n4389), .A(n7373), .ZN(P1_U3280) );
  INV_X1 U9054 ( .A(n7374), .ZN(n7375) );
  AOI21_X1 U9055 ( .B1(n7442), .B2(n7375), .A(n9743), .ZN(n7379) );
  NOR3_X1 U9056 ( .A1(n8552), .A2(n7376), .A3(n8129), .ZN(n7378) );
  OAI21_X1 U9057 ( .B1(n7379), .B2(n7378), .A(n7377), .ZN(n7383) );
  OAI22_X1 U9058 ( .A1(n9751), .A2(n8129), .B1(n9759), .B2(n7521), .ZN(n7380)
         );
  AOI211_X1 U9059 ( .C1(n8465), .C2(n8582), .A(n7381), .B(n7380), .ZN(n7382)
         );
  OAI211_X1 U9060 ( .C1(n9840), .C2(n9747), .A(n7383), .B(n7382), .ZN(P2_U3223) );
  NOR2_X1 U9061 ( .A1(n7389), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7385) );
  NOR2_X1 U9062 ( .A1(n7385), .A2(n7384), .ZN(n7387) );
  AOI22_X1 U9063 ( .A1(n7743), .A2(n8869), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7740), .ZN(n7386) );
  NOR2_X1 U9064 ( .A1(n7387), .A2(n7386), .ZN(n7739) );
  AOI21_X1 U9065 ( .B1(n7387), .B2(n7386), .A(n7739), .ZN(n7397) );
  AOI22_X1 U9066 ( .A1(n7743), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n5141), .B2(
        n7740), .ZN(n7391) );
  OAI21_X1 U9067 ( .B1(n7389), .B2(P2_REG1_REG_13__SCAN_IN), .A(n7388), .ZN(
        n7390) );
  NAND2_X1 U9068 ( .A1(n7391), .A2(n7390), .ZN(n7742) );
  OAI21_X1 U9069 ( .B1(n7391), .B2(n7390), .A(n7742), .ZN(n7392) );
  NAND2_X1 U9070 ( .A1(n7392), .A2(n9763), .ZN(n7396) );
  INV_X1 U9071 ( .A(n9760), .ZN(n9472) );
  INV_X1 U9072 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7393) );
  NAND2_X1 U9073 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7944) );
  OAI21_X1 U9074 ( .B1(n8655), .B2(n7393), .A(n7944), .ZN(n7394) );
  AOI21_X1 U9075 ( .B1(n9472), .B2(n7743), .A(n7394), .ZN(n7395) );
  OAI211_X1 U9076 ( .C1(n7397), .C2(n8633), .A(n7396), .B(n7395), .ZN(P2_U3259) );
  INV_X1 U9077 ( .A(n7398), .ZN(n7448) );
  AOI22_X1 U9078 ( .A1(n4388), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n7448), .B2(
        n8848), .ZN(n7399) );
  OAI21_X1 U9079 ( .B1(n7490), .B2(n8851), .A(n7399), .ZN(n7402) );
  NOR2_X1 U9080 ( .A1(n7400), .A2(n4388), .ZN(n7401) );
  AOI211_X1 U9081 ( .C1(n7403), .C2(n8834), .A(n7402), .B(n7401), .ZN(n7404)
         );
  OAI21_X1 U9082 ( .B1(n8862), .B2(n7405), .A(n7404), .ZN(P2_U3289) );
  INV_X1 U9083 ( .A(n7406), .ZN(n8418) );
  OAI222_X1 U9084 ( .A1(n8459), .A2(n7408), .B1(n4390), .B2(n8418), .C1(
        P2_U3152), .C2(n7407), .ZN(P2_U3336) );
  OR2_X1 U9085 ( .A1(n7409), .A2(n9535), .ZN(n9533) );
  NAND2_X1 U9086 ( .A1(n9533), .A2(n7410), .ZN(n7412) );
  XNOR2_X1 U9087 ( .A(n7412), .B(n7411), .ZN(n7566) );
  XNOR2_X1 U9088 ( .A(n7413), .B(n8266), .ZN(n7415) );
  AOI22_X1 U9089 ( .A1(n9526), .A2(n9120), .B1(n9524), .B2(n9119), .ZN(n7414)
         );
  OAI21_X1 U9090 ( .B1(n7415), .B2(n9657), .A(n7414), .ZN(n7416) );
  AOI21_X1 U9091 ( .B1(n7566), .B2(n7731), .A(n7416), .ZN(n7569) );
  INV_X1 U9092 ( .A(n7417), .ZN(n7478) );
  AOI21_X1 U9093 ( .B1(n7706), .B2(n9536), .A(n7478), .ZN(n7567) );
  NOR2_X1 U9094 ( .A1(n4689), .A2(n9370), .ZN(n7420) );
  OAI22_X1 U9095 ( .A1(n9665), .A2(n7418), .B1(n7703), .B2(n9629), .ZN(n7419)
         );
  AOI211_X1 U9096 ( .C1(n7567), .C2(n9337), .A(n7420), .B(n7419), .ZN(n7422)
         );
  NAND2_X1 U9097 ( .A1(n7566), .A2(n7737), .ZN(n7421) );
  OAI211_X1 U9098 ( .C1(n7569), .C2(n4389), .A(n7422), .B(n7421), .ZN(P1_U3278) );
  NAND2_X1 U9099 ( .A1(n7430), .A2(n6707), .ZN(n7427) );
  NAND2_X1 U9100 ( .A1(n8113), .A2(n9527), .ZN(n7426) );
  NAND2_X1 U9101 ( .A1(n7427), .A2(n7426), .ZN(n7428) );
  XNOR2_X1 U9102 ( .A(n7428), .B(n8062), .ZN(n7660) );
  NOR2_X1 U9103 ( .A1(n8101), .A2(n7671), .ZN(n7429) );
  AOI21_X1 U9104 ( .B1(n7430), .B2(n8113), .A(n7429), .ZN(n7661) );
  XNOR2_X1 U9105 ( .A(n7660), .B(n7661), .ZN(n7432) );
  AOI21_X1 U9106 ( .B1(n7431), .B2(n7432), .A(n9095), .ZN(n7433) );
  NAND2_X1 U9107 ( .A1(n7433), .A2(n7665), .ZN(n7439) );
  OAI22_X1 U9108 ( .A1(n9108), .A2(n7435), .B1(n7434), .B2(n9110), .ZN(n7436)
         );
  AOI211_X1 U9109 ( .C1(n9088), .C2(n9120), .A(n7437), .B(n7436), .ZN(n7438)
         );
  OAI211_X1 U9110 ( .C1(n7461), .C2(n9115), .A(n7439), .B(n7438), .ZN(P1_U3234) );
  AOI22_X1 U9111 ( .A1(n7440), .A2(n8523), .B1(P2_REG3_REG_7__SCAN_IN), .B2(
        P2_U3152), .ZN(n7441) );
  OAI21_X1 U9112 ( .B1(n7490), .B2(n9747), .A(n7441), .ZN(n7447) );
  INV_X1 U9113 ( .A(n7442), .ZN(n7443) );
  AOI211_X1 U9114 ( .C1(n7445), .C2(n7444), .A(n9743), .B(n7443), .ZN(n7446)
         );
  AOI211_X1 U9115 ( .C1(n8511), .C2(n7448), .A(n7447), .B(n7446), .ZN(n7449)
         );
  INV_X1 U9116 ( .A(n7449), .ZN(P2_U3215) );
  NAND2_X1 U9117 ( .A1(n7454), .A2(n7450), .ZN(n7452) );
  OAI211_X1 U9118 ( .C1(n7453), .C2(n8459), .A(n7452), .B(n7451), .ZN(P2_U3335) );
  NAND2_X1 U9119 ( .A1(n7454), .A2(n7710), .ZN(n7456) );
  NAND2_X1 U9120 ( .A1(n7455), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8417) );
  OAI211_X1 U9121 ( .C1(n7457), .C2(n8421), .A(n7456), .B(n8417), .ZN(P1_U3330) );
  INV_X1 U9122 ( .A(n7458), .ZN(n7484) );
  OAI222_X1 U9123 ( .A1(n8419), .A2(n7484), .B1(P1_U3084), .B2(n7460), .C1(
        n7459), .C2(n8421), .ZN(P1_U3329) );
  INV_X1 U9124 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7468) );
  OAI22_X1 U9125 ( .A1(n7462), .A2(n9705), .B1(n7461), .B2(n9718), .ZN(n7463)
         );
  INV_X1 U9126 ( .A(n7463), .ZN(n7464) );
  OAI211_X1 U9127 ( .C1(n9694), .C2(n7466), .A(n7465), .B(n7464), .ZN(n7469)
         );
  NAND2_X1 U9128 ( .A1(n7469), .A2(n9726), .ZN(n7467) );
  OAI21_X1 U9129 ( .B1(n9726), .B2(n7468), .A(n7467), .ZN(P1_U3487) );
  NAND2_X1 U9130 ( .A1(n7469), .A2(n9742), .ZN(n7470) );
  OAI21_X1 U9131 ( .B1(n9742), .B2(n6428), .A(n7470), .ZN(P1_U3534) );
  AOI21_X1 U9132 ( .B1(n7471), .B2(n8267), .A(n9657), .ZN(n7474) );
  OAI22_X1 U9133 ( .A1(n7700), .A2(n9660), .B1(n9662), .B2(n7975), .ZN(n7472)
         );
  AOI21_X1 U9134 ( .B1(n7474), .B2(n7473), .A(n7472), .ZN(n9557) );
  XOR2_X1 U9135 ( .A(n8267), .B(n7475), .Z(n9560) );
  NAND2_X1 U9136 ( .A1(n9560), .A2(n9540), .ZN(n7482) );
  INV_X1 U9137 ( .A(n7765), .ZN(n7476) );
  OAI22_X1 U9138 ( .A1(n9665), .A2(n7213), .B1(n7476), .B2(n9629), .ZN(n7480)
         );
  INV_X1 U9139 ( .A(n7769), .ZN(n9558) );
  INV_X1 U9140 ( .A(n7732), .ZN(n7477) );
  OAI211_X1 U9141 ( .C1(n9558), .C2(n7478), .A(n7477), .B(n9690), .ZN(n9556)
         );
  NOR2_X1 U9142 ( .A1(n9556), .A2(n9516), .ZN(n7479) );
  AOI211_X1 U9143 ( .C1(n9531), .C2(n7769), .A(n7480), .B(n7479), .ZN(n7481)
         );
  OAI211_X1 U9144 ( .C1(n4389), .C2(n9557), .A(n7482), .B(n7481), .ZN(P1_U3277) );
  OAI222_X1 U9145 ( .A1(P2_U3152), .A2(n7485), .B1(n4390), .B2(n7484), .C1(
        n7483), .C2(n8459), .ZN(P2_U3334) );
  INV_X1 U9146 ( .A(n7486), .ZN(n7489) );
  NAND2_X1 U9147 ( .A1(n7489), .A2(n7488), .ZN(n7782) );
  NAND2_X1 U9148 ( .A1(n8129), .A2(n7490), .ZN(n7583) );
  NAND2_X1 U9149 ( .A1(n7782), .A2(n7583), .ZN(n7576) );
  NAND2_X1 U9150 ( .A1(n8583), .A2(n7528), .ZN(n7491) );
  AND2_X1 U9151 ( .A1(n7514), .A2(n7491), .ZN(n7494) );
  AND2_X1 U9152 ( .A1(n7492), .A2(n7491), .ZN(n7577) );
  NAND2_X1 U9153 ( .A1(n7514), .A2(n7577), .ZN(n7493) );
  OAI21_X1 U9154 ( .B1(n7494), .B2(n7492), .A(n7493), .ZN(n7717) );
  INV_X1 U9155 ( .A(n7842), .ZN(n9827) );
  NAND3_X1 U9156 ( .A1(n7495), .A2(n7492), .A3(n7496), .ZN(n7497) );
  NAND2_X1 U9157 ( .A1(n7498), .A2(n7497), .ZN(n7499) );
  NAND2_X1 U9158 ( .A1(n7499), .A2(n9777), .ZN(n7502) );
  INV_X1 U9159 ( .A(n7687), .ZN(n8581) );
  NAND2_X1 U9160 ( .A1(n8581), .A2(n9774), .ZN(n7501) );
  NAND2_X1 U9161 ( .A1(n8583), .A2(n9772), .ZN(n7500) );
  AND2_X1 U9162 ( .A1(n7501), .A2(n7500), .ZN(n7551) );
  NAND2_X1 U9163 ( .A1(n7502), .A2(n7551), .ZN(n7503) );
  AOI21_X1 U9164 ( .B1(n7717), .B2(n9827), .A(n7503), .ZN(n7719) );
  INV_X1 U9165 ( .A(n7504), .ZN(n7505) );
  NAND2_X1 U9166 ( .A1(n8870), .A2(n7505), .ZN(n7861) );
  INV_X1 U9167 ( .A(n7861), .ZN(n7511) );
  OR2_X1 U9168 ( .A1(n7525), .A2(n7714), .ZN(n7506) );
  NAND2_X1 U9169 ( .A1(n7596), .A2(n7506), .ZN(n7715) );
  OAI22_X1 U9170 ( .A1(n8870), .A2(n7507), .B1(n7549), .B2(n9778), .ZN(n7508)
         );
  AOI21_X1 U9171 ( .B1(n8872), .B2(n6163), .A(n7508), .ZN(n7509) );
  OAI21_X1 U9172 ( .B1(n7715), .B2(n8874), .A(n7509), .ZN(n7510) );
  AOI21_X1 U9173 ( .B1(n7717), .B2(n7511), .A(n7510), .ZN(n7512) );
  OAI21_X1 U9174 ( .B1(n7719), .B2(n4388), .A(n7512), .ZN(P2_U3287) );
  NAND2_X1 U9175 ( .A1(n7576), .A2(n7575), .ZN(n7513) );
  INV_X1 U9176 ( .A(n9844), .ZN(n7531) );
  INV_X1 U9177 ( .A(n7495), .ZN(n7515) );
  AOI21_X1 U9178 ( .B1(n7517), .B2(n7516), .A(n7515), .ZN(n7520) );
  INV_X1 U9179 ( .A(n9777), .ZN(n8877) );
  AOI22_X1 U9180 ( .A1(n9772), .A2(n9775), .B1(n8582), .B2(n9774), .ZN(n7519)
         );
  NAND2_X1 U9181 ( .A1(n9844), .A2(n9827), .ZN(n7518) );
  OAI211_X1 U9182 ( .C1(n7520), .C2(n8877), .A(n7519), .B(n7518), .ZN(n9842)
         );
  NAND2_X1 U9183 ( .A1(n9842), .A2(n8870), .ZN(n7530) );
  OAI22_X1 U9184 ( .A1(n8870), .A2(n7522), .B1(n7521), .B2(n9778), .ZN(n7527)
         );
  NOR2_X1 U9185 ( .A1(n7523), .A2(n9840), .ZN(n7524) );
  OR2_X1 U9186 ( .A1(n7525), .A2(n7524), .ZN(n9841) );
  NOR2_X1 U9187 ( .A1(n9841), .A2(n8874), .ZN(n7526) );
  AOI211_X1 U9188 ( .C1(n8872), .C2(n7528), .A(n7527), .B(n7526), .ZN(n7529)
         );
  OAI211_X1 U9189 ( .C1(n7531), .C2(n7861), .A(n7530), .B(n7529), .ZN(P2_U3288) );
  INV_X1 U9190 ( .A(n7532), .ZN(n7564) );
  OAI222_X1 U9191 ( .A1(n8419), .A2(n7564), .B1(P1_U3084), .B2(n7534), .C1(
        n7533), .C2(n8421), .ZN(P1_U3327) );
  INV_X1 U9192 ( .A(n7535), .ZN(n7539) );
  OAI222_X1 U9193 ( .A1(n8459), .A2(n7537), .B1(n4390), .B2(n7539), .C1(
        P2_U3152), .C2(n7536), .ZN(P2_U3333) );
  OAI222_X1 U9194 ( .A1(n8421), .A2(n9958), .B1(n8419), .B2(n7539), .C1(n7538), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  INV_X1 U9195 ( .A(n7544), .ZN(n7541) );
  NOR3_X1 U9196 ( .A1(n7541), .A2(n7540), .A3(n9743), .ZN(n7547) );
  NAND3_X1 U9197 ( .A1(n8533), .A2(n7542), .A3(n8582), .ZN(n7543) );
  OAI21_X1 U9198 ( .B1(n7544), .B2(n9743), .A(n7543), .ZN(n7546) );
  MUX2_X1 U9199 ( .A(n7547), .B(n7546), .S(n7545), .Z(n7548) );
  INV_X1 U9200 ( .A(n7548), .ZN(n7555) );
  INV_X1 U9201 ( .A(n7549), .ZN(n7553) );
  OAI22_X1 U9202 ( .A1(n7551), .A2(n8508), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7550), .ZN(n7552) );
  AOI21_X1 U9203 ( .B1(n7553), .B2(n8511), .A(n7552), .ZN(n7554) );
  OAI211_X1 U9204 ( .C1(n7714), .C2(n9747), .A(n7555), .B(n7554), .ZN(P2_U3233) );
  XNOR2_X1 U9205 ( .A(n7557), .B(n7556), .ZN(n7562) );
  OAI21_X1 U9206 ( .B1(n9750), .B2(n7788), .A(n7558), .ZN(n7560) );
  OAI22_X1 U9207 ( .A1(n9751), .A2(n7593), .B1(n7594), .B2(n9759), .ZN(n7559)
         );
  AOI211_X1 U9208 ( .C1(n8565), .C2(n7779), .A(n7560), .B(n7559), .ZN(n7561)
         );
  OAI21_X1 U9209 ( .B1(n7562), .B2(n9743), .A(n7561), .ZN(P2_U3219) );
  OAI222_X1 U9210 ( .A1(P2_U3152), .A2(n7565), .B1(n4390), .B2(n7564), .C1(
        n7563), .C2(n8459), .ZN(P2_U3332) );
  INV_X1 U9211 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7572) );
  INV_X1 U9212 ( .A(n7566), .ZN(n7570) );
  AOI22_X1 U9213 ( .A1(n7567), .A2(n9690), .B1(n9689), .B2(n7706), .ZN(n7568)
         );
  OAI211_X1 U9214 ( .C1(n9694), .C2(n7570), .A(n7569), .B(n7568), .ZN(n7573)
         );
  NAND2_X1 U9215 ( .A1(n7573), .A2(n9726), .ZN(n7571) );
  OAI21_X1 U9216 ( .B1(n9726), .B2(n7572), .A(n7571), .ZN(P1_U3493) );
  NAND2_X1 U9217 ( .A1(n7573), .A2(n9742), .ZN(n7574) );
  OAI21_X1 U9218 ( .B1(n9742), .B2(n6413), .A(n7574), .ZN(P1_U3536) );
  AND2_X1 U9219 ( .A1(n7593), .A2(n7714), .ZN(n7578) );
  OR2_X1 U9220 ( .A1(n7575), .A2(n7578), .ZN(n7582) );
  OR2_X1 U9221 ( .A1(n7576), .A2(n7582), .ZN(n7581) );
  INV_X1 U9222 ( .A(n7577), .ZN(n7580) );
  NAND2_X1 U9223 ( .A1(n7581), .A2(n7586), .ZN(n7589) );
  INV_X1 U9224 ( .A(n7590), .ZN(n7585) );
  NOR2_X1 U9225 ( .A1(n7582), .A2(n7585), .ZN(n7584) );
  NAND2_X1 U9226 ( .A1(n7782), .A2(n7778), .ZN(n7865) );
  INV_X1 U9227 ( .A(n7865), .ZN(n7587) );
  NOR2_X1 U9228 ( .A1(n7587), .A2(n7780), .ZN(n7588) );
  OAI21_X1 U9229 ( .B1(n7589), .B2(n7590), .A(n7588), .ZN(n9846) );
  XNOR2_X1 U9230 ( .A(n7591), .B(n7590), .ZN(n7592) );
  OAI222_X1 U9231 ( .A1(n8882), .A2(n7788), .B1(n8880), .B2(n7593), .C1(n7592), 
        .C2(n8877), .ZN(n9848) );
  NAND2_X1 U9232 ( .A1(n9848), .A2(n8870), .ZN(n7601) );
  OAI22_X1 U9233 ( .A1(n8870), .A2(n7595), .B1(n7594), .B2(n9778), .ZN(n7599)
         );
  INV_X1 U9234 ( .A(n7596), .ZN(n7597) );
  OAI21_X1 U9235 ( .B1(n7597), .B2(n4702), .A(n7868), .ZN(n9847) );
  NOR2_X1 U9236 ( .A1(n9847), .A2(n8874), .ZN(n7598) );
  AOI211_X1 U9237 ( .C1(n8872), .C2(n7779), .A(n7599), .B(n7598), .ZN(n7600)
         );
  OAI211_X1 U9238 ( .C1(n9846), .C2(n8862), .A(n7601), .B(n7600), .ZN(P2_U3286) );
  NAND2_X1 U9239 ( .A1(n7676), .A2(n7710), .ZN(n7602) );
  OAI211_X1 U9240 ( .C1(n8421), .C2(n7603), .A(n7602), .B(n9180), .ZN(P1_U3326) );
  NOR2_X1 U9241 ( .A1(n7611), .A2(n7604), .ZN(n7606) );
  NAND2_X1 U9242 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n7805), .ZN(n7607) );
  OAI21_X1 U9243 ( .B1(n7805), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7607), .ZN(
        n7608) );
  AOI211_X1 U9244 ( .C1(n7609), .C2(n7608), .A(n7804), .B(n9598), .ZN(n7621)
         );
  NOR2_X1 U9245 ( .A1(n7611), .A2(n7610), .ZN(n7613) );
  NOR2_X1 U9246 ( .A1(n7613), .A2(n7612), .ZN(n7616) );
  INV_X1 U9247 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9555) );
  NOR2_X1 U9248 ( .A1(n7805), .A2(n9555), .ZN(n7614) );
  AOI21_X1 U9249 ( .B1(n7805), .B2(n9555), .A(n7614), .ZN(n7615) );
  NOR2_X1 U9250 ( .A1(n7616), .A2(n7615), .ZN(n7801) );
  AOI211_X1 U9251 ( .C1(n7616), .C2(n7615), .A(n7801), .B(n9608), .ZN(n7620)
         );
  INV_X1 U9252 ( .A(n9619), .ZN(n9146) );
  NAND2_X1 U9253 ( .A1(n9146), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7617) );
  NAND2_X1 U9254 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7974) );
  OAI211_X1 U9255 ( .C1(n7618), .C2(n9617), .A(n7617), .B(n7974), .ZN(n7619)
         );
  OR3_X1 U9256 ( .A1(n7621), .A2(n7620), .A3(n7619), .ZN(P1_U3257) );
  INV_X1 U9257 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10201) );
  NOR2_X1 U9258 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7622) );
  AOI21_X1 U9259 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7622), .ZN(n9882) );
  NOR2_X1 U9260 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7623) );
  AOI21_X1 U9261 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7623), .ZN(n9885) );
  NAND2_X1 U9262 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), 
        .ZN(n7624) );
  OAI21_X1 U9263 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7624), .ZN(n9894) );
  NOR2_X1 U9264 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7631) );
  XNOR2_X1 U9265 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10212) );
  NAND2_X1 U9266 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7629) );
  NOR2_X1 U9267 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n10124) );
  AOI21_X1 U9268 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10124), .ZN(n10210) );
  NAND2_X1 U9269 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7627) );
  XOR2_X1 U9270 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10208) );
  AOI21_X1 U9271 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9876) );
  INV_X1 U9272 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7625) );
  NAND3_X1 U9273 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9878) );
  OAI21_X1 U9274 ( .B1(n9876), .B2(n7625), .A(n9878), .ZN(n10207) );
  NAND2_X1 U9275 ( .A1(n10208), .A2(n10207), .ZN(n7626) );
  NAND2_X1 U9276 ( .A1(n7627), .A2(n7626), .ZN(n10209) );
  NAND2_X1 U9277 ( .A1(n10210), .A2(n10209), .ZN(n7628) );
  NAND2_X1 U9278 ( .A1(n7629), .A2(n7628), .ZN(n10211) );
  NOR2_X1 U9279 ( .A1(n10212), .A2(n10211), .ZN(n7630) );
  NOR2_X1 U9280 ( .A1(n7631), .A2(n7630), .ZN(n7632) );
  NOR2_X1 U9281 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7632), .ZN(n10197) );
  AND2_X1 U9282 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7632), .ZN(n10196) );
  NOR2_X1 U9283 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10196), .ZN(n7633) );
  NOR2_X1 U9284 ( .A1(n10197), .A2(n7633), .ZN(n7634) );
  NAND2_X1 U9285 ( .A1(n7634), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7636) );
  XOR2_X1 U9286 ( .A(n7634), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10195) );
  NAND2_X1 U9287 ( .A1(n10195), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7635) );
  NAND2_X1 U9288 ( .A1(n7636), .A2(n7635), .ZN(n7637) );
  NAND2_X1 U9289 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n7637), .ZN(n7639) );
  XOR2_X1 U9290 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n7637), .Z(n10194) );
  NAND2_X1 U9291 ( .A1(n10194), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n7638) );
  NAND2_X1 U9292 ( .A1(n7639), .A2(n7638), .ZN(n7640) );
  NAND2_X1 U9293 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n7640), .ZN(n7642) );
  XOR2_X1 U9294 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n7640), .Z(n10206) );
  NAND2_X1 U9295 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n10206), .ZN(n7641) );
  NAND2_X1 U9296 ( .A1(n7642), .A2(n7641), .ZN(n7643) );
  AND2_X1 U9297 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7643), .ZN(n7644) );
  XNOR2_X1 U9298 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7643), .ZN(n10204) );
  NOR2_X1 U9299 ( .A1(n10205), .A2(n10204), .ZN(n10203) );
  NAND2_X1 U9300 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7645) );
  OAI21_X1 U9301 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7645), .ZN(n9902) );
  AOI21_X1 U9302 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9901), .ZN(n9900) );
  NAND2_X1 U9303 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7646) );
  OAI21_X1 U9304 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7646), .ZN(n9899) );
  NOR2_X1 U9305 ( .A1(n9900), .A2(n9899), .ZN(n9898) );
  AOI21_X1 U9306 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9898), .ZN(n9897) );
  NOR2_X1 U9307 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7647) );
  AOI21_X1 U9308 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7647), .ZN(n9896) );
  NAND2_X1 U9309 ( .A1(n9897), .A2(n9896), .ZN(n9895) );
  OAI21_X1 U9310 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9895), .ZN(n9893) );
  NOR2_X1 U9311 ( .A1(n9894), .A2(n9893), .ZN(n9892) );
  AOI21_X1 U9312 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9892), .ZN(n9891) );
  NAND2_X1 U9313 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(P2_ADDR_REG_14__SCAN_IN), 
        .ZN(n7648) );
  OAI21_X1 U9314 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7648), .ZN(n9890) );
  NOR2_X1 U9315 ( .A1(n9891), .A2(n9890), .ZN(n9889) );
  AOI21_X1 U9316 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9889), .ZN(n9888) );
  NOR2_X1 U9317 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7649) );
  AOI21_X1 U9318 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7649), .ZN(n9887) );
  NAND2_X1 U9319 ( .A1(n9888), .A2(n9887), .ZN(n9886) );
  OAI21_X1 U9320 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9886), .ZN(n9884) );
  NAND2_X1 U9321 ( .A1(n9885), .A2(n9884), .ZN(n9883) );
  OAI21_X1 U9322 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9883), .ZN(n9881) );
  NAND2_X1 U9323 ( .A1(n9882), .A2(n9881), .ZN(n9880) );
  OAI21_X1 U9324 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9880), .ZN(n10200) );
  NOR2_X1 U9325 ( .A1(n10201), .A2(n10200), .ZN(n7650) );
  NAND2_X1 U9326 ( .A1(n10201), .A2(n10200), .ZN(n10199) );
  OAI21_X1 U9327 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7650), .A(n10199), .ZN(
        n7654) );
  NOR2_X1 U9328 ( .A1(n7652), .A2(n7651), .ZN(n7653) );
  XNOR2_X1 U9329 ( .A(n7654), .B(n7653), .ZN(ADD_1071_U4) );
  NAND2_X1 U9330 ( .A1(n9532), .A2(n6707), .ZN(n7656) );
  NAND2_X1 U9331 ( .A1(n8113), .A2(n9120), .ZN(n7655) );
  NAND2_X1 U9332 ( .A1(n7656), .A2(n7655), .ZN(n7657) );
  XNOR2_X1 U9333 ( .A(n7657), .B(n8062), .ZN(n7694) );
  NOR2_X1 U9334 ( .A1(n8101), .A2(n7658), .ZN(n7659) );
  AOI21_X1 U9335 ( .B1(n9532), .B2(n8113), .A(n7659), .ZN(n7693) );
  XNOR2_X1 U9336 ( .A(n7694), .B(n7693), .ZN(n7669) );
  INV_X1 U9337 ( .A(n7660), .ZN(n7663) );
  INV_X1 U9338 ( .A(n7661), .ZN(n7662) );
  NAND2_X1 U9339 ( .A1(n7663), .A2(n7662), .ZN(n7664) );
  INV_X1 U9340 ( .A(n7669), .ZN(n7666) );
  INV_X1 U9341 ( .A(n7696), .ZN(n7667) );
  AOI21_X1 U9342 ( .B1(n7669), .B2(n7668), .A(n7667), .ZN(n7675) );
  OAI21_X1 U9343 ( .B1(n9106), .B2(n7700), .A(n7670), .ZN(n7673) );
  OAI22_X1 U9344 ( .A1(n9108), .A2(n9529), .B1(n7671), .B2(n9110), .ZN(n7672)
         );
  AOI211_X1 U9345 ( .C1(n9532), .C2(n9100), .A(n7673), .B(n7672), .ZN(n7674)
         );
  OAI21_X1 U9346 ( .B1(n7675), .B2(n9095), .A(n7674), .ZN(P1_U3222) );
  INV_X1 U9347 ( .A(n7676), .ZN(n7678) );
  OAI222_X1 U9348 ( .A1(n8459), .A2(n7679), .B1(n4390), .B2(n7678), .C1(n7677), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  NOR3_X1 U9349 ( .A1(n7680), .A2(n7788), .A3(n8552), .ZN(n7681) );
  AOI21_X1 U9350 ( .B1(n7682), .B2(n8544), .A(n7681), .ZN(n7692) );
  AOI21_X1 U9351 ( .B1(n7685), .B2(n7684), .A(n7683), .ZN(n7691) );
  OAI22_X1 U9352 ( .A1(n9750), .A2(n7849), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7686), .ZN(n7689) );
  OAI22_X1 U9353 ( .A1(n9751), .A2(n7687), .B1(n7869), .B2(n9759), .ZN(n7688)
         );
  AOI211_X1 U9354 ( .C1(n8565), .C2(n8975), .A(n7689), .B(n7688), .ZN(n7690)
         );
  OAI21_X1 U9355 ( .B1(n7692), .B2(n7691), .A(n7690), .ZN(P2_U3238) );
  NAND2_X1 U9356 ( .A1(n7694), .A2(n7693), .ZN(n7695) );
  NAND2_X1 U9357 ( .A1(n7696), .A2(n7695), .ZN(n7758) );
  NAND2_X1 U9358 ( .A1(n7706), .A2(n6707), .ZN(n7698) );
  NAND2_X1 U9359 ( .A1(n8113), .A2(n9525), .ZN(n7697) );
  NAND2_X1 U9360 ( .A1(n7698), .A2(n7697), .ZN(n7699) );
  XNOR2_X1 U9361 ( .A(n7699), .B(n8062), .ZN(n7752) );
  NOR2_X1 U9362 ( .A1(n8101), .A2(n7700), .ZN(n7701) );
  AOI21_X1 U9363 ( .B1(n7706), .B2(n6846), .A(n7701), .ZN(n7753) );
  XNOR2_X1 U9364 ( .A(n7752), .B(n7753), .ZN(n7702) );
  XNOR2_X1 U9365 ( .A(n7758), .B(n7702), .ZN(n7709) );
  OAI22_X1 U9366 ( .A1(n9108), .A2(n7703), .B1(n7762), .B2(n9106), .ZN(n7704)
         );
  AOI211_X1 U9367 ( .C1(n7915), .C2(n9120), .A(n7705), .B(n7704), .ZN(n7708)
         );
  NAND2_X1 U9368 ( .A1(n7706), .A2(n9100), .ZN(n7707) );
  OAI211_X1 U9369 ( .C1(n7709), .C2(n9095), .A(n7708), .B(n7707), .ZN(P1_U3232) );
  NAND2_X1 U9370 ( .A1(n8457), .A2(n7710), .ZN(n7712) );
  OAI211_X1 U9371 ( .C1(n8421), .C2(n7713), .A(n7712), .B(n7711), .ZN(P1_U3325) );
  OAI22_X1 U9372 ( .A1(n7715), .A2(n9853), .B1(n7714), .B2(n9851), .ZN(n7716)
         );
  AOI21_X1 U9373 ( .B1(n7717), .B2(n9845), .A(n7716), .ZN(n7718) );
  AND2_X1 U9374 ( .A1(n7719), .A2(n7718), .ZN(n7721) );
  MUX2_X1 U9375 ( .A(n5353), .B(n7721), .S(n9861), .Z(n7720) );
  INV_X1 U9376 ( .A(n7720), .ZN(P2_U3478) );
  MUX2_X1 U9377 ( .A(n6811), .B(n7721), .S(n9875), .Z(n7722) );
  INV_X1 U9378 ( .A(n7722), .ZN(P2_U3529) );
  INV_X1 U9379 ( .A(n8269), .ZN(n7723) );
  XNOR2_X1 U9380 ( .A(n7724), .B(n7723), .ZN(n7817) );
  OAI21_X1 U9381 ( .B1(n8269), .B2(n7726), .A(n7725), .ZN(n7727) );
  NAND2_X1 U9382 ( .A1(n7727), .A2(n9635), .ZN(n7729) );
  AOI22_X1 U9383 ( .A1(n9524), .A2(n9118), .B1(n9526), .B2(n9119), .ZN(n7728)
         );
  NAND2_X1 U9384 ( .A1(n7729), .A2(n7728), .ZN(n7730) );
  AOI21_X1 U9385 ( .B1(n7817), .B2(n7731), .A(n7730), .ZN(n7819) );
  OR2_X1 U9386 ( .A1(n7732), .A2(n7918), .ZN(n7733) );
  NAND2_X1 U9387 ( .A1(n9513), .A2(n7733), .ZN(n7815) );
  AOI22_X1 U9388 ( .A1(n4389), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n7911), .B2(
        n9653), .ZN(n7735) );
  NAND2_X1 U9389 ( .A1(n7908), .A2(n9531), .ZN(n7734) );
  OAI211_X1 U9390 ( .C1(n7815), .C2(n9198), .A(n7735), .B(n7734), .ZN(n7736)
         );
  AOI21_X1 U9391 ( .B1(n7817), .B2(n7737), .A(n7736), .ZN(n7738) );
  OAI21_X1 U9392 ( .B1(n7819), .B2(n4389), .A(n7738), .ZN(P1_U3276) );
  AOI21_X1 U9393 ( .B1(n7740), .B2(n8869), .A(n7739), .ZN(n8596) );
  XNOR2_X1 U9394 ( .A(n8596), .B(n8597), .ZN(n7741) );
  NOR2_X1 U9395 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7741), .ZN(n8598) );
  AOI21_X1 U9396 ( .B1(n7741), .B2(P2_REG2_REG_15__SCAN_IN), .A(n8598), .ZN(
        n7751) );
  OAI21_X1 U9397 ( .B1(n7743), .B2(P2_REG1_REG_14__SCAN_IN), .A(n7742), .ZN(
        n8587) );
  XNOR2_X1 U9398 ( .A(n8587), .B(n8588), .ZN(n7745) );
  INV_X1 U9399 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7744) );
  NOR2_X1 U9400 ( .A1(n7744), .A2(n7745), .ZN(n8589) );
  AOI211_X1 U9401 ( .C1(n7745), .C2(n7744), .A(n8589), .B(n9761), .ZN(n7749)
         );
  NOR2_X1 U9402 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5117), .ZN(n7746) );
  AOI21_X1 U9403 ( .B1(n9766), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7746), .ZN(
        n7747) );
  OAI21_X1 U9404 ( .B1(n9760), .B2(n8588), .A(n7747), .ZN(n7748) );
  NOR2_X1 U9405 ( .A1(n7749), .A2(n7748), .ZN(n7750) );
  OAI21_X1 U9406 ( .B1(n7751), .B2(n8633), .A(n7750), .ZN(P2_U3260) );
  AND2_X1 U9407 ( .A1(n7752), .A2(n7753), .ZN(n7757) );
  INV_X1 U9408 ( .A(n7752), .ZN(n7755) );
  INV_X1 U9409 ( .A(n7753), .ZN(n7754) );
  NAND2_X1 U9410 ( .A1(n7755), .A2(n7754), .ZN(n7756) );
  NAND2_X1 U9411 ( .A1(n7769), .A2(n6707), .ZN(n7760) );
  NAND2_X1 U9412 ( .A1(n8113), .A2(n9119), .ZN(n7759) );
  NAND2_X1 U9413 ( .A1(n7760), .A2(n7759), .ZN(n7761) );
  XNOR2_X1 U9414 ( .A(n7761), .B(n8062), .ZN(n7899) );
  NOR2_X1 U9415 ( .A1(n8101), .A2(n7762), .ZN(n7763) );
  AOI21_X1 U9416 ( .B1(n7769), .B2(n6846), .A(n7763), .ZN(n7896) );
  INV_X1 U9417 ( .A(n7896), .ZN(n7900) );
  XNOR2_X1 U9418 ( .A(n7899), .B(n7900), .ZN(n7764) );
  XNOR2_X1 U9419 ( .A(n7898), .B(n7764), .ZN(n7771) );
  AOI22_X1 U9420 ( .A1(n9089), .A2(n7765), .B1(n7915), .B2(n9525), .ZN(n7767)
         );
  OAI211_X1 U9421 ( .C1(n7975), .C2(n9106), .A(n7767), .B(n7766), .ZN(n7768)
         );
  AOI21_X1 U9422 ( .B1(n7769), .B2(n9100), .A(n7768), .ZN(n7770) );
  OAI21_X1 U9423 ( .B1(n7771), .B2(n9095), .A(n7770), .ZN(P1_U3213) );
  XNOR2_X1 U9424 ( .A(n7772), .B(n7825), .ZN(n7777) );
  OAI21_X1 U9425 ( .B1(n9750), .B2(n8881), .A(n7773), .ZN(n7775) );
  OAI22_X1 U9426 ( .A1(n9751), .A2(n7788), .B1(n7790), .B2(n9759), .ZN(n7774)
         );
  AOI211_X1 U9427 ( .C1(n8565), .C2(n7837), .A(n7775), .B(n7774), .ZN(n7776)
         );
  OAI21_X1 U9428 ( .B1(n7777), .B2(n9743), .A(n7776), .ZN(P2_U3226) );
  AND2_X1 U9429 ( .A1(n7779), .A2(n8581), .ZN(n7781) );
  NAND2_X1 U9430 ( .A1(n8975), .A2(n8580), .ZN(n7836) );
  NAND2_X1 U9431 ( .A1(n4473), .A2(n7836), .ZN(n7783) );
  XNOR2_X1 U9432 ( .A(n7783), .B(n7834), .ZN(n9858) );
  INV_X1 U9433 ( .A(n9858), .ZN(n7796) );
  NAND2_X1 U9434 ( .A1(n7784), .A2(n7785), .ZN(n7786) );
  XNOR2_X1 U9435 ( .A(n7786), .B(n7834), .ZN(n7787) );
  OAI222_X1 U9436 ( .A1(n8882), .A2(n8881), .B1(n8880), .B2(n7788), .C1(n8877), 
        .C2(n7787), .ZN(n9855) );
  INV_X1 U9437 ( .A(n7837), .ZN(n9852) );
  INV_X1 U9438 ( .A(n7857), .ZN(n7789) );
  OAI21_X1 U9439 ( .B1(n9852), .B2(n7867), .A(n7789), .ZN(n9854) );
  OAI22_X1 U9440 ( .A1(n8870), .A2(n7791), .B1(n7790), .B2(n9778), .ZN(n7792)
         );
  AOI21_X1 U9441 ( .B1(n7837), .B2(n8872), .A(n7792), .ZN(n7793) );
  OAI21_X1 U9442 ( .B1(n9854), .B2(n8874), .A(n7793), .ZN(n7794) );
  AOI21_X1 U9443 ( .B1(n9855), .B2(n8870), .A(n7794), .ZN(n7795) );
  OAI21_X1 U9444 ( .B1(n8862), .B2(n7796), .A(n7795), .ZN(P2_U3284) );
  INV_X1 U9445 ( .A(n7797), .ZN(n7800) );
  OAI222_X1 U9446 ( .A1(n8419), .A2(n7800), .B1(n7799), .B2(P1_U3084), .C1(
        n7798), .C2(n8421), .ZN(P1_U3324) );
  OAI222_X1 U9447 ( .A1(n5091), .A2(P2_U3152), .B1(n4390), .B2(n7800), .C1(
        n10131), .C2(n8459), .ZN(P2_U3329) );
  INV_X1 U9448 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7814) );
  AOI21_X1 U9449 ( .B1(n7805), .B2(P1_REG1_REG_16__SCAN_IN), .A(n7801), .ZN(
        n7803) );
  XNOR2_X1 U9450 ( .A(n9163), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n7802) );
  NOR2_X1 U9451 ( .A1(n7803), .A2(n7802), .ZN(n9157) );
  AOI211_X1 U9452 ( .C1(n7803), .C2(n7802), .A(n9157), .B(n9608), .ZN(n7812)
         );
  NAND2_X1 U9453 ( .A1(n9163), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7806) );
  OAI21_X1 U9454 ( .B1(n9163), .B2(P1_REG2_REG_17__SCAN_IN), .A(n7806), .ZN(
        n7807) );
  AOI211_X1 U9455 ( .C1(n7808), .C2(n7807), .A(n9162), .B(n9598), .ZN(n7811)
         );
  NAND2_X1 U9456 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9045) );
  OAI21_X1 U9457 ( .B1(n9617), .B2(n7809), .A(n9045), .ZN(n7810) );
  NOR3_X1 U9458 ( .A1(n7812), .A2(n7811), .A3(n7810), .ZN(n7813) );
  OAI21_X1 U9459 ( .B1(n9619), .B2(n7814), .A(n7813), .ZN(P1_U3258) );
  INV_X1 U9460 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n7820) );
  INV_X1 U9461 ( .A(n9694), .ZN(n9687) );
  OAI22_X1 U9462 ( .A1(n7815), .A2(n9705), .B1(n7918), .B2(n9718), .ZN(n7816)
         );
  AOI21_X1 U9463 ( .B1(n7817), .B2(n9687), .A(n7816), .ZN(n7818) );
  AND2_X1 U9464 ( .A1(n7819), .A2(n7818), .ZN(n7822) );
  MUX2_X1 U9465 ( .A(n7820), .B(n7822), .S(n9726), .Z(n7821) );
  INV_X1 U9466 ( .A(n7821), .ZN(P1_U3499) );
  MUX2_X1 U9467 ( .A(n7823), .B(n7822), .S(n9742), .Z(n7824) );
  INV_X1 U9468 ( .A(n7824), .ZN(P1_U3538) );
  NAND2_X1 U9469 ( .A1(n7772), .A2(n7825), .ZN(n7827) );
  NAND2_X1 U9470 ( .A1(n7827), .A2(n7826), .ZN(n7829) );
  XNOR2_X1 U9471 ( .A(n7829), .B(n7828), .ZN(n7833) );
  OAI22_X1 U9472 ( .A1(n9750), .A2(n7999), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7243), .ZN(n7831) );
  OAI22_X1 U9473 ( .A1(n9751), .A2(n7849), .B1(n7854), .B2(n9759), .ZN(n7830)
         );
  AOI211_X1 U9474 ( .C1(n6166), .C2(n8565), .A(n7831), .B(n7830), .ZN(n7832)
         );
  OAI21_X1 U9475 ( .B1(n7833), .B2(n9743), .A(n7832), .ZN(P2_U3236) );
  INV_X1 U9476 ( .A(n7834), .ZN(n7835) );
  AND2_X1 U9477 ( .A1(n7836), .A2(n7835), .ZN(n7840) );
  OR2_X1 U9478 ( .A1(n7837), .A2(n8579), .ZN(n7838) );
  INV_X1 U9479 ( .A(n7838), .ZN(n7839) );
  OAI21_X1 U9480 ( .B1(n7841), .B2(n7847), .A(n7929), .ZN(n8971) );
  OR2_X1 U9481 ( .A1(n8971), .A2(n7842), .ZN(n7853) );
  NAND2_X1 U9482 ( .A1(n7843), .A2(n7846), .ZN(n7845) );
  NAND2_X1 U9483 ( .A1(n7845), .A2(n7844), .ZN(n8876) );
  NAND3_X1 U9484 ( .A1(n7843), .A2(n7847), .A3(n7846), .ZN(n7848) );
  NAND2_X1 U9485 ( .A1(n8876), .A2(n7848), .ZN(n7851) );
  OAI22_X1 U9486 ( .A1(n7849), .A2(n8880), .B1(n7999), .B2(n8882), .ZN(n7850)
         );
  AOI21_X1 U9487 ( .B1(n7851), .B2(n9777), .A(n7850), .ZN(n7852) );
  NAND2_X1 U9488 ( .A1(n7853), .A2(n7852), .ZN(n8973) );
  OAI22_X1 U9489 ( .A1(n8870), .A2(n7855), .B1(n7854), .B2(n9778), .ZN(n7856)
         );
  AOI21_X1 U9490 ( .B1(n6166), .B2(n8872), .A(n7856), .ZN(n7860) );
  INV_X1 U9491 ( .A(n6166), .ZN(n7928) );
  OR2_X1 U9492 ( .A1(n7857), .A2(n7928), .ZN(n7858) );
  AND2_X1 U9493 ( .A1(n8865), .A2(n7858), .ZN(n8969) );
  NAND2_X1 U9494 ( .A1(n8969), .A2(n8834), .ZN(n7859) );
  OAI211_X1 U9495 ( .C1(n8971), .C2(n7861), .A(n7860), .B(n7859), .ZN(n7862)
         );
  AOI21_X1 U9496 ( .B1(n8870), .B2(n8973), .A(n7862), .ZN(n7863) );
  INV_X1 U9497 ( .A(n7863), .ZN(P2_U3283) );
  NAND2_X1 U9498 ( .A1(n7865), .A2(n7864), .ZN(n7866) );
  XNOR2_X1 U9499 ( .A(n7866), .B(n7873), .ZN(n8979) );
  AOI21_X1 U9500 ( .B1(n8975), .B2(n7868), .A(n7867), .ZN(n8976) );
  INV_X1 U9501 ( .A(n7869), .ZN(n7870) );
  AOI22_X1 U9502 ( .A1(n4388), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7870), .B2(
        n8848), .ZN(n7871) );
  OAI21_X1 U9503 ( .B1(n4701), .B2(n8851), .A(n7871), .ZN(n7876) );
  XOR2_X1 U9504 ( .A(n7872), .B(n7873), .Z(n7874) );
  AOI222_X1 U9505 ( .A1(n9777), .A2(n7874), .B1(n8579), .B2(n9774), .C1(n8581), 
        .C2(n9772), .ZN(n8978) );
  NOR2_X1 U9506 ( .A1(n8978), .A2(n4388), .ZN(n7875) );
  AOI211_X1 U9507 ( .C1(n8976), .C2(n8834), .A(n7876), .B(n7875), .ZN(n7877)
         );
  OAI21_X1 U9508 ( .B1(n8862), .B2(n8979), .A(n7877), .ZN(P2_U3285) );
  NAND2_X1 U9509 ( .A1(n7772), .A2(n7878), .ZN(n7880) );
  AND2_X1 U9510 ( .A1(n7880), .A2(n7879), .ZN(n7882) );
  XNOR2_X1 U9511 ( .A(n7882), .B(n7881), .ZN(n7886) );
  OAI22_X1 U9512 ( .A1(n9750), .A2(n8859), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5425), .ZN(n7884) );
  OAI22_X1 U9513 ( .A1(n9751), .A2(n8858), .B1(n8847), .B2(n9759), .ZN(n7883)
         );
  AOI211_X1 U9514 ( .C1(n8960), .C2(n8565), .A(n7884), .B(n7883), .ZN(n7885)
         );
  OAI21_X1 U9515 ( .B1(n7886), .B2(n9743), .A(n7885), .ZN(P2_U3230) );
  XOR2_X1 U9516 ( .A(n8270), .B(n7887), .Z(n9442) );
  AOI211_X1 U9517 ( .C1(n9440), .C2(n9514), .A(n9705), .B(n9364), .ZN(n9439)
         );
  NOR2_X1 U9518 ( .A1(n7888), .A2(n9370), .ZN(n7891) );
  INV_X1 U9519 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n7889) );
  OAI22_X1 U9520 ( .A1(n9665), .A2(n7889), .B1(n9048), .B2(n9629), .ZN(n7890)
         );
  AOI211_X1 U9521 ( .C1(n9439), .C2(n9539), .A(n7891), .B(n7890), .ZN(n7895)
         );
  XNOR2_X1 U9522 ( .A(n7892), .B(n8270), .ZN(n7893) );
  OAI222_X1 U9523 ( .A1(n9662), .A2(n9047), .B1(n9660), .B2(n9046), .C1(n7893), 
        .C2(n9657), .ZN(n9438) );
  NAND2_X1 U9524 ( .A1(n9438), .A2(n9665), .ZN(n7894) );
  OAI211_X1 U9525 ( .C1(n9442), .C2(n9374), .A(n7895), .B(n7894), .ZN(P1_U3274) );
  NAND2_X1 U9526 ( .A1(n7899), .A2(n7896), .ZN(n7897) );
  NAND2_X1 U9527 ( .A1(n7898), .A2(n7897), .ZN(n7903) );
  INV_X1 U9528 ( .A(n7899), .ZN(n7901) );
  NAND2_X1 U9529 ( .A1(n7901), .A2(n7900), .ZN(n7902) );
  NAND2_X1 U9530 ( .A1(n7908), .A2(n6707), .ZN(n7905) );
  NAND2_X1 U9531 ( .A1(n8113), .A2(n9503), .ZN(n7904) );
  NAND2_X1 U9532 ( .A1(n7905), .A2(n7904), .ZN(n7906) );
  XNOR2_X1 U9533 ( .A(n7906), .B(n8062), .ZN(n7958) );
  NOR2_X1 U9534 ( .A1(n8101), .A2(n7975), .ZN(n7907) );
  AOI21_X1 U9535 ( .B1(n7908), .B2(n8113), .A(n7907), .ZN(n7959) );
  XNOR2_X1 U9536 ( .A(n7958), .B(n7959), .ZN(n7909) );
  XNOR2_X1 U9537 ( .A(n7957), .B(n7909), .ZN(n7910) );
  NAND2_X1 U9538 ( .A1(n7910), .A2(n9102), .ZN(n7917) );
  INV_X1 U9539 ( .A(n7911), .ZN(n7912) );
  OAI22_X1 U9540 ( .A1(n9108), .A2(n7912), .B1(n9046), .B2(n9106), .ZN(n7913)
         );
  AOI211_X1 U9541 ( .C1(n7915), .C2(n9119), .A(n7914), .B(n7913), .ZN(n7916)
         );
  OAI211_X1 U9542 ( .C1(n7918), .C2(n9115), .A(n7917), .B(n7916), .ZN(P1_U3239) );
  NAND2_X1 U9543 ( .A1(n8876), .A2(n7919), .ZN(n8885) );
  NAND2_X1 U9544 ( .A1(n8885), .A2(n7920), .ZN(n7925) );
  AND2_X1 U9545 ( .A1(n7922), .A2(n7921), .ZN(n7923) );
  OAI211_X1 U9546 ( .C1(n7925), .C2(n7924), .A(n7923), .B(n9777), .ZN(n7927)
         );
  INV_X1 U9547 ( .A(n8858), .ZN(n8575) );
  AOI22_X1 U9548 ( .A1(n9774), .A2(n8575), .B1(n8577), .B2(n9772), .ZN(n7926)
         );
  AND2_X1 U9549 ( .A1(n7927), .A2(n7926), .ZN(n8967) );
  NAND2_X1 U9550 ( .A1(n7930), .A2(n6170), .ZN(n7984) );
  OAI21_X1 U9551 ( .B1(n7930), .B2(n6170), .A(n7984), .ZN(n8963) );
  NAND2_X1 U9552 ( .A1(n8963), .A2(n9787), .ZN(n7936) );
  INV_X1 U9553 ( .A(n7987), .ZN(n7931) );
  AOI21_X1 U9554 ( .B1(n8964), .B2(n8867), .A(n7931), .ZN(n8965) );
  NOR2_X1 U9555 ( .A1(n4707), .A2(n8851), .ZN(n7934) );
  OAI22_X1 U9556 ( .A1(n8870), .A2(n7932), .B1(n8000), .B2(n9778), .ZN(n7933)
         );
  AOI211_X1 U9557 ( .C1(n8965), .C2(n8834), .A(n7934), .B(n7933), .ZN(n7935)
         );
  OAI211_X1 U9558 ( .C1(n4388), .C2(n8967), .A(n7936), .B(n7935), .ZN(P2_U3281) );
  NAND2_X1 U9559 ( .A1(n7772), .A2(n7937), .ZN(n7940) );
  NAND2_X1 U9560 ( .A1(n7940), .A2(n7938), .ZN(n7942) );
  AND2_X1 U9561 ( .A1(n7940), .A2(n7939), .ZN(n7941) );
  AOI21_X1 U9562 ( .B1(n7943), .B2(n7942), .A(n7941), .ZN(n7948) );
  OAI21_X1 U9563 ( .B1(n9750), .B2(n8883), .A(n7944), .ZN(n7946) );
  OAI22_X1 U9564 ( .A1(n9751), .A2(n8881), .B1(n8868), .B2(n9759), .ZN(n7945)
         );
  AOI211_X1 U9565 ( .C1(n9491), .C2(n8565), .A(n7946), .B(n7945), .ZN(n7947)
         );
  OAI21_X1 U9566 ( .B1(n7948), .B2(n9743), .A(n7947), .ZN(P2_U3217) );
  XNOR2_X1 U9567 ( .A(n7950), .B(n7949), .ZN(n7955) );
  INV_X1 U9568 ( .A(n7951), .ZN(n8835) );
  INV_X1 U9569 ( .A(n8830), .ZN(n8574) );
  AOI22_X1 U9570 ( .A1(n8511), .A2(n8835), .B1(n8554), .B2(n8574), .ZN(n7952)
         );
  NAND2_X1 U9571 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8623) );
  OAI211_X1 U9572 ( .C1(n8831), .C2(n9750), .A(n7952), .B(n8623), .ZN(n7953)
         );
  AOI21_X1 U9573 ( .B1(n8953), .B2(n8565), .A(n7953), .ZN(n7954) );
  OAI21_X1 U9574 ( .B1(n7955), .B2(n9743), .A(n7954), .ZN(P2_U3240) );
  NAND2_X1 U9575 ( .A1(n7958), .A2(n7959), .ZN(n7956) );
  INV_X1 U9576 ( .A(n7958), .ZN(n7961) );
  INV_X1 U9577 ( .A(n7959), .ZN(n7960) );
  NAND2_X1 U9578 ( .A1(n7961), .A2(n7960), .ZN(n7962) );
  NAND2_X1 U9579 ( .A1(n9549), .A2(n6707), .ZN(n7964) );
  NAND2_X1 U9580 ( .A1(n9118), .A2(n8113), .ZN(n7963) );
  NAND2_X1 U9581 ( .A1(n7964), .A2(n7963), .ZN(n7965) );
  XNOR2_X1 U9582 ( .A(n7965), .B(n6738), .ZN(n7971) );
  INV_X1 U9583 ( .A(n7971), .ZN(n7969) );
  NAND2_X1 U9584 ( .A1(n9549), .A2(n8113), .ZN(n7967) );
  NAND2_X1 U9585 ( .A1(n6764), .A2(n9118), .ZN(n7966) );
  NAND2_X1 U9586 ( .A1(n7967), .A2(n7966), .ZN(n7970) );
  INV_X1 U9587 ( .A(n7970), .ZN(n7968) );
  NAND2_X1 U9588 ( .A1(n7969), .A2(n7968), .ZN(n9041) );
  INV_X1 U9589 ( .A(n9041), .ZN(n7972) );
  AND2_X1 U9590 ( .A1(n7971), .A2(n7970), .ZN(n9040) );
  NOR2_X1 U9591 ( .A1(n7972), .A2(n9040), .ZN(n7973) );
  XNOR2_X1 U9592 ( .A(n8039), .B(n7973), .ZN(n7979) );
  OAI21_X1 U9593 ( .B1(n9110), .B2(n7975), .A(n7974), .ZN(n7977) );
  OAI22_X1 U9594 ( .A1(n9108), .A2(n9507), .B1(n9362), .B2(n9106), .ZN(n7976)
         );
  AOI211_X1 U9595 ( .C1(n9549), .C2(n9100), .A(n7977), .B(n7976), .ZN(n7978)
         );
  OAI21_X1 U9596 ( .B1(n7979), .B2(n9095), .A(n7978), .ZN(P1_U3224) );
  XOR2_X1 U9597 ( .A(n7986), .B(n7980), .Z(n7983) );
  NOR2_X1 U9598 ( .A1(n8830), .A2(n8882), .ZN(n7982) );
  NOR2_X1 U9599 ( .A1(n8883), .A2(n8880), .ZN(n7981) );
  OR2_X1 U9600 ( .A1(n7982), .A2(n7981), .ZN(n8524) );
  AOI21_X1 U9601 ( .B1(n7983), .B2(n9777), .A(n8524), .ZN(n9487) );
  INV_X1 U9602 ( .A(n8883), .ZN(n8576) );
  AOI21_X1 U9603 ( .B1(n7986), .B2(n7985), .A(n8434), .ZN(n9490) );
  AND2_X1 U9604 ( .A1(n7987), .A2(n8522), .ZN(n7988) );
  OR2_X1 U9605 ( .A1(n7988), .A2(n8843), .ZN(n9488) );
  OAI22_X1 U9606 ( .A1(n8870), .A2(n7989), .B1(n8527), .B2(n9778), .ZN(n7990)
         );
  AOI21_X1 U9607 ( .B1(n8522), .B2(n8872), .A(n7990), .ZN(n7991) );
  OAI21_X1 U9608 ( .B1(n9488), .B2(n8874), .A(n7991), .ZN(n7992) );
  AOI21_X1 U9609 ( .B1(n9490), .B2(n9787), .A(n7992), .ZN(n7993) );
  OAI21_X1 U9610 ( .B1(n4388), .B2(n9487), .A(n7993), .ZN(P2_U3280) );
  NAND2_X1 U9611 ( .A1(n8518), .A2(n8544), .ZN(n7998) );
  NAND2_X1 U9612 ( .A1(n8533), .A2(n8576), .ZN(n7997) );
  NAND2_X1 U9613 ( .A1(n7772), .A2(n7994), .ZN(n7996) );
  XNOR2_X1 U9614 ( .A(n8516), .B(n8517), .ZN(n8519) );
  MUX2_X1 U9615 ( .A(n7998), .B(n7997), .S(n8519), .Z(n8004) );
  OAI22_X1 U9616 ( .A1(n9751), .A2(n7999), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5117), .ZN(n8002) );
  OAI22_X1 U9617 ( .A1(n9750), .A2(n8858), .B1(n9759), .B2(n8000), .ZN(n8001)
         );
  AOI211_X1 U9618 ( .C1(n8964), .C2(n8565), .A(n8002), .B(n8001), .ZN(n8003)
         );
  NAND2_X1 U9619 ( .A1(n8004), .A2(n8003), .ZN(P2_U3243) );
  NOR4_X1 U9620 ( .A1(n8005), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n8006), .ZN(n8007) );
  AOI21_X1 U9621 ( .B1(n8008), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n8007), .ZN(
        n8009) );
  OAI21_X1 U9622 ( .B1(n8138), .B2(n8419), .A(n8009), .ZN(P1_U3322) );
  INV_X1 U9623 ( .A(n8010), .ZN(n8012) );
  NOR4_X1 U9624 ( .A1(n8012), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8011), .A4(
        P2_U3152), .ZN(n8013) );
  AOI21_X1 U9625 ( .B1(n8014), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8013), .ZN(
        n8015) );
  OAI21_X1 U9626 ( .B1(n8138), .B2(n4390), .A(n8015), .ZN(P2_U3327) );
  INV_X1 U9627 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8141) );
  INV_X1 U9628 ( .A(n8140), .ZN(n8432) );
  OAI222_X1 U9629 ( .A1(n8421), .A2(n8141), .B1(n8419), .B2(n8432), .C1(
        P1_U3084), .C2(n5737), .ZN(P1_U3323) );
  INV_X1 U9630 ( .A(n8960), .ZN(n8852) );
  NAND2_X1 U9631 ( .A1(n8843), .A2(n8852), .ZN(n8844) );
  NAND2_X1 U9632 ( .A1(n8897), .A2(n8656), .ZN(n8893) );
  NAND2_X1 U9633 ( .A1(n8017), .A2(P2_B_REG_SCAN_IN), .ZN(n8018) );
  AND2_X1 U9634 ( .A1(n9774), .A2(n8018), .ZN(n8450) );
  NAND2_X1 U9635 ( .A1(n8019), .A2(n8450), .ZN(n8895) );
  NOR2_X1 U9636 ( .A1(n8895), .A2(n4388), .ZN(n8658) );
  AOI21_X1 U9637 ( .B1(n4388), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8658), .ZN(
        n8021) );
  NAND2_X1 U9638 ( .A1(n8890), .A2(n8872), .ZN(n8020) );
  OAI211_X1 U9639 ( .C1(n8892), .C2(n8874), .A(n8021), .B(n8020), .ZN(P2_U3265) );
  INV_X1 U9640 ( .A(n8022), .ZN(n8023) );
  AOI211_X1 U9641 ( .C1(n8025), .C2(n8024), .A(n9743), .B(n8023), .ZN(n8030)
         );
  OAI22_X1 U9642 ( .A1(n8425), .A2(n8026), .B1(n9747), .B2(n9811), .ZN(n8029)
         );
  OAI22_X1 U9643 ( .A1(n8027), .A2(n9750), .B1(n9751), .B2(n7002), .ZN(n8028)
         );
  OR3_X1 U9644 ( .A1(n8030), .A2(n8029), .A3(n8028), .ZN(P2_U3239) );
  INV_X1 U9645 ( .A(n8770), .ZN(n8033) );
  OAI22_X1 U9646 ( .A1(n8746), .A2(n8882), .B1(n8562), .B2(n8880), .ZN(n8776)
         );
  AOI22_X1 U9647 ( .A1(n8776), .A2(n8523), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8032) );
  OAI21_X1 U9648 ( .B1(n8033), .B2(n9759), .A(n8032), .ZN(n8036) );
  NOR3_X1 U9649 ( .A1(n8034), .A2(n8572), .A3(n8552), .ZN(n8035) );
  AOI211_X1 U9650 ( .C1(n8565), .C2(n8932), .A(n8036), .B(n8035), .ZN(n8037)
         );
  OAI21_X1 U9651 ( .B1(n8031), .B2(n9743), .A(n8037), .ZN(P2_U3237) );
  NOR2_X1 U9652 ( .A1(n8101), .A2(n9269), .ZN(n8038) );
  AOI21_X1 U9653 ( .B1(n9408), .B2(n8113), .A(n8038), .ZN(n9011) );
  NAND2_X1 U9654 ( .A1(n9440), .A2(n6707), .ZN(n8041) );
  NAND2_X1 U9655 ( .A1(n9504), .A2(n8113), .ZN(n8040) );
  NAND2_X1 U9656 ( .A1(n8041), .A2(n8040), .ZN(n8042) );
  XNOR2_X1 U9657 ( .A(n8042), .B(n6738), .ZN(n8046) );
  INV_X1 U9658 ( .A(n8046), .ZN(n8044) );
  AND2_X1 U9659 ( .A1(n9504), .A2(n6764), .ZN(n8043) );
  AOI21_X1 U9660 ( .B1(n9440), .B2(n8113), .A(n8043), .ZN(n8045) );
  NAND2_X1 U9661 ( .A1(n8044), .A2(n8045), .ZN(n8048) );
  INV_X1 U9662 ( .A(n8048), .ZN(n8047) );
  XNOR2_X1 U9663 ( .A(n8046), .B(n8045), .ZN(n9044) );
  NOR2_X1 U9664 ( .A1(n8047), .A2(n9044), .ZN(n8050) );
  AND2_X1 U9665 ( .A1(n9041), .A2(n8048), .ZN(n8049) );
  NAND2_X1 U9666 ( .A1(n9435), .A2(n6707), .ZN(n8052) );
  NAND2_X1 U9667 ( .A1(n9346), .A2(n6846), .ZN(n8051) );
  NAND2_X1 U9668 ( .A1(n8052), .A2(n8051), .ZN(n8053) );
  XNOR2_X1 U9669 ( .A(n8053), .B(n8062), .ZN(n8057) );
  NAND2_X1 U9670 ( .A1(n9435), .A2(n8113), .ZN(n8055) );
  NAND2_X1 U9671 ( .A1(n9346), .A2(n6764), .ZN(n8054) );
  NAND2_X1 U9672 ( .A1(n8055), .A2(n8054), .ZN(n9093) );
  NAND2_X1 U9673 ( .A1(n9092), .A2(n9093), .ZN(n9091) );
  INV_X1 U9674 ( .A(n8056), .ZN(n8059) );
  INV_X1 U9675 ( .A(n8057), .ZN(n8058) );
  NAND2_X1 U9676 ( .A1(n8059), .A2(n8058), .ZN(n9096) );
  NAND2_X1 U9677 ( .A1(n9429), .A2(n6707), .ZN(n8061) );
  NAND2_X1 U9678 ( .A1(n8113), .A2(n9332), .ZN(n8060) );
  NAND2_X1 U9679 ( .A1(n8061), .A2(n8060), .ZN(n8063) );
  XNOR2_X1 U9680 ( .A(n8063), .B(n8062), .ZN(n8066) );
  NOR2_X1 U9681 ( .A1(n8101), .A2(n9363), .ZN(n8064) );
  AOI21_X1 U9682 ( .B1(n9429), .B2(n8113), .A(n8064), .ZN(n8065) );
  XNOR2_X1 U9683 ( .A(n8066), .B(n8065), .ZN(n9018) );
  NAND2_X1 U9684 ( .A1(n8066), .A2(n8065), .ZN(n8067) );
  NAND2_X1 U9685 ( .A1(n9423), .A2(n6707), .ZN(n8069) );
  NAND2_X1 U9686 ( .A1(n6846), .A2(n9347), .ZN(n8068) );
  NAND2_X1 U9687 ( .A1(n8069), .A2(n8068), .ZN(n8070) );
  XNOR2_X1 U9688 ( .A(n8070), .B(n6738), .ZN(n8072) );
  NOR2_X1 U9689 ( .A1(n8101), .A2(n9318), .ZN(n8071) );
  AOI21_X1 U9690 ( .B1(n9423), .B2(n6846), .A(n8071), .ZN(n8073) );
  XNOR2_X1 U9691 ( .A(n8072), .B(n8073), .ZN(n9072) );
  INV_X1 U9692 ( .A(n8072), .ZN(n8074) );
  NAND2_X1 U9693 ( .A1(n9420), .A2(n6707), .ZN(n8076) );
  NAND2_X1 U9694 ( .A1(n6846), .A2(n9333), .ZN(n8075) );
  NAND2_X1 U9695 ( .A1(n8076), .A2(n8075), .ZN(n8077) );
  XNOR2_X1 U9696 ( .A(n8077), .B(n6738), .ZN(n8079) );
  NOR2_X1 U9697 ( .A1(n8101), .A2(n9083), .ZN(n8078) );
  AOI21_X1 U9698 ( .B1(n9420), .B2(n6846), .A(n8078), .ZN(n8080) );
  XNOR2_X1 U9699 ( .A(n8079), .B(n8080), .ZN(n9025) );
  NAND2_X1 U9700 ( .A1(n9024), .A2(n9025), .ZN(n8083) );
  INV_X1 U9701 ( .A(n8079), .ZN(n8081) );
  NAND2_X1 U9702 ( .A1(n8081), .A2(n8080), .ZN(n8082) );
  NAND2_X1 U9703 ( .A1(n8083), .A2(n8082), .ZN(n8089) );
  NOR2_X1 U9704 ( .A1(n8101), .A2(n9319), .ZN(n8084) );
  AOI21_X1 U9705 ( .B1(n9413), .B2(n8113), .A(n8084), .ZN(n8088) );
  NAND2_X2 U9706 ( .A1(n8089), .A2(n8088), .ZN(n9077) );
  NAND2_X1 U9707 ( .A1(n9413), .A2(n6707), .ZN(n8086) );
  NAND2_X1 U9708 ( .A1(n8113), .A2(n9287), .ZN(n8085) );
  NAND2_X1 U9709 ( .A1(n8086), .A2(n8085), .ZN(n8087) );
  XNOR2_X1 U9710 ( .A(n8087), .B(n6738), .ZN(n9080) );
  NAND2_X1 U9711 ( .A1(n9408), .A2(n6707), .ZN(n8091) );
  NAND2_X1 U9712 ( .A1(n6846), .A2(n9905), .ZN(n8090) );
  NAND2_X1 U9713 ( .A1(n8091), .A2(n8090), .ZN(n8092) );
  XNOR2_X1 U9714 ( .A(n8092), .B(n6738), .ZN(n8093) );
  AOI22_X1 U9715 ( .A1(n9405), .A2(n6846), .B1(n6764), .B2(n9286), .ZN(n8097)
         );
  NAND2_X1 U9716 ( .A1(n9405), .A2(n6707), .ZN(n8095) );
  NAND2_X1 U9717 ( .A1(n8113), .A2(n9286), .ZN(n8094) );
  NAND2_X1 U9718 ( .A1(n8095), .A2(n8094), .ZN(n8096) );
  XNOR2_X1 U9719 ( .A(n8096), .B(n6738), .ZN(n8099) );
  XOR2_X1 U9720 ( .A(n8097), .B(n8099), .Z(n9054) );
  INV_X1 U9721 ( .A(n8097), .ZN(n8098) );
  NOR2_X1 U9722 ( .A1(n8101), .A2(n9268), .ZN(n8102) );
  AOI21_X1 U9723 ( .B1(n9398), .B2(n8113), .A(n8102), .ZN(n8104) );
  AOI22_X1 U9724 ( .A1(n9398), .A2(n6707), .B1(n6846), .B2(n9243), .ZN(n8103)
         );
  XNOR2_X1 U9725 ( .A(n8103), .B(n6738), .ZN(n8105) );
  XOR2_X1 U9726 ( .A(n8104), .B(n8105), .Z(n9032) );
  AOI22_X1 U9727 ( .A1(n9393), .A2(n8113), .B1(n6764), .B2(n9259), .ZN(n8108)
         );
  AOI22_X1 U9728 ( .A1(n9393), .A2(n6707), .B1(n6846), .B2(n9259), .ZN(n8106)
         );
  XNOR2_X1 U9729 ( .A(n8106), .B(n6738), .ZN(n8107) );
  XOR2_X1 U9730 ( .A(n8108), .B(n8107), .Z(n9104) );
  NAND2_X1 U9731 ( .A1(n9105), .A2(n9104), .ZN(n9103) );
  INV_X1 U9732 ( .A(n8108), .ZN(n8109) );
  AOI22_X1 U9733 ( .A1(n9388), .A2(n6707), .B1(n6846), .B2(n9244), .ZN(n8112)
         );
  XOR2_X1 U9734 ( .A(n6738), .B(n8112), .Z(n9003) );
  AOI22_X1 U9735 ( .A1(n9388), .A2(n8113), .B1(n6764), .B2(n9244), .ZN(n9002)
         );
  INV_X1 U9736 ( .A(n9002), .ZN(n8114) );
  AOI22_X1 U9737 ( .A1(n9383), .A2(n6707), .B1(n6846), .B2(n9117), .ZN(n8117)
         );
  AOI22_X1 U9738 ( .A1(n9383), .A2(n6846), .B1(n6764), .B2(n9117), .ZN(n8115)
         );
  XNOR2_X1 U9739 ( .A(n8115), .B(n6738), .ZN(n8116) );
  OAI22_X1 U9740 ( .A1(n9110), .A2(n9107), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8119), .ZN(n8121) );
  OAI22_X1 U9741 ( .A1(n9108), .A2(n9205), .B1(n8230), .B2(n9106), .ZN(n8120)
         );
  AOI211_X1 U9742 ( .C1(n9383), .C2(n9100), .A(n8121), .B(n8120), .ZN(n8122)
         );
  NAND3_X1 U9743 ( .A1(n8533), .A2(n8123), .A3(n9773), .ZN(n8124) );
  OAI21_X1 U9744 ( .B1(n9755), .B2(n9743), .A(n8124), .ZN(n8127) );
  INV_X1 U9745 ( .A(n8125), .ZN(n8126) );
  NAND2_X1 U9746 ( .A1(n8127), .A2(n8126), .ZN(n8134) );
  INV_X1 U9747 ( .A(n9779), .ZN(n8132) );
  OAI21_X1 U9748 ( .B1(n9747), .B2(n9785), .A(n8128), .ZN(n8131) );
  OAI22_X1 U9749 ( .A1(n8547), .A2(n9751), .B1(n9750), .B2(n8129), .ZN(n8130)
         );
  AOI211_X1 U9750 ( .C1(n8132), .C2(n8511), .A(n8131), .B(n8130), .ZN(n8133)
         );
  OAI211_X1 U9751 ( .C1(n9743), .C2(n8135), .A(n8134), .B(n8133), .ZN(P2_U3241) );
  INV_X1 U9752 ( .A(n8230), .ZN(n9212) );
  OR2_X1 U9753 ( .A1(n4387), .A2(n6808), .ZN(n8136) );
  NAND2_X1 U9754 ( .A1(n9375), .A2(n8231), .ZN(n8407) );
  NAND2_X1 U9755 ( .A1(n8140), .A2(n8139), .ZN(n8143) );
  OR2_X1 U9756 ( .A1(n4387), .A2(n8141), .ZN(n8142) );
  AND2_X1 U9757 ( .A1(n9194), .A2(n9116), .ZN(n8404) );
  NAND2_X1 U9758 ( .A1(n8404), .A2(n9375), .ZN(n8144) );
  NOR2_X1 U9759 ( .A1(n8354), .A2(n8236), .ZN(n8145) );
  MUX2_X1 U9760 ( .A(n9212), .B(n8145), .S(n8232), .Z(n8229) );
  NAND2_X1 U9761 ( .A1(n8394), .A2(n8388), .ZN(n8339) );
  NAND2_X1 U9762 ( .A1(n8339), .A2(n9255), .ZN(n8146) );
  AND2_X1 U9763 ( .A1(n8396), .A2(n8146), .ZN(n8150) );
  AND2_X1 U9764 ( .A1(n8394), .A2(n8147), .ZN(n8148) );
  NOR2_X1 U9765 ( .A1(n8343), .A2(n8148), .ZN(n8149) );
  MUX2_X1 U9766 ( .A(n8150), .B(n8149), .S(n4608), .Z(n8208) );
  NAND2_X1 U9767 ( .A1(n8293), .A2(n8168), .ZN(n8151) );
  AND2_X1 U9768 ( .A1(n8151), .A2(n8170), .ZN(n8174) );
  MUX2_X1 U9769 ( .A(n8152), .B(n9634), .S(n8232), .Z(n8159) );
  NAND2_X1 U9770 ( .A1(n8159), .A2(n8302), .ZN(n8155) );
  INV_X1 U9771 ( .A(n8158), .ZN(n8153) );
  NOR2_X1 U9772 ( .A1(n8154), .A2(n8153), .ZN(n8288) );
  NAND2_X1 U9773 ( .A1(n8155), .A2(n8288), .ZN(n8157) );
  NAND2_X1 U9774 ( .A1(n8159), .A2(n8158), .ZN(n8161) );
  NAND3_X1 U9775 ( .A1(n8161), .A2(n8160), .A3(n8302), .ZN(n8165) );
  NAND2_X1 U9776 ( .A1(n8176), .A2(n8162), .ZN(n8163) );
  NAND2_X1 U9777 ( .A1(n8166), .A2(n8176), .ZN(n8167) );
  AND2_X1 U9778 ( .A1(n8168), .A2(n8167), .ZN(n8287) );
  AND2_X1 U9779 ( .A1(n8170), .A2(n8169), .ZN(n8286) );
  AOI21_X1 U9780 ( .B1(n8172), .B2(n8286), .A(n8171), .ZN(n8173) );
  MUX2_X1 U9781 ( .A(n8174), .B(n8173), .S(n8232), .Z(n8186) );
  NAND2_X1 U9782 ( .A1(n8176), .A2(n8175), .ZN(n8305) );
  AOI21_X1 U9783 ( .B1(n8305), .B2(n8177), .A(n8232), .ZN(n8178) );
  NAND3_X1 U9784 ( .A1(n8179), .A2(n8286), .A3(n8178), .ZN(n8180) );
  NAND2_X1 U9785 ( .A1(n8180), .A2(n8269), .ZN(n8185) );
  MUX2_X1 U9786 ( .A(n9549), .B(n9118), .S(n8232), .Z(n8187) );
  INV_X1 U9787 ( .A(n8297), .ZN(n8181) );
  MUX2_X1 U9788 ( .A(n4725), .B(n8181), .S(n8232), .Z(n8182) );
  AOI21_X1 U9789 ( .B1(n8187), .B2(n8183), .A(n8182), .ZN(n8184) );
  OAI21_X1 U9790 ( .B1(n8186), .B2(n8185), .A(n8184), .ZN(n8191) );
  INV_X1 U9791 ( .A(n8187), .ZN(n8189) );
  NAND2_X1 U9792 ( .A1(n8189), .A2(n8188), .ZN(n8190) );
  NAND3_X1 U9793 ( .A1(n8191), .A2(n8270), .A3(n8190), .ZN(n8194) );
  AND2_X1 U9794 ( .A1(n9341), .A2(n8192), .ZN(n8283) );
  MUX2_X1 U9795 ( .A(n8283), .B(n8333), .S(n8232), .Z(n8193) );
  AND2_X1 U9796 ( .A1(n8326), .A2(n9341), .ZN(n8329) );
  AND2_X1 U9797 ( .A1(n8250), .A2(n8196), .ZN(n8330) );
  NAND3_X1 U9798 ( .A1(n8198), .A2(n8331), .A3(n8250), .ZN(n8197) );
  INV_X1 U9799 ( .A(n8198), .ZN(n8199) );
  NAND2_X1 U9800 ( .A1(n8331), .A2(n8200), .ZN(n8202) );
  AND2_X1 U9801 ( .A1(n8202), .A2(n8201), .ZN(n8204) );
  NAND2_X1 U9802 ( .A1(n9255), .A2(n8341), .ZN(n8364) );
  NOR2_X1 U9803 ( .A1(n8339), .A2(n8364), .ZN(n8205) );
  NAND2_X1 U9804 ( .A1(n8206), .A2(n8205), .ZN(n8207) );
  NAND2_X1 U9805 ( .A1(n8208), .A2(n8207), .ZN(n8218) );
  OAI21_X1 U9806 ( .B1(n9240), .B2(n8209), .A(n8348), .ZN(n8212) );
  NAND2_X1 U9807 ( .A1(n8398), .A2(n9259), .ZN(n8210) );
  NAND2_X1 U9808 ( .A1(n8346), .A2(n8210), .ZN(n8211) );
  MUX2_X1 U9809 ( .A(n8212), .B(n8211), .S(n8232), .Z(n8213) );
  OAI21_X1 U9810 ( .B1(n8218), .B2(n9227), .A(n8213), .ZN(n8221) );
  AND2_X1 U9811 ( .A1(n8396), .A2(n9228), .ZN(n8214) );
  AOI21_X1 U9812 ( .B1(n8218), .B2(n8214), .A(n8345), .ZN(n8215) );
  AOI21_X1 U9813 ( .B1(n8221), .B2(n8215), .A(n8351), .ZN(n8223) );
  INV_X1 U9814 ( .A(n8398), .ZN(n8216) );
  NOR2_X1 U9815 ( .A1(n9393), .A2(n8216), .ZN(n8217) );
  AOI21_X1 U9816 ( .B1(n8218), .B2(n8217), .A(n8397), .ZN(n8220) );
  INV_X1 U9817 ( .A(n8348), .ZN(n8219) );
  AOI21_X1 U9818 ( .B1(n8221), .B2(n8220), .A(n8219), .ZN(n8222) );
  MUX2_X1 U9819 ( .A(n8223), .B(n8222), .S(n8232), .Z(n8227) );
  MUX2_X1 U9820 ( .A(n8225), .B(n8224), .S(n8232), .Z(n8226) );
  AOI21_X1 U9821 ( .B1(n8227), .B2(n9211), .A(n8226), .ZN(n8240) );
  NAND2_X1 U9822 ( .A1(n9188), .A2(n9116), .ZN(n8228) );
  NAND2_X1 U9823 ( .A1(n9547), .A2(n8228), .ZN(n8237) );
  NAND3_X1 U9824 ( .A1(n8229), .A2(n8240), .A3(n8237), .ZN(n8245) );
  NAND2_X1 U9825 ( .A1(n8230), .A2(n8232), .ZN(n8239) );
  OR3_X1 U9826 ( .A1(n8354), .A2(n8236), .A3(n8239), .ZN(n8235) );
  OR2_X1 U9827 ( .A1(n9375), .A2(n8231), .ZN(n8360) );
  INV_X1 U9828 ( .A(n8237), .ZN(n8352) );
  NAND3_X1 U9829 ( .A1(n8407), .A2(n8352), .A3(n8232), .ZN(n8234) );
  NAND4_X1 U9830 ( .A1(n8237), .A2(n8236), .A3(n4608), .A4(n9212), .ZN(n8233)
         );
  AND4_X1 U9831 ( .A1(n8235), .A2(n8360), .A3(n8234), .A4(n8233), .ZN(n8244)
         );
  NAND3_X1 U9832 ( .A1(n8237), .A2(n4608), .A3(n8236), .ZN(n8238) );
  OAI21_X1 U9833 ( .B1(n8354), .B2(n8239), .A(n8238), .ZN(n8241) );
  NAND2_X1 U9834 ( .A1(n8241), .A2(n8240), .ZN(n8243) );
  NAND2_X1 U9835 ( .A1(n8354), .A2(n4608), .ZN(n8242) );
  NAND4_X1 U9836 ( .A1(n8245), .A2(n8244), .A3(n8243), .A4(n8242), .ZN(n8361)
         );
  OAI21_X1 U9837 ( .B1(n9194), .B2(n9116), .A(n8360), .ZN(n8408) );
  INV_X1 U9838 ( .A(n8407), .ZN(n8278) );
  INV_X1 U9839 ( .A(n8397), .ZN(n8342) );
  NAND2_X1 U9840 ( .A1(n8342), .A2(n8246), .ZN(n9241) );
  NOR2_X1 U9841 ( .A1(n8248), .A2(n8247), .ZN(n9301) );
  NAND2_X1 U9842 ( .A1(n8250), .A2(n8249), .ZN(n9331) );
  NOR3_X1 U9843 ( .A1(n8253), .A2(n8252), .A3(n8251), .ZN(n8254) );
  NAND4_X1 U9844 ( .A1(n8255), .A2(n8309), .A3(n8254), .A4(n8317), .ZN(n8260)
         );
  INV_X1 U9845 ( .A(n8315), .ZN(n8257) );
  NAND3_X1 U9846 ( .A1(n8322), .A2(n8257), .A3(n8256), .ZN(n8379) );
  NOR4_X1 U9847 ( .A1(n8260), .A2(n8259), .A3(n8379), .A4(n8258), .ZN(n8262)
         );
  NAND4_X1 U9848 ( .A1(n8264), .A2(n8263), .A3(n8262), .A4(n8261), .ZN(n8265)
         );
  NOR4_X1 U9849 ( .A1(n8267), .A2(n8266), .A3(n9522), .A4(n8265), .ZN(n8268)
         );
  NAND4_X1 U9850 ( .A1(n8270), .A2(n8269), .A3(n8268), .A4(n9510), .ZN(n8271)
         );
  NOR4_X1 U9851 ( .A1(n9331), .A2(n9342), .A3(n9360), .A4(n8271), .ZN(n8272)
         );
  NAND4_X1 U9852 ( .A1(n9284), .A2(n9301), .A3(n9306), .A4(n8272), .ZN(n8273)
         );
  NOR4_X1 U9853 ( .A1(n9241), .A2(n9257), .A3(n9266), .A4(n8273), .ZN(n8274)
         );
  NAND4_X1 U9854 ( .A1(n8276), .A2(n8275), .A3(n9211), .A4(n8274), .ZN(n8277)
         );
  NOR4_X1 U9855 ( .A1(n8408), .A2(n8278), .A3(n8404), .A4(n8277), .ZN(n8357)
         );
  OAI22_X1 U9856 ( .A1(n8361), .A2(n8279), .B1(n8367), .B2(n8357), .ZN(n8359)
         );
  INV_X1 U9857 ( .A(n8280), .ZN(n8282) );
  AND2_X1 U9858 ( .A1(n8282), .A2(n8281), .ZN(n8401) );
  INV_X1 U9859 ( .A(n8283), .ZN(n8285) );
  OR2_X1 U9860 ( .A1(n8285), .A2(n8284), .ZN(n8308) );
  INV_X1 U9861 ( .A(n8286), .ZN(n8306) );
  INV_X1 U9862 ( .A(n8287), .ZN(n8292) );
  INV_X1 U9863 ( .A(n8288), .ZN(n8289) );
  NAND2_X1 U9864 ( .A1(n8289), .A2(n8303), .ZN(n8290) );
  NOR2_X1 U9865 ( .A1(n8305), .A2(n8290), .ZN(n8291) );
  NOR2_X1 U9866 ( .A1(n8292), .A2(n8291), .ZN(n8294) );
  OAI21_X1 U9867 ( .B1(n8306), .B2(n8294), .A(n8293), .ZN(n8296) );
  NAND2_X1 U9868 ( .A1(n8296), .A2(n8295), .ZN(n8298) );
  OAI211_X1 U9869 ( .C1(n9549), .C2(n9046), .A(n8298), .B(n8297), .ZN(n8299)
         );
  INV_X1 U9870 ( .A(n8299), .ZN(n8300) );
  NOR2_X1 U9871 ( .A1(n8308), .A2(n8300), .ZN(n8382) );
  NAND3_X1 U9872 ( .A1(n8303), .A2(n8302), .A3(n8301), .ZN(n8304) );
  OR3_X1 U9873 ( .A1(n8306), .A2(n8305), .A3(n8304), .ZN(n8307) );
  OR3_X1 U9874 ( .A1(n8308), .A2(n4725), .A3(n8307), .ZN(n8385) );
  INV_X1 U9875 ( .A(n7157), .ZN(n8314) );
  INV_X1 U9876 ( .A(n8309), .ZN(n8310) );
  NAND2_X1 U9877 ( .A1(n8310), .A2(n8322), .ZN(n8312) );
  NAND2_X1 U9878 ( .A1(n8312), .A2(n8311), .ZN(n8376) );
  NAND2_X1 U9879 ( .A1(n8317), .A2(n8313), .ZN(n8365) );
  NOR3_X1 U9880 ( .A1(n8314), .A2(n8376), .A3(n8365), .ZN(n8325) );
  AOI21_X1 U9881 ( .B1(n8317), .B2(n8316), .A(n8315), .ZN(n8323) );
  INV_X1 U9882 ( .A(n8318), .ZN(n8321) );
  INV_X1 U9883 ( .A(n8319), .ZN(n8320) );
  NOR2_X1 U9884 ( .A1(n8379), .A2(n8320), .ZN(n8374) );
  AOI211_X1 U9885 ( .C1(n8323), .C2(n8322), .A(n8321), .B(n8374), .ZN(n8324)
         );
  NOR3_X1 U9886 ( .A1(n8385), .A2(n8325), .A3(n8324), .ZN(n8328) );
  INV_X1 U9887 ( .A(n8326), .ZN(n8327) );
  NOR2_X1 U9888 ( .A1(n4442), .A2(n8327), .ZN(n8387) );
  OAI21_X1 U9889 ( .B1(n8382), .B2(n8328), .A(n8387), .ZN(n8338) );
  INV_X1 U9890 ( .A(n8329), .ZN(n8332) );
  OAI211_X1 U9891 ( .C1(n8333), .C2(n8332), .A(n8331), .B(n8330), .ZN(n8334)
         );
  INV_X1 U9892 ( .A(n8334), .ZN(n8335) );
  OR2_X1 U9893 ( .A1(n4442), .A2(n8335), .ZN(n8337) );
  AND2_X1 U9894 ( .A1(n8337), .A2(n8336), .ZN(n8389) );
  NAND2_X1 U9895 ( .A1(n8338), .A2(n8389), .ZN(n8340) );
  AOI21_X1 U9896 ( .B1(n8341), .B2(n8340), .A(n8339), .ZN(n8344) );
  OAI211_X1 U9897 ( .C1(n8344), .C2(n8343), .A(n8342), .B(n8396), .ZN(n8350)
         );
  NAND2_X1 U9898 ( .A1(n8346), .A2(n8345), .ZN(n8347) );
  AND3_X1 U9899 ( .A1(n8349), .A2(n8348), .A3(n8347), .ZN(n8400) );
  OAI21_X1 U9900 ( .B1(n8351), .B2(n8350), .A(n8400), .ZN(n8353) );
  AOI211_X1 U9901 ( .C1(n8401), .C2(n8353), .A(n8363), .B(n8352), .ZN(n8355)
         );
  OAI21_X1 U9902 ( .B1(n8355), .B2(n8354), .A(n8360), .ZN(n8356) );
  MUX2_X1 U9903 ( .A(n8357), .B(n8356), .S(n8367), .Z(n8358) );
  AND4_X1 U9904 ( .A1(n8361), .A2(n8367), .A3(n8360), .A4(n6149), .ZN(n8362)
         );
  INV_X1 U9905 ( .A(n8363), .ZN(n8406) );
  INV_X1 U9906 ( .A(n8364), .ZN(n8393) );
  INV_X1 U9907 ( .A(n8365), .ZN(n8380) );
  NAND2_X1 U9908 ( .A1(n9130), .A2(n9671), .ZN(n8366) );
  NAND3_X1 U9909 ( .A1(n8368), .A2(n8367), .A3(n8366), .ZN(n8369) );
  NAND2_X1 U9910 ( .A1(n8370), .A2(n8369), .ZN(n8372) );
  OAI21_X1 U9911 ( .B1(n8373), .B2(n8372), .A(n8371), .ZN(n8375) );
  NAND2_X1 U9912 ( .A1(n8375), .A2(n8374), .ZN(n8378) );
  INV_X1 U9913 ( .A(n8376), .ZN(n8377) );
  OAI211_X1 U9914 ( .C1(n8380), .C2(n8379), .A(n8378), .B(n8377), .ZN(n8381)
         );
  INV_X1 U9915 ( .A(n8381), .ZN(n8384) );
  INV_X1 U9916 ( .A(n8382), .ZN(n8383) );
  OAI21_X1 U9917 ( .B1(n8385), .B2(n8384), .A(n8383), .ZN(n8386) );
  INV_X1 U9918 ( .A(n8386), .ZN(n8391) );
  INV_X1 U9919 ( .A(n8387), .ZN(n8390) );
  OAI211_X1 U9920 ( .C1(n8391), .C2(n8390), .A(n8389), .B(n8388), .ZN(n8392)
         );
  NAND2_X1 U9921 ( .A1(n8393), .A2(n8392), .ZN(n8395) );
  NAND3_X1 U9922 ( .A1(n8396), .A2(n8395), .A3(n8394), .ZN(n8399) );
  AOI211_X1 U9923 ( .C1(n8399), .C2(n8398), .A(n8397), .B(n9227), .ZN(n8403)
         );
  INV_X1 U9924 ( .A(n8400), .ZN(n8402) );
  OAI21_X1 U9925 ( .B1(n8403), .B2(n8402), .A(n8401), .ZN(n8405) );
  AOI21_X1 U9926 ( .B1(n8406), .B2(n8405), .A(n8404), .ZN(n8409) );
  OAI21_X1 U9927 ( .B1(n8409), .B2(n8408), .A(n8407), .ZN(n8410) );
  XNOR2_X1 U9928 ( .A(n8410), .B(n9350), .ZN(n8411) );
  NOR4_X1 U9929 ( .A1(n8414), .A2(n8413), .A3(n6068), .A4(n8412), .ZN(n8416)
         );
  OAI21_X1 U9930 ( .B1(n6146), .B2(n8417), .A(P1_B_REG_SCAN_IN), .ZN(n8415) );
  OAI222_X1 U9931 ( .A1(n8421), .A2(n8420), .B1(n8419), .B2(n8418), .C1(n6149), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  OAI22_X1 U9932 ( .A1(n8552), .A2(n8422), .B1(n9800), .B2(n9743), .ZN(n8424)
         );
  NAND2_X1 U9933 ( .A1(n8424), .A2(n8423), .ZN(n8429) );
  INV_X1 U9934 ( .A(n8425), .ZN(n8427) );
  AOI22_X1 U9935 ( .A1(n8427), .A2(P2_REG3_REG_0__SCAN_IN), .B1(n8565), .B2(
        n8426), .ZN(n8428) );
  OAI211_X1 U9936 ( .C1(n7002), .C2(n9750), .A(n8429), .B(n8428), .ZN(P2_U3234) );
  OAI222_X1 U9937 ( .A1(P2_U3152), .A2(n8430), .B1(n4390), .B2(n8432), .C1(
        n8431), .C2(n8459), .ZN(P2_U3328) );
  NAND2_X1 U9938 ( .A1(n8852), .A2(n8830), .ZN(n8435) );
  NAND2_X1 U9939 ( .A1(n8841), .A2(n8435), .ZN(n8826) );
  NAND2_X1 U9940 ( .A1(n8953), .A2(n8573), .ZN(n8436) );
  INV_X1 U9941 ( .A(n8953), .ZN(n8838) );
  NAND2_X1 U9942 ( .A1(n8787), .A2(n8562), .ZN(n8438) );
  INV_X1 U9943 ( .A(n8932), .ZN(n8772) );
  NAND2_X1 U9944 ( .A1(n8755), .A2(n8754), .ZN(n8753) );
  INV_X1 U9945 ( .A(n8927), .ZN(n8759) );
  INV_X1 U9946 ( .A(n8505), .ZN(n8763) );
  INV_X1 U9947 ( .A(n8687), .ZN(n8569) );
  NAND2_X1 U9948 ( .A1(n8682), .A2(n8681), .ZN(n8680) );
  NAND2_X1 U9949 ( .A1(n8680), .A2(n8441), .ZN(n8662) );
  NAND2_X1 U9950 ( .A1(n8662), .A2(n8669), .ZN(n8661) );
  INV_X1 U9951 ( .A(n8442), .ZN(n8695) );
  OR2_X1 U9952 ( .A1(n8902), .A2(n8695), .ZN(n8443) );
  AOI21_X1 U9953 ( .B1(n8898), .B2(n8444), .A(n8656), .ZN(n8899) );
  INV_X1 U9954 ( .A(n8898), .ZN(n8447) );
  AOI22_X1 U9955 ( .A1(n8445), .A2(n8848), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n4388), .ZN(n8446) );
  OAI21_X1 U9956 ( .B1(n8447), .B2(n8851), .A(n8446), .ZN(n8455) );
  OAI21_X1 U9957 ( .B1(n8901), .B2(n8862), .A(n8456), .ZN(P2_U3267) );
  INV_X1 U9958 ( .A(n8457), .ZN(n8458) );
  OAI222_X1 U9959 ( .A1(n8459), .A2(n10145), .B1(n4390), .B2(n8458), .C1(n5684), .C2(P2_U3152), .ZN(P2_U3330) );
  NOR2_X1 U9960 ( .A1(n8461), .A2(n8460), .ZN(n8464) );
  NAND3_X1 U9961 ( .A1(n8462), .A2(n8533), .A3(n8569), .ZN(n8463) );
  OAI21_X1 U9962 ( .B1(n8464), .B2(n9743), .A(n8463), .ZN(n8471) );
  AOI22_X1 U9963 ( .A1(n8695), .A2(n8465), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n8468) );
  INV_X1 U9964 ( .A(n8466), .ZN(n8685) );
  AOI22_X1 U9965 ( .A1(n8569), .A2(n8554), .B1(n8685), .B2(n8511), .ZN(n8467)
         );
  OAI211_X1 U9966 ( .C1(n4704), .C2(n9747), .A(n8468), .B(n8467), .ZN(n8469)
         );
  AOI21_X1 U9967 ( .B1(n8471), .B2(n8470), .A(n8469), .ZN(n8472) );
  INV_X1 U9968 ( .A(n8472), .ZN(P2_U3216) );
  INV_X1 U9969 ( .A(n8473), .ZN(n8474) );
  NAND2_X1 U9970 ( .A1(n8031), .A2(n8474), .ZN(n8476) );
  XNOR2_X1 U9971 ( .A(n8476), .B(n8475), .ZN(n8477) );
  NAND3_X1 U9972 ( .A1(n8477), .A2(n8533), .A3(n8571), .ZN(n8485) );
  INV_X1 U9973 ( .A(n8477), .ZN(n8479) );
  NAND3_X1 U9974 ( .A1(n8479), .A2(n8544), .A3(n8478), .ZN(n8484) );
  OAI22_X1 U9975 ( .A1(n9751), .A2(n8572), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9984), .ZN(n8482) );
  INV_X1 U9976 ( .A(n8757), .ZN(n8480) );
  OAI22_X1 U9977 ( .A1(n9750), .A2(n8505), .B1(n8480), .B2(n9759), .ZN(n8481)
         );
  AOI211_X1 U9978 ( .C1(n8927), .C2(n8565), .A(n8482), .B(n8481), .ZN(n8483)
         );
  NAND3_X1 U9979 ( .A1(n8485), .A2(n8484), .A3(n8483), .ZN(P2_U3218) );
  INV_X1 U9980 ( .A(n8486), .ZN(n8487) );
  AOI21_X1 U9981 ( .B1(n8489), .B2(n8488), .A(n8487), .ZN(n8493) );
  NOR2_X1 U9982 ( .A1(n9759), .A2(n8815), .ZN(n8491) );
  INV_X1 U9983 ( .A(n8496), .ZN(n8790) );
  AOI22_X1 U9984 ( .A1(n8790), .A2(n9774), .B1(n9772), .B2(n8573), .ZN(n8822)
         );
  NAND2_X1 U9985 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8652) );
  OAI21_X1 U9986 ( .B1(n8822), .B2(n8508), .A(n8652), .ZN(n8490) );
  AOI211_X1 U9987 ( .C1(n8949), .C2(n8565), .A(n8491), .B(n8490), .ZN(n8492)
         );
  OAI21_X1 U9988 ( .B1(n8493), .B2(n9743), .A(n8492), .ZN(P2_U3221) );
  XNOR2_X1 U9989 ( .A(n8495), .B(n8494), .ZN(n8500) );
  OAI22_X1 U9990 ( .A1(n9750), .A2(n8572), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10151), .ZN(n8498) );
  OAI22_X1 U9991 ( .A1(n9751), .A2(n8496), .B1(n8784), .B2(n9759), .ZN(n8497)
         );
  AOI211_X1 U9992 ( .C1(n8937), .C2(n8565), .A(n8498), .B(n8497), .ZN(n8499)
         );
  OAI21_X1 U9993 ( .B1(n8500), .B2(n9743), .A(n8499), .ZN(P2_U3225) );
  XNOR2_X1 U9994 ( .A(n8502), .B(n8501), .ZN(n8503) );
  XNOR2_X1 U9995 ( .A(n8504), .B(n8503), .ZN(n8513) );
  OAI22_X1 U9996 ( .A1(n8687), .A2(n8882), .B1(n8505), .B2(n8880), .ZN(n8506)
         );
  INV_X1 U9997 ( .A(n8506), .ZN(n8725) );
  OAI22_X1 U9998 ( .A1(n8725), .A2(n8508), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8507), .ZN(n8510) );
  NOR2_X1 U9999 ( .A1(n4759), .A2(n9747), .ZN(n8509) );
  AOI211_X1 U10000 ( .C1(n8511), .C2(n8730), .A(n8510), .B(n8509), .ZN(n8512)
         );
  OAI21_X1 U10001 ( .B1(n8513), .B2(n9743), .A(n8512), .ZN(P2_U3227) );
  NAND2_X1 U10002 ( .A1(n8515), .A2(n8514), .ZN(n8521) );
  OAI22_X1 U10003 ( .A1(n8519), .A2(n8518), .B1(n8517), .B2(n8516), .ZN(n8520)
         );
  XOR2_X1 U10004 ( .A(n8521), .B(n8520), .Z(n8532) );
  NAND2_X1 U10005 ( .A1(n8522), .A2(n9818), .ZN(n9486) );
  INV_X1 U10006 ( .A(n9486), .ZN(n8530) );
  NAND2_X1 U10007 ( .A1(n8524), .A2(n8523), .ZN(n8526) );
  NOR2_X1 U10008 ( .A1(n9982), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8595) );
  INV_X1 U10009 ( .A(n8595), .ZN(n8525) );
  OAI211_X1 U10010 ( .C1(n9759), .C2(n8527), .A(n8526), .B(n8525), .ZN(n8528)
         );
  AOI21_X1 U10011 ( .B1(n8530), .B2(n8529), .A(n8528), .ZN(n8531) );
  OAI21_X1 U10012 ( .B1(n8532), .B2(n9743), .A(n8531), .ZN(P2_U3228) );
  NAND2_X1 U10013 ( .A1(n8763), .A2(n8533), .ZN(n8537) );
  OR2_X1 U10014 ( .A1(n8534), .A2(n9743), .ZN(n8536) );
  MUX2_X1 U10015 ( .A(n8537), .B(n8536), .S(n8535), .Z(n8541) );
  OAI22_X1 U10016 ( .A1(n8747), .A2(n9750), .B1(n9759), .B2(n8738), .ZN(n8539)
         );
  OAI22_X1 U10017 ( .A1(n9751), .A2(n8746), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10109), .ZN(n8538) );
  NOR2_X1 U10018 ( .A1(n8539), .A2(n8538), .ZN(n8540) );
  OAI211_X1 U10019 ( .C1(n4761), .C2(n9747), .A(n8541), .B(n8540), .ZN(
        P2_U3231) );
  OAI21_X1 U10020 ( .B1(n8553), .B2(n8543), .A(n8542), .ZN(n8545) );
  NAND2_X1 U10021 ( .A1(n8545), .A2(n8544), .ZN(n8558) );
  OAI22_X1 U10022 ( .A1(n9750), .A2(n8547), .B1(n9759), .B2(n8546), .ZN(n8548)
         );
  AOI211_X1 U10023 ( .C1(n8565), .C2(n8550), .A(n8549), .B(n8548), .ZN(n8557)
         );
  NOR3_X1 U10024 ( .A1(n8553), .A2(n8552), .A3(n8551), .ZN(n8555) );
  OAI21_X1 U10025 ( .B1(n8555), .B2(n8554), .A(n8585), .ZN(n8556) );
  NAND3_X1 U10026 ( .A1(n8558), .A2(n8557), .A3(n8556), .ZN(P2_U3232) );
  XNOR2_X1 U10027 ( .A(n8560), .B(n8559), .ZN(n8567) );
  OAI22_X1 U10028 ( .A1(n9750), .A2(n8562), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8561), .ZN(n8564) );
  OAI22_X1 U10029 ( .A1(n9751), .A2(n8831), .B1(n8799), .B2(n9759), .ZN(n8563)
         );
  AOI211_X1 U10030 ( .C1(n8942), .C2(n8565), .A(n8564), .B(n8563), .ZN(n8566)
         );
  OAI21_X1 U10031 ( .B1(n8567), .B2(n9743), .A(n8566), .ZN(P2_U3235) );
  MUX2_X1 U10032 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8568), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U10033 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8671), .S(P2_U3966), .Z(
        P2_U3581) );
  MUX2_X1 U10034 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8695), .S(P2_U3966), .Z(
        P2_U3580) );
  MUX2_X1 U10035 ( .A(n8672), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8586), .Z(
        P2_U3579) );
  MUX2_X1 U10036 ( .A(n8569), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8586), .Z(
        P2_U3578) );
  MUX2_X1 U10037 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8570), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U10038 ( .A(n8763), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8586), .Z(
        P2_U3576) );
  MUX2_X1 U10039 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8571), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U10040 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8439), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U10041 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8807), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U10042 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8790), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U10043 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8806), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U10044 ( .A(n8573), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8586), .Z(
        P2_U3570) );
  MUX2_X1 U10045 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8574), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U10046 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8575), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10047 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8576), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10048 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8577), .S(P2_U3966), .Z(
        P2_U3566) );
  INV_X1 U10049 ( .A(n8881), .ZN(n8578) );
  MUX2_X1 U10050 ( .A(n8578), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8586), .Z(
        P2_U3565) );
  MUX2_X1 U10051 ( .A(n8579), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8586), .Z(
        P2_U3564) );
  MUX2_X1 U10052 ( .A(n8580), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8586), .Z(
        P2_U3563) );
  MUX2_X1 U10053 ( .A(n8581), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8586), .Z(
        P2_U3562) );
  MUX2_X1 U10054 ( .A(n8582), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8586), .Z(
        P2_U3561) );
  MUX2_X1 U10055 ( .A(n8583), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8586), .Z(
        P2_U3560) );
  MUX2_X1 U10056 ( .A(n9775), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8586), .Z(
        P2_U3559) );
  MUX2_X1 U10057 ( .A(n9748), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8586), .Z(
        P2_U3558) );
  MUX2_X1 U10058 ( .A(n9773), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8586), .Z(
        P2_U3557) );
  MUX2_X1 U10059 ( .A(n8584), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8586), .Z(
        P2_U3556) );
  MUX2_X1 U10060 ( .A(n8585), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8586), .Z(
        P2_U3555) );
  MUX2_X1 U10061 ( .A(n6158), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8586), .Z(
        P2_U3554) );
  MUX2_X1 U10062 ( .A(n6157), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8586), .Z(
        P2_U3553) );
  MUX2_X1 U10063 ( .A(n6209), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8586), .Z(
        P2_U3552) );
  NOR2_X1 U10064 ( .A1(n8588), .A2(n8587), .ZN(n8590) );
  NOR2_X1 U10065 ( .A1(n8590), .A2(n8589), .ZN(n8593) );
  MUX2_X1 U10066 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8591), .S(n8613), .Z(n8592) );
  NAND2_X1 U10067 ( .A1(n8592), .A2(n8593), .ZN(n8614) );
  OAI21_X1 U10068 ( .B1(n8593), .B2(n8592), .A(n8614), .ZN(n8594) );
  NAND2_X1 U10069 ( .A1(n8594), .A2(n9763), .ZN(n8606) );
  AOI21_X1 U10070 ( .B1(n9766), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8595), .ZN(
        n8605) );
  NOR2_X1 U10071 ( .A1(n8597), .A2(n8596), .ZN(n8599) );
  NOR2_X1 U10072 ( .A1(n8599), .A2(n8598), .ZN(n8602) );
  MUX2_X1 U10073 ( .A(n7989), .B(P2_REG2_REG_16__SCAN_IN), .S(n8613), .Z(n8600) );
  INV_X1 U10074 ( .A(n8600), .ZN(n8601) );
  NAND2_X1 U10075 ( .A1(n8601), .A2(n8602), .ZN(n8607) );
  OAI211_X1 U10076 ( .C1(n8602), .C2(n8601), .A(n9764), .B(n8607), .ZN(n8604)
         );
  NAND2_X1 U10077 ( .A1(n9472), .A2(n8613), .ZN(n8603) );
  NAND4_X1 U10078 ( .A1(n8606), .A2(n8605), .A3(n8604), .A4(n8603), .ZN(
        P2_U3261) );
  NAND2_X1 U10079 ( .A1(n8613), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8608) );
  NAND2_X1 U10080 ( .A1(n8608), .A2(n8607), .ZN(n8610) );
  XOR2_X1 U10081 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n8630), .Z(n8609) );
  NAND2_X1 U10082 ( .A1(n8609), .A2(n8610), .ZN(n8624) );
  OAI211_X1 U10083 ( .C1(n8610), .C2(n8609), .A(n9764), .B(n8624), .ZN(n8622)
         );
  NOR2_X1 U10084 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5425), .ZN(n8611) );
  AOI21_X1 U10085 ( .B1(n9766), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8611), .ZN(
        n8621) );
  OR2_X1 U10086 ( .A1(n9760), .A2(n8612), .ZN(n8620) );
  XNOR2_X1 U10087 ( .A(n8630), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8617) );
  OR2_X1 U10088 ( .A1(n8613), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8615) );
  NAND2_X1 U10089 ( .A1(n8615), .A2(n8614), .ZN(n8616) );
  NOR2_X1 U10090 ( .A1(n8617), .A2(n8616), .ZN(n8629) );
  AOI21_X1 U10091 ( .B1(n8617), .B2(n8616), .A(n8629), .ZN(n8618) );
  NAND2_X1 U10092 ( .A1(n9763), .A2(n8618), .ZN(n8619) );
  NAND4_X1 U10093 ( .A1(n8622), .A2(n8621), .A3(n8620), .A4(n8619), .ZN(
        P2_U3262) );
  OAI21_X1 U10094 ( .B1(n8655), .B2(n10201), .A(n8623), .ZN(n8636) );
  NAND2_X1 U10095 ( .A1(n8630), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8625) );
  NAND2_X1 U10096 ( .A1(n8625), .A2(n8624), .ZN(n8626) );
  NOR2_X1 U10097 ( .A1(n8626), .A2(n8643), .ZN(n8639) );
  AOI21_X1 U10098 ( .B1(n8643), .B2(n8626), .A(n8639), .ZN(n8627) );
  INV_X1 U10099 ( .A(n8627), .ZN(n8628) );
  NOR2_X1 U10100 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8628), .ZN(n8638) );
  AOI21_X1 U10101 ( .B1(n8628), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8638), .ZN(
        n8634) );
  XNOR2_X1 U10102 ( .A(n8643), .B(n8631), .ZN(n8642) );
  XOR2_X1 U10103 ( .A(n8641), .B(n8642), .Z(n8632) );
  OAI22_X1 U10104 ( .A1(n8634), .A2(n8633), .B1(n8632), .B2(n9761), .ZN(n8635)
         );
  AOI211_X1 U10105 ( .C1(n8643), .C2(n9472), .A(n8636), .B(n8635), .ZN(n8637)
         );
  INV_X1 U10106 ( .A(n8637), .ZN(P2_U3263) );
  INV_X1 U10107 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8654) );
  NOR2_X1 U10108 ( .A1(n8639), .A2(n8638), .ZN(n8640) );
  XOR2_X1 U10109 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8640), .Z(n8648) );
  INV_X1 U10110 ( .A(n8648), .ZN(n8646) );
  OR2_X1 U10111 ( .A1(n8643), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8644) );
  OAI21_X1 U10112 ( .B1(n8647), .B2(n9761), .A(n9760), .ZN(n8645) );
  AOI21_X1 U10113 ( .B1(n8646), .B2(n9764), .A(n8645), .ZN(n8651) );
  AOI22_X1 U10114 ( .A1(n8648), .A2(n9764), .B1(n8647), .B2(n9763), .ZN(n8650)
         );
  MUX2_X1 U10115 ( .A(n8651), .B(n8650), .S(n8649), .Z(n8653) );
  OAI211_X1 U10116 ( .C1(n8655), .C2(n8654), .A(n8653), .B(n8652), .ZN(
        P2_U3264) );
  INV_X1 U10117 ( .A(n8656), .ZN(n8657) );
  NAND2_X1 U10118 ( .A1(n4893), .A2(n8657), .ZN(n8894) );
  NAND3_X1 U10119 ( .A1(n8894), .A2(n8834), .A3(n8893), .ZN(n8660) );
  AOI21_X1 U10120 ( .B1(n4388), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8658), .ZN(
        n8659) );
  OAI211_X1 U10121 ( .C1(n8897), .C2(n8851), .A(n8660), .B(n8659), .ZN(
        P2_U3266) );
  OAI21_X1 U10122 ( .B1(n8662), .B2(n8669), .A(n8661), .ZN(n8663) );
  INV_X1 U10123 ( .A(n8663), .ZN(n8906) );
  INV_X1 U10124 ( .A(n8684), .ZN(n8665) );
  INV_X1 U10125 ( .A(n8444), .ZN(n8664) );
  AOI21_X1 U10126 ( .B1(n8902), .B2(n8665), .A(n8664), .ZN(n8903) );
  AOI22_X1 U10127 ( .A1(n8666), .A2(n8848), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n4388), .ZN(n8667) );
  OAI21_X1 U10128 ( .B1(n8668), .B2(n8851), .A(n8667), .ZN(n8678) );
  XNOR2_X1 U10129 ( .A(n8670), .B(n8669), .ZN(n8676) );
  NAND2_X1 U10130 ( .A1(n8672), .A2(n9772), .ZN(n8673) );
  AOI211_X1 U10131 ( .C1(n8903), .C2(n8834), .A(n8678), .B(n8677), .ZN(n8679)
         );
  OAI21_X1 U10132 ( .B1(n8906), .B2(n8862), .A(n8679), .ZN(P2_U3268) );
  OAI21_X1 U10133 ( .B1(n8682), .B2(n8681), .A(n8680), .ZN(n8683) );
  INV_X1 U10134 ( .A(n8683), .ZN(n8911) );
  AOI21_X1 U10135 ( .B1(n8907), .B2(n8711), .A(n8684), .ZN(n8908) );
  AOI22_X1 U10136 ( .A1(n8685), .A2(n8848), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n4388), .ZN(n8686) );
  OAI21_X1 U10137 ( .B1(n4704), .B2(n8851), .A(n8686), .ZN(n8697) );
  NOR2_X1 U10138 ( .A1(n8687), .A2(n8880), .ZN(n8694) );
  INV_X1 U10139 ( .A(n8688), .ZN(n8692) );
  AOI21_X1 U10140 ( .B1(n8690), .B2(n8689), .A(n4663), .ZN(n8691) );
  NOR3_X1 U10141 ( .A1(n8692), .A2(n8691), .A3(n8877), .ZN(n8693) );
  NOR2_X1 U10142 ( .A1(n8910), .A2(n4388), .ZN(n8696) );
  AOI211_X1 U10143 ( .C1(n8908), .C2(n8834), .A(n8697), .B(n8696), .ZN(n8698)
         );
  OAI21_X1 U10144 ( .B1(n8911), .B2(n8862), .A(n8698), .ZN(P2_U3269) );
  OAI21_X1 U10145 ( .B1(n8700), .B2(n8704), .A(n8699), .ZN(n8701) );
  INV_X1 U10146 ( .A(n8701), .ZN(n8916) );
  AOI22_X1 U10147 ( .A1(n8914), .A2(n8872), .B1(n4388), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8718) );
  NAND2_X1 U10148 ( .A1(n8702), .A2(n8703), .ZN(n8705) );
  NOR2_X1 U10149 ( .A1(n8747), .A2(n8880), .ZN(n8708) );
  INV_X1 U10150 ( .A(n8711), .ZN(n8712) );
  AOI211_X1 U10151 ( .C1(n8914), .C2(n8727), .A(n9853), .B(n8712), .ZN(n8913)
         );
  INV_X1 U10152 ( .A(n8913), .ZN(n8715) );
  OAI22_X1 U10153 ( .A1(n8715), .A2(n4385), .B1(n9778), .B2(n8713), .ZN(n8716)
         );
  OAI21_X1 U10154 ( .B1(n8912), .B2(n8716), .A(n8870), .ZN(n8717) );
  OAI211_X1 U10155 ( .C1(n8916), .C2(n8862), .A(n8718), .B(n8717), .ZN(
        P2_U3270) );
  OAI21_X1 U10156 ( .B1(n8721), .B2(n8720), .A(n8719), .ZN(n8722) );
  INV_X1 U10157 ( .A(n8722), .ZN(n8921) );
  OAI211_X1 U10158 ( .C1(n8724), .C2(n8723), .A(n8702), .B(n9777), .ZN(n8726)
         );
  NAND2_X1 U10159 ( .A1(n8726), .A2(n8725), .ZN(n8917) );
  INV_X1 U10160 ( .A(n8736), .ZN(n8729) );
  INV_X1 U10161 ( .A(n8727), .ZN(n8728) );
  AOI211_X1 U10162 ( .C1(n8919), .C2(n8729), .A(n9853), .B(n8728), .ZN(n8918)
         );
  NAND2_X1 U10163 ( .A1(n8918), .A2(n8854), .ZN(n8732) );
  AOI22_X1 U10164 ( .A1(n4388), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8730), .B2(
        n8848), .ZN(n8731) );
  OAI211_X1 U10165 ( .C1(n4759), .C2(n8851), .A(n8732), .B(n8731), .ZN(n8733)
         );
  AOI21_X1 U10166 ( .B1(n8917), .B2(n8870), .A(n8733), .ZN(n8734) );
  OAI21_X1 U10167 ( .B1(n8921), .B2(n8862), .A(n8734), .ZN(P2_U3271) );
  XOR2_X1 U10168 ( .A(n8742), .B(n8735), .Z(n8926) );
  INV_X1 U10169 ( .A(n8756), .ZN(n8737) );
  AOI21_X1 U10170 ( .B1(n8922), .B2(n8737), .A(n8736), .ZN(n8923) );
  INV_X1 U10171 ( .A(n8738), .ZN(n8739) );
  AOI22_X1 U10172 ( .A1(n4388), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8739), .B2(
        n8848), .ZN(n8740) );
  OAI21_X1 U10173 ( .B1(n4761), .B2(n8851), .A(n8740), .ZN(n8751) );
  INV_X1 U10174 ( .A(n8741), .ZN(n8745) );
  AOI21_X1 U10175 ( .B1(n8760), .B2(n8743), .A(n8742), .ZN(n8744) );
  NOR3_X1 U10176 ( .A1(n8745), .A2(n8744), .A3(n8877), .ZN(n8749) );
  OAI22_X1 U10177 ( .A1(n8747), .A2(n8882), .B1(n8746), .B2(n8880), .ZN(n8748)
         );
  NOR2_X1 U10178 ( .A1(n8749), .A2(n8748), .ZN(n8925) );
  NOR2_X1 U10179 ( .A1(n8925), .A2(n4388), .ZN(n8750) );
  AOI211_X1 U10180 ( .C1(n8923), .C2(n8834), .A(n8751), .B(n8750), .ZN(n8752)
         );
  OAI21_X1 U10181 ( .B1(n8862), .B2(n8926), .A(n8752), .ZN(P2_U3272) );
  OAI21_X1 U10182 ( .B1(n8755), .B2(n8754), .A(n8753), .ZN(n8931) );
  AOI21_X1 U10183 ( .B1(n8927), .B2(n8769), .A(n8756), .ZN(n8928) );
  AOI22_X1 U10184 ( .A1(n4388), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8757), .B2(
        n8848), .ZN(n8758) );
  OAI21_X1 U10185 ( .B1(n8759), .B2(n8851), .A(n8758), .ZN(n8766) );
  OAI21_X1 U10186 ( .B1(n8762), .B2(n8761), .A(n8760), .ZN(n8764) );
  AOI222_X1 U10187 ( .A1(n9777), .A2(n8764), .B1(n8439), .B2(n9772), .C1(n8763), .C2(n9774), .ZN(n8930) );
  NOR2_X1 U10188 ( .A1(n8930), .A2(n4388), .ZN(n8765) );
  AOI211_X1 U10189 ( .C1(n8928), .C2(n8834), .A(n8766), .B(n8765), .ZN(n8767)
         );
  OAI21_X1 U10190 ( .B1(n8862), .B2(n8931), .A(n8767), .ZN(P2_U3273) );
  XOR2_X1 U10191 ( .A(n8775), .B(n8768), .Z(n8936) );
  AOI21_X1 U10192 ( .B1(n8932), .B2(n8782), .A(n4697), .ZN(n8933) );
  AOI22_X1 U10193 ( .A1(n4388), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8770), .B2(
        n8848), .ZN(n8771) );
  OAI21_X1 U10194 ( .B1(n8772), .B2(n8851), .A(n8771), .ZN(n8779) );
  AOI211_X1 U10195 ( .C1(n8775), .C2(n8774), .A(n8877), .B(n8773), .ZN(n8777)
         );
  NOR2_X1 U10196 ( .A1(n8777), .A2(n8776), .ZN(n8935) );
  NOR2_X1 U10197 ( .A1(n8935), .A2(n4388), .ZN(n8778) );
  AOI211_X1 U10198 ( .C1(n8933), .C2(n8834), .A(n8779), .B(n8778), .ZN(n8780)
         );
  OAI21_X1 U10199 ( .B1(n8862), .B2(n8936), .A(n8780), .ZN(P2_U3274) );
  XNOR2_X1 U10200 ( .A(n8781), .B(n8788), .ZN(n8941) );
  INV_X1 U10201 ( .A(n8797), .ZN(n8783) );
  AOI21_X1 U10202 ( .B1(n8937), .B2(n8783), .A(n4694), .ZN(n8938) );
  INV_X1 U10203 ( .A(n8784), .ZN(n8785) );
  AOI22_X1 U10204 ( .A1(n4388), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8785), .B2(
        n8848), .ZN(n8786) );
  OAI21_X1 U10205 ( .B1(n8787), .B2(n8851), .A(n8786), .ZN(n8793) );
  XNOR2_X1 U10206 ( .A(n8789), .B(n8788), .ZN(n8791) );
  AOI222_X1 U10207 ( .A1(n9777), .A2(n8791), .B1(n8439), .B2(n9774), .C1(n8790), .C2(n9772), .ZN(n8940) );
  NOR2_X1 U10208 ( .A1(n8940), .A2(n4388), .ZN(n8792) );
  AOI211_X1 U10209 ( .C1(n8938), .C2(n8834), .A(n8793), .B(n8792), .ZN(n8794)
         );
  OAI21_X1 U10210 ( .B1(n8941), .B2(n8862), .A(n8794), .ZN(P2_U3275) );
  OAI21_X1 U10211 ( .B1(n8796), .B2(n8804), .A(n8795), .ZN(n8946) );
  INV_X1 U10212 ( .A(n8814), .ZN(n8798) );
  AOI21_X1 U10213 ( .B1(n8942), .B2(n8798), .A(n8797), .ZN(n8943) );
  INV_X1 U10214 ( .A(n8799), .ZN(n8800) );
  AOI22_X1 U10215 ( .A1(n4388), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8800), .B2(
        n8848), .ZN(n8801) );
  OAI21_X1 U10216 ( .B1(n8802), .B2(n8851), .A(n8801), .ZN(n8810) );
  NOR2_X1 U10217 ( .A1(n8819), .A2(n4652), .ZN(n8805) );
  XNOR2_X1 U10218 ( .A(n8805), .B(n8804), .ZN(n8808) );
  AOI222_X1 U10219 ( .A1(n9777), .A2(n8808), .B1(n8807), .B2(n9774), .C1(n8806), .C2(n9772), .ZN(n8945) );
  NOR2_X1 U10220 ( .A1(n8945), .A2(n4388), .ZN(n8809) );
  AOI211_X1 U10221 ( .C1(n8943), .C2(n8834), .A(n8810), .B(n8809), .ZN(n8811)
         );
  OAI21_X1 U10222 ( .B1(n8862), .B2(n8946), .A(n8811), .ZN(P2_U3276) );
  OAI21_X1 U10223 ( .B1(n8813), .B2(n8820), .A(n8812), .ZN(n8951) );
  AOI211_X1 U10224 ( .C1(n8949), .C2(n8832), .A(n9853), .B(n8814), .ZN(n8948)
         );
  NOR2_X1 U10225 ( .A1(n4696), .A2(n8851), .ZN(n8818) );
  OAI22_X1 U10226 ( .A1(n8870), .A2(n8816), .B1(n8815), .B2(n9778), .ZN(n8817)
         );
  AOI211_X1 U10227 ( .C1(n8948), .C2(n8854), .A(n8818), .B(n8817), .ZN(n8825)
         );
  AOI21_X1 U10228 ( .B1(n8821), .B2(n8820), .A(n8819), .ZN(n8823) );
  OAI21_X1 U10229 ( .B1(n8823), .B2(n8877), .A(n8822), .ZN(n8947) );
  NAND2_X1 U10230 ( .A1(n8947), .A2(n8870), .ZN(n8824) );
  OAI211_X1 U10231 ( .C1(n8951), .C2(n8862), .A(n8825), .B(n8824), .ZN(
        P2_U3277) );
  XOR2_X1 U10232 ( .A(n8826), .B(n8827), .Z(n8957) );
  AOI21_X1 U10233 ( .B1(n8828), .B2(n8827), .A(n4465), .ZN(n8829) );
  OAI222_X1 U10234 ( .A1(n8882), .A2(n8831), .B1(n8880), .B2(n8830), .C1(n8877), .C2(n8829), .ZN(n8952) );
  INV_X1 U10235 ( .A(n8832), .ZN(n8833) );
  AOI21_X1 U10236 ( .B1(n8953), .B2(n8844), .A(n8833), .ZN(n8954) );
  NAND2_X1 U10237 ( .A1(n8954), .A2(n8834), .ZN(n8837) );
  AOI22_X1 U10238 ( .A1(n4388), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8835), .B2(
        n8848), .ZN(n8836) );
  OAI211_X1 U10239 ( .C1(n8838), .C2(n8851), .A(n8837), .B(n8836), .ZN(n8839)
         );
  AOI21_X1 U10240 ( .B1(n8952), .B2(n8870), .A(n8839), .ZN(n8840) );
  OAI21_X1 U10241 ( .B1(n8957), .B2(n8862), .A(n8840), .ZN(P2_U3278) );
  OAI21_X1 U10242 ( .B1(n4468), .B2(n8855), .A(n8841), .ZN(n8842) );
  INV_X1 U10243 ( .A(n8842), .ZN(n8962) );
  INV_X1 U10244 ( .A(n8843), .ZN(n8846) );
  INV_X1 U10245 ( .A(n8844), .ZN(n8845) );
  AOI211_X1 U10246 ( .C1(n8960), .C2(n8846), .A(n9853), .B(n8845), .ZN(n8959)
         );
  INV_X1 U10247 ( .A(n8847), .ZN(n8849) );
  AOI22_X1 U10248 ( .A1(n4388), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8849), .B2(
        n8848), .ZN(n8850) );
  OAI21_X1 U10249 ( .B1(n8852), .B2(n8851), .A(n8850), .ZN(n8853) );
  AOI21_X1 U10250 ( .B1(n8959), .B2(n8854), .A(n8853), .ZN(n8861) );
  XNOR2_X1 U10251 ( .A(n8856), .B(n8855), .ZN(n8857) );
  OAI222_X1 U10252 ( .A1(n8882), .A2(n8859), .B1(n8880), .B2(n8858), .C1(n8857), .C2(n8877), .ZN(n8958) );
  NAND2_X1 U10253 ( .A1(n8958), .A2(n8870), .ZN(n8860) );
  OAI211_X1 U10254 ( .C1(n8962), .C2(n8862), .A(n8861), .B(n8860), .ZN(
        P2_U3279) );
  XNOR2_X1 U10255 ( .A(n8864), .B(n8863), .ZN(n9496) );
  NAND2_X1 U10256 ( .A1(n8865), .A2(n9491), .ZN(n8866) );
  NAND2_X1 U10257 ( .A1(n8867), .A2(n8866), .ZN(n9494) );
  OAI22_X1 U10258 ( .A1(n8870), .A2(n8869), .B1(n8868), .B2(n9778), .ZN(n8871)
         );
  AOI21_X1 U10259 ( .B1(n9491), .B2(n8872), .A(n8871), .ZN(n8873) );
  OAI21_X1 U10260 ( .B1(n9494), .B2(n8874), .A(n8873), .ZN(n8888) );
  NAND2_X1 U10261 ( .A1(n8876), .A2(n8875), .ZN(n8879) );
  AOI21_X1 U10262 ( .B1(n8879), .B2(n8878), .A(n8877), .ZN(n8886) );
  OAI22_X1 U10263 ( .A1(n8883), .A2(n8882), .B1(n8881), .B2(n8880), .ZN(n8884)
         );
  AOI21_X1 U10264 ( .B1(n8886), .B2(n8885), .A(n8884), .ZN(n9493) );
  NOR2_X1 U10265 ( .A1(n9493), .A2(n4388), .ZN(n8887) );
  AOI211_X1 U10266 ( .C1(n9496), .C2(n9787), .A(n8888), .B(n8887), .ZN(n8889)
         );
  INV_X1 U10267 ( .A(n8889), .ZN(P2_U3282) );
  NAND2_X1 U10268 ( .A1(n8890), .A2(n9818), .ZN(n8891) );
  OAI211_X1 U10269 ( .C1(n8892), .C2(n9853), .A(n8891), .B(n8895), .ZN(n8980)
         );
  MUX2_X1 U10270 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8980), .S(n9875), .Z(
        P2_U3551) );
  NAND3_X1 U10271 ( .A1(n8894), .A2(n9819), .A3(n8893), .ZN(n8896) );
  OAI211_X1 U10272 ( .C1(n8897), .C2(n9851), .A(n8896), .B(n8895), .ZN(n8981)
         );
  INV_X2 U10273 ( .A(n9873), .ZN(n9875) );
  MUX2_X1 U10274 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8981), .S(n9875), .Z(
        P2_U3550) );
  AOI22_X1 U10275 ( .A1(n8903), .A2(n9819), .B1(n9818), .B2(n8902), .ZN(n8904)
         );
  OAI211_X1 U10276 ( .C1(n8906), .C2(n9485), .A(n8905), .B(n8904), .ZN(n8983)
         );
  MUX2_X1 U10277 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8983), .S(n9875), .Z(
        P2_U3548) );
  AOI22_X1 U10278 ( .A1(n8908), .A2(n9819), .B1(n9818), .B2(n8907), .ZN(n8909)
         );
  OAI211_X1 U10279 ( .C1(n8911), .C2(n9485), .A(n8910), .B(n8909), .ZN(n8984)
         );
  MUX2_X1 U10280 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8984), .S(n9875), .Z(
        P2_U3547) );
  AOI211_X1 U10281 ( .C1(n9818), .C2(n8914), .A(n8913), .B(n8912), .ZN(n8915)
         );
  OAI21_X1 U10282 ( .B1(n9485), .B2(n8916), .A(n8915), .ZN(n8985) );
  MUX2_X1 U10283 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8985), .S(n9875), .Z(
        P2_U3546) );
  AOI211_X1 U10284 ( .C1(n9818), .C2(n8919), .A(n8918), .B(n8917), .ZN(n8920)
         );
  OAI21_X1 U10285 ( .B1(n8921), .B2(n9485), .A(n8920), .ZN(n8986) );
  MUX2_X1 U10286 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8986), .S(n9875), .Z(
        P2_U3545) );
  AOI22_X1 U10287 ( .A1(n8923), .A2(n9819), .B1(n9818), .B2(n8922), .ZN(n8924)
         );
  OAI211_X1 U10288 ( .C1(n8926), .C2(n9485), .A(n8925), .B(n8924), .ZN(n8987)
         );
  MUX2_X1 U10289 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8987), .S(n9875), .Z(
        P2_U3544) );
  AOI22_X1 U10290 ( .A1(n8928), .A2(n9819), .B1(n9818), .B2(n8927), .ZN(n8929)
         );
  OAI211_X1 U10291 ( .C1(n8931), .C2(n9485), .A(n8930), .B(n8929), .ZN(n8988)
         );
  MUX2_X1 U10292 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8988), .S(n9875), .Z(
        P2_U3543) );
  AOI22_X1 U10293 ( .A1(n8933), .A2(n9819), .B1(n9818), .B2(n8932), .ZN(n8934)
         );
  OAI211_X1 U10294 ( .C1(n8936), .C2(n9485), .A(n8935), .B(n8934), .ZN(n8989)
         );
  MUX2_X1 U10295 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8989), .S(n9875), .Z(
        P2_U3542) );
  AOI22_X1 U10296 ( .A1(n8938), .A2(n9819), .B1(n9818), .B2(n8937), .ZN(n8939)
         );
  OAI211_X1 U10297 ( .C1(n8941), .C2(n9485), .A(n8940), .B(n8939), .ZN(n8990)
         );
  MUX2_X1 U10298 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8990), .S(n9875), .Z(
        P2_U3541) );
  AOI22_X1 U10299 ( .A1(n8943), .A2(n9819), .B1(n9818), .B2(n8942), .ZN(n8944)
         );
  OAI211_X1 U10300 ( .C1(n8946), .C2(n9485), .A(n8945), .B(n8944), .ZN(n8991)
         );
  MUX2_X1 U10301 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8991), .S(n9875), .Z(
        P2_U3540) );
  AOI211_X1 U10302 ( .C1(n9818), .C2(n8949), .A(n8948), .B(n8947), .ZN(n8950)
         );
  OAI21_X1 U10303 ( .B1(n9485), .B2(n8951), .A(n8950), .ZN(n8992) );
  MUX2_X1 U10304 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8992), .S(n9875), .Z(
        P2_U3539) );
  INV_X1 U10305 ( .A(n8952), .ZN(n8956) );
  AOI22_X1 U10306 ( .A1(n8954), .A2(n9819), .B1(n9818), .B2(n8953), .ZN(n8955)
         );
  OAI211_X1 U10307 ( .C1(n8957), .C2(n9485), .A(n8956), .B(n8955), .ZN(n8993)
         );
  MUX2_X1 U10308 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8993), .S(n9875), .Z(
        P2_U3538) );
  AOI211_X1 U10309 ( .C1(n9818), .C2(n8960), .A(n8959), .B(n8958), .ZN(n8961)
         );
  OAI21_X1 U10310 ( .B1(n8962), .B2(n9485), .A(n8961), .ZN(n8994) );
  MUX2_X1 U10311 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8994), .S(n9875), .Z(
        P2_U3537) );
  INV_X1 U10312 ( .A(n8963), .ZN(n8968) );
  AOI22_X1 U10313 ( .A1(n8965), .A2(n9819), .B1(n9818), .B2(n8964), .ZN(n8966)
         );
  OAI211_X1 U10314 ( .C1(n8968), .C2(n9485), .A(n8967), .B(n8966), .ZN(n8995)
         );
  MUX2_X1 U10315 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8995), .S(n9875), .Z(
        P2_U3535) );
  AOI22_X1 U10316 ( .A1(n8969), .A2(n9819), .B1(n9818), .B2(n6166), .ZN(n8970)
         );
  OAI21_X1 U10317 ( .B1(n8971), .B2(n9824), .A(n8970), .ZN(n8972) );
  NOR2_X1 U10318 ( .A1(n8973), .A2(n8972), .ZN(n8996) );
  MUX2_X1 U10319 ( .A(n5158), .B(n8996), .S(n9875), .Z(n8974) );
  INV_X1 U10320 ( .A(n8974), .ZN(P2_U3533) );
  AOI22_X1 U10321 ( .A1(n8976), .A2(n9819), .B1(n9818), .B2(n8975), .ZN(n8977)
         );
  OAI211_X1 U10322 ( .C1(n9485), .C2(n8979), .A(n8978), .B(n8977), .ZN(n8999)
         );
  MUX2_X1 U10323 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n8999), .S(n9875), .Z(
        P2_U3531) );
  MUX2_X1 U10324 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8980), .S(n9861), .Z(
        P2_U3519) );
  INV_X2 U10325 ( .A(n9859), .ZN(n9861) );
  MUX2_X1 U10326 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8981), .S(n9861), .Z(
        P2_U3518) );
  MUX2_X1 U10327 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8983), .S(n9861), .Z(
        P2_U3516) );
  MUX2_X1 U10328 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8984), .S(n9861), .Z(
        P2_U3515) );
  MUX2_X1 U10329 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8985), .S(n9861), .Z(
        P2_U3514) );
  MUX2_X1 U10330 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8986), .S(n9861), .Z(
        P2_U3513) );
  MUX2_X1 U10331 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8987), .S(n9861), .Z(
        P2_U3512) );
  MUX2_X1 U10332 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8988), .S(n9861), .Z(
        P2_U3511) );
  MUX2_X1 U10333 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8989), .S(n9861), .Z(
        P2_U3510) );
  MUX2_X1 U10334 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8990), .S(n9861), .Z(
        P2_U3509) );
  MUX2_X1 U10335 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8991), .S(n9861), .Z(
        P2_U3508) );
  MUX2_X1 U10336 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8992), .S(n9861), .Z(
        P2_U3507) );
  MUX2_X1 U10337 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8993), .S(n9861), .Z(
        P2_U3505) );
  MUX2_X1 U10338 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8994), .S(n9861), .Z(
        P2_U3502) );
  MUX2_X1 U10339 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8995), .S(n9861), .Z(
        P2_U3496) );
  INV_X1 U10340 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8997) );
  MUX2_X1 U10341 ( .A(n8997), .B(n8996), .S(n9861), .Z(n8998) );
  INV_X1 U10342 ( .A(n8998), .ZN(P2_U3490) );
  MUX2_X1 U10343 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n8999), .S(n9861), .Z(
        P2_U3484) );
  MUX2_X1 U10344 ( .A(n9000), .B(n9765), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10345 ( .A(n9003), .B(n9002), .ZN(n9004) );
  XNOR2_X1 U10346 ( .A(n9001), .B(n9004), .ZN(n9009) );
  OAI22_X1 U10347 ( .A1(n9110), .A2(n9228), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9005), .ZN(n9007) );
  OAI22_X1 U10348 ( .A1(n9108), .A2(n9222), .B1(n9229), .B2(n9106), .ZN(n9006)
         );
  AOI211_X1 U10349 ( .C1(n9388), .C2(n9100), .A(n9007), .B(n9006), .ZN(n9008)
         );
  OAI21_X1 U10350 ( .B1(n9009), .B2(n9095), .A(n9008), .ZN(P1_U3212) );
  NAND2_X1 U10351 ( .A1(n4920), .A2(n9010), .ZN(n9012) );
  XNOR2_X1 U10352 ( .A(n9012), .B(n9011), .ZN(n9017) );
  OAI22_X1 U10353 ( .A1(n9106), .A2(n9034), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9013), .ZN(n9015) );
  OAI22_X1 U10354 ( .A1(n9108), .A2(n9280), .B1(n9319), .B2(n9110), .ZN(n9014)
         );
  AOI211_X1 U10355 ( .C1(n9408), .C2(n9100), .A(n9015), .B(n9014), .ZN(n9016)
         );
  OAI21_X1 U10356 ( .B1(n9017), .B2(n9095), .A(n9016), .ZN(P1_U3214) );
  XOR2_X1 U10357 ( .A(n9019), .B(n9018), .Z(n9023) );
  NAND2_X1 U10358 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9185) );
  OAI21_X1 U10359 ( .B1(n9106), .B2(n9318), .A(n9185), .ZN(n9021) );
  OAI22_X1 U10360 ( .A1(n9108), .A2(n9352), .B1(n9047), .B2(n9110), .ZN(n9020)
         );
  AOI211_X1 U10361 ( .C1(n9429), .C2(n9100), .A(n9021), .B(n9020), .ZN(n9022)
         );
  OAI21_X1 U10362 ( .B1(n9023), .B2(n9095), .A(n9022), .ZN(P1_U3217) );
  XOR2_X1 U10363 ( .A(n9024), .B(n9025), .Z(n9030) );
  INV_X1 U10364 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9026) );
  OAI22_X1 U10365 ( .A1(n9106), .A2(n9319), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9026), .ZN(n9028) );
  OAI22_X1 U10366 ( .A1(n9108), .A2(n9310), .B1(n9318), .B2(n9110), .ZN(n9027)
         );
  AOI211_X1 U10367 ( .C1(n9420), .C2(n9100), .A(n9028), .B(n9027), .ZN(n9029)
         );
  OAI21_X1 U10368 ( .B1(n9030), .B2(n9095), .A(n9029), .ZN(P1_U3221) );
  XNOR2_X1 U10369 ( .A(n9031), .B(n9032), .ZN(n9033) );
  NAND2_X1 U10370 ( .A1(n9033), .A2(n9102), .ZN(n9039) );
  OAI22_X1 U10371 ( .A1(n9108), .A2(n9251), .B1(n9034), .B2(n9110), .ZN(n9037)
         );
  OAI22_X1 U10372 ( .A1(n9106), .A2(n9228), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9035), .ZN(n9036) );
  NOR2_X1 U10373 ( .A1(n9037), .A2(n9036), .ZN(n9038) );
  OAI211_X1 U10374 ( .C1(n9254), .C2(n9115), .A(n9039), .B(n9038), .ZN(
        P1_U3223) );
  OR2_X1 U10375 ( .A1(n8039), .A2(n9040), .ZN(n9042) );
  NAND2_X1 U10376 ( .A1(n9042), .A2(n9041), .ZN(n9043) );
  XOR2_X1 U10377 ( .A(n9044), .B(n9043), .Z(n9052) );
  OAI21_X1 U10378 ( .B1(n9110), .B2(n9046), .A(n9045), .ZN(n9050) );
  OAI22_X1 U10379 ( .A1(n9108), .A2(n9048), .B1(n9047), .B2(n9106), .ZN(n9049)
         );
  AOI211_X1 U10380 ( .C1(n9440), .C2(n9100), .A(n9050), .B(n9049), .ZN(n9051)
         );
  OAI21_X1 U10381 ( .B1(n9052), .B2(n9095), .A(n9051), .ZN(P1_U3226) );
  XOR2_X1 U10382 ( .A(n9054), .B(n9053), .Z(n9059) );
  OAI22_X1 U10383 ( .A1(n9110), .A2(n9269), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9055), .ZN(n9057) );
  OAI22_X1 U10384 ( .A1(n9108), .A2(n9273), .B1(n9268), .B2(n9106), .ZN(n9056)
         );
  AOI211_X1 U10385 ( .C1(n9405), .C2(n9100), .A(n9057), .B(n9056), .ZN(n9058)
         );
  OAI21_X1 U10386 ( .B1(n9059), .B2(n9095), .A(n9058), .ZN(P1_U3227) );
  OAI211_X1 U10387 ( .C1(n9060), .C2(n9063), .A(n9062), .B(n9102), .ZN(n9070)
         );
  INV_X1 U10388 ( .A(n9064), .ZN(n9065) );
  AOI22_X1 U10389 ( .A1(n9089), .A2(n9065), .B1(n9088), .B2(n9126), .ZN(n9069)
         );
  AND2_X1 U10390 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9583) );
  NOR2_X1 U10391 ( .A1(n9110), .A2(n9066), .ZN(n9067) );
  AOI211_X1 U10392 ( .C1(n9100), .C2(n9688), .A(n9583), .B(n9067), .ZN(n9068)
         );
  NAND3_X1 U10393 ( .A1(n9070), .A2(n9069), .A3(n9068), .ZN(P1_U3228) );
  XOR2_X1 U10394 ( .A(n9071), .B(n9072), .Z(n9076) );
  OAI22_X1 U10395 ( .A1(n9106), .A2(n9083), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10029), .ZN(n9074) );
  OAI22_X1 U10396 ( .A1(n9108), .A2(n9326), .B1(n9363), .B2(n9110), .ZN(n9073)
         );
  AOI211_X1 U10397 ( .C1(n9423), .C2(n9100), .A(n9074), .B(n9073), .ZN(n9075)
         );
  OAI21_X1 U10398 ( .B1(n9076), .B2(n9095), .A(n9075), .ZN(P1_U3231) );
  INV_X1 U10399 ( .A(n9077), .ZN(n9079) );
  INV_X1 U10400 ( .A(n9080), .ZN(n9078) );
  OAI21_X1 U10401 ( .B1(n9081), .B2(n9079), .A(n9078), .ZN(n9082) );
  AOI22_X1 U10402 ( .A1(n9082), .A2(n4921), .B1(n9081), .B2(n9080), .ZN(n9087)
         );
  OAI22_X1 U10403 ( .A1(n9106), .A2(n9269), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9955), .ZN(n9085) );
  OAI22_X1 U10404 ( .A1(n9108), .A2(n9296), .B1(n9083), .B2(n9110), .ZN(n9084)
         );
  AOI211_X1 U10405 ( .C1(n9413), .C2(n9100), .A(n9085), .B(n9084), .ZN(n9086)
         );
  OAI21_X1 U10406 ( .B1(n9087), .B2(n9095), .A(n9086), .ZN(P1_U3233) );
  AOI22_X1 U10407 ( .A1(n9089), .A2(n9367), .B1(n9088), .B2(n9332), .ZN(n9090)
         );
  NAND2_X1 U10408 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9160) );
  OAI211_X1 U10409 ( .C1(n9362), .C2(n9110), .A(n9090), .B(n9160), .ZN(n9099)
         );
  INV_X1 U10410 ( .A(n9091), .ZN(n9097) );
  AOI21_X1 U10411 ( .B1(n9096), .B2(n9092), .A(n9093), .ZN(n9094) );
  AOI211_X1 U10412 ( .C1(n9097), .C2(n9096), .A(n9095), .B(n9094), .ZN(n9098)
         );
  AOI211_X1 U10413 ( .C1(n9100), .C2(n9435), .A(n9099), .B(n9098), .ZN(n9101)
         );
  INV_X1 U10414 ( .A(n9101), .ZN(P1_U3236) );
  OAI211_X1 U10415 ( .C1(n9105), .C2(n9104), .A(n9103), .B(n9102), .ZN(n9114)
         );
  OAI22_X1 U10416 ( .A1(n9108), .A2(n9237), .B1(n9107), .B2(n9106), .ZN(n9112)
         );
  OAI22_X1 U10417 ( .A1(n9110), .A2(n9268), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9109), .ZN(n9111) );
  NOR2_X1 U10418 ( .A1(n9112), .A2(n9111), .ZN(n9113) );
  OAI211_X1 U10419 ( .C1(n9240), .C2(n9115), .A(n9114), .B(n9113), .ZN(
        P1_U3238) );
  MUX2_X1 U10420 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9116), .S(n9904), .Z(
        P1_U3585) );
  MUX2_X1 U10421 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9212), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10422 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9117), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10423 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9244), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10424 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9259), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10425 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9243), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10426 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9286), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10427 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9287), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10428 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9333), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10429 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9347), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10430 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9332), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10431 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9346), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10432 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9504), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10433 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9118), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10434 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9503), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10435 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9119), .S(n9904), .Z(
        P1_U3569) );
  MUX2_X1 U10436 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9525), .S(n9904), .Z(
        P1_U3568) );
  MUX2_X1 U10437 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9120), .S(n9904), .Z(
        P1_U3567) );
  MUX2_X1 U10438 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9527), .S(n9904), .Z(
        P1_U3566) );
  MUX2_X1 U10439 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9121), .S(n9904), .Z(
        P1_U3565) );
  MUX2_X1 U10440 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9122), .S(n9904), .Z(
        P1_U3564) );
  MUX2_X1 U10441 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9123), .S(n9904), .Z(
        P1_U3563) );
  MUX2_X1 U10442 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9124), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10443 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9125), .S(n9904), .Z(
        P1_U3561) );
  MUX2_X1 U10444 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9126), .S(n9904), .Z(
        P1_U3560) );
  MUX2_X1 U10445 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9127), .S(n9904), .Z(
        P1_U3559) );
  MUX2_X1 U10446 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9128), .S(n9904), .Z(
        P1_U3558) );
  MUX2_X1 U10447 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9129), .S(n9904), .Z(
        P1_U3557) );
  MUX2_X1 U10448 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9130), .S(n9904), .Z(
        P1_U3556) );
  MUX2_X1 U10449 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6695), .S(n9904), .Z(
        P1_U3555) );
  NAND2_X1 U10450 ( .A1(n9146), .A2(P1_ADDR_REG_1__SCAN_IN), .ZN(n9141) );
  AOI22_X1 U10451 ( .A1(n9585), .A2(n9131), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        P1_U3084), .ZN(n9140) );
  OAI211_X1 U10452 ( .C1(n9134), .C2(n9133), .A(n9593), .B(n9132), .ZN(n9139)
         );
  OAI211_X1 U10453 ( .C1(n9137), .C2(n9136), .A(n9615), .B(n9135), .ZN(n9138)
         );
  NAND4_X1 U10454 ( .A1(n9141), .A2(n9140), .A3(n9139), .A4(n9138), .ZN(
        P1_U3242) );
  OAI21_X1 U10455 ( .B1(n9144), .B2(n9143), .A(n9142), .ZN(n9145) );
  AOI22_X1 U10456 ( .A1(n9146), .A2(P1_ADDR_REG_7__SCAN_IN), .B1(n9615), .B2(
        n9145), .ZN(n9155) );
  AOI21_X1 U10457 ( .B1(n9585), .B2(n9148), .A(n9147), .ZN(n9154) );
  OAI21_X1 U10458 ( .B1(n9151), .B2(n9150), .A(n9149), .ZN(n9152) );
  NAND2_X1 U10459 ( .A1(n9593), .A2(n9152), .ZN(n9153) );
  NAND3_X1 U10460 ( .A1(n9155), .A2(n9154), .A3(n9153), .ZN(P1_U3248) );
  INV_X1 U10461 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9170) );
  XNOR2_X1 U10462 ( .A(n9175), .B(n9156), .ZN(n9159) );
  AOI21_X1 U10463 ( .B1(n9163), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9157), .ZN(
        n9158) );
  NAND2_X1 U10464 ( .A1(n9159), .A2(n9158), .ZN(n9174) );
  OAI21_X1 U10465 ( .B1(n9159), .B2(n9158), .A(n9174), .ZN(n9168) );
  INV_X1 U10466 ( .A(n9175), .ZN(n9161) );
  OAI21_X1 U10467 ( .B1(n9617), .B2(n9161), .A(n9160), .ZN(n9167) );
  AOI21_X1 U10468 ( .B1(n9163), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9162), .ZN(
        n9165) );
  XNOR2_X1 U10469 ( .A(n9175), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n9164) );
  NOR2_X1 U10470 ( .A1(n9165), .A2(n9164), .ZN(n9171) );
  AOI211_X1 U10471 ( .C1(n9165), .C2(n9164), .A(n9171), .B(n9598), .ZN(n9166)
         );
  AOI211_X1 U10472 ( .C1(n9593), .C2(n9168), .A(n9167), .B(n9166), .ZN(n9169)
         );
  OAI21_X1 U10473 ( .B1(n9619), .B2(n9170), .A(n9169), .ZN(P1_U3259) );
  INV_X1 U10474 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9186) );
  AOI21_X1 U10475 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n9175), .A(n9171), .ZN(
        n9172) );
  XNOR2_X1 U10476 ( .A(n9173), .B(n9172), .ZN(n9179) );
  OAI21_X1 U10477 ( .B1(n9175), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9174), .ZN(
        n9177) );
  XNOR2_X1 U10478 ( .A(n9177), .B(n9176), .ZN(n9183) );
  OAI22_X1 U10479 ( .A1(n9179), .A2(n9598), .B1(n9183), .B2(n9608), .ZN(n9178)
         );
  INV_X1 U10480 ( .A(n9178), .ZN(n9184) );
  INV_X1 U10481 ( .A(n9179), .ZN(n9182) );
  NAND2_X1 U10482 ( .A1(n9194), .A2(n9193), .ZN(n9192) );
  XNOR2_X1 U10483 ( .A(n9192), .B(n9375), .ZN(n9377) );
  NOR2_X1 U10484 ( .A1(n9665), .A2(n9187), .ZN(n9190) );
  NAND2_X1 U10485 ( .A1(n9189), .A2(n9188), .ZN(n9543) );
  NOR2_X1 U10486 ( .A1(n4389), .A2(n9543), .ZN(n9195) );
  AOI211_X1 U10487 ( .C1(n9375), .C2(n9531), .A(n9190), .B(n9195), .ZN(n9191)
         );
  OAI21_X1 U10488 ( .B1(n9377), .B2(n9198), .A(n9191), .ZN(P1_U3261) );
  OAI21_X1 U10489 ( .B1(n9194), .B2(n9193), .A(n9192), .ZN(n9544) );
  NOR2_X1 U10490 ( .A1(n9665), .A2(n6067), .ZN(n9196) );
  AOI211_X1 U10491 ( .C1(n9547), .C2(n9531), .A(n9196), .B(n9195), .ZN(n9197)
         );
  OAI21_X1 U10492 ( .B1(n9198), .B2(n9544), .A(n9197), .ZN(P1_U3262) );
  AOI21_X1 U10493 ( .B1(n9211), .B2(n9200), .A(n9199), .ZN(n9201) );
  INV_X1 U10494 ( .A(n9201), .ZN(n9387) );
  INV_X1 U10495 ( .A(n9221), .ZN(n9204) );
  INV_X1 U10496 ( .A(n9202), .ZN(n9203) );
  AOI21_X1 U10497 ( .B1(n9383), .B2(n9204), .A(n9203), .ZN(n9384) );
  INV_X1 U10498 ( .A(n9205), .ZN(n9206) );
  AOI22_X1 U10499 ( .A1(n4389), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9206), .B2(
        n9653), .ZN(n9207) );
  OAI21_X1 U10500 ( .B1(n9208), .B2(n9370), .A(n9207), .ZN(n9218) );
  OAI21_X1 U10501 ( .B1(n9211), .B2(n9210), .A(n9209), .ZN(n9216) );
  NAND2_X1 U10502 ( .A1(n9212), .A2(n9524), .ZN(n9214) );
  NAND2_X1 U10503 ( .A1(n9244), .A2(n9526), .ZN(n9213) );
  NOR2_X1 U10504 ( .A1(n9386), .A2(n4389), .ZN(n9217) );
  AOI211_X1 U10505 ( .C1(n9384), .C2(n9337), .A(n9218), .B(n9217), .ZN(n9219)
         );
  OAI21_X1 U10506 ( .B1(n9387), .B2(n9374), .A(n9219), .ZN(P1_U3263) );
  XNOR2_X1 U10507 ( .A(n9220), .B(n9227), .ZN(n9392) );
  AOI21_X1 U10508 ( .B1(n9388), .B2(n9235), .A(n9221), .ZN(n9389) );
  INV_X1 U10509 ( .A(n9222), .ZN(n9223) );
  AOI22_X1 U10510 ( .A1(n4389), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9223), .B2(
        n9653), .ZN(n9224) );
  OAI21_X1 U10511 ( .B1(n4679), .B2(n9370), .A(n9224), .ZN(n9233) );
  AOI211_X1 U10512 ( .C1(n9227), .C2(n9226), .A(n9657), .B(n9225), .ZN(n9231)
         );
  OAI22_X1 U10513 ( .A1(n9229), .A2(n9662), .B1(n9660), .B2(n9228), .ZN(n9230)
         );
  NOR2_X1 U10514 ( .A1(n9231), .A2(n9230), .ZN(n9391) );
  NOR2_X1 U10515 ( .A1(n9391), .A2(n4389), .ZN(n9232) );
  AOI211_X1 U10516 ( .C1(n9337), .C2(n9389), .A(n9233), .B(n9232), .ZN(n9234)
         );
  OAI21_X1 U10517 ( .B1(n9392), .B2(n9374), .A(n9234), .ZN(P1_U3264) );
  XNOR2_X1 U10518 ( .A(n4417), .B(n9241), .ZN(n9397) );
  INV_X1 U10519 ( .A(n9235), .ZN(n9236) );
  AOI21_X1 U10520 ( .B1(n9393), .B2(n4681), .A(n9236), .ZN(n9394) );
  INV_X1 U10521 ( .A(n9237), .ZN(n9238) );
  AOI22_X1 U10522 ( .A1(n4389), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9238), .B2(
        n9653), .ZN(n9239) );
  OAI21_X1 U10523 ( .B1(n9240), .B2(n9370), .A(n9239), .ZN(n9247) );
  XNOR2_X1 U10524 ( .A(n9242), .B(n9241), .ZN(n9245) );
  AOI222_X1 U10525 ( .A1(n9635), .A2(n9245), .B1(n9244), .B2(n9524), .C1(n9243), .C2(n9526), .ZN(n9396) );
  NOR2_X1 U10526 ( .A1(n9396), .A2(n4389), .ZN(n9246) );
  AOI211_X1 U10527 ( .C1(n9394), .C2(n9337), .A(n9247), .B(n9246), .ZN(n9248)
         );
  OAI21_X1 U10528 ( .B1(n9397), .B2(n9374), .A(n9248), .ZN(P1_U3265) );
  XOR2_X1 U10529 ( .A(n9257), .B(n9249), .Z(n9402) );
  AOI21_X1 U10530 ( .B1(n9398), .B2(n9270), .A(n9250), .ZN(n9399) );
  INV_X1 U10531 ( .A(n9251), .ZN(n9252) );
  AOI22_X1 U10532 ( .A1(n4389), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9252), .B2(
        n9653), .ZN(n9253) );
  OAI21_X1 U10533 ( .B1(n9254), .B2(n9370), .A(n9253), .ZN(n9262) );
  INV_X1 U10534 ( .A(n9255), .ZN(n9256) );
  NOR2_X1 U10535 ( .A1(n4392), .A2(n9256), .ZN(n9258) );
  XNOR2_X1 U10536 ( .A(n9258), .B(n9257), .ZN(n9260) );
  AOI222_X1 U10537 ( .A1(n9635), .A2(n9260), .B1(n9259), .B2(n9524), .C1(n9286), .C2(n9526), .ZN(n9401) );
  NOR2_X1 U10538 ( .A1(n9401), .A2(n4389), .ZN(n9261) );
  AOI211_X1 U10539 ( .C1(n9399), .C2(n9337), .A(n9262), .B(n9261), .ZN(n9263)
         );
  OAI21_X1 U10540 ( .B1(n9402), .B2(n9374), .A(n9263), .ZN(P1_U3266) );
  XOR2_X1 U10541 ( .A(n9264), .B(n9266), .Z(n9407) );
  AOI22_X1 U10542 ( .A1(n9405), .A2(n9531), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n4389), .ZN(n9277) );
  AOI21_X1 U10543 ( .B1(n9266), .B2(n9265), .A(n4392), .ZN(n9267) );
  OAI222_X1 U10544 ( .A1(n9660), .A2(n9269), .B1(n9662), .B2(n9268), .C1(n9657), .C2(n9267), .ZN(n9403) );
  INV_X1 U10545 ( .A(n9279), .ZN(n9272) );
  INV_X1 U10546 ( .A(n9270), .ZN(n9271) );
  AOI211_X1 U10547 ( .C1(n9405), .C2(n9272), .A(n9705), .B(n9271), .ZN(n9404)
         );
  INV_X1 U10548 ( .A(n9404), .ZN(n9274) );
  OAI22_X1 U10549 ( .A1(n9274), .A2(n4486), .B1(n9629), .B2(n9273), .ZN(n9275)
         );
  OAI21_X1 U10550 ( .B1(n9403), .B2(n9275), .A(n9665), .ZN(n9276) );
  OAI211_X1 U10551 ( .C1(n9407), .C2(n9374), .A(n9277), .B(n9276), .ZN(
        P1_U3267) );
  XNOR2_X1 U10552 ( .A(n9278), .B(n9284), .ZN(n9412) );
  AOI21_X1 U10553 ( .B1(n9408), .B2(n9293), .A(n9279), .ZN(n9409) );
  INV_X1 U10554 ( .A(n9280), .ZN(n9281) );
  AOI22_X1 U10555 ( .A1(n4389), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9281), .B2(
        n9653), .ZN(n9282) );
  OAI21_X1 U10556 ( .B1(n9283), .B2(n9370), .A(n9282), .ZN(n9290) );
  XNOR2_X1 U10557 ( .A(n9285), .B(n9284), .ZN(n9288) );
  AOI222_X1 U10558 ( .A1(n9635), .A2(n9288), .B1(n9287), .B2(n9526), .C1(n9286), .C2(n9524), .ZN(n9411) );
  NOR2_X1 U10559 ( .A1(n9411), .A2(n4389), .ZN(n9289) );
  AOI211_X1 U10560 ( .C1(n9409), .C2(n9337), .A(n9290), .B(n9289), .ZN(n9291)
         );
  OAI21_X1 U10561 ( .B1(n9412), .B2(n9374), .A(n9291), .ZN(P1_U3268) );
  XOR2_X1 U10562 ( .A(n9301), .B(n9292), .Z(n9417) );
  INV_X1 U10563 ( .A(n9308), .ZN(n9295) );
  INV_X1 U10564 ( .A(n9293), .ZN(n9294) );
  AOI21_X1 U10565 ( .B1(n9413), .B2(n9295), .A(n9294), .ZN(n9414) );
  INV_X1 U10566 ( .A(n9296), .ZN(n9297) );
  AOI22_X1 U10567 ( .A1(n4389), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9297), .B2(
        n9653), .ZN(n9298) );
  OAI21_X1 U10568 ( .B1(n9299), .B2(n9370), .A(n9298), .ZN(n9304) );
  XOR2_X1 U10569 ( .A(n9301), .B(n9300), .Z(n9302) );
  AOI222_X1 U10570 ( .A1(n9635), .A2(n9302), .B1(n9333), .B2(n9526), .C1(n9905), .C2(n9524), .ZN(n9416) );
  NOR2_X1 U10571 ( .A1(n9416), .A2(n4389), .ZN(n9303) );
  AOI211_X1 U10572 ( .C1(n9414), .C2(n9337), .A(n9304), .B(n9303), .ZN(n9305)
         );
  OAI21_X1 U10573 ( .B1(n9374), .B2(n9417), .A(n9305), .ZN(P1_U3269) );
  XNOR2_X1 U10574 ( .A(n9307), .B(n9306), .ZN(n9422) );
  AOI211_X1 U10575 ( .C1(n9420), .C2(n9323), .A(n9705), .B(n9308), .ZN(n9419)
         );
  NOR2_X1 U10576 ( .A1(n9309), .A2(n9370), .ZN(n9313) );
  OAI22_X1 U10577 ( .A1(n9665), .A2(n9311), .B1(n9310), .B2(n9629), .ZN(n9312)
         );
  AOI211_X1 U10578 ( .C1(n9419), .C2(n9539), .A(n9313), .B(n9312), .ZN(n9321)
         );
  AOI21_X1 U10579 ( .B1(n9316), .B2(n9315), .A(n9314), .ZN(n9317) );
  OAI222_X1 U10580 ( .A1(n9662), .A2(n9319), .B1(n9660), .B2(n9318), .C1(n9657), .C2(n9317), .ZN(n9418) );
  NAND2_X1 U10581 ( .A1(n9418), .A2(n9665), .ZN(n9320) );
  OAI211_X1 U10582 ( .C1(n9422), .C2(n9374), .A(n9321), .B(n9320), .ZN(
        P1_U3270) );
  XOR2_X1 U10583 ( .A(n9322), .B(n9331), .Z(n9427) );
  INV_X1 U10584 ( .A(n9349), .ZN(n9325) );
  INV_X1 U10585 ( .A(n9323), .ZN(n9324) );
  AOI21_X1 U10586 ( .B1(n9423), .B2(n9325), .A(n9324), .ZN(n9424) );
  INV_X1 U10587 ( .A(n9326), .ZN(n9327) );
  AOI22_X1 U10588 ( .A1(n4389), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9327), .B2(
        n9653), .ZN(n9328) );
  OAI21_X1 U10589 ( .B1(n9329), .B2(n9370), .A(n9328), .ZN(n9336) );
  XOR2_X1 U10590 ( .A(n9331), .B(n9330), .Z(n9334) );
  AOI222_X1 U10591 ( .A1(n9635), .A2(n9334), .B1(n9333), .B2(n9524), .C1(n9332), .C2(n9526), .ZN(n9426) );
  NOR2_X1 U10592 ( .A1(n9426), .A2(n4389), .ZN(n9335) );
  AOI211_X1 U10593 ( .C1(n9424), .C2(n9337), .A(n9336), .B(n9335), .ZN(n9338)
         );
  OAI21_X1 U10594 ( .B1(n9427), .B2(n9374), .A(n9338), .ZN(P1_U3271) );
  XNOR2_X1 U10595 ( .A(n9340), .B(n9339), .ZN(n9432) );
  NAND2_X1 U10596 ( .A1(n9342), .A2(n9341), .ZN(n9344) );
  OAI21_X1 U10597 ( .B1(n9345), .B2(n9344), .A(n9343), .ZN(n9348) );
  AOI222_X1 U10598 ( .A1(n9635), .A2(n9348), .B1(n9347), .B2(n9524), .C1(n9346), .C2(n9526), .ZN(n9431) );
  AOI211_X1 U10599 ( .C1(n9429), .C2(n9365), .A(n9705), .B(n9349), .ZN(n9428)
         );
  NAND2_X1 U10600 ( .A1(n9428), .A2(n9350), .ZN(n9351) );
  OAI211_X1 U10601 ( .C1(n9629), .C2(n9352), .A(n9431), .B(n9351), .ZN(n9353)
         );
  NAND2_X1 U10602 ( .A1(n9353), .A2(n9665), .ZN(n9355) );
  AOI22_X1 U10603 ( .A1(n9429), .A2(n9531), .B1(P1_REG2_REG_19__SCAN_IN), .B2(
        n4389), .ZN(n9354) );
  OAI211_X1 U10604 ( .C1(n9432), .C2(n9374), .A(n9355), .B(n9354), .ZN(
        P1_U3272) );
  XNOR2_X1 U10605 ( .A(n9356), .B(n9360), .ZN(n9437) );
  NAND2_X1 U10606 ( .A1(n9358), .A2(n9357), .ZN(n9359) );
  XOR2_X1 U10607 ( .A(n9360), .B(n9359), .Z(n9361) );
  OAI222_X1 U10608 ( .A1(n9662), .A2(n9363), .B1(n9660), .B2(n9362), .C1(n9657), .C2(n9361), .ZN(n9433) );
  INV_X1 U10609 ( .A(n9365), .ZN(n9366) );
  AOI211_X1 U10610 ( .C1(n9435), .C2(n4684), .A(n9705), .B(n9366), .ZN(n9434)
         );
  NAND2_X1 U10611 ( .A1(n9434), .A2(n9539), .ZN(n9369) );
  AOI22_X1 U10612 ( .A1(n4389), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9367), .B2(
        n9653), .ZN(n9368) );
  OAI211_X1 U10613 ( .C1(n9371), .C2(n9370), .A(n9369), .B(n9368), .ZN(n9372)
         );
  AOI21_X1 U10614 ( .B1(n9433), .B2(n9665), .A(n9372), .ZN(n9373) );
  OAI21_X1 U10615 ( .B1(n9374), .B2(n9437), .A(n9373), .ZN(P1_U3273) );
  NAND2_X1 U10616 ( .A1(n9375), .A2(n9689), .ZN(n9376) );
  OAI211_X1 U10617 ( .C1(n9377), .C2(n9705), .A(n9543), .B(n9376), .ZN(n9443)
         );
  MUX2_X1 U10618 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9443), .S(n9742), .Z(
        P1_U3554) );
  AOI22_X1 U10619 ( .A1(n9381), .A2(n9690), .B1(n9689), .B2(n9380), .ZN(n9382)
         );
  AOI22_X1 U10620 ( .A1(n9384), .A2(n9690), .B1(n9689), .B2(n9383), .ZN(n9385)
         );
  OAI211_X1 U10621 ( .C1(n9387), .C2(n9710), .A(n9386), .B(n9385), .ZN(n9444)
         );
  MUX2_X1 U10622 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9444), .S(n9742), .Z(
        P1_U3551) );
  AOI22_X1 U10623 ( .A1(n9389), .A2(n9690), .B1(n9689), .B2(n9388), .ZN(n9390)
         );
  OAI211_X1 U10624 ( .C1(n9392), .C2(n9710), .A(n9391), .B(n9390), .ZN(n9445)
         );
  MUX2_X1 U10625 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9445), .S(n9742), .Z(
        P1_U3550) );
  AOI22_X1 U10626 ( .A1(n9394), .A2(n9690), .B1(n9689), .B2(n9393), .ZN(n9395)
         );
  OAI211_X1 U10627 ( .C1(n9397), .C2(n9710), .A(n9396), .B(n9395), .ZN(n9446)
         );
  MUX2_X1 U10628 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9446), .S(n9742), .Z(
        P1_U3549) );
  AOI22_X1 U10629 ( .A1(n9399), .A2(n9690), .B1(n9689), .B2(n9398), .ZN(n9400)
         );
  OAI211_X1 U10630 ( .C1(n9402), .C2(n9710), .A(n9401), .B(n9400), .ZN(n9447)
         );
  MUX2_X1 U10631 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9447), .S(n9742), .Z(
        P1_U3548) );
  AOI211_X1 U10632 ( .C1(n9689), .C2(n9405), .A(n9404), .B(n9403), .ZN(n9406)
         );
  OAI21_X1 U10633 ( .B1(n9407), .B2(n9710), .A(n9406), .ZN(n9448) );
  MUX2_X1 U10634 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9448), .S(n9742), .Z(
        P1_U3547) );
  AOI22_X1 U10635 ( .A1(n9409), .A2(n9690), .B1(n9689), .B2(n9408), .ZN(n9410)
         );
  OAI211_X1 U10636 ( .C1(n9412), .C2(n9710), .A(n9411), .B(n9410), .ZN(n9449)
         );
  MUX2_X1 U10637 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9449), .S(n9742), .Z(
        P1_U3546) );
  AOI22_X1 U10638 ( .A1(n9414), .A2(n9690), .B1(n9689), .B2(n9413), .ZN(n9415)
         );
  OAI211_X1 U10639 ( .C1(n9417), .C2(n9710), .A(n9416), .B(n9415), .ZN(n9450)
         );
  MUX2_X1 U10640 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9450), .S(n9742), .Z(
        P1_U3545) );
  AOI211_X1 U10641 ( .C1(n9689), .C2(n9420), .A(n9419), .B(n9418), .ZN(n9421)
         );
  OAI21_X1 U10642 ( .B1(n9710), .B2(n9422), .A(n9421), .ZN(n9451) );
  MUX2_X1 U10643 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9451), .S(n9742), .Z(
        P1_U3544) );
  AOI22_X1 U10644 ( .A1(n9424), .A2(n9690), .B1(n9689), .B2(n9423), .ZN(n9425)
         );
  OAI211_X1 U10645 ( .C1(n9427), .C2(n9710), .A(n9426), .B(n9425), .ZN(n9452)
         );
  MUX2_X1 U10646 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9452), .S(n9742), .Z(
        P1_U3543) );
  AOI21_X1 U10647 ( .B1(n9689), .B2(n9429), .A(n9428), .ZN(n9430) );
  OAI211_X1 U10648 ( .C1(n9432), .C2(n9710), .A(n9431), .B(n9430), .ZN(n9453)
         );
  MUX2_X1 U10649 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9453), .S(n9742), .Z(
        P1_U3542) );
  AOI211_X1 U10650 ( .C1(n9689), .C2(n9435), .A(n9434), .B(n9433), .ZN(n9436)
         );
  OAI21_X1 U10651 ( .B1(n9710), .B2(n9437), .A(n9436), .ZN(n9454) );
  MUX2_X1 U10652 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9454), .S(n9742), .Z(
        P1_U3541) );
  AOI211_X1 U10653 ( .C1(n9689), .C2(n9440), .A(n9439), .B(n9438), .ZN(n9441)
         );
  OAI21_X1 U10654 ( .B1(n9442), .B2(n9710), .A(n9441), .ZN(n9455) );
  MUX2_X1 U10655 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9455), .S(n9742), .Z(
        P1_U3540) );
  MUX2_X1 U10656 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9443), .S(n9726), .Z(
        P1_U3522) );
  MUX2_X1 U10657 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9444), .S(n9726), .Z(
        P1_U3519) );
  MUX2_X1 U10658 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9445), .S(n9726), .Z(
        P1_U3518) );
  MUX2_X1 U10659 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9446), .S(n9726), .Z(
        P1_U3517) );
  MUX2_X1 U10660 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9447), .S(n9726), .Z(
        P1_U3516) );
  MUX2_X1 U10661 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9448), .S(n9726), .Z(
        P1_U3515) );
  MUX2_X1 U10662 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9449), .S(n9726), .Z(
        P1_U3514) );
  MUX2_X1 U10663 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9450), .S(n9726), .Z(
        P1_U3513) );
  MUX2_X1 U10664 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9451), .S(n9726), .Z(
        P1_U3512) );
  MUX2_X1 U10665 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9452), .S(n9726), .Z(
        P1_U3511) );
  MUX2_X1 U10666 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9453), .S(n9726), .Z(
        P1_U3510) );
  MUX2_X1 U10667 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9454), .S(n9726), .Z(
        P1_U3508) );
  MUX2_X1 U10668 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9455), .S(n9726), .Z(
        P1_U3505) );
  AOI22_X1 U10669 ( .A1(n9766), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n9466) );
  AOI211_X1 U10670 ( .C1(n9458), .C2(n9457), .A(n9456), .B(n9761), .ZN(n9459)
         );
  AOI21_X1 U10671 ( .B1(n9472), .B2(n9460), .A(n9459), .ZN(n9465) );
  AND2_X1 U10672 ( .A1(n9765), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9463) );
  OAI211_X1 U10673 ( .C1(n9463), .C2(n9462), .A(n9764), .B(n9461), .ZN(n9464)
         );
  NAND3_X1 U10674 ( .A1(n9466), .A2(n9465), .A3(n9464), .ZN(P2_U3246) );
  AOI22_X1 U10675 ( .A1(n9766), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9478) );
  AOI211_X1 U10676 ( .C1(n9469), .C2(n9468), .A(n9467), .B(n9761), .ZN(n9470)
         );
  AOI21_X1 U10677 ( .B1(n9472), .B2(n9471), .A(n9470), .ZN(n9477) );
  OAI211_X1 U10678 ( .C1(n9475), .C2(n9474), .A(n9764), .B(n9473), .ZN(n9476)
         );
  NAND3_X1 U10679 ( .A1(n9478), .A2(n9477), .A3(n9476), .ZN(P2_U3247) );
  INV_X1 U10680 ( .A(n9710), .ZN(n9722) );
  OAI21_X1 U10681 ( .B1(n4687), .B2(n9718), .A(n9480), .ZN(n9482) );
  AOI211_X1 U10682 ( .C1(n9722), .C2(n9483), .A(n9482), .B(n9481), .ZN(n9484)
         );
  INV_X1 U10683 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10110) );
  AOI22_X1 U10684 ( .A1(n9726), .A2(n9484), .B1(n10110), .B2(n9724), .ZN(
        P1_U3484) );
  AOI22_X1 U10685 ( .A1(n9742), .A2(n9484), .B1(n5841), .B2(n9739), .ZN(
        P1_U3533) );
  INV_X1 U10686 ( .A(n9485), .ZN(n9857) );
  OAI211_X1 U10687 ( .C1(n9853), .C2(n9488), .A(n9487), .B(n9486), .ZN(n9489)
         );
  AOI21_X1 U10688 ( .B1(n9490), .B2(n9857), .A(n9489), .ZN(n9498) );
  AOI22_X1 U10689 ( .A1(n9875), .A2(n9498), .B1(n8591), .B2(n9873), .ZN(
        P2_U3536) );
  NAND2_X1 U10690 ( .A1(n9491), .A2(n9818), .ZN(n9492) );
  OAI211_X1 U10691 ( .C1(n9853), .C2(n9494), .A(n9493), .B(n9492), .ZN(n9495)
         );
  AOI21_X1 U10692 ( .B1(n9496), .B2(n9857), .A(n9495), .ZN(n9500) );
  AOI22_X1 U10693 ( .A1(n9875), .A2(n9500), .B1(n5141), .B2(n9873), .ZN(
        P2_U3534) );
  INV_X1 U10694 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9497) );
  AOI22_X1 U10695 ( .A1(n9861), .A2(n9498), .B1(n9497), .B2(n9859), .ZN(
        P2_U3499) );
  INV_X1 U10696 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9499) );
  AOI22_X1 U10697 ( .A1(n9861), .A2(n9500), .B1(n9499), .B2(n9859), .ZN(
        P2_U3493) );
  XNOR2_X1 U10698 ( .A(n9501), .B(n9510), .ZN(n9502) );
  NAND2_X1 U10699 ( .A1(n9502), .A2(n9635), .ZN(n9506) );
  AOI22_X1 U10700 ( .A1(n9504), .A2(n9524), .B1(n9526), .B2(n9503), .ZN(n9505)
         );
  AND2_X1 U10701 ( .A1(n9506), .A2(n9505), .ZN(n9551) );
  INV_X1 U10702 ( .A(n9507), .ZN(n9508) );
  AOI222_X1 U10703 ( .A1(n9549), .A2(n9531), .B1(P1_REG2_REG_16__SCAN_IN), 
        .B2(n4389), .C1(n9508), .C2(n9653), .ZN(n9519) );
  NAND2_X1 U10704 ( .A1(n9509), .A2(n9510), .ZN(n9511) );
  AND2_X1 U10705 ( .A1(n9512), .A2(n9511), .ZN(n9554) );
  AOI21_X1 U10706 ( .B1(n9513), .B2(n9549), .A(n9705), .ZN(n9515) );
  NAND2_X1 U10707 ( .A1(n9515), .A2(n9514), .ZN(n9550) );
  NOR2_X1 U10708 ( .A1(n9550), .A2(n9516), .ZN(n9517) );
  AOI21_X1 U10709 ( .B1(n9554), .B2(n9540), .A(n9517), .ZN(n9518) );
  OAI211_X1 U10710 ( .C1(n4389), .C2(n9551), .A(n9519), .B(n9518), .ZN(
        P1_U3275) );
  NAND2_X1 U10711 ( .A1(n9521), .A2(n9520), .ZN(n9523) );
  XNOR2_X1 U10712 ( .A(n9523), .B(n9522), .ZN(n9528) );
  AOI222_X1 U10713 ( .A1(n9635), .A2(n9528), .B1(n9527), .B2(n9526), .C1(n9525), .C2(n9524), .ZN(n9562) );
  INV_X1 U10714 ( .A(n9529), .ZN(n9530) );
  AOI222_X1 U10715 ( .A1(n9532), .A2(n9531), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n4389), .C1(n9653), .C2(n9530), .ZN(n9542) );
  INV_X1 U10716 ( .A(n9533), .ZN(n9534) );
  AOI21_X1 U10717 ( .B1(n9535), .B2(n7409), .A(n9534), .ZN(n9565) );
  OAI211_X1 U10718 ( .C1(n9537), .C2(n9563), .A(n9690), .B(n9536), .ZN(n9561)
         );
  INV_X1 U10719 ( .A(n9561), .ZN(n9538) );
  AOI22_X1 U10720 ( .A1(n9565), .A2(n9540), .B1(n9539), .B2(n9538), .ZN(n9541)
         );
  OAI211_X1 U10721 ( .C1(n4389), .C2(n9562), .A(n9542), .B(n9541), .ZN(
        P1_U3279) );
  INV_X1 U10722 ( .A(n9543), .ZN(n9546) );
  NOR2_X1 U10723 ( .A1(n9544), .A2(n9705), .ZN(n9545) );
  INV_X1 U10724 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9548) );
  AOI22_X1 U10725 ( .A1(n9742), .A2(n9567), .B1(n9548), .B2(n9739), .ZN(
        P1_U3553) );
  INV_X1 U10726 ( .A(n9549), .ZN(n9552) );
  OAI211_X1 U10727 ( .C1(n9552), .C2(n9718), .A(n9551), .B(n9550), .ZN(n9553)
         );
  AOI21_X1 U10728 ( .B1(n9554), .B2(n9722), .A(n9553), .ZN(n9569) );
  AOI22_X1 U10729 ( .A1(n9742), .A2(n9569), .B1(n9555), .B2(n9739), .ZN(
        P1_U3539) );
  OAI211_X1 U10730 ( .C1(n9558), .C2(n9718), .A(n9557), .B(n9556), .ZN(n9559)
         );
  AOI21_X1 U10731 ( .B1(n9560), .B2(n9722), .A(n9559), .ZN(n9570) );
  AOI22_X1 U10732 ( .A1(n9742), .A2(n9570), .B1(n6412), .B2(n9739), .ZN(
        P1_U3537) );
  OAI211_X1 U10733 ( .C1(n9563), .C2(n9718), .A(n9562), .B(n9561), .ZN(n9564)
         );
  AOI21_X1 U10734 ( .B1(n9565), .B2(n9722), .A(n9564), .ZN(n9572) );
  AOI22_X1 U10735 ( .A1(n9742), .A2(n9572), .B1(n6429), .B2(n9739), .ZN(
        P1_U3535) );
  INV_X1 U10736 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9566) );
  AOI22_X1 U10737 ( .A1(n9726), .A2(n9567), .B1(n9566), .B2(n9724), .ZN(
        P1_U3521) );
  INV_X1 U10738 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9568) );
  AOI22_X1 U10739 ( .A1(n9726), .A2(n9569), .B1(n9568), .B2(n9724), .ZN(
        P1_U3502) );
  INV_X1 U10740 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10172) );
  AOI22_X1 U10741 ( .A1(n9726), .A2(n9570), .B1(n10172), .B2(n9724), .ZN(
        P1_U3496) );
  INV_X1 U10742 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9571) );
  AOI22_X1 U10743 ( .A1(n9726), .A2(n9572), .B1(n9571), .B2(n9724), .ZN(
        P1_U3490) );
  XNOR2_X1 U10744 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X1 U10745 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9588) );
  AOI21_X1 U10746 ( .B1(n9575), .B2(n9574), .A(n9573), .ZN(n9580) );
  AOI21_X1 U10747 ( .B1(n9578), .B2(n9577), .A(n9576), .ZN(n9579) );
  OAI22_X1 U10748 ( .A1(n9608), .A2(n9580), .B1(n9579), .B2(n9598), .ZN(n9581)
         );
  INV_X1 U10749 ( .A(n9581), .ZN(n9587) );
  AOI211_X1 U10750 ( .C1(n9585), .C2(n9584), .A(n9583), .B(n9582), .ZN(n9586)
         );
  OAI211_X1 U10751 ( .C1(n9619), .C2(n9588), .A(n9587), .B(n9586), .ZN(
        P1_U3245) );
  XNOR2_X1 U10752 ( .A(n9590), .B(n9589), .ZN(n9592) );
  AOI21_X1 U10753 ( .B1(n9593), .B2(n9592), .A(n9591), .ZN(n9600) );
  AND2_X1 U10754 ( .A1(n9595), .A2(n9594), .ZN(n9596) );
  OR3_X1 U10755 ( .A1(n9598), .A2(n9597), .A3(n9596), .ZN(n9599) );
  AND2_X1 U10756 ( .A1(n9600), .A2(n9599), .ZN(n9604) );
  OAI22_X1 U10757 ( .A1(n9619), .A2(n10107), .B1(n9617), .B2(n9601), .ZN(n9602) );
  INV_X1 U10758 ( .A(n9602), .ZN(n9603) );
  NAND2_X1 U10759 ( .A1(n9604), .A2(n9603), .ZN(P1_U3247) );
  OAI21_X1 U10760 ( .B1(n9607), .B2(n9606), .A(n9605), .ZN(n9614) );
  AOI211_X1 U10761 ( .C1(n9611), .C2(n9610), .A(n9609), .B(n9608), .ZN(n9612)
         );
  AOI211_X1 U10762 ( .C1(n9615), .C2(n9614), .A(n9613), .B(n9612), .ZN(n9622)
         );
  INV_X1 U10763 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9618) );
  OAI22_X1 U10764 ( .A1(n9619), .A2(n9618), .B1(n9617), .B2(n9616), .ZN(n9620)
         );
  INV_X1 U10765 ( .A(n9620), .ZN(n9621) );
  NAND2_X1 U10766 ( .A1(n9622), .A2(n9621), .ZN(P1_U3249) );
  NAND2_X1 U10767 ( .A1(n9623), .A2(n9633), .ZN(n9624) );
  AND2_X1 U10768 ( .A1(n9625), .A2(n9624), .ZN(n9723) );
  OAI211_X1 U10769 ( .C1(n9627), .C2(n9719), .A(n9690), .B(n9626), .ZN(n9717)
         );
  NOR2_X1 U10770 ( .A1(n9629), .A2(n9628), .ZN(n9630) );
  AOI21_X1 U10771 ( .B1(n9631), .B2(n4487), .A(n9630), .ZN(n9632) );
  OAI21_X1 U10772 ( .B1(n9717), .B2(n4486), .A(n9632), .ZN(n9642) );
  XNOR2_X1 U10773 ( .A(n9634), .B(n9633), .ZN(n9636) );
  NAND2_X1 U10774 ( .A1(n9636), .A2(n9635), .ZN(n9641) );
  OAI22_X1 U10775 ( .A1(n9638), .A2(n9660), .B1(n9662), .B2(n9637), .ZN(n9639)
         );
  INV_X1 U10776 ( .A(n9639), .ZN(n9640) );
  NAND2_X1 U10777 ( .A1(n9641), .A2(n9640), .ZN(n9720) );
  AOI211_X1 U10778 ( .C1(n9723), .C2(n9664), .A(n9642), .B(n9720), .ZN(n9643)
         );
  AOI22_X1 U10779 ( .A1(n4389), .A2(n5828), .B1(n9643), .B2(n9665), .ZN(
        P1_U3283) );
  INV_X1 U10780 ( .A(n9644), .ZN(n9645) );
  INV_X1 U10781 ( .A(n9646), .ZN(n9647) );
  AOI21_X1 U10782 ( .B1(n9656), .B2(n9645), .A(n9647), .ZN(n9701) );
  AOI21_X1 U10783 ( .B1(n9648), .B2(n9651), .A(n9705), .ZN(n9650) );
  NAND2_X1 U10784 ( .A1(n9650), .A2(n9649), .ZN(n9697) );
  AOI22_X1 U10785 ( .A1(n9653), .A2(n9652), .B1(n4487), .B2(n9651), .ZN(n9654)
         );
  OAI21_X1 U10786 ( .B1(n9697), .B2(n4486), .A(n9654), .ZN(n9663) );
  XOR2_X1 U10787 ( .A(n9656), .B(n9655), .Z(n9658) );
  OAI222_X1 U10788 ( .A1(n9662), .A2(n9661), .B1(n9660), .B2(n9659), .C1(n9658), .C2(n9657), .ZN(n9699) );
  AOI211_X1 U10789 ( .C1(n9664), .C2(n9701), .A(n9663), .B(n9699), .ZN(n9666)
         );
  AOI22_X1 U10790 ( .A1(n4389), .A2(n6398), .B1(n9666), .B2(n9665), .ZN(
        P1_U3286) );
  AND2_X1 U10791 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9668), .ZN(P1_U3292) );
  AND2_X1 U10792 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9668), .ZN(P1_U3293) );
  AND2_X1 U10793 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9668), .ZN(P1_U3294) );
  AND2_X1 U10794 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9668), .ZN(P1_U3295) );
  INV_X1 U10795 ( .A(n9668), .ZN(n9667) );
  INV_X1 U10796 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10075) );
  NOR2_X1 U10797 ( .A1(n9667), .A2(n10075), .ZN(P1_U3296) );
  AND2_X1 U10798 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9668), .ZN(P1_U3297) );
  AND2_X1 U10799 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9668), .ZN(P1_U3298) );
  AND2_X1 U10800 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9668), .ZN(P1_U3299) );
  INV_X1 U10801 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10086) );
  NOR2_X1 U10802 ( .A1(n9667), .A2(n10086), .ZN(P1_U3300) );
  AND2_X1 U10803 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9668), .ZN(P1_U3301) );
  AND2_X1 U10804 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9668), .ZN(P1_U3302) );
  AND2_X1 U10805 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9668), .ZN(P1_U3303) );
  AND2_X1 U10806 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9668), .ZN(P1_U3304) );
  AND2_X1 U10807 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9668), .ZN(P1_U3305) );
  AND2_X1 U10808 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9668), .ZN(P1_U3306) );
  AND2_X1 U10809 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9668), .ZN(P1_U3307) );
  AND2_X1 U10810 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9668), .ZN(P1_U3308) );
  AND2_X1 U10811 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9668), .ZN(P1_U3309) );
  AND2_X1 U10812 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9668), .ZN(P1_U3310) );
  INV_X1 U10813 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10084) );
  NOR2_X1 U10814 ( .A1(n9667), .A2(n10084), .ZN(P1_U3311) );
  INV_X1 U10815 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10016) );
  NOR2_X1 U10816 ( .A1(n9667), .A2(n10016), .ZN(P1_U3312) );
  AND2_X1 U10817 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9668), .ZN(P1_U3313) );
  AND2_X1 U10818 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9668), .ZN(P1_U3314) );
  INV_X1 U10819 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10008) );
  NOR2_X1 U10820 ( .A1(n9667), .A2(n10008), .ZN(P1_U3315) );
  AND2_X1 U10821 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9668), .ZN(P1_U3316) );
  AND2_X1 U10822 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9668), .ZN(P1_U3317) );
  AND2_X1 U10823 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9668), .ZN(P1_U3318) );
  INV_X1 U10824 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10063) );
  NOR2_X1 U10825 ( .A1(n9667), .A2(n10063), .ZN(P1_U3319) );
  AND2_X1 U10826 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9668), .ZN(P1_U3320) );
  AND2_X1 U10827 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9668), .ZN(P1_U3321) );
  INV_X1 U10828 ( .A(n9669), .ZN(n9674) );
  OAI21_X1 U10829 ( .B1(n9671), .B2(n9718), .A(n9670), .ZN(n9673) );
  AOI211_X1 U10830 ( .C1(n9687), .C2(n9674), .A(n9673), .B(n9672), .ZN(n9728)
         );
  INV_X1 U10831 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10174) );
  AOI22_X1 U10832 ( .A1(n9726), .A2(n9728), .B1(n10174), .B2(n9724), .ZN(
        P1_U3457) );
  INV_X1 U10833 ( .A(n9675), .ZN(n9680) );
  OAI22_X1 U10834 ( .A1(n9677), .A2(n9705), .B1(n9718), .B2(n9676), .ZN(n9679)
         );
  AOI211_X1 U10835 ( .C1(n9687), .C2(n9680), .A(n9679), .B(n9678), .ZN(n9730)
         );
  INV_X1 U10836 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9971) );
  AOI22_X1 U10837 ( .A1(n9726), .A2(n9730), .B1(n9971), .B2(n9724), .ZN(
        P1_U3460) );
  NAND2_X1 U10838 ( .A1(n9681), .A2(n9690), .ZN(n9682) );
  OAI21_X1 U10839 ( .B1(n9683), .B2(n9718), .A(n9682), .ZN(n9685) );
  AOI211_X1 U10840 ( .C1(n9687), .C2(n9686), .A(n9685), .B(n9684), .ZN(n9731)
         );
  AOI22_X1 U10841 ( .A1(n9726), .A2(n9731), .B1(n5768), .B2(n9724), .ZN(
        P1_U3463) );
  AOI22_X1 U10842 ( .A1(n9691), .A2(n9690), .B1(n9689), .B2(n9688), .ZN(n9692)
         );
  OAI211_X1 U10843 ( .C1(n9695), .C2(n9694), .A(n9693), .B(n9692), .ZN(n9696)
         );
  INV_X1 U10844 ( .A(n9696), .ZN(n9733) );
  INV_X1 U10845 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10078) );
  AOI22_X1 U10846 ( .A1(n9726), .A2(n9733), .B1(n10078), .B2(n9724), .ZN(
        P1_U3466) );
  OAI21_X1 U10847 ( .B1(n9698), .B2(n9718), .A(n9697), .ZN(n9700) );
  AOI211_X1 U10848 ( .C1(n9701), .C2(n9722), .A(n9700), .B(n9699), .ZN(n9735)
         );
  INV_X1 U10849 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9702) );
  AOI22_X1 U10850 ( .A1(n9726), .A2(n9735), .B1(n9702), .B2(n9724), .ZN(
        P1_U3469) );
  INV_X1 U10851 ( .A(n9703), .ZN(n9704) );
  OAI21_X1 U10852 ( .B1(n9706), .B2(n9705), .A(n9704), .ZN(n9708) );
  AOI211_X1 U10853 ( .C1(n9709), .C2(n9722), .A(n9708), .B(n9707), .ZN(n9737)
         );
  INV_X1 U10854 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10134) );
  AOI22_X1 U10855 ( .A1(n9726), .A2(n9737), .B1(n10134), .B2(n9724), .ZN(
        P1_U3472) );
  NOR2_X1 U10856 ( .A1(n9711), .A2(n9710), .ZN(n9715) );
  NOR4_X1 U10857 ( .A1(n9715), .A2(n9714), .A3(n9713), .A4(n9712), .ZN(n9738)
         );
  INV_X1 U10858 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9716) );
  AOI22_X1 U10859 ( .A1(n9726), .A2(n9738), .B1(n9716), .B2(n9724), .ZN(
        P1_U3475) );
  OAI21_X1 U10860 ( .B1(n9719), .B2(n9718), .A(n9717), .ZN(n9721) );
  AOI211_X1 U10861 ( .C1(n9723), .C2(n9722), .A(n9721), .B(n9720), .ZN(n9741)
         );
  INV_X1 U10862 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9725) );
  AOI22_X1 U10863 ( .A1(n9726), .A2(n9741), .B1(n9725), .B2(n9724), .ZN(
        P1_U3478) );
  AOI22_X1 U10864 ( .A1(n9742), .A2(n9728), .B1(n9727), .B2(n9739), .ZN(
        P1_U3524) );
  AOI22_X1 U10865 ( .A1(n9742), .A2(n9730), .B1(n9729), .B2(n9739), .ZN(
        P1_U3525) );
  AOI22_X1 U10866 ( .A1(n9742), .A2(n9731), .B1(n5765), .B2(n9739), .ZN(
        P1_U3526) );
  AOI22_X1 U10867 ( .A1(n9742), .A2(n9733), .B1(n9732), .B2(n9739), .ZN(
        P1_U3527) );
  INV_X1 U10868 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9734) );
  AOI22_X1 U10869 ( .A1(n9742), .A2(n9735), .B1(n9734), .B2(n9739), .ZN(
        P1_U3528) );
  INV_X1 U10870 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9736) );
  AOI22_X1 U10871 ( .A1(n9742), .A2(n9737), .B1(n9736), .B2(n9739), .ZN(
        P1_U3529) );
  AOI22_X1 U10872 ( .A1(n9742), .A2(n9738), .B1(n5819), .B2(n9739), .ZN(
        P1_U3530) );
  INV_X1 U10873 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9740) );
  AOI22_X1 U10874 ( .A1(n9742), .A2(n9741), .B1(n9740), .B2(n9739), .ZN(
        P1_U3531) );
  AOI21_X1 U10875 ( .B1(n9745), .B2(n9744), .A(n9743), .ZN(n9756) );
  OAI22_X1 U10876 ( .A1(n9747), .A2(n9746), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10169), .ZN(n9754) );
  INV_X1 U10877 ( .A(n9748), .ZN(n9749) );
  OAI22_X1 U10878 ( .A1(n9752), .A2(n9751), .B1(n9750), .B2(n9749), .ZN(n9753)
         );
  AOI211_X1 U10879 ( .C1(n9756), .C2(n9755), .A(n9754), .B(n9753), .ZN(n9757)
         );
  OAI21_X1 U10880 ( .B1(n9759), .B2(n9758), .A(n9757), .ZN(P2_U3229) );
  INV_X1 U10881 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10060) );
  OAI211_X1 U10882 ( .C1(n9761), .C2(P2_REG1_REG_0__SCAN_IN), .A(n9760), .B(
        n9765), .ZN(n9762) );
  AOI21_X1 U10883 ( .B1(n9764), .B2(n5198), .A(n9762), .ZN(n9770) );
  AOI22_X1 U10884 ( .A1(n9764), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n9763), .B2(
        P2_REG1_REG_0__SCAN_IN), .ZN(n9769) );
  INV_X1 U10885 ( .A(n9765), .ZN(n9768) );
  AOI22_X1 U10886 ( .A1(n9766), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9767) );
  OAI221_X1 U10887 ( .B1(n9770), .B2(n9769), .C1(n9770), .C2(n9768), .A(n9767), 
        .ZN(P2_U3245) );
  XNOR2_X1 U10888 ( .A(n9771), .B(n9781), .ZN(n9776) );
  AOI222_X1 U10889 ( .A1(n9777), .A2(n9776), .B1(n9775), .B2(n9774), .C1(n9773), .C2(n9772), .ZN(n9836) );
  OAI22_X1 U10890 ( .A1(n6620), .A2(n8870), .B1(n9779), .B2(n9778), .ZN(n9780)
         );
  INV_X1 U10891 ( .A(n9780), .ZN(n9789) );
  XOR2_X1 U10892 ( .A(n9782), .B(n9781), .Z(n9839) );
  OAI211_X1 U10893 ( .C1(n9783), .C2(n9785), .A(n9819), .B(n4963), .ZN(n9784)
         );
  OAI21_X1 U10894 ( .B1(n9785), .B2(n9851), .A(n9784), .ZN(n9838) );
  AOI22_X1 U10895 ( .A1(n9839), .A2(n9787), .B1(n9838), .B2(n9786), .ZN(n9788)
         );
  OAI211_X1 U10896 ( .C1(n4388), .C2(n9836), .A(n9789), .B(n9788), .ZN(
        P2_U3290) );
  NOR2_X1 U10897 ( .A1(n9791), .A2(n9790), .ZN(n9792) );
  INV_X1 U10898 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n9928) );
  NOR2_X1 U10899 ( .A1(n9792), .A2(n9928), .ZN(P2_U3297) );
  AND2_X1 U10900 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9795), .ZN(P2_U3298) );
  INV_X1 U10901 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n9926) );
  NOR2_X1 U10902 ( .A1(n9792), .A2(n9926), .ZN(P2_U3299) );
  AND2_X1 U10903 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9795), .ZN(P2_U3300) );
  AND2_X1 U10904 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9795), .ZN(P2_U3301) );
  AND2_X1 U10905 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9795), .ZN(P2_U3302) );
  AND2_X1 U10906 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9795), .ZN(P2_U3303) );
  INV_X1 U10907 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n10087) );
  NOR2_X1 U10908 ( .A1(n9792), .A2(n10087), .ZN(P2_U3304) );
  AND2_X1 U10909 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9795), .ZN(P2_U3305) );
  AND2_X1 U10910 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9795), .ZN(P2_U3306) );
  INV_X1 U10911 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n10025) );
  NOR2_X1 U10912 ( .A1(n9792), .A2(n10025), .ZN(P2_U3307) );
  INV_X1 U10913 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n9917) );
  NOR2_X1 U10914 ( .A1(n9792), .A2(n9917), .ZN(P2_U3308) );
  AND2_X1 U10915 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9795), .ZN(P2_U3309) );
  AND2_X1 U10916 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9795), .ZN(P2_U3310) );
  AND2_X1 U10917 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9795), .ZN(P2_U3311) );
  AND2_X1 U10918 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9795), .ZN(P2_U3312) );
  AND2_X1 U10919 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9795), .ZN(P2_U3313) );
  INV_X1 U10920 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n9942) );
  NOR2_X1 U10921 ( .A1(n9792), .A2(n9942), .ZN(P2_U3314) );
  AND2_X1 U10922 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9795), .ZN(P2_U3315) );
  AND2_X1 U10923 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9795), .ZN(P2_U3316) );
  INV_X1 U10924 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n10170) );
  NOR2_X1 U10925 ( .A1(n9792), .A2(n10170), .ZN(P2_U3317) );
  AND2_X1 U10926 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9795), .ZN(P2_U3318) );
  AND2_X1 U10927 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9795), .ZN(P2_U3319) );
  AND2_X1 U10928 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9795), .ZN(P2_U3320) );
  AND2_X1 U10929 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9795), .ZN(P2_U3321) );
  AND2_X1 U10930 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9795), .ZN(P2_U3322) );
  AND2_X1 U10931 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9795), .ZN(P2_U3323) );
  AND2_X1 U10932 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9795), .ZN(P2_U3324) );
  AND2_X1 U10933 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9795), .ZN(P2_U3325) );
  AND2_X1 U10934 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9795), .ZN(P2_U3326) );
  AOI22_X1 U10935 ( .A1(n9794), .A2(n9795), .B1(n9798), .B2(n9793), .ZN(
        P2_U3437) );
  AOI22_X1 U10936 ( .A1(n9798), .A2(n9797), .B1(n9796), .B2(n9795), .ZN(
        P2_U3438) );
  OAI21_X1 U10937 ( .B1(n9801), .B2(n9800), .A(n9799), .ZN(n9802) );
  AOI21_X1 U10938 ( .B1(n9857), .B2(n9803), .A(n9802), .ZN(n9862) );
  INV_X1 U10939 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9804) );
  AOI22_X1 U10940 ( .A1(n9861), .A2(n9862), .B1(n9804), .B2(n9859), .ZN(
        P2_U3451) );
  INV_X1 U10941 ( .A(n9805), .ZN(n9809) );
  INV_X1 U10942 ( .A(n9806), .ZN(n9807) );
  AOI211_X1 U10943 ( .C1(n9857), .C2(n9809), .A(n9808), .B(n9807), .ZN(n9863)
         );
  AOI22_X1 U10944 ( .A1(n9861), .A2(n9863), .B1(n5187), .B2(n9859), .ZN(
        P2_U3454) );
  INV_X1 U10945 ( .A(n9810), .ZN(n9816) );
  OAI22_X1 U10946 ( .A1(n9812), .A2(n9853), .B1(n9811), .B2(n9851), .ZN(n9815)
         );
  INV_X1 U10947 ( .A(n9813), .ZN(n9814) );
  AOI211_X1 U10948 ( .C1(n9857), .C2(n9816), .A(n9815), .B(n9814), .ZN(n9865)
         );
  AOI22_X1 U10949 ( .A1(n9861), .A2(n9865), .B1(n5212), .B2(n9859), .ZN(
        P2_U3457) );
  AOI22_X1 U10950 ( .A1(n9820), .A2(n9819), .B1(n9818), .B2(n9817), .ZN(n9821)
         );
  OAI211_X1 U10951 ( .C1(n9824), .C2(n9823), .A(n9822), .B(n9821), .ZN(n9825)
         );
  AOI21_X1 U10952 ( .B1(n9827), .B2(n9826), .A(n9825), .ZN(n9866) );
  INV_X1 U10953 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9828) );
  AOI22_X1 U10954 ( .A1(n9861), .A2(n9866), .B1(n9828), .B2(n9859), .ZN(
        P2_U3460) );
  NAND2_X1 U10955 ( .A1(n9829), .A2(n9857), .ZN(n9835) );
  OAI22_X1 U10956 ( .A1(n9831), .A2(n9853), .B1(n9830), .B2(n9851), .ZN(n9832)
         );
  INV_X1 U10957 ( .A(n9832), .ZN(n9833) );
  AND3_X1 U10958 ( .A1(n9835), .A2(n9834), .A3(n9833), .ZN(n9867) );
  AOI22_X1 U10959 ( .A1(n9861), .A2(n9867), .B1(n5254), .B2(n9859), .ZN(
        P2_U3463) );
  INV_X1 U10960 ( .A(n9836), .ZN(n9837) );
  AOI211_X1 U10961 ( .C1(n9839), .C2(n9857), .A(n9838), .B(n9837), .ZN(n9869)
         );
  INV_X1 U10962 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9959) );
  AOI22_X1 U10963 ( .A1(n9861), .A2(n9869), .B1(n9959), .B2(n9859), .ZN(
        P2_U3469) );
  OAI22_X1 U10964 ( .A1(n9841), .A2(n9853), .B1(n9840), .B2(n9851), .ZN(n9843)
         );
  AOI211_X1 U10965 ( .C1(n9845), .C2(n9844), .A(n9843), .B(n9842), .ZN(n9871)
         );
  AOI22_X1 U10966 ( .A1(n9861), .A2(n9871), .B1(n5333), .B2(n9859), .ZN(
        P2_U3475) );
  INV_X1 U10967 ( .A(n9846), .ZN(n9850) );
  OAI22_X1 U10968 ( .A1(n9847), .A2(n9853), .B1(n4702), .B2(n9851), .ZN(n9849)
         );
  AOI211_X1 U10969 ( .C1(n9850), .C2(n9857), .A(n9849), .B(n9848), .ZN(n9872)
         );
  AOI22_X1 U10970 ( .A1(n9861), .A2(n9872), .B1(n5376), .B2(n9859), .ZN(
        P2_U3481) );
  OAI22_X1 U10971 ( .A1(n9854), .A2(n9853), .B1(n9852), .B2(n9851), .ZN(n9856)
         );
  AOI211_X1 U10972 ( .C1(n9858), .C2(n9857), .A(n9856), .B(n9855), .ZN(n9874)
         );
  INV_X1 U10973 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9860) );
  AOI22_X1 U10974 ( .A1(n9861), .A2(n9874), .B1(n9860), .B2(n9859), .ZN(
        P2_U3487) );
  AOI22_X1 U10975 ( .A1(n9875), .A2(n9862), .B1(n10060), .B2(n9873), .ZN(
        P2_U3520) );
  AOI22_X1 U10976 ( .A1(n9875), .A2(n9863), .B1(n6565), .B2(n9873), .ZN(
        P2_U3521) );
  INV_X1 U10977 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9864) );
  AOI22_X1 U10978 ( .A1(n9875), .A2(n9865), .B1(n9864), .B2(n9873), .ZN(
        P2_U3522) );
  AOI22_X1 U10979 ( .A1(n9875), .A2(n9866), .B1(n6567), .B2(n9873), .ZN(
        P2_U3523) );
  AOI22_X1 U10980 ( .A1(n9875), .A2(n9867), .B1(n6564), .B2(n9873), .ZN(
        P2_U3524) );
  INV_X1 U10981 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9868) );
  AOI22_X1 U10982 ( .A1(n9875), .A2(n9869), .B1(n9868), .B2(n9873), .ZN(
        P2_U3526) );
  INV_X1 U10983 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9870) );
  AOI22_X1 U10984 ( .A1(n9875), .A2(n9871), .B1(n9870), .B2(n9873), .ZN(
        P2_U3528) );
  AOI22_X1 U10985 ( .A1(n9875), .A2(n9872), .B1(n6879), .B2(n9873), .ZN(
        P2_U3530) );
  AOI22_X1 U10986 ( .A1(n9875), .A2(n9874), .B1(n7079), .B2(n9873), .ZN(
        P2_U3532) );
  INV_X1 U10987 ( .A(n9876), .ZN(n9877) );
  NAND2_X1 U10988 ( .A1(n9878), .A2(n9877), .ZN(n9879) );
  XNOR2_X1 U10989 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9879), .ZN(ADD_1071_U5) );
  XOR2_X1 U10990 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U10991 ( .B1(n9882), .B2(n9881), .A(n9880), .ZN(ADD_1071_U56) );
  OAI21_X1 U10992 ( .B1(n9885), .B2(n9884), .A(n9883), .ZN(ADD_1071_U57) );
  OAI21_X1 U10993 ( .B1(n9888), .B2(n9887), .A(n9886), .ZN(ADD_1071_U58) );
  AOI21_X1 U10994 ( .B1(n9891), .B2(n9890), .A(n9889), .ZN(ADD_1071_U59) );
  AOI21_X1 U10995 ( .B1(n9894), .B2(n9893), .A(n9892), .ZN(ADD_1071_U60) );
  OAI21_X1 U10996 ( .B1(n9897), .B2(n9896), .A(n9895), .ZN(ADD_1071_U61) );
  AOI21_X1 U10997 ( .B1(n9900), .B2(n9899), .A(n9898), .ZN(ADD_1071_U62) );
  AOI21_X1 U10998 ( .B1(n9903), .B2(n9902), .A(n9901), .ZN(ADD_1071_U63) );
  MUX2_X1 U10999 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9905), .S(n9904), .Z(
        n10105) );
  AOI22_X1 U11000 ( .A1(n10110), .A2(keyinput49), .B1(keyinput70), .B2(n10109), 
        .ZN(n9906) );
  OAI221_X1 U11001 ( .B1(n10110), .B2(keyinput49), .C1(n10109), .C2(keyinput70), .A(n9906), .ZN(n9914) );
  AOI22_X1 U11002 ( .A1(n9908), .A2(keyinput100), .B1(keyinput123), .B2(n5748), 
        .ZN(n9907) );
  OAI221_X1 U11003 ( .B1(n9908), .B2(keyinput100), .C1(n5748), .C2(keyinput123), .A(n9907), .ZN(n9913) );
  AOI22_X1 U11004 ( .A1(n6023), .A2(keyinput45), .B1(n10137), .B2(keyinput95), 
        .ZN(n9909) );
  OAI221_X1 U11005 ( .B1(n6023), .B2(keyinput45), .C1(n10137), .C2(keyinput95), 
        .A(n9909), .ZN(n9912) );
  AOI22_X1 U11006 ( .A1(n7393), .A2(keyinput65), .B1(n6871), .B2(keyinput29), 
        .ZN(n9910) );
  OAI221_X1 U11007 ( .B1(n7393), .B2(keyinput65), .C1(n6871), .C2(keyinput29), 
        .A(n9910), .ZN(n9911) );
  NOR4_X1 U11008 ( .A1(n9914), .A2(n9913), .A3(n9912), .A4(n9911), .ZN(n9952)
         );
  AOI22_X1 U11009 ( .A1(n6200), .A2(keyinput6), .B1(keyinput9), .B2(n6067), 
        .ZN(n9915) );
  OAI221_X1 U11010 ( .B1(n6200), .B2(keyinput6), .C1(n6067), .C2(keyinput9), 
        .A(n9915), .ZN(n9924) );
  AOI22_X1 U11011 ( .A1(n10138), .A2(keyinput60), .B1(keyinput113), .B2(n9917), 
        .ZN(n9916) );
  OAI221_X1 U11012 ( .B1(n10138), .B2(keyinput60), .C1(n9917), .C2(keyinput113), .A(n9916), .ZN(n9923) );
  AOI22_X1 U11013 ( .A1(n7932), .A2(keyinput30), .B1(n6620), .B2(keyinput94), 
        .ZN(n9918) );
  OAI221_X1 U11014 ( .B1(n7932), .B2(keyinput30), .C1(n6620), .C2(keyinput94), 
        .A(n9918), .ZN(n9922) );
  XOR2_X1 U11015 ( .A(n7244), .B(keyinput122), .Z(n9920) );
  XNOR2_X1 U11016 ( .A(P1_RD_REG_SCAN_IN), .B(keyinput3), .ZN(n9919) );
  NAND2_X1 U11017 ( .A1(n9920), .A2(n9919), .ZN(n9921) );
  NOR4_X1 U11018 ( .A1(n9924), .A2(n9923), .A3(n9922), .A4(n9921), .ZN(n9951)
         );
  INV_X1 U11019 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10108) );
  AOI22_X1 U11020 ( .A1(n9926), .A2(keyinput0), .B1(keyinput23), .B2(n10108), 
        .ZN(n9925) );
  OAI221_X1 U11021 ( .B1(n9926), .B2(keyinput0), .C1(n10108), .C2(keyinput23), 
        .A(n9925), .ZN(n9936) );
  AOI22_X1 U11022 ( .A1(n5068), .A2(keyinput88), .B1(keyinput31), .B2(n9928), 
        .ZN(n9927) );
  OAI221_X1 U11023 ( .B1(n5068), .B2(keyinput88), .C1(n9928), .C2(keyinput31), 
        .A(n9927), .ZN(n9935) );
  XOR2_X1 U11024 ( .A(n6057), .B(keyinput33), .Z(n9933) );
  INV_X1 U11025 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n9929) );
  XOR2_X1 U11026 ( .A(n9929), .B(keyinput77), .Z(n9932) );
  XNOR2_X1 U11027 ( .A(P2_IR_REG_17__SCAN_IN), .B(keyinput119), .ZN(n9931) );
  XNOR2_X1 U11028 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput108), .ZN(n9930) );
  NAND4_X1 U11029 ( .A1(n9933), .A2(n9932), .A3(n9931), .A4(n9930), .ZN(n9934)
         );
  NOR3_X1 U11030 ( .A1(n9936), .A2(n9935), .A3(n9934), .ZN(n9950) );
  INV_X1 U11031 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n9938) );
  AOI22_X1 U11032 ( .A1(n9939), .A2(keyinput20), .B1(keyinput115), .B2(n9938), 
        .ZN(n9937) );
  OAI221_X1 U11033 ( .B1(n9939), .B2(keyinput20), .C1(n9938), .C2(keyinput115), 
        .A(n9937), .ZN(n9948) );
  AOI22_X1 U11034 ( .A1(n10129), .A2(keyinput104), .B1(keyinput112), .B2(
        n10134), .ZN(n9940) );
  OAI221_X1 U11035 ( .B1(n10129), .B2(keyinput104), .C1(n10134), .C2(
        keyinput112), .A(n9940), .ZN(n9947) );
  AOI22_X1 U11036 ( .A1(n10131), .A2(keyinput71), .B1(n9942), .B2(keyinput22), 
        .ZN(n9941) );
  OAI221_X1 U11037 ( .B1(n10131), .B2(keyinput71), .C1(n9942), .C2(keyinput22), 
        .A(n9941), .ZN(n9946) );
  XNOR2_X1 U11038 ( .A(P1_REG3_REG_8__SCAN_IN), .B(keyinput18), .ZN(n9944) );
  XNOR2_X1 U11039 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput50), .ZN(n9943) );
  NAND2_X1 U11040 ( .A1(n9944), .A2(n9943), .ZN(n9945) );
  NOR4_X1 U11041 ( .A1(n9948), .A2(n9947), .A3(n9946), .A4(n9945), .ZN(n9949)
         );
  NAND4_X1 U11042 ( .A1(n9952), .A2(n9951), .A3(n9950), .A4(n9949), .ZN(n10103) );
  INV_X1 U11043 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n9954) );
  AOI22_X1 U11044 ( .A1(n9955), .A2(keyinput102), .B1(keyinput97), .B2(n9954), 
        .ZN(n9953) );
  OAI221_X1 U11045 ( .B1(n9955), .B2(keyinput102), .C1(n9954), .C2(keyinput97), 
        .A(n9953), .ZN(n9966) );
  AOI22_X1 U11046 ( .A1(n9958), .A2(keyinput47), .B1(keyinput35), .B2(n9957), 
        .ZN(n9956) );
  OAI221_X1 U11047 ( .B1(n9958), .B2(keyinput47), .C1(n9957), .C2(keyinput35), 
        .A(n9956), .ZN(n9965) );
  XOR2_X1 U11048 ( .A(n5080), .B(keyinput58), .Z(n9963) );
  XOR2_X1 U11049 ( .A(n9959), .B(keyinput1), .Z(n9962) );
  XNOR2_X1 U11050 ( .A(SI_0_), .B(keyinput121), .ZN(n9961) );
  XNOR2_X1 U11051 ( .A(P2_IR_REG_6__SCAN_IN), .B(keyinput7), .ZN(n9960) );
  NAND4_X1 U11052 ( .A1(n9963), .A2(n9962), .A3(n9961), .A4(n9960), .ZN(n9964)
         );
  NOR3_X1 U11053 ( .A1(n9966), .A2(n9965), .A3(n9964), .ZN(n10003) );
  INV_X1 U11054 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n10127) );
  AOI22_X1 U11055 ( .A1(n9968), .A2(keyinput64), .B1(keyinput36), .B2(n10127), 
        .ZN(n9967) );
  OAI221_X1 U11056 ( .B1(n9968), .B2(keyinput64), .C1(n10127), .C2(keyinput36), 
        .A(n9967), .ZN(n9979) );
  AOI22_X1 U11057 ( .A1(n9971), .A2(keyinput37), .B1(n9970), .B2(keyinput93), 
        .ZN(n9969) );
  OAI221_X1 U11058 ( .B1(n9971), .B2(keyinput37), .C1(n9970), .C2(keyinput93), 
        .A(n9969), .ZN(n9978) );
  AOI22_X1 U11059 ( .A1(n10151), .A2(keyinput55), .B1(n9973), .B2(keyinput13), 
        .ZN(n9972) );
  OAI221_X1 U11060 ( .B1(n10151), .B2(keyinput55), .C1(n9973), .C2(keyinput13), 
        .A(n9972), .ZN(n9977) );
  XNOR2_X1 U11061 ( .A(P1_REG3_REG_6__SCAN_IN), .B(keyinput99), .ZN(n9975) );
  XNOR2_X1 U11062 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput79), .ZN(n9974) );
  NAND2_X1 U11063 ( .A1(n9975), .A2(n9974), .ZN(n9976) );
  NOR4_X1 U11064 ( .A1(n9979), .A2(n9978), .A3(n9977), .A4(n9976), .ZN(n10002)
         );
  AOI22_X1 U11065 ( .A1(n6427), .A2(keyinput73), .B1(n10152), .B2(keyinput83), 
        .ZN(n9980) );
  OAI221_X1 U11066 ( .B1(n6427), .B2(keyinput73), .C1(n10152), .C2(keyinput83), 
        .A(n9980), .ZN(n9990) );
  AOI22_X1 U11067 ( .A1(n10150), .A2(keyinput72), .B1(keyinput117), .B2(n9982), 
        .ZN(n9981) );
  OAI221_X1 U11068 ( .B1(n10150), .B2(keyinput72), .C1(n9982), .C2(keyinput117), .A(n9981), .ZN(n9989) );
  AOI22_X1 U11069 ( .A1(n9985), .A2(keyinput12), .B1(n9984), .B2(keyinput17), 
        .ZN(n9983) );
  OAI221_X1 U11070 ( .B1(n9985), .B2(keyinput12), .C1(n9984), .C2(keyinput17), 
        .A(n9983), .ZN(n9988) );
  AOI22_X1 U11071 ( .A1(n6413), .A2(keyinput68), .B1(n10155), .B2(keyinput106), 
        .ZN(n9986) );
  OAI221_X1 U11072 ( .B1(n6413), .B2(keyinput68), .C1(n10155), .C2(keyinput106), .A(n9986), .ZN(n9987) );
  NOR4_X1 U11073 ( .A1(n9990), .A2(n9989), .A3(n9988), .A4(n9987), .ZN(n10001)
         );
  AOI22_X1 U11074 ( .A1(n6429), .A2(keyinput57), .B1(keyinput14), .B2(n10154), 
        .ZN(n9991) );
  OAI221_X1 U11075 ( .B1(n6429), .B2(keyinput57), .C1(n10154), .C2(keyinput14), 
        .A(n9991), .ZN(n9999) );
  AOI22_X1 U11076 ( .A1(n10153), .A2(keyinput126), .B1(keyinput92), .B2(n6032), 
        .ZN(n9992) );
  OAI221_X1 U11077 ( .B1(n10153), .B2(keyinput126), .C1(n6032), .C2(keyinput92), .A(n9992), .ZN(n9998) );
  AOI22_X1 U11078 ( .A1(n9994), .A2(keyinput59), .B1(keyinput118), .B2(n6565), 
        .ZN(n9993) );
  OAI221_X1 U11079 ( .B1(n9994), .B2(keyinput59), .C1(n6565), .C2(keyinput118), 
        .A(n9993), .ZN(n9997) );
  INV_X1 U11080 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10107) );
  AOI22_X1 U11081 ( .A1(n10107), .A2(keyinput105), .B1(n10145), .B2(keyinput39), .ZN(n9995) );
  OAI221_X1 U11082 ( .B1(n10107), .B2(keyinput105), .C1(n10145), .C2(
        keyinput39), .A(n9995), .ZN(n9996) );
  NOR4_X1 U11083 ( .A1(n9999), .A2(n9998), .A3(n9997), .A4(n9996), .ZN(n10000)
         );
  NAND4_X1 U11084 ( .A1(n10003), .A2(n10002), .A3(n10001), .A4(n10000), .ZN(
        n10102) );
  INV_X1 U11085 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n10112) );
  AOI22_X1 U11086 ( .A1(n10112), .A2(keyinput82), .B1(keyinput40), .B2(n7305), 
        .ZN(n10004) );
  OAI221_X1 U11087 ( .B1(n10112), .B2(keyinput82), .C1(n7305), .C2(keyinput40), 
        .A(n10004), .ZN(n10013) );
  AOI22_X1 U11088 ( .A1(n6069), .A2(keyinput96), .B1(keyinput34), .B2(n7791), 
        .ZN(n10005) );
  OAI221_X1 U11089 ( .B1(n6069), .B2(keyinput96), .C1(n7791), .C2(keyinput34), 
        .A(n10005), .ZN(n10012) );
  AOI22_X1 U11090 ( .A1(n5701), .A2(keyinput63), .B1(keyinput66), .B2(n8816), 
        .ZN(n10006) );
  OAI221_X1 U11091 ( .B1(n5701), .B2(keyinput63), .C1(n8816), .C2(keyinput66), 
        .A(n10006), .ZN(n10011) );
  AOI22_X1 U11092 ( .A1(n10009), .A2(keyinput52), .B1(n10008), .B2(keyinput24), 
        .ZN(n10007) );
  OAI221_X1 U11093 ( .B1(n10009), .B2(keyinput52), .C1(n10008), .C2(keyinput24), .A(n10007), .ZN(n10010) );
  NOR4_X1 U11094 ( .A1(n10013), .A2(n10012), .A3(n10011), .A4(n10010), .ZN(
        n10048) );
  AOI22_X1 U11095 ( .A1(n5623), .A2(keyinput114), .B1(keyinput28), .B2(n6564), 
        .ZN(n10014) );
  OAI221_X1 U11096 ( .B1(n5623), .B2(keyinput114), .C1(n6564), .C2(keyinput28), 
        .A(n10014), .ZN(n10023) );
  AOI22_X1 U11097 ( .A1(n10119), .A2(keyinput43), .B1(keyinput27), .B2(n10016), 
        .ZN(n10015) );
  OAI221_X1 U11098 ( .B1(n10119), .B2(keyinput43), .C1(n10016), .C2(keyinput27), .A(n10015), .ZN(n10022) );
  AOI22_X1 U11099 ( .A1(n6879), .A2(keyinput110), .B1(n10144), .B2(keyinput54), 
        .ZN(n10017) );
  OAI221_X1 U11100 ( .B1(n6879), .B2(keyinput110), .C1(n10144), .C2(keyinput54), .A(n10017), .ZN(n10021) );
  XOR2_X1 U11101 ( .A(n5850), .B(keyinput80), .Z(n10019) );
  XNOR2_X1 U11102 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput69), .ZN(n10018) );
  NAND2_X1 U11103 ( .A1(n10019), .A2(n10018), .ZN(n10020) );
  NOR4_X1 U11104 ( .A1(n10023), .A2(n10022), .A3(n10021), .A4(n10020), .ZN(
        n10047) );
  INV_X1 U11105 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10193) );
  AOI22_X1 U11106 ( .A1(n10025), .A2(keyinput103), .B1(keyinput53), .B2(n10193), .ZN(n10024) );
  OAI221_X1 U11107 ( .B1(n10025), .B2(keyinput103), .C1(n10193), .C2(
        keyinput53), .A(n10024), .ZN(n10035) );
  INV_X1 U11108 ( .A(SI_24_), .ZN(n10027) );
  AOI22_X1 U11109 ( .A1(n9311), .A2(keyinput85), .B1(n10027), .B2(keyinput86), 
        .ZN(n10026) );
  OAI221_X1 U11110 ( .B1(n9311), .B2(keyinput85), .C1(n10027), .C2(keyinput86), 
        .A(n10026), .ZN(n10034) );
  AOI22_X1 U11111 ( .A1(n5251), .A2(keyinput16), .B1(n10029), .B2(keyinput44), 
        .ZN(n10028) );
  OAI221_X1 U11112 ( .B1(n5251), .B2(keyinput16), .C1(n10029), .C2(keyinput44), 
        .A(n10028), .ZN(n10033) );
  XNOR2_X1 U11113 ( .A(P1_REG3_REG_16__SCAN_IN), .B(keyinput78), .ZN(n10031)
         );
  XNOR2_X1 U11114 ( .A(SI_1_), .B(keyinput48), .ZN(n10030) );
  NAND2_X1 U11115 ( .A1(n10031), .A2(n10030), .ZN(n10032) );
  NOR4_X1 U11116 ( .A1(n10035), .A2(n10034), .A3(n10033), .A4(n10032), .ZN(
        n10046) );
  AOI22_X1 U11117 ( .A1(n6928), .A2(keyinput26), .B1(n5158), .B2(keyinput124), 
        .ZN(n10036) );
  OAI221_X1 U11118 ( .B1(n6928), .B2(keyinput26), .C1(n5158), .C2(keyinput124), 
        .A(n10036), .ZN(n10044) );
  AOI22_X1 U11119 ( .A1(n10171), .A2(keyinput19), .B1(keyinput91), .B2(n10170), 
        .ZN(n10037) );
  OAI221_X1 U11120 ( .B1(n10171), .B2(keyinput19), .C1(n10170), .C2(keyinput91), .A(n10037), .ZN(n10043) );
  AOI22_X1 U11121 ( .A1(n10039), .A2(keyinput87), .B1(n10169), .B2(keyinput42), 
        .ZN(n10038) );
  OAI221_X1 U11122 ( .B1(n10039), .B2(keyinput87), .C1(n10169), .C2(keyinput42), .A(n10038), .ZN(n10042) );
  AOI22_X1 U11123 ( .A1(n10174), .A2(keyinput32), .B1(n10175), .B2(keyinput127), .ZN(n10040) );
  OAI221_X1 U11124 ( .B1(n10174), .B2(keyinput32), .C1(n10175), .C2(
        keyinput127), .A(n10040), .ZN(n10041) );
  NOR4_X1 U11125 ( .A1(n10044), .A2(n10043), .A3(n10042), .A4(n10041), .ZN(
        n10045) );
  NAND4_X1 U11126 ( .A1(n10048), .A2(n10047), .A3(n10046), .A4(n10045), .ZN(
        n10101) );
  AOI22_X1 U11127 ( .A1(n10172), .A2(keyinput101), .B1(keyinput10), .B2(n5141), 
        .ZN(n10049) );
  OAI221_X1 U11128 ( .B1(n10172), .B2(keyinput101), .C1(n5141), .C2(keyinput10), .A(n10049), .ZN(n10058) );
  AOI22_X1 U11129 ( .A1(n10051), .A2(keyinput111), .B1(n6412), .B2(keyinput120), .ZN(n10050) );
  OAI221_X1 U11130 ( .B1(n10051), .B2(keyinput111), .C1(n6412), .C2(
        keyinput120), .A(n10050), .ZN(n10057) );
  AOI22_X1 U11131 ( .A1(n7229), .A2(keyinput107), .B1(n5917), .B2(keyinput51), 
        .ZN(n10052) );
  OAI221_X1 U11132 ( .B1(n7229), .B2(keyinput107), .C1(n5917), .C2(keyinput51), 
        .A(n10052), .ZN(n10056) );
  XNOR2_X1 U11133 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(keyinput74), .ZN(n10054)
         );
  XNOR2_X1 U11134 ( .A(P2_REG0_REG_20__SCAN_IN), .B(keyinput75), .ZN(n10053)
         );
  NAND2_X1 U11135 ( .A1(n10054), .A2(n10053), .ZN(n10055) );
  NOR4_X1 U11136 ( .A1(n10058), .A2(n10057), .A3(n10056), .A4(n10055), .ZN(
        n10099) );
  INV_X1 U11137 ( .A(SI_5_), .ZN(n10061) );
  AOI22_X1 U11138 ( .A1(n10061), .A2(keyinput8), .B1(keyinput109), .B2(n10060), 
        .ZN(n10059) );
  OAI221_X1 U11139 ( .B1(n10061), .B2(keyinput8), .C1(n10060), .C2(keyinput109), .A(n10059), .ZN(n10071) );
  AOI22_X1 U11140 ( .A1(n10064), .A2(keyinput90), .B1(n10063), .B2(keyinput4), 
        .ZN(n10062) );
  OAI221_X1 U11141 ( .B1(n10064), .B2(keyinput90), .C1(n10063), .C2(keyinput4), 
        .A(n10062), .ZN(n10070) );
  AOI22_X1 U11142 ( .A1(n10178), .A2(keyinput116), .B1(keyinput11), .B2(n10176), .ZN(n10065) );
  OAI221_X1 U11143 ( .B1(n10178), .B2(keyinput116), .C1(n10176), .C2(
        keyinput11), .A(n10065), .ZN(n10069) );
  XNOR2_X1 U11144 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput46), .ZN(n10067) );
  XNOR2_X1 U11145 ( .A(P2_IR_REG_27__SCAN_IN), .B(keyinput38), .ZN(n10066) );
  NAND2_X1 U11146 ( .A1(n10067), .A2(n10066), .ZN(n10068) );
  NOR4_X1 U11147 ( .A1(n10071), .A2(n10070), .A3(n10069), .A4(n10068), .ZN(
        n10098) );
  AOI22_X1 U11148 ( .A1(n5117), .A2(keyinput62), .B1(keyinput81), .B2(n5568), 
        .ZN(n10072) );
  OAI221_X1 U11149 ( .B1(n5117), .B2(keyinput62), .C1(n5568), .C2(keyinput81), 
        .A(n10072), .ZN(n10082) );
  AOI22_X1 U11150 ( .A1(n10075), .A2(keyinput5), .B1(keyinput2), .B2(n10074), 
        .ZN(n10073) );
  OAI221_X1 U11151 ( .B1(n10075), .B2(keyinput5), .C1(n10074), .C2(keyinput2), 
        .A(n10073), .ZN(n10081) );
  INV_X1 U11152 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n10164) );
  AOI22_X1 U11153 ( .A1(n9618), .A2(keyinput61), .B1(n10164), .B2(keyinput21), 
        .ZN(n10076) );
  OAI221_X1 U11154 ( .B1(n9618), .B2(keyinput61), .C1(n10164), .C2(keyinput21), 
        .A(n10076), .ZN(n10080) );
  INV_X1 U11155 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n10162) );
  AOI22_X1 U11156 ( .A1(n10162), .A2(keyinput98), .B1(n10078), .B2(keyinput15), 
        .ZN(n10077) );
  OAI221_X1 U11157 ( .B1(n10162), .B2(keyinput98), .C1(n10078), .C2(keyinput15), .A(n10077), .ZN(n10079) );
  NOR4_X1 U11158 ( .A1(n10082), .A2(n10081), .A3(n10080), .A4(n10079), .ZN(
        n10097) );
  INV_X1 U11159 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n10163) );
  AOI22_X1 U11160 ( .A1(n10084), .A2(keyinput125), .B1(keyinput56), .B2(n10163), .ZN(n10083) );
  OAI221_X1 U11161 ( .B1(n10084), .B2(keyinput125), .C1(n10163), .C2(
        keyinput56), .A(n10083), .ZN(n10095) );
  AOI22_X1 U11162 ( .A1(n10087), .A2(keyinput84), .B1(n10086), .B2(keyinput41), 
        .ZN(n10085) );
  OAI221_X1 U11163 ( .B1(n10087), .B2(keyinput84), .C1(n10086), .C2(keyinput41), .A(n10085), .ZN(n10094) );
  AOI22_X1 U11164 ( .A1(n10089), .A2(keyinput76), .B1(n10161), .B2(keyinput25), 
        .ZN(n10088) );
  OAI221_X1 U11165 ( .B1(n10089), .B2(keyinput76), .C1(n10161), .C2(keyinput25), .A(n10088), .ZN(n10093) );
  XNOR2_X1 U11166 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput89), .ZN(n10091) );
  XNOR2_X1 U11167 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput67), .ZN(n10090)
         );
  NAND2_X1 U11168 ( .A1(n10091), .A2(n10090), .ZN(n10092) );
  NOR4_X1 U11169 ( .A1(n10095), .A2(n10094), .A3(n10093), .A4(n10092), .ZN(
        n10096) );
  NAND4_X1 U11170 ( .A1(n10099), .A2(n10098), .A3(n10097), .A4(n10096), .ZN(
        n10100) );
  NOR4_X1 U11171 ( .A1(n10103), .A2(n10102), .A3(n10101), .A4(n10100), .ZN(
        n10104) );
  XNOR2_X1 U11172 ( .A(n10105), .B(n10104), .ZN(n10192) );
  NOR2_X1 U11173 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), 
        .ZN(n10125) );
  OR4_X1 U11174 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(n10106), .A3(n5850), .A4(
        n5917), .ZN(n10122) );
  NOR4_X1 U11175 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .A3(
        P2_ADDR_REG_16__SCAN_IN), .A4(P2_ADDR_REG_14__SCAN_IN), .ZN(n10116) );
  NOR4_X1 U11176 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .A3(n10108), .A4(n10107), .ZN(n10115) );
  NOR4_X1 U11177 ( .A1(SI_12_), .A2(P1_REG2_REG_0__SCAN_IN), .A3(n10110), .A4(
        n10109), .ZN(n10114) );
  NOR4_X1 U11178 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_22__SCAN_IN), 
        .A3(n10112), .A4(n10111), .ZN(n10113) );
  NAND4_X1 U11179 ( .A1(n10116), .A2(n10115), .A3(n10114), .A4(n10113), .ZN(
        n10121) );
  NAND4_X1 U11180 ( .A1(n10119), .A2(n10118), .A3(n10117), .A4(
        P1_IR_REG_16__SCAN_IN), .ZN(n10120) );
  NOR3_X1 U11181 ( .A1(n10122), .A2(n10121), .A3(n10120), .ZN(n10123) );
  NAND4_X1 U11182 ( .A1(n10126), .A2(n10125), .A3(n10124), .A4(n10123), .ZN(
        n10190) );
  OR4_X1 U11183 ( .A1(SI_21_), .A2(SI_10_), .A3(P1_REG0_REG_2__SCAN_IN), .A4(
        n10127), .ZN(n10133) );
  NOR4_X1 U11184 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(P1_DATAO_REG_20__SCAN_IN), .A3(P2_IR_REG_6__SCAN_IN), .A4(P2_REG0_REG_6__SCAN_IN), .ZN(n10128) );
  NAND3_X1 U11185 ( .A1(n9942), .A2(n10129), .A3(n10128), .ZN(n10130) );
  NOR4_X1 U11186 ( .A1(n10133), .A2(n10132), .A3(n10131), .A4(n10130), .ZN(
        n10136) );
  NOR4_X1 U11187 ( .A1(SI_0_), .A2(P2_REG3_REG_14__SCAN_IN), .A3(
        P2_IR_REG_30__SCAN_IN), .A4(n10134), .ZN(n10135) );
  NAND2_X1 U11188 ( .A1(n10136), .A2(n10135), .ZN(n10189) );
  NAND4_X1 U11189 ( .A1(P2_D_REG_31__SCAN_IN), .A2(SI_31_), .A3(n5068), .A4(
        n6067), .ZN(n10143) );
  NAND4_X1 U11190 ( .A1(P1_REG2_REG_26__SCAN_IN), .A2(P2_REG2_REG_15__SCAN_IN), 
        .A3(n10137), .A4(n6871), .ZN(n10142) );
  NAND4_X1 U11191 ( .A1(P1_RD_REG_SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_REG2_REG_6__SCAN_IN), .A4(n10138), .ZN(n10141) );
  NAND4_X1 U11192 ( .A1(n10139), .A2(P1_REG2_REG_29__SCAN_IN), .A3(
        P2_REG2_REG_29__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n10140) );
  OR4_X1 U11193 ( .A1(n10143), .A2(n10142), .A3(n10141), .A4(n10140), .ZN(
        n10188) );
  NAND4_X1 U11194 ( .A1(SI_25_), .A2(n8816), .A3(n10144), .A4(n6879), .ZN(
        n10149) );
  NAND4_X1 U11195 ( .A1(P1_B_REG_SCAN_IN), .A2(n7305), .A3(n10145), .A4(n7791), 
        .ZN(n10148) );
  NAND4_X1 U11196 ( .A1(P2_D_REG_21__SCAN_IN), .A2(SI_1_), .A3(
        P2_REG1_REG_13__SCAN_IN), .A4(n5251), .ZN(n10147) );
  NAND4_X1 U11197 ( .A1(SI_24_), .A2(P1_REG2_REG_21__SCAN_IN), .A3(
        P2_REG3_REG_28__SCAN_IN), .A4(P2_REG1_REG_4__SCAN_IN), .ZN(n10146) );
  NOR4_X1 U11198 ( .A1(n10149), .A2(n10148), .A3(n10147), .A4(n10146), .ZN(
        n10186) );
  NAND4_X1 U11199 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .A3(P2_REG1_REG_28__SCAN_IN), .A4(n10150), .ZN(n10159) );
  NAND4_X1 U11200 ( .A1(P2_DATAO_REG_5__SCAN_IN), .A2(P1_REG1_REG_9__SCAN_IN), 
        .A3(n10152), .A4(n10151), .ZN(n10158) );
  NAND4_X1 U11201 ( .A1(P1_REG2_REG_27__SCAN_IN), .A2(P2_B_REG_SCAN_IN), .A3(
        P2_REG1_REG_1__SCAN_IN), .A4(n10153), .ZN(n10157) );
  NAND4_X1 U11202 ( .A1(P1_REG1_REG_13__SCAN_IN), .A2(P1_REG1_REG_12__SCAN_IN), 
        .A3(n10155), .A4(n10154), .ZN(n10156) );
  NOR4_X1 U11203 ( .A1(n10159), .A2(n10158), .A3(n10157), .A4(n10156), .ZN(
        n10185) );
  NAND4_X1 U11204 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), 
        .A3(P2_REG2_REG_25__SCAN_IN), .A4(n5117), .ZN(n10168) );
  NAND4_X1 U11205 ( .A1(P1_D_REG_4__SCAN_IN), .A2(SI_19_), .A3(SI_5_), .A4(
        P2_REG1_REG_0__SCAN_IN), .ZN(n10167) );
  NAND4_X1 U11206 ( .A1(P1_REG2_REG_24__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), 
        .A3(n10161), .A4(n10160), .ZN(n10166) );
  NAND4_X1 U11207 ( .A1(P1_REG0_REG_4__SCAN_IN), .A2(n10164), .A3(n10163), 
        .A4(n10162), .ZN(n10165) );
  NOR4_X1 U11208 ( .A1(n10168), .A2(n10167), .A3(n10166), .A4(n10165), .ZN(
        n10184) );
  NAND4_X1 U11209 ( .A1(P2_REG0_REG_27__SCAN_IN), .A2(n10171), .A3(n10170), 
        .A4(n10169), .ZN(n10182) );
  NAND4_X1 U11210 ( .A1(P1_REG1_REG_14__SCAN_IN), .A2(n5141), .A3(n10172), 
        .A4(n7229), .ZN(n10181) );
  NAND4_X1 U11211 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(n10175), .A3(n10174), 
        .A4(n10173), .ZN(n10180) );
  NAND4_X1 U11212 ( .A1(n10178), .A2(n10177), .A3(n10176), .A4(
        P2_IR_REG_31__SCAN_IN), .ZN(n10179) );
  NOR4_X1 U11213 ( .A1(n10182), .A2(n10181), .A3(n10180), .A4(n10179), .ZN(
        n10183) );
  NAND4_X1 U11214 ( .A1(n10186), .A2(n10185), .A3(n10184), .A4(n10183), .ZN(
        n10187) );
  NOR4_X1 U11215 ( .A1(n10190), .A2(n10189), .A3(n10188), .A4(n10187), .ZN(
        n10191) );
  XNOR2_X1 U11216 ( .A(n10192), .B(n10191), .ZN(P1_U3578) );
  XNOR2_X1 U11217 ( .A(n10194), .B(n10193), .ZN(ADD_1071_U49) );
  XOR2_X1 U11218 ( .A(n10195), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11219 ( .A1(n10197), .A2(n10196), .ZN(n10198) );
  XOR2_X1 U11220 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10198), .Z(ADD_1071_U51) );
  OAI21_X1 U11221 ( .B1(n10201), .B2(n10200), .A(n10199), .ZN(n10202) );
  XNOR2_X1 U11222 ( .A(n10202), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11223 ( .B1(n10205), .B2(n10204), .A(n10203), .ZN(ADD_1071_U47) );
  XNOR2_X1 U11224 ( .A(n10206), .B(n9618), .ZN(ADD_1071_U48) );
  XOR2_X1 U11225 ( .A(n10208), .B(n10207), .Z(ADD_1071_U54) );
  XOR2_X1 U11226 ( .A(n10210), .B(n10209), .Z(ADD_1071_U53) );
  XNOR2_X1 U11227 ( .A(n10212), .B(n10211), .ZN(ADD_1071_U52) );
  INV_X2 U5072 ( .A(n4386), .ZN(n5797) );
  CLKBUF_X1 U4893 ( .A(n5964), .Z(n4386) );
  CLKBUF_X1 U4899 ( .A(n6850), .Z(n8101) );
  CLKBUF_X1 U4917 ( .A(n8714), .Z(n4385) );
  CLKBUF_X1 U4928 ( .A(n5213), .Z(n6195) );
endmodule

