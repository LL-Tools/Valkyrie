

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4378, n4379, n4380, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10279;

  AND2_X1 U4881 ( .A1(n8208), .A2(n8402), .ZN(n8394) );
  NAND2_X1 U4882 ( .A1(n6071), .A2(n6070), .ZN(n8696) );
  INV_X2 U4883 ( .A(n5057), .ZN(n5791) );
  XNOR2_X1 U4884 ( .A(n5830), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5837) );
  INV_X1 U4886 ( .A(n8163), .ZN(n8152) );
  OR2_X1 U4887 ( .A1(n7185), .A2(n7384), .ZN(n7396) );
  OAI21_X1 U4888 ( .B1(n6076), .B2(n4732), .A(n4734), .ZN(n8522) );
  OR2_X1 U4889 ( .A1(n7931), .A2(n7764), .ZN(n6278) );
  AND2_X1 U4890 ( .A1(n4799), .A2(n9109), .ZN(n9255) );
  INV_X1 U4891 ( .A(n6975), .ZN(n6718) );
  INV_X1 U4892 ( .A(n8148), .ZN(n8162) );
  AND2_X1 U4893 ( .A1(n6316), .A2(n6313), .ZN(n8539) );
  BUF_X1 U4894 ( .A(n5058), .Z(n5534) );
  AND3_X1 U4895 ( .A1(n5027), .A2(n5026), .A3(n4599), .ZN(n6975) );
  NAND2_X1 U4896 ( .A1(n5990), .A2(n5989), .ZN(n7931) );
  NAND2_X1 U4897 ( .A1(n5976), .A2(n5975), .ZN(n7823) );
  AND2_X1 U4898 ( .A1(n4489), .A2(n6873), .ZN(n9868) );
  INV_X2 U4899 ( .A(n5091), .ZN(n5634) );
  AND3_X1 U4900 ( .A1(n6397), .A2(n4539), .A3(n4538), .ZN(n6420) );
  MUX2_X1 U4901 ( .A(n9150), .B(n9149), .S(n9148), .Z(n9155) );
  OAI22_X2 U4903 ( .A1(n7993), .A2(n7992), .B1(n8716), .B2(n8316), .ZN(n7994)
         );
  NAND2_X2 U4904 ( .A1(n4602), .A2(n4992), .ZN(n5798) );
  AOI22_X2 U4907 ( .A1(n8823), .A2(n4889), .B1(n4888), .B2(n4891), .ZN(n4887)
         );
  OAI21_X2 U4908 ( .B1(n8762), .B2(n8764), .A(n8761), .ZN(n8823) );
  NOR2_X2 U4909 ( .A1(n8674), .A2(n8515), .ZN(n8499) );
  AOI211_X2 U4910 ( .C1(n9564), .C2(n9563), .A(n9562), .B(n9561), .ZN(n9584)
         );
  AND2_X4 U4914 ( .A1(n8180), .A2(n8749), .ZN(n5915) );
  NAND2_X1 U4915 ( .A1(n4652), .A2(n4996), .ZN(n4380) );
  NAND2_X1 U4916 ( .A1(n4652), .A2(n4996), .ZN(n6466) );
  NAND2_X1 U4917 ( .A1(n4473), .A2(n4790), .ZN(n9285) );
  NAND2_X1 U4918 ( .A1(n9336), .A2(n9335), .ZN(n9334) );
  INV_X1 U4919 ( .A(n9168), .ZN(n7478) );
  INV_X2 U4920 ( .A(n7246), .ZN(n7436) );
  NAND2_X1 U4921 ( .A1(n5777), .A2(n7489), .ZN(n6982) );
  NAND2_X1 U4922 ( .A1(n4994), .A2(n4995), .ZN(n6688) );
  NAND2_X1 U4923 ( .A1(n5011), .A2(n5010), .ZN(n9317) );
  INV_X1 U4924 ( .A(n5837), .ZN(n8180) );
  INV_X2 U4925 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NOR2_X1 U4926 ( .A1(n9451), .A2(n4924), .ZN(n9452) );
  AOI211_X1 U4927 ( .C1(n9414), .C2(n9461), .A(n8134), .B(n8133), .ZN(n8135)
         );
  OAI21_X1 U4928 ( .B1(n9069), .B2(n9136), .A(n4587), .ZN(n4586) );
  AOI21_X1 U4929 ( .B1(n4469), .B2(n4799), .A(n4467), .ZN(n9463) );
  NOR2_X1 U4930 ( .A1(n9285), .A2(n9284), .ZN(n9283) );
  AOI211_X1 U4931 ( .C1(n9868), .C2(n9557), .A(n9556), .B(n9555), .ZN(n9559)
         );
  OR2_X1 U4932 ( .A1(n4936), .A2(n4750), .ZN(n4749) );
  AOI21_X1 U4933 ( .B1(n8226), .B2(n8223), .A(n8225), .ZN(n8145) );
  NOR2_X1 U4934 ( .A1(n4890), .A2(n5706), .ZN(n4889) );
  NAND2_X1 U4935 ( .A1(n8276), .A2(n4922), .ZN(n8144) );
  XNOR2_X1 U4936 ( .A(n6216), .B(n6215), .ZN(n9545) );
  NAND2_X1 U4937 ( .A1(n6175), .A2(n6174), .ZN(n8641) );
  NAND2_X1 U4938 ( .A1(n5719), .A2(n5718), .ZN(n9460) );
  OAI21_X1 U4939 ( .B1(n6201), .B2(n6200), .A(n6199), .ZN(n6211) );
  XNOR2_X1 U4940 ( .A(n6184), .B(n6183), .ZN(n8007) );
  NAND2_X1 U4941 ( .A1(n5250), .A2(n5249), .ZN(n7653) );
  OAI21_X1 U4942 ( .B1(n4783), .B2(n4780), .A(n4778), .ZN(n8127) );
  NAND2_X1 U4943 ( .A1(n5636), .A2(n5635), .ZN(n9478) );
  NAND2_X1 U4944 ( .A1(n7809), .A2(n8999), .ZN(n7851) );
  NAND2_X1 U4945 ( .A1(n4404), .A2(n6316), .ZN(n4736) );
  OR2_X1 U4946 ( .A1(n9486), .A2(n9337), .ZN(n8117) );
  NAND2_X1 U4947 ( .A1(n6098), .A2(n6097), .ZN(n8679) );
  OAI21_X1 U4948 ( .B1(n7590), .B2(n8987), .A(n8981), .ZN(n7613) );
  NAND2_X1 U4949 ( .A1(n6079), .A2(n6078), .ZN(n8693) );
  OR2_X1 U4950 ( .A1(n8686), .A2(n8555), .ZN(n6316) );
  NAND2_X1 U4951 ( .A1(n5509), .A2(n5508), .ZN(n9501) );
  NAND2_X1 U4952 ( .A1(n4474), .A2(n8924), .ZN(n7590) );
  AND2_X1 U4953 ( .A1(n6298), .A2(n6293), .ZN(n8587) );
  OR2_X1 U4954 ( .A1(n8703), .A2(n8618), .ZN(n6298) );
  NAND2_X1 U4955 ( .A1(n5480), .A2(n5479), .ZN(n9509) );
  NOR3_X2 U4956 ( .A1(n7685), .A2(n8711), .A3(n4644), .ZN(n4641) );
  NAND2_X1 U4957 ( .A1(n6059), .A2(n6058), .ZN(n8703) );
  AND2_X1 U4958 ( .A1(n6287), .A2(n6286), .ZN(n7992) );
  NAND2_X1 U4959 ( .A1(n6035), .A2(n6034), .ZN(n8711) );
  NAND2_X1 U4960 ( .A1(n5264), .A2(n5263), .ZN(n7664) );
  NAND2_X1 U4961 ( .A1(n5953), .A2(n5952), .ZN(n7840) );
  NAND2_X1 U4962 ( .A1(n9817), .A2(n9808), .ZN(n8626) );
  INV_X2 U4963 ( .A(n9817), .ZN(n8600) );
  AND2_X2 U4964 ( .A1(n7290), .A2(n9425), .ZN(n9404) );
  OAI21_X1 U4965 ( .B1(n4664), .B2(n4388), .A(n5283), .ZN(n5309) );
  OAI21_X1 U4966 ( .B1(n5222), .B2(n5221), .A(n5223), .ZN(n5251) );
  INV_X1 U4967 ( .A(n6924), .ZN(n9807) );
  AND2_X1 U4968 ( .A1(n5914), .A2(n4528), .ZN(n6924) );
  AND2_X2 U4969 ( .A1(n6690), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  NAND2_X1 U4970 ( .A1(n5154), .A2(n5153), .ZN(n5176) );
  CLKBUF_X3 U4971 ( .A(n5028), .Z(n5753) );
  OAI211_X1 U4972 ( .C1(n5155), .C2(n6478), .A(n5129), .B(n5128), .ZN(n7213)
         );
  AND2_X1 U4973 ( .A1(n6982), .A2(n5000), .ZN(n5028) );
  NAND4_X2 U4974 ( .A1(n5022), .A2(n5021), .A3(n5020), .A4(n5019), .ZN(n6974)
         );
  CLKBUF_X1 U4975 ( .A(n5000), .Z(n6430) );
  INV_X1 U4976 ( .A(n4384), .ZN(n4386) );
  OAI21_X1 U4977 ( .B1(n5069), .B2(n4999), .A(n4998), .ZN(n7348) );
  CLKBUF_X1 U4978 ( .A(n5776), .Z(n9071) );
  AND2_X2 U4979 ( .A1(n4962), .A2(n4961), .ZN(n5098) );
  AND2_X1 U4980 ( .A1(n7489), .A2(n9317), .ZN(n5787) );
  AND3_X1 U4981 ( .A1(n5090), .A2(n4788), .A3(n4786), .ZN(n5122) );
  INV_X1 U4982 ( .A(n8220), .ZN(n4961) );
  XNOR2_X1 U4983 ( .A(n5005), .B(n5004), .ZN(n5776) );
  XNOR2_X1 U4984 ( .A(n4988), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5770) );
  NAND2_X1 U4985 ( .A1(n4987), .A2(n4983), .ZN(n7944) );
  NAND2_X2 U4986 ( .A1(n6851), .A2(n6850), .ZN(n8163) );
  AND2_X1 U4987 ( .A1(n4976), .A2(n5003), .ZN(n5777) );
  NAND2_X1 U4988 ( .A1(n6557), .A2(n5091), .ZN(n5921) );
  AND2_X2 U4989 ( .A1(n8180), .A2(n5849), .ZN(n6179) );
  NAND2_X1 U4990 ( .A1(n5003), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5005) );
  NAND2_X1 U4991 ( .A1(n4987), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4988) );
  NAND2_X1 U4992 ( .A1(n4603), .A2(n4991), .ZN(n4602) );
  XNOR2_X1 U4993 ( .A(n4986), .B(n4985), .ZN(n7839) );
  NAND2_X1 U4994 ( .A1(n4959), .A2(n4958), .ZN(n8047) );
  NAND2_X1 U4995 ( .A1(n4981), .A2(n4980), .ZN(n4987) );
  NAND2_X1 U4996 ( .A1(n4958), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4956) );
  OAI21_X1 U4997 ( .B1(n4993), .B2(n9546), .A(P1_IR_REG_28__SCAN_IN), .ZN(
        n4603) );
  OR2_X1 U4998 ( .A1(n4979), .A2(n9546), .ZN(n4981) );
  MUX2_X1 U4999 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5856), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n5859) );
  AND2_X1 U5000 ( .A1(n4971), .A2(n4972), .ZN(n5006) );
  XNOR2_X1 U5001 ( .A(n5073), .B(P1_IR_REG_3__SCAN_IN), .ZN(n8061) );
  AND2_X1 U5002 ( .A1(n4544), .A2(n4543), .ZN(n5083) );
  XNOR2_X1 U5003 ( .A(n5862), .B(n5861), .ZN(n8212) );
  INV_X2 U5004 ( .A(n9954), .ZN(n8747) );
  NAND2_X2 U5005 ( .A1(n5634), .A2(P1_U3084), .ZN(n9550) );
  AND4_X1 U5006 ( .A1(n4864), .A2(n5844), .A3(n5845), .A4(n4776), .ZN(n5854)
         );
  AND4_X1 U5007 ( .A1(n6401), .A2(n4863), .A3(n5827), .A4(n5825), .ZN(n4864)
         );
  NAND2_X1 U5008 ( .A1(n4990), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4991) );
  AND3_X1 U5009 ( .A1(n6409), .A2(n6398), .A3(n6412), .ZN(n6401) );
  AND2_X1 U5010 ( .A1(n5828), .A2(n5861), .ZN(n4776) );
  AND4_X1 U5011 ( .A1(n5823), .A2(n5822), .A3(n5821), .A4(n5820), .ZN(n5845)
         );
  NOR2_X1 U5012 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4942) );
  INV_X1 U5013 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n4972) );
  INV_X1 U5014 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6412) );
  INV_X1 U5015 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6409) );
  INV_X1 U5016 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6398) );
  INV_X1 U5017 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4955) );
  INV_X1 U5018 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5260) );
  INV_X1 U5019 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5004) );
  INV_X1 U5020 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10225) );
  INV_X1 U5021 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n10138) );
  INV_X1 U5022 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5229) );
  INV_X1 U5023 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5365) );
  NOR2_X1 U5024 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5863) );
  INV_X1 U5025 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9214) );
  NOR2_X2 U5026 ( .A1(n8445), .A2(n8652), .ZN(n4647) );
  AND2_X2 U5027 ( .A1(n4971), .A2(n4951), .ZN(n5771) );
  NOR2_X4 U5028 ( .A1(n5227), .A2(n4945), .ZN(n4971) );
  XNOR2_X2 U5029 ( .A(n6974), .B(n6975), .ZN(n9077) );
  OAI21_X2 U5030 ( .B1(n7653), .B2(n5276), .A(n5275), .ZN(n7786) );
  INV_X1 U5031 ( .A(n7211), .ZN(n4382) );
  INV_X1 U5032 ( .A(n4382), .ZN(n4383) );
  NOR3_X2 U5033 ( .A1(n7599), .A2(n4606), .A3(n9524), .ZN(n7856) );
  NAND2_X1 U5034 ( .A1(n5406), .A2(n5380), .ZN(n8026) );
  NOR2_X2 U5035 ( .A1(n7253), .A2(n9807), .ZN(n7256) );
  NAND2_X1 U5036 ( .A1(n4640), .A2(n7085), .ZN(n7253) );
  INV_X4 U5037 ( .A(n5629), .ZN(n5747) );
  INV_X1 U5038 ( .A(n6852), .ZN(n4384) );
  INV_X1 U5039 ( .A(n4384), .ZN(n4385) );
  AND2_X1 U5040 ( .A1(n9557), .A2(n4650), .ZN(n6351) );
  INV_X1 U5041 ( .A(n8311), .ZN(n4650) );
  OR2_X1 U5042 ( .A1(n8438), .A2(n6160), .ZN(n6166) );
  NAND2_X1 U5043 ( .A1(n4547), .A2(n6298), .ZN(n4546) );
  INV_X1 U5044 ( .A(n4548), .ZN(n4547) );
  AOI21_X1 U5045 ( .B1(n6297), .B2(n6296), .A(n8187), .ZN(n4548) );
  INV_X1 U5046 ( .A(n8992), .ZN(n4584) );
  INV_X1 U5047 ( .A(n4575), .ZN(n4568) );
  AND2_X1 U5048 ( .A1(n4573), .A2(n9011), .ZN(n4572) );
  NAND2_X1 U5049 ( .A1(n6307), .A2(n6345), .ZN(n4559) );
  AND2_X1 U5050 ( .A1(n4951), .A2(n4405), .ZN(n4560) );
  INV_X1 U5051 ( .A(n7870), .ZN(n4810) );
  INV_X1 U5052 ( .A(n6332), .ZN(n4756) );
  OR2_X1 U5053 ( .A1(n8674), .A2(n8229), .ZN(n6304) );
  OR2_X1 U5054 ( .A1(n8716), .A2(n7991), .ZN(n6287) );
  OR2_X1 U5055 ( .A1(n8711), .A2(n8616), .ZN(n6290) );
  OAI21_X1 U5056 ( .B1(n6878), .B2(n6835), .A(n6836), .ZN(n6959) );
  INV_X1 U5057 ( .A(n6882), .ZN(n6835) );
  AOI21_X1 U5058 ( .B1(n9820), .B2(n6809), .A(n6808), .ZN(n7008) );
  INV_X1 U5059 ( .A(n7976), .ZN(n6806) );
  INV_X1 U5060 ( .A(n8047), .ZN(n4962) );
  AND2_X1 U5061 ( .A1(n9450), .A2(n9156), .ZN(n9060) );
  OR2_X1 U5062 ( .A1(n9455), .A2(n9242), .ZN(n9074) );
  NAND2_X1 U5063 ( .A1(n5688), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5739) );
  INV_X1 U5064 ( .A(n5690), .ZN(n5688) );
  OR2_X1 U5065 ( .A1(n9478), .A2(n8767), .ZN(n9132) );
  OR2_X1 U5066 ( .A1(n9486), .A2(n9370), .ZN(n9035) );
  XNOR2_X1 U5067 ( .A(n6211), .B(n6210), .ZN(n6208) );
  NAND2_X1 U5068 ( .A1(n4688), .A2(n4687), .ZN(n6201) );
  AOI21_X1 U5069 ( .B1(n4689), .B2(n4691), .A(n4456), .ZN(n4687) );
  NAND2_X1 U5070 ( .A1(n5716), .A2(n4689), .ZN(n4688) );
  AOI21_X1 U5071 ( .B1(n4695), .B2(n4397), .A(n4694), .ZN(n4693) );
  INV_X1 U5072 ( .A(n4659), .ZN(n5362) );
  AOI21_X1 U5073 ( .B1(n5251), .B2(n4661), .A(n4660), .ZN(n4659) );
  OAI21_X1 U5074 ( .B1(n4662), .B2(n4667), .A(n5337), .ZN(n4660) );
  NAND2_X1 U5075 ( .A1(n6393), .A2(n4830), .ZN(n6851) );
  NOR2_X1 U5076 ( .A1(n9812), .A2(n7581), .ZN(n4830) );
  AND2_X1 U5077 ( .A1(n6393), .A2(n7581), .ZN(n6862) );
  XNOR2_X1 U5078 ( .A(n6226), .B(n6225), .ZN(n7010) );
  OAI21_X1 U5079 ( .B1(n6363), .B2(n4657), .A(n4655), .ZN(n6395) );
  NAND2_X1 U5080 ( .A1(n4656), .A2(n4416), .ZN(n4655) );
  OR2_X1 U5081 ( .A1(n8652), .A2(n8423), .ZN(n8200) );
  AND2_X1 U5082 ( .A1(n6153), .A2(n4775), .ZN(n4774) );
  OR2_X1 U5083 ( .A1(n8662), .A2(n8254), .ZN(n6228) );
  NAND2_X1 U5084 ( .A1(n8468), .A2(n8450), .ZN(n8445) );
  OR2_X1 U5085 ( .A1(n4880), .A2(n4878), .ZN(n4877) );
  INV_X1 U5086 ( .A(n8198), .ZN(n4878) );
  NAND2_X1 U5087 ( .A1(n8198), .A2(n8498), .ZN(n4879) );
  OR2_X1 U5088 ( .A1(n8674), .A2(n8525), .ZN(n4881) );
  OAI211_X1 U5089 ( .C1(n4845), .C2(n4841), .A(n8194), .B(n4839), .ZN(n8196)
         );
  OAI21_X1 U5090 ( .B1(n7707), .B2(n4873), .A(n4871), .ZN(n7679) );
  INV_X1 U5091 ( .A(n4872), .ZN(n4871) );
  NAND2_X1 U5092 ( .A1(n7707), .A2(n4400), .ZN(n7677) );
  NAND2_X1 U5093 ( .A1(n7632), .A2(n7631), .ZN(n7709) );
  NAND2_X1 U5094 ( .A1(n6825), .A2(n6824), .ZN(n8585) );
  NAND2_X1 U5095 ( .A1(n5831), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5830) );
  INV_X1 U5096 ( .A(n9338), .ZN(n8767) );
  INV_X1 U5097 ( .A(n5155), .ZN(n4601) );
  AND2_X1 U5098 ( .A1(n5013), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n5014) );
  NAND2_X1 U5099 ( .A1(n5002), .A2(n5001), .ZN(n4516) );
  OR2_X1 U5100 ( .A1(n9445), .A2(n9219), .ZN(n9139) );
  INV_X1 U5101 ( .A(n5142), .ZN(n5792) );
  XNOR2_X1 U5102 ( .A(n4499), .B(n4498), .ZN(n9211) );
  INV_X1 U5103 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n4498) );
  NOR2_X1 U5104 ( .A1(n9740), .A2(n4500), .ZN(n4499) );
  AND2_X1 U5105 ( .A1(n9205), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4500) );
  NAND2_X1 U5106 ( .A1(n9268), .A2(n9250), .ZN(n9246) );
  NAND2_X1 U5107 ( .A1(n9292), .A2(n4720), .ZN(n4719) );
  NOR2_X1 U5108 ( .A1(n4721), .A2(n8124), .ZN(n4720) );
  INV_X1 U5109 ( .A(n8122), .ZN(n4721) );
  AOI21_X1 U5110 ( .B1(n4724), .B2(n4728), .A(n4426), .ZN(n4723) );
  NAND2_X1 U5111 ( .A1(n7851), .A2(n4784), .ZN(n4783) );
  AND2_X1 U5112 ( .A1(n9013), .A2(n9004), .ZN(n4784) );
  NAND2_X1 U5113 ( .A1(n4717), .A2(n4715), .ZN(n7979) );
  INV_X1 U5114 ( .A(n4716), .ZN(n4715) );
  OAI22_X1 U5115 ( .A1(n9007), .A2(n4402), .B1(n7855), .B2(n8030), .ZN(n4716)
         );
  INV_X1 U5116 ( .A(n9091), .ZN(n7586) );
  NAND2_X1 U5117 ( .A1(n7330), .A2(n4420), .ZN(n7407) );
  NAND2_X1 U5118 ( .A1(n5069), .A2(n5634), .ZN(n5155) );
  NOR2_X1 U5119 ( .A1(n4993), .A2(n5634), .ZN(n4710) );
  INV_X1 U5120 ( .A(n5069), .ZN(n5507) );
  NAND2_X2 U5121 ( .A1(n5798), .A2(n6688), .ZN(n5069) );
  CLKBUF_X1 U5122 ( .A(n5777), .Z(n9140) );
  NOR2_X1 U5123 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(n4970), .ZN(n4973) );
  INV_X1 U5124 ( .A(n5007), .ZN(n4970) );
  INV_X1 U5125 ( .A(SI_3_), .ZN(n4542) );
  NAND3_X1 U5126 ( .A1(n9214), .A2(n4654), .A3(n4653), .ZN(n4652) );
  INV_X1 U5127 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4804) );
  OR2_X1 U5128 ( .A1(n8345), .A2(n8344), .ZN(n4625) );
  OAI21_X1 U5129 ( .B1(n8383), .B2(n9792), .A(n4637), .ZN(n4636) );
  AOI21_X1 U5130 ( .B1(n8385), .B2(n9790), .A(n8384), .ZN(n4637) );
  INV_X1 U5131 ( .A(n7489), .ZN(n9148) );
  NAND2_X1 U5132 ( .A1(n6309), .A2(n6293), .ZN(n4551) );
  INV_X1 U5133 ( .A(n9011), .ZN(n4567) );
  OAI22_X1 U5134 ( .A1(n4584), .A2(n9070), .B1(n4578), .B2(n4577), .ZN(n8993)
         );
  OR2_X1 U5135 ( .A1(n8990), .A2(n8994), .ZN(n4577) );
  AND2_X1 U5136 ( .A1(n4579), .A2(n8991), .ZN(n4578) );
  AND2_X1 U5137 ( .A1(n9021), .A2(n4574), .ZN(n4573) );
  NAND2_X1 U5138 ( .A1(n4403), .A2(n9020), .ZN(n4574) );
  NAND2_X1 U5139 ( .A1(n4403), .A2(n4576), .ZN(n4575) );
  INV_X1 U5140 ( .A(n9010), .ZN(n4576) );
  INV_X1 U5141 ( .A(n9036), .ZN(n4594) );
  NOR2_X1 U5142 ( .A1(n9041), .A2(n9040), .ZN(n4597) );
  OAI21_X1 U5143 ( .B1(n9039), .B2(n9038), .A(n9037), .ZN(n4598) );
  AOI21_X1 U5144 ( .B1(n9039), .B2(n9362), .A(n9033), .ZN(n4595) );
  INV_X1 U5145 ( .A(n5336), .ZN(n4906) );
  INV_X1 U5146 ( .A(n7899), .ZN(n4903) );
  INV_X1 U5147 ( .A(n5304), .ZN(n4519) );
  INV_X1 U5148 ( .A(n4690), .ZN(n4689) );
  INV_X1 U5149 ( .A(SI_13_), .ZN(n9970) );
  NAND2_X1 U5150 ( .A1(n5311), .A2(n5310), .ZN(n5337) );
  INV_X1 U5151 ( .A(n7537), .ZN(n4827) );
  NAND2_X1 U5152 ( .A1(n4755), .A2(n6386), .ZN(n4750) );
  INV_X1 U5153 ( .A(n4752), .ZN(n4748) );
  INV_X1 U5154 ( .A(n8565), .ZN(n4845) );
  INV_X1 U5155 ( .A(n8551), .ZN(n4739) );
  OR2_X1 U5156 ( .A1(n5992), .A2(n5991), .ZN(n6008) );
  NAND2_X1 U5157 ( .A1(n5967), .A2(n5966), .ZN(n5977) );
  AND2_X1 U5158 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n5966) );
  NAND2_X1 U5159 ( .A1(n6374), .A2(n4743), .ZN(n4742) );
  INV_X1 U5160 ( .A(n6375), .ZN(n4743) );
  NOR2_X1 U5161 ( .A1(n4535), .A2(n4745), .ZN(n4744) );
  INV_X1 U5162 ( .A(n6264), .ZN(n4745) );
  AND2_X1 U5163 ( .A1(n7258), .A2(n6369), .ZN(n6235) );
  NAND2_X1 U5164 ( .A1(n6924), .A2(n8325), .ZN(n6369) );
  INV_X1 U5165 ( .A(n6961), .ZN(n6367) );
  NAND2_X1 U5166 ( .A1(n8328), .A2(n9859), .ZN(n6251) );
  AND2_X1 U5167 ( .A1(n5845), .A2(n4932), .ZN(n5846) );
  OR2_X1 U5168 ( .A1(n7479), .A2(n4913), .ZN(n4912) );
  INV_X1 U5169 ( .A(n7145), .ZN(n4913) );
  NOR2_X1 U5170 ( .A1(n8799), .A2(n8800), .ZN(n4901) );
  NOR2_X1 U5171 ( .A1(n8791), .A2(n4897), .ZN(n4896) );
  INV_X1 U5172 ( .A(n8824), .ZN(n4897) );
  INV_X1 U5173 ( .A(n9136), .ZN(n4589) );
  NAND2_X1 U5174 ( .A1(n9063), .A2(n8994), .ZN(n9064) );
  AND2_X1 U5175 ( .A1(n8957), .A2(n9066), .ZN(n9138) );
  NAND2_X1 U5176 ( .A1(n9445), .A2(n9219), .ZN(n9066) );
  NAND2_X1 U5177 ( .A1(n4512), .A2(n4455), .ZN(n4510) );
  INV_X1 U5178 ( .A(n9668), .ZN(n4512) );
  NAND2_X1 U5179 ( .A1(n9656), .A2(n4513), .ZN(n4511) );
  NOR2_X1 U5180 ( .A1(n4514), .A2(n9668), .ZN(n4513) );
  INV_X1 U5181 ( .A(n9657), .ZN(n4514) );
  OR2_X1 U5182 ( .A1(n5739), .A2(n5738), .ZN(n5790) );
  AND2_X1 U5183 ( .A1(n9109), .A2(n9049), .ZN(n9228) );
  AND2_X1 U5184 ( .A1(n4615), .A2(n4614), .ZN(n4613) );
  OR2_X1 U5185 ( .A1(n9465), .A2(n8794), .ZN(n8131) );
  NOR2_X1 U5186 ( .A1(n9318), .A2(n4793), .ZN(n4792) );
  INV_X1 U5187 ( .A(n8897), .ZN(n4793) );
  NAND2_X1 U5188 ( .A1(n8130), .A2(n9042), .ZN(n9296) );
  NOR2_X1 U5189 ( .A1(n9478), .A2(n9481), .ZN(n4615) );
  OR2_X1 U5190 ( .A1(n9493), .A2(n8854), .ZN(n9034) );
  AND2_X1 U5191 ( .A1(n9013), .A2(n9014), .ZN(n9007) );
  OR2_X1 U5192 ( .A1(n7906), .A2(n9161), .ZN(n7799) );
  OR2_X1 U5193 ( .A1(n9573), .A2(n7889), .ZN(n4931) );
  INV_X1 U5194 ( .A(n8996), .ZN(n4466) );
  NAND2_X1 U5195 ( .A1(n5165), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5207) );
  INV_X1 U5196 ( .A(n5167), .ZN(n5165) );
  NOR2_X1 U5197 ( .A1(n9113), .A2(n4591), .ZN(n4590) );
  INV_X1 U5198 ( .A(n8913), .ZN(n4591) );
  NAND2_X1 U5199 ( .A1(n8914), .A2(n8913), .ZN(n4718) );
  INV_X1 U5200 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4946) );
  OAI21_X1 U5201 ( .B1(n5633), .B2(n4445), .A(n4701), .ZN(n5708) );
  INV_X1 U5202 ( .A(n4702), .ZN(n4701) );
  OAI21_X1 U5203 ( .B1(n4705), .B2(n4445), .A(n5679), .ZN(n4702) );
  NOR2_X1 U5204 ( .A1(n5604), .A2(n4685), .ZN(n4684) );
  INV_X1 U5205 ( .A(n5572), .ZN(n4685) );
  INV_X1 U5206 ( .A(n5569), .ZN(n4686) );
  OR2_X1 U5207 ( .A1(n4975), .A2(n4974), .ZN(n4976) );
  AOI21_X1 U5208 ( .B1(n4671), .B2(n4673), .A(n4669), .ZN(n4668) );
  INV_X1 U5209 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5450) );
  INV_X1 U5210 ( .A(n5384), .ZN(n4697) );
  INV_X1 U5211 ( .A(n4696), .ZN(n4695) );
  OAI21_X1 U5212 ( .B1(n4699), .B2(n4397), .A(n5418), .ZN(n4696) );
  AOI21_X1 U5213 ( .B1(n4388), .B2(n4667), .A(n4429), .ZN(n4665) );
  OR2_X1 U5214 ( .A1(n5282), .A2(n5281), .ZN(n5283) );
  AND2_X1 U5215 ( .A1(n5280), .A2(n5279), .ZN(n5281) );
  NOR2_X1 U5216 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n4941) );
  INV_X1 U5217 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4939) );
  AND2_X1 U5218 ( .A1(n5280), .A2(n5226), .ZN(n5277) );
  AOI21_X1 U5219 ( .B1(n5195), .B2(n4679), .A(n4427), .ZN(n4678) );
  NAND2_X1 U5220 ( .A1(n4380), .A2(n5067), .ZN(n4543) );
  NOR2_X2 U5221 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5044) );
  NAND2_X1 U5222 ( .A1(n4813), .A2(n4479), .ZN(n4478) );
  INV_X1 U5223 ( .A(n8155), .ZN(n4479) );
  NAND2_X1 U5224 ( .A1(n4806), .A2(n4411), .ZN(n8011) );
  INV_X1 U5225 ( .A(n7877), .ZN(n4805) );
  NAND2_X1 U5226 ( .A1(n4490), .A2(n7731), .ZN(n4806) );
  AND2_X1 U5227 ( .A1(n4809), .A2(n7730), .ZN(n4490) );
  NOR2_X1 U5228 ( .A1(n8144), .A2(n8143), .ZN(n8225) );
  AOI21_X1 U5229 ( .B1(n4815), .B2(n4814), .A(n8151), .ZN(n4813) );
  INV_X1 U5230 ( .A(n4444), .ZN(n4814) );
  OAI21_X1 U5231 ( .B1(n8013), .B2(n4487), .A(n4485), .ZN(n8081) );
  AND2_X1 U5232 ( .A1(n8012), .A2(n8014), .ZN(n4487) );
  AND2_X1 U5233 ( .A1(n8039), .A2(n4486), .ZN(n4485) );
  OR2_X1 U5234 ( .A1(n8012), .A2(n8014), .ZN(n4486) );
  OR2_X1 U5235 ( .A1(n6112), .A2(n6111), .ZN(n6124) );
  NOR2_X1 U5236 ( .A1(n7502), .A2(n4827), .ZN(n4825) );
  INV_X1 U5237 ( .A(n7621), .ZN(n4826) );
  OR2_X1 U5238 ( .A1(n7123), .A2(n7124), .ZN(n4821) );
  INV_X1 U5239 ( .A(n8251), .ZN(n4818) );
  OR2_X1 U5240 ( .A1(n6865), .A2(n9819), .ZN(n6874) );
  AND2_X1 U5241 ( .A1(n6142), .A2(n6141), .ZN(n8254) );
  OR2_X1 U5242 ( .A1(n6414), .A2(n7836), .ZN(n6869) );
  AND4_X1 U5243 ( .A1(n6029), .A2(n6028), .A3(n6027), .A4(n6026), .ZN(n7991)
         );
  OR2_X1 U5244 ( .A1(n6627), .A2(n6626), .ZN(n4620) );
  NOR2_X1 U5245 ( .A1(n6784), .A2(n4457), .ZN(n6786) );
  AOI21_X1 U5246 ( .B1(n4755), .B2(n8429), .A(n4753), .ZN(n4752) );
  INV_X1 U5247 ( .A(n6336), .ZN(n4753) );
  OR2_X1 U5248 ( .A1(n4936), .A2(n4754), .ZN(n4751) );
  OR2_X1 U5249 ( .A1(n8646), .A2(n8434), .ZN(n8201) );
  NAND2_X1 U5250 ( .A1(n4647), .A2(n4646), .ZN(n8416) );
  NAND2_X1 U5251 ( .A1(n4876), .A2(n4875), .ZN(n8458) );
  AOI21_X1 U5252 ( .B1(n4877), .B2(n4879), .A(n6143), .ZN(n4875) );
  OR2_X1 U5253 ( .A1(n8461), .A2(n8460), .ZN(n8463) );
  AND2_X1 U5254 ( .A1(n8488), .A2(n4881), .ZN(n4880) );
  AND2_X1 U5255 ( .A1(n6315), .A2(n8504), .ZN(n8523) );
  NAND2_X1 U5256 ( .A1(n8192), .A2(n4391), .ZN(n4842) );
  NAND2_X1 U5257 ( .A1(n8192), .A2(n4443), .ZN(n4840) );
  AND3_X1 U5258 ( .A1(n6096), .A2(n6095), .A3(n6094), .ZN(n8555) );
  OR2_X1 U5259 ( .A1(n8696), .A2(n8554), .ZN(n6301) );
  NAND2_X1 U5260 ( .A1(n6076), .A2(n4401), .ZN(n8549) );
  INV_X1 U5261 ( .A(n6067), .ZN(n4769) );
  INV_X1 U5262 ( .A(n6298), .ZN(n4770) );
  AND2_X1 U5263 ( .A1(n6301), .A2(n6309), .ZN(n8564) );
  NAND2_X1 U5264 ( .A1(n8614), .A2(n6067), .ZN(n8586) );
  AND2_X1 U5265 ( .A1(n8610), .A2(n8185), .ZN(n4862) );
  INV_X1 U5266 ( .A(n7929), .ZN(n4860) );
  NAND2_X1 U5267 ( .A1(n6000), .A2(n4765), .ZN(n7963) );
  AND4_X1 U5268 ( .A1(n6013), .A2(n6012), .A3(n6011), .A4(n6010), .ZN(n7965)
         );
  INV_X1 U5269 ( .A(n7710), .ZN(n7633) );
  NOR2_X1 U5270 ( .A1(n5931), .A2(n5930), .ZN(n5941) );
  OR2_X1 U5271 ( .A1(n7384), .A2(n8323), .ZN(n4870) );
  NOR2_X1 U5272 ( .A1(n7385), .A2(n4869), .ZN(n4868) );
  INV_X1 U5273 ( .A(n7178), .ZN(n4869) );
  NAND2_X1 U5274 ( .A1(n4867), .A2(n4865), .ZN(n7632) );
  NOR2_X1 U5275 ( .A1(n7391), .A2(n4866), .ZN(n4865) );
  INV_X1 U5276 ( .A(n4870), .ZN(n4866) );
  AND2_X1 U5277 ( .A1(n6261), .A2(n6260), .ZN(n7385) );
  NAND2_X1 U5278 ( .A1(n7256), .A2(n9876), .ZN(n7185) );
  OR2_X1 U5279 ( .A1(n6827), .A2(n6826), .ZN(n8617) );
  INV_X1 U5280 ( .A(n8591), .ZN(n8615) );
  NAND2_X1 U5281 ( .A1(n6834), .A2(n4386), .ZN(n4861) );
  AND2_X1 U5282 ( .A1(n6895), .A2(n9847), .ZN(n6892) );
  NAND2_X1 U5283 ( .A1(n6190), .A2(n6189), .ZN(n8636) );
  NAND2_X1 U5284 ( .A1(n6046), .A2(n6045), .ZN(n8706) );
  AND2_X1 U5285 ( .A1(n6807), .A2(n6806), .ZN(n9820) );
  INV_X1 U5286 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5827) );
  NAND2_X1 U5287 ( .A1(n6400), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6410) );
  NAND2_X1 U5288 ( .A1(n5847), .A2(n4836), .ZN(n4835) );
  NAND2_X1 U5289 ( .A1(n5844), .A2(n5846), .ZN(n6068) );
  AND2_X1 U5290 ( .A1(n5913), .A2(n5926), .ZN(n6578) );
  NAND2_X1 U5291 ( .A1(n7100), .A2(n4915), .ZN(n4914) );
  INV_X1 U5292 ( .A(n4916), .ZN(n4915) );
  NAND2_X1 U5293 ( .A1(n4909), .A2(n4907), .ZN(n8830) );
  AOI21_X1 U5294 ( .B1(n8775), .B2(n5524), .A(n4908), .ZN(n4907) );
  INV_X1 U5295 ( .A(n8832), .ZN(n4908) );
  OR2_X1 U5296 ( .A1(n5579), .A2(n8852), .ZN(n5619) );
  OAI21_X1 U5297 ( .B1(n8791), .B2(n4895), .A(n5678), .ZN(n4894) );
  INV_X1 U5298 ( .A(n4929), .ZN(n4895) );
  NAND2_X1 U5299 ( .A1(n8823), .A2(n4896), .ZN(n4893) );
  NAND2_X1 U5300 ( .A1(n9656), .A2(n9657), .ZN(n9654) );
  OAI21_X1 U5301 ( .B1(n9701), .B2(n4504), .A(n4503), .ZN(n9710) );
  NAND2_X1 U5302 ( .A1(n4507), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4504) );
  NAND2_X1 U5303 ( .A1(n9196), .A2(n4507), .ZN(n4503) );
  INV_X1 U5304 ( .A(n9711), .ZN(n4507) );
  OR2_X1 U5305 ( .A1(n9701), .A2(n9700), .ZN(n4506) );
  NAND2_X1 U5306 ( .A1(n8885), .A2(n8884), .ZN(n9450) );
  NOR2_X1 U5307 ( .A1(n9056), .A2(n9060), .ZN(n9237) );
  AND2_X1 U5308 ( .A1(n9074), .A2(n9236), .ZN(n9264) );
  NAND2_X1 U5309 ( .A1(n9157), .A2(n9438), .ZN(n4468) );
  NAND2_X1 U5310 ( .A1(n4614), .A2(n9315), .ZN(n8122) );
  NAND2_X1 U5311 ( .A1(n8131), .A2(n9048), .ZN(n9284) );
  NAND2_X1 U5312 ( .A1(n5637), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5665) );
  INV_X1 U5313 ( .A(n5639), .ZN(n5637) );
  NAND2_X1 U5314 ( .A1(n9334), .A2(n4792), .ZN(n4795) );
  OAI21_X1 U5315 ( .B1(n8119), .B2(n9101), .A(n4707), .ZN(n9294) );
  AOI21_X1 U5316 ( .B1(n9318), .B2(n4708), .A(n4422), .ZN(n4707) );
  INV_X1 U5317 ( .A(n8962), .ZN(n4708) );
  OR2_X1 U5318 ( .A1(n9481), .A2(n9314), .ZN(n8897) );
  INV_X1 U5319 ( .A(n9354), .ZN(n9314) );
  OAI21_X1 U5320 ( .B1(n8854), .B2(n9377), .A(n9360), .ZN(n9344) );
  OR2_X1 U5321 ( .A1(n9496), .A2(n9368), .ZN(n9362) );
  INV_X1 U5322 ( .A(n4801), .ZN(n4800) );
  NAND2_X1 U5323 ( .A1(n4803), .A2(n9418), .ZN(n4802) );
  NAND2_X1 U5324 ( .A1(n9431), .A2(n4729), .ZN(n4728) );
  INV_X1 U5325 ( .A(n8115), .ZN(n4729) );
  NAND2_X1 U5326 ( .A1(n9509), .A2(n9410), .ZN(n4730) );
  OR2_X1 U5327 ( .A1(n9514), .A2(n9436), .ZN(n8113) );
  OR2_X1 U5328 ( .A1(n8816), .A2(n8803), .ZN(n4927) );
  OR2_X1 U5329 ( .A1(n9417), .A2(n9418), .ZN(n4731) );
  NAND2_X1 U5330 ( .A1(n4782), .A2(n9013), .ZN(n4781) );
  NAND2_X1 U5331 ( .A1(n4777), .A2(n9014), .ZN(n4782) );
  NAND2_X1 U5332 ( .A1(n9094), .A2(n9004), .ZN(n4777) );
  INV_X1 U5333 ( .A(n9007), .ZN(n9095) );
  INV_X1 U5334 ( .A(n9159), .ZN(n8030) );
  NAND2_X1 U5335 ( .A1(n7800), .A2(n7799), .ZN(n7850) );
  INV_X1 U5336 ( .A(n9160), .ZN(n8904) );
  AND2_X1 U5337 ( .A1(n8921), .A2(n8905), .ZN(n9091) );
  AOI21_X1 U5338 ( .B1(n7448), .B2(n7334), .A(n7333), .ZN(n7335) );
  NAND2_X1 U5339 ( .A1(n7335), .A2(n9087), .ZN(n7585) );
  AND2_X1 U5340 ( .A1(n8924), .A2(n8983), .ZN(n9085) );
  NAND2_X1 U5341 ( .A1(n7217), .A2(n7216), .ZN(n7330) );
  OR2_X1 U5342 ( .A1(n6997), .A2(n6996), .ZN(n9371) );
  INV_X1 U5343 ( .A(n6982), .ZN(n6984) );
  INV_X1 U5344 ( .A(n9369), .ZN(n9437) );
  INV_X1 U5345 ( .A(n9389), .ZN(n9433) );
  INV_X1 U5346 ( .A(n9371), .ZN(n9438) );
  NAND2_X1 U5347 ( .A1(n5578), .A2(n5577), .ZN(n9486) );
  OR2_X1 U5348 ( .A1(n7072), .A2(n5787), .ZN(n9774) );
  NAND2_X1 U5349 ( .A1(n6718), .A2(n7348), .ZN(n6987) );
  INV_X1 U5350 ( .A(n9774), .ZN(n9564) );
  XNOR2_X1 U5351 ( .A(n5681), .B(n5680), .ZN(n7943) );
  NAND2_X1 U5352 ( .A1(n4704), .A2(n5657), .ZN(n5681) );
  NAND2_X1 U5353 ( .A1(n4698), .A2(n5384), .ZN(n5420) );
  NAND4_X1 U5354 ( .A1(n4944), .A2(n10225), .A3(n5260), .A4(n5229), .ZN(n4945)
         );
  INV_X1 U5355 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n4944) );
  OR2_X1 U5356 ( .A1(n5285), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5314) );
  INV_X1 U5357 ( .A(n8486), .ZN(n8669) );
  AND4_X1 U5358 ( .A1(n6041), .A2(n6040), .A3(n6039), .A4(n6038), .ZN(n8616)
         );
  NAND2_X1 U5359 ( .A1(n6133), .A2(n6132), .ZN(n8662) );
  NAND2_X1 U5360 ( .A1(n6110), .A2(n6109), .ZN(n8674) );
  NOR4_X1 U5361 ( .A1(n6389), .A2(n6388), .A3(n8210), .A4(n6387), .ZN(n6390)
         );
  NAND2_X1 U5362 ( .A1(n4389), .A2(n4460), .ZN(n4538) );
  AOI21_X1 U5363 ( .B1(n6218), .B2(n6355), .A(n6356), .ZN(n6219) );
  NAND2_X1 U5364 ( .A1(n6395), .A2(n4462), .ZN(n4540) );
  OR2_X1 U5365 ( .A1(n6395), .A2(n6396), .ZN(n4541) );
  INV_X1 U5366 ( .A(n8229), .ZN(n8525) );
  NAND2_X1 U5367 ( .A1(n6662), .A2(n4632), .ZN(n4631) );
  NAND2_X1 U5368 ( .A1(n6655), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4632) );
  AND2_X1 U5369 ( .A1(n4631), .A2(n4630), .ZN(n6610) );
  INV_X1 U5370 ( .A(n6611), .ZN(n4630) );
  OR2_X1 U5371 ( .A1(n6575), .A2(n6574), .ZN(n4622) );
  AND2_X1 U5372 ( .A1(n4622), .A2(n4621), .ZN(n6627) );
  NAND2_X1 U5373 ( .A1(n6623), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4621) );
  NOR2_X1 U5374 ( .A1(n8341), .A2(n4626), .ZN(n8345) );
  NOR2_X1 U5375 ( .A1(n4628), .A2(n4627), .ZN(n4626) );
  INV_X1 U5376 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n4627) );
  INV_X1 U5377 ( .A(n4623), .ZN(n8374) );
  AND2_X1 U5378 ( .A1(n8216), .A2(n8215), .ZN(n8639) );
  NAND2_X1 U5379 ( .A1(n8211), .A2(n8585), .ZN(n8216) );
  NAND2_X1 U5380 ( .A1(n8204), .A2(n8405), .ZN(n4853) );
  OAI21_X1 U5381 ( .B1(n4413), .B2(n8204), .A(n4852), .ZN(n4851) );
  NAND2_X1 U5382 ( .A1(n8432), .A2(n6332), .ZN(n8420) );
  INV_X1 U5383 ( .A(n6227), .ZN(n9812) );
  AND2_X1 U5384 ( .A1(n8629), .A2(n6832), .ZN(n8606) );
  INV_X1 U5385 ( .A(n9157), .ZN(n9242) );
  NAND2_X1 U5386 ( .A1(n5369), .A2(n5368), .ZN(n9524) );
  NAND2_X1 U5387 ( .A1(n5735), .A2(n5734), .ZN(n9455) );
  INV_X1 U5388 ( .A(n9167), .ZN(n7694) );
  NAND2_X1 U5389 ( .A1(n4601), .A2(n4600), .ZN(n4599) );
  NAND2_X1 U5390 ( .A1(n8065), .A2(n8064), .ZN(n8798) );
  INV_X1 U5391 ( .A(n9282), .ZN(n9229) );
  AOI21_X1 U5392 ( .B1(n4585), .B2(n4934), .A(n9147), .ZN(n9149) );
  XNOR2_X1 U5393 ( .A(n4586), .B(n9071), .ZN(n4585) );
  NAND2_X1 U5394 ( .A1(n5697), .A2(n5696), .ZN(n9299) );
  NAND2_X1 U5395 ( .A1(n5098), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n4966) );
  NOR2_X1 U5396 ( .A1(n9210), .A2(n9751), .ZN(n4501) );
  NOR2_X1 U5397 ( .A1(n9211), .A2(n9741), .ZN(n4497) );
  NAND2_X1 U5398 ( .A1(n9212), .A2(n7289), .ZN(n4502) );
  NAND2_X1 U5399 ( .A1(n8878), .A2(n8877), .ZN(n9563) );
  OR2_X1 U5400 ( .A1(n9776), .A2(n6981), .ZN(n9425) );
  OAI211_X1 U5401 ( .C1(n5155), .C2(n8049), .A(n5075), .B(n5074), .ZN(n7380)
         );
  NOR2_X1 U5402 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n4954) );
  INV_X1 U5403 ( .A(n6266), .ZN(n4534) );
  NAND2_X1 U5404 ( .A1(n4532), .A2(n4536), .ZN(n4531) );
  NAND2_X1 U5405 ( .A1(n4537), .A2(n4533), .ZN(n4532) );
  INV_X1 U5406 ( .A(n6272), .ZN(n4537) );
  NAND2_X1 U5407 ( .A1(n6273), .A2(n4423), .ZN(n4533) );
  NAND2_X1 U5408 ( .A1(n4583), .A2(n4582), .ZN(n8986) );
  NAND2_X1 U5409 ( .A1(n8977), .A2(n8994), .ZN(n4583) );
  NAND2_X1 U5410 ( .A1(n8978), .A2(n9070), .ZN(n4582) );
  OAI21_X1 U5411 ( .B1(n8986), .B2(n8985), .A(n4580), .ZN(n4579) );
  NOR2_X1 U5412 ( .A1(n7591), .A2(n4581), .ZN(n4580) );
  INV_X1 U5413 ( .A(n8983), .ZN(n4581) );
  AOI21_X1 U5414 ( .B1(n4546), .B2(n6360), .A(n6299), .ZN(n4545) );
  AOI21_X1 U5415 ( .B1(n6292), .B2(n8587), .A(n4551), .ZN(n4550) );
  NAND2_X1 U5416 ( .A1(n4569), .A2(n4565), .ZN(n9028) );
  AND2_X1 U5417 ( .A1(n4573), .A2(n4566), .ZN(n4565) );
  NAND2_X1 U5418 ( .A1(n4568), .A2(n4567), .ZN(n4566) );
  NAND2_X1 U5419 ( .A1(n4571), .A2(n4570), .ZN(n9026) );
  AOI21_X1 U5420 ( .B1(n4573), .B2(n4575), .A(n4430), .ZN(n4570) );
  NAND2_X1 U5421 ( .A1(n4553), .A2(n6153), .ZN(n4552) );
  NAND2_X1 U5422 ( .A1(n4556), .A2(n6325), .ZN(n4555) );
  NAND2_X1 U5423 ( .A1(n4596), .A2(n4592), .ZN(n9046) );
  OAI21_X1 U5424 ( .B1(n4595), .B2(n9038), .A(n4593), .ZN(n4592) );
  NOR2_X1 U5425 ( .A1(n4594), .A2(n9070), .ZN(n4593) );
  NAND2_X1 U5426 ( .A1(n7032), .A2(n6364), .ZN(n6243) );
  INV_X1 U5427 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4952) );
  INV_X1 U5428 ( .A(n5731), .ZN(n4691) );
  INV_X1 U5429 ( .A(n5657), .ZN(n4703) );
  INV_X1 U5430 ( .A(n5551), .ZN(n4669) );
  INV_X1 U5431 ( .A(n5441), .ZN(n4694) );
  INV_X1 U5432 ( .A(n5338), .ZN(n4663) );
  INV_X1 U5433 ( .A(n5178), .ZN(n4679) );
  AND2_X1 U5434 ( .A1(n6834), .A2(n8148), .ZN(n6856) );
  XNOR2_X1 U5435 ( .A(n8163), .B(n4386), .ZN(n6855) );
  INV_X1 U5436 ( .A(n6362), .ZN(n4656) );
  OR2_X1 U5437 ( .A1(n8636), .A2(n8168), .ZN(n6349) );
  AOI21_X1 U5438 ( .B1(n8405), .B2(n4855), .A(n4407), .ZN(n4854) );
  INV_X1 U5439 ( .A(n8201), .ZN(n4855) );
  NAND2_X1 U5440 ( .A1(n8460), .A2(n6228), .ZN(n4775) );
  INV_X1 U5441 ( .A(n4842), .ZN(n4841) );
  NAND2_X1 U5442 ( .A1(n4840), .A2(n4842), .ZN(n4839) );
  NOR2_X1 U5443 ( .A1(n8693), .A2(n8696), .ZN(n4649) );
  NAND2_X1 U5444 ( .A1(n6085), .A2(n6084), .ZN(n6092) );
  INV_X1 U5445 ( .A(n6083), .ZN(n6085) );
  INV_X1 U5446 ( .A(n8587), .ZN(n8187) );
  NAND2_X1 U5447 ( .A1(n7961), .A2(n4645), .ZN(n4644) );
  NOR2_X1 U5448 ( .A1(n8722), .A2(n7931), .ZN(n4645) );
  INV_X1 U5449 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5991) );
  INV_X1 U5450 ( .A(n7676), .ZN(n4873) );
  OAI21_X1 U5451 ( .B1(n4400), .B2(n4873), .A(n7745), .ZN(n4872) );
  OR2_X1 U5452 ( .A1(n5977), .A2(n7625), .ZN(n5992) );
  NAND2_X1 U5453 ( .A1(n6227), .A2(n7010), .ZN(n6873) );
  NAND2_X1 U5454 ( .A1(n6243), .A2(n6365), .ZN(n6881) );
  INV_X1 U5455 ( .A(n4835), .ZN(n4833) );
  NAND2_X1 U5456 ( .A1(n5138), .A2(n4461), .ZN(n4916) );
  INV_X1 U5457 ( .A(n7101), .ZN(n4526) );
  NAND2_X1 U5458 ( .A1(n4911), .A2(n4916), .ZN(n4910) );
  XNOR2_X1 U5459 ( .A(n5132), .B(n5049), .ZN(n5133) );
  AND2_X1 U5460 ( .A1(n4902), .A2(n4518), .ZN(n4517) );
  NAND2_X1 U5461 ( .A1(n4904), .A2(n4519), .ZN(n4518) );
  AOI21_X1 U5462 ( .B1(n4904), .B2(n7887), .A(n4903), .ZN(n4902) );
  OR3_X1 U5463 ( .A1(n8947), .A2(n9044), .A3(n9050), .ZN(n9134) );
  AND2_X1 U5464 ( .A1(n4511), .A2(n4509), .ZN(n9192) );
  AND2_X1 U5465 ( .A1(n4510), .A2(n4459), .ZN(n4509) );
  NOR2_X1 U5466 ( .A1(n8116), .A2(n4727), .ZN(n4724) );
  NAND2_X1 U5467 ( .A1(n8816), .A2(n4611), .ZN(n4610) );
  NOR2_X1 U5468 ( .A1(n9509), .A2(n4610), .ZN(n4609) );
  NOR2_X1 U5469 ( .A1(n9007), .A2(n4425), .ZN(n4712) );
  INV_X1 U5470 ( .A(n7799), .ZN(n4713) );
  INV_X1 U5471 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5395) );
  NAND2_X1 U5472 ( .A1(n4393), .A2(n7608), .ZN(n4606) );
  AND2_X1 U5473 ( .A1(n7593), .A2(n8988), .ZN(n8981) );
  OR2_X1 U5474 ( .A1(n7664), .A2(n7594), .ZN(n7592) );
  NAND2_X1 U5475 ( .A1(n5139), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5167) );
  NAND2_X1 U5476 ( .A1(n7311), .A2(n4379), .ZN(n7308) );
  NAND2_X1 U5477 ( .A1(n4562), .A2(n4561), .ZN(n4994) );
  NAND2_X1 U5478 ( .A1(n4953), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4561) );
  NAND2_X1 U5479 ( .A1(n4564), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4563) );
  AND2_X1 U5480 ( .A1(n5731), .A2(n5714), .ZN(n5715) );
  AND2_X1 U5481 ( .A1(n5709), .A2(n5685), .ZN(n5707) );
  AND2_X1 U5482 ( .A1(n10082), .A2(n4985), .ZN(n4917) );
  INV_X1 U5483 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4980) );
  NOR2_X1 U5484 ( .A1(n5653), .A2(n4706), .ZN(n4705) );
  INV_X1 U5485 ( .A(n5632), .ZN(n4706) );
  INV_X1 U5486 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n10082) );
  NAND2_X1 U5487 ( .A1(n4975), .A2(n4974), .ZN(n5003) );
  NOR2_X1 U5488 ( .A1(n5526), .A2(n4675), .ZN(n4674) );
  INV_X1 U5489 ( .A(n5502), .ZN(n4675) );
  AND2_X1 U5490 ( .A1(n5446), .A2(n4969), .ZN(n5007) );
  INV_X1 U5491 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5447) );
  NOR2_X1 U5492 ( .A1(n5385), .A2(n4700), .ZN(n4699) );
  INV_X1 U5493 ( .A(n5363), .ZN(n4700) );
  INV_X1 U5494 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4654) );
  AOI21_X1 U5495 ( .B1(n4809), .B2(n4808), .A(n4424), .ZN(n4807) );
  INV_X1 U5496 ( .A(n7762), .ZN(n4808) );
  OR2_X1 U5497 ( .A1(n6092), .A2(n8106), .ZN(n6100) );
  OR2_X1 U5498 ( .A1(n6036), .A2(n10068), .ZN(n6049) );
  NOR2_X1 U5499 ( .A1(n4529), .A2(n4415), .ZN(n4528) );
  NOR2_X1 U5500 ( .A1(n6557), .A2(n6619), .ZN(n4529) );
  OAI22_X1 U5501 ( .A1(n7465), .A2(n7464), .B1(n7463), .B2(n7462), .ZN(n7491)
         );
  NAND2_X1 U5502 ( .A1(n4828), .A2(n7502), .ZN(n7538) );
  INV_X1 U5503 ( .A(n7505), .ZN(n4828) );
  AND2_X1 U5504 ( .A1(n4928), .A2(n8080), .ZN(n4831) );
  INV_X1 U5505 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6089) );
  NAND2_X1 U5506 ( .A1(n6099), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6112) );
  INV_X1 U5507 ( .A(n6100), .ZN(n6099) );
  NAND2_X1 U5508 ( .A1(n6857), .A2(n6948), .ZN(n4820) );
  NAND2_X1 U5509 ( .A1(n8328), .A2(n8148), .ZN(n6904) );
  NAND2_X1 U5510 ( .A1(n4817), .A2(n4444), .ZN(n4816) );
  INV_X1 U5511 ( .A(n8250), .ZN(n4817) );
  OR2_X1 U5512 ( .A1(n8013), .A2(n8012), .ZN(n4829) );
  NAND2_X1 U5513 ( .A1(n6403), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6399) );
  NAND2_X1 U5514 ( .A1(n6358), .A2(n6357), .ZN(n6388) );
  INV_X1 U5515 ( .A(n6355), .ZN(n6389) );
  AOI21_X1 U5516 ( .B1(n6359), .B2(n8390), .A(n6351), .ZN(n6355) );
  NAND2_X1 U5517 ( .A1(n6393), .A2(n9812), .ZN(n6825) );
  AND2_X1 U5518 ( .A1(n6118), .A2(n6117), .ZN(n8229) );
  AND4_X1 U5519 ( .A1(n6054), .A2(n6053), .A3(n6052), .A4(n6051), .ZN(n8262)
         );
  AND4_X1 U5520 ( .A1(n5997), .A2(n5996), .A3(n5995), .A4(n5994), .ZN(n7764)
         );
  NOR2_X1 U5521 ( .A1(n6786), .A2(n6787), .ZN(n4639) );
  NAND2_X1 U5522 ( .A1(n7426), .A2(n4618), .ZN(n7428) );
  OR2_X1 U5523 ( .A1(n7427), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4618) );
  NAND2_X1 U5524 ( .A1(n7428), .A2(n7429), .ZN(n7527) );
  NAND2_X1 U5525 ( .A1(n7527), .A2(n4617), .ZN(n7529) );
  OR2_X1 U5526 ( .A1(n7528), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4617) );
  NAND2_X1 U5527 ( .A1(n7529), .A2(n7530), .ZN(n7917) );
  NAND2_X1 U5528 ( .A1(n4625), .A2(n4624), .ZN(n4623) );
  NAND2_X1 U5529 ( .A1(n8366), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4624) );
  AOI21_X1 U5530 ( .B1(n6386), .B2(n4748), .A(n4747), .ZN(n4746) );
  INV_X1 U5531 ( .A(n6337), .ZN(n4747) );
  NAND2_X1 U5532 ( .A1(n6349), .A2(n6350), .ZN(n8210) );
  NOR2_X1 U5533 ( .A1(n8204), .A2(n4850), .ZN(n4849) );
  INV_X1 U5534 ( .A(n4854), .ZN(n4850) );
  NAND2_X1 U5535 ( .A1(n8204), .A2(n4854), .ZN(n4852) );
  OR2_X1 U5536 ( .A1(n6147), .A2(n6146), .ZN(n6158) );
  INV_X1 U5537 ( .A(n4736), .ZN(n4732) );
  INV_X1 U5538 ( .A(n8523), .ZN(n4735) );
  NAND2_X1 U5539 ( .A1(n8596), .A2(n4649), .ZN(n8556) );
  AND2_X1 U5540 ( .A1(n8596), .A2(n4392), .ZN(n8542) );
  NAND2_X1 U5541 ( .A1(n4844), .A2(n4846), .ZN(n8548) );
  NAND2_X1 U5542 ( .A1(n4845), .A2(n4443), .ZN(n4844) );
  AND2_X1 U5543 ( .A1(n8622), .A2(n8603), .ZN(n8596) );
  NAND2_X1 U5544 ( .A1(n8596), .A2(n8571), .ZN(n8566) );
  NAND2_X1 U5545 ( .A1(n8582), .A2(n8189), .ZN(n8565) );
  NAND2_X1 U5546 ( .A1(n6047), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6060) );
  INV_X1 U5547 ( .A(n6049), .ZN(n6047) );
  NOR2_X2 U5548 ( .A1(n8623), .A2(n8706), .ZN(n8622) );
  NAND2_X1 U5549 ( .A1(n6042), .A2(n6290), .ZN(n8611) );
  NAND2_X1 U5550 ( .A1(n8186), .A2(n8185), .ZN(n8608) );
  NAND2_X1 U5551 ( .A1(n6042), .A2(n4771), .ZN(n8614) );
  INV_X1 U5552 ( .A(n6287), .ZN(n4764) );
  AOI21_X1 U5553 ( .B1(n4858), .B2(n7930), .A(n4451), .ZN(n4857) );
  NOR2_X1 U5554 ( .A1(n7685), .A2(n4643), .ZN(n7957) );
  INV_X1 U5555 ( .A(n4645), .ZN(n4643) );
  AOI21_X1 U5556 ( .B1(n7389), .B2(n4410), .A(n4741), .ZN(n4937) );
  OAI21_X1 U5557 ( .B1(n4742), .B2(n6269), .A(n6373), .ZN(n4741) );
  INV_X1 U5558 ( .A(n7745), .ZN(n5983) );
  NAND2_X1 U5559 ( .A1(n4740), .A2(n4742), .ZN(n7637) );
  NAND2_X1 U5560 ( .A1(n7389), .A2(n4744), .ZN(n4740) );
  AND4_X1 U5561 ( .A1(n5982), .A2(n5981), .A3(n5980), .A4(n5979), .ZN(n7739)
         );
  AND2_X1 U5562 ( .A1(n6375), .A2(n6374), .ZN(n7710) );
  NAND2_X1 U5563 ( .A1(n7389), .A2(n6264), .ZN(n7704) );
  AND4_X1 U5564 ( .A1(n5946), .A2(n5945), .A3(n5944), .A4(n5943), .ZN(n7706)
         );
  AND4_X1 U5565 ( .A1(n5972), .A2(n5971), .A3(n5970), .A4(n5969), .ZN(n7705)
         );
  INV_X1 U5566 ( .A(n5901), .ZN(n6217) );
  INV_X1 U5567 ( .A(n6557), .ZN(n6077) );
  INV_X1 U5568 ( .A(n6370), .ZN(n4759) );
  AND4_X1 U5569 ( .A1(n5898), .A2(n5897), .A3(n5896), .A4(n5895), .ZN(n7262)
         );
  AND4_X1 U5570 ( .A1(n5920), .A2(n5919), .A3(n5918), .A4(n5917), .ZN(n7263)
         );
  INV_X1 U5571 ( .A(n6967), .ZN(n4640) );
  OAI21_X1 U5572 ( .B1(n6881), .B2(n6882), .A(n6250), .ZN(n6960) );
  AND2_X1 U5573 ( .A1(n6862), .A2(n6826), .ZN(n8591) );
  CLKBUF_X1 U5574 ( .A(n6833), .Z(n6893) );
  OR2_X1 U5575 ( .A1(n6821), .A2(n7006), .ZN(n6841) );
  NAND2_X1 U5576 ( .A1(n4489), .A2(n4488), .ZN(n8148) );
  INV_X1 U5577 ( .A(n6873), .ZN(n4488) );
  NAND2_X1 U5578 ( .A1(n4651), .A2(n6202), .ZN(n9557) );
  NAND2_X1 U5579 ( .A1(n8876), .A2(n5947), .ZN(n4651) );
  INV_X1 U5580 ( .A(n7026), .ZN(n7009) );
  OR3_X1 U5581 ( .A1(n7008), .A2(n7007), .A3(n7006), .ZN(n7027) );
  NAND2_X1 U5582 ( .A1(n4834), .A2(n4832), .ZN(n6403) );
  AND2_X1 U5583 ( .A1(n4833), .A2(n6221), .ZN(n4832) );
  INV_X1 U5584 ( .A(n6068), .ZN(n4834) );
  INV_X1 U5585 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6221) );
  NAND2_X1 U5586 ( .A1(n4491), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6223) );
  AND2_X1 U5587 ( .A1(n6032), .A2(n6019), .ZN(n7918) );
  AND2_X1 U5588 ( .A1(n5961), .A2(n5973), .ZN(n7115) );
  AND2_X1 U5589 ( .A1(n5951), .A2(n5987), .ZN(n6785) );
  INV_X1 U5590 ( .A(n4896), .ZN(n4890) );
  INV_X1 U5591 ( .A(n4892), .ZN(n4888) );
  NAND2_X1 U5592 ( .A1(n5028), .A2(n7346), .ZN(n5629) );
  INV_X1 U5593 ( .A(n6467), .ZN(n4600) );
  NAND2_X1 U5594 ( .A1(n4521), .A2(n4406), .ZN(n4520) );
  INV_X1 U5595 ( .A(n4901), .ZN(n4521) );
  NAND2_X1 U5596 ( .A1(n8067), .A2(n4899), .ZN(n4523) );
  NOR2_X1 U5597 ( .A1(n4901), .A2(n4900), .ZN(n4899) );
  INV_X1 U5598 ( .A(n8068), .ZN(n4900) );
  NAND2_X1 U5599 ( .A1(n5417), .A2(n4898), .ZN(n4522) );
  NOR2_X1 U5600 ( .A1(n4901), .A2(n5415), .ZN(n4898) );
  NAND2_X1 U5601 ( .A1(n5617), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5639) );
  INV_X1 U5602 ( .A(n5619), .ZN(n5617) );
  XNOR2_X1 U5603 ( .A(n5107), .B(n5750), .ZN(n5108) );
  XNOR2_X1 U5604 ( .A(n5246), .B(n5247), .ZN(n7780) );
  NAND2_X1 U5605 ( .A1(n5535), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5557) );
  INV_X1 U5606 ( .A(n5537), .ZN(n5535) );
  OR2_X1 U5607 ( .A1(n5511), .A2(n5510), .ZN(n5537) );
  OR2_X1 U5608 ( .A1(n5557), .A2(n8785), .ZN(n5579) );
  INV_X1 U5609 ( .A(n9388), .ZN(n8854) );
  INV_X1 U5610 ( .A(n5494), .ZN(n5495) );
  NOR2_X1 U5611 ( .A1(n4894), .A2(n6421), .ZN(n4892) );
  INV_X1 U5612 ( .A(n4588), .ZN(n4587) );
  OAI22_X1 U5613 ( .A1(n9068), .A2(n4589), .B1(n9138), .B2(n9070), .ZN(n4588)
         );
  OAI21_X1 U5614 ( .B1(n9108), .B2(n9107), .A(n9106), .ZN(n9145) );
  OR2_X1 U5615 ( .A1(n5142), .A2(n9961), .ZN(n7043) );
  NAND2_X1 U5616 ( .A1(n6693), .A2(n6436), .ZN(n8054) );
  XNOR2_X1 U5617 ( .A(n8061), .B(n7374), .ZN(n8053) );
  AND2_X1 U5618 ( .A1(n8054), .A2(n8053), .ZN(n8056) );
  NAND2_X1 U5619 ( .A1(n9641), .A2(n9642), .ZN(n9640) );
  OR2_X1 U5620 ( .A1(n6441), .A2(n6440), .ZN(n4494) );
  AND2_X1 U5621 ( .A1(n4494), .A2(n4493), .ZN(n6733) );
  NAND2_X1 U5622 ( .A1(n6731), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4493) );
  NOR2_X1 U5623 ( .A1(n4515), .A2(n4455), .ZN(n9669) );
  INV_X1 U5624 ( .A(n9654), .ZN(n4515) );
  NOR2_X1 U5625 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5446) );
  NAND2_X1 U5626 ( .A1(n4798), .A2(n4796), .ZN(n9239) );
  AOI21_X1 U5627 ( .B1(n4399), .B2(n9103), .A(n4797), .ZN(n4796) );
  INV_X1 U5628 ( .A(n9236), .ZN(n4797) );
  AND2_X1 U5629 ( .A1(n5740), .A2(n5790), .ZN(n9270) );
  NOR2_X1 U5630 ( .A1(n9269), .A2(n9455), .ZN(n9268) );
  NAND2_X1 U5631 ( .A1(n4791), .A2(n8130), .ZN(n4790) );
  NAND2_X1 U5632 ( .A1(n9334), .A2(n4417), .ZN(n4473) );
  INV_X1 U5633 ( .A(n4794), .ZN(n4791) );
  AND2_X1 U5634 ( .A1(n4613), .A2(n9281), .ZN(n4612) );
  OR2_X1 U5635 ( .A1(n5665), .A2(n5664), .ZN(n5690) );
  NOR2_X1 U5636 ( .A1(n9296), .A2(n9297), .ZN(n4794) );
  NAND2_X1 U5637 ( .A1(n9345), .A2(n4615), .ZN(n9308) );
  NAND2_X1 U5638 ( .A1(n8119), .A2(n8962), .ZN(n9319) );
  NAND2_X1 U5639 ( .A1(n9345), .A2(n9333), .ZN(n9327) );
  OR2_X1 U5640 ( .A1(n7948), .A2(n4608), .ZN(n9398) );
  NAND2_X1 U5641 ( .A1(n4609), .A2(n9406), .ZN(n4608) );
  NAND2_X1 U5642 ( .A1(n5483), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5511) );
  INV_X1 U5643 ( .A(n5484), .ZN(n5483) );
  NOR2_X1 U5644 ( .A1(n7948), .A2(n4610), .ZN(n9420) );
  NOR2_X1 U5645 ( .A1(n7948), .A2(n4607), .ZN(n9421) );
  INV_X1 U5646 ( .A(n4609), .ZN(n4607) );
  NOR2_X1 U5647 ( .A1(n9432), .A2(n9431), .ZN(n9435) );
  OR2_X1 U5648 ( .A1(n5456), .A2(n5455), .ZN(n5484) );
  INV_X1 U5649 ( .A(n4779), .ZN(n4778) );
  OAI21_X1 U5650 ( .B1(n4781), .B2(n4780), .A(n9017), .ZN(n4779) );
  INV_X1 U5651 ( .A(n9018), .ZN(n4780) );
  AND2_X1 U5652 ( .A1(n9519), .A2(n9158), .ZN(n7978) );
  OR2_X1 U5653 ( .A1(n5396), .A2(n5395), .ZN(n5430) );
  NAND2_X1 U5654 ( .A1(n5429), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5456) );
  INV_X1 U5655 ( .A(n5430), .ZN(n5429) );
  NOR2_X1 U5656 ( .A1(n7948), .A2(n9519), .ZN(n7983) );
  NAND2_X1 U5657 ( .A1(n4785), .A2(n9004), .ZN(n7951) );
  OR2_X1 U5658 ( .A1(n7851), .A2(n9094), .ZN(n4785) );
  NAND2_X1 U5659 ( .A1(n5370), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5396) );
  INV_X1 U5660 ( .A(n5371), .ZN(n5370) );
  OR2_X1 U5661 ( .A1(n5348), .A2(n5347), .ZN(n5371) );
  NAND2_X1 U5662 ( .A1(n4465), .A2(n4463), .ZN(n7809) );
  INV_X1 U5663 ( .A(n9092), .ZN(n4464) );
  AND2_X1 U5664 ( .A1(n9003), .A2(n8999), .ZN(n9092) );
  INV_X1 U5665 ( .A(n9161), .ZN(n7889) );
  NOR2_X1 U5666 ( .A1(n7599), .A2(n7794), .ZN(n7606) );
  NOR3_X1 U5667 ( .A1(n7599), .A2(n7894), .A3(n7794), .ZN(n7816) );
  NAND2_X1 U5668 ( .A1(n5320), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5348) );
  INV_X1 U5669 ( .A(n5321), .ZN(n5320) );
  OR2_X1 U5670 ( .A1(n9579), .A2(n7658), .ZN(n4921) );
  NAND2_X1 U5671 ( .A1(n5289), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5321) );
  INV_X1 U5672 ( .A(n5291), .ZN(n5289) );
  INV_X1 U5673 ( .A(n9163), .ZN(n7658) );
  OR2_X1 U5674 ( .A1(n5265), .A2(n9986), .ZN(n5291) );
  NAND2_X1 U5675 ( .A1(n5206), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5235) );
  INV_X1 U5676 ( .A(n5207), .ZN(n5206) );
  INV_X1 U5677 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5234) );
  OR2_X1 U5678 ( .A1(n5235), .A2(n5234), .ZN(n5265) );
  NAND2_X1 U5679 ( .A1(n7402), .A2(n8975), .ZN(n4474) );
  AND2_X1 U5680 ( .A1(n7412), .A2(n7411), .ZN(n7453) );
  NOR2_X1 U5681 ( .A1(n7318), .A2(n7485), .ZN(n7412) );
  NAND2_X1 U5682 ( .A1(n7245), .A2(n7202), .ZN(n7317) );
  OR2_X1 U5683 ( .A1(n7317), .A2(n4383), .ZN(n7318) );
  OR2_X1 U5684 ( .A1(n7375), .A2(n7380), .ZN(n7377) );
  NOR2_X1 U5685 ( .A1(n7377), .A2(n7246), .ZN(n7245) );
  NAND2_X1 U5686 ( .A1(n7164), .A2(n8913), .ZN(n9119) );
  INV_X1 U5687 ( .A(n9170), .ZN(n7368) );
  NAND2_X1 U5688 ( .A1(n6974), .A2(n6718), .ZN(n7047) );
  NAND2_X1 U5689 ( .A1(n7052), .A2(n6718), .ZN(n7053) );
  INV_X1 U5690 ( .A(n4718), .ZN(n9075) );
  NAND2_X1 U5691 ( .A1(n5556), .A2(n5555), .ZN(n9493) );
  NAND2_X1 U5692 ( .A1(n5092), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4711) );
  OR2_X1 U5693 ( .A1(n5757), .A2(n7974), .ZN(n9755) );
  XNOR2_X1 U5694 ( .A(n6208), .B(SI_30_), .ZN(n8876) );
  XNOR2_X1 U5695 ( .A(n6201), .B(n6188), .ZN(n8883) );
  NAND2_X1 U5696 ( .A1(n5732), .A2(n5731), .ZN(n6184) );
  AOI21_X1 U5697 ( .B1(n4684), .B2(n4686), .A(n4683), .ZN(n4682) );
  INV_X1 U5698 ( .A(n5603), .ZN(n4683) );
  AND2_X1 U5699 ( .A1(n5632), .A2(n5610), .ZN(n5611) );
  OAI21_X1 U5700 ( .B1(n5568), .B2(n4686), .A(n5572), .ZN(n5605) );
  AOI21_X1 U5701 ( .B1(n4674), .B2(n5498), .A(n4672), .ZN(n4671) );
  INV_X1 U5702 ( .A(n5525), .ZN(n4672) );
  INV_X1 U5703 ( .A(n4674), .ZN(n4673) );
  NAND2_X1 U5704 ( .A1(n4676), .A2(n5502), .ZN(n5527) );
  NAND2_X1 U5705 ( .A1(n5500), .A2(n5499), .ZN(n4676) );
  OAI21_X1 U5706 ( .B1(n5364), .B2(n4397), .A(n4695), .ZN(n5442) );
  NAND2_X1 U5707 ( .A1(n4421), .A2(n4665), .ZN(n5339) );
  AND2_X1 U5708 ( .A1(n5286), .A2(n5314), .ZN(n9185) );
  INV_X1 U5709 ( .A(n5251), .ZN(n4664) );
  INV_X1 U5710 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4940) );
  NAND2_X1 U5711 ( .A1(n4680), .A2(n5178), .ZN(n5196) );
  NAND2_X1 U5712 ( .A1(n5176), .A2(n5175), .ZN(n4680) );
  OR2_X1 U5713 ( .A1(n5089), .A2(n5088), .ZN(n5090) );
  OR2_X1 U5714 ( .A1(n5093), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5147) );
  NAND2_X1 U5715 ( .A1(n4508), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5071) );
  INV_X1 U5716 ( .A(n5044), .ZN(n4508) );
  NAND2_X1 U5717 ( .A1(n4484), .A2(n4482), .ZN(n7465) );
  AOI21_X1 U5718 ( .B1(n7124), .B2(n4387), .A(n4483), .ZN(n4482) );
  NAND2_X1 U5719 ( .A1(n7123), .A2(n4387), .ZN(n4484) );
  INV_X1 U5720 ( .A(n7192), .ZN(n4483) );
  OAI21_X1 U5721 ( .B1(n8250), .B2(n4478), .A(n4476), .ZN(n4481) );
  INV_X1 U5722 ( .A(n4477), .ZN(n4476) );
  OAI21_X1 U5723 ( .B1(n4815), .B2(n4478), .A(n8298), .ZN(n4477) );
  NAND2_X1 U5724 ( .A1(n4806), .A2(n4807), .ZN(n7876) );
  NAND2_X1 U5725 ( .A1(n7538), .A2(n7537), .ZN(n7622) );
  NAND2_X1 U5726 ( .A1(n8250), .A2(n4815), .ZN(n4475) );
  AND4_X1 U5727 ( .A1(n5958), .A2(n5957), .A3(n5956), .A4(n5955), .ZN(n7638)
         );
  NAND2_X1 U5728 ( .A1(n4819), .A2(n6859), .ZN(n6947) );
  INV_X1 U5729 ( .A(n4820), .ZN(n4819) );
  AND2_X1 U5730 ( .A1(n6859), .A2(n6857), .ZN(n6949) );
  NAND2_X1 U5731 ( .A1(n6145), .A2(n6144), .ZN(n8657) );
  NAND2_X1 U5732 ( .A1(n8081), .A2(n8080), .ZN(n8236) );
  AOI21_X1 U5733 ( .B1(n5904), .B2(n5886), .A(n5885), .ZN(n6942) );
  NAND3_X1 U5734 ( .A1(n5884), .A2(n5883), .A3(n5882), .ZN(n5885) );
  NAND2_X1 U5735 ( .A1(n7763), .A2(n7762), .ZN(n4811) );
  AOI21_X1 U5736 ( .B1(n4826), .B2(n4825), .A(n4824), .ZN(n4823) );
  NOR2_X1 U5737 ( .A1(n7620), .A2(n7619), .ZN(n4824) );
  AND2_X1 U5738 ( .A1(n6921), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8293) );
  NAND2_X1 U5739 ( .A1(n4821), .A2(n4387), .ZN(n7193) );
  NAND2_X1 U5740 ( .A1(n4821), .A2(n7129), .ZN(n7134) );
  AND4_X1 U5741 ( .A1(n5936), .A2(n5935), .A3(n5934), .A4(n5933), .ZN(n7469)
         );
  AOI21_X1 U5742 ( .B1(n6863), .B2(n9808), .A(n9810), .ZN(n8247) );
  NAND2_X1 U5743 ( .A1(n4816), .A2(n4815), .ZN(n8299) );
  INV_X1 U5744 ( .A(n8296), .ZN(n8298) );
  INV_X1 U5745 ( .A(n8293), .ZN(n8301) );
  INV_X1 U5746 ( .A(n8247), .ZN(n8308) );
  INV_X1 U5747 ( .A(n8255), .ZN(n8423) );
  OR2_X1 U5748 ( .A1(n6869), .A2(n9844), .ZN(n8314) );
  NAND4_X1 U5749 ( .A1(n5869), .A2(n5868), .A3(n5867), .A4(n5866), .ZN(n6895)
         );
  NOR2_X1 U5750 ( .A1(n6610), .A2(n4450), .ZN(n6601) );
  INV_X1 U5751 ( .A(n4620), .ZN(n6743) );
  NAND2_X1 U5752 ( .A1(n6744), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4619) );
  INV_X1 U5753 ( .A(n4639), .ZN(n7114) );
  NOR2_X1 U5754 ( .A1(n4639), .A2(n4638), .ZN(n7118) );
  AND2_X1 U5755 ( .A1(n7115), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4638) );
  AND2_X1 U5756 ( .A1(n6555), .A2(n6416), .ZN(n8384) );
  XNOR2_X1 U5757 ( .A(n4623), .B(n8373), .ZN(n8369) );
  OAI21_X1 U5758 ( .B1(n8388), .B2(n4653), .A(n8387), .ZN(n4634) );
  INV_X1 U5759 ( .A(n9557), .ZN(n8395) );
  NAND2_X1 U5760 ( .A1(n4751), .A2(n4752), .ZN(n8406) );
  NAND2_X1 U5761 ( .A1(n8400), .A2(n8405), .ZN(n8399) );
  NAND2_X1 U5762 ( .A1(n6156), .A2(n6155), .ZN(n8652) );
  NAND2_X1 U5763 ( .A1(n8463), .A2(n6228), .ZN(n8452) );
  NAND2_X1 U5764 ( .A1(n4874), .A2(n4877), .ZN(n8459) );
  OR2_X1 U5765 ( .A1(n8497), .A2(n4879), .ZN(n4874) );
  AND2_X1 U5766 ( .A1(n6122), .A2(n6121), .ZN(n8486) );
  NAND2_X1 U5767 ( .A1(n4882), .A2(n4880), .ZN(n8479) );
  OR2_X1 U5768 ( .A1(n8497), .A2(n8503), .ZN(n4882) );
  INV_X1 U5769 ( .A(n8679), .ZN(n8521) );
  NAND2_X1 U5770 ( .A1(n4838), .A2(n4842), .ZN(n8514) );
  NAND2_X1 U5771 ( .A1(n4845), .A2(n4843), .ZN(n4838) );
  INV_X1 U5772 ( .A(n4840), .ZN(n4843) );
  NAND2_X1 U5773 ( .A1(n6076), .A2(n6301), .ZN(n8552) );
  NAND2_X1 U5774 ( .A1(n7963), .A2(n6031), .ZN(n7967) );
  AND2_X1 U5775 ( .A1(n4859), .A2(n4408), .ZN(n7933) );
  NAND2_X1 U5776 ( .A1(n4859), .A2(n4858), .ZN(n7955) );
  NAND2_X1 U5777 ( .A1(n4860), .A2(n7682), .ZN(n4859) );
  NAND2_X1 U5778 ( .A1(n7677), .A2(n7676), .ZN(n7744) );
  NAND2_X1 U5779 ( .A1(n4867), .A2(n4870), .ZN(n7387) );
  NAND2_X1 U5780 ( .A1(n7179), .A2(n7178), .ZN(n7386) );
  OR2_X1 U5781 ( .A1(n5901), .A2(n6477), .ZN(n5864) );
  OR2_X1 U5782 ( .A1(n9819), .A2(n6864), .ZN(n8469) );
  OR2_X1 U5783 ( .A1(n6841), .A2(n8148), .ZN(n8475) );
  NAND2_X1 U5784 ( .A1(n5831), .A2(n5836), .ZN(n8749) );
  NAND2_X1 U5785 ( .A1(n5835), .A2(n5834), .ZN(n5836) );
  NAND2_X1 U5786 ( .A1(n5833), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5834) );
  XNOR2_X1 U5787 ( .A(n6407), .B(n5828), .ZN(n7976) );
  INV_X1 U5788 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n10086) );
  INV_X1 U5789 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7835) );
  XNOR2_X1 U5790 ( .A(n6413), .B(n6412), .ZN(n7836) );
  INV_X1 U5791 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7729) );
  INV_X1 U5792 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n10066) );
  XNOR2_X1 U5793 ( .A(n5848), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7581) );
  OR2_X1 U5794 ( .A1(n6068), .A2(n4835), .ZN(n6220) );
  INV_X1 U5795 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7353) );
  INV_X1 U5796 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n9999) );
  INV_X1 U5797 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10188) );
  INV_X1 U5798 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6742) );
  INV_X1 U5799 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6739) );
  INV_X1 U5800 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6683) );
  INV_X1 U5801 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6540) );
  INV_X1 U5802 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6537) );
  INV_X1 U5803 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6509) );
  INV_X1 U5804 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10193) );
  XNOR2_X1 U5805 ( .A(n5878), .B(n4629), .ZN(n6580) );
  NAND2_X1 U5806 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4629) );
  NAND2_X1 U5807 ( .A1(n4914), .A2(n7145), .ZN(n7480) );
  NAND2_X1 U5808 ( .A1(n4914), .A2(n4911), .ZN(n7482) );
  AOI22_X1 U5809 ( .A1(n6974), .A2(n5747), .B1(n5752), .B2(n6718), .ZN(n6717)
         );
  AND2_X1 U5810 ( .A1(n9151), .A2(n5807), .ZN(n8868) );
  NAND2_X1 U5811 ( .A1(n8773), .A2(n5524), .ZN(n8831) );
  NAND2_X1 U5812 ( .A1(n5533), .A2(n5532), .ZN(n9496) );
  INV_X1 U5813 ( .A(n6708), .ZN(n7357) );
  INV_X1 U5814 ( .A(n8819), .ZN(n8870) );
  NAND2_X1 U5815 ( .A1(n4893), .A2(n4527), .ZN(n6422) );
  INV_X1 U5816 ( .A(n4894), .ZN(n4527) );
  NAND2_X1 U5817 ( .A1(n8067), .A2(n8068), .ZN(n8065) );
  AND2_X1 U5818 ( .A1(n5800), .A2(n5779), .ZN(n8850) );
  NAND2_X1 U5819 ( .A1(n5417), .A2(n5416), .ZN(n8064) );
  NAND2_X1 U5820 ( .A1(n5394), .A2(n5393), .ZN(n8073) );
  AND2_X1 U5821 ( .A1(n5789), .A2(n7150), .ZN(n8872) );
  AND3_X1 U5822 ( .A1(n6527), .A2(n6526), .A3(n6525), .ZN(n9219) );
  NAND2_X1 U5823 ( .A1(n5645), .A2(n5644), .ZN(n9338) );
  OAI21_X1 U5824 ( .B1(n9347), .B2(n5692), .A(n5584), .ZN(n9337) );
  NAND2_X1 U5825 ( .A1(n6695), .A2(n6694), .ZN(n6693) );
  NOR2_X1 U5826 ( .A1(n8056), .A2(n4492), .ZN(n9600) );
  AND2_X1 U5827 ( .A1(n8061), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4492) );
  NAND2_X1 U5828 ( .A1(n9640), .A2(n4495), .ZN(n6441) );
  OR2_X1 U5829 ( .A1(n9650), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4495) );
  INV_X1 U5830 ( .A(n4494), .ZN(n6730) );
  INV_X1 U5831 ( .A(n4506), .ZN(n9699) );
  INV_X1 U5832 ( .A(n9196), .ZN(n4505) );
  NAND2_X1 U5833 ( .A1(n8880), .A2(n8879), .ZN(n9445) );
  NAND2_X1 U5834 ( .A1(n9545), .A2(n8882), .ZN(n8880) );
  XNOR2_X1 U5835 ( .A(n4605), .B(n4604), .ZN(n9447) );
  INV_X1 U5836 ( .A(n9445), .ZN(n4604) );
  NOR2_X1 U5837 ( .A1(n9246), .A2(n9563), .ZN(n4605) );
  INV_X1 U5838 ( .A(n9450), .ZN(n9250) );
  OR2_X1 U5839 ( .A1(n9272), .A2(n9242), .ZN(n9233) );
  AND2_X1 U5840 ( .A1(n9267), .A2(n9266), .ZN(n9454) );
  NAND2_X1 U5841 ( .A1(n4453), .A2(n4468), .ZN(n4467) );
  AOI21_X1 U5842 ( .B1(n8132), .B2(n9103), .A(n9389), .ZN(n4469) );
  NAND2_X1 U5843 ( .A1(n4719), .A2(n8123), .ZN(n9227) );
  NAND2_X1 U5844 ( .A1(n9292), .A2(n8122), .ZN(n9276) );
  NAND2_X1 U5845 ( .A1(n9334), .A2(n8897), .ZN(n9312) );
  AND2_X1 U5846 ( .A1(n9356), .A2(n9355), .ZN(n9489) );
  NAND2_X1 U5847 ( .A1(n4725), .A2(n4726), .ZN(n9381) );
  OR2_X1 U5848 ( .A1(n9417), .A2(n4728), .ZN(n4725) );
  AND2_X1 U5849 ( .A1(n4731), .A2(n4730), .ZN(n9397) );
  NAND2_X1 U5850 ( .A1(n4783), .A2(n4781), .ZN(n7980) );
  AND2_X1 U5851 ( .A1(n4714), .A2(n4402), .ZN(n7947) );
  OR2_X1 U5852 ( .A1(n4926), .A2(n7850), .ZN(n4714) );
  NAND2_X1 U5853 ( .A1(n5346), .A2(n5345), .ZN(n7906) );
  NAND2_X1 U5854 ( .A1(n7585), .A2(n7584), .ZN(n7587) );
  NAND2_X1 U5855 ( .A1(n7330), .A2(n7329), .ZN(n7405) );
  NAND2_X1 U5856 ( .A1(n9379), .A2(n7170), .ZN(n9423) );
  NAND2_X1 U5857 ( .A1(n5069), .A2(n9552), .ZN(n4998) );
  INV_X1 U5858 ( .A(n9423), .ZN(n9321) );
  INV_X1 U5859 ( .A(n9247), .ZN(n9414) );
  AOI21_X1 U5860 ( .B1(n9564), .B2(n6718), .A(n7076), .ZN(n7077) );
  AND2_X1 U5861 ( .A1(n6430), .A2(n5775), .ZN(n9756) );
  MUX2_X1 U5862 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4957), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n4959) );
  NAND2_X1 U5863 ( .A1(n4992), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4957) );
  INV_X1 U5864 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7554) );
  INV_X1 U5865 ( .A(n9140), .ZN(n9106) );
  INV_X1 U5866 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7488) );
  NAND2_X1 U5867 ( .A1(n5010), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4978) );
  INV_X1 U5868 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7355) );
  AND2_X1 U5869 ( .A1(n5452), .A2(n5477), .ZN(n9202) );
  INV_X1 U5870 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6955) );
  INV_X1 U5871 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10015) );
  INV_X1 U5872 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6542) );
  INV_X1 U5873 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6536) );
  INV_X1 U5874 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6507) );
  INV_X1 U5875 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6491) );
  NAND2_X1 U5876 ( .A1(n5064), .A2(n5063), .ZN(n5086) );
  XNOR2_X1 U5877 ( .A(n5071), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6692) );
  INV_X1 U5878 ( .A(n4631), .ZN(n6612) );
  INV_X1 U5879 ( .A(n4622), .ZN(n6622) );
  INV_X1 U5880 ( .A(n4625), .ZN(n8365) );
  OAI211_X1 U5881 ( .C1(n8386), .C2(n9812), .A(n4635), .B(n4633), .ZN(P2_U3264) );
  INV_X1 U5882 ( .A(n4634), .ZN(n4633) );
  NAND2_X1 U5883 ( .A1(n4636), .A2(n9812), .ZN(n4635) );
  NOR2_X1 U5884 ( .A1(n8639), .A2(n8600), .ZN(n8217) );
  NAND2_X1 U5885 ( .A1(n4502), .A2(n4496), .ZN(n9216) );
  OAI21_X1 U5886 ( .B1(n4501), .B2(n4497), .A(n9317), .ZN(n4496) );
  CLKBUF_X3 U5887 ( .A(n4601), .Z(n8882) );
  AND2_X1 U5888 ( .A1(n7132), .A2(n7129), .ZN(n4387) );
  INV_X1 U5889 ( .A(n6466), .ZN(n5091) );
  NAND2_X1 U5890 ( .A1(n5277), .A2(n5278), .ZN(n4388) );
  NAND2_X1 U5891 ( .A1(n4665), .A2(n4663), .ZN(n4662) );
  AND2_X1 U5892 ( .A1(n6278), .A2(n6277), .ZN(n7930) );
  XOR2_X1 U5893 ( .A(n6219), .B(n9812), .Z(n4389) );
  AND4_X1 U5894 ( .A1(n4941), .A2(n4940), .A3(n4939), .A4(n10138), .ZN(n4390)
         );
  OR2_X1 U5895 ( .A1(n8193), .A2(n4847), .ZN(n4391) );
  OR2_X1 U5896 ( .A1(n8772), .A2(n8775), .ZN(n8773) );
  AND2_X1 U5897 ( .A1(n4649), .A2(n4648), .ZN(n4392) );
  AND2_X1 U5898 ( .A1(n9573), .A2(n9579), .ZN(n4393) );
  NAND2_X1 U5899 ( .A1(n5454), .A2(n5453), .ZN(n9514) );
  AND2_X1 U5900 ( .A1(n5193), .A2(n5214), .ZN(n4394) );
  AND2_X1 U5901 ( .A1(n4816), .A2(n4446), .ZN(n4395) );
  AND2_X1 U5902 ( .A1(n8300), .A2(n4446), .ZN(n4815) );
  AND2_X1 U5903 ( .A1(n4811), .A2(n4812), .ZN(n7871) );
  NAND2_X1 U5904 ( .A1(n5305), .A2(n5304), .ZN(n7884) );
  OR2_X1 U5905 ( .A1(n7599), .A2(n4606), .ZN(n4396) );
  NAND2_X1 U5906 ( .A1(n7099), .A2(n7101), .ZN(n7100) );
  XNOR2_X1 U5907 ( .A(n5079), .B(n5080), .ZN(n6758) );
  INV_X1 U5909 ( .A(n5904), .ZN(n6160) );
  NAND2_X2 U5910 ( .A1(n9072), .A2(n6982), .ZN(n5049) );
  NAND2_X2 U5911 ( .A1(n6557), .A2(n5634), .ZN(n5901) );
  XNOR2_X1 U5912 ( .A(n6399), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6393) );
  OR2_X1 U5913 ( .A1(n9460), .A2(n9229), .ZN(n9109) );
  OR2_X1 U5914 ( .A1(n5419), .A2(n4697), .ZN(n4397) );
  AOI22_X1 U5915 ( .A1(n9545), .A2(n5947), .B1(P1_DATAO_REG_31__SCAN_IN), .B2(
        n6217), .ZN(n6359) );
  NOR2_X1 U5916 ( .A1(n9390), .A2(n9391), .ZN(n9361) );
  NAND2_X1 U5917 ( .A1(n9319), .A2(n9318), .ZN(n9320) );
  AND2_X1 U5918 ( .A1(n4722), .A2(n4723), .ZN(n4398) );
  AND2_X1 U5919 ( .A1(n9264), .A2(n9109), .ZN(n4399) );
  NAND2_X1 U5920 ( .A1(n5319), .A2(n5318), .ZN(n7894) );
  OAI211_X1 U5921 ( .C1(n5155), .C2(n6476), .A(n5046), .B(n4711), .ZN(n6708)
         );
  AND2_X1 U5922 ( .A1(n7636), .A2(n7635), .ZN(n4400) );
  OR2_X1 U5923 ( .A1(n9472), .A2(n9315), .ZN(n8130) );
  AND2_X1 U5924 ( .A1(n4739), .A2(n6301), .ZN(n4401) );
  NAND2_X1 U5925 ( .A1(n9524), .A2(n9160), .ZN(n4402) );
  OR2_X1 U5926 ( .A1(n8073), .A2(n8030), .ZN(n9013) );
  AND2_X1 U5927 ( .A1(n9098), .A2(n9019), .ZN(n4403) );
  AND2_X1 U5928 ( .A1(n5863), .A2(n4837), .ZN(n5899) );
  OR2_X1 U5929 ( .A1(n8190), .A2(n6300), .ZN(n4404) );
  AND2_X1 U5930 ( .A1(n4917), .A2(n4920), .ZN(n4405) );
  AND2_X1 U5931 ( .A1(n8799), .A2(n8800), .ZN(n4406) );
  AND2_X1 U5932 ( .A1(n8203), .A2(n8202), .ZN(n4407) );
  NAND2_X1 U5933 ( .A1(n9132), .A2(n8887), .ZN(n9318) );
  AND2_X1 U5934 ( .A1(n5771), .A2(n4917), .ZN(n4979) );
  OR2_X1 U5935 ( .A1(n7931), .A2(n8318), .ZN(n4408) );
  AND2_X1 U5936 ( .A1(n4620), .A2(n4619), .ZN(n4409) );
  NAND2_X1 U5937 ( .A1(n5616), .A2(n5615), .ZN(n9481) );
  AND2_X1 U5938 ( .A1(n4744), .A2(n6372), .ZN(n4410) );
  AND4_X1 U5939 ( .A1(n5877), .A2(n5876), .A3(n5875), .A4(n5874), .ZN(n7033)
         );
  AND2_X1 U5940 ( .A1(n4807), .A2(n4805), .ZN(n4411) );
  OR2_X1 U5941 ( .A1(n6355), .A2(n6360), .ZN(n4412) );
  INV_X1 U5942 ( .A(n5706), .ZN(n4891) );
  AND2_X1 U5943 ( .A1(n5705), .A2(n5704), .ZN(n5706) );
  AND2_X1 U5944 ( .A1(n4854), .A2(n6386), .ZN(n4413) );
  INV_X1 U5945 ( .A(n4647), .ZN(n8436) );
  NAND2_X1 U5946 ( .A1(n6337), .A2(n6343), .ZN(n8405) );
  NAND2_X1 U5947 ( .A1(n6005), .A2(n6004), .ZN(n8722) );
  AND2_X1 U5948 ( .A1(n4405), .A2(n4953), .ZN(n4414) );
  NOR2_X1 U5949 ( .A1(n5901), .A2(n6479), .ZN(n4415) );
  OR2_X1 U5950 ( .A1(n6359), .A2(n6361), .ZN(n4416) );
  NAND2_X1 U5951 ( .A1(n9345), .A2(n4613), .ZN(n4616) );
  AND2_X1 U5952 ( .A1(n6304), .A2(n6318), .ZN(n8503) );
  AND2_X1 U5953 ( .A1(n8130), .A2(n4792), .ZN(n4417) );
  AND3_X1 U5954 ( .A1(n4531), .A2(n4530), .A3(n6281), .ZN(n4418) );
  AND2_X1 U5955 ( .A1(n4882), .A2(n4881), .ZN(n4419) );
  INV_X1 U5956 ( .A(n4727), .ZN(n4726) );
  OAI22_X1 U5957 ( .A1(n8115), .A2(n4730), .B1(n9406), .B2(n8866), .ZN(n4727)
         );
  AND2_X1 U5958 ( .A1(n7331), .A2(n7329), .ZN(n4420) );
  INV_X1 U5959 ( .A(n4662), .ZN(n4661) );
  INV_X1 U5960 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9546) );
  OR2_X1 U5961 ( .A1(n5251), .A2(n4666), .ZN(n4421) );
  NOR2_X1 U5962 ( .A1(n8120), .A2(n8767), .ZN(n4422) );
  OR2_X1 U5963 ( .A1(n4535), .A2(n4534), .ZN(n4423) );
  INV_X1 U5964 ( .A(n4847), .ZN(n4846) );
  NOR2_X1 U5965 ( .A1(n8571), .A2(n8554), .ZN(n4847) );
  AND2_X1 U5966 ( .A1(n7874), .A2(n7873), .ZN(n4424) );
  OR2_X1 U5967 ( .A1(n4926), .A2(n4713), .ZN(n4425) );
  NOR2_X1 U5968 ( .A1(n9496), .A2(n9409), .ZN(n4426) );
  AND2_X1 U5969 ( .A1(n5197), .A2(SI_7_), .ZN(n4427) );
  INV_X1 U5970 ( .A(n4667), .ZN(n4666) );
  AND2_X1 U5971 ( .A1(n5283), .A2(n5306), .ZN(n4667) );
  AND4_X1 U5972 ( .A1(n5853), .A2(n5852), .A3(n5851), .A4(n5850), .ZN(n6860)
         );
  INV_X1 U5973 ( .A(n6860), .ZN(n8328) );
  NAND2_X1 U5974 ( .A1(n4795), .A2(n4794), .ZN(n4428) );
  AND2_X1 U5975 ( .A1(n5308), .A2(SI_11_), .ZN(n4429) );
  INV_X1 U5976 ( .A(n4755), .ZN(n4754) );
  NOR2_X1 U5977 ( .A1(n8421), .A2(n4756), .ZN(n4755) );
  AND2_X1 U5978 ( .A1(n9023), .A2(n8964), .ZN(n9418) );
  INV_X1 U5979 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4977) );
  AND2_X1 U5980 ( .A1(n6296), .A2(n8588), .ZN(n8609) );
  NAND2_X1 U5981 ( .A1(n9022), .A2(n9023), .ZN(n4430) );
  OR2_X1 U5982 ( .A1(n8641), .A2(n8202), .ZN(n6337) );
  AND2_X1 U5983 ( .A1(n9103), .A2(n8123), .ZN(n4431) );
  NOR2_X1 U5984 ( .A1(n9082), .A2(n7214), .ZN(n4432) );
  NAND2_X1 U5985 ( .A1(n4893), .A2(n4892), .ZN(n4433) );
  AND2_X1 U5986 ( .A1(n6262), .A2(n7391), .ZN(n4434) );
  NOR2_X1 U5987 ( .A1(n7621), .A2(n4827), .ZN(n4435) );
  AND2_X1 U5988 ( .A1(n6230), .A2(n6323), .ZN(n8197) );
  INV_X1 U5989 ( .A(n8197), .ZN(n8488) );
  AND2_X1 U5990 ( .A1(n5195), .A2(n5175), .ZN(n4436) );
  NOR2_X1 U5991 ( .A1(n4938), .A2(n4810), .ZN(n4809) );
  AND2_X1 U5992 ( .A1(n7586), .A2(n7584), .ZN(n4437) );
  NAND2_X1 U5993 ( .A1(n5687), .A2(n5686), .ZN(n9465) );
  AND2_X1 U5994 ( .A1(n5467), .A2(n4520), .ZN(n4438) );
  AND2_X1 U5995 ( .A1(n4392), .A2(n8521), .ZN(n4439) );
  AND2_X1 U5996 ( .A1(n7932), .A2(n4408), .ZN(n4858) );
  INV_X1 U5997 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5861) );
  INV_X1 U5998 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4985) );
  INV_X1 U5999 ( .A(n4766), .ZN(n4765) );
  NAND2_X1 U6000 ( .A1(n4767), .A2(n6278), .ZN(n4766) );
  INV_X1 U6001 ( .A(n4761), .ZN(n4760) );
  NAND2_X1 U6002 ( .A1(n6366), .A2(n6239), .ZN(n4761) );
  INV_X1 U6003 ( .A(n4738), .ZN(n4737) );
  NAND2_X1 U6004 ( .A1(n4401), .A2(n6316), .ZN(n4738) );
  INV_X1 U6005 ( .A(n4772), .ZN(n4771) );
  NAND2_X1 U6006 ( .A1(n8609), .A2(n6290), .ZN(n4772) );
  INV_X1 U6007 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5833) );
  INV_X1 U6008 ( .A(n4905), .ZN(n4904) );
  OR2_X1 U6009 ( .A1(n7898), .A2(n4906), .ZN(n4905) );
  INV_X1 U6010 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4836) );
  INV_X1 U6011 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4953) );
  NAND2_X1 U6012 ( .A1(n6984), .A2(n5000), .ZN(n5630) );
  NAND2_X1 U6013 ( .A1(n5663), .A2(n5662), .ZN(n9472) );
  INV_X1 U6014 ( .A(n9472), .ZN(n4614) );
  NAND2_X1 U6015 ( .A1(n4937), .A2(n5983), .ZN(n7680) );
  AND3_X1 U6016 ( .A1(n4829), .A2(n8014), .A3(n8038), .ZN(n4440) );
  XOR2_X1 U6017 ( .A(n8662), .B(n8163), .Z(n4441) );
  OR2_X1 U6018 ( .A1(n7685), .A2(n7931), .ZN(n4442) );
  OR2_X1 U6019 ( .A1(n8696), .A2(n8589), .ZN(n4443) );
  OR2_X1 U6020 ( .A1(n8147), .A2(n8251), .ZN(n4444) );
  OR2_X1 U6021 ( .A1(n5680), .A2(n4703), .ZN(n4445) );
  NAND2_X1 U6022 ( .A1(n5844), .A2(n5845), .ZN(n6043) );
  OR2_X1 U6023 ( .A1(n8252), .A2(n4818), .ZN(n4446) );
  OAI21_X1 U6024 ( .B1(n7613), .B2(n7612), .A(n8921), .ZN(n7804) );
  NOR2_X1 U6025 ( .A1(n9435), .A2(n8128), .ZN(n9407) );
  NAND2_X1 U6026 ( .A1(n7885), .A2(n5336), .ZN(n7897) );
  OAI21_X1 U6027 ( .B1(n6042), .B2(n4769), .A(n4768), .ZN(n8572) );
  NAND2_X1 U6028 ( .A1(n5288), .A2(n5287), .ZN(n7794) );
  NAND2_X1 U6029 ( .A1(n6169), .A2(n6168), .ZN(n8646) );
  INV_X1 U6030 ( .A(n8646), .ZN(n4646) );
  NAND2_X1 U6031 ( .A1(n8013), .A2(n8012), .ZN(n8038) );
  OR2_X1 U6032 ( .A1(n7884), .A2(n7887), .ZN(n7885) );
  INV_X1 U6033 ( .A(n5498), .ZN(n5499) );
  AND2_X1 U6034 ( .A1(n6000), .A2(n6278), .ZN(n4447) );
  NAND2_X1 U6035 ( .A1(n8235), .A2(n8234), .ZN(n4448) );
  AND2_X1 U6036 ( .A1(n4506), .A2(n4505), .ZN(n4449) );
  AND2_X1 U6037 ( .A1(n6578), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4450) );
  AND2_X1 U6038 ( .A1(n8722), .A2(n8317), .ZN(n4451) );
  INV_X1 U6039 ( .A(n4642), .ZN(n7996) );
  NOR2_X1 U6040 ( .A1(n7685), .A2(n4644), .ZN(n4642) );
  NAND2_X1 U6041 ( .A1(n8580), .A2(n8188), .ZN(n8582) );
  NAND2_X1 U6042 ( .A1(n5448), .A2(n5447), .ZN(n4452) );
  NAND2_X1 U6043 ( .A1(n9299), .A2(n9437), .ZN(n4453) );
  AND2_X1 U6044 ( .A1(n7707), .A2(n7635), .ZN(n4454) );
  OR2_X1 U6045 ( .A1(n6393), .A2(n7581), .ZN(n6394) );
  INV_X1 U6046 ( .A(n6394), .ZN(n4489) );
  AND2_X1 U6047 ( .A1(n9661), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4455) );
  AND2_X1 U6048 ( .A1(n6186), .A2(n6185), .ZN(n4456) );
  OAI21_X1 U6049 ( .B1(n5894), .B2(n4758), .A(n4757), .ZN(n7090) );
  NAND2_X1 U6050 ( .A1(n5428), .A2(n5427), .ZN(n9519) );
  INV_X1 U6051 ( .A(n9519), .ZN(n4611) );
  NAND2_X1 U6052 ( .A1(n5894), .A2(n6239), .ZN(n6822) );
  INV_X1 U6053 ( .A(n7932), .ZN(n4767) );
  NAND2_X1 U6054 ( .A1(n6091), .A2(n6090), .ZN(n8686) );
  INV_X1 U6055 ( .A(n8686), .ZN(n4648) );
  INV_X1 U6056 ( .A(n5915), .ZN(n6172) );
  AND2_X1 U6057 ( .A1(n5137), .A2(n5138), .ZN(n7099) );
  NAND2_X1 U6058 ( .A1(n7731), .A2(n7730), .ZN(n7763) );
  NAND2_X1 U6059 ( .A1(n5894), .A2(n4760), .ZN(n7257) );
  AND2_X1 U6060 ( .A1(n6785), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4457) );
  AND2_X1 U6061 ( .A1(n4511), .A2(n4510), .ZN(n4458) );
  NAND2_X1 U6062 ( .A1(n9191), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4459) );
  INV_X1 U6063 ( .A(n8342), .ZN(n4628) );
  NAND2_X1 U6064 ( .A1(n5859), .A2(n5858), .ZN(n6416) );
  OAI21_X1 U6065 ( .B1(n6910), .B2(n6909), .A(n6908), .ZN(n6929) );
  NAND2_X1 U6066 ( .A1(n6833), .A2(n6892), .ZN(n6891) );
  NAND2_X1 U6067 ( .A1(n7048), .A2(n7047), .ZN(n7049) );
  NAND2_X1 U6068 ( .A1(n8148), .A2(n6824), .ZN(n4460) );
  NAND2_X1 U6069 ( .A1(n5161), .A2(n5162), .ZN(n4461) );
  INV_X1 U6070 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5347) );
  NAND2_X1 U6071 ( .A1(n6394), .A2(n6825), .ZN(n4462) );
  INV_X1 U6072 ( .A(n7320), .ZN(n4472) );
  INV_X1 U6073 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4653) );
  OR2_X2 U6074 ( .A1(n6393), .A2(n6229), .ZN(n6360) );
  OAI21_X1 U6075 ( .B1(n7804), .B2(n4466), .A(n8989), .ZN(n7810) );
  AOI21_X1 U6076 ( .B1(n4466), .B2(n8989), .A(n4464), .ZN(n4463) );
  NAND2_X1 U6077 ( .A1(n7804), .A2(n8989), .ZN(n4465) );
  OR2_X2 U6078 ( .A1(n8132), .A2(n9103), .ZN(n4799) );
  INV_X4 U6079 ( .A(n5098), .ZN(n5692) );
  NAND3_X1 U6080 ( .A1(n5146), .A2(n4470), .A3(n5144), .ZN(n9168) );
  AND2_X1 U6081 ( .A1(n5145), .A2(n4471), .ZN(n4470) );
  NAND2_X1 U6082 ( .A1(n5098), .A2(n4472), .ZN(n4471) );
  AND2_X2 U6083 ( .A1(n5771), .A2(n4414), .ZN(n4993) );
  NAND4_X1 U6084 ( .A1(n4414), .A2(n4971), .A3(n4951), .A4(n4990), .ZN(n4992)
         );
  NAND2_X1 U6085 ( .A1(n4475), .A2(n4813), .ZN(n8156) );
  NAND2_X1 U6086 ( .A1(n8177), .A2(n4480), .ZN(n8161) );
  INV_X1 U6087 ( .A(n4481), .ZN(n4480) );
  NAND3_X1 U6088 ( .A1(n5844), .A2(n5846), .A3(n4836), .ZN(n4491) );
  XNOR2_X1 U6089 ( .A(n9195), .B(n9194), .ZN(n9701) );
  INV_X1 U6090 ( .A(n4516), .ZN(n5012) );
  OAI21_X1 U6091 ( .B1(n6637), .B2(n4516), .A(n6638), .ZN(n6685) );
  NAND2_X1 U6092 ( .A1(n6637), .A2(n4516), .ZN(n6638) );
  OAI21_X1 U6093 ( .B1(n5305), .B2(n4905), .A(n4517), .ZN(n5406) );
  OAI21_X2 U6094 ( .B1(n5010), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n4975) );
  NAND3_X1 U6095 ( .A1(n4523), .A2(n4522), .A3(n4438), .ZN(n8811) );
  NAND3_X1 U6096 ( .A1(n4523), .A2(n4522), .A3(n4520), .ZN(n8810) );
  NAND2_X1 U6097 ( .A1(n7099), .A2(n4525), .ZN(n4524) );
  NAND3_X1 U6098 ( .A1(n4524), .A2(n4910), .A3(n5193), .ZN(n5219) );
  NAND3_X1 U6099 ( .A1(n4524), .A2(n4910), .A3(n4394), .ZN(n7695) );
  NOR2_X1 U6100 ( .A1(n4912), .A2(n4526), .ZN(n4525) );
  NAND4_X1 U6101 ( .A1(n6263), .A2(n4536), .A3(n6273), .A4(n4434), .ZN(n4530)
         );
  INV_X1 U6102 ( .A(n6374), .ZN(n4535) );
  INV_X1 U6103 ( .A(n6282), .ZN(n4536) );
  NAND3_X1 U6104 ( .A1(n4541), .A2(n4540), .A3(n7010), .ZN(n4539) );
  XNOR2_X1 U6105 ( .A(n5083), .B(n4542), .ZN(n5088) );
  NAND2_X1 U6106 ( .A1(n5091), .A2(n6484), .ZN(n4544) );
  NAND2_X1 U6107 ( .A1(n4549), .A2(n4545), .ZN(n6308) );
  OR2_X1 U6108 ( .A1(n4550), .A2(n6360), .ZN(n4549) );
  AOI21_X1 U6109 ( .B1(n4555), .B2(n4554), .A(n4552), .ZN(n6335) );
  NAND2_X1 U6110 ( .A1(n6326), .A2(n6360), .ZN(n4553) );
  NAND2_X1 U6111 ( .A1(n6324), .A2(n6360), .ZN(n4554) );
  OAI22_X1 U6112 ( .A1(n6321), .A2(n4557), .B1(n6360), .B2(n6322), .ZN(n4556)
         );
  NAND2_X1 U6113 ( .A1(n4559), .A2(n4558), .ZN(n4557) );
  NAND2_X1 U6114 ( .A1(n8489), .A2(n6360), .ZN(n4558) );
  NAND2_X1 U6115 ( .A1(n4560), .A2(n4971), .ZN(n4564) );
  NAND2_X1 U6116 ( .A1(n4563), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n4562) );
  OR2_X1 U6117 ( .A1(n9012), .A2(n4575), .ZN(n4569) );
  NAND2_X1 U6118 ( .A1(n9012), .A2(n4572), .ZN(n4571) );
  NAND2_X1 U6119 ( .A1(n7164), .A2(n4590), .ZN(n7240) );
  NAND2_X1 U6120 ( .A1(n7240), .A2(n7221), .ZN(n7165) );
  AOI21_X1 U6121 ( .B1(n4598), .B2(n9070), .A(n4597), .ZN(n4596) );
  NOR2_X2 U6122 ( .A1(n6718), .A2(n7348), .ZN(n7058) );
  NAND2_X1 U6123 ( .A1(n9345), .A2(n4612), .ZN(n9277) );
  INV_X1 U6124 ( .A(n4616), .ZN(n9302) );
  OR2_X1 U6125 ( .A1(n6467), .A2(n5921), .ZN(n5879) );
  NAND2_X2 U6126 ( .A1(n6416), .A2(n8212), .ZN(n6557) );
  INV_X1 U6127 ( .A(n4641), .ZN(n8623) );
  NOR2_X2 U6128 ( .A1(n8480), .A2(n8662), .ZN(n8468) );
  NAND2_X1 U6129 ( .A1(n8596), .A2(n4439), .ZN(n8515) );
  NAND2_X1 U6130 ( .A1(n4658), .A2(n4412), .ZN(n4657) );
  NAND2_X1 U6131 ( .A1(n6388), .A2(n6360), .ZN(n4658) );
  OAI21_X1 U6132 ( .B1(n5500), .B2(n4673), .A(n4671), .ZN(n5552) );
  NAND2_X1 U6133 ( .A1(n4670), .A2(n4668), .ZN(n5554) );
  NAND2_X1 U6134 ( .A1(n5500), .A2(n4671), .ZN(n4670) );
  NAND2_X1 U6135 ( .A1(n5176), .A2(n4436), .ZN(n4677) );
  NAND2_X1 U6136 ( .A1(n4677), .A2(n4678), .ZN(n5222) );
  NAND2_X1 U6137 ( .A1(n5568), .A2(n4684), .ZN(n4681) );
  NAND2_X1 U6138 ( .A1(n4681), .A2(n4682), .ZN(n5612) );
  NAND2_X1 U6139 ( .A1(n5716), .A2(n5715), .ZN(n5732) );
  OAI21_X1 U6140 ( .B1(n5715), .B2(n4691), .A(n6183), .ZN(n4690) );
  NAND2_X1 U6141 ( .A1(n5364), .A2(n4695), .ZN(n4692) );
  NAND2_X1 U6142 ( .A1(n4692), .A2(n4693), .ZN(n5444) );
  NAND2_X1 U6143 ( .A1(n5364), .A2(n4699), .ZN(n4698) );
  NAND2_X1 U6144 ( .A1(n5364), .A2(n5363), .ZN(n5386) );
  NAND2_X1 U6145 ( .A1(n5633), .A2(n4705), .ZN(n4704) );
  NAND2_X1 U6146 ( .A1(n5633), .A2(n5632), .ZN(n5654) );
  OAI21_X2 U6147 ( .B1(n5476), .B2(n5475), .A(n5474), .ZN(n5500) );
  INV_X1 U6148 ( .A(n9146), .ZN(n9147) );
  XNOR2_X1 U6149 ( .A(n5065), .B(SI_2_), .ZN(n5063) );
  AND2_X1 U6150 ( .A1(n5084), .A2(n5087), .ZN(n5085) );
  NAND2_X1 U6151 ( .A1(n5612), .A2(n5611), .ZN(n5633) );
  NAND2_X1 U6152 ( .A1(n5444), .A2(n5443), .ZN(n5476) );
  NAND2_X1 U6153 ( .A1(n5554), .A2(n5553), .ZN(n5568) );
  NAND2_X1 U6154 ( .A1(n5362), .A2(n4933), .ZN(n5364) );
  INV_X1 U6155 ( .A(n9294), .ZN(n8121) );
  OAI21_X1 U6156 ( .B1(n5798), .B2(n5634), .A(n4709), .ZN(n5092) );
  NAND2_X1 U6157 ( .A1(n4994), .A2(n4710), .ZN(n4709) );
  NAND2_X1 U6158 ( .A1(n7800), .A2(n4712), .ZN(n4717) );
  NAND2_X1 U6159 ( .A1(n7357), .A2(n6719), .ZN(n8914) );
  NAND3_X1 U6160 ( .A1(n4718), .A2(n7047), .A3(n7048), .ZN(n7156) );
  NAND2_X1 U6161 ( .A1(n9077), .A2(n6976), .ZN(n7048) );
  NAND2_X1 U6162 ( .A1(n7585), .A2(n4437), .ZN(n7605) );
  NAND2_X1 U6163 ( .A1(n4719), .A2(n4431), .ZN(n9263) );
  NAND2_X1 U6164 ( .A1(n9417), .A2(n4724), .ZN(n4722) );
  INV_X1 U6165 ( .A(n4731), .ZN(n9416) );
  NAND2_X1 U6166 ( .A1(n6251), .A2(n6250), .ZN(n6882) );
  NAND2_X1 U6167 ( .A1(n6953), .A2(n9847), .ZN(n7032) );
  NAND2_X1 U6168 ( .A1(n4733), .A2(n4736), .ZN(n8524) );
  NAND2_X1 U6169 ( .A1(n6076), .A2(n4737), .ZN(n4733) );
  AOI21_X1 U6170 ( .B1(n4736), .B2(n4738), .A(n4735), .ZN(n4734) );
  AND2_X2 U6171 ( .A1(n4749), .A2(n4746), .ZN(n8209) );
  NAND2_X1 U6172 ( .A1(n4936), .A2(n6167), .ZN(n8432) );
  AOI21_X1 U6173 ( .B1(n4761), .B2(n6235), .A(n4759), .ZN(n4757) );
  INV_X1 U6174 ( .A(n6235), .ZN(n4758) );
  OAI21_X2 U6175 ( .B1(n6000), .B2(n4763), .A(n4762), .ZN(n8000) );
  AOI21_X1 U6176 ( .B1(n6031), .B2(n4766), .A(n4764), .ZN(n4762) );
  INV_X1 U6177 ( .A(n6031), .ZN(n4763) );
  AOI21_X1 U6178 ( .B1(n4772), .B2(n6067), .A(n4770), .ZN(n4768) );
  NAND2_X1 U6179 ( .A1(n4773), .A2(n4774), .ZN(n6154) );
  NAND2_X1 U6180 ( .A1(n8461), .A2(n6228), .ZN(n4773) );
  NAND4_X1 U6181 ( .A1(n4864), .A2(n5844), .A3(n5845), .A4(n5828), .ZN(n5860)
         );
  NAND3_X1 U6182 ( .A1(n4864), .A2(n5844), .A3(n5845), .ZN(n6405) );
  NAND2_X1 U6183 ( .A1(n5042), .A2(n5041), .ZN(n5064) );
  NAND2_X1 U6184 ( .A1(n4787), .A2(n5042), .ZN(n4786) );
  AND2_X1 U6185 ( .A1(n5085), .A2(n5041), .ZN(n4787) );
  NAND2_X1 U6186 ( .A1(n4789), .A2(n5085), .ZN(n4788) );
  INV_X1 U6187 ( .A(n5063), .ZN(n4789) );
  INV_X1 U6188 ( .A(n4795), .ZN(n9311) );
  NAND2_X1 U6189 ( .A1(n8132), .A2(n4399), .ZN(n4798) );
  NAND2_X1 U6190 ( .A1(n4799), .A2(n4399), .ZN(n9256) );
  OAI21_X2 U6191 ( .B1(n9432), .B2(n4802), .A(n4800), .ZN(n9390) );
  OAI21_X1 U6192 ( .B1(n9408), .B2(n8964), .A(n9025), .ZN(n4801) );
  INV_X1 U6193 ( .A(n9408), .ZN(n4803) );
  NAND3_X1 U6194 ( .A1(n4804), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4996) );
  INV_X1 U6195 ( .A(n4938), .ZN(n4812) );
  NAND2_X1 U6196 ( .A1(n4820), .A2(n6859), .ZN(n6910) );
  NAND2_X1 U6197 ( .A1(n7505), .A2(n4435), .ZN(n4822) );
  NAND2_X1 U6198 ( .A1(n4822), .A2(n4823), .ZN(n7731) );
  NAND2_X1 U6199 ( .A1(n4829), .A2(n8038), .ZN(n8015) );
  NAND2_X1 U6200 ( .A1(n8081), .A2(n4831), .ZN(n8235) );
  NOR2_X1 U6201 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4837) );
  NAND2_X1 U6202 ( .A1(n8413), .A2(n4849), .ZN(n4848) );
  NAND2_X1 U6203 ( .A1(n8413), .A2(n8201), .ZN(n8400) );
  OAI211_X1 U6204 ( .C1(n8413), .C2(n4853), .A(n4851), .B(n4848), .ZN(n8640)
         );
  NAND2_X1 U6205 ( .A1(n7929), .A2(n4858), .ZN(n4856) );
  NAND2_X1 U6206 ( .A1(n4856), .A2(n4857), .ZN(n7993) );
  NAND2_X1 U6207 ( .A1(n6891), .A2(n4861), .ZN(n6878) );
  NAND2_X1 U6208 ( .A1(n8186), .A2(n4862), .ZN(n8580) );
  AND2_X1 U6209 ( .A1(n5824), .A2(n5826), .ZN(n4863) );
  NAND2_X1 U6210 ( .A1(n7179), .A2(n4868), .ZN(n4867) );
  NAND2_X1 U6211 ( .A1(n8497), .A2(n4877), .ZN(n4876) );
  NAND2_X1 U6212 ( .A1(n4886), .A2(n4885), .ZN(n6770) );
  OAI211_X1 U6213 ( .C1(n4886), .C2(n4884), .A(n4883), .B(n5133), .ZN(n5137)
         );
  NAND2_X1 U6214 ( .A1(n6769), .A2(n5134), .ZN(n4883) );
  INV_X1 U6215 ( .A(n5134), .ZN(n4884) );
  INV_X1 U6216 ( .A(n6769), .ZN(n4885) );
  INV_X1 U6217 ( .A(n6768), .ZN(n4886) );
  INV_X1 U6218 ( .A(n4887), .ZN(n8754) );
  AOI21_X1 U6219 ( .B1(n8823), .B2(n8824), .A(n4929), .ZN(n8790) );
  NAND2_X1 U6220 ( .A1(n8772), .A2(n5524), .ZN(n4909) );
  INV_X1 U6221 ( .A(n4912), .ZN(n4911) );
  NAND2_X1 U6222 ( .A1(n7100), .A2(n5138), .ZN(n7144) );
  NAND2_X1 U6223 ( .A1(n5771), .A2(n10082), .ZN(n4984) );
  NAND2_X1 U6224 ( .A1(n8118), .A2(n4925), .ZN(n9326) );
  NAND2_X1 U6225 ( .A1(n9344), .A2(n8117), .ZN(n8118) );
  NAND2_X1 U6226 ( .A1(n9256), .A2(n4919), .ZN(n9261) );
  NAND2_X1 U6227 ( .A1(n4433), .A2(n6423), .ZN(n6429) );
  OAI222_X1 U6228 ( .A1(P2_U3152), .A2(n8180), .B1(n8747), .B2(n8221), .C1(
        n8179), .C2(n7728), .ZN(P2_U3328) );
  NAND2_X1 U6229 ( .A1(n6834), .A2(n9852), .ZN(n6365) );
  OAI21_X1 U6230 ( .B1(n5857), .B2(n5832), .A(P2_IR_REG_29__SCAN_IN), .ZN(
        n5835) );
  OR2_X1 U6231 ( .A1(n6394), .A2(n9953), .ZN(n9900) );
  OR2_X1 U6232 ( .A1(n5069), .A2(n5045), .ZN(n5046) );
  INV_X1 U6233 ( .A(n7181), .ZN(n7182) );
  NAND2_X1 U6234 ( .A1(n7033), .A2(n4386), .ZN(n6364) );
  NAND2_X1 U6235 ( .A1(n4993), .A2(n4954), .ZN(n4958) );
  OR2_X1 U6236 ( .A1(n8145), .A2(n4441), .ZN(n8146) );
  OR2_X1 U6237 ( .A1(n7455), .A2(n7664), .ZN(n7599) );
  INV_X1 U6238 ( .A(n6179), .ZN(n6194) );
  NAND2_X1 U6239 ( .A1(n6705), .A2(n5056), .ZN(n6760) );
  INV_X1 U6240 ( .A(n8641), .ZN(n8203) );
  OR2_X1 U6241 ( .A1(n9449), .A2(n9776), .ZN(n4918) );
  OR2_X1 U6242 ( .A1(n9255), .A2(n9264), .ZN(n4919) );
  INV_X1 U6243 ( .A(n9786), .ZN(n9787) );
  AND2_X1 U6244 ( .A1(n4980), .A2(n4952), .ZN(n4920) );
  OR2_X1 U6245 ( .A1(n8142), .A2(n8141), .ZN(n4922) );
  NAND2_X1 U6246 ( .A1(n8842), .A2(n5594), .ZN(n8844) );
  INV_X1 U6247 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4999) );
  OR2_X1 U6248 ( .A1(n9216), .A2(n9215), .ZN(P1_U3260) );
  NAND2_X1 U6249 ( .A1(n4918), .A2(n4930), .ZN(n4924) );
  OR2_X1 U6250 ( .A1(n9350), .A2(n9370), .ZN(n4925) );
  AND2_X1 U6251 ( .A1(n7849), .A2(n8904), .ZN(n4926) );
  NOR2_X1 U6252 ( .A1(n8237), .A2(n8094), .ZN(n4928) );
  AND2_X1 U6253 ( .A1(n5651), .A2(n5650), .ZN(n4929) );
  OR2_X1 U6254 ( .A1(n9250), .A2(n9774), .ZN(n4930) );
  AOI21_X1 U6255 ( .B1(n8403), .B2(n5904), .A(n6182), .ZN(n8202) );
  NOR2_X1 U6256 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n4932) );
  AND2_X1 U6257 ( .A1(n5363), .A2(n5343), .ZN(n4933) );
  AND2_X1 U6258 ( .A1(n9139), .A2(n9073), .ZN(n4934) );
  NAND2_X1 U6259 ( .A1(n5671), .A2(n5670), .ZN(n9288) );
  INV_X1 U6260 ( .A(n9288), .ZN(n9315) );
  NAND2_X1 U6261 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n4935) );
  NAND2_X1 U6262 ( .A1(n5032), .A2(n5033), .ZN(n6714) );
  AND2_X1 U6263 ( .A1(n6154), .A2(n6327), .ZN(n4936) );
  INV_X1 U6264 ( .A(n9085), .ZN(n7331) );
  INV_X1 U6265 ( .A(n8073), .ZN(n7855) );
  INV_X1 U6266 ( .A(n8125), .ZN(n9269) );
  NOR2_X1 U6267 ( .A1(n9277), .A2(n9460), .ZN(n8125) );
  AOI21_X1 U6268 ( .B1(n8104), .B2(n8105), .A(n8098), .ZN(n8139) );
  NOR2_X1 U6269 ( .A1(n7761), .A2(n7760), .ZN(n4938) );
  INV_X1 U6270 ( .A(n9922), .ZN(n9919) );
  OR3_X1 U6271 ( .A1(n6874), .A2(n6862), .A3(n9868), .ZN(n8296) );
  AND2_X1 U6272 ( .A1(n9059), .A2(n9109), .ZN(n9055) );
  INV_X1 U6273 ( .A(n5218), .ZN(n5214) );
  INV_X1 U6274 ( .A(n9062), .ZN(n9063) );
  INV_X1 U6275 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4990) );
  AND2_X1 U6276 ( .A1(n7223), .A2(n7221), .ZN(n9120) );
  INV_X1 U6277 ( .A(n6008), .ZN(n6006) );
  INV_X1 U6278 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5930) );
  INV_X1 U6279 ( .A(n6261), .ZN(n5937) );
  INV_X1 U6280 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5340) );
  INV_X1 U6281 ( .A(n6124), .ZN(n6123) );
  INV_X1 U6282 ( .A(n8460), .ZN(n6143) );
  NAND2_X1 U6283 ( .A1(n6006), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6024) );
  INV_X1 U6284 ( .A(n8429), .ZN(n6167) );
  INV_X1 U6285 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5828) );
  INV_X1 U6286 ( .A(n5053), .ZN(n5051) );
  AND2_X1 U6287 ( .A1(n9072), .A2(n9140), .ZN(n9073) );
  INV_X1 U6288 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9986) );
  OR2_X1 U6289 ( .A1(n5069), .A2(n6510), .ZN(n5026) );
  INV_X1 U6290 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4974) );
  INV_X1 U6291 ( .A(SI_9_), .ZN(n10074) );
  INV_X1 U6292 ( .A(n6158), .ZN(n6157) );
  AND2_X1 U6293 ( .A1(n8097), .A2(n8096), .ZN(n8098) );
  OR2_X1 U6294 ( .A1(n6135), .A2(n6134), .ZN(n6147) );
  INV_X1 U6295 ( .A(n7504), .ZN(n7502) );
  INV_X1 U6296 ( .A(n8016), .ZN(n8014) );
  OR3_X1 U6297 ( .A1(n6177), .A2(n8157), .A3(n6176), .ZN(n6191) );
  NAND2_X1 U6298 ( .A1(n6123), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6135) );
  INV_X1 U6299 ( .A(n8749), .ZN(n5849) );
  OR2_X1 U6300 ( .A1(n8657), .A2(n8433), .ZN(n8199) );
  AND2_X1 U6301 ( .A1(n5941), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5967) );
  AND3_X1 U6302 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n5916) );
  INV_X1 U6303 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5829) );
  NAND2_X1 U6304 ( .A1(n5855), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5856) );
  INV_X1 U6305 ( .A(n8813), .ZN(n5467) );
  NAND2_X1 U6306 ( .A1(n8811), .A2(n5470), .ZN(n5493) );
  OR2_X1 U6307 ( .A1(n5677), .A2(n5676), .ZN(n5678) );
  NAND2_X1 U6308 ( .A1(n5778), .A2(n9140), .ZN(n6997) );
  NAND2_X1 U6309 ( .A1(n5422), .A2(n5421), .ZN(n5443) );
  NAND2_X1 U6310 ( .A1(n5341), .A2(n9970), .ZN(n5363) );
  NAND2_X1 U6311 ( .A1(n6157), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6177) );
  INV_X1 U6312 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8346) );
  OR2_X1 U6313 ( .A1(n6060), .A2(n8346), .ZN(n6083) );
  INV_X1 U6314 ( .A(n7133), .ZN(n7132) );
  AND2_X1 U6315 ( .A1(n6178), .A2(n6191), .ZN(n8403) );
  INV_X1 U6316 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7625) );
  INV_X1 U6317 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10068) );
  INV_X1 U6318 ( .A(n8589), .ZN(n8554) );
  NAND2_X1 U6319 ( .A1(n7634), .A2(n7633), .ZN(n7707) );
  AND2_X1 U6320 ( .A1(n6265), .A2(n6264), .ZN(n7391) );
  OAI21_X1 U6321 ( .B1(n7252), .B2(n7089), .A(n7088), .ZN(n7176) );
  NAND2_X1 U6322 ( .A1(n6239), .A2(n6234), .ZN(n6961) );
  INV_X1 U6323 ( .A(n9900), .ZN(n9869) );
  NOR2_X1 U6324 ( .A1(n9900), .A2(n6227), .ZN(n7007) );
  INV_X1 U6325 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6222) );
  OR2_X1 U6326 ( .A1(n5950), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5987) );
  OR2_X1 U6327 ( .A1(n5912), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5926) );
  AND2_X1 U6328 ( .A1(n8752), .A2(n8850), .ZN(n5785) );
  AND2_X1 U6329 ( .A1(n5602), .A2(n5601), .ZN(n8846) );
  AND2_X1 U6330 ( .A1(n5055), .A2(n5056), .ZN(n6707) );
  INV_X1 U6331 ( .A(n5776), .ZN(n5778) );
  AND2_X1 U6332 ( .A1(n5690), .A2(n5666), .ZN(n9303) );
  INV_X1 U6333 ( .A(n6506), .ZN(n6731) );
  OR3_X1 U6334 ( .A1(n9741), .A2(n9740), .A3(n9739), .ZN(n9743) );
  INV_X1 U6335 ( .A(n9337), .ZN(n9370) );
  INV_X1 U6336 ( .A(n9514), .ZN(n8816) );
  NAND2_X1 U6337 ( .A1(n7856), .A2(n7855), .ZN(n7948) );
  AND2_X1 U6338 ( .A1(n7894), .A2(n9162), .ZN(n7797) );
  INV_X1 U6339 ( .A(n9317), .ZN(n7289) );
  INV_X1 U6340 ( .A(n9776), .ZN(n9502) );
  INV_X1 U6341 ( .A(n7906), .ZN(n9573) );
  OR2_X1 U6342 ( .A1(n6997), .A2(n5798), .ZN(n9369) );
  AND2_X1 U6343 ( .A1(n6994), .A2(n6993), .ZN(n9389) );
  AND2_X1 U6344 ( .A1(n5553), .A2(n5531), .ZN(n5551) );
  AND2_X1 U6345 ( .A1(n5443), .A2(n5424), .ZN(n5441) );
  INV_X1 U6346 ( .A(n8469), .ZN(n9810) );
  OR2_X1 U6347 ( .A1(n8170), .A2(n8617), .ZN(n8304) );
  AND2_X1 U6348 ( .A1(n6166), .A2(n6165), .ZN(n8255) );
  AND4_X1 U6349 ( .A1(n6065), .A2(n6064), .A3(n6063), .A4(n6062), .ZN(n8618)
         );
  AND2_X1 U6350 ( .A1(n6559), .A2(n6558), .ZN(n9790) );
  INV_X1 U6351 ( .A(n9792), .ZN(n9791) );
  INV_X1 U6352 ( .A(n8210), .ZN(n8204) );
  INV_X1 U6353 ( .A(n8503), .ZN(n8498) );
  INV_X1 U6354 ( .A(n8617), .ZN(n8590) );
  INV_X1 U6355 ( .A(n8475), .ZN(n8632) );
  NAND2_X1 U6356 ( .A1(n6811), .A2(n9841), .ZN(n7026) );
  AND2_X1 U6357 ( .A1(n9805), .A2(n9883), .ZN(n8720) );
  INV_X1 U6358 ( .A(n8720), .ZN(n9904) );
  NAND2_X1 U6359 ( .A1(n6869), .A2(n6415), .ZN(n9819) );
  NAND2_X1 U6360 ( .A1(n5857), .A2(n5833), .ZN(n5831) );
  NAND2_X1 U6361 ( .A1(n5725), .A2(n5724), .ZN(n9282) );
  NAND4_X1 U6362 ( .A1(n7046), .A2(n7045), .A3(n7044), .A4(n7043), .ZN(n6719)
         );
  INV_X1 U6363 ( .A(n9745), .ZN(n9714) );
  INV_X1 U6364 ( .A(n9228), .ZN(n9103) );
  AND2_X1 U6365 ( .A1(n9035), .A2(n9036), .ZN(n9352) );
  AND2_X1 U6366 ( .A1(n8963), .A2(n8888), .ZN(n9098) );
  OR2_X1 U6367 ( .A1(n7447), .A2(n7591), .ZN(n9086) );
  OR2_X1 U6368 ( .A1(n7072), .A2(n9148), .ZN(n9776) );
  AND2_X1 U6369 ( .A1(n9340), .A2(n9339), .ZN(n9484) );
  INV_X1 U6370 ( .A(n9771), .ZN(n9526) );
  NAND2_X1 U6371 ( .A1(n7815), .A2(n9571), .ZN(n9771) );
  OR2_X1 U6372 ( .A1(n7041), .A2(n7040), .ZN(n7064) );
  INV_X1 U6373 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10190) );
  INV_X1 U6374 ( .A(n8388), .ZN(n9797) );
  OR2_X1 U6375 ( .A1(n8170), .A2(n8615), .ZN(n8302) );
  OR2_X1 U6376 ( .A1(n6418), .A2(n6417), .ZN(n6419) );
  INV_X1 U6377 ( .A(n8254), .ZN(n8492) );
  INV_X1 U6378 ( .A(n9790), .ZN(n9795) );
  NAND2_X1 U6379 ( .A1(n6841), .A2(n8469), .ZN(n9817) );
  NOR2_X1 U6380 ( .A1(n7027), .A2(n7026), .ZN(n9922) );
  INV_X1 U6381 ( .A(n9908), .ZN(n9906) );
  NOR2_X1 U6382 ( .A1(n9820), .A2(n9819), .ZN(n9831) );
  CLKBUF_X1 U6383 ( .A(n9831), .Z(n9845) );
  INV_X1 U6384 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7651) );
  INV_X1 U6385 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6957) );
  INV_X1 U6386 ( .A(n9486), .ZN(n9350) );
  INV_X1 U6387 ( .A(n8850), .ZN(n8874) );
  NAND2_X1 U6388 ( .A1(n5746), .A2(n5745), .ZN(n9157) );
  NAND2_X1 U6389 ( .A1(n5625), .A2(n5624), .ZN(n9354) );
  OR2_X1 U6390 ( .A1(P1_U3083), .A2(n6690), .ZN(n9754) );
  AOI21_X1 U6391 ( .B1(n9261), .B2(n9433), .A(n9260), .ZN(n9458) );
  NAND2_X1 U6392 ( .A1(n9379), .A2(n7162), .ZN(n9444) );
  INV_X1 U6393 ( .A(n7442), .ZN(n7822) );
  INV_X1 U6394 ( .A(n9787), .ZN(n9528) );
  INV_X1 U6395 ( .A(n9782), .ZN(n9783) );
  INV_X1 U6396 ( .A(n9772), .ZN(n9782) );
  INV_X1 U6397 ( .A(n9758), .ZN(n9757) );
  AND2_X1 U6398 ( .A1(n9756), .A2(n9755), .ZN(n9758) );
  INV_X1 U6399 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10223) );
  INV_X1 U6400 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10230) );
  INV_X1 U6401 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10131) );
  INV_X1 U6402 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10194) );
  INV_X1 U6403 ( .A(n9548), .ZN(n8222) );
  NAND2_X1 U6404 ( .A1(n6429), .A2(n6428), .ZN(P1_U3238) );
  INV_X2 U6405 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NAND2_X1 U6406 ( .A1(n5044), .A2(n4942), .ZN(n5093) );
  INV_X1 U6407 ( .A(n5093), .ZN(n4943) );
  NAND2_X1 U6408 ( .A1(n4390), .A2(n4943), .ZN(n5227) );
  NOR2_X1 U6409 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n4948) );
  NOR2_X1 U6410 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4947) );
  NAND4_X1 U6411 ( .A1(n4948), .A2(n4947), .A3(n4946), .A4(n4974), .ZN(n4950)
         );
  NAND4_X1 U6412 ( .A1(n4972), .A2(n5365), .A3(n5450), .A4(n5004), .ZN(n4949)
         );
  NOR2_X1 U6413 ( .A1(n4950), .A2(n4949), .ZN(n4951) );
  XNOR2_X2 U6414 ( .A(n4956), .B(n4955), .ZN(n8220) );
  NAND2_X4 U6415 ( .A1(n4961), .A2(n8047), .ZN(n5142) );
  INV_X1 U6416 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n4960) );
  OR2_X1 U6417 ( .A1(n5142), .A2(n4960), .ZN(n4967) );
  NAND2_X1 U6418 ( .A1(n5058), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4965) );
  INV_X1 U6420 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n4963) );
  OR2_X1 U6421 ( .A1(n5057), .A2(n4963), .ZN(n4964) );
  NAND4_X2 U6422 ( .A1(n4967), .A2(n4966), .A3(n4965), .A4(n4964), .ZN(n6680)
         );
  NOR2_X1 U6423 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n4968) );
  AND2_X1 U6424 ( .A1(n4968), .A2(n5447), .ZN(n4969) );
  NAND2_X1 U6425 ( .A1(n4973), .A2(n5006), .ZN(n5010) );
  XNOR2_X2 U6426 ( .A(n4978), .B(n4977), .ZN(n7489) );
  INV_X1 U6427 ( .A(n4981), .ZN(n4982) );
  NAND2_X1 U6428 ( .A1(n4982), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4983) );
  NAND2_X1 U6429 ( .A1(n4984), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4986) );
  NOR2_X1 U6430 ( .A1(n7944), .A2(n7839), .ZN(n4989) );
  NAND2_X1 U6431 ( .A1(n4989), .A2(n5770), .ZN(n5000) );
  NAND2_X1 U6432 ( .A1(n6680), .A2(n5699), .ZN(n5002) );
  INV_X1 U6433 ( .A(n4993), .ZN(n4995) );
  NAND2_X1 U6434 ( .A1(n5634), .A2(SI_0_), .ZN(n4997) );
  XNOR2_X1 U6435 ( .A(n4997), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9552) );
  INV_X1 U6436 ( .A(n6430), .ZN(n5013) );
  AOI22_X1 U6437 ( .A1(n7348), .A2(n5028), .B1(P1_REG1_REG_0__SCAN_IN), .B2(
        n5013), .ZN(n5001) );
  NAND2_X1 U6438 ( .A1(n5006), .A2(n5007), .ZN(n5008) );
  NAND2_X1 U6439 ( .A1(n5008), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5009) );
  MUX2_X1 U6440 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5009), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n5011) );
  NAND2_X1 U6441 ( .A1(n5778), .A2(n9317), .ZN(n9072) );
  NAND2_X1 U6442 ( .A1(n5012), .A2(n5049), .ZN(n5017) );
  NAND2_X1 U6443 ( .A1(n5776), .A2(n5787), .ZN(n7346) );
  NAND2_X1 U6444 ( .A1(n6680), .A2(n5747), .ZN(n5016) );
  INV_X1 U6445 ( .A(n5630), .ZN(n5699) );
  AOI21_X1 U6446 ( .B1(n5699), .B2(n7348), .A(n5014), .ZN(n5015) );
  AND2_X1 U6447 ( .A1(n5016), .A2(n5015), .ZN(n6637) );
  AND2_X1 U6448 ( .A1(n5017), .A2(n6638), .ZN(n5032) );
  INV_X1 U6449 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7002) );
  OR2_X1 U6450 ( .A1(n5142), .A2(n7002), .ZN(n5022) );
  NAND2_X1 U6451 ( .A1(n5098), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5021) );
  INV_X1 U6452 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5018) );
  OR2_X1 U6453 ( .A1(n5057), .A2(n5018), .ZN(n5020) );
  NAND2_X1 U6454 ( .A1(n5058), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5019) );
  NAND2_X1 U6455 ( .A1(n6974), .A2(n5699), .ZN(n5030) );
  AND2_X1 U6456 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5023) );
  NAND2_X1 U6457 ( .A1(n5091), .A2(n5023), .ZN(n5872) );
  NAND3_X1 U6458 ( .A1(n4380), .A2(SI_0_), .A3(P2_DATAO_REG_0__SCAN_IN), .ZN(
        n5024) );
  NAND2_X1 U6459 ( .A1(n5872), .A2(n5024), .ZN(n5040) );
  INV_X1 U6460 ( .A(SI_1_), .ZN(n10210) );
  XNOR2_X1 U6461 ( .A(n5040), .B(n10210), .ZN(n5039) );
  MUX2_X1 U6462 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4380), .Z(n5038) );
  XNOR2_X1 U6463 ( .A(n5039), .B(n5038), .ZN(n6467) );
  NAND2_X1 U6464 ( .A1(n5092), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5027) );
  NAND2_X1 U6465 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5025) );
  XNOR2_X1 U6466 ( .A(n5025), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6463) );
  NAND2_X1 U6467 ( .A1(n6718), .A2(n5753), .ZN(n5029) );
  NAND2_X1 U6468 ( .A1(n5030), .A2(n5029), .ZN(n5031) );
  XNOR2_X1 U6469 ( .A(n5031), .B(n5049), .ZN(n5033) );
  INV_X2 U6470 ( .A(n5630), .ZN(n5752) );
  NAND2_X1 U6471 ( .A1(n6714), .A2(n6717), .ZN(n5036) );
  INV_X1 U6472 ( .A(n5032), .ZN(n5035) );
  INV_X1 U6473 ( .A(n5033), .ZN(n5034) );
  NAND2_X1 U6474 ( .A1(n5035), .A2(n5034), .ZN(n6715) );
  NAND2_X1 U6475 ( .A1(n5036), .A2(n6715), .ZN(n6706) );
  NAND2_X1 U6476 ( .A1(n5098), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n7046) );
  NAND2_X1 U6477 ( .A1(n5058), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7045) );
  INV_X1 U6478 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5037) );
  OR2_X1 U6479 ( .A1(n5057), .A2(n5037), .ZN(n7044) );
  INV_X1 U6480 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9961) );
  NAND2_X1 U6481 ( .A1(n6719), .A2(n5699), .ZN(n5048) );
  NAND2_X1 U6482 ( .A1(n5039), .A2(n5038), .ZN(n5042) );
  NAND2_X1 U6483 ( .A1(n5040), .A2(SI_1_), .ZN(n5041) );
  INV_X1 U6484 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6477) );
  INV_X1 U6485 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n5043) );
  MUX2_X1 U6486 ( .A(n6477), .B(n5043), .S(n6466), .Z(n5065) );
  XNOR2_X1 U6487 ( .A(n5064), .B(n5063), .ZN(n6476) );
  INV_X1 U6488 ( .A(n6692), .ZN(n5045) );
  NAND2_X1 U6489 ( .A1(n6708), .A2(n5753), .ZN(n5047) );
  NAND2_X1 U6490 ( .A1(n5048), .A2(n5047), .ZN(n5050) );
  INV_X4 U6491 ( .A(n5049), .ZN(n5750) );
  XNOR2_X1 U6492 ( .A(n5050), .B(n5750), .ZN(n5054) );
  INV_X1 U6493 ( .A(n5054), .ZN(n5052) );
  AOI22_X1 U6494 ( .A1(n6719), .A2(n5747), .B1(n5752), .B2(n6708), .ZN(n5053)
         );
  NAND2_X1 U6495 ( .A1(n5052), .A2(n5051), .ZN(n5055) );
  NAND2_X1 U6496 ( .A1(n5054), .A2(n5053), .ZN(n5056) );
  NAND2_X1 U6497 ( .A1(n6706), .A2(n6707), .ZN(n6705) );
  OR2_X1 U6498 ( .A1(n5692), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5062) );
  NAND2_X1 U6499 ( .A1(n5791), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5061) );
  NAND2_X1 U6500 ( .A1(n5058), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5060) );
  INV_X1 U6501 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7374) );
  OR2_X1 U6502 ( .A1(n5142), .A2(n7374), .ZN(n5059) );
  NAND4_X2 U6503 ( .A1(n5062), .A2(n5061), .A3(n5060), .A4(n5059), .ZN(n7157)
         );
  NAND2_X1 U6504 ( .A1(n7157), .A2(n5752), .ZN(n5077) );
  INV_X1 U6505 ( .A(n5065), .ZN(n5066) );
  NAND2_X1 U6506 ( .A1(n5066), .A2(SI_2_), .ZN(n5084) );
  NAND2_X1 U6507 ( .A1(n5086), .A2(n5084), .ZN(n5068) );
  INV_X1 U6508 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6484) );
  INV_X1 U6509 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5067) );
  XNOR2_X1 U6510 ( .A(n5068), .B(n5088), .ZN(n8049) );
  NAND2_X1 U6511 ( .A1(n5092), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5075) );
  INV_X1 U6512 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5070) );
  NAND2_X1 U6513 ( .A1(n5071), .A2(n5070), .ZN(n5072) );
  NAND2_X1 U6514 ( .A1(n5072), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5073) );
  NAND2_X1 U6515 ( .A1(n5507), .A2(n8061), .ZN(n5074) );
  NAND2_X1 U6516 ( .A1(n7380), .A2(n5753), .ZN(n5076) );
  NAND2_X1 U6517 ( .A1(n5077), .A2(n5076), .ZN(n5078) );
  XNOR2_X1 U6518 ( .A(n5078), .B(n5049), .ZN(n5079) );
  AOI22_X1 U6519 ( .A1(n7157), .A2(n5747), .B1(n5752), .B2(n7380), .ZN(n5080)
         );
  NAND2_X1 U6520 ( .A1(n6760), .A2(n6758), .ZN(n6759) );
  INV_X1 U6521 ( .A(n5079), .ZN(n5081) );
  NAND2_X1 U6522 ( .A1(n5081), .A2(n5080), .ZN(n5082) );
  NAND2_X1 U6523 ( .A1(n6759), .A2(n5082), .ZN(n6768) );
  NAND2_X1 U6524 ( .A1(n5083), .A2(SI_3_), .ZN(n5087) );
  INV_X1 U6525 ( .A(n5087), .ZN(n5089) );
  MUX2_X1 U6526 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n4380), .Z(n5123) );
  INV_X1 U6527 ( .A(SI_4_), .ZN(n10209) );
  XNOR2_X1 U6528 ( .A(n5123), .B(n10209), .ZN(n5121) );
  XNOR2_X1 U6529 ( .A(n5122), .B(n5121), .ZN(n6482) );
  CLKBUF_X3 U6530 ( .A(n5092), .Z(n5614) );
  NAND2_X1 U6531 ( .A1(n5614), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5097) );
  NAND2_X1 U6532 ( .A1(n5093), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5094) );
  MUX2_X1 U6533 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5094), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5095) );
  AND2_X1 U6534 ( .A1(n5095), .A2(n5147), .ZN(n9603) );
  NAND2_X1 U6535 ( .A1(n5507), .A2(n9603), .ZN(n5096) );
  OAI211_X1 U6536 ( .C1(n5155), .C2(n6482), .A(n5097), .B(n5096), .ZN(n7246)
         );
  NAND2_X1 U6537 ( .A1(n7246), .A2(n5753), .ZN(n5106) );
  NAND2_X1 U6538 ( .A1(n5058), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5104) );
  INV_X1 U6539 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5099) );
  XNOR2_X1 U6540 ( .A(n5099), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n6773) );
  NAND2_X1 U6541 ( .A1(n5098), .A2(n6773), .ZN(n5103) );
  INV_X1 U6542 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5100) );
  OR2_X1 U6543 ( .A1(n5057), .A2(n5100), .ZN(n5102) );
  INV_X1 U6544 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7438) );
  OR2_X1 U6545 ( .A1(n5142), .A2(n7438), .ZN(n5101) );
  NAND4_X1 U6546 ( .A1(n5104), .A2(n5103), .A3(n5102), .A4(n5101), .ZN(n9170)
         );
  NAND2_X1 U6547 ( .A1(n9170), .A2(n5752), .ZN(n5105) );
  NAND2_X1 U6548 ( .A1(n5106), .A2(n5105), .ZN(n5107) );
  AOI22_X1 U6549 ( .A1(n9170), .A2(n5747), .B1(n5752), .B2(n7246), .ZN(n5109)
         );
  XNOR2_X1 U6550 ( .A(n5108), .B(n5109), .ZN(n6769) );
  INV_X1 U6551 ( .A(n5108), .ZN(n5111) );
  INV_X1 U6552 ( .A(n5109), .ZN(n5110) );
  NAND2_X1 U6553 ( .A1(n5111), .A2(n5110), .ZN(n5134) );
  NAND2_X1 U6554 ( .A1(n5058), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5120) );
  NAND3_X1 U6555 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5140) );
  INV_X1 U6556 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5113) );
  NAND2_X1 U6557 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5112) );
  NAND2_X1 U6558 ( .A1(n5113), .A2(n5112), .ZN(n5114) );
  AND2_X1 U6559 ( .A1(n5140), .A2(n5114), .ZN(n7105) );
  NAND2_X1 U6560 ( .A1(n5098), .A2(n7105), .ZN(n5119) );
  INV_X1 U6561 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5115) );
  OR2_X1 U6562 ( .A1(n5057), .A2(n5115), .ZN(n5118) );
  INV_X1 U6563 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5116) );
  OR2_X1 U6564 ( .A1(n5142), .A2(n5116), .ZN(n5117) );
  NAND4_X1 U6565 ( .A1(n5120), .A2(n5119), .A3(n5118), .A4(n5117), .ZN(n9169)
         );
  NAND2_X1 U6566 ( .A1(n9169), .A2(n5699), .ZN(n5131) );
  NAND2_X1 U6567 ( .A1(n5122), .A2(n5121), .ZN(n5125) );
  NAND2_X1 U6568 ( .A1(n5123), .A2(SI_4_), .ZN(n5124) );
  NAND2_X1 U6569 ( .A1(n5125), .A2(n5124), .ZN(n5150) );
  INV_X1 U6570 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6479) );
  INV_X1 U6571 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n5126) );
  MUX2_X1 U6572 ( .A(n6479), .B(n5126), .S(n4380), .Z(n5151) );
  XNOR2_X1 U6573 ( .A(n5151), .B(SI_5_), .ZN(n5149) );
  XNOR2_X1 U6574 ( .A(n5150), .B(n5149), .ZN(n6478) );
  NAND2_X1 U6575 ( .A1(n5614), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5129) );
  NAND2_X1 U6576 ( .A1(n5147), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5127) );
  XNOR2_X1 U6577 ( .A(n5127), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9618) );
  NAND2_X1 U6578 ( .A1(n5507), .A2(n9618), .ZN(n5128) );
  NAND2_X1 U6579 ( .A1(n4379), .A2(n5753), .ZN(n5130) );
  NAND2_X1 U6580 ( .A1(n5131), .A2(n5130), .ZN(n5132) );
  INV_X1 U6581 ( .A(n5133), .ZN(n5135) );
  AND2_X1 U6582 ( .A1(n5135), .A2(n5134), .ZN(n5136) );
  NAND2_X1 U6583 ( .A1(n6770), .A2(n5136), .ZN(n5138) );
  AOI22_X1 U6584 ( .A1(n9169), .A2(n5747), .B1(n5699), .B2(n4379), .ZN(n7101)
         );
  INV_X1 U6585 ( .A(n5140), .ZN(n5139) );
  INV_X1 U6586 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n10071) );
  NAND2_X1 U6587 ( .A1(n5140), .A2(n10071), .ZN(n5141) );
  NAND2_X1 U6588 ( .A1(n5167), .A2(n5141), .ZN(n7320) );
  NAND2_X1 U6589 ( .A1(n5058), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5146) );
  NAND2_X1 U6590 ( .A1(n5792), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5145) );
  INV_X1 U6591 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5143) );
  OR2_X1 U6592 ( .A1(n5057), .A2(n5143), .ZN(n5144) );
  NAND2_X1 U6593 ( .A1(n9168), .A2(n5752), .ZN(n5159) );
  NOR2_X1 U6594 ( .A1(n5147), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5180) );
  OR2_X1 U6595 ( .A1(n5180), .A2(n9546), .ZN(n5148) );
  INV_X1 U6596 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5179) );
  XNOR2_X1 U6597 ( .A(n5148), .B(n5179), .ZN(n9635) );
  NAND2_X1 U6598 ( .A1(n5150), .A2(n5149), .ZN(n5154) );
  INV_X1 U6599 ( .A(n5151), .ZN(n5152) );
  NAND2_X1 U6600 ( .A1(n5152), .A2(SI_5_), .ZN(n5153) );
  MUX2_X1 U6601 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n4380), .Z(n5177) );
  XNOR2_X1 U6602 ( .A(n5177), .B(SI_6_), .ZN(n5174) );
  XNOR2_X1 U6603 ( .A(n5176), .B(n5174), .ZN(n6474) );
  NAND2_X1 U6604 ( .A1(n6474), .A2(n8882), .ZN(n5157) );
  NAND2_X1 U6605 ( .A1(n5614), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n5156) );
  OAI211_X1 U6606 ( .C1(n5069), .C2(n9635), .A(n5157), .B(n5156), .ZN(n7211)
         );
  NAND2_X1 U6607 ( .A1(n4383), .A2(n5753), .ZN(n5158) );
  NAND2_X1 U6608 ( .A1(n5159), .A2(n5158), .ZN(n5160) );
  XNOR2_X1 U6609 ( .A(n5160), .B(n5750), .ZN(n5161) );
  AOI22_X1 U6610 ( .A1(n9168), .A2(n5747), .B1(n5699), .B2(n4383), .ZN(n5162)
         );
  INV_X1 U6611 ( .A(n5161), .ZN(n5164) );
  INV_X1 U6612 ( .A(n5162), .ZN(n5163) );
  NAND2_X1 U6613 ( .A1(n5164), .A2(n5163), .ZN(n7145) );
  INV_X1 U6614 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U6615 ( .A1(n5167), .A2(n5166), .ZN(n5168) );
  NAND2_X1 U6616 ( .A1(n5207), .A2(n5168), .ZN(n7291) );
  OR2_X1 U6617 ( .A1(n5692), .A2(n7291), .ZN(n5173) );
  NAND2_X1 U6618 ( .A1(n5534), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5172) );
  NAND2_X1 U6619 ( .A1(n5791), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5171) );
  INV_X1 U6620 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n5169) );
  OR2_X1 U6621 ( .A1(n5142), .A2(n5169), .ZN(n5170) );
  NAND4_X1 U6622 ( .A1(n5173), .A2(n5172), .A3(n5171), .A4(n5170), .ZN(n9167)
         );
  NAND2_X1 U6623 ( .A1(n9167), .A2(n5752), .ZN(n5185) );
  INV_X1 U6624 ( .A(n5174), .ZN(n5175) );
  NAND2_X1 U6625 ( .A1(n5177), .A2(SI_6_), .ZN(n5178) );
  MUX2_X1 U6626 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4380), .Z(n5197) );
  XNOR2_X1 U6627 ( .A(n5197), .B(SI_7_), .ZN(n5194) );
  XNOR2_X1 U6628 ( .A(n5196), .B(n5194), .ZN(n6485) );
  NAND2_X1 U6629 ( .A1(n6485), .A2(n8882), .ZN(n5183) );
  NAND2_X1 U6630 ( .A1(n5180), .A2(n5179), .ZN(n5202) );
  NAND2_X1 U6631 ( .A1(n5202), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5181) );
  XNOR2_X1 U6632 ( .A(n5181), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6501) );
  AOI22_X1 U6633 ( .A1(n5614), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5507), .B2(
        n6501), .ZN(n5182) );
  NAND2_X1 U6634 ( .A1(n5183), .A2(n5182), .ZN(n7485) );
  NAND2_X1 U6635 ( .A1(n7485), .A2(n5753), .ZN(n5184) );
  NAND2_X1 U6636 ( .A1(n5185), .A2(n5184), .ZN(n5186) );
  XNOR2_X1 U6637 ( .A(n5186), .B(n5049), .ZN(n5189) );
  NAND2_X1 U6638 ( .A1(n9167), .A2(n5747), .ZN(n5188) );
  NAND2_X1 U6639 ( .A1(n7485), .A2(n5752), .ZN(n5187) );
  NAND2_X1 U6640 ( .A1(n5188), .A2(n5187), .ZN(n5190) );
  XNOR2_X1 U6641 ( .A(n5189), .B(n5190), .ZN(n7479) );
  INV_X1 U6642 ( .A(n5189), .ZN(n5192) );
  INV_X1 U6643 ( .A(n5190), .ZN(n5191) );
  NAND2_X1 U6644 ( .A1(n5192), .A2(n5191), .ZN(n5193) );
  INV_X1 U6645 ( .A(n5194), .ZN(n5195) );
  MUX2_X1 U6646 ( .A(n10193), .B(n6491), .S(n5634), .Z(n5199) );
  INV_X1 U6647 ( .A(SI_8_), .ZN(n5198) );
  NAND2_X1 U6648 ( .A1(n5199), .A2(n5198), .ZN(n5223) );
  INV_X1 U6649 ( .A(n5199), .ZN(n5200) );
  NAND2_X1 U6650 ( .A1(n5200), .A2(SI_8_), .ZN(n5201) );
  NAND2_X1 U6651 ( .A1(n5223), .A2(n5201), .ZN(n5221) );
  XNOR2_X1 U6652 ( .A(n5222), .B(n5221), .ZN(n6489) );
  NAND2_X1 U6653 ( .A1(n6489), .A2(n8882), .ZN(n5205) );
  OAI21_X1 U6654 ( .B1(n5202), .B2(P1_IR_REG_7__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5203) );
  XNOR2_X1 U6655 ( .A(n5203), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9650) );
  AOI22_X1 U6656 ( .A1(n5614), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5507), .B2(
        n9650), .ZN(n5204) );
  NAND2_X1 U6657 ( .A1(n5205), .A2(n5204), .ZN(n7702) );
  NAND2_X1 U6658 ( .A1(n5534), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5213) );
  INV_X1 U6659 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10219) );
  NAND2_X1 U6660 ( .A1(n5207), .A2(n10219), .ZN(n5208) );
  AND2_X1 U6661 ( .A1(n5235), .A2(n5208), .ZN(n7691) );
  NAND2_X1 U6662 ( .A1(n5098), .A2(n7691), .ZN(n5212) );
  INV_X1 U6663 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5209) );
  OR2_X1 U6664 ( .A1(n5057), .A2(n5209), .ZN(n5211) );
  INV_X1 U6665 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7415) );
  OR2_X1 U6666 ( .A1(n5142), .A2(n7415), .ZN(n5210) );
  NAND4_X1 U6667 ( .A1(n5213), .A2(n5212), .A3(n5211), .A4(n5210), .ZN(n9166)
         );
  AOI22_X1 U6668 ( .A1(n7702), .A2(n5752), .B1(n5747), .B2(n9166), .ZN(n5218)
         );
  NAND2_X1 U6669 ( .A1(n7702), .A2(n5753), .ZN(n5216) );
  NAND2_X1 U6670 ( .A1(n9166), .A2(n5699), .ZN(n5215) );
  NAND2_X1 U6671 ( .A1(n5216), .A2(n5215), .ZN(n5217) );
  XNOR2_X1 U6672 ( .A(n5217), .B(n5750), .ZN(n7697) );
  NAND2_X1 U6673 ( .A1(n7695), .A2(n7697), .ZN(n5220) );
  NAND2_X1 U6674 ( .A1(n5219), .A2(n5218), .ZN(n7696) );
  NAND2_X1 U6675 ( .A1(n5220), .A2(n7696), .ZN(n7779) );
  MUX2_X1 U6676 ( .A(n6509), .B(n6507), .S(n4380), .Z(n5224) );
  NAND2_X1 U6677 ( .A1(n5224), .A2(n10074), .ZN(n5280) );
  INV_X1 U6678 ( .A(n5224), .ZN(n5225) );
  NAND2_X1 U6679 ( .A1(n5225), .A2(SI_9_), .ZN(n5226) );
  XNOR2_X1 U6680 ( .A(n5251), .B(n5277), .ZN(n6505) );
  NAND2_X1 U6681 ( .A1(n6505), .A2(n8882), .ZN(n5233) );
  NAND2_X1 U6682 ( .A1(n5227), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5228) );
  MUX2_X1 U6683 ( .A(n5228), .B(P1_IR_REG_31__SCAN_IN), .S(n5229), .Z(n5231)
         );
  INV_X1 U6684 ( .A(n5227), .ZN(n5230) );
  NAND2_X1 U6685 ( .A1(n5230), .A2(n5229), .ZN(n5259) );
  NAND2_X1 U6686 ( .A1(n5231), .A2(n5259), .ZN(n6506) );
  AOI22_X1 U6687 ( .A1(n5614), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5507), .B2(
        n6731), .ZN(n5232) );
  NAND2_X1 U6688 ( .A1(n5233), .A2(n5232), .ZN(n7784) );
  NAND2_X1 U6689 ( .A1(n7784), .A2(n5753), .ZN(n5243) );
  NAND2_X1 U6690 ( .A1(n5235), .A2(n5234), .ZN(n5236) );
  NAND2_X1 U6691 ( .A1(n5265), .A2(n5236), .ZN(n7774) );
  OR2_X1 U6692 ( .A1(n5692), .A2(n7774), .ZN(n5241) );
  NAND2_X1 U6693 ( .A1(n5534), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5240) );
  INV_X1 U6694 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n5237) );
  OR2_X1 U6695 ( .A1(n5057), .A2(n5237), .ZN(n5239) );
  INV_X1 U6696 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7452) );
  OR2_X1 U6697 ( .A1(n5142), .A2(n7452), .ZN(n5238) );
  NAND4_X1 U6698 ( .A1(n5241), .A2(n5240), .A3(n5239), .A4(n5238), .ZN(n9165)
         );
  NAND2_X1 U6699 ( .A1(n9165), .A2(n5752), .ZN(n5242) );
  NAND2_X1 U6700 ( .A1(n5243), .A2(n5242), .ZN(n5244) );
  XNOR2_X1 U6701 ( .A(n5244), .B(n5049), .ZN(n5246) );
  AND2_X1 U6702 ( .A1(n9165), .A2(n5747), .ZN(n5245) );
  AOI21_X1 U6703 ( .B1(n7784), .B2(n5752), .A(n5245), .ZN(n5247) );
  NAND2_X1 U6704 ( .A1(n7779), .A2(n7780), .ZN(n5250) );
  INV_X1 U6705 ( .A(n5246), .ZN(n5248) );
  NAND2_X1 U6706 ( .A1(n5248), .A2(n5247), .ZN(n5249) );
  NAND2_X1 U6707 ( .A1(n5251), .A2(n5277), .ZN(n5252) );
  NAND2_X1 U6708 ( .A1(n5252), .A2(n5280), .ZN(n5257) );
  MUX2_X1 U6709 ( .A(n6537), .B(n6536), .S(n4380), .Z(n5254) );
  INV_X1 U6710 ( .A(SI_10_), .ZN(n5253) );
  NAND2_X1 U6711 ( .A1(n5254), .A2(n5253), .ZN(n5279) );
  INV_X1 U6712 ( .A(n5254), .ZN(n5255) );
  NAND2_X1 U6713 ( .A1(n5255), .A2(SI_10_), .ZN(n5278) );
  AND2_X1 U6714 ( .A1(n5279), .A2(n5278), .ZN(n5256) );
  XNOR2_X1 U6715 ( .A(n5257), .B(n5256), .ZN(n6535) );
  NAND2_X1 U6716 ( .A1(n6535), .A2(n8882), .ZN(n5264) );
  NAND2_X1 U6717 ( .A1(n5259), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5258) );
  MUX2_X1 U6718 ( .A(n5258), .B(P1_IR_REG_31__SCAN_IN), .S(n5260), .Z(n5262)
         );
  INV_X1 U6719 ( .A(n5259), .ZN(n5261) );
  NAND2_X1 U6720 ( .A1(n5261), .A2(n5260), .ZN(n5285) );
  NAND2_X1 U6721 ( .A1(n5262), .A2(n5285), .ZN(n6794) );
  INV_X1 U6722 ( .A(n6794), .ZN(n6799) );
  AOI22_X1 U6723 ( .A1(n5614), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5507), .B2(
        n6799), .ZN(n5263) );
  NAND2_X1 U6724 ( .A1(n7664), .A2(n5753), .ZN(n5272) );
  NAND2_X1 U6725 ( .A1(n5265), .A2(n9986), .ZN(n5266) );
  NAND2_X1 U6726 ( .A1(n5291), .A2(n5266), .ZN(n7662) );
  OR2_X1 U6727 ( .A1(n5692), .A2(n7662), .ZN(n5270) );
  NAND2_X1 U6728 ( .A1(n5791), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5269) );
  NAND2_X1 U6729 ( .A1(n5534), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5268) );
  INV_X1 U6730 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7339) );
  OR2_X1 U6731 ( .A1(n5142), .A2(n7339), .ZN(n5267) );
  NAND4_X1 U6732 ( .A1(n5270), .A2(n5269), .A3(n5268), .A4(n5267), .ZN(n9164)
         );
  NAND2_X1 U6733 ( .A1(n9164), .A2(n5752), .ZN(n5271) );
  NAND2_X1 U6734 ( .A1(n5272), .A2(n5271), .ZN(n5273) );
  XNOR2_X1 U6735 ( .A(n5273), .B(n5750), .ZN(n7655) );
  AND2_X1 U6736 ( .A1(n9164), .A2(n5747), .ZN(n5274) );
  AOI21_X1 U6737 ( .B1(n7664), .B2(n5752), .A(n5274), .ZN(n7654) );
  AND2_X1 U6738 ( .A1(n7655), .A2(n7654), .ZN(n5276) );
  OR2_X1 U6739 ( .A1(n7655), .A2(n7654), .ZN(n5275) );
  INV_X1 U6740 ( .A(n5278), .ZN(n5282) );
  MUX2_X1 U6741 ( .A(n6540), .B(n6542), .S(n5634), .Z(n5307) );
  XNOR2_X1 U6742 ( .A(n5307), .B(SI_11_), .ZN(n5306) );
  XNOR2_X1 U6743 ( .A(n5309), .B(n5306), .ZN(n6539) );
  NAND2_X1 U6744 ( .A1(n6539), .A2(n8882), .ZN(n5288) );
  NAND2_X1 U6745 ( .A1(n5285), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5284) );
  MUX2_X1 U6746 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5284), .S(
        P1_IR_REG_11__SCAN_IN), .Z(n5286) );
  AOI22_X1 U6747 ( .A1(n5614), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5507), .B2(
        n9185), .ZN(n5287) );
  NAND2_X1 U6748 ( .A1(n7794), .A2(n5753), .ZN(n5298) );
  INV_X1 U6749 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5290) );
  NAND2_X1 U6750 ( .A1(n5291), .A2(n5290), .ZN(n5292) );
  NAND2_X1 U6751 ( .A1(n5321), .A2(n5292), .ZN(n7792) );
  OR2_X1 U6752 ( .A1(n5692), .A2(n7792), .ZN(n5296) );
  NAND2_X1 U6753 ( .A1(n5534), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5295) );
  NAND2_X1 U6754 ( .A1(n5791), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5294) );
  INV_X1 U6755 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7598) );
  OR2_X1 U6756 ( .A1(n5142), .A2(n7598), .ZN(n5293) );
  NAND4_X1 U6757 ( .A1(n5296), .A2(n5295), .A3(n5294), .A4(n5293), .ZN(n9163)
         );
  NAND2_X1 U6758 ( .A1(n9163), .A2(n5752), .ZN(n5297) );
  NAND2_X1 U6759 ( .A1(n5298), .A2(n5297), .ZN(n5299) );
  XNOR2_X1 U6760 ( .A(n5299), .B(n5049), .ZN(n5303) );
  AND2_X1 U6761 ( .A1(n9163), .A2(n5747), .ZN(n5300) );
  AOI21_X1 U6762 ( .B1(n7794), .B2(n5752), .A(n5300), .ZN(n5301) );
  XNOR2_X1 U6763 ( .A(n5303), .B(n5301), .ZN(n7787) );
  NAND2_X1 U6764 ( .A1(n7786), .A2(n7787), .ZN(n5305) );
  INV_X1 U6765 ( .A(n5301), .ZN(n5302) );
  NAND2_X1 U6766 ( .A1(n5303), .A2(n5302), .ZN(n5304) );
  INV_X1 U6767 ( .A(n5307), .ZN(n5308) );
  MUX2_X1 U6768 ( .A(n6683), .B(n10194), .S(n5634), .Z(n5311) );
  INV_X1 U6769 ( .A(SI_12_), .ZN(n5310) );
  INV_X1 U6770 ( .A(n5311), .ZN(n5312) );
  NAND2_X1 U6771 ( .A1(n5312), .A2(SI_12_), .ZN(n5313) );
  NAND2_X1 U6772 ( .A1(n5337), .A2(n5313), .ZN(n5338) );
  XNOR2_X1 U6773 ( .A(n5339), .B(n5338), .ZN(n6682) );
  NAND2_X1 U6774 ( .A1(n6682), .A2(n8882), .ZN(n5319) );
  NAND2_X1 U6775 ( .A1(n5314), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5315) );
  MUX2_X1 U6776 ( .A(n5315), .B(P1_IR_REG_31__SCAN_IN), .S(n10225), .Z(n5317)
         );
  INV_X1 U6777 ( .A(n4971), .ZN(n5316) );
  NAND2_X1 U6778 ( .A1(n5317), .A2(n5316), .ZN(n9189) );
  INV_X1 U6779 ( .A(n9189), .ZN(n9661) );
  AOI22_X1 U6780 ( .A1(n5614), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5507), .B2(
        n9661), .ZN(n5318) );
  NAND2_X1 U6781 ( .A1(n7894), .A2(n5753), .ZN(n5328) );
  INV_X1 U6782 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7888) );
  NAND2_X1 U6783 ( .A1(n5321), .A2(n7888), .ZN(n5322) );
  NAND2_X1 U6784 ( .A1(n5348), .A2(n5322), .ZN(n7892) );
  OR2_X1 U6785 ( .A1(n5692), .A2(n7892), .ZN(n5326) );
  NAND2_X1 U6786 ( .A1(n5791), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5325) );
  NAND2_X1 U6787 ( .A1(n5534), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5324) );
  INV_X1 U6788 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7609) );
  OR2_X1 U6789 ( .A1(n5142), .A2(n7609), .ZN(n5323) );
  NAND4_X1 U6790 ( .A1(n5326), .A2(n5325), .A3(n5324), .A4(n5323), .ZN(n9162)
         );
  NAND2_X1 U6791 ( .A1(n9162), .A2(n5752), .ZN(n5327) );
  NAND2_X1 U6792 ( .A1(n5328), .A2(n5327), .ZN(n5329) );
  XNOR2_X1 U6793 ( .A(n5329), .B(n5750), .ZN(n5331) );
  AND2_X1 U6794 ( .A1(n9162), .A2(n5747), .ZN(n5330) );
  AOI21_X1 U6795 ( .B1(n7894), .B2(n5752), .A(n5330), .ZN(n5332) );
  NAND2_X1 U6796 ( .A1(n5331), .A2(n5332), .ZN(n5336) );
  INV_X1 U6797 ( .A(n5331), .ZN(n5334) );
  INV_X1 U6798 ( .A(n5332), .ZN(n5333) );
  NAND2_X1 U6799 ( .A1(n5334), .A2(n5333), .ZN(n5335) );
  NAND2_X1 U6800 ( .A1(n5336), .A2(n5335), .ZN(n7887) );
  MUX2_X1 U6801 ( .A(n6739), .B(n5340), .S(n5634), .Z(n5341) );
  INV_X1 U6802 ( .A(n5341), .ZN(n5342) );
  NAND2_X1 U6803 ( .A1(n5342), .A2(SI_13_), .ZN(n5343) );
  XNOR2_X1 U6804 ( .A(n5362), .B(n4933), .ZN(n6703) );
  NAND2_X1 U6805 ( .A1(n6703), .A2(n8882), .ZN(n5346) );
  OR2_X1 U6806 ( .A1(n4971), .A2(n9546), .ZN(n5344) );
  XNOR2_X1 U6807 ( .A(n5344), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9191) );
  AOI22_X1 U6808 ( .A1(n5614), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5507), .B2(
        n9191), .ZN(n5345) );
  NAND2_X1 U6809 ( .A1(n7906), .A2(n5753), .ZN(n5355) );
  NAND2_X1 U6810 ( .A1(n5348), .A2(n5347), .ZN(n5349) );
  NAND2_X1 U6811 ( .A1(n5371), .A2(n5349), .ZN(n7904) );
  OR2_X1 U6812 ( .A1(n5692), .A2(n7904), .ZN(n5353) );
  NAND2_X1 U6813 ( .A1(n5534), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5352) );
  NAND2_X1 U6814 ( .A1(n5791), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5351) );
  INV_X1 U6815 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9190) );
  OR2_X1 U6816 ( .A1(n5142), .A2(n9190), .ZN(n5350) );
  NAND4_X1 U6817 ( .A1(n5353), .A2(n5352), .A3(n5351), .A4(n5350), .ZN(n9161)
         );
  NAND2_X1 U6818 ( .A1(n9161), .A2(n5752), .ZN(n5354) );
  NAND2_X1 U6819 ( .A1(n5355), .A2(n5354), .ZN(n5356) );
  XNOR2_X1 U6820 ( .A(n5356), .B(n5750), .ZN(n5358) );
  AND2_X1 U6821 ( .A1(n9161), .A2(n5747), .ZN(n5357) );
  AOI21_X1 U6822 ( .B1(n7906), .B2(n5752), .A(n5357), .ZN(n5359) );
  AND2_X1 U6823 ( .A1(n5358), .A2(n5359), .ZN(n7898) );
  INV_X1 U6824 ( .A(n5358), .ZN(n5361) );
  INV_X1 U6825 ( .A(n5359), .ZN(n5360) );
  NAND2_X1 U6826 ( .A1(n5361), .A2(n5360), .ZN(n7899) );
  MUX2_X1 U6827 ( .A(n6742), .B(n10015), .S(n5634), .Z(n5382) );
  XNOR2_X1 U6828 ( .A(n5382), .B(SI_14_), .ZN(n5381) );
  XNOR2_X1 U6829 ( .A(n5386), .B(n5381), .ZN(n6740) );
  NAND2_X1 U6830 ( .A1(n6740), .A2(n8882), .ZN(n5369) );
  OR2_X1 U6831 ( .A1(n5006), .A2(n9546), .ZN(n5366) );
  NAND2_X1 U6832 ( .A1(n5366), .A2(n5365), .ZN(n5391) );
  OAI21_X1 U6833 ( .B1(n5366), .B2(n5365), .A(n5391), .ZN(n9690) );
  INV_X1 U6834 ( .A(n9690), .ZN(n5367) );
  AOI22_X1 U6835 ( .A1(n5614), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5507), .B2(
        n5367), .ZN(n5368) );
  NAND2_X1 U6836 ( .A1(n9524), .A2(n5753), .ZN(n5378) );
  INV_X1 U6837 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8029) );
  NAND2_X1 U6838 ( .A1(n5371), .A2(n8029), .ZN(n5372) );
  NAND2_X1 U6839 ( .A1(n5396), .A2(n5372), .ZN(n8033) );
  OR2_X1 U6840 ( .A1(n5692), .A2(n8033), .ZN(n5376) );
  NAND2_X1 U6841 ( .A1(n5534), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5375) );
  NAND2_X1 U6842 ( .A1(n5791), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5374) );
  INV_X1 U6843 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7801) );
  OR2_X1 U6844 ( .A1(n5142), .A2(n7801), .ZN(n5373) );
  NAND4_X1 U6845 ( .A1(n5376), .A2(n5375), .A3(n5374), .A4(n5373), .ZN(n9160)
         );
  NAND2_X1 U6846 ( .A1(n9160), .A2(n5752), .ZN(n5377) );
  NAND2_X1 U6847 ( .A1(n5378), .A2(n5377), .ZN(n5379) );
  XNOR2_X1 U6848 ( .A(n5379), .B(n5750), .ZN(n5407) );
  INV_X1 U6849 ( .A(n5407), .ZN(n5380) );
  INV_X1 U6850 ( .A(n5381), .ZN(n5385) );
  INV_X1 U6851 ( .A(n5382), .ZN(n5383) );
  NAND2_X1 U6852 ( .A1(n5383), .A2(SI_14_), .ZN(n5384) );
  MUX2_X1 U6853 ( .A(n6957), .B(n6955), .S(n5634), .Z(n5388) );
  INV_X1 U6854 ( .A(SI_15_), .ZN(n5387) );
  NAND2_X1 U6855 ( .A1(n5388), .A2(n5387), .ZN(n5418) );
  INV_X1 U6856 ( .A(n5388), .ZN(n5389) );
  NAND2_X1 U6857 ( .A1(n5389), .A2(SI_15_), .ZN(n5390) );
  NAND2_X1 U6858 ( .A1(n5418), .A2(n5390), .ZN(n5419) );
  XNOR2_X1 U6859 ( .A(n5420), .B(n5419), .ZN(n6954) );
  NAND2_X1 U6860 ( .A1(n6954), .A2(n8882), .ZN(n5394) );
  NAND2_X1 U6861 ( .A1(n5391), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5392) );
  XNOR2_X1 U6862 ( .A(n5392), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9704) );
  AOI22_X1 U6863 ( .A1(n5614), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5507), .B2(
        n9704), .ZN(n5393) );
  NAND2_X1 U6864 ( .A1(n8073), .A2(n5753), .ZN(n5404) );
  NAND2_X1 U6865 ( .A1(n5396), .A2(n5395), .ZN(n5397) );
  AND2_X1 U6866 ( .A1(n5430), .A2(n5397), .ZN(n8069) );
  NAND2_X1 U6867 ( .A1(n5098), .A2(n8069), .ZN(n5402) );
  NAND2_X1 U6868 ( .A1(n5534), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5401) );
  INV_X1 U6869 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n5398) );
  OR2_X1 U6870 ( .A1(n5057), .A2(n5398), .ZN(n5400) );
  OR2_X1 U6871 ( .A1(n5142), .A2(n9700), .ZN(n5399) );
  NAND4_X1 U6872 ( .A1(n5402), .A2(n5401), .A3(n5400), .A4(n5399), .ZN(n9159)
         );
  NAND2_X1 U6873 ( .A1(n9159), .A2(n5752), .ZN(n5403) );
  NAND2_X1 U6874 ( .A1(n5404), .A2(n5403), .ZN(n5405) );
  XNOR2_X1 U6875 ( .A(n5405), .B(n5750), .ZN(n5415) );
  AND2_X1 U6876 ( .A1(n8026), .A2(n5415), .ZN(n5411) );
  INV_X1 U6877 ( .A(n5406), .ZN(n5408) );
  NAND2_X1 U6878 ( .A1(n5408), .A2(n5407), .ZN(n8025) );
  NAND2_X1 U6879 ( .A1(n9524), .A2(n5752), .ZN(n5410) );
  NAND2_X1 U6880 ( .A1(n9160), .A2(n5747), .ZN(n5409) );
  NAND2_X1 U6881 ( .A1(n5410), .A2(n5409), .ZN(n8028) );
  NAND2_X1 U6882 ( .A1(n8025), .A2(n8028), .ZN(n5414) );
  NAND2_X1 U6883 ( .A1(n5411), .A2(n5414), .ZN(n8067) );
  NAND2_X1 U6884 ( .A1(n8073), .A2(n5752), .ZN(n5413) );
  NAND2_X1 U6885 ( .A1(n9159), .A2(n5747), .ZN(n5412) );
  NAND2_X1 U6886 ( .A1(n5413), .A2(n5412), .ZN(n8068) );
  NAND2_X1 U6887 ( .A1(n5414), .A2(n8026), .ZN(n5417) );
  INV_X1 U6888 ( .A(n5415), .ZN(n5416) );
  MUX2_X1 U6889 ( .A(n10188), .B(n10131), .S(n5634), .Z(n5422) );
  INV_X1 U6890 ( .A(SI_16_), .ZN(n5421) );
  INV_X1 U6891 ( .A(n5422), .ZN(n5423) );
  NAND2_X1 U6892 ( .A1(n5423), .A2(SI_16_), .ZN(n5424) );
  XNOR2_X1 U6893 ( .A(n5442), .B(n5441), .ZN(n7004) );
  NAND2_X1 U6894 ( .A1(n7004), .A2(n8882), .ZN(n5428) );
  NAND2_X1 U6895 ( .A1(n5006), .A2(n5446), .ZN(n5425) );
  NAND2_X1 U6896 ( .A1(n5425), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5426) );
  XNOR2_X1 U6897 ( .A(n5426), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9715) );
  AOI22_X1 U6898 ( .A1(n5614), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5507), .B2(
        n9715), .ZN(n5427) );
  NAND2_X1 U6899 ( .A1(n9519), .A2(n5753), .ZN(n5437) );
  INV_X1 U6900 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8802) );
  NAND2_X1 U6901 ( .A1(n5430), .A2(n8802), .ZN(n5431) );
  NAND2_X1 U6902 ( .A1(n5456), .A2(n5431), .ZN(n8806) );
  OR2_X1 U6903 ( .A1(n5692), .A2(n8806), .ZN(n5435) );
  NAND2_X1 U6904 ( .A1(n5791), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5434) );
  NAND2_X1 U6905 ( .A1(n5534), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5433) );
  INV_X1 U6906 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9197) );
  OR2_X1 U6907 ( .A1(n5142), .A2(n9197), .ZN(n5432) );
  NAND4_X1 U6908 ( .A1(n5435), .A2(n5434), .A3(n5433), .A4(n5432), .ZN(n9158)
         );
  NAND2_X1 U6909 ( .A1(n9158), .A2(n5752), .ZN(n5436) );
  NAND2_X1 U6910 ( .A1(n5437), .A2(n5436), .ZN(n5438) );
  XNOR2_X1 U6911 ( .A(n5438), .B(n5049), .ZN(n8799) );
  NAND2_X1 U6912 ( .A1(n9519), .A2(n5752), .ZN(n5440) );
  NAND2_X1 U6913 ( .A1(n9158), .A2(n5747), .ZN(n5439) );
  NAND2_X1 U6914 ( .A1(n5440), .A2(n5439), .ZN(n8800) );
  INV_X1 U6915 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5445) );
  MUX2_X1 U6916 ( .A(n9999), .B(n5445), .S(n5634), .Z(n5472) );
  XNOR2_X1 U6917 ( .A(n5472), .B(SI_17_), .ZN(n5471) );
  XNOR2_X1 U6918 ( .A(n5476), .B(n5471), .ZN(n7024) );
  NAND2_X1 U6919 ( .A1(n7024), .A2(n8882), .ZN(n5454) );
  AND2_X1 U6920 ( .A1(n5006), .A2(n5446), .ZN(n5448) );
  NAND2_X1 U6921 ( .A1(n4452), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5451) );
  INV_X1 U6922 ( .A(n5451), .ZN(n5449) );
  NAND2_X1 U6923 ( .A1(n5449), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U6924 ( .A1(n5451), .A2(n5450), .ZN(n5477) );
  AOI22_X1 U6925 ( .A1(n5614), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5507), .B2(
        n9202), .ZN(n5453) );
  NAND2_X1 U6926 ( .A1(n9514), .A2(n5753), .ZN(n5464) );
  NAND2_X1 U6927 ( .A1(n5534), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5462) );
  INV_X1 U6928 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5455) );
  NAND2_X1 U6929 ( .A1(n5456), .A2(n5455), .ZN(n5457) );
  AND2_X1 U6930 ( .A1(n5484), .A2(n5457), .ZN(n8820) );
  NAND2_X1 U6931 ( .A1(n5098), .A2(n8820), .ZN(n5461) );
  INV_X1 U6932 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n5458) );
  OR2_X1 U6933 ( .A1(n5057), .A2(n5458), .ZN(n5460) );
  INV_X1 U6934 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9199) );
  OR2_X1 U6935 ( .A1(n5142), .A2(n9199), .ZN(n5459) );
  NAND4_X1 U6936 ( .A1(n5462), .A2(n5461), .A3(n5460), .A4(n5459), .ZN(n9436)
         );
  NAND2_X1 U6937 ( .A1(n9436), .A2(n5752), .ZN(n5463) );
  NAND2_X1 U6938 ( .A1(n5464), .A2(n5463), .ZN(n5465) );
  XNOR2_X1 U6939 ( .A(n5465), .B(n5750), .ZN(n5469) );
  AND2_X1 U6940 ( .A1(n9436), .A2(n5747), .ZN(n5466) );
  AOI21_X1 U6941 ( .B1(n9514), .B2(n5752), .A(n5466), .ZN(n5468) );
  XNOR2_X1 U6942 ( .A(n5469), .B(n5468), .ZN(n8813) );
  NAND2_X1 U6943 ( .A1(n5469), .A2(n5468), .ZN(n5470) );
  INV_X1 U6944 ( .A(n5471), .ZN(n5475) );
  INV_X1 U6945 ( .A(n5472), .ZN(n5473) );
  NAND2_X1 U6946 ( .A1(n5473), .A2(SI_17_), .ZN(n5474) );
  MUX2_X1 U6947 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5634), .Z(n5501) );
  XNOR2_X1 U6948 ( .A(n5501), .B(SI_18_), .ZN(n5498) );
  XNOR2_X1 U6949 ( .A(n5500), .B(n5498), .ZN(n7285) );
  NAND2_X1 U6950 ( .A1(n7285), .A2(n8882), .ZN(n5480) );
  NAND2_X1 U6951 ( .A1(n5477), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5478) );
  XNOR2_X1 U6952 ( .A(n5478), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9205) );
  AOI22_X1 U6953 ( .A1(n5614), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5507), .B2(
        n9205), .ZN(n5479) );
  NAND2_X1 U6954 ( .A1(n9509), .A2(n5753), .ZN(n5489) );
  INV_X1 U6955 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9427) );
  NAND2_X1 U6956 ( .A1(n5534), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5482) );
  NAND2_X1 U6957 ( .A1(n5791), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5481) );
  AND2_X1 U6958 ( .A1(n5482), .A2(n5481), .ZN(n5487) );
  INV_X1 U6959 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n10012) );
  NAND2_X1 U6960 ( .A1(n5484), .A2(n10012), .ZN(n5485) );
  NAND2_X1 U6961 ( .A1(n5511), .A2(n5485), .ZN(n9426) );
  OR2_X1 U6962 ( .A1(n9426), .A2(n5692), .ZN(n5486) );
  OAI211_X1 U6963 ( .C1(n5142), .C2(n9427), .A(n5487), .B(n5486), .ZN(n9410)
         );
  NAND2_X1 U6964 ( .A1(n9410), .A2(n5752), .ZN(n5488) );
  NAND2_X1 U6965 ( .A1(n5489), .A2(n5488), .ZN(n5490) );
  XNOR2_X1 U6966 ( .A(n5490), .B(n5750), .ZN(n5494) );
  NAND2_X1 U6967 ( .A1(n5493), .A2(n5494), .ZN(n8861) );
  NAND2_X1 U6968 ( .A1(n9509), .A2(n5752), .ZN(n5492) );
  NAND2_X1 U6969 ( .A1(n9410), .A2(n5747), .ZN(n5491) );
  NAND2_X1 U6970 ( .A1(n5492), .A2(n5491), .ZN(n8864) );
  NAND2_X1 U6971 ( .A1(n8861), .A2(n8864), .ZN(n5497) );
  INV_X1 U6972 ( .A(n5493), .ZN(n5496) );
  NAND2_X1 U6973 ( .A1(n5496), .A2(n5495), .ZN(n8862) );
  NAND2_X1 U6974 ( .A1(n5497), .A2(n8862), .ZN(n8772) );
  NAND2_X1 U6975 ( .A1(n5501), .A2(SI_18_), .ZN(n5502) );
  MUX2_X1 U6976 ( .A(n7353), .B(n7355), .S(n5634), .Z(n5504) );
  INV_X1 U6977 ( .A(SI_19_), .ZN(n5503) );
  NAND2_X1 U6978 ( .A1(n5504), .A2(n5503), .ZN(n5525) );
  INV_X1 U6979 ( .A(n5504), .ZN(n5505) );
  NAND2_X1 U6980 ( .A1(n5505), .A2(SI_19_), .ZN(n5506) );
  NAND2_X1 U6981 ( .A1(n5525), .A2(n5506), .ZN(n5526) );
  XNOR2_X1 U6982 ( .A(n5527), .B(n5526), .ZN(n7352) );
  NAND2_X1 U6983 ( .A1(n7352), .A2(n8882), .ZN(n5509) );
  AOI22_X1 U6984 ( .A1(n5614), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5507), .B2(
        n7289), .ZN(n5508) );
  NAND2_X1 U6985 ( .A1(n9501), .A2(n5753), .ZN(n5516) );
  INV_X1 U6986 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U6987 ( .A1(n5511), .A2(n5510), .ZN(n5512) );
  NAND2_X1 U6988 ( .A1(n5537), .A2(n5512), .ZN(n9401) );
  AOI22_X1 U6989 ( .A1(n5534), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n5791), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n5514) );
  NAND2_X1 U6990 ( .A1(n5792), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5513) );
  OAI211_X1 U6991 ( .C1(n9401), .C2(n5692), .A(n5514), .B(n5513), .ZN(n9439)
         );
  NAND2_X1 U6992 ( .A1(n9439), .A2(n5752), .ZN(n5515) );
  NAND2_X1 U6993 ( .A1(n5516), .A2(n5515), .ZN(n5517) );
  XNOR2_X1 U6994 ( .A(n5517), .B(n5750), .ZN(n5519) );
  AND2_X1 U6995 ( .A1(n9439), .A2(n5747), .ZN(n5518) );
  AOI21_X1 U6996 ( .B1(n9501), .B2(n5752), .A(n5518), .ZN(n5520) );
  NAND2_X1 U6997 ( .A1(n5519), .A2(n5520), .ZN(n5524) );
  INV_X1 U6998 ( .A(n5519), .ZN(n5522) );
  INV_X1 U6999 ( .A(n5520), .ZN(n5521) );
  NAND2_X1 U7000 ( .A1(n5522), .A2(n5521), .ZN(n5523) );
  NAND2_X1 U7001 ( .A1(n5524), .A2(n5523), .ZN(n8775) );
  MUX2_X1 U7002 ( .A(n6089), .B(n7488), .S(n5634), .Z(n5529) );
  INV_X1 U7003 ( .A(SI_20_), .ZN(n5528) );
  NAND2_X1 U7004 ( .A1(n5529), .A2(n5528), .ZN(n5553) );
  INV_X1 U7005 ( .A(n5529), .ZN(n5530) );
  NAND2_X1 U7006 ( .A1(n5530), .A2(SI_20_), .ZN(n5531) );
  XNOR2_X1 U7007 ( .A(n5552), .B(n5551), .ZN(n9955) );
  NAND2_X1 U7008 ( .A1(n9955), .A2(n8882), .ZN(n5533) );
  NAND2_X1 U7009 ( .A1(n5614), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U7010 ( .A1(n9496), .A2(n5753), .ZN(n5543) );
  INV_X1 U7011 ( .A(n5534), .ZN(n5795) );
  INV_X1 U7012 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5541) );
  INV_X1 U7013 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5536) );
  NAND2_X1 U7014 ( .A1(n5537), .A2(n5536), .ZN(n5538) );
  NAND2_X1 U7015 ( .A1(n5557), .A2(n5538), .ZN(n9384) );
  OR2_X1 U7016 ( .A1(n9384), .A2(n5692), .ZN(n5540) );
  AOI22_X1 U7017 ( .A1(n5792), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n5791), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n5539) );
  OAI211_X1 U7018 ( .C1(n5795), .C2(n5541), .A(n5540), .B(n5539), .ZN(n9409)
         );
  NAND2_X1 U7019 ( .A1(n9409), .A2(n5752), .ZN(n5542) );
  NAND2_X1 U7020 ( .A1(n5543), .A2(n5542), .ZN(n5544) );
  XNOR2_X1 U7021 ( .A(n5544), .B(n5049), .ZN(n5547) );
  NAND2_X1 U7022 ( .A1(n9496), .A2(n5752), .ZN(n5546) );
  NAND2_X1 U7023 ( .A1(n9409), .A2(n5747), .ZN(n5545) );
  NAND2_X1 U7024 ( .A1(n5546), .A2(n5545), .ZN(n5548) );
  NAND2_X1 U7025 ( .A1(n5547), .A2(n5548), .ZN(n8832) );
  INV_X1 U7026 ( .A(n5547), .ZN(n5550) );
  INV_X1 U7027 ( .A(n5548), .ZN(n5549) );
  NAND2_X1 U7028 ( .A1(n5550), .A2(n5549), .ZN(n8834) );
  NAND2_X1 U7029 ( .A1(n8830), .A2(n8834), .ZN(n8781) );
  MUX2_X1 U7030 ( .A(n10066), .B(n7554), .S(n5634), .Z(n5570) );
  XNOR2_X1 U7031 ( .A(n5570), .B(SI_21_), .ZN(n5569) );
  XNOR2_X1 U7032 ( .A(n5568), .B(n5569), .ZN(n7553) );
  NAND2_X1 U7033 ( .A1(n7553), .A2(n8882), .ZN(n5556) );
  NAND2_X1 U7034 ( .A1(n5614), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5555) );
  NAND2_X1 U7035 ( .A1(n9493), .A2(n5753), .ZN(n5565) );
  INV_X1 U7036 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8785) );
  NAND2_X1 U7037 ( .A1(n5557), .A2(n8785), .ZN(n5558) );
  NAND2_X1 U7038 ( .A1(n5579), .A2(n5558), .ZN(n9373) );
  OR2_X1 U7039 ( .A1(n9373), .A2(n5692), .ZN(n5563) );
  INV_X1 U7040 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n10203) );
  NAND2_X1 U7041 ( .A1(n5791), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5560) );
  NAND2_X1 U7042 ( .A1(n5534), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5559) );
  OAI211_X1 U7043 ( .C1(n5142), .C2(n10203), .A(n5560), .B(n5559), .ZN(n5561)
         );
  INV_X1 U7044 ( .A(n5561), .ZN(n5562) );
  NAND2_X1 U7045 ( .A1(n5563), .A2(n5562), .ZN(n9388) );
  NAND2_X1 U7046 ( .A1(n9388), .A2(n5699), .ZN(n5564) );
  NAND2_X1 U7047 ( .A1(n5565), .A2(n5564), .ZN(n5566) );
  XNOR2_X1 U7048 ( .A(n5566), .B(n5049), .ZN(n5590) );
  AND2_X1 U7049 ( .A1(n9388), .A2(n5747), .ZN(n5567) );
  AOI21_X1 U7050 ( .B1(n9493), .B2(n5752), .A(n5567), .ZN(n5591) );
  XNOR2_X1 U7051 ( .A(n5590), .B(n5591), .ZN(n8783) );
  INV_X1 U7052 ( .A(n5570), .ZN(n5571) );
  NAND2_X1 U7053 ( .A1(n5571), .A2(SI_21_), .ZN(n5572) );
  MUX2_X1 U7054 ( .A(n7651), .B(n10230), .S(n5634), .Z(n5574) );
  INV_X1 U7055 ( .A(SI_22_), .ZN(n5573) );
  NAND2_X1 U7056 ( .A1(n5574), .A2(n5573), .ZN(n5603) );
  INV_X1 U7057 ( .A(n5574), .ZN(n5575) );
  NAND2_X1 U7058 ( .A1(n5575), .A2(SI_22_), .ZN(n5576) );
  NAND2_X1 U7059 ( .A1(n5603), .A2(n5576), .ZN(n5604) );
  XNOR2_X1 U7060 ( .A(n5605), .B(n5604), .ZN(n7649) );
  NAND2_X1 U7061 ( .A1(n7649), .A2(n8882), .ZN(n5578) );
  NAND2_X1 U7062 ( .A1(n5614), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5577) );
  INV_X1 U7063 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8852) );
  NAND2_X1 U7064 ( .A1(n5579), .A2(n8852), .ZN(n5580) );
  NAND2_X1 U7065 ( .A1(n5619), .A2(n5580), .ZN(n9347) );
  INV_X1 U7066 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n10055) );
  NAND2_X1 U7067 ( .A1(n5792), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U7068 ( .A1(n5791), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5581) );
  OAI211_X1 U7069 ( .C1(n5795), .C2(n10055), .A(n5582), .B(n5581), .ZN(n5583)
         );
  INV_X1 U7070 ( .A(n5583), .ZN(n5584) );
  AND2_X1 U7071 ( .A1(n9337), .A2(n5747), .ZN(n5585) );
  AOI21_X1 U7072 ( .B1(n9486), .B2(n5752), .A(n5585), .ZN(n5597) );
  AND2_X1 U7073 ( .A1(n8783), .A2(n5597), .ZN(n5586) );
  NAND2_X1 U7074 ( .A1(n8781), .A2(n5586), .ZN(n8842) );
  NAND2_X1 U7075 ( .A1(n9486), .A2(n5753), .ZN(n5588) );
  NAND2_X1 U7076 ( .A1(n9337), .A2(n5752), .ZN(n5587) );
  NAND2_X1 U7077 ( .A1(n5588), .A2(n5587), .ZN(n5589) );
  XNOR2_X1 U7078 ( .A(n5589), .B(n5049), .ZN(n8845) );
  INV_X1 U7079 ( .A(n5597), .ZN(n5593) );
  INV_X1 U7080 ( .A(n5590), .ZN(n5592) );
  NAND2_X1 U7081 ( .A1(n5592), .A2(n5591), .ZN(n5595) );
  OR2_X1 U7082 ( .A1(n5593), .A2(n5595), .ZN(n8841) );
  AND2_X1 U7083 ( .A1(n8845), .A2(n8841), .ZN(n5594) );
  INV_X1 U7084 ( .A(n5595), .ZN(n5596) );
  OR2_X1 U7085 ( .A1(n5597), .A2(n5596), .ZN(n5600) );
  INV_X1 U7086 ( .A(n5600), .ZN(n5598) );
  AND2_X1 U7087 ( .A1(n8834), .A2(n5598), .ZN(n5599) );
  NAND2_X1 U7088 ( .A1(n8830), .A2(n5599), .ZN(n5602) );
  OR2_X1 U7089 ( .A1(n5600), .A2(n8783), .ZN(n5601) );
  INV_X1 U7090 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5606) );
  MUX2_X1 U7091 ( .A(n7729), .B(n5606), .S(n5634), .Z(n5608) );
  INV_X1 U7092 ( .A(SI_23_), .ZN(n5607) );
  NAND2_X1 U7093 ( .A1(n5608), .A2(n5607), .ZN(n5632) );
  INV_X1 U7094 ( .A(n5608), .ZN(n5609) );
  NAND2_X1 U7095 ( .A1(n5609), .A2(SI_23_), .ZN(n5610) );
  OR2_X1 U7096 ( .A1(n5612), .A2(n5611), .ZN(n5613) );
  NAND2_X1 U7097 ( .A1(n5633), .A2(n5613), .ZN(n7725) );
  NAND2_X1 U7098 ( .A1(n7725), .A2(n8882), .ZN(n5616) );
  NAND2_X1 U7099 ( .A1(n5614), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5615) );
  NAND2_X1 U7100 ( .A1(n9481), .A2(n5753), .ZN(n5627) );
  INV_X1 U7101 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U7102 ( .A1(n5619), .A2(n5618), .ZN(n5620) );
  NAND2_X1 U7103 ( .A1(n5639), .A2(n5620), .ZN(n9330) );
  OR2_X1 U7104 ( .A1(n9330), .A2(n5692), .ZN(n5625) );
  INV_X1 U7105 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10069) );
  NAND2_X1 U7106 ( .A1(n5058), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5622) );
  NAND2_X1 U7107 ( .A1(n5792), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5621) );
  OAI211_X1 U7108 ( .C1(n5057), .C2(n10069), .A(n5622), .B(n5621), .ZN(n5623)
         );
  INV_X1 U7109 ( .A(n5623), .ZN(n5624) );
  NAND2_X1 U7110 ( .A1(n9354), .A2(n5752), .ZN(n5626) );
  NAND2_X1 U7111 ( .A1(n5627), .A2(n5626), .ZN(n5628) );
  XNOR2_X1 U7112 ( .A(n5628), .B(n5750), .ZN(n5631) );
  AOI21_X2 U7113 ( .B1(n8844), .B2(n8846), .A(n5631), .ZN(n8762) );
  INV_X1 U7114 ( .A(n9481), .ZN(n9333) );
  OAI22_X1 U7115 ( .A1(n9333), .A2(n5630), .B1(n9314), .B2(n5629), .ZN(n8764)
         );
  NAND3_X1 U7116 ( .A1(n8844), .A2(n5631), .A3(n8846), .ZN(n8761) );
  INV_X1 U7117 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7838) );
  MUX2_X1 U7118 ( .A(n7835), .B(n7838), .S(n5634), .Z(n5655) );
  XNOR2_X1 U7119 ( .A(n5655), .B(SI_24_), .ZN(n5652) );
  XNOR2_X1 U7120 ( .A(n5654), .B(n5652), .ZN(n7834) );
  NAND2_X1 U7121 ( .A1(n7834), .A2(n8882), .ZN(n5636) );
  NAND2_X1 U7122 ( .A1(n5614), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5635) );
  NAND2_X1 U7123 ( .A1(n9478), .A2(n5753), .ZN(n5647) );
  INV_X1 U7124 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U7125 ( .A1(n5639), .A2(n5638), .ZN(n5640) );
  NAND2_X1 U7126 ( .A1(n5665), .A2(n5640), .ZN(n9310) );
  OR2_X1 U7127 ( .A1(n9310), .A2(n5692), .ZN(n5645) );
  INV_X1 U7128 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n10014) );
  NAND2_X1 U7129 ( .A1(n5058), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5642) );
  NAND2_X1 U7130 ( .A1(n5791), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5641) );
  OAI211_X1 U7131 ( .C1(n10014), .C2(n5142), .A(n5642), .B(n5641), .ZN(n5643)
         );
  INV_X1 U7132 ( .A(n5643), .ZN(n5644) );
  NAND2_X1 U7133 ( .A1(n9338), .A2(n5699), .ZN(n5646) );
  NAND2_X1 U7134 ( .A1(n5647), .A2(n5646), .ZN(n5648) );
  XNOR2_X1 U7135 ( .A(n5648), .B(n5049), .ZN(n5649) );
  AOI22_X1 U7136 ( .A1(n9478), .A2(n5752), .B1(n5747), .B2(n9338), .ZN(n5650)
         );
  XNOR2_X1 U7137 ( .A(n5649), .B(n5650), .ZN(n8824) );
  INV_X1 U7138 ( .A(n5649), .ZN(n5651) );
  INV_X1 U7139 ( .A(n5652), .ZN(n5653) );
  INV_X1 U7140 ( .A(n5655), .ZN(n5656) );
  NAND2_X1 U7141 ( .A1(n5656), .A2(SI_24_), .ZN(n5657) );
  MUX2_X1 U7142 ( .A(n10086), .B(n10223), .S(n5634), .Z(n5659) );
  INV_X1 U7143 ( .A(SI_25_), .ZN(n5658) );
  NAND2_X1 U7144 ( .A1(n5659), .A2(n5658), .ZN(n5679) );
  INV_X1 U7145 ( .A(n5659), .ZN(n5660) );
  NAND2_X1 U7146 ( .A1(n5660), .A2(SI_25_), .ZN(n5661) );
  NAND2_X1 U7147 ( .A1(n5679), .A2(n5661), .ZN(n5680) );
  NAND2_X1 U7148 ( .A1(n7943), .A2(n8882), .ZN(n5663) );
  NAND2_X1 U7149 ( .A1(n5614), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5662) );
  INV_X1 U7150 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5664) );
  NAND2_X1 U7151 ( .A1(n5665), .A2(n5664), .ZN(n5666) );
  NAND2_X1 U7152 ( .A1(n9303), .A2(n5098), .ZN(n5671) );
  INV_X1 U7153 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n10052) );
  NAND2_X1 U7154 ( .A1(n5792), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5668) );
  NAND2_X1 U7155 ( .A1(n5791), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5667) );
  OAI211_X1 U7156 ( .C1(n5795), .C2(n10052), .A(n5668), .B(n5667), .ZN(n5669)
         );
  INV_X1 U7157 ( .A(n5669), .ZN(n5670) );
  AOI22_X1 U7158 ( .A1(n9472), .A2(n5752), .B1(n5747), .B2(n9288), .ZN(n5675)
         );
  NAND2_X1 U7159 ( .A1(n9472), .A2(n5753), .ZN(n5673) );
  NAND2_X1 U7160 ( .A1(n9288), .A2(n5752), .ZN(n5672) );
  NAND2_X1 U7161 ( .A1(n5673), .A2(n5672), .ZN(n5674) );
  XNOR2_X1 U7162 ( .A(n5674), .B(n5049), .ZN(n5677) );
  XOR2_X1 U7163 ( .A(n5675), .B(n5677), .Z(n8791) );
  INV_X1 U7164 ( .A(n5675), .ZN(n5676) );
  INV_X1 U7165 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7977) );
  INV_X1 U7166 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7973) );
  MUX2_X1 U7167 ( .A(n7977), .B(n7973), .S(n5634), .Z(n5683) );
  INV_X1 U7168 ( .A(SI_26_), .ZN(n5682) );
  NAND2_X1 U7169 ( .A1(n5683), .A2(n5682), .ZN(n5709) );
  INV_X1 U7170 ( .A(n5683), .ZN(n5684) );
  NAND2_X1 U7171 ( .A1(n5684), .A2(SI_26_), .ZN(n5685) );
  XNOR2_X1 U7172 ( .A(n5708), .B(n5707), .ZN(n7972) );
  NAND2_X1 U7173 ( .A1(n7972), .A2(n8882), .ZN(n5687) );
  NAND2_X1 U7174 ( .A1(n5614), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5686) );
  INV_X1 U7175 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5689) );
  NAND2_X1 U7176 ( .A1(n5690), .A2(n5689), .ZN(n5691) );
  NAND2_X1 U7177 ( .A1(n5739), .A2(n5691), .ZN(n6424) );
  OR2_X1 U7178 ( .A1(n6424), .A2(n5692), .ZN(n5697) );
  INV_X1 U7179 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10143) );
  NAND2_X1 U7180 ( .A1(n5534), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5694) );
  NAND2_X1 U7181 ( .A1(n5792), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5693) );
  OAI211_X1 U7182 ( .C1(n5057), .C2(n10143), .A(n5694), .B(n5693), .ZN(n5695)
         );
  INV_X1 U7183 ( .A(n5695), .ZN(n5696) );
  AND2_X1 U7184 ( .A1(n9299), .A2(n5747), .ZN(n5698) );
  AOI21_X1 U7185 ( .B1(n9465), .B2(n5699), .A(n5698), .ZN(n5703) );
  NAND2_X1 U7186 ( .A1(n9465), .A2(n5753), .ZN(n5701) );
  NAND2_X1 U7187 ( .A1(n9299), .A2(n5699), .ZN(n5700) );
  NAND2_X1 U7188 ( .A1(n5701), .A2(n5700), .ZN(n5702) );
  XNOR2_X1 U7189 ( .A(n5702), .B(n5049), .ZN(n5705) );
  XOR2_X1 U7190 ( .A(n5703), .B(n5705), .Z(n6421) );
  INV_X1 U7191 ( .A(n5703), .ZN(n5704) );
  NAND2_X1 U7192 ( .A1(n5708), .A2(n5707), .ZN(n5710) );
  NAND2_X1 U7193 ( .A1(n5710), .A2(n5709), .ZN(n5716) );
  INV_X1 U7194 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8006) );
  INV_X1 U7195 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5711) );
  MUX2_X1 U7196 ( .A(n8006), .B(n5711), .S(n5634), .Z(n5712) );
  INV_X1 U7197 ( .A(SI_27_), .ZN(n10125) );
  NAND2_X1 U7198 ( .A1(n5712), .A2(n10125), .ZN(n5731) );
  INV_X1 U7199 ( .A(n5712), .ZN(n5713) );
  NAND2_X1 U7200 ( .A1(n5713), .A2(SI_27_), .ZN(n5714) );
  OR2_X1 U7201 ( .A1(n5716), .A2(n5715), .ZN(n5717) );
  NAND2_X1 U7202 ( .A1(n5732), .A2(n5717), .ZN(n7989) );
  NAND2_X1 U7203 ( .A1(n7989), .A2(n8882), .ZN(n5719) );
  NAND2_X1 U7204 ( .A1(n5614), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5718) );
  NAND2_X1 U7205 ( .A1(n9460), .A2(n5753), .ZN(n5727) );
  XNOR2_X1 U7206 ( .A(n5739), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U7207 ( .A1(n8755), .A2(n5098), .ZN(n5725) );
  INV_X1 U7208 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n5722) );
  NAND2_X1 U7209 ( .A1(n5058), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5721) );
  NAND2_X1 U7210 ( .A1(n5791), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5720) );
  OAI211_X1 U7211 ( .C1(n5722), .C2(n5142), .A(n5721), .B(n5720), .ZN(n5723)
         );
  INV_X1 U7212 ( .A(n5723), .ZN(n5724) );
  NAND2_X1 U7213 ( .A1(n9282), .A2(n5699), .ZN(n5726) );
  NAND2_X1 U7214 ( .A1(n5727), .A2(n5726), .ZN(n5728) );
  XNOR2_X1 U7215 ( .A(n5728), .B(n5049), .ZN(n5781) );
  NAND2_X1 U7216 ( .A1(n9460), .A2(n5699), .ZN(n5730) );
  NAND2_X1 U7217 ( .A1(n9282), .A2(n5747), .ZN(n5729) );
  NAND2_X1 U7218 ( .A1(n5730), .A2(n5729), .ZN(n5782) );
  NAND2_X1 U7219 ( .A1(n5781), .A2(n5782), .ZN(n8751) );
  NAND2_X1 U7220 ( .A1(n8754), .A2(n8751), .ZN(n5816) );
  INV_X1 U7221 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n10144) );
  INV_X1 U7222 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5733) );
  MUX2_X1 U7223 ( .A(n10144), .B(n5733), .S(n5634), .Z(n6186) );
  XNOR2_X1 U7224 ( .A(n6186), .B(SI_28_), .ZN(n6183) );
  NAND2_X1 U7225 ( .A1(n8007), .A2(n8882), .ZN(n5735) );
  NAND2_X1 U7226 ( .A1(n5614), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5734) );
  NAND2_X1 U7227 ( .A1(n9455), .A2(n5752), .ZN(n5749) );
  INV_X1 U7228 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5737) );
  INV_X1 U7229 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5736) );
  OAI21_X1 U7230 ( .B1(n5739), .B2(n5737), .A(n5736), .ZN(n5740) );
  NAND2_X1 U7231 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5738) );
  NAND2_X1 U7232 ( .A1(n9270), .A2(n5098), .ZN(n5746) );
  INV_X1 U7233 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5743) );
  NAND2_X1 U7234 ( .A1(n5792), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5742) );
  NAND2_X1 U7235 ( .A1(n5791), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5741) );
  OAI211_X1 U7236 ( .C1(n5795), .C2(n5743), .A(n5742), .B(n5741), .ZN(n5744)
         );
  INV_X1 U7237 ( .A(n5744), .ZN(n5745) );
  NAND2_X1 U7238 ( .A1(n9157), .A2(n5747), .ZN(n5748) );
  NAND2_X1 U7239 ( .A1(n5749), .A2(n5748), .ZN(n5751) );
  XNOR2_X1 U7240 ( .A(n5751), .B(n5750), .ZN(n5755) );
  AOI22_X1 U7241 ( .A1(n9455), .A2(n5753), .B1(n5752), .B2(n9157), .ZN(n5754)
         );
  XNOR2_X1 U7242 ( .A(n5755), .B(n5754), .ZN(n5810) );
  INV_X1 U7243 ( .A(n5810), .ZN(n5780) );
  NAND3_X1 U7244 ( .A1(n7944), .A2(P1_B_REG_SCAN_IN), .A3(n7839), .ZN(n5756)
         );
  OAI21_X1 U7245 ( .B1(P1_B_REG_SCAN_IN), .B2(n7839), .A(n5756), .ZN(n5757) );
  INV_X1 U7246 ( .A(n5770), .ZN(n7974) );
  INV_X1 U7247 ( .A(n7839), .ZN(n5758) );
  OAI22_X1 U7248 ( .A1(n9755), .A2(P1_D_REG_0__SCAN_IN), .B1(n5770), .B2(n5758), .ZN(n6978) );
  INV_X1 U7249 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10096) );
  INV_X1 U7250 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10081) );
  INV_X1 U7251 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10132) );
  INV_X1 U7252 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n9996) );
  NAND4_X1 U7253 ( .A1(n10096), .A2(n10081), .A3(n10132), .A4(n9996), .ZN(
        n5759) );
  NOR3_X1 U7254 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        n5759), .ZN(n10236) );
  NOR4_X1 U7255 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n5761) );
  NOR4_X1 U7256 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n5760) );
  NAND3_X1 U7257 ( .A1(n10236), .A2(n5761), .A3(n5760), .ZN(n5767) );
  NOR4_X1 U7258 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n5765) );
  NOR4_X1 U7259 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5764) );
  NOR4_X1 U7260 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5763) );
  NOR4_X1 U7261 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n5762) );
  NAND4_X1 U7262 ( .A1(n5765), .A2(n5764), .A3(n5763), .A4(n5762), .ZN(n5766)
         );
  NOR2_X1 U7263 ( .A1(n5767), .A2(n5766), .ZN(n5768) );
  NOR2_X1 U7264 ( .A1(n9755), .A2(n5768), .ZN(n6977) );
  OR2_X1 U7265 ( .A1(n6978), .A2(n6977), .ZN(n7042) );
  INV_X1 U7266 ( .A(n7944), .ZN(n5769) );
  OAI22_X1 U7267 ( .A1(n9755), .A2(P1_D_REG_1__SCAN_IN), .B1(n5770), .B2(n5769), .ZN(n7039) );
  NOR2_X1 U7268 ( .A1(n7042), .A2(n7039), .ZN(n5807) );
  INV_X1 U7269 ( .A(n5771), .ZN(n5772) );
  NAND2_X1 U7270 ( .A1(n5772), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5773) );
  MUX2_X1 U7271 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5773), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n5774) );
  NAND2_X1 U7272 ( .A1(n5774), .A2(n4984), .ZN(n6431) );
  AND2_X1 U7273 ( .A1(n6431), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5775) );
  AND2_X1 U7274 ( .A1(n5807), .A2(n9756), .ZN(n5800) );
  NAND2_X1 U7275 ( .A1(n9071), .A2(n9106), .ZN(n7072) );
  AND2_X1 U7276 ( .A1(n9774), .A2(n6997), .ZN(n5779) );
  NAND2_X1 U7277 ( .A1(n5780), .A2(n8850), .ZN(n5815) );
  INV_X1 U7278 ( .A(n5781), .ZN(n5784) );
  INV_X1 U7279 ( .A(n5782), .ZN(n5783) );
  NAND2_X1 U7280 ( .A1(n5784), .A2(n5783), .ZN(n8752) );
  AND2_X1 U7281 ( .A1(n5810), .A2(n5785), .ZN(n5786) );
  NAND2_X1 U7282 ( .A1(n5816), .A2(n5786), .ZN(n5814) );
  OR2_X1 U7283 ( .A1(n6997), .A2(n5787), .ZN(n5801) );
  NAND2_X1 U7284 ( .A1(n5801), .A2(n9756), .ZN(n7041) );
  NOR2_X1 U7285 ( .A1(n7041), .A2(n9774), .ZN(n5789) );
  INV_X1 U7286 ( .A(n5807), .ZN(n5802) );
  AND2_X1 U7287 ( .A1(n5802), .A2(n9756), .ZN(n5788) );
  OR2_X1 U7288 ( .A1(n7072), .A2(n7489), .ZN(n7169) );
  NAND2_X1 U7289 ( .A1(n5788), .A2(n7170), .ZN(n7150) );
  INV_X1 U7290 ( .A(n5790), .ZN(n9248) );
  INV_X1 U7291 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5796) );
  NAND2_X1 U7292 ( .A1(n5791), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U7293 ( .A1(n5792), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5793) );
  OAI211_X1 U7294 ( .C1(n5796), .C2(n5795), .A(n5794), .B(n5793), .ZN(n5797)
         );
  AOI21_X1 U7295 ( .B1(n9248), .B2(n5098), .A(n5797), .ZN(n9156) );
  OR2_X1 U7296 ( .A1(n9072), .A2(n6982), .ZN(n7161) );
  INV_X1 U7297 ( .A(n5798), .ZN(n6996) );
  NOR2_X1 U7298 ( .A1(n7161), .A2(n6996), .ZN(n5799) );
  NAND2_X1 U7299 ( .A1(n5800), .A2(n5799), .ZN(n8865) );
  AND3_X1 U7300 ( .A1(n5801), .A2(n6431), .A3(n6430), .ZN(n5803) );
  NAND2_X1 U7301 ( .A1(n9774), .A2(n5802), .ZN(n6639) );
  NAND2_X1 U7302 ( .A1(n5803), .A2(n6639), .ZN(n5804) );
  NAND2_X1 U7303 ( .A1(n5804), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5805) );
  NAND2_X1 U7304 ( .A1(n5805), .A2(n7150), .ZN(n8819) );
  AOI22_X1 U7305 ( .A1(n9270), .A2(n8819), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n5809) );
  NAND2_X1 U7306 ( .A1(n9756), .A2(n6996), .ZN(n5806) );
  NOR2_X1 U7307 ( .A1(n7161), .A2(n5806), .ZN(n9151) );
  NAND2_X1 U7308 ( .A1(n9282), .A2(n8868), .ZN(n5808) );
  OAI211_X1 U7309 ( .C1(n9156), .C2(n8865), .A(n5809), .B(n5808), .ZN(n5812)
         );
  NOR3_X1 U7310 ( .A1(n5810), .A2(n8874), .A3(n8752), .ZN(n5811) );
  AOI211_X1 U7311 ( .C1(n8872), .C2(n9455), .A(n5812), .B(n5811), .ZN(n5813)
         );
  OAI211_X1 U7312 ( .C1(n5816), .C2(n5815), .A(n5814), .B(n5813), .ZN(P1_U3218) );
  NOR2_X1 U7313 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5818) );
  NOR2_X1 U7314 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5817) );
  AND2_X1 U7315 ( .A1(n5818), .A2(n5817), .ZN(n5819) );
  AND2_X2 U7316 ( .A1(n5899), .A2(n5819), .ZN(n5844) );
  NOR2_X1 U7317 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5823) );
  NOR2_X1 U7318 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5822) );
  NOR2_X1 U7319 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5821) );
  NOR2_X1 U7320 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5820) );
  NOR2_X1 U7321 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5826) );
  NOR2_X1 U7322 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5825) );
  NOR2_X1 U7323 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n5824) );
  AND2_X2 U7324 ( .A1(n5854), .A2(n5829), .ZN(n5857) );
  INV_X1 U7325 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5832) );
  INV_X1 U7326 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n5840) );
  NAND2_X1 U7327 ( .A1(n4378), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U7328 ( .A1(n5915), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5838) );
  OAI211_X1 U7329 ( .C1(n6194), .C2(n5840), .A(n5839), .B(n5838), .ZN(n8311)
         );
  NAND2_X1 U7330 ( .A1(n6179), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5843) );
  NAND2_X1 U7331 ( .A1(n4378), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n5842) );
  NAND2_X1 U7332 ( .A1(n5915), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5841) );
  AND3_X1 U7333 ( .A1(n5843), .A2(n5842), .A3(n5841), .ZN(n6361) );
  NOR2_X1 U7334 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5847) );
  NAND2_X1 U7335 ( .A1(n6220), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5848) );
  NAND2_X1 U7336 ( .A1(n6361), .A2(n7581), .ZN(n6203) );
  NAND2_X1 U7337 ( .A1(n4378), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5853) );
  AND2_X2 U7338 ( .A1(n5837), .A2(n5849), .ZN(n5904) );
  NAND2_X1 U7339 ( .A1(n5904), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5852) );
  NAND2_X1 U7340 ( .A1(n6179), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5851) );
  NAND2_X1 U7341 ( .A1(n5915), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5850) );
  INV_X1 U7342 ( .A(n5854), .ZN(n5855) );
  INV_X1 U7343 ( .A(n5857), .ZN(n5858) );
  NAND2_X1 U7344 ( .A1(n5860), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5862) );
  OR2_X1 U7345 ( .A1(n5863), .A2(n5832), .ZN(n5888) );
  INV_X1 U7346 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5887) );
  XNOR2_X1 U7347 ( .A(n5888), .B(n5887), .ZN(n6653) );
  OR2_X1 U7348 ( .A1(n5921), .A2(n6476), .ZN(n5865) );
  OAI211_X1 U7349 ( .C1(n6557), .C2(n6653), .A(n5865), .B(n5864), .ZN(n6889)
         );
  NAND2_X1 U7350 ( .A1(n6860), .A2(n6889), .ZN(n6250) );
  INV_X1 U7351 ( .A(n6889), .ZN(n9859) );
  NAND2_X1 U7352 ( .A1(n5915), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5869) );
  NAND2_X1 U7353 ( .A1(n4378), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U7354 ( .A1(n5904), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5867) );
  NAND2_X1 U7355 ( .A1(n6179), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5866) );
  INV_X1 U7356 ( .A(n6895), .ZN(n6953) );
  INV_X1 U7357 ( .A(SI_0_), .ZN(n5871) );
  INV_X1 U7358 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5870) );
  OAI21_X1 U7359 ( .B1(n5634), .B2(n5871), .A(n5870), .ZN(n5873) );
  AND2_X1 U7360 ( .A1(n5873), .A2(n5872), .ZN(n8750) );
  MUX2_X1 U7361 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8750), .S(n6557), .Z(n9847) );
  NAND2_X1 U7362 ( .A1(n6179), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5877) );
  NAND2_X1 U7363 ( .A1(n5915), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5876) );
  NAND2_X1 U7364 ( .A1(n4378), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U7365 ( .A1(n5904), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5874) );
  INV_X1 U7366 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5878) );
  INV_X1 U7367 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6468) );
  OR2_X1 U7368 ( .A1(n5901), .A2(n6468), .ZN(n5880) );
  OAI211_X1 U7369 ( .C1(n6557), .C2(n6580), .A(n5880), .B(n5879), .ZN(n6852)
         );
  INV_X1 U7370 ( .A(n7033), .ZN(n6834) );
  INV_X1 U7371 ( .A(n4386), .ZN(n9852) );
  INV_X1 U7372 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5886) );
  NAND2_X1 U7373 ( .A1(n6179), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5884) );
  NAND2_X1 U7374 ( .A1(n5915), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5883) );
  NAND2_X1 U7375 ( .A1(n4378), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5882) );
  NAND2_X1 U7376 ( .A1(n5888), .A2(n5887), .ZN(n5889) );
  NAND2_X1 U7377 ( .A1(n5889), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5891) );
  INV_X1 U7378 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5890) );
  XNOR2_X1 U7379 ( .A(n5891), .B(n5890), .ZN(n6679) );
  OR2_X1 U7380 ( .A1(n5921), .A2(n8049), .ZN(n5893) );
  OR2_X1 U7381 ( .A1(n5901), .A2(n6484), .ZN(n5892) );
  OAI211_X1 U7382 ( .C1(n6557), .C2(n6679), .A(n5893), .B(n5892), .ZN(n7012)
         );
  NAND2_X1 U7383 ( .A1(n6942), .A2(n7012), .ZN(n6239) );
  INV_X1 U7384 ( .A(n6942), .ZN(n8327) );
  INV_X1 U7385 ( .A(n7012), .ZN(n6970) );
  NAND2_X1 U7386 ( .A1(n8327), .A2(n6970), .ZN(n6234) );
  NAND2_X1 U7387 ( .A1(n6960), .A2(n6367), .ZN(n5894) );
  NAND2_X1 U7388 ( .A1(n5915), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5898) );
  NAND2_X1 U7389 ( .A1(n4378), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5897) );
  XNOR2_X1 U7390 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6843) );
  INV_X1 U7391 ( .A(n6843), .ZN(n6939) );
  NAND2_X1 U7392 ( .A1(n5904), .A2(n6939), .ZN(n5896) );
  NAND2_X1 U7393 ( .A1(n6179), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5895) );
  OR2_X1 U7394 ( .A1(n5899), .A2(n5832), .ZN(n5900) );
  XNOR2_X1 U7395 ( .A(n5900), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6655) );
  INV_X1 U7396 ( .A(n6655), .ZN(n6667) );
  OR2_X1 U7397 ( .A1(n5921), .A2(n6482), .ZN(n5903) );
  INV_X1 U7398 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6483) );
  OR2_X1 U7399 ( .A1(n5901), .A2(n6483), .ZN(n5902) );
  OAI211_X1 U7400 ( .C1(n6557), .C2(n6667), .A(n5903), .B(n5902), .ZN(n9867)
         );
  NAND2_X1 U7401 ( .A1(n7262), .A2(n9867), .ZN(n6366) );
  INV_X1 U7402 ( .A(n7262), .ZN(n8326) );
  INV_X1 U7403 ( .A(n9867), .ZN(n7085) );
  NAND2_X1 U7404 ( .A1(n8326), .A2(n7085), .ZN(n7258) );
  NAND2_X1 U7405 ( .A1(n5915), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5909) );
  NAND2_X1 U7406 ( .A1(n4378), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5908) );
  AOI21_X1 U7407 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5905) );
  NOR2_X1 U7408 ( .A1(n5905), .A2(n5916), .ZN(n9809) );
  NAND2_X1 U7409 ( .A1(n5904), .A2(n9809), .ZN(n5907) );
  NAND2_X1 U7410 ( .A1(n6179), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5906) );
  NAND4_X1 U7411 ( .A1(n5909), .A2(n5908), .A3(n5907), .A4(n5906), .ZN(n8325)
         );
  INV_X1 U7412 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5910) );
  NAND2_X1 U7413 ( .A1(n5899), .A2(n5910), .ZN(n5912) );
  NAND2_X1 U7414 ( .A1(n5912), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5911) );
  MUX2_X1 U7415 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5911), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5913) );
  INV_X1 U7416 ( .A(n6578), .ZN(n6619) );
  OR2_X1 U7417 ( .A1(n6478), .A2(n5921), .ZN(n5914) );
  INV_X1 U7418 ( .A(n8325), .ZN(n7140) );
  NAND2_X1 U7419 ( .A1(n7140), .A2(n9807), .ZN(n6370) );
  NAND2_X1 U7420 ( .A1(n5915), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5920) );
  NAND2_X1 U7421 ( .A1(n4378), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U7422 ( .A1(n5916), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5931) );
  OAI21_X1 U7423 ( .B1(n5916), .B2(P2_REG3_REG_6__SCAN_IN), .A(n5931), .ZN(
        n7095) );
  INV_X1 U7424 ( .A(n7095), .ZN(n7137) );
  NAND2_X1 U7425 ( .A1(n5904), .A2(n7137), .ZN(n5918) );
  NAND2_X1 U7426 ( .A1(n6179), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5917) );
  INV_X2 U7427 ( .A(n5921), .ZN(n5947) );
  NAND2_X1 U7428 ( .A1(n6474), .A2(n5947), .ZN(n5924) );
  NAND2_X1 U7429 ( .A1(n5926), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5922) );
  XNOR2_X1 U7430 ( .A(n5922), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6577) );
  AOI22_X1 U7431 ( .A1(n6217), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6077), .B2(
        n6577), .ZN(n5923) );
  NAND2_X1 U7432 ( .A1(n5924), .A2(n5923), .ZN(n7177) );
  NAND2_X1 U7433 ( .A1(n7263), .A2(n7177), .ZN(n6259) );
  INV_X1 U7434 ( .A(n7177), .ZN(n9876) );
  INV_X1 U7435 ( .A(n7263), .ZN(n8324) );
  NAND2_X1 U7436 ( .A1(n9876), .A2(n8324), .ZN(n6254) );
  NAND2_X1 U7437 ( .A1(n6259), .A2(n6254), .ZN(n7175) );
  INV_X1 U7438 ( .A(n7175), .ZN(n7091) );
  INV_X1 U7439 ( .A(n6259), .ZN(n5925) );
  AOI21_X1 U7440 ( .B1(n7090), .B2(n7091), .A(n5925), .ZN(n7181) );
  NAND2_X1 U7441 ( .A1(n6485), .A2(n5947), .ZN(n5929) );
  OAI21_X1 U7442 ( .B1(n5926), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5927) );
  XNOR2_X1 U7443 ( .A(n5927), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6623) );
  AOI22_X1 U7444 ( .A1(n6217), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6077), .B2(
        n6623), .ZN(n5928) );
  NAND2_X1 U7445 ( .A1(n5929), .A2(n5928), .ZN(n7384) );
  NAND2_X1 U7446 ( .A1(n4378), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5936) );
  NAND2_X1 U7447 ( .A1(n5915), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5935) );
  AND2_X1 U7448 ( .A1(n5931), .A2(n5930), .ZN(n5932) );
  NOR2_X1 U7449 ( .A1(n5941), .A2(n5932), .ZN(n7194) );
  NAND2_X1 U7450 ( .A1(n5904), .A2(n7194), .ZN(n5934) );
  NAND2_X1 U7451 ( .A1(n6179), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5933) );
  NAND2_X1 U7452 ( .A1(n7384), .A2(n7469), .ZN(n6260) );
  OR2_X1 U7453 ( .A1(n7469), .A2(n7384), .ZN(n6261) );
  AOI21_X1 U7454 ( .B1(n7181), .B2(n6260), .A(n5937), .ZN(n7390) );
  NAND2_X1 U7455 ( .A1(n6489), .A2(n5947), .ZN(n5940) );
  OR2_X1 U7456 ( .A1(n5844), .A2(n5832), .ZN(n5938) );
  XNOR2_X1 U7457 ( .A(n5938), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6744) );
  AOI22_X1 U7458 ( .A1(n6217), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6077), .B2(
        n6744), .ZN(n5939) );
  NAND2_X1 U7459 ( .A1(n5940), .A2(n5939), .ZN(n7630) );
  NAND2_X1 U7460 ( .A1(n5915), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U7461 ( .A1(n4378), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5945) );
  NOR2_X1 U7462 ( .A1(n5941), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5942) );
  OR2_X1 U7463 ( .A1(n5967), .A2(n5942), .ZN(n7395) );
  INV_X1 U7464 ( .A(n7395), .ZN(n7466) );
  NAND2_X1 U7465 ( .A1(n5904), .A2(n7466), .ZN(n5944) );
  NAND2_X1 U7466 ( .A1(n6179), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5943) );
  OR2_X1 U7467 ( .A1(n7630), .A2(n7706), .ZN(n6265) );
  NAND2_X1 U7468 ( .A1(n7630), .A2(n7706), .ZN(n6264) );
  NAND2_X1 U7469 ( .A1(n7390), .A2(n7391), .ZN(n7389) );
  NAND2_X1 U7470 ( .A1(n6505), .A2(n5947), .ZN(n5953) );
  INV_X1 U7471 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U7472 ( .A1(n5844), .A2(n5948), .ZN(n5950) );
  NAND2_X1 U7473 ( .A1(n5950), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5949) );
  MUX2_X1 U7474 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5949), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n5951) );
  AOI22_X1 U7475 ( .A1(n6217), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6077), .B2(
        n6785), .ZN(n5952) );
  NAND2_X1 U7476 ( .A1(n4378), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5958) );
  NAND2_X1 U7477 ( .A1(n6179), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5957) );
  INV_X1 U7478 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5954) );
  XNOR2_X1 U7479 ( .A(n5967), .B(n5954), .ZN(n7716) );
  NAND2_X1 U7480 ( .A1(n5904), .A2(n7716), .ZN(n5956) );
  NAND2_X1 U7481 ( .A1(n5915), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5955) );
  OR2_X1 U7482 ( .A1(n7840), .A2(n7638), .ZN(n6375) );
  NAND2_X1 U7483 ( .A1(n7840), .A2(n7638), .ZN(n6374) );
  NAND2_X1 U7484 ( .A1(n6535), .A2(n5947), .ZN(n5963) );
  NAND2_X1 U7485 ( .A1(n5987), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5960) );
  INV_X1 U7486 ( .A(n5960), .ZN(n5959) );
  NAND2_X1 U7487 ( .A1(n5959), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5961) );
  INV_X1 U7488 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5985) );
  NAND2_X1 U7489 ( .A1(n5960), .A2(n5985), .ZN(n5973) );
  AOI22_X1 U7490 ( .A1(n6217), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6077), .B2(
        n7115), .ZN(n5962) );
  NAND2_X1 U7491 ( .A1(n5963), .A2(n5962), .ZN(n7675) );
  NAND2_X1 U7492 ( .A1(n4378), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U7493 ( .A1(n5915), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5971) );
  NAND2_X1 U7494 ( .A1(n5967), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5965) );
  INV_X1 U7495 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U7496 ( .A1(n5965), .A2(n5964), .ZN(n5968) );
  AND2_X1 U7497 ( .A1(n5968), .A2(n5977), .ZN(n7643) );
  NAND2_X1 U7498 ( .A1(n5904), .A2(n7643), .ZN(n5970) );
  NAND2_X1 U7499 ( .A1(n6179), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U7500 ( .A1(n7675), .A2(n7705), .ZN(n6372) );
  OR2_X1 U7501 ( .A1(n7675), .A2(n7705), .ZN(n6373) );
  NAND2_X1 U7502 ( .A1(n6539), .A2(n5947), .ZN(n5976) );
  NAND2_X1 U7503 ( .A1(n5973), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5974) );
  XNOR2_X1 U7504 ( .A(n5974), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7277) );
  AOI22_X1 U7505 ( .A1(n6217), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6077), .B2(
        n7277), .ZN(n5975) );
  NAND2_X1 U7506 ( .A1(n4378), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U7507 ( .A1(n6179), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7508 ( .A1(n5977), .A2(n7625), .ZN(n5978) );
  NAND2_X1 U7509 ( .A1(n5992), .A2(n5978), .ZN(n7824) );
  INV_X1 U7510 ( .A(n7824), .ZN(n7623) );
  NAND2_X1 U7511 ( .A1(n5904), .A2(n7623), .ZN(n5980) );
  NAND2_X1 U7512 ( .A1(n5915), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5979) );
  OR2_X1 U7513 ( .A1(n7823), .A2(n7739), .ZN(n6274) );
  NAND2_X1 U7514 ( .A1(n7823), .A2(n7739), .ZN(n7681) );
  NAND2_X1 U7515 ( .A1(n6274), .A2(n7681), .ZN(n7745) );
  NAND2_X1 U7516 ( .A1(n6682), .A2(n5947), .ZN(n5990) );
  INV_X1 U7517 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5984) );
  NAND2_X1 U7518 ( .A1(n5985), .A2(n5984), .ZN(n5986) );
  NOR2_X1 U7519 ( .A1(n5987), .A2(n5986), .ZN(n6002) );
  OR2_X1 U7520 ( .A1(n6002), .A2(n5832), .ZN(n5988) );
  XNOR2_X1 U7521 ( .A(n5988), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7427) );
  AOI22_X1 U7522 ( .A1(n6217), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6077), .B2(
        n7427), .ZN(n5989) );
  NAND2_X1 U7523 ( .A1(n5915), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5997) );
  NAND2_X1 U7524 ( .A1(n4378), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5996) );
  NAND2_X1 U7525 ( .A1(n5992), .A2(n5991), .ZN(n5993) );
  AND2_X1 U7526 ( .A1(n6008), .A2(n5993), .ZN(n7736) );
  NAND2_X1 U7527 ( .A1(n5904), .A2(n7736), .ZN(n5995) );
  NAND2_X1 U7528 ( .A1(n6179), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5994) );
  NAND2_X1 U7529 ( .A1(n7931), .A2(n7764), .ZN(n6277) );
  INV_X1 U7530 ( .A(n7930), .ZN(n7682) );
  INV_X1 U7531 ( .A(n7681), .ZN(n5998) );
  NOR2_X1 U7532 ( .A1(n7682), .A2(n5998), .ZN(n5999) );
  NAND2_X1 U7533 ( .A1(n7680), .A2(n5999), .ZN(n6000) );
  NAND2_X1 U7534 ( .A1(n6703), .A2(n5947), .ZN(n6005) );
  INV_X1 U7535 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U7536 ( .A1(n6002), .A2(n6001), .ZN(n6003) );
  NAND2_X1 U7537 ( .A1(n6003), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6015) );
  XNOR2_X1 U7538 ( .A(n6015), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7528) );
  AOI22_X1 U7539 ( .A1(n6217), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6077), .B2(
        n7528), .ZN(n6004) );
  NAND2_X1 U7540 ( .A1(n4378), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6013) );
  NAND2_X1 U7541 ( .A1(n6179), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6012) );
  INV_X1 U7542 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7543 ( .A1(n6008), .A2(n6007), .ZN(n6009) );
  AND2_X1 U7544 ( .A1(n6024), .A2(n6009), .ZN(n7937) );
  NAND2_X1 U7545 ( .A1(n5904), .A2(n7937), .ZN(n6011) );
  NAND2_X1 U7546 ( .A1(n5915), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6010) );
  OR2_X1 U7547 ( .A1(n8722), .A2(n7965), .ZN(n6283) );
  NAND2_X1 U7548 ( .A1(n8722), .A2(n7965), .ZN(n7962) );
  NAND2_X1 U7549 ( .A1(n6283), .A2(n7962), .ZN(n7932) );
  NAND2_X1 U7550 ( .A1(n6740), .A2(n5947), .ZN(n6021) );
  INV_X1 U7551 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U7552 ( .A1(n6015), .A2(n6014), .ZN(n6016) );
  NAND2_X1 U7553 ( .A1(n6016), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6018) );
  INV_X1 U7554 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7555 ( .A1(n6018), .A2(n6017), .ZN(n6032) );
  OR2_X1 U7556 ( .A1(n6018), .A2(n6017), .ZN(n6019) );
  AOI22_X1 U7557 ( .A1(n6217), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6077), .B2(
        n7918), .ZN(n6020) );
  NAND2_X2 U7558 ( .A1(n6021), .A2(n6020), .ZN(n8716) );
  NAND2_X1 U7559 ( .A1(n5915), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6029) );
  NAND2_X1 U7560 ( .A1(n4378), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6028) );
  INV_X1 U7561 ( .A(n6024), .ZN(n6022) );
  NAND2_X1 U7562 ( .A1(n6022), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6036) );
  INV_X1 U7563 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U7564 ( .A1(n6024), .A2(n6023), .ZN(n6025) );
  AND2_X1 U7565 ( .A1(n6036), .A2(n6025), .ZN(n7959) );
  NAND2_X1 U7566 ( .A1(n5904), .A2(n7959), .ZN(n6027) );
  NAND2_X1 U7567 ( .A1(n6179), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6026) );
  NAND2_X1 U7568 ( .A1(n8716), .A2(n7991), .ZN(n6286) );
  INV_X1 U7569 ( .A(n7992), .ZN(n7956) );
  INV_X1 U7570 ( .A(n7962), .ZN(n6030) );
  NOR2_X1 U7571 ( .A1(n7956), .A2(n6030), .ZN(n6031) );
  NAND2_X1 U7572 ( .A1(n6954), .A2(n5947), .ZN(n6035) );
  NAND2_X1 U7573 ( .A1(n6032), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6033) );
  XNOR2_X1 U7574 ( .A(n6033), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8336) );
  AOI22_X1 U7575 ( .A1(n6217), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8336), .B2(
        n6077), .ZN(n6034) );
  NAND2_X1 U7576 ( .A1(n5915), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6041) );
  NAND2_X1 U7577 ( .A1(n4378), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U7578 ( .A1(n6036), .A2(n10068), .ZN(n6037) );
  AND2_X1 U7579 ( .A1(n6049), .A2(n6037), .ZN(n8017) );
  NAND2_X1 U7580 ( .A1(n5904), .A2(n8017), .ZN(n6039) );
  NAND2_X1 U7581 ( .A1(n6179), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6038) );
  NAND2_X1 U7582 ( .A1(n8711), .A2(n8616), .ZN(n6295) );
  NAND2_X1 U7583 ( .A1(n6290), .A2(n6295), .ZN(n7999) );
  INV_X1 U7584 ( .A(n7999), .ZN(n6380) );
  NAND2_X1 U7585 ( .A1(n8000), .A2(n6380), .ZN(n6042) );
  NAND2_X1 U7586 ( .A1(n7004), .A2(n5947), .ZN(n6046) );
  NAND2_X1 U7587 ( .A1(n6043), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6044) );
  XNOR2_X1 U7588 ( .A(n6044), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8342) );
  AOI22_X1 U7589 ( .A1(n6217), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6077), .B2(
        n8342), .ZN(n6045) );
  NAND2_X1 U7590 ( .A1(n4378), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6054) );
  NAND2_X1 U7591 ( .A1(n5915), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6053) );
  INV_X1 U7592 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6048) );
  NAND2_X1 U7593 ( .A1(n6049), .A2(n6048), .ZN(n6050) );
  AND2_X1 U7594 ( .A1(n6060), .A2(n6050), .ZN(n8624) );
  NAND2_X1 U7595 ( .A1(n5904), .A2(n8624), .ZN(n6052) );
  NAND2_X1 U7596 ( .A1(n6179), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6051) );
  OR2_X1 U7597 ( .A1(n8706), .A2(n8262), .ZN(n6296) );
  NAND2_X1 U7598 ( .A1(n8706), .A2(n8262), .ZN(n8588) );
  INV_X1 U7599 ( .A(n8609), .ZN(n8610) );
  NAND2_X1 U7600 ( .A1(n7024), .A2(n5947), .ZN(n6059) );
  OR2_X1 U7601 ( .A1(n6043), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n6055) );
  NAND2_X1 U7602 ( .A1(n6055), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6056) );
  MUX2_X1 U7603 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6056), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n6057) );
  NAND2_X1 U7604 ( .A1(n6057), .A2(n6068), .ZN(n8357) );
  INV_X1 U7605 ( .A(n8357), .ZN(n8366) );
  AOI22_X1 U7606 ( .A1(n6217), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6077), .B2(
        n8366), .ZN(n6058) );
  NAND2_X1 U7607 ( .A1(n5915), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7608 ( .A1(n4378), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7609 ( .A1(n6060), .A2(n8346), .ZN(n6061) );
  AND2_X1 U7610 ( .A1(n6083), .A2(n6061), .ZN(n8599) );
  NAND2_X1 U7611 ( .A1(n5904), .A2(n8599), .ZN(n6063) );
  NAND2_X1 U7612 ( .A1(n6179), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7613 ( .A1(n8703), .A2(n8618), .ZN(n6293) );
  INV_X1 U7614 ( .A(n8588), .ZN(n6066) );
  NOR2_X1 U7615 ( .A1(n8187), .A2(n6066), .ZN(n6067) );
  NAND2_X1 U7616 ( .A1(n7285), .A2(n5947), .ZN(n6071) );
  NAND2_X1 U7617 ( .A1(n6068), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6069) );
  XNOR2_X1 U7618 ( .A(n6069), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8367) );
  AOI22_X1 U7619 ( .A1(n6217), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6077), .B2(
        n8367), .ZN(n6070) );
  XNOR2_X1 U7620 ( .A(n6083), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n8569) );
  NAND2_X1 U7621 ( .A1(n8569), .A2(n5904), .ZN(n6075) );
  NAND2_X1 U7622 ( .A1(n5915), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U7623 ( .A1(n4378), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U7624 ( .A1(n6179), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6072) );
  NAND4_X1 U7625 ( .A1(n6075), .A2(n6074), .A3(n6073), .A4(n6072), .ZN(n8589)
         );
  NAND2_X1 U7626 ( .A1(n8696), .A2(n8554), .ZN(n6309) );
  NAND2_X1 U7627 ( .A1(n8572), .A2(n8564), .ZN(n6076) );
  NAND2_X1 U7628 ( .A1(n7352), .A2(n5947), .ZN(n6079) );
  XNOR2_X1 U7629 ( .A(n6223), .B(n6222), .ZN(n6227) );
  AOI22_X1 U7630 ( .A1(n6217), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6077), .B2(
        n9812), .ZN(n6078) );
  INV_X1 U7631 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n10222) );
  NAND2_X1 U7632 ( .A1(n4378), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U7633 ( .A1(n5915), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6080) );
  AND2_X1 U7634 ( .A1(n6081), .A2(n6080), .ZN(n6088) );
  INV_X1 U7635 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10228) );
  INV_X1 U7636 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6082) );
  OAI21_X1 U7637 ( .B1(n6083), .B2(n10228), .A(n6082), .ZN(n6086) );
  AND2_X1 U7638 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n6084) );
  NAND2_X1 U7639 ( .A1(n6086), .A2(n6092), .ZN(n8244) );
  OR2_X1 U7640 ( .A1(n8244), .A2(n6160), .ZN(n6087) );
  OAI211_X1 U7641 ( .C1(n6194), .C2(n10222), .A(n6088), .B(n6087), .ZN(n8575)
         );
  INV_X1 U7642 ( .A(n8575), .ZN(n8291) );
  OR2_X1 U7643 ( .A1(n8693), .A2(n8291), .ZN(n6310) );
  NAND2_X1 U7644 ( .A1(n8693), .A2(n8291), .ZN(n8531) );
  NAND2_X1 U7645 ( .A1(n6310), .A2(n8531), .ZN(n8551) );
  NAND2_X1 U7646 ( .A1(n9955), .A2(n5947), .ZN(n6091) );
  OR2_X1 U7647 ( .A1(n5901), .A2(n6089), .ZN(n6090) );
  INV_X1 U7648 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8106) );
  NAND2_X1 U7649 ( .A1(n6092), .A2(n8106), .ZN(n6093) );
  AND2_X1 U7650 ( .A1(n6100), .A2(n6093), .ZN(n8543) );
  NAND2_X1 U7651 ( .A1(n8543), .A2(n5904), .ZN(n6096) );
  AOI22_X1 U7652 ( .A1(n6179), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n4378), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U7653 ( .A1(n5915), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U7654 ( .A1(n8686), .A2(n8555), .ZN(n6313) );
  INV_X1 U7655 ( .A(n8539), .ZN(n8190) );
  INV_X1 U7656 ( .A(n8531), .ZN(n6300) );
  NAND2_X1 U7657 ( .A1(n7553), .A2(n5947), .ZN(n6098) );
  OR2_X1 U7658 ( .A1(n5901), .A2(n10066), .ZN(n6097) );
  INV_X1 U7659 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8099) );
  NAND2_X1 U7660 ( .A1(n6100), .A2(n8099), .ZN(n6101) );
  NAND2_X1 U7661 ( .A1(n6112), .A2(n6101), .ZN(n8518) );
  OR2_X1 U7662 ( .A1(n8518), .A2(n6160), .ZN(n6108) );
  INV_X1 U7663 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U7664 ( .A1(n5915), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7665 ( .A1(n6179), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6102) );
  OAI211_X1 U7666 ( .C1(n10279), .C2(n6104), .A(n6103), .B(n6102), .ZN(n6106)
         );
  INV_X1 U7667 ( .A(n6106), .ZN(n6107) );
  NAND2_X1 U7668 ( .A1(n6108), .A2(n6107), .ZN(n8533) );
  INV_X1 U7669 ( .A(n8533), .ZN(n8507) );
  OR2_X1 U7670 ( .A1(n8679), .A2(n8507), .ZN(n6315) );
  NAND2_X1 U7671 ( .A1(n8679), .A2(n8507), .ZN(n8504) );
  NAND2_X1 U7672 ( .A1(n7649), .A2(n5947), .ZN(n6110) );
  OR2_X1 U7673 ( .A1(n5901), .A2(n7651), .ZN(n6109) );
  INV_X1 U7674 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U7675 ( .A1(n6112), .A2(n6111), .ZN(n6113) );
  AND2_X1 U7676 ( .A1(n6124), .A2(n6113), .ZN(n8500) );
  NAND2_X1 U7677 ( .A1(n8500), .A2(n5904), .ZN(n6118) );
  INV_X1 U7678 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n10128) );
  NAND2_X1 U7679 ( .A1(n4378), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U7680 ( .A1(n5915), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6114) );
  OAI211_X1 U7681 ( .C1(n6194), .C2(n10128), .A(n6115), .B(n6114), .ZN(n6116)
         );
  INV_X1 U7682 ( .A(n6116), .ZN(n6117) );
  NAND2_X1 U7683 ( .A1(n8674), .A2(n8229), .ZN(n6318) );
  INV_X1 U7684 ( .A(n8504), .ZN(n6119) );
  NOR2_X1 U7685 ( .A1(n8498), .A2(n6119), .ZN(n6120) );
  NAND2_X1 U7686 ( .A1(n8522), .A2(n6120), .ZN(n8487) );
  NAND2_X1 U7687 ( .A1(n7725), .A2(n5947), .ZN(n6122) );
  OR2_X1 U7688 ( .A1(n5901), .A2(n7729), .ZN(n6121) );
  INV_X1 U7689 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8228) );
  NAND2_X1 U7690 ( .A1(n6124), .A2(n8228), .ZN(n6125) );
  NAND2_X1 U7691 ( .A1(n6135), .A2(n6125), .ZN(n8483) );
  OR2_X1 U7692 ( .A1(n8483), .A2(n6160), .ZN(n6130) );
  INV_X1 U7693 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n10072) );
  NAND2_X1 U7694 ( .A1(n5915), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U7695 ( .A1(n4378), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6126) );
  OAI211_X1 U7696 ( .C1(n10072), .C2(n6194), .A(n6127), .B(n6126), .ZN(n6128)
         );
  INV_X1 U7697 ( .A(n6128), .ZN(n6129) );
  NAND2_X1 U7698 ( .A1(n6130), .A2(n6129), .ZN(n8313) );
  NAND2_X1 U7699 ( .A1(n8486), .A2(n8313), .ZN(n6230) );
  INV_X1 U7700 ( .A(n8313), .ZN(n8508) );
  NAND2_X1 U7701 ( .A1(n8669), .A2(n8508), .ZN(n6323) );
  INV_X1 U7702 ( .A(n6304), .ZN(n8489) );
  NOR2_X1 U7703 ( .A1(n8488), .A2(n8489), .ZN(n6131) );
  NAND2_X1 U7704 ( .A1(n8487), .A2(n6131), .ZN(n8490) );
  NAND2_X1 U7705 ( .A1(n8490), .A2(n6323), .ZN(n8461) );
  NAND2_X1 U7706 ( .A1(n7834), .A2(n5947), .ZN(n6133) );
  OR2_X1 U7707 ( .A1(n5901), .A2(n7835), .ZN(n6132) );
  INV_X1 U7708 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6134) );
  NAND2_X1 U7709 ( .A1(n6135), .A2(n6134), .ZN(n6136) );
  NAND2_X1 U7710 ( .A1(n6147), .A2(n6136), .ZN(n8470) );
  OR2_X1 U7711 ( .A1(n8470), .A2(n6160), .ZN(n6142) );
  INV_X1 U7712 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n6139) );
  NAND2_X1 U7713 ( .A1(n5915), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U7714 ( .A1(n4378), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6137) );
  OAI211_X1 U7715 ( .C1(n6139), .C2(n6194), .A(n6138), .B(n6137), .ZN(n6140)
         );
  INV_X1 U7716 ( .A(n6140), .ZN(n6141) );
  NAND2_X1 U7717 ( .A1(n8662), .A2(n8254), .ZN(n6325) );
  NAND2_X1 U7718 ( .A1(n6228), .A2(n6325), .ZN(n8460) );
  NAND2_X1 U7719 ( .A1(n7943), .A2(n5947), .ZN(n6145) );
  OR2_X1 U7720 ( .A1(n5901), .A2(n10086), .ZN(n6144) );
  INV_X1 U7721 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6146) );
  NAND2_X1 U7722 ( .A1(n6147), .A2(n6146), .ZN(n6148) );
  NAND2_X1 U7723 ( .A1(n6158), .A2(n6148), .ZN(n8257) );
  INV_X1 U7724 ( .A(n8257), .ZN(n8448) );
  INV_X1 U7725 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7726 ( .A1(n5915), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U7727 ( .A1(n4378), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6149) );
  OAI211_X1 U7728 ( .C1(n6151), .C2(n6194), .A(n6150), .B(n6149), .ZN(n6152)
         );
  AOI21_X1 U7729 ( .B1(n8448), .B2(n5904), .A(n6152), .ZN(n8303) );
  OR2_X1 U7730 ( .A1(n8657), .A2(n8303), .ZN(n6327) );
  NAND2_X1 U7731 ( .A1(n8657), .A2(n8303), .ZN(n6328) );
  NAND2_X1 U7732 ( .A1(n6327), .A2(n6328), .ZN(n8451) );
  INV_X1 U7733 ( .A(n8451), .ZN(n6153) );
  NAND2_X1 U7734 ( .A1(n7972), .A2(n5947), .ZN(n6156) );
  OR2_X1 U7735 ( .A1(n5901), .A2(n7977), .ZN(n6155) );
  INV_X1 U7736 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10169) );
  NAND2_X1 U7737 ( .A1(n6158), .A2(n10169), .ZN(n6159) );
  NAND2_X1 U7738 ( .A1(n6177), .A2(n6159), .ZN(n8438) );
  INV_X1 U7739 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U7740 ( .A1(n5915), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U7741 ( .A1(n4378), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6161) );
  OAI211_X1 U7742 ( .C1(n6163), .C2(n6194), .A(n6162), .B(n6161), .ZN(n6164)
         );
  INV_X1 U7743 ( .A(n6164), .ZN(n6165) );
  OR2_X1 U7744 ( .A1(n8652), .A2(n8255), .ZN(n6331) );
  NAND2_X1 U7745 ( .A1(n8652), .A2(n8255), .ZN(n6332) );
  NAND2_X1 U7746 ( .A1(n6331), .A2(n6332), .ZN(n8429) );
  NAND2_X1 U7747 ( .A1(n7989), .A2(n5947), .ZN(n6169) );
  OR2_X1 U7748 ( .A1(n5901), .A2(n8006), .ZN(n6168) );
  XNOR2_X1 U7749 ( .A(n6177), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8418) );
  INV_X1 U7750 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n10129) );
  NAND2_X1 U7751 ( .A1(n6179), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U7752 ( .A1(n4378), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6170) );
  OAI211_X1 U7753 ( .C1(n6172), .C2(n10129), .A(n6171), .B(n6170), .ZN(n6173)
         );
  AOI21_X1 U7754 ( .B1(n8418), .B2(n5904), .A(n6173), .ZN(n8305) );
  XNOR2_X1 U7755 ( .A(n8646), .B(n8305), .ZN(n8421) );
  OR2_X1 U7756 ( .A1(n8646), .A2(n8305), .ZN(n6336) );
  NAND2_X1 U7757 ( .A1(n8007), .A2(n5947), .ZN(n6175) );
  OR2_X1 U7758 ( .A1(n5901), .A2(n10144), .ZN(n6174) );
  INV_X1 U7759 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8157) );
  INV_X1 U7760 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6176) );
  OAI21_X1 U7761 ( .B1(n6177), .B2(n8157), .A(n6176), .ZN(n6178) );
  INV_X1 U7762 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n10088) );
  NAND2_X1 U7763 ( .A1(n6179), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6181) );
  NAND2_X1 U7764 ( .A1(n4378), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6180) );
  OAI211_X1 U7765 ( .C1(n6172), .C2(n10088), .A(n6181), .B(n6180), .ZN(n6182)
         );
  NAND2_X1 U7766 ( .A1(n8641), .A2(n8202), .ZN(n6343) );
  INV_X1 U7767 ( .A(n8405), .ZN(n6386) );
  INV_X1 U7768 ( .A(SI_28_), .ZN(n6185) );
  MUX2_X1 U7769 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n5634), .Z(n6198) );
  INV_X1 U7770 ( .A(SI_29_), .ZN(n6187) );
  XNOR2_X1 U7771 ( .A(n6198), .B(n6187), .ZN(n6188) );
  NAND2_X1 U7772 ( .A1(n8883), .A2(n5947), .ZN(n6190) );
  INV_X1 U7773 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8745) );
  OR2_X1 U7774 ( .A1(n5901), .A2(n8745), .ZN(n6189) );
  INV_X1 U7775 ( .A(n6191), .ZN(n8206) );
  INV_X1 U7776 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U7777 ( .A1(n4378), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6193) );
  NAND2_X1 U7778 ( .A1(n5915), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6192) );
  OAI211_X1 U7779 ( .C1(n6195), .C2(n6194), .A(n6193), .B(n6192), .ZN(n6196)
         );
  AOI21_X1 U7780 ( .B1(n8206), .B2(n5904), .A(n6196), .ZN(n8168) );
  NAND2_X1 U7781 ( .A1(n8636), .A2(n8168), .ZN(n6350) );
  INV_X1 U7782 ( .A(n6350), .ZN(n6197) );
  AOI21_X1 U7783 ( .B1(n8209), .B2(n8204), .A(n6197), .ZN(n6204) );
  AOI21_X1 U7784 ( .B1(n8311), .B2(n6203), .A(n6204), .ZN(n6207) );
  NOR2_X1 U7785 ( .A1(n6198), .A2(SI_29_), .ZN(n6200) );
  NAND2_X1 U7786 ( .A1(n6198), .A2(SI_29_), .ZN(n6199) );
  MUX2_X1 U7787 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n5634), .Z(n6210) );
  INV_X1 U7788 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8179) );
  OR2_X1 U7789 ( .A1(n5901), .A2(n8179), .ZN(n6202) );
  INV_X1 U7790 ( .A(n6203), .ZN(n6206) );
  INV_X1 U7791 ( .A(n6204), .ZN(n6205) );
  OAI22_X1 U7792 ( .A1(n6207), .A2(n9557), .B1(n6206), .B2(n6205), .ZN(n6218)
         );
  INV_X1 U7793 ( .A(n6208), .ZN(n6209) );
  NAND2_X1 U7794 ( .A1(n6209), .A2(SI_30_), .ZN(n6213) );
  NAND2_X1 U7795 ( .A1(n6211), .A2(n6210), .ZN(n6212) );
  NAND2_X1 U7796 ( .A1(n6213), .A2(n6212), .ZN(n6216) );
  MUX2_X1 U7797 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n5634), .Z(n6214) );
  XNOR2_X1 U7798 ( .A(n6214), .B(SI_31_), .ZN(n6215) );
  INV_X1 U7799 ( .A(n6361), .ZN(n8390) );
  NOR2_X1 U7800 ( .A1(n6359), .A2(n8390), .ZN(n6356) );
  NAND2_X1 U7801 ( .A1(n6223), .A2(n6222), .ZN(n6224) );
  NAND2_X1 U7802 ( .A1(n6224), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6226) );
  INV_X1 U7803 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6225) );
  INV_X1 U7804 ( .A(n7010), .ZN(n9953) );
  NAND2_X1 U7805 ( .A1(n7581), .A2(n9953), .ZN(n6824) );
  INV_X1 U7806 ( .A(n6228), .ZN(n6326) );
  NAND2_X1 U7807 ( .A1(n7581), .A2(n9812), .ZN(n6229) );
  INV_X1 U7808 ( .A(n6230), .ZN(n6231) );
  NOR2_X1 U7809 ( .A1(n8460), .A2(n6231), .ZN(n6322) );
  AND2_X1 U7810 ( .A1(n6366), .A2(n6370), .ZN(n6232) );
  INV_X1 U7811 ( .A(n6360), .ZN(n6345) );
  MUX2_X1 U7812 ( .A(n6235), .B(n6232), .S(n6345), .Z(n6246) );
  INV_X1 U7813 ( .A(n6246), .ZN(n6233) );
  NAND2_X1 U7814 ( .A1(n6233), .A2(n6369), .ZN(n6238) );
  NAND2_X1 U7815 ( .A1(n6235), .A2(n6234), .ZN(n6237) );
  INV_X1 U7816 ( .A(n6254), .ZN(n6236) );
  AOI21_X1 U7817 ( .B1(n6238), .B2(n6237), .A(n6236), .ZN(n6257) );
  NAND2_X1 U7818 ( .A1(n6366), .A2(n6239), .ZN(n6241) );
  NAND2_X1 U7819 ( .A1(n6370), .A2(n6259), .ZN(n6240) );
  AOI21_X1 U7820 ( .B1(n6246), .B2(n6241), .A(n6240), .ZN(n6248) );
  INV_X1 U7821 ( .A(n9847), .ZN(n7034) );
  NAND2_X1 U7822 ( .A1(n6895), .A2(n7034), .ZN(n7030) );
  AND2_X1 U7823 ( .A1(n7030), .A2(n7581), .ZN(n6242) );
  OAI211_X1 U7824 ( .C1(n6243), .C2(n6242), .A(n6251), .B(n6365), .ZN(n6244)
         );
  NAND3_X1 U7825 ( .A1(n6244), .A2(n6360), .A3(n6250), .ZN(n6245) );
  NAND3_X1 U7826 ( .A1(n6246), .A2(n6367), .A3(n6245), .ZN(n6247) );
  OAI21_X1 U7827 ( .B1(n6248), .B2(n6345), .A(n6247), .ZN(n6255) );
  NAND2_X1 U7828 ( .A1(n7030), .A2(n6365), .ZN(n6249) );
  NAND3_X1 U7829 ( .A1(n6364), .A2(n6250), .A3(n6249), .ZN(n6252) );
  NAND3_X1 U7830 ( .A1(n6252), .A2(n6345), .A3(n6251), .ZN(n6253) );
  NAND3_X1 U7831 ( .A1(n6255), .A2(n6254), .A3(n6253), .ZN(n6256) );
  OAI21_X1 U7832 ( .B1(n6257), .B2(n6360), .A(n6256), .ZN(n6258) );
  OAI211_X1 U7833 ( .C1(n6259), .C2(n6360), .A(n6258), .B(n7385), .ZN(n6263)
         );
  MUX2_X1 U7834 ( .A(n6261), .B(n6260), .S(n6360), .Z(n6262) );
  MUX2_X1 U7835 ( .A(n6265), .B(n6264), .S(n6345), .Z(n6266) );
  AND2_X1 U7836 ( .A1(n6372), .A2(n6374), .ZN(n6268) );
  AND2_X1 U7837 ( .A1(n6373), .A2(n6375), .ZN(n6267) );
  MUX2_X1 U7838 ( .A(n6268), .B(n6267), .S(n6345), .Z(n6273) );
  NAND2_X1 U7839 ( .A1(n7681), .A2(n6372), .ZN(n6271) );
  INV_X1 U7840 ( .A(n6372), .ZN(n6269) );
  OAI211_X1 U7841 ( .C1(n6269), .C2(n6375), .A(n6274), .B(n6373), .ZN(n6270)
         );
  MUX2_X1 U7842 ( .A(n6271), .B(n6270), .S(n6360), .Z(n6272) );
  NAND2_X1 U7843 ( .A1(n6277), .A2(n7681), .ZN(n6276) );
  NAND2_X1 U7844 ( .A1(n6278), .A2(n6274), .ZN(n6275) );
  MUX2_X1 U7845 ( .A(n6276), .B(n6275), .S(n6345), .Z(n6282) );
  NOR2_X1 U7846 ( .A1(n6277), .A2(n6360), .ZN(n6279) );
  MUX2_X1 U7847 ( .A(n6360), .B(n6279), .S(n6278), .Z(n6280) );
  NOR2_X1 U7848 ( .A1(n7932), .A2(n6280), .ZN(n6281) );
  NAND2_X1 U7849 ( .A1(n6287), .A2(n6283), .ZN(n6285) );
  NAND2_X1 U7850 ( .A1(n6286), .A2(n7962), .ZN(n6284) );
  MUX2_X1 U7851 ( .A(n6285), .B(n6284), .S(n6360), .Z(n6289) );
  MUX2_X1 U7852 ( .A(n6287), .B(n6286), .S(n6345), .Z(n6288) );
  OAI211_X1 U7853 ( .C1(n4418), .C2(n6289), .A(n6380), .B(n6288), .ZN(n6294)
         );
  NAND3_X1 U7854 ( .A1(n8609), .A2(n6290), .A3(n6294), .ZN(n6291) );
  NAND2_X1 U7855 ( .A1(n6291), .A2(n8588), .ZN(n6292) );
  NAND3_X1 U7856 ( .A1(n8609), .A2(n6295), .A3(n6294), .ZN(n6297) );
  INV_X1 U7857 ( .A(n6301), .ZN(n6299) );
  AOI21_X1 U7858 ( .B1(n6308), .B2(n6301), .A(n6300), .ZN(n6303) );
  NAND2_X1 U7859 ( .A1(n6316), .A2(n6310), .ZN(n6302) );
  OAI211_X1 U7860 ( .C1(n6303), .C2(n6302), .A(n8504), .B(n6313), .ZN(n6305)
         );
  NAND3_X1 U7861 ( .A1(n6305), .A2(n6304), .A3(n6315), .ZN(n6306) );
  NAND2_X1 U7862 ( .A1(n6306), .A2(n6318), .ZN(n6307) );
  INV_X1 U7863 ( .A(n6308), .ZN(n6312) );
  INV_X1 U7864 ( .A(n6309), .ZN(n6311) );
  OAI21_X1 U7865 ( .B1(n6312), .B2(n6311), .A(n6310), .ZN(n6314) );
  NAND3_X1 U7866 ( .A1(n6314), .A2(n8531), .A3(n6313), .ZN(n6317) );
  NAND3_X1 U7867 ( .A1(n6317), .A2(n6316), .A3(n6315), .ZN(n6319) );
  NAND4_X1 U7868 ( .A1(n6319), .A2(n6360), .A3(n6318), .A4(n8504), .ZN(n6320)
         );
  NAND2_X1 U7869 ( .A1(n8197), .A2(n6320), .ZN(n6321) );
  NAND2_X1 U7870 ( .A1(n6325), .A2(n6323), .ZN(n6324) );
  NAND2_X1 U7871 ( .A1(n6331), .A2(n6327), .ZN(n6330) );
  NAND2_X1 U7872 ( .A1(n6332), .A2(n6328), .ZN(n6329) );
  MUX2_X1 U7873 ( .A(n6330), .B(n6329), .S(n6360), .Z(n6334) );
  MUX2_X1 U7874 ( .A(n6332), .B(n6331), .S(n6360), .Z(n6333) );
  INV_X1 U7875 ( .A(n8421), .ZN(n6384) );
  OAI211_X1 U7876 ( .C1(n6335), .C2(n6334), .A(n6333), .B(n6384), .ZN(n6341)
         );
  AND2_X1 U7877 ( .A1(n6337), .A2(n6336), .ZN(n6339) );
  NAND2_X1 U7878 ( .A1(n8646), .A2(n8305), .ZN(n6338) );
  MUX2_X1 U7879 ( .A(n6339), .B(n6338), .S(n6360), .Z(n6340) );
  NAND3_X1 U7880 ( .A1(n6341), .A2(n6340), .A3(n6343), .ZN(n6344) );
  AOI21_X1 U7881 ( .B1(n6344), .B2(n8202), .A(n8210), .ZN(n6348) );
  INV_X1 U7882 ( .A(n6349), .ZN(n6342) );
  NOR2_X1 U7883 ( .A1(n6342), .A2(n6360), .ZN(n6347) );
  OAI211_X1 U7884 ( .C1(n6345), .C2(n8641), .A(n6344), .B(n6343), .ZN(n6346)
         );
  OAI21_X1 U7885 ( .B1(n6348), .B2(n6347), .A(n6346), .ZN(n6354) );
  MUX2_X1 U7886 ( .A(n6350), .B(n6349), .S(n6360), .Z(n6353) );
  NAND2_X1 U7887 ( .A1(n8395), .A2(n8311), .ZN(n6357) );
  INV_X1 U7888 ( .A(n6357), .ZN(n6352) );
  AOI211_X1 U7889 ( .C1(n6354), .C2(n6353), .A(n6352), .B(n6351), .ZN(n6363)
         );
  INV_X1 U7890 ( .A(n6356), .ZN(n6358) );
  MUX2_X1 U7891 ( .A(n6359), .B(n6361), .S(n6360), .Z(n6362) );
  INV_X1 U7892 ( .A(n8564), .ZN(n8573) );
  NAND2_X1 U7893 ( .A1(n7032), .A2(n7030), .ZN(n9848) );
  NAND2_X1 U7894 ( .A1(n6365), .A2(n6364), .ZN(n6833) );
  NOR4_X1 U7895 ( .A1(n6882), .A2(n9848), .A3(n6893), .A4(n7010), .ZN(n6368)
         );
  NAND2_X1 U7896 ( .A1(n6366), .A2(n7258), .ZN(n6838) );
  INV_X1 U7897 ( .A(n6838), .ZN(n6823) );
  NAND3_X1 U7898 ( .A1(n6368), .A2(n6367), .A3(n6823), .ZN(n6371) );
  INV_X1 U7899 ( .A(n7385), .ZN(n7180) );
  NAND2_X1 U7900 ( .A1(n6370), .A2(n6369), .ZN(n7260) );
  NOR4_X1 U7901 ( .A1(n6371), .A2(n7180), .A3(n7175), .A4(n7260), .ZN(n6377)
         );
  NAND2_X1 U7902 ( .A1(n6373), .A2(n6372), .ZN(n7636) );
  INV_X1 U7903 ( .A(n7636), .ZN(n6376) );
  NAND4_X1 U7904 ( .A1(n6377), .A2(n7391), .A3(n6376), .A4(n7710), .ZN(n6378)
         );
  NOR4_X1 U7905 ( .A1(n7932), .A2(n7682), .A3(n7745), .A4(n6378), .ZN(n6379)
         );
  NAND4_X1 U7906 ( .A1(n8609), .A2(n6380), .A3(n7992), .A4(n6379), .ZN(n6381)
         );
  NOR4_X1 U7907 ( .A1(n8551), .A2(n8573), .A3(n8187), .A4(n6381), .ZN(n6382)
         );
  NAND4_X1 U7908 ( .A1(n8197), .A2(n8539), .A3(n8523), .A4(n6382), .ZN(n6383)
         );
  NOR4_X1 U7909 ( .A1(n8451), .A2(n8460), .A3(n8498), .A4(n6383), .ZN(n6385)
         );
  NAND4_X1 U7910 ( .A1(n6386), .A2(n6167), .A3(n6385), .A4(n6384), .ZN(n6387)
         );
  XNOR2_X1 U7911 ( .A(n6390), .B(n9812), .ZN(n6391) );
  AOI211_X1 U7912 ( .C1(n7010), .C2(n6395), .A(n7581), .B(n6391), .ZN(n6392)
         );
  INV_X1 U7913 ( .A(n6392), .ZN(n6397) );
  INV_X1 U7914 ( .A(n6825), .ZN(n6396) );
  NAND2_X1 U7915 ( .A1(n6399), .A2(n6398), .ZN(n6400) );
  XNOR2_X1 U7916 ( .A(n6410), .B(n6409), .ZN(n6866) );
  OR2_X1 U7917 ( .A1(n6866), .A2(P2_U3152), .ZN(n7726) );
  INV_X1 U7918 ( .A(n6401), .ZN(n6402) );
  OAI21_X1 U7919 ( .B1(n6403), .B2(n6402), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6404) );
  MUX2_X1 U7920 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6404), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6406) );
  NAND2_X1 U7921 ( .A1(n6406), .A2(n6405), .ZN(n7945) );
  INV_X1 U7922 ( .A(n7945), .ZN(n6408) );
  NAND2_X1 U7923 ( .A1(n6405), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6407) );
  NAND2_X1 U7924 ( .A1(n6408), .A2(n6806), .ZN(n6414) );
  NAND2_X1 U7925 ( .A1(n6410), .A2(n6409), .ZN(n6411) );
  NAND2_X1 U7926 ( .A1(n6411), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6413) );
  NAND2_X1 U7927 ( .A1(n6866), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9844) );
  INV_X1 U7928 ( .A(n9844), .ZN(n6415) );
  INV_X1 U7929 ( .A(n6416), .ZN(n6826) );
  AND2_X1 U7930 ( .A1(n6862), .A2(n6873), .ZN(n6868) );
  NOR4_X1 U7931 ( .A1(n9819), .A2(n8615), .A3(n6868), .A4(n8212), .ZN(n6418)
         );
  OAI21_X1 U7932 ( .B1(n7726), .B2(n6393), .A(P2_B_REG_SCAN_IN), .ZN(n6417) );
  OAI21_X1 U7933 ( .B1(n6420), .B2(n7726), .A(n6419), .ZN(P2_U3244) );
  AOI21_X1 U7934 ( .B1(n6422), .B2(n6421), .A(n8874), .ZN(n6423) );
  INV_X1 U7935 ( .A(n6424), .ZN(n9279) );
  AOI22_X1 U7936 ( .A1(n9279), .A2(n8819), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n6426) );
  NAND2_X1 U7937 ( .A1(n9288), .A2(n8868), .ZN(n6425) );
  OAI211_X1 U7938 ( .C1(n9229), .C2(n8865), .A(n6426), .B(n6425), .ZN(n6427)
         );
  AOI21_X1 U7939 ( .B1(n9465), .B2(n8872), .A(n6427), .ZN(n6428) );
  INV_X1 U7940 ( .A(n6431), .ZN(n7722) );
  NOR2_X1 U7941 ( .A1(n6430), .A2(n7722), .ZN(n6690) );
  NAND2_X1 U7942 ( .A1(n6997), .A2(n6430), .ZN(n6432) );
  NAND2_X1 U7943 ( .A1(n6432), .A2(n6431), .ZN(n9206) );
  NAND2_X1 U7944 ( .A1(n9206), .A2(n5069), .ZN(n9590) );
  NAND2_X1 U7945 ( .A1(n9590), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X2 U7946 ( .A(n8314), .ZN(P2_U3966) );
  AND2_X1 U7947 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7773) );
  INV_X1 U7948 ( .A(n9650), .ZN(n6490) );
  AOI22_X1 U7949 ( .A1(n9650), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7415), .B2(
        n6490), .ZN(n9642) );
  INV_X1 U7950 ( .A(n6501), .ZN(n6486) );
  AOI22_X1 U7951 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6501), .B1(n6486), .B2(
        n5169), .ZN(n6494) );
  INV_X1 U7952 ( .A(n9635), .ZN(n6451) );
  INV_X1 U7953 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6433) );
  MUX2_X1 U7954 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6433), .S(n9635), .Z(n9631)
         );
  NOR2_X1 U7955 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n9618), .ZN(n6434) );
  AOI21_X1 U7956 ( .B1(n9618), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6434), .ZN(
        n9620) );
  MUX2_X1 U7957 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n7002), .S(n6463), .Z(n6513)
         );
  NAND2_X1 U7958 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6686) );
  INV_X1 U7959 ( .A(n6686), .ZN(n6512) );
  NAND2_X1 U7960 ( .A1(n6513), .A2(n6512), .ZN(n6511) );
  NAND2_X1 U7961 ( .A1(n6463), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6435) );
  NAND2_X1 U7962 ( .A1(n6511), .A2(n6435), .ZN(n6694) );
  XNOR2_X1 U7963 ( .A(n6692), .B(n9961), .ZN(n6695) );
  NAND2_X1 U7964 ( .A1(n6692), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6436) );
  XNOR2_X1 U7965 ( .A(n9603), .B(n7438), .ZN(n9601) );
  NAND2_X1 U7966 ( .A1(n9600), .A2(n9601), .ZN(n9599) );
  OAI21_X1 U7967 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n9603), .A(n9599), .ZN(
        n9621) );
  NAND2_X1 U7968 ( .A1(n9620), .A2(n9621), .ZN(n9619) );
  OAI21_X1 U7969 ( .B1(n9618), .B2(P1_REG2_REG_5__SCAN_IN), .A(n9619), .ZN(
        n9630) );
  NOR2_X1 U7970 ( .A1(n9631), .A2(n9630), .ZN(n9629) );
  AOI21_X1 U7971 ( .B1(n6451), .B2(P1_REG2_REG_6__SCAN_IN), .A(n9629), .ZN(
        n6495) );
  NAND2_X1 U7972 ( .A1(n6494), .A2(n6495), .ZN(n6493) );
  OAI21_X1 U7973 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6501), .A(n6493), .ZN(
        n9641) );
  NAND2_X1 U7974 ( .A1(n6731), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6437) );
  OAI21_X1 U7975 ( .B1(n6731), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6437), .ZN(
        n6440) );
  NOR2_X1 U7976 ( .A1(n6688), .A2(P1_U3084), .ZN(n9207) );
  INV_X1 U7977 ( .A(n9207), .ZN(n6438) );
  NOR2_X1 U7978 ( .A1(n6438), .A2(n5798), .ZN(n6439) );
  NAND2_X1 U7979 ( .A1(n9206), .A2(n6439), .ZN(n9741) );
  AOI211_X1 U7980 ( .C1(n6441), .C2(n6440), .A(n6730), .B(n9741), .ZN(n6460)
         );
  NAND2_X1 U7981 ( .A1(n9650), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6453) );
  OR2_X1 U7982 ( .A1(n6501), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6452) );
  NOR2_X1 U7983 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6501), .ZN(n6442) );
  AOI21_X1 U7984 ( .B1(n6501), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6442), .ZN(
        n6498) );
  INV_X1 U7985 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6443) );
  MUX2_X1 U7986 ( .A(n6443), .B(P1_REG1_REG_6__SCAN_IN), .S(n9635), .Z(n9627)
         );
  INV_X1 U7987 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10041) );
  MUX2_X1 U7988 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10041), .S(n6692), .Z(n6698)
         );
  INV_X1 U7989 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10155) );
  MUX2_X1 U7990 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10155), .S(n6463), .Z(n6516)
         );
  AND2_X1 U7991 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6515) );
  NAND2_X1 U7992 ( .A1(n6516), .A2(n6515), .ZN(n6514) );
  NAND2_X1 U7993 ( .A1(n6463), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6444) );
  NAND2_X1 U7994 ( .A1(n6514), .A2(n6444), .ZN(n6697) );
  NAND2_X1 U7995 ( .A1(n6698), .A2(n6697), .ZN(n6696) );
  NAND2_X1 U7996 ( .A1(n6692), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6445) );
  NAND2_X1 U7997 ( .A1(n6696), .A2(n6445), .ZN(n8051) );
  INV_X1 U7998 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6446) );
  XNOR2_X1 U7999 ( .A(n8061), .B(n6446), .ZN(n8052) );
  NAND2_X1 U8000 ( .A1(n8051), .A2(n8052), .ZN(n8050) );
  NAND2_X1 U8001 ( .A1(n8061), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6447) );
  NAND2_X1 U8002 ( .A1(n8050), .A2(n6447), .ZN(n9606) );
  INV_X1 U8003 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10106) );
  MUX2_X1 U8004 ( .A(n10106), .B(P1_REG1_REG_4__SCAN_IN), .S(n9603), .Z(n9605)
         );
  NOR2_X1 U8005 ( .A1(n9606), .A2(n9605), .ZN(n9604) );
  NOR2_X1 U8006 ( .A1(n9603), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6448) );
  OR2_X1 U8007 ( .A1(n9604), .A2(n6448), .ZN(n9615) );
  OR2_X1 U8008 ( .A1(n9618), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6450) );
  NAND2_X1 U8009 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n9618), .ZN(n6449) );
  NAND2_X1 U8010 ( .A1(n6450), .A2(n6449), .ZN(n9614) );
  NOR2_X1 U8011 ( .A1(n9615), .A2(n9614), .ZN(n9613) );
  AOI21_X1 U8012 ( .B1(n9618), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9613), .ZN(
        n9628) );
  NAND2_X1 U8013 ( .A1(n9627), .A2(n9628), .ZN(n9626) );
  OAI21_X1 U8014 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n6451), .A(n9626), .ZN(
        n6497) );
  NAND2_X1 U8015 ( .A1(n6498), .A2(n6497), .ZN(n6496) );
  NAND2_X1 U8016 ( .A1(n6452), .A2(n6496), .ZN(n9648) );
  NOR2_X1 U8017 ( .A1(n9650), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9644) );
  AOI21_X1 U8018 ( .B1(n6453), .B2(n9648), .A(n9644), .ZN(n9643) );
  INV_X1 U8019 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9788) );
  AOI22_X1 U8020 ( .A1(n6731), .A2(n9788), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6506), .ZN(n6454) );
  NOR2_X1 U8021 ( .A1(n9643), .A2(n6454), .ZN(n6726) );
  AOI21_X1 U8022 ( .B1(n9643), .B2(n6454), .A(n6726), .ZN(n6456) );
  NOR2_X1 U8023 ( .A1(n5798), .A2(P1_U3084), .ZN(n8008) );
  AND2_X1 U8024 ( .A1(n6688), .A2(n8008), .ZN(n6455) );
  NAND2_X1 U8025 ( .A1(n9206), .A2(n6455), .ZN(n9751) );
  NOR2_X1 U8026 ( .A1(n6456), .A2(n9751), .ZN(n6459) );
  INV_X1 U8027 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10264) );
  AND2_X1 U8028 ( .A1(n5798), .A2(n9207), .ZN(n6457) );
  NAND2_X1 U8029 ( .A1(n9206), .A2(n6457), .ZN(n9745) );
  OAI22_X1 U8030 ( .A1(n9754), .A2(n10264), .B1(n6506), .B2(n9745), .ZN(n6458)
         );
  OR4_X1 U8031 ( .A1(n7773), .A2(n6460), .A3(n6459), .A4(n6458), .ZN(P1_U3250)
         );
  NOR2_X1 U8032 ( .A1(n5634), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9548) );
  AOI22_X1 U8033 ( .A1(n9548), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n6692), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6461) );
  OAI21_X1 U8034 ( .B1(n6476), .B2(n9550), .A(n6461), .ZN(P1_U3351) );
  AOI22_X1 U8035 ( .A1(n9603), .A2(P1_STATE_REG_SCAN_IN), .B1(n9548), .B2(
        P2_DATAO_REG_4__SCAN_IN), .ZN(n6462) );
  OAI21_X1 U8036 ( .B1(n6482), .B2(n9550), .A(n6462), .ZN(P1_U3349) );
  INV_X1 U8037 ( .A(n6463), .ZN(n6510) );
  INV_X1 U8038 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6464) );
  OAI222_X1 U8039 ( .A1(n6510), .A2(P1_U3084), .B1(n9550), .B2(n6467), .C1(
        n6464), .C2(n8222), .ZN(P1_U3352) );
  AOI22_X1 U8040 ( .A1(n9618), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9548), .ZN(n6465) );
  OAI21_X1 U8041 ( .B1(n6478), .B2(n9550), .A(n6465), .ZN(P1_U3348) );
  AND2_X1 U8042 ( .A1(n5634), .A2(P2_U3152), .ZN(n9952) );
  INV_X2 U8043 ( .A(n9952), .ZN(n7728) );
  NOR2_X1 U8044 ( .A1(n5634), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9954) );
  OAI222_X1 U8045 ( .A1(n7728), .A2(n6468), .B1(n8747), .B2(n6467), .C1(
        P2_U3152), .C2(n6580), .ZN(P2_U3357) );
  INV_X1 U8046 ( .A(n9756), .ZN(n6470) );
  NAND2_X1 U8047 ( .A1(n6470), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6469) );
  OAI21_X1 U8048 ( .B1(n6978), .B2(n6470), .A(n6469), .ZN(P1_U3440) );
  INV_X1 U8049 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6473) );
  INV_X1 U8050 ( .A(n7039), .ZN(n6471) );
  NAND2_X1 U8051 ( .A1(n6471), .A2(n9756), .ZN(n6472) );
  OAI21_X1 U8052 ( .B1(n9756), .B2(n6473), .A(n6472), .ZN(P1_U3441) );
  INV_X1 U8053 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6475) );
  INV_X1 U8054 ( .A(n6474), .ZN(n6480) );
  OAI222_X1 U8055 ( .A1(n8222), .A2(n6475), .B1(n9550), .B2(n6480), .C1(
        P1_U3084), .C2(n9635), .ZN(P1_U3347) );
  OAI222_X1 U8056 ( .A1(n7728), .A2(n6477), .B1(n8747), .B2(n6476), .C1(
        P2_U3152), .C2(n6653), .ZN(P2_U3356) );
  OAI222_X1 U8057 ( .A1(n7728), .A2(n6479), .B1(n8747), .B2(n6478), .C1(
        P2_U3152), .C2(n6619), .ZN(P2_U3353) );
  INV_X1 U8058 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6481) );
  INV_X1 U8059 ( .A(n6577), .ZN(n6607) );
  OAI222_X1 U8060 ( .A1(n7728), .A2(n6481), .B1(n8747), .B2(n6480), .C1(
        P2_U3152), .C2(n6607), .ZN(P2_U3352) );
  OAI222_X1 U8061 ( .A1(n7728), .A2(n6483), .B1(n8747), .B2(n6482), .C1(
        P2_U3152), .C2(n6667), .ZN(P2_U3354) );
  OAI222_X1 U8062 ( .A1(n7728), .A2(n6484), .B1(n8747), .B2(n8049), .C1(
        P2_U3152), .C2(n6679), .ZN(P2_U3355) );
  INV_X1 U8063 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10089) );
  INV_X1 U8064 ( .A(n6485), .ZN(n6487) );
  OAI222_X1 U8065 ( .A1(n8222), .A2(n10089), .B1(n9550), .B2(n6487), .C1(
        P1_U3084), .C2(n6486), .ZN(P1_U3346) );
  INV_X1 U8066 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6488) );
  INV_X1 U8067 ( .A(n6623), .ZN(n6630) );
  OAI222_X1 U8068 ( .A1(n7728), .A2(n6488), .B1(n8747), .B2(n6487), .C1(
        P2_U3152), .C2(n6630), .ZN(P2_U3351) );
  INV_X1 U8069 ( .A(n6489), .ZN(n6492) );
  OAI222_X1 U8070 ( .A1(n8222), .A2(n6491), .B1(n9550), .B2(n6492), .C1(
        P1_U3084), .C2(n6490), .ZN(P1_U3345) );
  INV_X1 U8071 ( .A(n6744), .ZN(n6749) );
  OAI222_X1 U8072 ( .A1(n7728), .A2(n10193), .B1(n8747), .B2(n6492), .C1(
        P2_U3152), .C2(n6749), .ZN(P2_U3350) );
  INV_X1 U8073 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6504) );
  INV_X1 U8074 ( .A(n9741), .ZN(n9655) );
  OAI21_X1 U8075 ( .B1(n6495), .B2(n6494), .A(n6493), .ZN(n6500) );
  INV_X1 U8076 ( .A(n9751), .ZN(n9731) );
  OAI21_X1 U8077 ( .B1(n6498), .B2(n6497), .A(n6496), .ZN(n6499) );
  AOI22_X1 U8078 ( .A1(n9655), .A2(n6500), .B1(n9731), .B2(n6499), .ZN(n6503)
         );
  NOR2_X1 U8079 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5166), .ZN(n7474) );
  AOI21_X1 U8080 ( .B1(n9714), .B2(n6501), .A(n7474), .ZN(n6502) );
  OAI211_X1 U8081 ( .C1(n9754), .C2(n6504), .A(n6503), .B(n6502), .ZN(P1_U3248) );
  INV_X1 U8082 ( .A(n6505), .ZN(n6508) );
  OAI222_X1 U8083 ( .A1(n8222), .A2(n6507), .B1(n9550), .B2(n6508), .C1(n6506), 
        .C2(P1_U3084), .ZN(P1_U3344) );
  INV_X1 U8084 ( .A(n6785), .ZN(n6755) );
  OAI222_X1 U8085 ( .A1(n7728), .A2(n6509), .B1(n8747), .B2(n6508), .C1(n6755), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U8086 ( .A(n9754), .ZN(n9623) );
  INV_X1 U8087 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6989) );
  OAI22_X1 U8088 ( .A1(n9745), .A2(n6510), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6989), .ZN(n6520) );
  OAI21_X1 U8089 ( .B1(n6513), .B2(n6512), .A(n6511), .ZN(n6518) );
  OAI21_X1 U8090 ( .B1(n6516), .B2(n6515), .A(n6514), .ZN(n6517) );
  OAI22_X1 U8091 ( .A1(n9741), .A2(n6518), .B1(n9751), .B2(n6517), .ZN(n6519)
         );
  AOI211_X1 U8092 ( .C1(n9623), .C2(P1_ADDR_REG_1__SCAN_IN), .A(n6520), .B(
        n6519), .ZN(n6521) );
  INV_X1 U8093 ( .A(n6521), .ZN(P1_U3242) );
  INV_X1 U8094 ( .A(n6862), .ZN(n6827) );
  OAI21_X1 U8095 ( .B1(n9819), .B2(n6827), .A(n6557), .ZN(n6523) );
  NAND2_X1 U8096 ( .A1(n9819), .A2(n7726), .ZN(n6522) );
  NAND2_X1 U8097 ( .A1(n6523), .A2(n6522), .ZN(n8388) );
  NOR2_X1 U8098 ( .A1(n9797), .A2(P2_U3966), .ZN(P2_U3151) );
  NAND2_X1 U8099 ( .A1(n5058), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6527) );
  INV_X1 U8100 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9220) );
  OR2_X1 U8101 ( .A1(n5142), .A2(n9220), .ZN(n6526) );
  INV_X1 U8102 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6524) );
  OR2_X1 U8103 ( .A1(n5057), .A2(n6524), .ZN(n6525) );
  INV_X1 U8104 ( .A(P1_U4006), .ZN(n6534) );
  NAND2_X1 U8105 ( .A1(n6534), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n6528) );
  OAI21_X1 U8106 ( .B1(n9219), .B2(n6534), .A(n6528), .ZN(P1_U3586) );
  NAND2_X1 U8107 ( .A1(n5058), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6532) );
  INV_X1 U8108 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9224) );
  OR2_X1 U8109 ( .A1(n5142), .A2(n9224), .ZN(n6531) );
  INV_X1 U8110 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n6529) );
  OR2_X1 U8111 ( .A1(n5057), .A2(n6529), .ZN(n6530) );
  AND3_X1 U8112 ( .A1(n6532), .A2(n6531), .A3(n6530), .ZN(n9240) );
  NAND2_X1 U8113 ( .A1(n6534), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6533) );
  OAI21_X1 U8114 ( .B1(n9240), .B2(n6534), .A(n6533), .ZN(P1_U3585) );
  INV_X1 U8115 ( .A(n6535), .ZN(n6538) );
  OAI222_X1 U8116 ( .A1(n8222), .A2(n6536), .B1(n9550), .B2(n6538), .C1(n6794), 
        .C2(P1_U3084), .ZN(P1_U3343) );
  INV_X1 U8117 ( .A(n7115), .ZN(n6792) );
  OAI222_X1 U8118 ( .A1(P2_U3152), .A2(n6792), .B1(n8747), .B2(n6538), .C1(
        n6537), .C2(n7728), .ZN(P2_U3348) );
  INV_X1 U8119 ( .A(n6539), .ZN(n6541) );
  INV_X1 U8120 ( .A(n7277), .ZN(n7272) );
  OAI222_X1 U8121 ( .A1(n7728), .A2(n6540), .B1(n8747), .B2(n6541), .C1(n7272), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U8122 ( .A(n9185), .ZN(n9173) );
  OAI222_X1 U8123 ( .A1(n8222), .A2(n6542), .B1(n9550), .B2(n6541), .C1(n9173), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  INV_X1 U8124 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6544) );
  NAND2_X1 U8125 ( .A1(P2_U3966), .A2(n6895), .ZN(n6543) );
  OAI21_X1 U8126 ( .B1(P2_U3966), .B2(n6544), .A(n6543), .ZN(P2_U3552) );
  INV_X1 U8127 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U8128 ( .A1(n8390), .A2(P2_U3966), .ZN(n6545) );
  OAI21_X1 U8129 ( .B1(P2_U3966), .B2(n6546), .A(n6545), .ZN(P2_U3583) );
  NAND2_X1 U8130 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n6554) );
  INV_X1 U8131 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6899) );
  XNOR2_X1 U8132 ( .A(n6580), .B(n6899), .ZN(n6553) );
  INV_X1 U8133 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6547) );
  INV_X1 U8134 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9800) );
  OR3_X1 U8135 ( .A1(n6553), .A2(n6547), .A3(n9800), .ZN(n6566) );
  INV_X1 U8136 ( .A(n6566), .ZN(n6552) );
  OAI21_X1 U8137 ( .B1(n6869), .B2(P2_U3152), .A(n7726), .ZN(n6548) );
  INV_X1 U8138 ( .A(n6548), .ZN(n6549) );
  OAI21_X1 U8139 ( .B1(n9819), .B2(n6862), .A(n6549), .ZN(n6559) );
  NAND2_X1 U8140 ( .A1(n6559), .A2(n6557), .ZN(n6550) );
  NAND2_X1 U8141 ( .A1(n6550), .A2(n8314), .ZN(n6555) );
  NOR2_X1 U8142 ( .A1(n6416), .A2(n8212), .ZN(n6551) );
  NAND2_X1 U8143 ( .A1(n6555), .A2(n6551), .ZN(n9792) );
  AOI211_X1 U8144 ( .C1(n6554), .C2(n6553), .A(n6552), .B(n9792), .ZN(n6565)
         );
  INV_X1 U8145 ( .A(n8384), .ZN(n9794) );
  AOI22_X1 U8146 ( .A1(n9797), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n6563) );
  AND2_X1 U8147 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(
        n6561) );
  INV_X1 U8148 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6556) );
  MUX2_X1 U8149 ( .A(n6556), .B(P2_REG1_REG_1__SCAN_IN), .S(n6580), .Z(n6560)
         );
  AND2_X1 U8150 ( .A1(n6557), .A2(n8212), .ZN(n6558) );
  NAND2_X1 U8151 ( .A1(n6560), .A2(n6561), .ZN(n6582) );
  OAI211_X1 U8152 ( .C1(n6561), .C2(n6560), .A(n9790), .B(n6582), .ZN(n6562)
         );
  OAI211_X1 U8153 ( .C1(n9794), .C2(n6580), .A(n6563), .B(n6562), .ZN(n6564)
         );
  OR2_X1 U8154 ( .A1(n6565), .A2(n6564), .ZN(P2_U3246) );
  INV_X1 U8155 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6567) );
  INV_X1 U8156 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6885) );
  OAI21_X1 U8157 ( .B1(n6899), .B2(n6580), .A(n6566), .ZN(n6649) );
  XNOR2_X1 U8158 ( .A(n6653), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n6650) );
  NAND2_X1 U8159 ( .A1(n6649), .A2(n6650), .ZN(n6648) );
  OAI21_X1 U8160 ( .B1(n6885), .B2(n6653), .A(n6648), .ZN(n6675) );
  XNOR2_X1 U8161 ( .A(n6679), .B(P2_REG2_REG_3__SCAN_IN), .ZN(n6676) );
  NAND2_X1 U8162 ( .A1(n6675), .A2(n6676), .ZN(n6674) );
  OAI21_X1 U8163 ( .B1(n6567), .B2(n6679), .A(n6674), .ZN(n6663) );
  NAND2_X1 U8164 ( .A1(n6655), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6568) );
  OAI21_X1 U8165 ( .B1(n6655), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6568), .ZN(
        n6569) );
  INV_X1 U8166 ( .A(n6569), .ZN(n6664) );
  NAND2_X1 U8167 ( .A1(n6663), .A2(n6664), .ZN(n6662) );
  INV_X1 U8168 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6570) );
  MUX2_X1 U8169 ( .A(n6570), .B(P2_REG2_REG_5__SCAN_IN), .S(n6578), .Z(n6611)
         );
  INV_X1 U8170 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6571) );
  MUX2_X1 U8171 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6571), .S(n6577), .Z(n6572)
         );
  INV_X1 U8172 ( .A(n6572), .ZN(n6600) );
  NOR2_X1 U8173 ( .A1(n6601), .A2(n6600), .ZN(n6599) );
  AOI21_X1 U8174 ( .B1(n6577), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6599), .ZN(
        n6575) );
  NAND2_X1 U8175 ( .A1(n6623), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6573) );
  OAI21_X1 U8176 ( .B1(n6623), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6573), .ZN(
        n6574) );
  AOI211_X1 U8177 ( .C1(n6575), .C2(n6574), .A(n6622), .B(n9792), .ZN(n6598)
         );
  NOR2_X1 U8178 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5930), .ZN(n6576) );
  AOI21_X1 U8179 ( .B1(n9797), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6576), .ZN(
        n6596) );
  INV_X1 U8180 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9915) );
  MUX2_X1 U8181 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9915), .S(n6577), .Z(n6603)
         );
  NAND2_X1 U8182 ( .A1(n6578), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6591) );
  INV_X1 U8183 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6579) );
  MUX2_X1 U8184 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6579), .S(n6578), .Z(n6615)
         );
  XNOR2_X1 U8185 ( .A(n6653), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n6642) );
  OR2_X1 U8186 ( .A1(n6580), .A2(n6556), .ZN(n6581) );
  NAND2_X1 U8187 ( .A1(n6582), .A2(n6581), .ZN(n6643) );
  NAND2_X1 U8188 ( .A1(n6642), .A2(n6643), .ZN(n6585) );
  INV_X1 U8189 ( .A(n6653), .ZN(n6583) );
  NAND2_X1 U8190 ( .A1(n6583), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6584) );
  NAND2_X1 U8191 ( .A1(n6585), .A2(n6584), .ZN(n6668) );
  INV_X1 U8192 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6586) );
  MUX2_X1 U8193 ( .A(n6586), .B(P2_REG1_REG_3__SCAN_IN), .S(n6679), .Z(n6587)
         );
  AND2_X1 U8194 ( .A1(n6668), .A2(n6587), .ZN(n6669) );
  NOR2_X1 U8195 ( .A1(n6679), .A2(n6586), .ZN(n6654) );
  INV_X1 U8196 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6588) );
  MUX2_X1 U8197 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6588), .S(n6655), .Z(n6589)
         );
  OAI21_X1 U8198 ( .B1(n6669), .B2(n6654), .A(n6589), .ZN(n6660) );
  NAND2_X1 U8199 ( .A1(n6655), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6590) );
  NAND2_X1 U8200 ( .A1(n6660), .A2(n6590), .ZN(n6616) );
  NAND2_X1 U8201 ( .A1(n6615), .A2(n6616), .ZN(n6614) );
  NAND2_X1 U8202 ( .A1(n6591), .A2(n6614), .ZN(n6604) );
  NAND2_X1 U8203 ( .A1(n6603), .A2(n6604), .ZN(n6602) );
  OAI21_X1 U8204 ( .B1(n6607), .B2(n9915), .A(n6602), .ZN(n6594) );
  INV_X1 U8205 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6592) );
  MUX2_X1 U8206 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6592), .S(n6623), .Z(n6593)
         );
  NAND2_X1 U8207 ( .A1(n6593), .A2(n6594), .ZN(n6629) );
  OAI211_X1 U8208 ( .C1(n6594), .C2(n6593), .A(n9790), .B(n6629), .ZN(n6595)
         );
  OAI211_X1 U8209 ( .C1(n9794), .C2(n6630), .A(n6596), .B(n6595), .ZN(n6597)
         );
  OR2_X1 U8210 ( .A1(n6598), .A2(n6597), .ZN(P2_U3252) );
  AOI211_X1 U8211 ( .C1(n6601), .C2(n6600), .A(n6599), .B(n9792), .ZN(n6609)
         );
  INV_X1 U8212 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9982) );
  NOR2_X1 U8213 ( .A1(n9982), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7136) );
  AOI21_X1 U8214 ( .B1(n9797), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n7136), .ZN(
        n6606) );
  OAI211_X1 U8215 ( .C1(n6604), .C2(n6603), .A(n9790), .B(n6602), .ZN(n6605)
         );
  OAI211_X1 U8216 ( .C1(n9794), .C2(n6607), .A(n6606), .B(n6605), .ZN(n6608)
         );
  OR2_X1 U8217 ( .A1(n6609), .A2(n6608), .ZN(P2_U3251) );
  AOI211_X1 U8218 ( .C1(n6612), .C2(n6611), .A(n6610), .B(n9792), .ZN(n6621)
         );
  INV_X1 U8219 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6923) );
  NOR2_X1 U8220 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6923), .ZN(n6613) );
  AOI21_X1 U8221 ( .B1(n9797), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6613), .ZN(
        n6618) );
  OAI211_X1 U8222 ( .C1(n6616), .C2(n6615), .A(n9790), .B(n6614), .ZN(n6617)
         );
  OAI211_X1 U8223 ( .C1(n9794), .C2(n6619), .A(n6618), .B(n6617), .ZN(n6620)
         );
  OR2_X1 U8224 ( .A1(n6621), .A2(n6620), .ZN(P2_U3250) );
  INV_X1 U8225 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6624) );
  MUX2_X1 U8226 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n6624), .S(n6744), .Z(n6625)
         );
  INV_X1 U8227 ( .A(n6625), .ZN(n6626) );
  AOI211_X1 U8228 ( .C1(n6627), .C2(n6626), .A(n6743), .B(n9792), .ZN(n6636)
         );
  NAND2_X1 U8229 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n7468) );
  INV_X1 U8230 ( .A(n7468), .ZN(n6628) );
  AOI21_X1 U8231 ( .B1(n9797), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6628), .ZN(
        n6634) );
  OAI21_X1 U8232 ( .B1(n6630), .B2(n6592), .A(n6629), .ZN(n6632) );
  MUX2_X1 U8233 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10141), .S(n6744), .Z(n6631)
         );
  NAND2_X1 U8234 ( .A1(n6631), .A2(n6632), .ZN(n6748) );
  OAI211_X1 U8235 ( .C1(n6632), .C2(n6631), .A(n9790), .B(n6748), .ZN(n6633)
         );
  OAI211_X1 U8236 ( .C1(n9794), .C2(n6749), .A(n6634), .B(n6633), .ZN(n6635)
         );
  OR2_X1 U8237 ( .A1(n6636), .A2(n6635), .ZN(P2_U3253) );
  INV_X1 U8238 ( .A(n8872), .ZN(n8860) );
  INV_X1 U8239 ( .A(n7348), .ZN(n7073) );
  NAND2_X1 U8240 ( .A1(n6685), .A2(n8850), .ZN(n6641) );
  INV_X1 U8241 ( .A(n8865), .ZN(n8857) );
  INV_X1 U8242 ( .A(n7041), .ZN(n7151) );
  NAND3_X1 U8243 ( .A1(n7150), .A2(n7151), .A3(n6639), .ZN(n6720) );
  AOI22_X1 U8244 ( .A1(n8857), .A2(n6974), .B1(n6720), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n6640) );
  OAI211_X1 U8245 ( .C1(n8860), .C2(n7073), .A(n6641), .B(n6640), .ZN(P1_U3230) );
  XOR2_X1 U8246 ( .A(n6643), .B(n6642), .Z(n6647) );
  INV_X1 U8247 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6645) );
  INV_X1 U8248 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6644) );
  OAI22_X1 U8249 ( .A1(n8388), .A2(n6645), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6644), .ZN(n6646) );
  AOI21_X1 U8250 ( .B1(n9790), .B2(n6647), .A(n6646), .ZN(n6652) );
  OAI211_X1 U8251 ( .C1(n6650), .C2(n6649), .A(n9791), .B(n6648), .ZN(n6651)
         );
  OAI211_X1 U8252 ( .C1(n9794), .C2(n6653), .A(n6652), .B(n6651), .ZN(P2_U3247) );
  INV_X1 U8253 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10166) );
  NOR2_X1 U8254 ( .A1(n10166), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6938) );
  INV_X1 U8255 ( .A(n6669), .ZN(n6658) );
  INV_X1 U8256 ( .A(n6654), .ZN(n6657) );
  MUX2_X1 U8257 ( .A(n6588), .B(P2_REG1_REG_4__SCAN_IN), .S(n6655), .Z(n6656)
         );
  NAND3_X1 U8258 ( .A1(n6658), .A2(n6657), .A3(n6656), .ZN(n6659) );
  AND3_X1 U8259 ( .A1(n9790), .A2(n6660), .A3(n6659), .ZN(n6661) );
  AOI211_X1 U8260 ( .C1(n9797), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6938), .B(
        n6661), .ZN(n6666) );
  OAI211_X1 U8261 ( .C1(n6664), .C2(n6663), .A(n9791), .B(n6662), .ZN(n6665)
         );
  OAI211_X1 U8262 ( .C1(n9794), .C2(n6667), .A(n6666), .B(n6665), .ZN(P2_U3249) );
  NOR2_X1 U8263 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5886), .ZN(n6673) );
  INV_X1 U8264 ( .A(n6668), .ZN(n6671) );
  MUX2_X1 U8265 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6586), .S(n6679), .Z(n6670)
         );
  AOI211_X1 U8266 ( .C1(n6671), .C2(n6670), .A(n6669), .B(n9795), .ZN(n6672)
         );
  AOI211_X1 U8267 ( .C1(n9797), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n6673), .B(
        n6672), .ZN(n6678) );
  OAI211_X1 U8268 ( .C1(n6676), .C2(n6675), .A(n9791), .B(n6674), .ZN(n6677)
         );
  OAI211_X1 U8269 ( .C1(n9794), .C2(n6679), .A(n6678), .B(n6677), .ZN(P2_U3248) );
  NAND2_X1 U8270 ( .A1(n6680), .A2(P1_U4006), .ZN(n6681) );
  OAI21_X1 U8271 ( .B1(P1_U4006), .B2(n5870), .A(n6681), .ZN(P1_U3555) );
  INV_X1 U8272 ( .A(n6682), .ZN(n6684) );
  INV_X1 U8273 ( .A(n7427), .ZN(n7422) );
  OAI222_X1 U8274 ( .A1(n7728), .A2(n6683), .B1(n8747), .B2(n6684), .C1(
        P2_U3152), .C2(n7422), .ZN(P2_U3346) );
  OAI222_X1 U8275 ( .A1(n8222), .A2(n10194), .B1(n9550), .B2(n6684), .C1(
        P1_U3084), .C2(n9189), .ZN(P1_U3341) );
  INV_X1 U8276 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7560) );
  INV_X1 U8277 ( .A(n6685), .ZN(n6687) );
  INV_X1 U8278 ( .A(n6688), .ZN(n9217) );
  AOI21_X1 U8279 ( .B1(n9217), .B2(n6686), .A(n5798), .ZN(n9592) );
  OAI21_X1 U8280 ( .B1(n6687), .B2(n9217), .A(n9592), .ZN(n6691) );
  OAI21_X1 U8281 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n6688), .A(n6996), .ZN(
        n6689) );
  AOI21_X1 U8282 ( .B1(n6689), .B2(n4999), .A(P1_U3084), .ZN(n9593) );
  NAND3_X1 U8283 ( .A1(n6691), .A2(n6690), .A3(n9593), .ZN(n9607) );
  AOI22_X1 U8284 ( .A1(n9714), .A2(n6692), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        P1_U3084), .ZN(n6701) );
  OAI211_X1 U8285 ( .C1(n6695), .C2(n6694), .A(n9655), .B(n6693), .ZN(n6700)
         );
  OAI211_X1 U8286 ( .C1(n6698), .C2(n6697), .A(n9731), .B(n6696), .ZN(n6699)
         );
  AND3_X1 U8287 ( .A1(n6701), .A2(n6700), .A3(n6699), .ZN(n6702) );
  OAI211_X1 U8288 ( .C1(n7560), .C2(n9754), .A(n9607), .B(n6702), .ZN(P1_U3243) );
  INV_X1 U8289 ( .A(n6703), .ZN(n6738) );
  AOI22_X1 U8290 ( .A1(n9191), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9548), .ZN(n6704) );
  OAI21_X1 U8291 ( .B1(n6738), .B2(n9550), .A(n6704), .ZN(P1_U3340) );
  OAI21_X1 U8292 ( .B1(n6707), .B2(n6706), .A(n6705), .ZN(n6712) );
  INV_X1 U8293 ( .A(n7157), .ZN(n7238) );
  AOI22_X1 U8294 ( .A1(n8857), .A2(n7157), .B1(n8868), .B2(n6974), .ZN(n6710)
         );
  NAND2_X1 U8295 ( .A1(n6720), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6709) );
  OAI211_X1 U8296 ( .C1(n7357), .C2(n8860), .A(n6710), .B(n6709), .ZN(n6711)
         );
  AOI21_X1 U8297 ( .B1(n6712), .B2(n8850), .A(n6711), .ZN(n6713) );
  INV_X1 U8298 ( .A(n6713), .ZN(P1_U3235) );
  NAND2_X1 U8299 ( .A1(n6714), .A2(n6715), .ZN(n6716) );
  XOR2_X1 U8300 ( .A(n6717), .B(n6716), .Z(n6724) );
  AOI22_X1 U8301 ( .A1(n8857), .A2(n6719), .B1(n8868), .B2(n6680), .ZN(n6722)
         );
  NAND2_X1 U8302 ( .A1(n6720), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6721) );
  OAI211_X1 U8303 ( .C1(n6975), .C2(n8860), .A(n6722), .B(n6721), .ZN(n6723)
         );
  AOI21_X1 U8304 ( .B1(n6724), .B2(n8850), .A(n6723), .ZN(n6725) );
  INV_X1 U8305 ( .A(n6725), .ZN(P1_U3220) );
  NOR2_X1 U8306 ( .A1(n6731), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6727) );
  NOR2_X1 U8307 ( .A1(n6727), .A2(n6726), .ZN(n6729) );
  INV_X1 U8308 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7517) );
  AOI22_X1 U8309 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n6794), .B1(n6799), .B2(
        n7517), .ZN(n6728) );
  NOR2_X1 U8310 ( .A1(n6729), .A2(n6728), .ZN(n6793) );
  AOI21_X1 U8311 ( .B1(n6729), .B2(n6728), .A(n6793), .ZN(n6737) );
  NAND2_X1 U8312 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7657) );
  OAI21_X1 U8313 ( .B1(n9745), .B2(n6794), .A(n7657), .ZN(n6735) );
  MUX2_X1 U8314 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n7339), .S(n6794), .Z(n6732)
         );
  NOR2_X1 U8315 ( .A1(n6733), .A2(n6732), .ZN(n6798) );
  AOI211_X1 U8316 ( .C1(n6733), .C2(n6732), .A(n6798), .B(n9741), .ZN(n6734)
         );
  AOI211_X1 U8317 ( .C1(P1_ADDR_REG_10__SCAN_IN), .C2(n9623), .A(n6735), .B(
        n6734), .ZN(n6736) );
  OAI21_X1 U8318 ( .B1(n6737), .B2(n9751), .A(n6736), .ZN(P1_U3251) );
  INV_X1 U8319 ( .A(n7528), .ZN(n7523) );
  OAI222_X1 U8320 ( .A1(n7728), .A2(n6739), .B1(n8747), .B2(n6738), .C1(n7523), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8321 ( .A(n6740), .ZN(n6741) );
  OAI222_X1 U8322 ( .A1(n8222), .A2(n10015), .B1(n9550), .B2(n6741), .C1(n9690), .C2(P1_U3084), .ZN(P1_U3339) );
  INV_X1 U8323 ( .A(n7918), .ZN(n7911) );
  OAI222_X1 U8324 ( .A1(n7728), .A2(n6742), .B1(n8747), .B2(n6741), .C1(n7911), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  NAND2_X1 U8325 ( .A1(n6785), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6745) );
  OAI21_X1 U8326 ( .B1(n6785), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6745), .ZN(
        n6746) );
  NOR2_X1 U8327 ( .A1(n4409), .A2(n6746), .ZN(n6784) );
  AOI211_X1 U8328 ( .C1(n4409), .C2(n6746), .A(n6784), .B(n9792), .ZN(n6757)
         );
  NAND2_X1 U8329 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7506) );
  INV_X1 U8330 ( .A(n7506), .ZN(n6747) );
  AOI21_X1 U8331 ( .B1(n9797), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n6747), .ZN(
        n6754) );
  INV_X1 U8332 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10141) );
  OAI21_X1 U8333 ( .B1(n6749), .B2(n10141), .A(n6748), .ZN(n6752) );
  INV_X1 U8334 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6750) );
  MUX2_X1 U8335 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n6750), .S(n6785), .Z(n6751)
         );
  NAND2_X1 U8336 ( .A1(n6751), .A2(n6752), .ZN(n6778) );
  OAI211_X1 U8337 ( .C1(n6752), .C2(n6751), .A(n9790), .B(n6778), .ZN(n6753)
         );
  OAI211_X1 U8338 ( .C1(n9794), .C2(n6755), .A(n6754), .B(n6753), .ZN(n6756)
         );
  OR2_X1 U8339 ( .A1(n6757), .A2(n6756), .ZN(P2_U3254) );
  OAI21_X1 U8340 ( .B1(n6758), .B2(n6760), .A(n6759), .ZN(n6761) );
  NAND2_X1 U8341 ( .A1(n6761), .A2(n8850), .ZN(n6767) );
  NAND2_X1 U8342 ( .A1(n8868), .A2(n6719), .ZN(n6763) );
  AND2_X1 U8343 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8060) );
  INV_X1 U8344 ( .A(n8060), .ZN(n6762) );
  OAI211_X1 U8345 ( .C1(n7368), .C2(n8865), .A(n6763), .B(n6762), .ZN(n6765)
         );
  NOR2_X1 U8346 ( .A1(n8870), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6764) );
  AOI211_X1 U8347 ( .C1(n8872), .C2(n7380), .A(n6765), .B(n6764), .ZN(n6766)
         );
  NAND2_X1 U8348 ( .A1(n6767), .A2(n6766), .ZN(P1_U3216) );
  AOI21_X1 U8349 ( .B1(n6768), .B2(n6769), .A(n8874), .ZN(n6771) );
  NAND2_X1 U8350 ( .A1(n6771), .A2(n6770), .ZN(n6777) );
  INV_X1 U8351 ( .A(n9169), .ZN(n7311) );
  NAND2_X1 U8352 ( .A1(n8868), .A2(n7157), .ZN(n6772) );
  OAI211_X1 U8353 ( .C1(n7311), .C2(n8865), .A(n6772), .B(n4935), .ZN(n6775)
         );
  INV_X1 U8354 ( .A(n6773), .ZN(n7437) );
  NOR2_X1 U8355 ( .A1(n8870), .A2(n7437), .ZN(n6774) );
  AOI211_X1 U8356 ( .C1(n8872), .C2(n7246), .A(n6775), .B(n6774), .ZN(n6776)
         );
  NAND2_X1 U8357 ( .A1(n6777), .A2(n6776), .ZN(P1_U3228) );
  NAND2_X1 U8358 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n7539) );
  INV_X1 U8359 ( .A(n7539), .ZN(n6783) );
  INV_X1 U8360 ( .A(n6778), .ZN(n6779) );
  AOI21_X1 U8361 ( .B1(n6785), .B2(P2_REG1_REG_9__SCAN_IN), .A(n6779), .ZN(
        n6781) );
  INV_X1 U8362 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9981) );
  MUX2_X1 U8363 ( .A(n9981), .B(P2_REG1_REG_10__SCAN_IN), .S(n7115), .Z(n6780)
         );
  NOR2_X1 U8364 ( .A1(n6780), .A2(n6781), .ZN(n7110) );
  AOI211_X1 U8365 ( .C1(n6781), .C2(n6780), .A(n7110), .B(n9795), .ZN(n6782)
         );
  AOI211_X1 U8366 ( .C1(n9797), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n6783), .B(
        n6782), .ZN(n6791) );
  XOR2_X1 U8367 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7115), .Z(n6789) );
  INV_X1 U8368 ( .A(n6786), .ZN(n6788) );
  INV_X1 U8369 ( .A(n6789), .ZN(n6787) );
  OAI211_X1 U8370 ( .C1(n6789), .C2(n6788), .A(n9791), .B(n7114), .ZN(n6790)
         );
  OAI211_X1 U8371 ( .C1(n9794), .C2(n6792), .A(n6791), .B(n6790), .ZN(P2_U3255) );
  AOI21_X1 U8372 ( .B1(n7517), .B2(n6794), .A(n6793), .ZN(n6797) );
  INV_X1 U8373 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6795) );
  MUX2_X1 U8374 ( .A(n6795), .B(P1_REG1_REG_11__SCAN_IN), .S(n9185), .Z(n6796)
         );
  NOR2_X1 U8375 ( .A1(n6797), .A2(n6796), .ZN(n9172) );
  AOI21_X1 U8376 ( .B1(n6797), .B2(n6796), .A(n9172), .ZN(n6804) );
  XNOR2_X1 U8377 ( .A(n9185), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n9184) );
  AOI21_X1 U8378 ( .B1(n6799), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6798), .ZN(
        n9187) );
  XNOR2_X1 U8379 ( .A(n9184), .B(n9187), .ZN(n6801) );
  NAND2_X1 U8380 ( .A1(n9714), .A2(n9185), .ZN(n6800) );
  NAND2_X1 U8381 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7788) );
  OAI211_X1 U8382 ( .C1(n6801), .C2(n9741), .A(n6800), .B(n7788), .ZN(n6802)
         );
  AOI21_X1 U8383 ( .B1(n9623), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n6802), .ZN(
        n6803) );
  OAI21_X1 U8384 ( .B1(n6804), .B2(n9751), .A(n6803), .ZN(P1_U3252) );
  XNOR2_X1 U8385 ( .A(n7836), .B(P2_B_REG_SCAN_IN), .ZN(n6805) );
  NAND2_X1 U8386 ( .A1(n6805), .A2(n7945), .ZN(n6807) );
  INV_X1 U8387 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6809) );
  NAND2_X1 U8388 ( .A1(n7945), .A2(n7976), .ZN(n9843) );
  INV_X1 U8389 ( .A(n9843), .ZN(n6808) );
  INV_X1 U8390 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6810) );
  NAND2_X1 U8391 ( .A1(n9820), .A2(n6810), .ZN(n6811) );
  NAND2_X1 U8392 ( .A1(n7836), .A2(n7976), .ZN(n9841) );
  NAND2_X1 U8393 ( .A1(n7008), .A2(n7026), .ZN(n6821) );
  NOR4_X1 U8394 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n6818) );
  INV_X1 U8395 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n9987) );
  INV_X1 U8396 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n9973) );
  INV_X1 U8397 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10105) );
  INV_X1 U8398 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n9971) );
  NAND4_X1 U8399 ( .A1(n9987), .A2(n9973), .A3(n10105), .A4(n9971), .ZN(n10201) );
  NOR4_X1 U8400 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6815) );
  NOR4_X1 U8401 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6814) );
  NOR4_X1 U8402 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n6813) );
  NOR4_X1 U8403 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6812) );
  NAND4_X1 U8404 ( .A1(n6815), .A2(n6814), .A3(n6813), .A4(n6812), .ZN(n6816)
         );
  NOR4_X1 U8405 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        n10201), .A4(n6816), .ZN(n6817) );
  NOR4_X1 U8406 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n10191) );
  NAND3_X1 U8407 ( .A1(n6818), .A2(n6817), .A3(n10191), .ZN(n6819) );
  NAND2_X1 U8408 ( .A1(n9820), .A2(n6819), .ZN(n6861) );
  NOR2_X1 U8409 ( .A1(n9819), .A2(n6868), .ZN(n6820) );
  NAND2_X1 U8410 ( .A1(n6861), .A2(n6820), .ZN(n7006) );
  INV_X1 U8411 ( .A(n7007), .ZN(n6864) );
  XNOR2_X1 U8412 ( .A(n6822), .B(n6823), .ZN(n6830) );
  NAND2_X1 U8413 ( .A1(n8325), .A2(n8590), .ZN(n6828) );
  OAI21_X1 U8414 ( .B1(n6942), .B2(n8615), .A(n6828), .ZN(n6829) );
  AOI21_X1 U8415 ( .B1(n6830), .B2(n8585), .A(n6829), .ZN(n9873) );
  NAND2_X1 U8416 ( .A1(n7581), .A2(n7010), .ZN(n6850) );
  NOR2_X1 U8417 ( .A1(n6850), .A2(n6227), .ZN(n9802) );
  NAND2_X1 U8418 ( .A1(n9817), .A2(n9802), .ZN(n8629) );
  XNOR2_X1 U8419 ( .A(n6393), .B(n6850), .ZN(n6831) );
  NAND2_X1 U8420 ( .A1(n6831), .A2(n6227), .ZN(n9805) );
  INV_X1 U8421 ( .A(n9805), .ZN(n8621) );
  NAND2_X1 U8422 ( .A1(n9817), .A2(n8621), .ZN(n6832) );
  INV_X1 U8423 ( .A(n8606), .ZN(n8541) );
  NAND2_X1 U8424 ( .A1(n6860), .A2(n9859), .ZN(n6836) );
  NAND2_X1 U8425 ( .A1(n6959), .A2(n6961), .ZN(n6958) );
  NAND2_X1 U8426 ( .A1(n6942), .A2(n6970), .ZN(n6837) );
  NAND2_X1 U8427 ( .A1(n6958), .A2(n6837), .ZN(n6839) );
  NAND2_X1 U8428 ( .A1(n6839), .A2(n6838), .ZN(n7087) );
  OR2_X1 U8429 ( .A1(n6839), .A2(n6838), .ZN(n6840) );
  NAND2_X1 U8430 ( .A1(n7087), .A2(n6840), .ZN(n9866) );
  NOR2_X1 U8431 ( .A1(n6394), .A2(n7010), .ZN(n9808) );
  NOR2_X1 U8432 ( .A1(n4385), .A2(n9847), .ZN(n6879) );
  AND2_X1 U8433 ( .A1(n6879), .A2(n9859), .ZN(n6965) );
  NAND2_X1 U8434 ( .A1(n6965), .A2(n6970), .ZN(n6967) );
  NAND2_X1 U8435 ( .A1(n6967), .A2(n9867), .ZN(n6842) );
  AND2_X1 U8436 ( .A1(n7253), .A2(n6842), .ZN(n9870) );
  NOR2_X1 U8437 ( .A1(n8469), .A2(n6843), .ZN(n6844) );
  AOI21_X1 U8438 ( .B1(n8632), .B2(n9870), .A(n6844), .ZN(n6847) );
  INV_X1 U8439 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6845) );
  OR2_X1 U8440 ( .A1(n9817), .A2(n6845), .ZN(n6846) );
  OAI211_X1 U8441 ( .C1(n7085), .C2(n8626), .A(n6847), .B(n6846), .ZN(n6848)
         );
  AOI21_X1 U8442 ( .B1(n8541), .B2(n9866), .A(n6848), .ZN(n6849) );
  OAI21_X1 U8443 ( .B1(n8600), .B2(n9873), .A(n6849), .ZN(P2_U3292) );
  INV_X1 U8444 ( .A(n6855), .ZN(n6854) );
  INV_X1 U8445 ( .A(n6856), .ZN(n6853) );
  NAND2_X1 U8446 ( .A1(n6854), .A2(n6853), .ZN(n6859) );
  NAND2_X1 U8447 ( .A1(n6856), .A2(n6855), .ZN(n6857) );
  NOR2_X1 U8448 ( .A1(n8163), .A2(n9847), .ZN(n6858) );
  AOI21_X1 U8449 ( .B1(n6892), .B2(n8148), .A(n6858), .ZN(n6948) );
  XNOR2_X1 U8450 ( .A(n9859), .B(n8163), .ZN(n6905) );
  XNOR2_X1 U8451 ( .A(n6904), .B(n6905), .ZN(n6909) );
  XNOR2_X1 U8452 ( .A(n6910), .B(n6909), .ZN(n6877) );
  NAND3_X1 U8453 ( .A1(n7009), .A2(n7008), .A3(n6861), .ZN(n6865) );
  INV_X1 U8454 ( .A(n6874), .ZN(n6863) );
  NAND2_X1 U8455 ( .A1(n6865), .A2(n6864), .ZN(n6872) );
  INV_X1 U8456 ( .A(n6866), .ZN(n6867) );
  NOR2_X1 U8457 ( .A1(n6868), .A2(n6867), .ZN(n6870) );
  AND2_X1 U8458 ( .A1(n6870), .A2(n6869), .ZN(n6871) );
  NAND2_X1 U8459 ( .A1(n6872), .A2(n6871), .ZN(n6921) );
  OR2_X1 U8460 ( .A1(n6921), .A2(P2_U3152), .ZN(n7037) );
  AOI22_X1 U8461 ( .A1(n8308), .A2(n6889), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n7037), .ZN(n6876) );
  OR2_X1 U8462 ( .A1(n6874), .A2(n6873), .ZN(n8170) );
  INV_X1 U8463 ( .A(n8302), .ZN(n8280) );
  INV_X1 U8464 ( .A(n8304), .ZN(n8281) );
  AOI22_X1 U8465 ( .A1(n8280), .A2(n6834), .B1(n8281), .B2(n8327), .ZN(n6875)
         );
  OAI211_X1 U8466 ( .C1(n6877), .C2(n8296), .A(n6876), .B(n6875), .ZN(P2_U3239) );
  XNOR2_X1 U8467 ( .A(n6878), .B(n6882), .ZN(n9858) );
  INV_X1 U8468 ( .A(n8626), .ZN(n8473) );
  NOR2_X1 U8469 ( .A1(n6879), .A2(n9859), .ZN(n6880) );
  OR2_X1 U8470 ( .A1(n6965), .A2(n6880), .ZN(n9860) );
  XNOR2_X1 U8471 ( .A(n6882), .B(n6881), .ZN(n6884) );
  OAI22_X1 U8472 ( .A1(n7033), .A2(n8615), .B1(n6942), .B2(n8617), .ZN(n6883)
         );
  AOI21_X1 U8473 ( .B1(n6884), .B2(n8585), .A(n6883), .ZN(n9861) );
  MUX2_X1 U8474 ( .A(n6885), .B(n9861), .S(n9817), .Z(n6887) );
  NAND2_X1 U8475 ( .A1(n9810), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6886) );
  OAI211_X1 U8476 ( .C1(n8475), .C2(n9860), .A(n6887), .B(n6886), .ZN(n6888)
         );
  AOI21_X1 U8477 ( .B1(n8473), .B2(n6889), .A(n6888), .ZN(n6890) );
  OAI21_X1 U8478 ( .B1(n8606), .B2(n9858), .A(n6890), .ZN(P2_U3294) );
  OAI21_X1 U8479 ( .B1(n6893), .B2(n6892), .A(n6891), .ZN(n9851) );
  XNOR2_X1 U8480 ( .A(n6893), .B(n7032), .ZN(n6894) );
  NAND2_X1 U8481 ( .A1(n6894), .A2(n8585), .ZN(n6897) );
  AOI22_X1 U8482 ( .A1(n8328), .A2(n8590), .B1(n8591), .B2(n6895), .ZN(n6896)
         );
  NAND2_X1 U8483 ( .A1(n6897), .A2(n6896), .ZN(n9854) );
  NAND2_X1 U8484 ( .A1(n9817), .A2(n9854), .ZN(n6898) );
  OAI21_X1 U8485 ( .B1(n9817), .B2(n6899), .A(n6898), .ZN(n6902) );
  XNOR2_X1 U8486 ( .A(n4386), .B(n9847), .ZN(n9853) );
  INV_X1 U8487 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6900) );
  OAI22_X1 U8488 ( .A1(n8475), .A2(n9853), .B1(n6900), .B2(n8469), .ZN(n6901)
         );
  AOI211_X1 U8489 ( .C1(n8473), .C2(n4386), .A(n6902), .B(n6901), .ZN(n6903)
         );
  OAI21_X1 U8490 ( .B1(n8606), .B2(n9851), .A(n6903), .ZN(P2_U3295) );
  INV_X1 U8491 ( .A(n6904), .ZN(n6907) );
  INV_X1 U8492 ( .A(n6905), .ZN(n6906) );
  NAND2_X1 U8493 ( .A1(n6907), .A2(n6906), .ZN(n6908) );
  OR2_X1 U8494 ( .A1(n6942), .A2(n8162), .ZN(n6913) );
  XNOR2_X1 U8495 ( .A(n8163), .B(n7012), .ZN(n6911) );
  XNOR2_X1 U8496 ( .A(n6913), .B(n6911), .ZN(n6930) );
  INV_X1 U8497 ( .A(n6911), .ZN(n6912) );
  NOR2_X1 U8498 ( .A1(n6913), .A2(n6912), .ZN(n6914) );
  AOI21_X1 U8499 ( .B1(n6929), .B2(n6930), .A(n6914), .ZN(n6935) );
  NOR2_X1 U8500 ( .A1(n7262), .A2(n8162), .ZN(n6915) );
  XNOR2_X1 U8501 ( .A(n8163), .B(n9867), .ZN(n6916) );
  NAND2_X1 U8502 ( .A1(n6915), .A2(n6916), .ZN(n6919) );
  INV_X1 U8503 ( .A(n6915), .ZN(n6918) );
  INV_X1 U8504 ( .A(n6916), .ZN(n6917) );
  NAND2_X1 U8505 ( .A1(n6918), .A2(n6917), .ZN(n6920) );
  AND2_X1 U8506 ( .A1(n6919), .A2(n6920), .ZN(n6937) );
  NAND2_X1 U8507 ( .A1(n6935), .A2(n6937), .ZN(n6936) );
  NAND2_X1 U8508 ( .A1(n6936), .A2(n6920), .ZN(n7123) );
  XNOR2_X1 U8509 ( .A(n8152), .B(n9807), .ZN(n7126) );
  NAND2_X1 U8510 ( .A1(n8325), .A2(n8148), .ZN(n7125) );
  XNOR2_X1 U8511 ( .A(n7126), .B(n7125), .ZN(n7124) );
  XNOR2_X1 U8512 ( .A(n7123), .B(n7124), .ZN(n6928) );
  NAND2_X1 U8513 ( .A1(n8293), .A2(n9809), .ZN(n6922) );
  OAI21_X1 U8514 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n6923), .A(n6922), .ZN(n6926) );
  OAI22_X1 U8515 ( .A1(n8247), .A2(n6924), .B1(n7263), .B2(n8304), .ZN(n6925)
         );
  AOI211_X1 U8516 ( .C1(n8280), .C2(n8326), .A(n6926), .B(n6925), .ZN(n6927)
         );
  OAI21_X1 U8517 ( .B1(n6928), .B2(n8296), .A(n6927), .ZN(P2_U3229) );
  XNOR2_X1 U8518 ( .A(n6929), .B(n6930), .ZN(n6934) );
  OAI22_X1 U8519 ( .A1(n8301), .A2(P2_REG3_REG_3__SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(n5886), .ZN(n6932) );
  OAI22_X1 U8520 ( .A1(n8247), .A2(n6970), .B1(n7262), .B2(n8304), .ZN(n6931)
         );
  AOI211_X1 U8521 ( .C1(n8280), .C2(n8328), .A(n6932), .B(n6931), .ZN(n6933)
         );
  OAI21_X1 U8522 ( .B1(n8296), .B2(n6934), .A(n6933), .ZN(P2_U3220) );
  OAI21_X1 U8523 ( .B1(n6935), .B2(n6937), .A(n6936), .ZN(n6945) );
  INV_X1 U8524 ( .A(n6938), .ZN(n6941) );
  NAND2_X1 U8525 ( .A1(n8293), .A2(n6939), .ZN(n6940) );
  OAI211_X1 U8526 ( .C1(n8302), .C2(n6942), .A(n6941), .B(n6940), .ZN(n6944)
         );
  OAI22_X1 U8527 ( .A1(n8247), .A2(n7085), .B1(n7140), .B2(n8304), .ZN(n6943)
         );
  AOI211_X1 U8528 ( .C1(n8298), .C2(n6945), .A(n6944), .B(n6943), .ZN(n6946)
         );
  INV_X1 U8529 ( .A(n6946), .ZN(P2_U3232) );
  AOI22_X1 U8530 ( .A1(n8308), .A2(n4386), .B1(n8281), .B2(n8328), .ZN(n6952)
         );
  OAI21_X1 U8531 ( .B1(n6949), .B2(n6948), .A(n6947), .ZN(n6950) );
  AOI22_X1 U8532 ( .A1(n8298), .A2(n6950), .B1(n7037), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n6951) );
  OAI211_X1 U8533 ( .C1(n6953), .C2(n8302), .A(n6952), .B(n6951), .ZN(P2_U3224) );
  INV_X1 U8534 ( .A(n6954), .ZN(n6956) );
  INV_X1 U8535 ( .A(n9704), .ZN(n9194) );
  OAI222_X1 U8536 ( .A1(n8222), .A2(n6955), .B1(n9550), .B2(n6956), .C1(
        P1_U3084), .C2(n9194), .ZN(P1_U3338) );
  INV_X1 U8537 ( .A(n8336), .ZN(n7919) );
  OAI222_X1 U8538 ( .A1(n7728), .A2(n6957), .B1(n8747), .B2(n6956), .C1(
        P2_U3152), .C2(n7919), .ZN(P2_U3343) );
  OAI21_X1 U8539 ( .B1(n6959), .B2(n6961), .A(n6958), .ZN(n6969) );
  XNOR2_X1 U8540 ( .A(n6961), .B(n6960), .ZN(n6963) );
  INV_X1 U8541 ( .A(n8585), .ZN(n8612) );
  AOI22_X1 U8542 ( .A1(n8591), .A2(n8328), .B1(n8326), .B2(n8590), .ZN(n6962)
         );
  OAI21_X1 U8543 ( .B1(n6963), .B2(n8612), .A(n6962), .ZN(n6964) );
  AOI21_X1 U8544 ( .B1(n8621), .B2(n6969), .A(n6964), .ZN(n7015) );
  OR2_X1 U8545 ( .A1(n6965), .A2(n6970), .ZN(n6966) );
  AND2_X1 U8546 ( .A1(n6967), .A2(n6966), .ZN(n7013) );
  INV_X1 U8547 ( .A(n7013), .ZN(n6968) );
  OAI22_X1 U8548 ( .A1(n8475), .A2(n6968), .B1(n8469), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n6972) );
  INV_X1 U8549 ( .A(n6969), .ZN(n7016) );
  OAI22_X1 U8550 ( .A1(n7016), .A2(n8629), .B1(n6970), .B2(n8626), .ZN(n6971)
         );
  AOI211_X1 U8551 ( .C1(P2_REG2_REG_3__SCAN_IN), .C2(n8600), .A(n6972), .B(
        n6971), .ZN(n6973) );
  OAI21_X1 U8552 ( .B1(n8600), .B2(n7015), .A(n6973), .ZN(P2_U3293) );
  AND2_X1 U8553 ( .A1(n6680), .A2(n7348), .ZN(n6976) );
  OAI21_X1 U8554 ( .B1(n9077), .B2(n6976), .A(n7048), .ZN(n7079) );
  INV_X1 U8555 ( .A(n6977), .ZN(n6979) );
  NAND2_X1 U8556 ( .A1(n6979), .A2(n6978), .ZN(n7063) );
  NOR2_X1 U8557 ( .A1(n7063), .A2(n7039), .ZN(n6980) );
  NAND2_X1 U8558 ( .A1(n7151), .A2(n6980), .ZN(n7290) );
  NAND2_X1 U8559 ( .A1(n9756), .A2(n7289), .ZN(n6981) );
  NOR2_X1 U8560 ( .A1(n6982), .A2(n9317), .ZN(n6983) );
  AND2_X1 U8561 ( .A1(n9379), .A2(n6983), .ZN(n7442) );
  OR2_X1 U8562 ( .A1(n6984), .A2(n9072), .ZN(n6986) );
  OR2_X1 U8563 ( .A1(n7346), .A2(n9106), .ZN(n6985) );
  AND2_X1 U8564 ( .A1(n6986), .A2(n6985), .ZN(n7815) );
  NAND2_X1 U8565 ( .A1(n9502), .A2(n6987), .ZN(n6988) );
  NOR2_X1 U8566 ( .A1(n6988), .A2(n7058), .ZN(n7076) );
  OAI22_X1 U8567 ( .A1(n9425), .A2(n6989), .B1(n6975), .B2(n7169), .ZN(n6990)
         );
  AOI21_X1 U8568 ( .B1(n7076), .B2(n9317), .A(n6990), .ZN(n6991) );
  OAI21_X1 U8569 ( .B1(n7079), .B2(n7815), .A(n6991), .ZN(n7000) );
  NOR2_X1 U8570 ( .A1(n6680), .A2(n7073), .ZN(n7068) );
  INV_X1 U8571 ( .A(n7068), .ZN(n6992) );
  XNOR2_X1 U8572 ( .A(n6992), .B(n9077), .ZN(n6995) );
  OR2_X1 U8573 ( .A1(n9071), .A2(n9317), .ZN(n6994) );
  NAND2_X1 U8574 ( .A1(n9140), .A2(n9148), .ZN(n6993) );
  NAND2_X1 U8575 ( .A1(n6995), .A2(n9433), .ZN(n6999) );
  AOI22_X1 U8576 ( .A1(n9437), .A2(n6680), .B1(n6719), .B2(n9438), .ZN(n6998)
         );
  NAND2_X1 U8577 ( .A1(n6999), .A2(n6998), .ZN(n7075) );
  NOR2_X1 U8578 ( .A1(n7000), .A2(n7075), .ZN(n7001) );
  MUX2_X1 U8579 ( .A(n7002), .B(n7001), .S(n9379), .Z(n7003) );
  OAI21_X1 U8580 ( .B1(n7079), .B2(n7822), .A(n7003), .ZN(P1_U3290) );
  INV_X1 U8581 ( .A(n7004), .ZN(n7005) );
  OAI222_X1 U8582 ( .A1(n7728), .A2(n10188), .B1(n8747), .B2(n7005), .C1(n4628), .C2(P2_U3152), .ZN(P2_U3342) );
  INV_X1 U8583 ( .A(n9715), .ZN(n9181) );
  OAI222_X1 U8584 ( .A1(n8222), .A2(n10131), .B1(n9550), .B2(n7005), .C1(n9181), .C2(P1_U3084), .ZN(P1_U3337) );
  NOR2_X4 U8585 ( .A1(n7027), .A2(n7009), .ZN(n9908) );
  INV_X1 U8586 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7018) );
  INV_X1 U8587 ( .A(n6393), .ZN(n7650) );
  AND2_X1 U8588 ( .A1(n7010), .A2(n9812), .ZN(n7011) );
  NAND2_X1 U8589 ( .A1(n7650), .A2(n7011), .ZN(n9883) );
  AOI22_X1 U8590 ( .A1(n7013), .A2(n9869), .B1(n9868), .B2(n7012), .ZN(n7014)
         );
  OAI211_X1 U8591 ( .C1(n7016), .C2(n9883), .A(n7015), .B(n7014), .ZN(n7028)
         );
  NAND2_X1 U8592 ( .A1(n7028), .A2(n9908), .ZN(n7017) );
  OAI21_X1 U8593 ( .B1(n9908), .B2(n7018), .A(n7017), .ZN(P2_U3460) );
  INV_X1 U8594 ( .A(n9848), .ZN(n7023) );
  AOI21_X1 U8595 ( .B1(n8626), .B2(n8475), .A(n7034), .ZN(n7021) );
  AOI22_X1 U8596 ( .A1(n9848), .A2(n8585), .B1(n8590), .B2(n6834), .ZN(n9850)
         );
  INV_X1 U8597 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7019) );
  OAI22_X1 U8598 ( .A1(n8600), .A2(n9850), .B1(n7019), .B2(n8469), .ZN(n7020)
         );
  AOI211_X1 U8599 ( .C1(n8600), .C2(P2_REG2_REG_0__SCAN_IN), .A(n7021), .B(
        n7020), .ZN(n7022) );
  OAI21_X1 U8600 ( .B1(n7023), .B2(n8606), .A(n7022), .ZN(P2_U3296) );
  INV_X1 U8601 ( .A(n7024), .ZN(n7067) );
  AOI22_X1 U8602 ( .A1(n9202), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9548), .ZN(n7025) );
  OAI21_X1 U8603 ( .B1(n7067), .B2(n9550), .A(n7025), .ZN(P1_U3336) );
  INV_X2 U8604 ( .A(n9919), .ZN(n9914) );
  NAND2_X1 U8605 ( .A1(n7028), .A2(n9914), .ZN(n7029) );
  OAI21_X1 U8606 ( .B1(n9914), .B2(n6586), .A(n7029), .ZN(P2_U3523) );
  MUX2_X1 U8607 ( .A(n7030), .B(n7034), .S(n8162), .Z(n7031) );
  AOI21_X1 U8608 ( .B1(n7032), .B2(n7031), .A(n8296), .ZN(n7036) );
  OAI22_X1 U8609 ( .A1(n8247), .A2(n7034), .B1(n7033), .B2(n8304), .ZN(n7035)
         );
  AOI211_X1 U8610 ( .C1(P2_REG3_REG_0__SCAN_IN), .C2(n7037), .A(n7036), .B(
        n7035), .ZN(n7038) );
  INV_X1 U8611 ( .A(n7038), .ZN(P2_U3234) );
  OAI21_X1 U8612 ( .B1(n9776), .B2(n9317), .A(n7039), .ZN(n7040) );
  NOR2_X4 U8613 ( .A1(n7064), .A2(n7042), .ZN(n9786) );
  AND4_X1 U8614 ( .A1(n7046), .A2(n7045), .A3(n7044), .A4(n7043), .ZN(n7369)
         );
  NAND2_X1 U8615 ( .A1(n7369), .A2(n6708), .ZN(n8913) );
  INV_X1 U8616 ( .A(n7156), .ZN(n7050) );
  AOI21_X1 U8617 ( .B1(n9075), .B2(n7049), .A(n7050), .ZN(n7361) );
  NAND2_X1 U8618 ( .A1(n9071), .A2(n7289), .ZN(n9070) );
  OR2_X1 U8619 ( .A1(n9070), .A2(n9148), .ZN(n9571) );
  INV_X1 U8620 ( .A(n9077), .ZN(n7051) );
  NAND2_X1 U8621 ( .A1(n7051), .A2(n7068), .ZN(n7054) );
  INV_X1 U8622 ( .A(n6974), .ZN(n7052) );
  NAND2_X1 U8623 ( .A1(n7054), .A2(n7053), .ZN(n7163) );
  XNOR2_X1 U8624 ( .A(n7163), .B(n9075), .ZN(n7057) );
  AOI22_X1 U8625 ( .A1(n9437), .A2(n6974), .B1(n7157), .B2(n9438), .ZN(n7055)
         );
  OAI21_X1 U8626 ( .B1(n7361), .B2(n7815), .A(n7055), .ZN(n7056) );
  AOI21_X1 U8627 ( .B1(n7057), .B2(n9433), .A(n7056), .ZN(n7365) );
  INV_X1 U8628 ( .A(n7058), .ZN(n7060) );
  NAND2_X1 U8629 ( .A1(n7058), .A2(n7357), .ZN(n7375) );
  INV_X1 U8630 ( .A(n7375), .ZN(n7059) );
  AOI21_X1 U8631 ( .B1(n6708), .B2(n7060), .A(n7059), .ZN(n7360) );
  AOI22_X1 U8632 ( .A1(n7360), .A2(n9502), .B1(n9564), .B2(n6708), .ZN(n7061)
         );
  OAI211_X1 U8633 ( .C1(n7361), .C2(n9571), .A(n7365), .B(n7061), .ZN(n7065)
         );
  NAND2_X1 U8634 ( .A1(n7065), .A2(n9786), .ZN(n7062) );
  OAI21_X1 U8635 ( .B1(n9528), .B2(n10041), .A(n7062), .ZN(P1_U3525) );
  NOR2_X4 U8636 ( .A1(n7064), .A2(n7063), .ZN(n9772) );
  NAND2_X1 U8637 ( .A1(n7065), .A2(n9783), .ZN(n7066) );
  OAI21_X1 U8638 ( .B1(n9772), .B2(n5037), .A(n7066), .ZN(P1_U3460) );
  OAI222_X1 U8639 ( .A1(n7728), .A2(n9999), .B1(n8747), .B2(n7067), .C1(n8357), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U8640 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9595) );
  AND2_X1 U8641 ( .A1(n6680), .A2(n7073), .ZN(n8909) );
  NOR2_X1 U8642 ( .A1(n7068), .A2(n8909), .ZN(n9076) );
  INV_X1 U8643 ( .A(n7161), .ZN(n7070) );
  INV_X1 U8644 ( .A(n7072), .ZN(n7069) );
  NOR3_X1 U8645 ( .A1(n9076), .A2(n7070), .A3(n7069), .ZN(n7071) );
  AOI21_X1 U8646 ( .B1(n9438), .B2(n6974), .A(n7071), .ZN(n7351) );
  OAI21_X1 U8647 ( .B1(n7073), .B2(n7072), .A(n7351), .ZN(n7083) );
  NAND2_X1 U8648 ( .A1(n7083), .A2(n9528), .ZN(n7074) );
  OAI21_X1 U8649 ( .B1(n9786), .B2(n9595), .A(n7074), .ZN(P1_U3523) );
  INV_X1 U8650 ( .A(n7075), .ZN(n7078) );
  OAI211_X1 U8651 ( .C1(n9526), .C2(n7079), .A(n7078), .B(n7077), .ZN(n7081)
         );
  NAND2_X1 U8652 ( .A1(n7081), .A2(n9528), .ZN(n7080) );
  OAI21_X1 U8653 ( .B1(n9528), .B2(n10155), .A(n7080), .ZN(P1_U3524) );
  NAND2_X1 U8654 ( .A1(n7081), .A2(n9772), .ZN(n7082) );
  OAI21_X1 U8655 ( .B1(n9772), .B2(n5018), .A(n7082), .ZN(P1_U3457) );
  NAND2_X1 U8656 ( .A1(n7083), .A2(n9772), .ZN(n7084) );
  OAI21_X1 U8657 ( .B1(n9772), .B2(n4963), .A(n7084), .ZN(P1_U3454) );
  NAND2_X1 U8658 ( .A1(n7262), .A2(n7085), .ZN(n7086) );
  NAND2_X1 U8659 ( .A1(n7087), .A2(n7086), .ZN(n7252) );
  NOR2_X1 U8660 ( .A1(n8325), .A2(n9807), .ZN(n7089) );
  OR2_X1 U8661 ( .A1(n7260), .A2(n7140), .ZN(n7088) );
  XNOR2_X1 U8662 ( .A(n7176), .B(n7175), .ZN(n9875) );
  XNOR2_X1 U8663 ( .A(n7090), .B(n7091), .ZN(n7094) );
  NAND2_X1 U8664 ( .A1(n8325), .A2(n8591), .ZN(n7092) );
  OAI21_X1 U8665 ( .B1(n7469), .B2(n8617), .A(n7092), .ZN(n7093) );
  AOI21_X1 U8666 ( .B1(n7094), .B2(n8585), .A(n7093), .ZN(n9878) );
  MUX2_X1 U8667 ( .A(n6571), .B(n9878), .S(n9817), .Z(n7098) );
  OAI21_X1 U8668 ( .B1(n7256), .B2(n9876), .A(n7185), .ZN(n9877) );
  OAI22_X1 U8669 ( .A1(n9877), .A2(n8475), .B1(n7095), .B2(n8469), .ZN(n7096)
         );
  AOI21_X1 U8670 ( .B1(n8473), .B2(n7177), .A(n7096), .ZN(n7097) );
  OAI211_X1 U8671 ( .C1(n8606), .C2(n9875), .A(n7098), .B(n7097), .ZN(P2_U3290) );
  OAI21_X1 U8672 ( .B1(n7101), .B2(n7099), .A(n7100), .ZN(n7102) );
  NAND2_X1 U8673 ( .A1(n7102), .A2(n8850), .ZN(n7109) );
  NAND2_X1 U8674 ( .A1(n8868), .A2(n9170), .ZN(n7104) );
  AND2_X1 U8675 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9617) );
  INV_X1 U8676 ( .A(n9617), .ZN(n7103) );
  OAI211_X1 U8677 ( .C1(n7478), .C2(n8865), .A(n7104), .B(n7103), .ZN(n7107)
         );
  INV_X1 U8678 ( .A(n7105), .ZN(n7167) );
  NOR2_X1 U8679 ( .A1(n8870), .A2(n7167), .ZN(n7106) );
  AOI211_X1 U8680 ( .C1(n8872), .C2(n4379), .A(n7107), .B(n7106), .ZN(n7108)
         );
  NAND2_X1 U8681 ( .A1(n7109), .A2(n7108), .ZN(P1_U3225) );
  NOR2_X1 U8682 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7625), .ZN(n7113) );
  AOI21_X1 U8683 ( .B1(n7115), .B2(P2_REG1_REG_10__SCAN_IN), .A(n7110), .ZN(
        n7270) );
  INV_X1 U8684 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7754) );
  MUX2_X1 U8685 ( .A(n7754), .B(P2_REG1_REG_11__SCAN_IN), .S(n7277), .Z(n7269)
         );
  XNOR2_X1 U8686 ( .A(n7270), .B(n7269), .ZN(n7111) );
  NOR2_X1 U8687 ( .A1(n9795), .A2(n7111), .ZN(n7112) );
  AOI211_X1 U8688 ( .C1(n9797), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n7113), .B(
        n7112), .ZN(n7121) );
  NOR2_X1 U8689 ( .A1(n7277), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7116) );
  AOI21_X1 U8690 ( .B1(n7277), .B2(P2_REG2_REG_11__SCAN_IN), .A(n7116), .ZN(
        n7117) );
  NAND2_X1 U8691 ( .A1(n7118), .A2(n7117), .ZN(n7276) );
  OAI21_X1 U8692 ( .B1(n7118), .B2(n7117), .A(n7276), .ZN(n7119) );
  NAND2_X1 U8693 ( .A1(n9791), .A2(n7119), .ZN(n7120) );
  OAI211_X1 U8694 ( .C1(n9794), .C2(n7272), .A(n7121), .B(n7120), .ZN(P2_U3256) );
  INV_X1 U8695 ( .A(n8305), .ZN(n8434) );
  NAND2_X1 U8696 ( .A1(n8434), .A2(P2_U3966), .ZN(n7122) );
  OAI21_X1 U8697 ( .B1(P2_U3966), .B2(n5711), .A(n7122), .ZN(P2_U3579) );
  INV_X1 U8698 ( .A(n7125), .ZN(n7128) );
  INV_X1 U8699 ( .A(n7126), .ZN(n7127) );
  NAND2_X1 U8700 ( .A1(n7128), .A2(n7127), .ZN(n7129) );
  OR2_X1 U8701 ( .A1(n7263), .A2(n8162), .ZN(n7131) );
  XNOR2_X1 U8702 ( .A(n7177), .B(n8152), .ZN(n7130) );
  NAND2_X1 U8703 ( .A1(n7131), .A2(n7130), .ZN(n7192) );
  OAI21_X1 U8704 ( .B1(n7131), .B2(n7130), .A(n7192), .ZN(n7133) );
  NAND2_X1 U8705 ( .A1(n7134), .A2(n7133), .ZN(n7135) );
  AOI21_X1 U8706 ( .B1(n7193), .B2(n7135), .A(n8296), .ZN(n7143) );
  OAI22_X1 U8707 ( .A1(n8247), .A2(n9876), .B1(n7469), .B2(n8304), .ZN(n7142)
         );
  INV_X1 U8708 ( .A(n7136), .ZN(n7139) );
  NAND2_X1 U8709 ( .A1(n8293), .A2(n7137), .ZN(n7138) );
  OAI211_X1 U8710 ( .C1(n8302), .C2(n7140), .A(n7139), .B(n7138), .ZN(n7141)
         );
  OR3_X1 U8711 ( .A1(n7143), .A2(n7142), .A3(n7141), .ZN(P2_U3241) );
  NAND2_X1 U8712 ( .A1(n4461), .A2(n7145), .ZN(n7146) );
  XNOR2_X1 U8713 ( .A(n7144), .B(n7146), .ZN(n7154) );
  INV_X1 U8714 ( .A(n8868), .ZN(n8853) );
  NOR2_X1 U8715 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10071), .ZN(n9633) );
  AOI21_X1 U8716 ( .B1(n8857), .B2(n9167), .A(n9633), .ZN(n7148) );
  NAND2_X1 U8717 ( .A1(n8819), .A2(n4472), .ZN(n7147) );
  OAI211_X1 U8718 ( .C1(n8853), .C2(n7311), .A(n7148), .B(n7147), .ZN(n7149)
         );
  INV_X1 U8719 ( .A(n7149), .ZN(n7153) );
  AND2_X1 U8720 ( .A1(n9564), .A2(n4383), .ZN(n9765) );
  NAND3_X1 U8721 ( .A1(n9765), .A2(n7151), .A3(n7150), .ZN(n7152) );
  OAI211_X1 U8722 ( .C1(n7154), .C2(n8874), .A(n7153), .B(n7152), .ZN(P1_U3237) );
  INV_X1 U8723 ( .A(n7213), .ZN(n7202) );
  NAND2_X1 U8724 ( .A1(n9169), .A2(n7202), .ZN(n9111) );
  AND2_X1 U8725 ( .A1(n7308), .A2(n9111), .ZN(n9082) );
  NAND2_X1 U8726 ( .A1(n7369), .A2(n7357), .ZN(n7155) );
  NAND2_X1 U8727 ( .A1(n7156), .A2(n7155), .ZN(n7367) );
  NAND2_X1 U8728 ( .A1(n7238), .A2(n7380), .ZN(n8916) );
  INV_X1 U8729 ( .A(n7380), .ZN(n9759) );
  NAND2_X1 U8730 ( .A1(n7157), .A2(n9759), .ZN(n7239) );
  NAND2_X1 U8731 ( .A1(n8916), .A2(n7239), .ZN(n9078) );
  NAND2_X1 U8732 ( .A1(n7367), .A2(n9078), .ZN(n7366) );
  NAND2_X1 U8733 ( .A1(n7238), .A2(n9759), .ZN(n7158) );
  NAND2_X1 U8734 ( .A1(n7366), .A2(n7158), .ZN(n7237) );
  NAND2_X1 U8735 ( .A1(n7368), .A2(n7246), .ZN(n7222) );
  NAND2_X1 U8736 ( .A1(n9170), .A2(n7436), .ZN(n9110) );
  NAND2_X1 U8737 ( .A1(n7222), .A2(n9110), .ZN(n9079) );
  NAND2_X1 U8738 ( .A1(n7237), .A2(n9079), .ZN(n7236) );
  NAND2_X1 U8739 ( .A1(n7368), .A2(n7436), .ZN(n7159) );
  NAND2_X1 U8740 ( .A1(n7236), .A2(n7159), .ZN(n7210) );
  OR2_X1 U8741 ( .A1(n7210), .A2(n9082), .ZN(n7314) );
  INV_X1 U8742 ( .A(n7314), .ZN(n7160) );
  AOI21_X1 U8743 ( .B1(n9082), .B2(n7210), .A(n7160), .ZN(n7205) );
  INV_X1 U8744 ( .A(n7205), .ZN(n7173) );
  INV_X2 U8745 ( .A(n9404), .ZN(n9379) );
  AND2_X1 U8746 ( .A1(n7161), .A2(n5049), .ZN(n7162) );
  NAND2_X1 U8747 ( .A1(n7163), .A2(n9075), .ZN(n7164) );
  INV_X1 U8748 ( .A(n8916), .ZN(n9113) );
  AND2_X1 U8749 ( .A1(n7239), .A2(n9110), .ZN(n7221) );
  NAND2_X1 U8750 ( .A1(n7165), .A2(n7222), .ZN(n7307) );
  XOR2_X1 U8751 ( .A(n9082), .B(n7307), .Z(n7166) );
  OAI222_X1 U8752 ( .A1(n9371), .A2(n7478), .B1(n9369), .B2(n7368), .C1(n7166), 
        .C2(n9389), .ZN(n7203) );
  OAI211_X1 U8753 ( .C1(n7245), .C2(n7202), .A(n7317), .B(n9502), .ZN(n7201)
         );
  OAI22_X1 U8754 ( .A1(n7201), .A2(n7289), .B1(n9425), .B2(n7167), .ZN(n7168)
         );
  OAI21_X1 U8755 ( .B1(n7203), .B2(n7168), .A(n9379), .ZN(n7172) );
  INV_X1 U8756 ( .A(n7169), .ZN(n7170) );
  AOI22_X1 U8757 ( .A1(n9321), .A2(n4379), .B1(P1_REG2_REG_5__SCAN_IN), .B2(
        n9404), .ZN(n7171) );
  OAI211_X1 U8758 ( .C1(n7173), .C2(n9444), .A(n7172), .B(n7171), .ZN(P1_U3286) );
  NAND2_X1 U8759 ( .A1(n9282), .A2(P1_U4006), .ZN(n7174) );
  OAI21_X1 U8760 ( .B1(P1_U4006), .B2(n8006), .A(n7174), .ZN(P1_U3582) );
  NAND2_X1 U8761 ( .A1(n7176), .A2(n7175), .ZN(n7179) );
  NAND2_X1 U8762 ( .A1(n8324), .A2(n7177), .ZN(n7178) );
  XNOR2_X1 U8763 ( .A(n7386), .B(n7180), .ZN(n7302) );
  XNOR2_X1 U8764 ( .A(n7182), .B(n7385), .ZN(n7183) );
  INV_X1 U8765 ( .A(n7706), .ZN(n8322) );
  AOI222_X1 U8766 ( .A1(n8585), .A2(n7183), .B1(n8322), .B2(n8590), .C1(n8324), 
        .C2(n8591), .ZN(n7301) );
  OR2_X1 U8767 ( .A1(n7301), .A2(n8600), .ZN(n7191) );
  INV_X1 U8768 ( .A(n7396), .ZN(n7184) );
  AOI21_X1 U8769 ( .B1(n7384), .B2(n7185), .A(n7184), .ZN(n7299) );
  INV_X1 U8770 ( .A(n7384), .ZN(n7196) );
  NOR2_X1 U8771 ( .A1(n8626), .A2(n7196), .ZN(n7189) );
  INV_X1 U8772 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7187) );
  INV_X1 U8773 ( .A(n7194), .ZN(n7186) );
  OAI22_X1 U8774 ( .A1(n9817), .A2(n7187), .B1(n7186), .B2(n8469), .ZN(n7188)
         );
  AOI211_X1 U8775 ( .C1(n7299), .C2(n8632), .A(n7189), .B(n7188), .ZN(n7190)
         );
  OAI211_X1 U8776 ( .C1(n8606), .C2(n7302), .A(n7191), .B(n7190), .ZN(P2_U3289) );
  XNOR2_X1 U8777 ( .A(n7384), .B(n8163), .ZN(n7460) );
  NOR2_X1 U8778 ( .A1(n7469), .A2(n8162), .ZN(n7461) );
  XNOR2_X1 U8779 ( .A(n7460), .B(n7461), .ZN(n7464) );
  XNOR2_X1 U8780 ( .A(n7465), .B(n7464), .ZN(n7200) );
  NAND2_X1 U8781 ( .A1(n8293), .A2(n7194), .ZN(n7195) );
  OAI21_X1 U8782 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n5930), .A(n7195), .ZN(n7198) );
  OAI22_X1 U8783 ( .A1(n8247), .A2(n7196), .B1(n7706), .B2(n8304), .ZN(n7197)
         );
  AOI211_X1 U8784 ( .C1(n8280), .C2(n8324), .A(n7198), .B(n7197), .ZN(n7199)
         );
  OAI21_X1 U8785 ( .B1(n7200), .B2(n8296), .A(n7199), .ZN(P2_U3215) );
  INV_X1 U8786 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7207) );
  OAI21_X1 U8787 ( .B1(n7202), .B2(n9774), .A(n7201), .ZN(n7204) );
  AOI211_X1 U8788 ( .C1(n7205), .C2(n9771), .A(n7204), .B(n7203), .ZN(n7208)
         );
  OR2_X1 U8789 ( .A1(n7208), .A2(n9787), .ZN(n7206) );
  OAI21_X1 U8790 ( .B1(n9528), .B2(n7207), .A(n7206), .ZN(P1_U3528) );
  OR2_X1 U8791 ( .A1(n7208), .A2(n9782), .ZN(n7209) );
  OAI21_X1 U8792 ( .B1(n9772), .B2(n5115), .A(n7209), .ZN(P1_U3469) );
  INV_X1 U8793 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7232) );
  INV_X1 U8794 ( .A(n7210), .ZN(n7212) );
  AND2_X1 U8795 ( .A1(n7478), .A2(n4382), .ZN(n7214) );
  NAND2_X1 U8796 ( .A1(n7212), .A2(n4432), .ZN(n7217) );
  NAND2_X1 U8797 ( .A1(n7478), .A2(n7211), .ZN(n8969) );
  NAND2_X1 U8798 ( .A1(n9168), .A2(n4382), .ZN(n9117) );
  NAND2_X1 U8799 ( .A1(n8969), .A2(n9117), .ZN(n8973) );
  NAND2_X1 U8800 ( .A1(n9169), .A2(n4379), .ZN(n7312) );
  AND2_X1 U8801 ( .A1(n8973), .A2(n7312), .ZN(n7313) );
  OR2_X1 U8802 ( .A1(n7214), .A2(n7313), .ZN(n7215) );
  AND2_X1 U8803 ( .A1(n7217), .A2(n7215), .ZN(n7218) );
  NAND2_X1 U8804 ( .A1(n7694), .A2(n7485), .ZN(n8968) );
  INV_X1 U8805 ( .A(n7485), .ZN(n7328) );
  NAND2_X1 U8806 ( .A1(n7328), .A2(n9167), .ZN(n8972) );
  NAND2_X1 U8807 ( .A1(n8968), .A2(n8972), .ZN(n7226) );
  AND2_X1 U8808 ( .A1(n7226), .A2(n7215), .ZN(n7216) );
  OAI21_X1 U8809 ( .B1(n7218), .B2(n7226), .A(n7330), .ZN(n7219) );
  INV_X1 U8810 ( .A(n7219), .ZN(n7298) );
  NAND2_X1 U8811 ( .A1(n9117), .A2(n9111), .ZN(n7220) );
  NAND2_X1 U8812 ( .A1(n8969), .A2(n7220), .ZN(n7223) );
  NAND2_X1 U8813 ( .A1(n7240), .A2(n9120), .ZN(n7227) );
  NAND2_X1 U8814 ( .A1(n8969), .A2(n7308), .ZN(n9114) );
  INV_X1 U8815 ( .A(n7222), .ZN(n9112) );
  OR2_X1 U8816 ( .A1(n9114), .A2(n9112), .ZN(n7224) );
  NAND2_X1 U8817 ( .A1(n7224), .A2(n7223), .ZN(n8919) );
  NAND2_X1 U8818 ( .A1(n7227), .A2(n8919), .ZN(n7225) );
  INV_X1 U8819 ( .A(n7226), .ZN(n9081) );
  NAND2_X1 U8820 ( .A1(n7225), .A2(n9081), .ZN(n7402) );
  NAND3_X1 U8821 ( .A1(n7227), .A2(n8919), .A3(n7226), .ZN(n7228) );
  NAND2_X1 U8822 ( .A1(n7402), .A2(n7228), .ZN(n7229) );
  AOI222_X1 U8823 ( .A1(n9433), .A2(n7229), .B1(n9166), .B2(n9438), .C1(n9168), 
        .C2(n9437), .ZN(n7293) );
  AOI211_X1 U8824 ( .C1(n7485), .C2(n7318), .A(n9776), .B(n7412), .ZN(n7296)
         );
  AOI21_X1 U8825 ( .B1(n9564), .B2(n7485), .A(n7296), .ZN(n7230) );
  OAI211_X1 U8826 ( .C1(n7298), .C2(n9526), .A(n7293), .B(n7230), .ZN(n7233)
         );
  NAND2_X1 U8827 ( .A1(n7233), .A2(n9786), .ZN(n7231) );
  OAI21_X1 U8828 ( .B1(n9528), .B2(n7232), .A(n7231), .ZN(P1_U3530) );
  INV_X1 U8829 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7235) );
  NAND2_X1 U8830 ( .A1(n7233), .A2(n9783), .ZN(n7234) );
  OAI21_X1 U8831 ( .B1(n9772), .B2(n7235), .A(n7234), .ZN(P1_U3475) );
  OAI21_X1 U8832 ( .B1(n7237), .B2(n9079), .A(n7236), .ZN(n7443) );
  INV_X1 U8833 ( .A(n7443), .ZN(n7248) );
  INV_X1 U8834 ( .A(n7815), .ZN(n7371) );
  OAI22_X1 U8835 ( .A1(n7238), .A2(n9369), .B1(n7311), .B2(n9371), .ZN(n7244)
         );
  NAND2_X1 U8836 ( .A1(n7240), .A2(n7239), .ZN(n7241) );
  XOR2_X1 U8837 ( .A(n9079), .B(n7241), .Z(n7242) );
  NOR2_X1 U8838 ( .A1(n7242), .A2(n9389), .ZN(n7243) );
  AOI211_X1 U8839 ( .C1(n7371), .C2(n7443), .A(n7244), .B(n7243), .ZN(n7446)
         );
  AOI21_X1 U8840 ( .B1(n7246), .B2(n7377), .A(n7245), .ZN(n7441) );
  AOI22_X1 U8841 ( .A1(n7441), .A2(n9502), .B1(n9564), .B2(n7246), .ZN(n7247)
         );
  OAI211_X1 U8842 ( .C1(n7248), .C2(n9571), .A(n7446), .B(n7247), .ZN(n7250)
         );
  NAND2_X1 U8843 ( .A1(n7250), .A2(n9772), .ZN(n7249) );
  OAI21_X1 U8844 ( .B1(n9772), .B2(n5100), .A(n7249), .ZN(P1_U3466) );
  NAND2_X1 U8845 ( .A1(n7250), .A2(n9528), .ZN(n7251) );
  OAI21_X1 U8846 ( .B1(n9528), .B2(n10106), .A(n7251), .ZN(P1_U3527) );
  INV_X1 U8847 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7266) );
  XOR2_X1 U8848 ( .A(n7260), .B(n7252), .Z(n9803) );
  NAND2_X1 U8849 ( .A1(n7253), .A2(n9807), .ZN(n7254) );
  NAND2_X1 U8850 ( .A1(n7254), .A2(n9869), .ZN(n7255) );
  NOR2_X1 U8851 ( .A1(n7256), .A2(n7255), .ZN(n9806) );
  NAND2_X1 U8852 ( .A1(n7257), .A2(n7258), .ZN(n7259) );
  XOR2_X1 U8853 ( .A(n7260), .B(n7259), .Z(n7261) );
  OAI222_X1 U8854 ( .A1(n8617), .A2(n7263), .B1(n8615), .B2(n7262), .C1(n8612), 
        .C2(n7261), .ZN(n9815) );
  AOI211_X1 U8855 ( .C1(n9868), .C2(n9807), .A(n9806), .B(n9815), .ZN(n7264)
         );
  OAI21_X1 U8856 ( .B1(n8720), .B2(n9803), .A(n7264), .ZN(n7267) );
  NAND2_X1 U8857 ( .A1(n7267), .A2(n9908), .ZN(n7265) );
  OAI21_X1 U8858 ( .B1(n9908), .B2(n7266), .A(n7265), .ZN(P2_U3466) );
  NAND2_X1 U8859 ( .A1(n7267), .A2(n9914), .ZN(n7268) );
  OAI21_X1 U8860 ( .B1(n9914), .B2(n6579), .A(n7268), .ZN(P2_U3525) );
  INV_X1 U8861 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9920) );
  AOI22_X1 U8862 ( .A1(n7427), .A2(n9920), .B1(P2_REG1_REG_12__SCAN_IN), .B2(
        n7422), .ZN(n7274) );
  OR2_X1 U8863 ( .A1(n7270), .A2(n7269), .ZN(n7271) );
  OAI21_X1 U8864 ( .B1(n7754), .B2(n7272), .A(n7271), .ZN(n7273) );
  NOR2_X1 U8865 ( .A1(n7274), .A2(n7273), .ZN(n7421) );
  AOI21_X1 U8866 ( .B1(n7274), .B2(n7273), .A(n7421), .ZN(n7284) );
  NOR2_X1 U8867 ( .A1(n7427), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7275) );
  AOI21_X1 U8868 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7427), .A(n7275), .ZN(
        n7279) );
  OAI21_X1 U8869 ( .B1(n7277), .B2(P2_REG2_REG_11__SCAN_IN), .A(n7276), .ZN(
        n7278) );
  NAND2_X1 U8870 ( .A1(n7279), .A2(n7278), .ZN(n7426) );
  OAI21_X1 U8871 ( .B1(n7279), .B2(n7278), .A(n7426), .ZN(n7280) );
  NAND2_X1 U8872 ( .A1(n7280), .A2(n9791), .ZN(n7283) );
  INV_X1 U8873 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n10152) );
  NAND2_X1 U8874 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7737) );
  OAI21_X1 U8875 ( .B1(n8388), .B2(n10152), .A(n7737), .ZN(n7281) );
  AOI21_X1 U8876 ( .B1(n8384), .B2(n7427), .A(n7281), .ZN(n7282) );
  OAI211_X1 U8877 ( .C1(n7284), .C2(n9795), .A(n7283), .B(n7282), .ZN(P2_U3257) );
  INV_X1 U8878 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7286) );
  INV_X1 U8879 ( .A(n7285), .ZN(n7287) );
  INV_X1 U8880 ( .A(n9205), .ZN(n9744) );
  OAI222_X1 U8881 ( .A1(n8222), .A2(n7286), .B1(n9550), .B2(n7287), .C1(
        P1_U3084), .C2(n9744), .ZN(P1_U3335) );
  INV_X1 U8882 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7288) );
  INV_X1 U8883 ( .A(n8367), .ZN(n8373) );
  OAI222_X1 U8884 ( .A1(n7728), .A2(n7288), .B1(n8747), .B2(n7287), .C1(
        P2_U3152), .C2(n8373), .ZN(P2_U3340) );
  NOR2_X1 U8885 ( .A1(n7290), .A2(n7289), .ZN(n9430) );
  INV_X1 U8886 ( .A(n7291), .ZN(n7475) );
  INV_X1 U8887 ( .A(n9425), .ZN(n9402) );
  AOI22_X1 U8888 ( .A1(n9404), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7475), .B2(
        n9402), .ZN(n7292) );
  OAI21_X1 U8889 ( .B1(n7328), .B2(n9423), .A(n7292), .ZN(n7295) );
  NOR2_X1 U8890 ( .A1(n7293), .A2(n9404), .ZN(n7294) );
  AOI211_X1 U8891 ( .C1(n7296), .C2(n9430), .A(n7295), .B(n7294), .ZN(n7297)
         );
  OAI21_X1 U8892 ( .B1(n7298), .B2(n9444), .A(n7297), .ZN(P1_U3284) );
  INV_X1 U8893 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7304) );
  AOI22_X1 U8894 ( .A1(n7299), .A2(n9869), .B1(n9868), .B2(n7384), .ZN(n7300)
         );
  OAI211_X1 U8895 ( .C1(n8720), .C2(n7302), .A(n7301), .B(n7300), .ZN(n7305)
         );
  NAND2_X1 U8896 ( .A1(n7305), .A2(n9908), .ZN(n7303) );
  OAI21_X1 U8897 ( .B1(n9908), .B2(n7304), .A(n7303), .ZN(P2_U3472) );
  NAND2_X1 U8898 ( .A1(n7305), .A2(n9914), .ZN(n7306) );
  OAI21_X1 U8899 ( .B1(n9914), .B2(n6592), .A(n7306), .ZN(P2_U3527) );
  NAND2_X1 U8900 ( .A1(n7307), .A2(n9082), .ZN(n7309) );
  NAND2_X1 U8901 ( .A1(n7309), .A2(n7308), .ZN(n8974) );
  XNOR2_X1 U8902 ( .A(n8974), .B(n8973), .ZN(n7310) );
  OAI222_X1 U8903 ( .A1(n9371), .A2(n7694), .B1(n9369), .B2(n7311), .C1(n7310), 
        .C2(n9389), .ZN(n9768) );
  INV_X1 U8904 ( .A(n9768), .ZN(n7327) );
  AND2_X1 U8905 ( .A1(n7314), .A2(n7312), .ZN(n7316) );
  NAND2_X1 U8906 ( .A1(n7314), .A2(n7313), .ZN(n7315) );
  OAI21_X1 U8907 ( .B1(n7316), .B2(n8973), .A(n7315), .ZN(n9770) );
  INV_X1 U8908 ( .A(n9444), .ZN(n7325) );
  AOI21_X1 U8909 ( .B1(n7317), .B2(n4383), .A(n9776), .ZN(n7319) );
  NAND2_X1 U8910 ( .A1(n7319), .A2(n7318), .ZN(n9767) );
  INV_X1 U8911 ( .A(n9430), .ZN(n7323) );
  OAI22_X1 U8912 ( .A1(n9379), .A2(n6433), .B1(n7320), .B2(n9425), .ZN(n7321)
         );
  AOI21_X1 U8913 ( .B1(n9321), .B2(n4383), .A(n7321), .ZN(n7322) );
  OAI21_X1 U8914 ( .B1(n9767), .B2(n7323), .A(n7322), .ZN(n7324) );
  AOI21_X1 U8915 ( .B1(n9770), .B2(n7325), .A(n7324), .ZN(n7326) );
  OAI21_X1 U8916 ( .B1(n7327), .B2(n9404), .A(n7326), .ZN(P1_U3285) );
  NAND2_X1 U8917 ( .A1(n7694), .A2(n7328), .ZN(n7329) );
  INV_X1 U8918 ( .A(n9166), .ZN(n7778) );
  OR2_X1 U8919 ( .A1(n7778), .A2(n7702), .ZN(n8924) );
  NAND2_X1 U8920 ( .A1(n7702), .A2(n7778), .ZN(n8983) );
  NAND2_X1 U8921 ( .A1(n7702), .A2(n9166), .ZN(n7332) );
  NAND2_X1 U8922 ( .A1(n7407), .A2(n7332), .ZN(n7448) );
  OR2_X1 U8923 ( .A1(n7784), .A2(n9165), .ZN(n7334) );
  AND2_X1 U8924 ( .A1(n7784), .A2(n9165), .ZN(n7333) );
  INV_X1 U8925 ( .A(n9164), .ZN(n7594) );
  NAND2_X1 U8926 ( .A1(n7664), .A2(n7594), .ZN(n8988) );
  NAND2_X1 U8927 ( .A1(n7592), .A2(n8988), .ZN(n9087) );
  OAI21_X1 U8928 ( .B1(n7335), .B2(n9087), .A(n7585), .ZN(n7336) );
  INV_X1 U8929 ( .A(n7336), .ZN(n7515) );
  INV_X1 U8930 ( .A(n7702), .ZN(n7411) );
  INV_X1 U8931 ( .A(n7784), .ZN(n9775) );
  NAND2_X1 U8932 ( .A1(n7453), .A2(n9775), .ZN(n7455) );
  INV_X1 U8933 ( .A(n7599), .ZN(n7337) );
  AOI211_X1 U8934 ( .C1(n7664), .C2(n7455), .A(n9776), .B(n7337), .ZN(n7513)
         );
  INV_X1 U8935 ( .A(n7664), .ZN(n7338) );
  NOR2_X1 U8936 ( .A1(n7338), .A2(n9423), .ZN(n7341) );
  OAI22_X1 U8937 ( .A1(n9379), .A2(n7339), .B1(n7662), .B2(n9425), .ZN(n7340)
         );
  AOI211_X1 U8938 ( .C1(n7513), .C2(n9430), .A(n7341), .B(n7340), .ZN(n7345)
         );
  INV_X1 U8939 ( .A(n9165), .ZN(n7404) );
  AND2_X1 U8940 ( .A1(n8983), .A2(n8968), .ZN(n8975) );
  OR2_X1 U8941 ( .A1(n7784), .A2(n7404), .ZN(n7589) );
  INV_X1 U8942 ( .A(n7589), .ZN(n7447) );
  AND2_X1 U8943 ( .A1(n7784), .A2(n7404), .ZN(n7591) );
  INV_X1 U8944 ( .A(n7591), .ZN(n8984) );
  OAI21_X1 U8945 ( .B1(n7590), .B2(n7447), .A(n8984), .ZN(n7342) );
  XNOR2_X1 U8946 ( .A(n7342), .B(n9087), .ZN(n7343) );
  OAI222_X1 U8947 ( .A1(n9371), .A2(n7658), .B1(n9369), .B2(n7404), .C1(n7343), 
        .C2(n9389), .ZN(n7512) );
  NAND2_X1 U8948 ( .A1(n7512), .A2(n9379), .ZN(n7344) );
  OAI211_X1 U8949 ( .C1(n7515), .C2(n9444), .A(n7345), .B(n7344), .ZN(P1_U3281) );
  AOI22_X1 U8950 ( .A1(n9404), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n9402), .ZN(n7350) );
  NOR2_X1 U8951 ( .A1(n7346), .A2(n9140), .ZN(n7347) );
  NAND2_X1 U8952 ( .A1(n9379), .A2(n7347), .ZN(n9247) );
  OAI21_X1 U8953 ( .B1(n9414), .B2(n9321), .A(n7348), .ZN(n7349) );
  OAI211_X1 U8954 ( .C1(n7351), .C2(n9404), .A(n7350), .B(n7349), .ZN(P1_U3291) );
  INV_X1 U8955 ( .A(n7352), .ZN(n7354) );
  OAI222_X1 U8956 ( .A1(n7728), .A2(n7353), .B1(n8747), .B2(n7354), .C1(
        P2_U3152), .C2(n6227), .ZN(P2_U3339) );
  OAI222_X1 U8957 ( .A1(n8222), .A2(n7355), .B1(n9550), .B2(n7354), .C1(n9317), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  INV_X1 U8958 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7356) );
  OAI22_X1 U8959 ( .A1(n9379), .A2(n9961), .B1(n7356), .B2(n9425), .ZN(n7359)
         );
  NOR2_X1 U8960 ( .A1(n9423), .A2(n7357), .ZN(n7358) );
  AOI211_X1 U8961 ( .C1(n7360), .C2(n9414), .A(n7359), .B(n7358), .ZN(n7364)
         );
  INV_X1 U8962 ( .A(n7361), .ZN(n7362) );
  NAND2_X1 U8963 ( .A1(n7362), .A2(n7442), .ZN(n7363) );
  OAI211_X1 U8964 ( .C1(n7365), .C2(n9404), .A(n7364), .B(n7363), .ZN(P1_U3289) );
  OAI21_X1 U8965 ( .B1(n7367), .B2(n9078), .A(n7366), .ZN(n9763) );
  INV_X1 U8966 ( .A(n9763), .ZN(n7383) );
  XNOR2_X1 U8967 ( .A(n9119), .B(n9078), .ZN(n7373) );
  OAI22_X1 U8968 ( .A1(n7369), .A2(n9369), .B1(n7368), .B2(n9371), .ZN(n7370)
         );
  AOI21_X1 U8969 ( .B1(n9763), .B2(n7371), .A(n7370), .ZN(n7372) );
  OAI21_X1 U8970 ( .B1(n9389), .B2(n7373), .A(n7372), .ZN(n9761) );
  NAND2_X1 U8971 ( .A1(n9761), .A2(n9379), .ZN(n7382) );
  OAI22_X1 U8972 ( .A1(n9379), .A2(n7374), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9425), .ZN(n7379) );
  NAND2_X1 U8973 ( .A1(n7375), .A2(n7380), .ZN(n7376) );
  NAND2_X1 U8974 ( .A1(n7377), .A2(n7376), .ZN(n9760) );
  NOR2_X1 U8975 ( .A1(n9247), .A2(n9760), .ZN(n7378) );
  AOI211_X1 U8976 ( .C1(n9321), .C2(n7380), .A(n7379), .B(n7378), .ZN(n7381)
         );
  OAI211_X1 U8977 ( .C1(n7383), .C2(n7822), .A(n7382), .B(n7381), .ZN(P1_U3288) );
  INV_X1 U8978 ( .A(n7469), .ZN(n8323) );
  NAND2_X1 U8979 ( .A1(n7387), .A2(n7391), .ZN(n7388) );
  NAND2_X1 U8980 ( .A1(n7632), .A2(n7388), .ZN(n9884) );
  OAI21_X1 U8981 ( .B1(n7391), .B2(n7390), .A(n7389), .ZN(n7393) );
  OAI22_X1 U8982 ( .A1(n7469), .A2(n8615), .B1(n7638), .B2(n8617), .ZN(n7392)
         );
  AOI21_X1 U8983 ( .B1(n7393), .B2(n8585), .A(n7392), .ZN(n7394) );
  OAI21_X1 U8984 ( .B1(n9884), .B2(n9805), .A(n7394), .ZN(n9887) );
  NAND2_X1 U8985 ( .A1(n9887), .A2(n9817), .ZN(n7401) );
  OAI22_X1 U8986 ( .A1(n9817), .A2(n6624), .B1(n7395), .B2(n8469), .ZN(n7399)
         );
  OR2_X2 U8987 ( .A1(n7396), .A2(n7630), .ZN(n7715) );
  NAND2_X1 U8988 ( .A1(n7396), .A2(n7630), .ZN(n7397) );
  NAND2_X1 U8989 ( .A1(n7715), .A2(n7397), .ZN(n9886) );
  NOR2_X1 U8990 ( .A1(n9886), .A2(n8475), .ZN(n7398) );
  AOI211_X1 U8991 ( .C1(n8473), .C2(n7630), .A(n7399), .B(n7398), .ZN(n7400)
         );
  OAI211_X1 U8992 ( .C1(n9884), .C2(n8629), .A(n7401), .B(n7400), .ZN(P2_U3288) );
  NAND2_X1 U8993 ( .A1(n7402), .A2(n8968), .ZN(n7403) );
  XNOR2_X1 U8994 ( .A(n7403), .B(n9085), .ZN(n7410) );
  OAI22_X1 U8995 ( .A1(n7694), .A2(n9369), .B1(n7404), .B2(n9371), .ZN(n7409)
         );
  NAND2_X1 U8996 ( .A1(n7405), .A2(n9085), .ZN(n7406) );
  NAND2_X1 U8997 ( .A1(n7407), .A2(n7406), .ZN(n7549) );
  NOR2_X1 U8998 ( .A1(n7549), .A2(n7815), .ZN(n7408) );
  AOI211_X1 U8999 ( .C1(n7410), .C2(n9433), .A(n7409), .B(n7408), .ZN(n7548)
         );
  INV_X1 U9000 ( .A(n7549), .ZN(n7419) );
  NOR2_X1 U9001 ( .A1(n7412), .A2(n7411), .ZN(n7413) );
  OR2_X1 U9002 ( .A1(n7453), .A2(n7413), .ZN(n7545) );
  INV_X1 U9003 ( .A(n7691), .ZN(n7414) );
  OAI22_X1 U9004 ( .A1(n9379), .A2(n7415), .B1(n7414), .B2(n9425), .ZN(n7416)
         );
  AOI21_X1 U9005 ( .B1(n9321), .B2(n7702), .A(n7416), .ZN(n7417) );
  OAI21_X1 U9006 ( .B1(n7545), .B2(n9247), .A(n7417), .ZN(n7418) );
  AOI21_X1 U9007 ( .B1(n7419), .B2(n7442), .A(n7418), .ZN(n7420) );
  OAI21_X1 U9008 ( .B1(n7548), .B2(n9404), .A(n7420), .ZN(P1_U3283) );
  AOI21_X1 U9009 ( .B1(n7422), .B2(n9920), .A(n7421), .ZN(n7424) );
  INV_X1 U9010 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7522) );
  AOI22_X1 U9011 ( .A1(n7528), .A2(n7522), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7523), .ZN(n7423) );
  NOR2_X1 U9012 ( .A1(n7424), .A2(n7423), .ZN(n7521) );
  AOI21_X1 U9013 ( .B1(n7424), .B2(n7423), .A(n7521), .ZN(n7435) );
  INV_X1 U9014 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7425) );
  AOI22_X1 U9015 ( .A1(n7528), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7425), .B2(
        n7523), .ZN(n7429) );
  OAI21_X1 U9016 ( .B1(n7429), .B2(n7428), .A(n7527), .ZN(n7430) );
  NAND2_X1 U9017 ( .A1(n7430), .A2(n9791), .ZN(n7434) );
  INV_X1 U9018 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7431) );
  NAND2_X1 U9019 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7768) );
  OAI21_X1 U9020 ( .B1(n8388), .B2(n7431), .A(n7768), .ZN(n7432) );
  AOI21_X1 U9021 ( .B1(n8384), .B2(n7528), .A(n7432), .ZN(n7433) );
  OAI211_X1 U9022 ( .C1(n7435), .C2(n9795), .A(n7434), .B(n7433), .ZN(P2_U3258) );
  NOR2_X1 U9023 ( .A1(n9423), .A2(n7436), .ZN(n7440) );
  OAI22_X1 U9024 ( .A1(n9379), .A2(n7438), .B1(n7437), .B2(n9425), .ZN(n7439)
         );
  AOI211_X1 U9025 ( .C1(n7441), .C2(n9414), .A(n7440), .B(n7439), .ZN(n7445)
         );
  NAND2_X1 U9026 ( .A1(n7443), .A2(n7442), .ZN(n7444) );
  OAI211_X1 U9027 ( .C1(n7446), .C2(n9404), .A(n7445), .B(n7444), .ZN(P1_U3287) );
  XNOR2_X1 U9028 ( .A(n7448), .B(n9086), .ZN(n9773) );
  XNOR2_X1 U9029 ( .A(n7590), .B(n9086), .ZN(n7450) );
  OAI22_X1 U9030 ( .A1(n7594), .A2(n9371), .B1(n7778), .B2(n9369), .ZN(n7449)
         );
  AOI21_X1 U9031 ( .B1(n7450), .B2(n9433), .A(n7449), .ZN(n7451) );
  OAI21_X1 U9032 ( .B1(n9773), .B2(n7815), .A(n7451), .ZN(n9778) );
  NAND2_X1 U9033 ( .A1(n9778), .A2(n9379), .ZN(n7459) );
  OAI22_X1 U9034 ( .A1(n9379), .A2(n7452), .B1(n7774), .B2(n9425), .ZN(n7457)
         );
  OR2_X1 U9035 ( .A1(n7453), .A2(n9775), .ZN(n7454) );
  NAND2_X1 U9036 ( .A1(n7455), .A2(n7454), .ZN(n9777) );
  NOR2_X1 U9037 ( .A1(n9777), .A2(n9247), .ZN(n7456) );
  AOI211_X1 U9038 ( .C1(n9321), .C2(n7784), .A(n7457), .B(n7456), .ZN(n7458)
         );
  OAI211_X1 U9039 ( .C1(n9773), .C2(n7822), .A(n7459), .B(n7458), .ZN(P1_U3282) );
  INV_X1 U9040 ( .A(n7460), .ZN(n7463) );
  INV_X1 U9041 ( .A(n7461), .ZN(n7462) );
  XNOR2_X1 U9042 ( .A(n7630), .B(n8152), .ZN(n7492) );
  NOR2_X1 U9043 ( .A1(n7706), .A2(n8162), .ZN(n7493) );
  XNOR2_X1 U9044 ( .A(n7492), .B(n7493), .ZN(n7490) );
  XOR2_X1 U9045 ( .A(n7491), .B(n7490), .Z(n7472) );
  INV_X1 U9046 ( .A(n7630), .ZN(n9885) );
  OAI22_X1 U9047 ( .A1(n8247), .A2(n9885), .B1(n7638), .B2(n8304), .ZN(n7471)
         );
  NAND2_X1 U9048 ( .A1(n8293), .A2(n7466), .ZN(n7467) );
  OAI211_X1 U9049 ( .C1(n8302), .C2(n7469), .A(n7468), .B(n7467), .ZN(n7470)
         );
  AOI211_X1 U9050 ( .C1(n7472), .C2(n8298), .A(n7471), .B(n7470), .ZN(n7473)
         );
  INV_X1 U9051 ( .A(n7473), .ZN(P2_U3223) );
  AOI21_X1 U9052 ( .B1(n8857), .B2(n9166), .A(n7474), .ZN(n7477) );
  NAND2_X1 U9053 ( .A1(n8819), .A2(n7475), .ZN(n7476) );
  OAI211_X1 U9054 ( .C1(n8853), .C2(n7478), .A(n7477), .B(n7476), .ZN(n7484)
         );
  NAND2_X1 U9055 ( .A1(n7480), .A2(n7479), .ZN(n7481) );
  AOI21_X1 U9056 ( .B1(n7482), .B2(n7481), .A(n8874), .ZN(n7483) );
  AOI211_X1 U9057 ( .C1(n8872), .C2(n7485), .A(n7484), .B(n7483), .ZN(n7486)
         );
  INV_X1 U9058 ( .A(n7486), .ZN(P1_U3211) );
  INV_X1 U9059 ( .A(n9955), .ZN(n7487) );
  OAI222_X1 U9060 ( .A1(P1_U3084), .A2(n7489), .B1(n8222), .B2(n7488), .C1(
        n9550), .C2(n7487), .ZN(P1_U3333) );
  NAND2_X1 U9061 ( .A1(n7491), .A2(n7490), .ZN(n7496) );
  INV_X1 U9062 ( .A(n7492), .ZN(n7494) );
  NAND2_X1 U9063 ( .A1(n7494), .A2(n7493), .ZN(n7495) );
  NAND2_X1 U9064 ( .A1(n7496), .A2(n7495), .ZN(n7505) );
  XNOR2_X1 U9065 ( .A(n7840), .B(n8152), .ZN(n7497) );
  OR2_X1 U9066 ( .A1(n7638), .A2(n8162), .ZN(n7498) );
  NAND2_X1 U9067 ( .A1(n7497), .A2(n7498), .ZN(n7537) );
  INV_X1 U9068 ( .A(n7497), .ZN(n7500) );
  INV_X1 U9069 ( .A(n7498), .ZN(n7499) );
  NAND2_X1 U9070 ( .A1(n7500), .A2(n7499), .ZN(n7501) );
  NAND2_X1 U9071 ( .A1(n7537), .A2(n7501), .ZN(n7504) );
  INV_X1 U9072 ( .A(n7538), .ZN(n7503) );
  AOI21_X1 U9073 ( .B1(n7505), .B2(n7504), .A(n7503), .ZN(n7511) );
  OAI22_X1 U9074 ( .A1(n7706), .A2(n8302), .B1(n8304), .B2(n7705), .ZN(n7509)
         );
  INV_X1 U9075 ( .A(n7716), .ZN(n7507) );
  OAI21_X1 U9076 ( .B1(n8301), .B2(n7507), .A(n7506), .ZN(n7508) );
  AOI211_X1 U9077 ( .C1(n7840), .C2(n8308), .A(n7509), .B(n7508), .ZN(n7510)
         );
  OAI21_X1 U9078 ( .B1(n7511), .B2(n8296), .A(n7510), .ZN(P2_U3233) );
  AOI211_X1 U9079 ( .C1(n9564), .C2(n7664), .A(n7513), .B(n7512), .ZN(n7514)
         );
  OAI21_X1 U9080 ( .B1(n7515), .B2(n9526), .A(n7514), .ZN(n7518) );
  NAND2_X1 U9081 ( .A1(n7518), .A2(n9528), .ZN(n7516) );
  OAI21_X1 U9082 ( .B1(n9528), .B2(n7517), .A(n7516), .ZN(P1_U3533) );
  INV_X1 U9083 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7520) );
  NAND2_X1 U9084 ( .A1(n7518), .A2(n9772), .ZN(n7519) );
  OAI21_X1 U9085 ( .B1(n9772), .B2(n7520), .A(n7519), .ZN(P1_U3484) );
  AOI21_X1 U9086 ( .B1(n7523), .B2(n7522), .A(n7521), .ZN(n7525) );
  INV_X1 U9087 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7910) );
  AOI22_X1 U9088 ( .A1(n7918), .A2(n7910), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n7911), .ZN(n7524) );
  NOR2_X1 U9089 ( .A1(n7525), .A2(n7524), .ZN(n7909) );
  AOI21_X1 U9090 ( .B1(n7525), .B2(n7524), .A(n7909), .ZN(n7536) );
  NOR2_X1 U9091 ( .A1(n7918), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7526) );
  AOI21_X1 U9092 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n7918), .A(n7526), .ZN(
        n7530) );
  OAI21_X1 U9093 ( .B1(n7530), .B2(n7529), .A(n7917), .ZN(n7534) );
  INV_X1 U9094 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7532) );
  NAND2_X1 U9095 ( .A1(n8384), .A2(n7918), .ZN(n7531) );
  NAND2_X1 U9096 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7878) );
  OAI211_X1 U9097 ( .C1(n7532), .C2(n8388), .A(n7531), .B(n7878), .ZN(n7533)
         );
  AOI21_X1 U9098 ( .B1(n7534), .B2(n9791), .A(n7533), .ZN(n7535) );
  OAI21_X1 U9099 ( .B1(n7536), .B2(n9795), .A(n7535), .ZN(P2_U3259) );
  XNOR2_X1 U9100 ( .A(n7675), .B(n8163), .ZN(n7617) );
  NOR2_X1 U9101 ( .A1(n7705), .A2(n8162), .ZN(n7618) );
  XNOR2_X1 U9102 ( .A(n7617), .B(n7618), .ZN(n7621) );
  XNOR2_X1 U9103 ( .A(n7622), .B(n7621), .ZN(n7544) );
  NAND2_X1 U9104 ( .A1(n8293), .A2(n7643), .ZN(n7540) );
  NAND2_X1 U9105 ( .A1(n7540), .A2(n7539), .ZN(n7542) );
  OAI22_X1 U9106 ( .A1(n7638), .A2(n8302), .B1(n8304), .B2(n7739), .ZN(n7541)
         );
  AOI211_X1 U9107 ( .C1(n7675), .C2(n8308), .A(n7542), .B(n7541), .ZN(n7543)
         );
  OAI21_X1 U9108 ( .B1(n7544), .B2(n8296), .A(n7543), .ZN(P2_U3219) );
  INV_X1 U9109 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9649) );
  INV_X1 U9110 ( .A(n7545), .ZN(n7546) );
  AOI22_X1 U9111 ( .A1(n7546), .A2(n9502), .B1(n9564), .B2(n7702), .ZN(n7547)
         );
  OAI211_X1 U9112 ( .C1(n9571), .C2(n7549), .A(n7548), .B(n7547), .ZN(n7551)
         );
  NAND2_X1 U9113 ( .A1(n7551), .A2(n9786), .ZN(n7550) );
  OAI21_X1 U9114 ( .B1(n9528), .B2(n9649), .A(n7550), .ZN(P1_U3531) );
  NAND2_X1 U9115 ( .A1(n7551), .A2(n9783), .ZN(n7552) );
  OAI21_X1 U9116 ( .B1(n9772), .B2(n5209), .A(n7552), .ZN(P1_U3478) );
  INV_X1 U9117 ( .A(n7553), .ZN(n7583) );
  OAI222_X1 U9118 ( .A1(n9550), .A2(n7583), .B1(P1_U3084), .B2(n9106), .C1(
        n7554), .C2(n8222), .ZN(P1_U3332) );
  INV_X1 U9119 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10258) );
  NOR2_X1 U9120 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7555) );
  AOI21_X1 U9121 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7555), .ZN(n9930) );
  NOR2_X1 U9122 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7556) );
  AOI21_X1 U9123 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7556), .ZN(n9933) );
  NOR2_X1 U9124 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7557) );
  AOI21_X1 U9125 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7557), .ZN(n9936) );
  NOR2_X1 U9126 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7558) );
  AOI21_X1 U9127 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7558), .ZN(n9939) );
  NOR2_X1 U9128 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7559) );
  AOI21_X1 U9129 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7559), .ZN(n9942) );
  INV_X1 U9130 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10262) );
  INV_X1 U9131 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10270) );
  INV_X1 U9132 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10269) );
  NOR2_X1 U9133 ( .A1(n10270), .A2(n10269), .ZN(n10268) );
  NOR2_X1 U9134 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(P1_ADDR_REG_4__SCAN_IN), 
        .ZN(n7566) );
  INV_X1 U9135 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9612) );
  AOI22_X1 U9136 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n9612), .B1(
        P1_ADDR_REG_4__SCAN_IN), .B2(n10190), .ZN(n10276) );
  NAND2_X1 U9137 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7564) );
  XOR2_X1 U9138 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10274) );
  NAND2_X1 U9139 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7562) );
  XNOR2_X1 U9140 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n7560), .ZN(n10267) );
  AOI21_X1 U9141 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9923) );
  INV_X1 U9142 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9927) );
  NAND3_X1 U9143 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9925) );
  OAI21_X1 U9144 ( .B1(n9923), .B2(n9927), .A(n9925), .ZN(n10266) );
  NAND2_X1 U9145 ( .A1(n10267), .A2(n10266), .ZN(n7561) );
  NAND2_X1 U9146 ( .A1(n7562), .A2(n7561), .ZN(n10273) );
  NAND2_X1 U9147 ( .A1(n10274), .A2(n10273), .ZN(n7563) );
  NAND2_X1 U9148 ( .A1(n7564), .A2(n7563), .ZN(n10275) );
  NOR2_X1 U9149 ( .A1(n10276), .A2(n10275), .ZN(n7565) );
  NOR2_X1 U9150 ( .A1(n7566), .A2(n7565), .ZN(n7567) );
  NOR2_X1 U9151 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7567), .ZN(n10254) );
  AND2_X1 U9152 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7567), .ZN(n10253) );
  NOR2_X1 U9153 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10253), .ZN(n7568) );
  NOR2_X1 U9154 ( .A1(n10254), .A2(n7568), .ZN(n7569) );
  NAND2_X1 U9155 ( .A1(n7569), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7571) );
  XOR2_X1 U9156 ( .A(n7569), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10252) );
  NAND2_X1 U9157 ( .A1(n10252), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7570) );
  NAND2_X1 U9158 ( .A1(n7571), .A2(n7570), .ZN(n7572) );
  NAND2_X1 U9159 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7572), .ZN(n7574) );
  XOR2_X1 U9160 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7572), .Z(n10251) );
  NAND2_X1 U9161 ( .A1(n10251), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7573) );
  NAND2_X1 U9162 ( .A1(n7574), .A2(n7573), .ZN(n10271) );
  OAI22_X1 U9163 ( .A1(n10268), .A2(n10271), .B1(P2_ADDR_REG_8__SCAN_IN), .B2(
        P1_ADDR_REG_8__SCAN_IN), .ZN(n10263) );
  NOR2_X1 U9164 ( .A1(n10262), .A2(n10263), .ZN(n7575) );
  NAND2_X1 U9165 ( .A1(n10262), .A2(n10263), .ZN(n10261) );
  OAI21_X1 U9166 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n7575), .A(n10261), .ZN(
        n9951) );
  NAND2_X1 U9167 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7576) );
  OAI21_X1 U9168 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7576), .ZN(n9950) );
  NOR2_X1 U9169 ( .A1(n9951), .A2(n9950), .ZN(n9949) );
  AOI21_X1 U9170 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9949), .ZN(n9948) );
  NAND2_X1 U9171 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7577) );
  OAI21_X1 U9172 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7577), .ZN(n9947) );
  NOR2_X1 U9173 ( .A1(n9948), .A2(n9947), .ZN(n9946) );
  AOI21_X1 U9174 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9946), .ZN(n9945) );
  INV_X1 U9175 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10038) );
  NOR2_X1 U9176 ( .A1(n10038), .A2(n10152), .ZN(n10192) );
  AOI21_X1 U9177 ( .B1(n10038), .B2(n10152), .A(n10192), .ZN(n9944) );
  NAND2_X1 U9178 ( .A1(n9945), .A2(n9944), .ZN(n9943) );
  OAI21_X1 U9179 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9943), .ZN(n9941) );
  NAND2_X1 U9180 ( .A1(n9942), .A2(n9941), .ZN(n9940) );
  OAI21_X1 U9181 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9940), .ZN(n9938) );
  NAND2_X1 U9182 ( .A1(n9939), .A2(n9938), .ZN(n9937) );
  OAI21_X1 U9183 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9937), .ZN(n9935) );
  NAND2_X1 U9184 ( .A1(n9936), .A2(n9935), .ZN(n9934) );
  OAI21_X1 U9185 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9934), .ZN(n9932) );
  NAND2_X1 U9186 ( .A1(n9933), .A2(n9932), .ZN(n9931) );
  OAI21_X1 U9187 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9931), .ZN(n9929) );
  NAND2_X1 U9188 ( .A1(n9930), .A2(n9929), .ZN(n9928) );
  OAI21_X1 U9189 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9928), .ZN(n10257) );
  NOR2_X1 U9190 ( .A1(n10258), .A2(n10257), .ZN(n7578) );
  NAND2_X1 U9191 ( .A1(n10258), .A2(n10257), .ZN(n10256) );
  OAI21_X1 U9192 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7578), .A(n10256), .ZN(
        n7580) );
  XNOR2_X1 U9193 ( .A(n9214), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7579) );
  XNOR2_X1 U9194 ( .A(n7580), .B(n7579), .ZN(ADD_1071_U4) );
  INV_X1 U9195 ( .A(n7581), .ZN(n7582) );
  OAI222_X1 U9196 ( .A1(n7728), .A2(n10066), .B1(n8747), .B2(n7583), .C1(n7582), .C2(P2_U3152), .ZN(P2_U3337) );
  OR2_X1 U9197 ( .A1(n7664), .A2(n9164), .ZN(n7584) );
  OR2_X1 U9198 ( .A1(n7794), .A2(n7658), .ZN(n8921) );
  NAND2_X1 U9199 ( .A1(n7794), .A2(n7658), .ZN(n8905) );
  NAND2_X1 U9200 ( .A1(n7587), .A2(n9091), .ZN(n7588) );
  NAND2_X1 U9201 ( .A1(n7605), .A2(n7588), .ZN(n9578) );
  NAND2_X1 U9202 ( .A1(n7592), .A2(n7589), .ZN(n8987) );
  NAND2_X1 U9203 ( .A1(n7592), .A2(n7591), .ZN(n7593) );
  XNOR2_X1 U9204 ( .A(n7613), .B(n9091), .ZN(n7596) );
  INV_X1 U9205 ( .A(n9162), .ZN(n7811) );
  OAI22_X1 U9206 ( .A1(n7594), .A2(n9369), .B1(n7811), .B2(n9371), .ZN(n7595)
         );
  AOI21_X1 U9207 ( .B1(n7596), .B2(n9433), .A(n7595), .ZN(n7597) );
  OAI21_X1 U9208 ( .B1(n9578), .B2(n7815), .A(n7597), .ZN(n9581) );
  NAND2_X1 U9209 ( .A1(n9581), .A2(n9379), .ZN(n7604) );
  OAI22_X1 U9210 ( .A1(n9379), .A2(n7598), .B1(n7792), .B2(n9425), .ZN(n7602)
         );
  AND2_X1 U9211 ( .A1(n7599), .A2(n7794), .ZN(n7600) );
  OR2_X1 U9212 ( .A1(n7600), .A2(n7606), .ZN(n9580) );
  NOR2_X1 U9213 ( .A1(n9580), .A2(n9247), .ZN(n7601) );
  AOI211_X1 U9214 ( .C1(n9321), .C2(n7794), .A(n7602), .B(n7601), .ZN(n7603)
         );
  OAI211_X1 U9215 ( .C1(n9578), .C2(n7822), .A(n7604), .B(n7603), .ZN(P1_U3280) );
  INV_X1 U9216 ( .A(n7794), .ZN(n9579) );
  NAND2_X1 U9217 ( .A1(n7605), .A2(n4921), .ZN(n7798) );
  OR2_X1 U9218 ( .A1(n7894), .A2(n7811), .ZN(n8996) );
  NAND2_X1 U9219 ( .A1(n7894), .A2(n7811), .ZN(n8989) );
  NAND2_X1 U9220 ( .A1(n8996), .A2(n8989), .ZN(n8980) );
  XNOR2_X1 U9221 ( .A(n7798), .B(n8980), .ZN(n7670) );
  INV_X1 U9222 ( .A(n7606), .ZN(n7607) );
  INV_X1 U9223 ( .A(n7894), .ZN(n7608) );
  AOI211_X1 U9224 ( .C1(n7894), .C2(n7607), .A(n9776), .B(n7816), .ZN(n7668)
         );
  NOR2_X1 U9225 ( .A1(n7608), .A2(n9423), .ZN(n7611) );
  OAI22_X1 U9226 ( .A1(n9379), .A2(n7609), .B1(n7892), .B2(n9425), .ZN(n7610)
         );
  AOI211_X1 U9227 ( .C1(n7668), .C2(n9430), .A(n7611), .B(n7610), .ZN(n7616)
         );
  INV_X1 U9228 ( .A(n8905), .ZN(n7612) );
  INV_X1 U9229 ( .A(n8980), .ZN(n9090) );
  XNOR2_X1 U9230 ( .A(n7804), .B(n9090), .ZN(n7614) );
  OAI222_X1 U9231 ( .A1(n9369), .A2(n7658), .B1(n9371), .B2(n7889), .C1(n9389), 
        .C2(n7614), .ZN(n7667) );
  NAND2_X1 U9232 ( .A1(n7667), .A2(n9379), .ZN(n7615) );
  OAI211_X1 U9233 ( .C1(n7670), .C2(n9444), .A(n7616), .B(n7615), .ZN(P1_U3279) );
  INV_X1 U9234 ( .A(n7617), .ZN(n7620) );
  INV_X1 U9235 ( .A(n7618), .ZN(n7619) );
  XNOR2_X1 U9236 ( .A(n7823), .B(n8152), .ZN(n7732) );
  NOR2_X1 U9237 ( .A1(n7739), .A2(n8162), .ZN(n7733) );
  XNOR2_X1 U9238 ( .A(n7732), .B(n7733), .ZN(n7730) );
  XNOR2_X1 U9239 ( .A(n7731), .B(n7730), .ZN(n7629) );
  NAND2_X1 U9240 ( .A1(n8293), .A2(n7623), .ZN(n7624) );
  OAI21_X1 U9241 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n7625), .A(n7624), .ZN(n7627) );
  OAI22_X1 U9242 ( .A1(n7705), .A2(n8302), .B1(n8304), .B2(n7764), .ZN(n7626)
         );
  AOI211_X1 U9243 ( .C1(n7823), .C2(n8308), .A(n7627), .B(n7626), .ZN(n7628)
         );
  OAI21_X1 U9244 ( .B1(n7629), .B2(n8296), .A(n7628), .ZN(P2_U3238) );
  NAND2_X1 U9245 ( .A1(n7630), .A2(n8322), .ZN(n7631) );
  INV_X1 U9246 ( .A(n7709), .ZN(n7634) );
  INV_X1 U9247 ( .A(n7638), .ZN(n8321) );
  OR2_X1 U9248 ( .A1(n7840), .A2(n8321), .ZN(n7635) );
  OAI21_X1 U9249 ( .B1(n4454), .B2(n7636), .A(n7677), .ZN(n9891) );
  XNOR2_X1 U9250 ( .A(n7637), .B(n7636), .ZN(n7640) );
  OAI22_X1 U9251 ( .A1(n7638), .A2(n8615), .B1(n7739), .B2(n8617), .ZN(n7639)
         );
  AOI21_X1 U9252 ( .B1(n7640), .B2(n8585), .A(n7639), .ZN(n7641) );
  OAI21_X1 U9253 ( .B1(n9891), .B2(n9805), .A(n7641), .ZN(n9894) );
  NAND2_X1 U9254 ( .A1(n9894), .A2(n9817), .ZN(n7648) );
  NOR2_X2 U9255 ( .A1(n7715), .A2(n7840), .ZN(n7714) );
  INV_X1 U9256 ( .A(n7675), .ZN(n9892) );
  NAND2_X1 U9257 ( .A1(n7714), .A2(n9892), .ZN(n7748) );
  OR2_X1 U9258 ( .A1(n7714), .A2(n9892), .ZN(n7642) );
  NAND2_X1 U9259 ( .A1(n7748), .A2(n7642), .ZN(n9893) );
  INV_X1 U9260 ( .A(n9893), .ZN(n7646) );
  AOI22_X1 U9261 ( .A1(n8600), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n7643), .B2(
        n9810), .ZN(n7644) );
  OAI21_X1 U9262 ( .B1(n9892), .B2(n8626), .A(n7644), .ZN(n7645) );
  AOI21_X1 U9263 ( .B1(n7646), .B2(n8632), .A(n7645), .ZN(n7647) );
  OAI211_X1 U9264 ( .C1(n9891), .C2(n8629), .A(n7648), .B(n7647), .ZN(P2_U3286) );
  INV_X1 U9265 ( .A(n7649), .ZN(n7652) );
  OAI222_X1 U9266 ( .A1(n7728), .A2(n7651), .B1(n8747), .B2(n7652), .C1(
        P2_U3152), .C2(n7650), .ZN(P2_U3336) );
  OAI222_X1 U9267 ( .A1(n9071), .A2(P1_U3084), .B1(n9550), .B2(n7652), .C1(
        n10230), .C2(n8222), .ZN(P1_U3331) );
  XNOR2_X1 U9268 ( .A(n7655), .B(n7654), .ZN(n7656) );
  XNOR2_X1 U9269 ( .A(n7653), .B(n7656), .ZN(n7666) );
  INV_X1 U9270 ( .A(n7657), .ZN(n7660) );
  NOR2_X1 U9271 ( .A1(n8865), .A2(n7658), .ZN(n7659) );
  AOI211_X1 U9272 ( .C1(n8868), .C2(n9165), .A(n7660), .B(n7659), .ZN(n7661)
         );
  OAI21_X1 U9273 ( .B1(n8870), .B2(n7662), .A(n7661), .ZN(n7663) );
  AOI21_X1 U9274 ( .B1(n8872), .B2(n7664), .A(n7663), .ZN(n7665) );
  OAI21_X1 U9275 ( .B1(n7666), .B2(n8874), .A(n7665), .ZN(P1_U3215) );
  INV_X1 U9276 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7672) );
  AOI211_X1 U9277 ( .C1(n9564), .C2(n7894), .A(n7668), .B(n7667), .ZN(n7669)
         );
  OAI21_X1 U9278 ( .B1(n7670), .B2(n9526), .A(n7669), .ZN(n7673) );
  NAND2_X1 U9279 ( .A1(n7673), .A2(n9772), .ZN(n7671) );
  OAI21_X1 U9280 ( .B1(n9772), .B2(n7672), .A(n7671), .ZN(P1_U3490) );
  INV_X1 U9281 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9174) );
  NAND2_X1 U9282 ( .A1(n7673), .A2(n9786), .ZN(n7674) );
  OAI21_X1 U9283 ( .B1(n9528), .B2(n9174), .A(n7674), .ZN(P1_U3535) );
  INV_X1 U9284 ( .A(n7705), .ZN(n8320) );
  NAND2_X1 U9285 ( .A1(n7675), .A2(n8320), .ZN(n7676) );
  INV_X1 U9286 ( .A(n7739), .ZN(n8319) );
  NAND2_X1 U9287 ( .A1(n7823), .A2(n8319), .ZN(n7678) );
  NAND2_X1 U9288 ( .A1(n7679), .A2(n7678), .ZN(n7929) );
  XNOR2_X1 U9289 ( .A(n7929), .B(n7930), .ZN(n9905) );
  INV_X1 U9290 ( .A(n9905), .ZN(n7690) );
  NAND2_X1 U9291 ( .A1(n7680), .A2(n7681), .ZN(n7683) );
  XNOR2_X1 U9292 ( .A(n7683), .B(n7682), .ZN(n7684) );
  OAI222_X1 U9293 ( .A1(n8617), .A2(n7965), .B1(n8615), .B2(n7739), .C1(n7684), 
        .C2(n8612), .ZN(n9902) );
  INV_X1 U9294 ( .A(n7931), .ZN(n9899) );
  OR2_X2 U9295 ( .A1(n7748), .A2(n7823), .ZN(n7685) );
  INV_X1 U9296 ( .A(n7685), .ZN(n7747) );
  OAI21_X1 U9297 ( .B1(n9899), .B2(n7747), .A(n4442), .ZN(n9901) );
  AOI22_X1 U9298 ( .A1(n8600), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7736), .B2(
        n9810), .ZN(n7687) );
  NAND2_X1 U9299 ( .A1(n7931), .A2(n8473), .ZN(n7686) );
  OAI211_X1 U9300 ( .C1(n9901), .C2(n8475), .A(n7687), .B(n7686), .ZN(n7688)
         );
  AOI21_X1 U9301 ( .B1(n9902), .B2(n9817), .A(n7688), .ZN(n7689) );
  OAI21_X1 U9302 ( .B1(n8606), .B2(n7690), .A(n7689), .ZN(P2_U3284) );
  NOR2_X1 U9303 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10219), .ZN(n9646) );
  AOI21_X1 U9304 ( .B1(n8857), .B2(n9165), .A(n9646), .ZN(n7693) );
  NAND2_X1 U9305 ( .A1(n8819), .A2(n7691), .ZN(n7692) );
  OAI211_X1 U9306 ( .C1(n8853), .C2(n7694), .A(n7693), .B(n7692), .ZN(n7701)
         );
  NAND2_X1 U9307 ( .A1(n7695), .A2(n7696), .ZN(n7698) );
  XNOR2_X1 U9308 ( .A(n7698), .B(n7697), .ZN(n7699) );
  NOR2_X1 U9309 ( .A1(n7699), .A2(n8874), .ZN(n7700) );
  AOI211_X1 U9310 ( .C1(n8872), .C2(n7702), .A(n7701), .B(n7700), .ZN(n7703)
         );
  INV_X1 U9311 ( .A(n7703), .ZN(P1_U3219) );
  XNOR2_X1 U9312 ( .A(n7704), .B(n7710), .ZN(n7713) );
  OAI22_X1 U9313 ( .A1(n7706), .A2(n8615), .B1(n7705), .B2(n8617), .ZN(n7712)
         );
  INV_X1 U9314 ( .A(n7707), .ZN(n7708) );
  AOI21_X1 U9315 ( .B1(n7710), .B2(n7709), .A(n7708), .ZN(n7844) );
  NOR2_X1 U9316 ( .A1(n7844), .A2(n9805), .ZN(n7711) );
  AOI211_X1 U9317 ( .C1(n7713), .C2(n8585), .A(n7712), .B(n7711), .ZN(n7843)
         );
  AOI21_X1 U9318 ( .B1(n7840), .B2(n7715), .A(n7714), .ZN(n7841) );
  INV_X1 U9319 ( .A(n7840), .ZN(n7718) );
  AOI22_X1 U9320 ( .A1(n8600), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7716), .B2(
        n9810), .ZN(n7717) );
  OAI21_X1 U9321 ( .B1(n7718), .B2(n8626), .A(n7717), .ZN(n7720) );
  NOR2_X1 U9322 ( .A1(n7844), .A2(n8629), .ZN(n7719) );
  AOI211_X1 U9323 ( .C1(n7841), .C2(n8632), .A(n7720), .B(n7719), .ZN(n7721)
         );
  OAI21_X1 U9324 ( .B1(n7843), .B2(n8600), .A(n7721), .ZN(P2_U3287) );
  INV_X1 U9325 ( .A(n7725), .ZN(n7724) );
  NAND2_X1 U9326 ( .A1(n9548), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7723) );
  NAND2_X1 U9327 ( .A1(n7722), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9154) );
  OAI211_X1 U9328 ( .C1(n7724), .C2(n9550), .A(n7723), .B(n9154), .ZN(P1_U3330) );
  NAND2_X1 U9329 ( .A1(n7725), .A2(n9954), .ZN(n7727) );
  OAI211_X1 U9330 ( .C1(n7729), .C2(n7728), .A(n7727), .B(n7726), .ZN(P2_U3335) );
  INV_X1 U9331 ( .A(n7732), .ZN(n7734) );
  NAND2_X1 U9332 ( .A1(n7734), .A2(n7733), .ZN(n7758) );
  NAND2_X1 U9333 ( .A1(n7763), .A2(n7758), .ZN(n7735) );
  XNOR2_X1 U9334 ( .A(n7931), .B(n8152), .ZN(n7755) );
  NOR2_X1 U9335 ( .A1(n7764), .A2(n8162), .ZN(n7756) );
  XNOR2_X1 U9336 ( .A(n7755), .B(n7756), .ZN(n7760) );
  XNOR2_X1 U9337 ( .A(n7735), .B(n7760), .ZN(n7743) );
  NAND2_X1 U9338 ( .A1(n8293), .A2(n7736), .ZN(n7738) );
  NAND2_X1 U9339 ( .A1(n7738), .A2(n7737), .ZN(n7741) );
  OAI22_X1 U9340 ( .A1(n7739), .A2(n8302), .B1(n8304), .B2(n7965), .ZN(n7740)
         );
  AOI211_X1 U9341 ( .C1(n7931), .C2(n8308), .A(n7741), .B(n7740), .ZN(n7742)
         );
  OAI21_X1 U9342 ( .B1(n7743), .B2(n8296), .A(n7742), .ZN(P2_U3226) );
  INV_X1 U9343 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7751) );
  XNOR2_X1 U9344 ( .A(n7744), .B(n7745), .ZN(n7833) );
  OAI21_X1 U9345 ( .B1(n4937), .B2(n5983), .A(n7680), .ZN(n7746) );
  INV_X1 U9346 ( .A(n7764), .ZN(n8318) );
  AOI222_X1 U9347 ( .A1(n8585), .A2(n7746), .B1(n8318), .B2(n8590), .C1(n8320), 
        .C2(n8591), .ZN(n7828) );
  AOI21_X1 U9348 ( .B1(n7823), .B2(n7748), .A(n7747), .ZN(n7831) );
  AOI22_X1 U9349 ( .A1(n7831), .A2(n9869), .B1(n9868), .B2(n7823), .ZN(n7749)
         );
  OAI211_X1 U9350 ( .C1(n8720), .C2(n7833), .A(n7828), .B(n7749), .ZN(n7752)
         );
  NAND2_X1 U9351 ( .A1(n7752), .A2(n9908), .ZN(n7750) );
  OAI21_X1 U9352 ( .B1(n9908), .B2(n7751), .A(n7750), .ZN(P2_U3484) );
  NAND2_X1 U9353 ( .A1(n7752), .A2(n9914), .ZN(n7753) );
  OAI21_X1 U9354 ( .B1(n9914), .B2(n7754), .A(n7753), .ZN(P2_U3531) );
  INV_X1 U9355 ( .A(n7755), .ZN(n7757) );
  NAND2_X1 U9356 ( .A1(n7757), .A2(n7756), .ZN(n7759) );
  AND2_X1 U9357 ( .A1(n7758), .A2(n7759), .ZN(n7762) );
  INV_X1 U9358 ( .A(n7759), .ZN(n7761) );
  XNOR2_X1 U9359 ( .A(n8722), .B(n8152), .ZN(n7872) );
  NOR2_X1 U9360 ( .A1(n7965), .A2(n8162), .ZN(n7873) );
  XNOR2_X1 U9361 ( .A(n7872), .B(n7873), .ZN(n7870) );
  XNOR2_X1 U9362 ( .A(n7871), .B(n7870), .ZN(n7772) );
  INV_X1 U9363 ( .A(n7937), .ZN(n7769) );
  INV_X1 U9364 ( .A(n8170), .ZN(n8271) );
  OR2_X1 U9365 ( .A1(n7991), .A2(n8617), .ZN(n7766) );
  OR2_X1 U9366 ( .A1(n7764), .A2(n8615), .ZN(n7765) );
  NAND2_X1 U9367 ( .A1(n7766), .A2(n7765), .ZN(n7935) );
  NAND2_X1 U9368 ( .A1(n8271), .A2(n7935), .ZN(n7767) );
  OAI211_X1 U9369 ( .C1(n8301), .C2(n7769), .A(n7768), .B(n7767), .ZN(n7770)
         );
  AOI21_X1 U9370 ( .B1(n8722), .B2(n8308), .A(n7770), .ZN(n7771) );
  OAI21_X1 U9371 ( .B1(n7772), .B2(n8296), .A(n7771), .ZN(P2_U3236) );
  AOI21_X1 U9372 ( .B1(n8857), .B2(n9164), .A(n7773), .ZN(n7777) );
  INV_X1 U9373 ( .A(n7774), .ZN(n7775) );
  NAND2_X1 U9374 ( .A1(n8819), .A2(n7775), .ZN(n7776) );
  OAI211_X1 U9375 ( .C1(n8853), .C2(n7778), .A(n7777), .B(n7776), .ZN(n7783)
         );
  XOR2_X1 U9376 ( .A(n7779), .B(n7780), .Z(n7781) );
  NOR2_X1 U9377 ( .A1(n7781), .A2(n8874), .ZN(n7782) );
  AOI211_X1 U9378 ( .C1(n8872), .C2(n7784), .A(n7783), .B(n7782), .ZN(n7785)
         );
  INV_X1 U9379 ( .A(n7785), .ZN(P1_U3229) );
  XNOR2_X1 U9380 ( .A(n7786), .B(n7787), .ZN(n7796) );
  INV_X1 U9381 ( .A(n7788), .ZN(n7790) );
  NOR2_X1 U9382 ( .A1(n8865), .A2(n7811), .ZN(n7789) );
  AOI211_X1 U9383 ( .C1(n8868), .C2(n9164), .A(n7790), .B(n7789), .ZN(n7791)
         );
  OAI21_X1 U9384 ( .B1(n8870), .B2(n7792), .A(n7791), .ZN(n7793) );
  AOI21_X1 U9385 ( .B1(n8872), .B2(n7794), .A(n7793), .ZN(n7795) );
  OAI21_X1 U9386 ( .B1(n7796), .B2(n8874), .A(n7795), .ZN(P1_U3234) );
  AOI21_X1 U9387 ( .B1(n7798), .B2(n8980), .A(n7797), .ZN(n7808) );
  NAND2_X1 U9388 ( .A1(n7808), .A2(n4931), .ZN(n7800) );
  XNOR2_X1 U9389 ( .A(n9524), .B(n8904), .ZN(n9094) );
  XOR2_X1 U9390 ( .A(n7850), .B(n9094), .Z(n9527) );
  INV_X1 U9391 ( .A(n7856), .ZN(n7857) );
  AOI211_X1 U9392 ( .C1(n9524), .C2(n4396), .A(n9776), .B(n7856), .ZN(n9523)
         );
  INV_X1 U9393 ( .A(n9524), .ZN(n7849) );
  NOR2_X1 U9394 ( .A1(n7849), .A2(n9423), .ZN(n7803) );
  OAI22_X1 U9395 ( .A1(n9379), .A2(n7801), .B1(n8033), .B2(n9425), .ZN(n7802)
         );
  AOI211_X1 U9396 ( .C1(n9523), .C2(n9430), .A(n7803), .B(n7802), .ZN(n7807)
         );
  OR2_X1 U9397 ( .A1(n7906), .A2(n7889), .ZN(n9003) );
  NAND2_X1 U9398 ( .A1(n7906), .A2(n7889), .ZN(n8999) );
  XNOR2_X1 U9399 ( .A(n7851), .B(n9094), .ZN(n7805) );
  OAI222_X1 U9400 ( .A1(n9371), .A2(n8030), .B1(n9369), .B2(n7889), .C1(n9389), 
        .C2(n7805), .ZN(n9522) );
  NAND2_X1 U9401 ( .A1(n9522), .A2(n9379), .ZN(n7806) );
  OAI211_X1 U9402 ( .C1(n9527), .C2(n9444), .A(n7807), .B(n7806), .ZN(P1_U3277) );
  XNOR2_X1 U9403 ( .A(n7808), .B(n9092), .ZN(n9572) );
  OAI21_X1 U9404 ( .B1(n9092), .B2(n7810), .A(n7809), .ZN(n7813) );
  OAI22_X1 U9405 ( .A1(n7811), .A2(n9369), .B1(n8904), .B2(n9371), .ZN(n7812)
         );
  AOI21_X1 U9406 ( .B1(n7813), .B2(n9433), .A(n7812), .ZN(n7814) );
  OAI21_X1 U9407 ( .B1(n9572), .B2(n7815), .A(n7814), .ZN(n9575) );
  NAND2_X1 U9408 ( .A1(n9575), .A2(n9379), .ZN(n7821) );
  OAI22_X1 U9409 ( .A1(n9379), .A2(n9190), .B1(n7904), .B2(n9425), .ZN(n7819)
         );
  OR2_X1 U9410 ( .A1(n7816), .A2(n9573), .ZN(n7817) );
  NAND2_X1 U9411 ( .A1(n4396), .A2(n7817), .ZN(n9574) );
  NOR2_X1 U9412 ( .A1(n9574), .A2(n9247), .ZN(n7818) );
  AOI211_X1 U9413 ( .C1(n9321), .C2(n7906), .A(n7819), .B(n7818), .ZN(n7820)
         );
  OAI211_X1 U9414 ( .C1(n9572), .C2(n7822), .A(n7821), .B(n7820), .ZN(P1_U3278) );
  INV_X1 U9415 ( .A(n7823), .ZN(n7827) );
  NOR2_X1 U9416 ( .A1(n8469), .A2(n7824), .ZN(n7825) );
  AOI21_X1 U9417 ( .B1(n8600), .B2(P2_REG2_REG_11__SCAN_IN), .A(n7825), .ZN(
        n7826) );
  OAI21_X1 U9418 ( .B1(n7827), .B2(n8626), .A(n7826), .ZN(n7830) );
  NOR2_X1 U9419 ( .A1(n7828), .A2(n8600), .ZN(n7829) );
  AOI211_X1 U9420 ( .C1(n7831), .C2(n8632), .A(n7830), .B(n7829), .ZN(n7832)
         );
  OAI21_X1 U9421 ( .B1(n8606), .B2(n7833), .A(n7832), .ZN(P2_U3285) );
  INV_X1 U9422 ( .A(n7834), .ZN(n7837) );
  OAI222_X1 U9423 ( .A1(P2_U3152), .A2(n7836), .B1(n8747), .B2(n7837), .C1(
        n7835), .C2(n7728), .ZN(P2_U3334) );
  OAI222_X1 U9424 ( .A1(n7839), .A2(P1_U3084), .B1(n8222), .B2(n7838), .C1(
        n9550), .C2(n7837), .ZN(P1_U3329) );
  INV_X1 U9425 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7846) );
  AOI22_X1 U9426 ( .A1(n7841), .A2(n9869), .B1(n9868), .B2(n7840), .ZN(n7842)
         );
  OAI211_X1 U9427 ( .C1(n7844), .C2(n9883), .A(n7843), .B(n7842), .ZN(n7847)
         );
  NAND2_X1 U9428 ( .A1(n7847), .A2(n9908), .ZN(n7845) );
  OAI21_X1 U9429 ( .B1(n9908), .B2(n7846), .A(n7845), .ZN(P2_U3478) );
  NAND2_X1 U9430 ( .A1(n7847), .A2(n9914), .ZN(n7848) );
  OAI21_X1 U9431 ( .B1(n9914), .B2(n6750), .A(n7848), .ZN(P2_U3529) );
  NAND2_X1 U9432 ( .A1(n8073), .A2(n8030), .ZN(n9014) );
  XNOR2_X1 U9433 ( .A(n7947), .B(n9095), .ZN(n9569) );
  INV_X1 U9434 ( .A(n9569), .ZN(n7864) );
  OR2_X1 U9435 ( .A1(n9524), .A2(n8904), .ZN(n9004) );
  XNOR2_X1 U9436 ( .A(n7951), .B(n9095), .ZN(n7852) );
  NAND2_X1 U9437 ( .A1(n7852), .A2(n9433), .ZN(n7854) );
  AOI22_X1 U9438 ( .A1(n9437), .A2(n9160), .B1(n9158), .B2(n9438), .ZN(n7853)
         );
  NAND2_X1 U9439 ( .A1(n7854), .A2(n7853), .ZN(n9568) );
  NAND2_X1 U9440 ( .A1(n7857), .A2(n8073), .ZN(n7858) );
  NAND2_X1 U9441 ( .A1(n7948), .A2(n7858), .ZN(n9566) );
  INV_X1 U9442 ( .A(n8069), .ZN(n7859) );
  OAI22_X1 U9443 ( .A1(n9379), .A2(n9700), .B1(n7859), .B2(n9425), .ZN(n7860)
         );
  AOI21_X1 U9444 ( .B1(n8073), .B2(n9321), .A(n7860), .ZN(n7861) );
  OAI21_X1 U9445 ( .B1(n9566), .B2(n9247), .A(n7861), .ZN(n7862) );
  AOI21_X1 U9446 ( .B1(n9568), .B2(n9379), .A(n7862), .ZN(n7863) );
  OAI21_X1 U9447 ( .B1(n7864), .B2(n9444), .A(n7863), .ZN(P1_U3276) );
  XNOR2_X1 U9448 ( .A(n8716), .B(n8152), .ZN(n7865) );
  OR2_X1 U9449 ( .A1(n7991), .A2(n8162), .ZN(n7866) );
  NAND2_X1 U9450 ( .A1(n7865), .A2(n7866), .ZN(n8010) );
  INV_X1 U9451 ( .A(n7865), .ZN(n7868) );
  INV_X1 U9452 ( .A(n7866), .ZN(n7867) );
  NAND2_X1 U9453 ( .A1(n7868), .A2(n7867), .ZN(n7869) );
  NAND2_X1 U9454 ( .A1(n8010), .A2(n7869), .ZN(n7877) );
  INV_X1 U9455 ( .A(n7872), .ZN(n7874) );
  INV_X1 U9456 ( .A(n8011), .ZN(n7875) );
  AOI21_X1 U9457 ( .B1(n7877), .B2(n7876), .A(n7875), .ZN(n7883) );
  INV_X1 U9458 ( .A(n7959), .ZN(n7880) );
  INV_X1 U9459 ( .A(n8616), .ZN(n8315) );
  INV_X1 U9460 ( .A(n7965), .ZN(n8317) );
  AOI22_X1 U9461 ( .A1(n8281), .A2(n8315), .B1(n8280), .B2(n8317), .ZN(n7879)
         );
  OAI211_X1 U9462 ( .C1(n7880), .C2(n8301), .A(n7879), .B(n7878), .ZN(n7881)
         );
  AOI21_X1 U9463 ( .B1(n8716), .B2(n8308), .A(n7881), .ZN(n7882) );
  OAI21_X1 U9464 ( .B1(n7883), .B2(n8296), .A(n7882), .ZN(P2_U3217) );
  INV_X1 U9465 ( .A(n7885), .ZN(n7886) );
  AOI21_X1 U9466 ( .B1(n7887), .B2(n7884), .A(n7886), .ZN(n7896) );
  NOR2_X1 U9467 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7888), .ZN(n9660) );
  NOR2_X1 U9468 ( .A1(n8865), .A2(n7889), .ZN(n7890) );
  AOI211_X1 U9469 ( .C1(n8868), .C2(n9163), .A(n9660), .B(n7890), .ZN(n7891)
         );
  OAI21_X1 U9470 ( .B1(n8870), .B2(n7892), .A(n7891), .ZN(n7893) );
  AOI21_X1 U9471 ( .B1(n7894), .B2(n8872), .A(n7893), .ZN(n7895) );
  OAI21_X1 U9472 ( .B1(n7896), .B2(n8874), .A(n7895), .ZN(P1_U3222) );
  INV_X1 U9473 ( .A(n7898), .ZN(n7900) );
  NAND2_X1 U9474 ( .A1(n7900), .A2(n7899), .ZN(n7901) );
  XNOR2_X1 U9475 ( .A(n7897), .B(n7901), .ZN(n7908) );
  NOR2_X1 U9476 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5347), .ZN(n9672) );
  NOR2_X1 U9477 ( .A1(n8865), .A2(n8904), .ZN(n7902) );
  AOI211_X1 U9478 ( .C1(n8868), .C2(n9162), .A(n9672), .B(n7902), .ZN(n7903)
         );
  OAI21_X1 U9479 ( .B1(n8870), .B2(n7904), .A(n7903), .ZN(n7905) );
  AOI21_X1 U9480 ( .B1(n7906), .B2(n8872), .A(n7905), .ZN(n7907) );
  OAI21_X1 U9481 ( .B1(n7908), .B2(n8874), .A(n7907), .ZN(P1_U3232) );
  AOI21_X1 U9482 ( .B1(n7911), .B2(n7910), .A(n7909), .ZN(n7912) );
  NAND2_X1 U9483 ( .A1(n8336), .A2(n7912), .ZN(n7913) );
  XNOR2_X1 U9484 ( .A(n7912), .B(n7919), .ZN(n8330) );
  NAND2_X1 U9485 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8330), .ZN(n8329) );
  NAND2_X1 U9486 ( .A1(n7913), .A2(n8329), .ZN(n7915) );
  XNOR2_X1 U9487 ( .A(n8342), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n7914) );
  NOR2_X1 U9488 ( .A1(n7914), .A2(n7915), .ZN(n8348) );
  AOI21_X1 U9489 ( .B1(n7915), .B2(n7914), .A(n8348), .ZN(n7928) );
  AND2_X1 U9490 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8043) );
  AOI21_X1 U9491 ( .B1(n9797), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8043), .ZN(
        n7916) );
  INV_X1 U9492 ( .A(n7916), .ZN(n7926) );
  OAI21_X1 U9493 ( .B1(n7918), .B2(P2_REG2_REG_14__SCAN_IN), .A(n7917), .ZN(
        n7920) );
  NAND2_X1 U9494 ( .A1(n7919), .A2(n7920), .ZN(n7921) );
  XNOR2_X1 U9495 ( .A(n7920), .B(n8336), .ZN(n8333) );
  INV_X1 U9496 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8332) );
  NAND2_X1 U9497 ( .A1(n8333), .A2(n8332), .ZN(n8331) );
  NAND2_X1 U9498 ( .A1(n7921), .A2(n8331), .ZN(n7924) );
  NAND2_X1 U9499 ( .A1(n8342), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7922) );
  OAI21_X1 U9500 ( .B1(n8342), .B2(P2_REG2_REG_16__SCAN_IN), .A(n7922), .ZN(
        n7923) );
  NOR2_X1 U9501 ( .A1(n7923), .A2(n7924), .ZN(n8341) );
  AOI211_X1 U9502 ( .C1(n7924), .C2(n7923), .A(n8341), .B(n9792), .ZN(n7925)
         );
  AOI211_X1 U9503 ( .C1(n8384), .C2(n8342), .A(n7926), .B(n7925), .ZN(n7927)
         );
  OAI21_X1 U9504 ( .B1(n7928), .B2(n9795), .A(n7927), .ZN(P2_U3261) );
  OAI21_X1 U9505 ( .B1(n4447), .B2(n4767), .A(n7963), .ZN(n7936) );
  OAI21_X1 U9506 ( .B1(n7933), .B2(n7932), .A(n7955), .ZN(n8726) );
  NOR2_X1 U9507 ( .A1(n8726), .A2(n9805), .ZN(n7934) );
  AOI211_X1 U9508 ( .C1(n8585), .C2(n7936), .A(n7935), .B(n7934), .ZN(n8725)
         );
  INV_X1 U9509 ( .A(n8722), .ZN(n7939) );
  AOI21_X1 U9510 ( .B1(n8722), .B2(n4442), .A(n7957), .ZN(n8723) );
  AOI22_X1 U9511 ( .A1(n8600), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7937), .B2(
        n9810), .ZN(n7938) );
  OAI21_X1 U9512 ( .B1(n7939), .B2(n8626), .A(n7938), .ZN(n7941) );
  NOR2_X1 U9513 ( .A1(n8726), .A2(n8629), .ZN(n7940) );
  AOI211_X1 U9514 ( .C1(n8723), .C2(n8632), .A(n7941), .B(n7940), .ZN(n7942)
         );
  OAI21_X1 U9515 ( .B1(n8725), .B2(n8600), .A(n7942), .ZN(P2_U3283) );
  INV_X1 U9516 ( .A(n7943), .ZN(n7946) );
  OAI222_X1 U9517 ( .A1(P1_U3084), .A2(n7944), .B1(n9550), .B2(n7946), .C1(
        n10223), .C2(n8222), .ZN(P1_U3328) );
  OAI222_X1 U9518 ( .A1(n7728), .A2(n10086), .B1(n8747), .B2(n7946), .C1(
        P2_U3152), .C2(n7945), .ZN(P2_U3333) );
  INV_X1 U9519 ( .A(n9158), .ZN(n7982) );
  OR2_X1 U9520 ( .A1(n9519), .A2(n7982), .ZN(n9018) );
  NAND2_X1 U9521 ( .A1(n9519), .A2(n7982), .ZN(n9017) );
  NAND2_X1 U9522 ( .A1(n9018), .A2(n9017), .ZN(n9096) );
  XNOR2_X1 U9523 ( .A(n7979), .B(n9096), .ZN(n9521) );
  AOI211_X1 U9524 ( .C1(n9519), .C2(n7948), .A(n9776), .B(n7983), .ZN(n9518)
         );
  NOR2_X1 U9525 ( .A1(n4611), .A2(n9423), .ZN(n7950) );
  OAI22_X1 U9526 ( .A1(n9379), .A2(n9197), .B1(n8806), .B2(n9425), .ZN(n7949)
         );
  AOI211_X1 U9527 ( .C1(n9518), .C2(n9430), .A(n7950), .B(n7949), .ZN(n7954)
         );
  INV_X1 U9528 ( .A(n9436), .ZN(n8803) );
  XNOR2_X1 U9529 ( .A(n7980), .B(n9096), .ZN(n7952) );
  OAI222_X1 U9530 ( .A1(n9369), .A2(n8030), .B1(n9371), .B2(n8803), .C1(n9389), 
        .C2(n7952), .ZN(n9517) );
  NAND2_X1 U9531 ( .A1(n9517), .A2(n9379), .ZN(n7953) );
  OAI211_X1 U9532 ( .C1(n9521), .C2(n9444), .A(n7954), .B(n7953), .ZN(P1_U3275) );
  XNOR2_X1 U9533 ( .A(n7993), .B(n7956), .ZN(n8721) );
  INV_X1 U9534 ( .A(n7957), .ZN(n7958) );
  INV_X1 U9535 ( .A(n8716), .ZN(n7961) );
  AOI21_X1 U9536 ( .B1(n8716), .B2(n7958), .A(n4642), .ZN(n8717) );
  AOI22_X1 U9537 ( .A1(n8600), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7959), .B2(
        n9810), .ZN(n7960) );
  OAI21_X1 U9538 ( .B1(n7961), .B2(n8626), .A(n7960), .ZN(n7970) );
  AOI21_X1 U9539 ( .B1(n7963), .B2(n7962), .A(n7992), .ZN(n7964) );
  NOR2_X1 U9540 ( .A1(n7964), .A2(n8612), .ZN(n7968) );
  OAI22_X1 U9541 ( .A1(n8616), .A2(n8617), .B1(n7965), .B2(n8615), .ZN(n7966)
         );
  AOI21_X1 U9542 ( .B1(n7968), .B2(n7967), .A(n7966), .ZN(n8719) );
  NOR2_X1 U9543 ( .A1(n8719), .A2(n8600), .ZN(n7969) );
  AOI211_X1 U9544 ( .C1(n8717), .C2(n8632), .A(n7970), .B(n7969), .ZN(n7971)
         );
  OAI21_X1 U9545 ( .B1(n8606), .B2(n8721), .A(n7971), .ZN(P2_U3282) );
  INV_X1 U9546 ( .A(n7972), .ZN(n7975) );
  OAI222_X1 U9547 ( .A1(n7974), .A2(P1_U3084), .B1(n9550), .B2(n7975), .C1(
        n7973), .C2(n8222), .ZN(P1_U3327) );
  OAI222_X1 U9548 ( .A1(n7728), .A2(n7977), .B1(P2_U3152), .B2(n7976), .C1(
        n7975), .C2(n8747), .ZN(P2_U3332) );
  AOI21_X1 U9549 ( .B1(n7979), .B2(n9096), .A(n7978), .ZN(n8112) );
  AND2_X1 U9550 ( .A1(n9514), .A2(n8803), .ZN(n8902) );
  INV_X1 U9551 ( .A(n8902), .ZN(n8963) );
  OR2_X1 U9552 ( .A1(n9514), .A2(n8803), .ZN(n8888) );
  XNOR2_X1 U9553 ( .A(n8112), .B(n9098), .ZN(n9516) );
  INV_X1 U9554 ( .A(n9410), .ZN(n8815) );
  XOR2_X1 U9555 ( .A(n8127), .B(n9098), .Z(n7981) );
  OAI222_X1 U9556 ( .A1(n9369), .A2(n7982), .B1(n9371), .B2(n8815), .C1(n7981), 
        .C2(n9389), .ZN(n9512) );
  INV_X1 U9557 ( .A(n7983), .ZN(n7984) );
  AOI211_X1 U9558 ( .C1(n9514), .C2(n7984), .A(n9776), .B(n9420), .ZN(n9513)
         );
  NAND2_X1 U9559 ( .A1(n9513), .A2(n9430), .ZN(n7986) );
  AOI22_X1 U9560 ( .A1(n9404), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n8820), .B2(
        n9402), .ZN(n7985) );
  OAI211_X1 U9561 ( .C1(n8816), .C2(n9423), .A(n7986), .B(n7985), .ZN(n7987)
         );
  AOI21_X1 U9562 ( .B1(n9512), .B2(n9379), .A(n7987), .ZN(n7988) );
  OAI21_X1 U9563 ( .B1(n9516), .B2(n9444), .A(n7988), .ZN(P1_U3274) );
  INV_X1 U9564 ( .A(n7989), .ZN(n8005) );
  AOI21_X1 U9565 ( .B1(n9548), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n9207), .ZN(
        n7990) );
  OAI21_X1 U9566 ( .B1(n8005), .B2(n9550), .A(n7990), .ZN(P1_U3326) );
  INV_X1 U9567 ( .A(n7991), .ZN(n8316) );
  NAND2_X1 U9568 ( .A1(n7994), .A2(n7999), .ZN(n8186) );
  OAI21_X1 U9569 ( .B1(n7994), .B2(n7999), .A(n8186), .ZN(n7995) );
  INV_X1 U9570 ( .A(n7995), .ZN(n8715) );
  AOI21_X1 U9571 ( .B1(n8711), .B2(n7996), .A(n4641), .ZN(n8712) );
  INV_X1 U9572 ( .A(n8711), .ZN(n7998) );
  AOI22_X1 U9573 ( .A1(n8600), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8017), .B2(
        n9810), .ZN(n7997) );
  OAI21_X1 U9574 ( .B1(n7998), .B2(n8626), .A(n7997), .ZN(n8003) );
  XNOR2_X1 U9575 ( .A(n8000), .B(n7999), .ZN(n8001) );
  INV_X1 U9576 ( .A(n8262), .ZN(n8592) );
  AOI222_X1 U9577 ( .A1(n8585), .A2(n8001), .B1(n8316), .B2(n8591), .C1(n8592), 
        .C2(n8590), .ZN(n8714) );
  NOR2_X1 U9578 ( .A1(n8714), .A2(n8600), .ZN(n8002) );
  AOI211_X1 U9579 ( .C1(n8712), .C2(n8632), .A(n8003), .B(n8002), .ZN(n8004)
         );
  OAI21_X1 U9580 ( .B1(n8606), .B2(n8715), .A(n8004), .ZN(P2_U3281) );
  OAI222_X1 U9581 ( .A1(n7728), .A2(n8006), .B1(n8747), .B2(n8005), .C1(
        P2_U3152), .C2(n8212), .ZN(P2_U3331) );
  INV_X1 U9582 ( .A(n8007), .ZN(n8024) );
  AOI21_X1 U9583 ( .B1(n9548), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n8008), .ZN(
        n8009) );
  OAI21_X1 U9584 ( .B1(n8024), .B2(n9550), .A(n8009), .ZN(P1_U3325) );
  NOR2_X1 U9585 ( .A1(n8616), .A2(n8162), .ZN(n8016) );
  NAND2_X1 U9586 ( .A1(n8011), .A2(n8010), .ZN(n8013) );
  XNOR2_X1 U9587 ( .A(n8711), .B(n8152), .ZN(n8012) );
  AOI21_X1 U9588 ( .B1(n8016), .B2(n8015), .A(n4440), .ZN(n8023) );
  INV_X1 U9589 ( .A(n8017), .ZN(n8020) );
  AOI22_X1 U9590 ( .A1(n8281), .A2(n8592), .B1(n8280), .B2(n8316), .ZN(n8019)
         );
  NOR2_X1 U9591 ( .A1(n10068), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8335) );
  INV_X1 U9592 ( .A(n8335), .ZN(n8018) );
  OAI211_X1 U9593 ( .C1(n8020), .C2(n8301), .A(n8019), .B(n8018), .ZN(n8021)
         );
  AOI21_X1 U9594 ( .B1(n8711), .B2(n8308), .A(n8021), .ZN(n8022) );
  OAI21_X1 U9595 ( .B1(n8023), .B2(n8296), .A(n8022), .ZN(P2_U3243) );
  OAI222_X1 U9596 ( .A1(n6416), .A2(P2_U3152), .B1(n8747), .B2(n8024), .C1(
        n10144), .C2(n7728), .ZN(P2_U3330) );
  NAND2_X1 U9597 ( .A1(n8025), .A2(n8026), .ZN(n8027) );
  XOR2_X1 U9598 ( .A(n8028), .B(n8027), .Z(n8036) );
  NOR2_X1 U9599 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8029), .ZN(n9687) );
  NOR2_X1 U9600 ( .A1(n8865), .A2(n8030), .ZN(n8031) );
  AOI211_X1 U9601 ( .C1(n8868), .C2(n9161), .A(n9687), .B(n8031), .ZN(n8032)
         );
  OAI21_X1 U9602 ( .B1(n8870), .B2(n8033), .A(n8032), .ZN(n8034) );
  AOI21_X1 U9603 ( .B1(n9524), .B2(n8872), .A(n8034), .ZN(n8035) );
  OAI21_X1 U9604 ( .B1(n8036), .B2(n8874), .A(n8035), .ZN(P1_U3213) );
  INV_X1 U9605 ( .A(n8706), .ZN(n8627) );
  INV_X1 U9606 ( .A(n8038), .ZN(n8037) );
  XNOR2_X1 U9607 ( .A(n8706), .B(n8152), .ZN(n8079) );
  NOR2_X1 U9608 ( .A1(n8262), .A2(n8162), .ZN(n8077) );
  XNOR2_X1 U9609 ( .A(n8079), .B(n8077), .ZN(n8039) );
  NOR3_X1 U9610 ( .A1(n4440), .A2(n8037), .A3(n8039), .ZN(n8041) );
  INV_X1 U9611 ( .A(n8081), .ZN(n8040) );
  OAI21_X1 U9612 ( .B1(n8041), .B2(n8040), .A(n8298), .ZN(n8045) );
  OAI22_X1 U9613 ( .A1(n8616), .A2(n8302), .B1(n8304), .B2(n8618), .ZN(n8042)
         );
  AOI211_X1 U9614 ( .C1(n8624), .C2(n8293), .A(n8043), .B(n8042), .ZN(n8044)
         );
  OAI211_X1 U9615 ( .C1(n8627), .C2(n8247), .A(n8045), .B(n8044), .ZN(P2_U3228) );
  INV_X1 U9616 ( .A(n8883), .ZN(n8746) );
  INV_X1 U9617 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8046) );
  OAI222_X1 U9618 ( .A1(n9550), .A2(n8746), .B1(P1_U3084), .B2(n8047), .C1(
        n8046), .C2(n8222), .ZN(P1_U3324) );
  AOI22_X1 U9619 ( .A1(n8061), .A2(P1_STATE_REG_SCAN_IN), .B1(n9548), .B2(
        P2_DATAO_REG_3__SCAN_IN), .ZN(n8048) );
  OAI21_X1 U9620 ( .B1(n8049), .B2(n9550), .A(n8048), .ZN(P1_U3350) );
  INV_X1 U9621 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n8063) );
  OAI21_X1 U9622 ( .B1(n8052), .B2(n8051), .A(n8050), .ZN(n8058) );
  NOR2_X1 U9623 ( .A1(n8054), .A2(n8053), .ZN(n8055) );
  OR3_X1 U9624 ( .A1(n9741), .A2(n8056), .A3(n8055), .ZN(n8057) );
  OAI21_X1 U9625 ( .B1(n9751), .B2(n8058), .A(n8057), .ZN(n8059) );
  AOI211_X1 U9626 ( .C1(n9714), .C2(n8061), .A(n8060), .B(n8059), .ZN(n8062)
         );
  OAI21_X1 U9627 ( .B1(n8063), .B2(n9754), .A(n8062), .ZN(P1_U3244) );
  INV_X1 U9628 ( .A(n8064), .ZN(n8066) );
  OAI21_X1 U9629 ( .B1(n8066), .B2(n8065), .A(n8850), .ZN(n8076) );
  AOI21_X1 U9630 ( .B1(n8064), .B2(n8067), .A(n8068), .ZN(n8075) );
  AND2_X1 U9631 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9703) );
  AOI21_X1 U9632 ( .B1(n8857), .B2(n9158), .A(n9703), .ZN(n8071) );
  NAND2_X1 U9633 ( .A1(n8819), .A2(n8069), .ZN(n8070) );
  OAI211_X1 U9634 ( .C1(n8853), .C2(n8904), .A(n8071), .B(n8070), .ZN(n8072)
         );
  AOI21_X1 U9635 ( .B1(n8073), .B2(n8872), .A(n8072), .ZN(n8074) );
  OAI21_X1 U9636 ( .B1(n8076), .B2(n8075), .A(n8074), .ZN(P1_U3239) );
  INV_X1 U9637 ( .A(n8077), .ZN(n8078) );
  NAND2_X1 U9638 ( .A1(n8079), .A2(n8078), .ZN(n8080) );
  XNOR2_X1 U9639 ( .A(n8703), .B(n8163), .ZN(n8087) );
  NOR2_X1 U9640 ( .A1(n8618), .A2(n8162), .ZN(n8086) );
  XNOR2_X1 U9641 ( .A(n8087), .B(n8086), .ZN(n8286) );
  XNOR2_X1 U9642 ( .A(n8696), .B(n8163), .ZN(n8091) );
  NAND2_X1 U9643 ( .A1(n8589), .A2(n8148), .ZN(n8089) );
  XNOR2_X1 U9644 ( .A(n8091), .B(n8089), .ZN(n8289) );
  INV_X1 U9645 ( .A(n8289), .ZN(n8088) );
  OR2_X1 U9646 ( .A1(n8286), .A2(n8088), .ZN(n8237) );
  XNOR2_X1 U9647 ( .A(n8693), .B(n8152), .ZN(n8082) );
  NAND2_X1 U9648 ( .A1(n8575), .A2(n8148), .ZN(n8083) );
  NAND2_X1 U9649 ( .A1(n8082), .A2(n8083), .ZN(n8241) );
  INV_X1 U9650 ( .A(n8241), .ZN(n8094) );
  INV_X1 U9651 ( .A(n8082), .ZN(n8085) );
  INV_X1 U9652 ( .A(n8083), .ZN(n8084) );
  NAND2_X1 U9653 ( .A1(n8085), .A2(n8084), .ZN(n8243) );
  NAND2_X1 U9654 ( .A1(n8087), .A2(n8086), .ZN(n8287) );
  OR2_X1 U9655 ( .A1(n8088), .A2(n8287), .ZN(n8093) );
  INV_X1 U9656 ( .A(n8089), .ZN(n8090) );
  NAND2_X1 U9657 ( .A1(n8091), .A2(n8090), .ZN(n8092) );
  AND2_X1 U9658 ( .A1(n8093), .A2(n8092), .ZN(n8238) );
  OR2_X1 U9659 ( .A1(n8094), .A2(n8238), .ZN(n8234) );
  AND2_X1 U9660 ( .A1(n8243), .A2(n8234), .ZN(n8095) );
  NAND2_X1 U9661 ( .A1(n8235), .A2(n8095), .ZN(n8104) );
  NOR2_X1 U9662 ( .A1(n8555), .A2(n8162), .ZN(n8096) );
  XNOR2_X1 U9663 ( .A(n8686), .B(n8163), .ZN(n8097) );
  XOR2_X1 U9664 ( .A(n8096), .B(n8097), .Z(n8105) );
  XNOR2_X1 U9665 ( .A(n8521), .B(n8163), .ZN(n8137) );
  NAND2_X1 U9666 ( .A1(n8533), .A2(n8148), .ZN(n8136) );
  XNOR2_X1 U9667 ( .A(n8137), .B(n8136), .ZN(n8138) );
  XNOR2_X1 U9668 ( .A(n8139), .B(n8138), .ZN(n8103) );
  OAI22_X1 U9669 ( .A1(n8301), .A2(n8518), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8099), .ZN(n8101) );
  OAI22_X1 U9670 ( .A1(n8229), .A2(n8304), .B1(n8302), .B2(n8555), .ZN(n8100)
         );
  AOI211_X1 U9671 ( .C1(n8679), .C2(n8308), .A(n8101), .B(n8100), .ZN(n8102)
         );
  OAI21_X1 U9672 ( .B1(n8103), .B2(n8296), .A(n8102), .ZN(P2_U3225) );
  XNOR2_X1 U9673 ( .A(n8104), .B(n8105), .ZN(n8111) );
  INV_X1 U9674 ( .A(n8543), .ZN(n8107) );
  OAI22_X1 U9675 ( .A1(n8301), .A2(n8107), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8106), .ZN(n8109) );
  OAI22_X1 U9676 ( .A1(n8291), .A2(n8302), .B1(n8304), .B2(n8507), .ZN(n8108)
         );
  AOI211_X1 U9677 ( .C1(n8686), .C2(n8308), .A(n8109), .B(n8108), .ZN(n8110)
         );
  OAI21_X1 U9678 ( .B1(n8111), .B2(n8296), .A(n8110), .ZN(P2_U3235) );
  INV_X1 U9679 ( .A(n9493), .ZN(n9377) );
  NAND2_X1 U9680 ( .A1(n8112), .A2(n4927), .ZN(n8114) );
  NAND2_X1 U9681 ( .A1(n8114), .A2(n8113), .ZN(n9417) );
  OR2_X1 U9682 ( .A1(n9509), .A2(n8815), .ZN(n9023) );
  NAND2_X1 U9683 ( .A1(n9509), .A2(n8815), .ZN(n8964) );
  NOR2_X1 U9684 ( .A1(n9501), .A2(n9439), .ZN(n8115) );
  INV_X1 U9685 ( .A(n9439), .ZN(n8866) );
  INV_X1 U9686 ( .A(n9501), .ZN(n9406) );
  INV_X1 U9687 ( .A(n9496), .ZN(n9387) );
  INV_X1 U9688 ( .A(n9409), .ZN(n9368) );
  NOR2_X1 U9689 ( .A1(n9387), .A2(n9368), .ZN(n8116) );
  NAND2_X1 U9690 ( .A1(n9493), .A2(n8854), .ZN(n8892) );
  NAND2_X1 U9691 ( .A1(n9034), .A2(n8892), .ZN(n9366) );
  NAND2_X1 U9692 ( .A1(n4398), .A2(n9366), .ZN(n9360) );
  OAI21_X1 U9693 ( .B1(n9481), .B2(n9354), .A(n9326), .ZN(n8119) );
  NAND2_X1 U9694 ( .A1(n9481), .A2(n9354), .ZN(n8962) );
  NAND2_X1 U9695 ( .A1(n9478), .A2(n8767), .ZN(n8887) );
  INV_X1 U9696 ( .A(n9478), .ZN(n8120) );
  NAND2_X1 U9697 ( .A1(n9472), .A2(n9315), .ZN(n9042) );
  NAND2_X1 U9698 ( .A1(n8121), .A2(n9296), .ZN(n9292) );
  NOR2_X1 U9699 ( .A1(n9465), .A2(n9299), .ZN(n8124) );
  NAND2_X1 U9700 ( .A1(n9465), .A2(n9299), .ZN(n8123) );
  NAND2_X1 U9701 ( .A1(n9460), .A2(n9229), .ZN(n9049) );
  XNOR2_X1 U9702 ( .A(n9227), .B(n9103), .ZN(n9464) );
  INV_X1 U9703 ( .A(n9465), .ZN(n9281) );
  INV_X1 U9704 ( .A(n9509), .ZN(n9424) );
  OR2_X2 U9705 ( .A1(n9398), .A2(n9496), .ZN(n9382) );
  NOR2_X2 U9706 ( .A1(n9382), .A2(n9493), .ZN(n9372) );
  AND2_X2 U9707 ( .A1(n9372), .A2(n9350), .ZN(n9345) );
  AOI21_X1 U9708 ( .B1(n9460), .B2(n9277), .A(n8125), .ZN(n9461) );
  INV_X1 U9709 ( .A(n9460), .ZN(n9230) );
  AOI22_X1 U9710 ( .A1(n8755), .A2(n9402), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9404), .ZN(n8126) );
  OAI21_X1 U9711 ( .B1(n9230), .B2(n9423), .A(n8126), .ZN(n8134) );
  OAI21_X2 U9712 ( .B1(n8127), .B2(n8902), .A(n8888), .ZN(n9432) );
  INV_X1 U9713 ( .A(n9418), .ZN(n9431) );
  INV_X1 U9714 ( .A(n8964), .ZN(n8128) );
  OR2_X1 U9715 ( .A1(n9501), .A2(n8866), .ZN(n9022) );
  NAND2_X1 U9716 ( .A1(n9501), .A2(n8866), .ZN(n9025) );
  NAND2_X1 U9717 ( .A1(n9022), .A2(n9025), .ZN(n9408) );
  NAND2_X1 U9718 ( .A1(n9496), .A2(n9368), .ZN(n9024) );
  NAND2_X1 U9719 ( .A1(n9362), .A2(n9024), .ZN(n9391) );
  INV_X1 U9720 ( .A(n9362), .ZN(n8129) );
  NOR3_X1 U9721 ( .A1(n9361), .A2(n8129), .A3(n9366), .ZN(n9364) );
  INV_X1 U9722 ( .A(n8892), .ZN(n9033) );
  NOR2_X1 U9723 ( .A1(n9364), .A2(n9033), .ZN(n9353) );
  NAND2_X1 U9724 ( .A1(n9486), .A2(n9370), .ZN(n9036) );
  NAND2_X1 U9725 ( .A1(n9353), .A2(n9352), .ZN(n9351) );
  NAND2_X1 U9726 ( .A1(n9351), .A2(n9035), .ZN(n9336) );
  NAND2_X1 U9727 ( .A1(n9481), .A2(n9314), .ZN(n9127) );
  NAND2_X1 U9728 ( .A1(n8897), .A2(n9127), .ZN(n9325) );
  INV_X1 U9729 ( .A(n9325), .ZN(n9335) );
  INV_X1 U9730 ( .A(n8887), .ZN(n9297) );
  INV_X1 U9731 ( .A(n8130), .ZN(n9044) );
  INV_X1 U9732 ( .A(n9299), .ZN(n8794) );
  NAND2_X1 U9733 ( .A1(n9465), .A2(n8794), .ZN(n9048) );
  INV_X1 U9734 ( .A(n8131), .ZN(n9050) );
  NOR2_X2 U9735 ( .A1(n9283), .A2(n9050), .ZN(n8132) );
  NOR2_X1 U9736 ( .A1(n9463), .A2(n9404), .ZN(n8133) );
  OAI21_X1 U9737 ( .B1(n9464), .B2(n9444), .A(n8135), .ZN(P1_U3264) );
  NOR2_X1 U9738 ( .A1(n8508), .A2(n8162), .ZN(n8226) );
  OAI22_X1 U9739 ( .A1(n8139), .A2(n8138), .B1(n8137), .B2(n8136), .ZN(n8142)
         );
  XNOR2_X1 U9740 ( .A(n8674), .B(n8163), .ZN(n8141) );
  INV_X1 U9741 ( .A(n8141), .ZN(n8140) );
  XNOR2_X1 U9742 ( .A(n8142), .B(n8140), .ZN(n8278) );
  NAND2_X1 U9743 ( .A1(n8525), .A2(n8148), .ZN(n8277) );
  NAND2_X1 U9744 ( .A1(n8278), .A2(n8277), .ZN(n8276) );
  XNOR2_X1 U9745 ( .A(n8486), .B(n8163), .ZN(n8143) );
  NAND2_X1 U9746 ( .A1(n8144), .A2(n8143), .ZN(n8223) );
  XNOR2_X1 U9747 ( .A(n8145), .B(n4441), .ZN(n8268) );
  NAND2_X1 U9748 ( .A1(n8492), .A2(n8148), .ZN(n8267) );
  OAI21_X2 U9749 ( .B1(n8268), .B2(n8267), .A(n8146), .ZN(n8250) );
  XNOR2_X1 U9750 ( .A(n8657), .B(n8163), .ZN(n8252) );
  INV_X1 U9751 ( .A(n8303), .ZN(n8433) );
  NAND2_X1 U9752 ( .A1(n8433), .A2(n8148), .ZN(n8251) );
  INV_X1 U9753 ( .A(n8252), .ZN(n8147) );
  XNOR2_X1 U9754 ( .A(n8652), .B(n8152), .ZN(n8150) );
  NAND2_X1 U9755 ( .A1(n8423), .A2(n8148), .ZN(n8149) );
  NOR2_X1 U9756 ( .A1(n8150), .A2(n8149), .ZN(n8151) );
  AOI21_X1 U9757 ( .B1(n8150), .B2(n8149), .A(n8151), .ZN(n8300) );
  XNOR2_X1 U9758 ( .A(n8646), .B(n8152), .ZN(n8154) );
  OR2_X1 U9759 ( .A1(n8305), .A2(n8162), .ZN(n8153) );
  NOR2_X1 U9760 ( .A1(n8154), .A2(n8153), .ZN(n8167) );
  AOI21_X1 U9761 ( .B1(n8154), .B2(n8153), .A(n8167), .ZN(n8155) );
  NAND2_X1 U9762 ( .A1(n8156), .A2(n8155), .ZN(n8177) );
  NOR2_X1 U9763 ( .A1(n8157), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8159) );
  OAI22_X1 U9764 ( .A1(n8202), .A2(n8304), .B1(n8255), .B2(n8302), .ZN(n8158)
         );
  AOI211_X1 U9765 ( .C1(n8293), .C2(n8418), .A(n8159), .B(n8158), .ZN(n8160)
         );
  OAI211_X1 U9766 ( .C1(n4646), .C2(n8247), .A(n8161), .B(n8160), .ZN(P2_U3216) );
  OR2_X1 U9767 ( .A1(n8202), .A2(n8162), .ZN(n8164) );
  XNOR2_X1 U9768 ( .A(n8164), .B(n8163), .ZN(n8165) );
  XNOR2_X1 U9769 ( .A(n8641), .B(n8165), .ZN(n8171) );
  INV_X1 U9770 ( .A(n8171), .ZN(n8166) );
  NAND2_X1 U9771 ( .A1(n8166), .A2(n8298), .ZN(n8178) );
  INV_X1 U9772 ( .A(n8167), .ZN(n8172) );
  NAND4_X1 U9773 ( .A1(n8177), .A2(n8298), .A3(n8172), .A4(n8171), .ZN(n8176)
         );
  INV_X1 U9774 ( .A(n8168), .ZN(n8312) );
  AOI22_X1 U9775 ( .A1(n8434), .A2(n8591), .B1(n8312), .B2(n8590), .ZN(n8407)
         );
  AOI22_X1 U9776 ( .A1(n8403), .A2(n8293), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n8169) );
  OAI21_X1 U9777 ( .B1(n8407), .B2(n8170), .A(n8169), .ZN(n8174) );
  NOR3_X1 U9778 ( .A1(n8172), .A2(n8171), .A3(n8296), .ZN(n8173) );
  AOI211_X1 U9779 ( .C1(n8641), .C2(n8308), .A(n8174), .B(n8173), .ZN(n8175)
         );
  OAI211_X1 U9780 ( .C1(n8178), .C2(n8177), .A(n8176), .B(n8175), .ZN(P2_U3222) );
  INV_X1 U9781 ( .A(n8876), .ZN(n8221) );
  INV_X1 U9782 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8181) );
  NAND3_X1 U9783 ( .A1(n8181), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n8184) );
  NAND2_X1 U9784 ( .A1(n9545), .A2(n9954), .ZN(n8183) );
  NAND2_X1 U9785 ( .A1(n9952), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8182) );
  OAI211_X1 U9786 ( .C1(n5831), .C2(n8184), .A(n8183), .B(n8182), .ZN(P2_U3327) );
  OR2_X1 U9787 ( .A1(n8711), .A2(n8315), .ZN(n8185) );
  NAND2_X1 U9788 ( .A1(n8706), .A2(n8592), .ZN(n8581) );
  AND2_X1 U9789 ( .A1(n8581), .A2(n8187), .ZN(n8188) );
  INV_X1 U9790 ( .A(n8618), .ZN(n8574) );
  OR2_X1 U9791 ( .A1(n8703), .A2(n8574), .ZN(n8189) );
  INV_X1 U9792 ( .A(n8696), .ZN(n8571) );
  AND2_X1 U9793 ( .A1(n8693), .A2(n8575), .ZN(n8535) );
  INV_X1 U9794 ( .A(n8555), .ZN(n8526) );
  AND2_X1 U9795 ( .A1(n8686), .A2(n8526), .ZN(n8191) );
  OR2_X1 U9796 ( .A1(n8535), .A2(n8191), .ZN(n8193) );
  OR2_X1 U9797 ( .A1(n8693), .A2(n8575), .ZN(n8537) );
  AND2_X1 U9798 ( .A1(n8537), .A2(n8190), .ZN(n8536) );
  OR2_X1 U9799 ( .A1(n8191), .A2(n8536), .ZN(n8192) );
  OR2_X1 U9800 ( .A1(n8679), .A2(n8533), .ZN(n8194) );
  NAND2_X1 U9801 ( .A1(n8679), .A2(n8533), .ZN(n8195) );
  NAND2_X1 U9802 ( .A1(n8196), .A2(n8195), .ZN(n8497) );
  NAND2_X1 U9803 ( .A1(n8669), .A2(n8313), .ZN(n8198) );
  OAI21_X1 U9804 ( .B1(n8492), .B2(n8662), .A(n8458), .ZN(n8443) );
  NAND2_X1 U9805 ( .A1(n8443), .A2(n8451), .ZN(n8442) );
  NAND2_X1 U9806 ( .A1(n8442), .A2(n8199), .ZN(n8430) );
  NAND2_X1 U9807 ( .A1(n8430), .A2(n8429), .ZN(n8428) );
  NAND2_X1 U9808 ( .A1(n8428), .A2(n8200), .ZN(n8414) );
  NAND2_X1 U9809 ( .A1(n8414), .A2(n8421), .ZN(n8413) );
  INV_X1 U9810 ( .A(n8202), .ZN(n8422) );
  INV_X1 U9811 ( .A(n8657), .ZN(n8450) );
  INV_X1 U9812 ( .A(n8703), .ZN(n8603) );
  NAND2_X1 U9813 ( .A1(n8499), .A2(n8486), .ZN(n8480) );
  NOR2_X2 U9814 ( .A1(n8641), .A2(n8416), .ZN(n8402) );
  INV_X1 U9815 ( .A(n8402), .ZN(n8205) );
  INV_X1 U9816 ( .A(n8636), .ZN(n8208) );
  AOI21_X1 U9817 ( .B1(n8636), .B2(n8205), .A(n8394), .ZN(n8637) );
  AOI22_X1 U9818 ( .A1(n8206), .A2(n9810), .B1(n8600), .B2(
        P2_REG2_REG_29__SCAN_IN), .ZN(n8207) );
  OAI21_X1 U9819 ( .B1(n8208), .B2(n8626), .A(n8207), .ZN(n8218) );
  XOR2_X1 U9820 ( .A(n8210), .B(n8209), .Z(n8211) );
  INV_X1 U9821 ( .A(n8212), .ZN(n8213) );
  AND2_X1 U9822 ( .A1(n8213), .A2(P2_B_REG_SCAN_IN), .ZN(n8214) );
  NOR2_X1 U9823 ( .A1(n8617), .A2(n8214), .ZN(n8389) );
  AOI22_X1 U9824 ( .A1(n8422), .A2(n8591), .B1(n8389), .B2(n8311), .ZN(n8215)
         );
  AOI211_X1 U9825 ( .C1(n8637), .C2(n8632), .A(n8218), .B(n8217), .ZN(n8219)
         );
  OAI21_X1 U9826 ( .B1(n8640), .B2(n8606), .A(n8219), .ZN(P2_U3267) );
  INV_X1 U9827 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10075) );
  OAI222_X1 U9828 ( .A1(n8222), .A2(n10075), .B1(n9550), .B2(n8221), .C1(n8220), .C2(P1_U3084), .ZN(P1_U3323) );
  INV_X1 U9829 ( .A(n8223), .ZN(n8224) );
  NOR2_X1 U9830 ( .A1(n8225), .A2(n8224), .ZN(n8227) );
  XNOR2_X1 U9831 ( .A(n8227), .B(n8226), .ZN(n8233) );
  OAI22_X1 U9832 ( .A1(n8301), .A2(n8483), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8228), .ZN(n8231) );
  OAI22_X1 U9833 ( .A1(n8254), .A2(n8304), .B1(n8302), .B2(n8229), .ZN(n8230)
         );
  AOI211_X1 U9834 ( .C1(n8669), .C2(n8308), .A(n8231), .B(n8230), .ZN(n8232)
         );
  OAI21_X1 U9835 ( .B1(n8233), .B2(n8296), .A(n8232), .ZN(P2_U3218) );
  OR2_X1 U9836 ( .A1(n8236), .A2(n8237), .ZN(n8239) );
  NAND2_X1 U9837 ( .A1(n8239), .A2(n8238), .ZN(n8240) );
  AOI21_X1 U9838 ( .B1(n8243), .B2(n8241), .A(n8240), .ZN(n8242) );
  AOI211_X1 U9839 ( .C1(n4448), .C2(n8243), .A(n8296), .B(n8242), .ZN(n8249)
         );
  INV_X1 U9840 ( .A(n8693), .ZN(n8561) );
  INV_X1 U9841 ( .A(n8244), .ZN(n8558) );
  AOI22_X1 U9842 ( .A1(n8293), .A2(n8558), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3152), .ZN(n8246) );
  AOI22_X1 U9843 ( .A1(n8280), .A2(n8589), .B1(n8281), .B2(n8526), .ZN(n8245)
         );
  OAI211_X1 U9844 ( .C1(n8561), .C2(n8247), .A(n8246), .B(n8245), .ZN(n8248)
         );
  OR2_X1 U9845 ( .A1(n8249), .A2(n8248), .ZN(P2_U3221) );
  XNOR2_X1 U9846 ( .A(n8252), .B(n8251), .ZN(n8253) );
  XNOR2_X1 U9847 ( .A(n8250), .B(n8253), .ZN(n8260) );
  OAI22_X1 U9848 ( .A1(n8255), .A2(n8617), .B1(n8254), .B2(n8615), .ZN(n8453)
         );
  AOI22_X1 U9849 ( .A1(n8453), .A2(n8271), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8256) );
  OAI21_X1 U9850 ( .B1(n8257), .B2(n8301), .A(n8256), .ZN(n8258) );
  AOI21_X1 U9851 ( .B1(n8657), .B2(n8308), .A(n8258), .ZN(n8259) );
  OAI21_X1 U9852 ( .B1(n8260), .B2(n8296), .A(n8259), .ZN(P2_U3227) );
  XNOR2_X1 U9853 ( .A(n8236), .B(n8286), .ZN(n8266) );
  INV_X1 U9854 ( .A(n8599), .ZN(n8261) );
  OAI22_X1 U9855 ( .A1(n8301), .A2(n8261), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8346), .ZN(n8264) );
  OAI22_X1 U9856 ( .A1(n8262), .A2(n8302), .B1(n8304), .B2(n8554), .ZN(n8263)
         );
  AOI211_X1 U9857 ( .C1(n8703), .C2(n8308), .A(n8264), .B(n8263), .ZN(n8265)
         );
  OAI21_X1 U9858 ( .B1(n8266), .B2(n8296), .A(n8265), .ZN(P2_U3230) );
  XNOR2_X1 U9859 ( .A(n8268), .B(n8267), .ZN(n8275) );
  OR2_X1 U9860 ( .A1(n8303), .A2(n8617), .ZN(n8270) );
  NAND2_X1 U9861 ( .A1(n8313), .A2(n8591), .ZN(n8269) );
  NAND2_X1 U9862 ( .A1(n8270), .A2(n8269), .ZN(n8464) );
  AOI22_X1 U9863 ( .A1(n8464), .A2(n8271), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n8272) );
  OAI21_X1 U9864 ( .B1(n8470), .B2(n8301), .A(n8272), .ZN(n8273) );
  AOI21_X1 U9865 ( .B1(n8662), .B2(n8308), .A(n8273), .ZN(n8274) );
  OAI21_X1 U9866 ( .B1(n8275), .B2(n8296), .A(n8274), .ZN(P2_U3231) );
  OAI21_X1 U9867 ( .B1(n8278), .B2(n8277), .A(n8276), .ZN(n8279) );
  NAND2_X1 U9868 ( .A1(n8279), .A2(n8298), .ZN(n8285) );
  AOI22_X1 U9869 ( .A1(n8293), .A2(n8500), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8284) );
  AOI22_X1 U9870 ( .A1(n8281), .A2(n8313), .B1(n8280), .B2(n8533), .ZN(n8283)
         );
  NAND2_X1 U9871 ( .A1(n8674), .A2(n8308), .ZN(n8282) );
  NAND4_X1 U9872 ( .A1(n8285), .A2(n8284), .A3(n8283), .A4(n8282), .ZN(
        P2_U3237) );
  OR2_X1 U9873 ( .A1(n8236), .A2(n8286), .ZN(n8288) );
  NAND2_X1 U9874 ( .A1(n8288), .A2(n8287), .ZN(n8290) );
  XNOR2_X1 U9875 ( .A(n8290), .B(n8289), .ZN(n8297) );
  AND2_X1 U9876 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8364) );
  OAI22_X1 U9877 ( .A1(n8618), .A2(n8302), .B1(n8304), .B2(n8291), .ZN(n8292)
         );
  AOI211_X1 U9878 ( .C1(n8293), .C2(n8569), .A(n8364), .B(n8292), .ZN(n8295)
         );
  NAND2_X1 U9879 ( .A1(n8696), .A2(n8308), .ZN(n8294) );
  OAI211_X1 U9880 ( .C1(n8297), .C2(n8296), .A(n8295), .B(n8294), .ZN(P2_U3240) );
  OAI211_X1 U9881 ( .C1(n4395), .C2(n8300), .A(n8299), .B(n8298), .ZN(n8310)
         );
  OAI22_X1 U9882 ( .A1(n8301), .A2(n8438), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10169), .ZN(n8307) );
  OAI22_X1 U9883 ( .A1(n8305), .A2(n8304), .B1(n8303), .B2(n8302), .ZN(n8306)
         );
  AOI211_X1 U9884 ( .C1(n8652), .C2(n8308), .A(n8307), .B(n8306), .ZN(n8309)
         );
  NAND2_X1 U9885 ( .A1(n8310), .A2(n8309), .ZN(P2_U3242) );
  MUX2_X1 U9886 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8311), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9887 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8312), .S(P2_U3966), .Z(
        P2_U3581) );
  MUX2_X1 U9888 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8422), .S(P2_U3966), .Z(
        P2_U3580) );
  MUX2_X1 U9889 ( .A(n8423), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8314), .Z(
        P2_U3578) );
  MUX2_X1 U9890 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8433), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U9891 ( .A(n8492), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8314), .Z(
        P2_U3576) );
  MUX2_X1 U9892 ( .A(n8313), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8314), .Z(
        P2_U3575) );
  MUX2_X1 U9893 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8525), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9894 ( .A(n8533), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8314), .Z(
        P2_U3573) );
  MUX2_X1 U9895 ( .A(n8526), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8314), .Z(
        P2_U3572) );
  MUX2_X1 U9896 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8575), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9897 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8589), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9898 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8574), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9899 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8592), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9900 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8315), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9901 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8316), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9902 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8317), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9903 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8318), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U9904 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8319), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U9905 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8320), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U9906 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8321), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U9907 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8322), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U9908 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8323), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U9909 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8324), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U9910 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8325), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U9911 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8326), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U9912 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8327), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U9913 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8328), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U9914 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n6834), .S(P2_U3966), .Z(
        P2_U3553) );
  OAI211_X1 U9915 ( .C1(n8330), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9790), .B(
        n8329), .ZN(n8340) );
  OAI21_X1 U9916 ( .B1(n8333), .B2(n8332), .A(n8331), .ZN(n8334) );
  NAND2_X1 U9917 ( .A1(n8334), .A2(n9791), .ZN(n8339) );
  AOI21_X1 U9918 ( .B1(n9797), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8335), .ZN(
        n8338) );
  NAND2_X1 U9919 ( .A1(n8384), .A2(n8336), .ZN(n8337) );
  NAND4_X1 U9920 ( .A1(n8340), .A2(n8339), .A3(n8338), .A4(n8337), .ZN(
        P2_U3260) );
  NAND2_X1 U9921 ( .A1(n8366), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8343) );
  OAI21_X1 U9922 ( .B1(n8366), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8343), .ZN(
        n8344) );
  AOI211_X1 U9923 ( .C1(n8345), .C2(n8344), .A(n8365), .B(n9792), .ZN(n8355)
         );
  NOR2_X1 U9924 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8346), .ZN(n8347) );
  AOI21_X1 U9925 ( .B1(n9797), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8347), .ZN(
        n8353) );
  INV_X1 U9926 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8349) );
  AOI21_X1 U9927 ( .B1(n4628), .B2(n8349), .A(n8348), .ZN(n8351) );
  XNOR2_X1 U9928 ( .A(n8357), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8350) );
  NAND2_X1 U9929 ( .A1(n8350), .A2(n8351), .ZN(n8356) );
  OAI211_X1 U9930 ( .C1(n8351), .C2(n8350), .A(n9790), .B(n8356), .ZN(n8352)
         );
  OAI211_X1 U9931 ( .C1(n9794), .C2(n8357), .A(n8353), .B(n8352), .ZN(n8354)
         );
  OR2_X1 U9932 ( .A1(n8355), .A2(n8354), .ZN(P2_U3262) );
  INV_X1 U9933 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8358) );
  OAI21_X1 U9934 ( .B1(n8358), .B2(n8357), .A(n8356), .ZN(n8361) );
  INV_X1 U9935 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8359) );
  NAND2_X1 U9936 ( .A1(n8373), .A2(n8359), .ZN(n8378) );
  OAI21_X1 U9937 ( .B1(n8373), .B2(n8359), .A(n8378), .ZN(n8360) );
  NOR2_X1 U9938 ( .A1(n8360), .A2(n8361), .ZN(n8380) );
  AOI21_X1 U9939 ( .B1(n8361), .B2(n8360), .A(n8380), .ZN(n8362) );
  NOR2_X1 U9940 ( .A1(n9795), .A2(n8362), .ZN(n8363) );
  AOI211_X1 U9941 ( .C1(n9797), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n8364), .B(
        n8363), .ZN(n8372) );
  INV_X1 U9942 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8368) );
  NAND2_X1 U9943 ( .A1(n8369), .A2(n8368), .ZN(n8376) );
  OAI21_X1 U9944 ( .B1(n8369), .B2(n8368), .A(n8376), .ZN(n8370) );
  NAND2_X1 U9945 ( .A1(n9791), .A2(n8370), .ZN(n8371) );
  OAI211_X1 U9946 ( .C1(n9794), .C2(n8373), .A(n8372), .B(n8371), .ZN(P2_U3263) );
  NAND2_X1 U9947 ( .A1(n8374), .A2(n8373), .ZN(n8375) );
  NAND2_X1 U9948 ( .A1(n8376), .A2(n8375), .ZN(n8377) );
  XNOR2_X1 U9949 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8377), .ZN(n8383) );
  INV_X1 U9950 ( .A(n8378), .ZN(n8379) );
  NOR2_X1 U9951 ( .A1(n8380), .A2(n8379), .ZN(n8381) );
  XNOR2_X1 U9952 ( .A(n8381), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8385) );
  INV_X1 U9953 ( .A(n8385), .ZN(n8382) );
  AOI22_X1 U9954 ( .A1(n8383), .A2(n9791), .B1(n8382), .B2(n9790), .ZN(n8386)
         );
  NAND2_X1 U9955 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8387) );
  NAND2_X1 U9956 ( .A1(n8395), .A2(n8394), .ZN(n8393) );
  XNOR2_X1 U9957 ( .A(n6359), .B(n8393), .ZN(n8634) );
  NAND2_X1 U9958 ( .A1(n8634), .A2(n8632), .ZN(n8392) );
  NAND2_X1 U9959 ( .A1(n8390), .A2(n8389), .ZN(n9553) );
  NOR2_X1 U9960 ( .A1(n8600), .A2(n9553), .ZN(n8397) );
  AOI21_X1 U9961 ( .B1(n8600), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8397), .ZN(
        n8391) );
  OAI211_X1 U9962 ( .C1(n6359), .C2(n8626), .A(n8392), .B(n8391), .ZN(P2_U3265) );
  OAI21_X1 U9963 ( .B1(n8395), .B2(n8394), .A(n8393), .ZN(n9554) );
  NOR2_X1 U9964 ( .A1(n8395), .A2(n8626), .ZN(n8396) );
  AOI211_X1 U9965 ( .C1(n8600), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8397), .B(
        n8396), .ZN(n8398) );
  OAI21_X1 U9966 ( .B1(n8475), .B2(n9554), .A(n8398), .ZN(P2_U3266) );
  OAI21_X1 U9967 ( .B1(n8400), .B2(n8405), .A(n8399), .ZN(n8401) );
  INV_X1 U9968 ( .A(n8401), .ZN(n8645) );
  AOI21_X1 U9969 ( .B1(n8641), .B2(n8416), .A(n8402), .ZN(n8642) );
  AOI22_X1 U9970 ( .A1(n8403), .A2(n9810), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n8600), .ZN(n8404) );
  OAI21_X1 U9971 ( .B1(n8203), .B2(n8626), .A(n8404), .ZN(n8411) );
  XNOR2_X1 U9972 ( .A(n8406), .B(n8405), .ZN(n8409) );
  INV_X1 U9973 ( .A(n8407), .ZN(n8408) );
  AOI21_X1 U9974 ( .B1(n8409), .B2(n8585), .A(n8408), .ZN(n8644) );
  NOR2_X1 U9975 ( .A1(n8644), .A2(n8600), .ZN(n8410) );
  AOI211_X1 U9976 ( .C1(n8642), .C2(n8632), .A(n8411), .B(n8410), .ZN(n8412)
         );
  OAI21_X1 U9977 ( .B1(n8645), .B2(n8606), .A(n8412), .ZN(P2_U3268) );
  OAI21_X1 U9978 ( .B1(n8414), .B2(n8421), .A(n8413), .ZN(n8415) );
  INV_X1 U9979 ( .A(n8415), .ZN(n8650) );
  INV_X1 U9980 ( .A(n8416), .ZN(n8417) );
  AOI21_X1 U9981 ( .B1(n8646), .B2(n8436), .A(n8417), .ZN(n8647) );
  AOI22_X1 U9982 ( .A1(n8418), .A2(n9810), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n8600), .ZN(n8419) );
  OAI21_X1 U9983 ( .B1(n4646), .B2(n8626), .A(n8419), .ZN(n8426) );
  XOR2_X1 U9984 ( .A(n8421), .B(n8420), .Z(n8424) );
  AOI222_X1 U9985 ( .A1(n8585), .A2(n8424), .B1(n8423), .B2(n8591), .C1(n8422), 
        .C2(n8590), .ZN(n8649) );
  NOR2_X1 U9986 ( .A1(n8649), .A2(n8600), .ZN(n8425) );
  AOI211_X1 U9987 ( .C1(n8647), .C2(n8632), .A(n8426), .B(n8425), .ZN(n8427)
         );
  OAI21_X1 U9988 ( .B1(n8650), .B2(n8606), .A(n8427), .ZN(P2_U3269) );
  OAI21_X1 U9989 ( .B1(n8430), .B2(n8429), .A(n8428), .ZN(n8431) );
  INV_X1 U9990 ( .A(n8431), .ZN(n8655) );
  AOI22_X1 U9991 ( .A1(n8652), .A2(n8473), .B1(n8600), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8441) );
  OAI21_X1 U9992 ( .B1(n4936), .B2(n6167), .A(n8432), .ZN(n8435) );
  AOI222_X1 U9993 ( .A1(n8585), .A2(n8435), .B1(n8434), .B2(n8590), .C1(n8433), 
        .C2(n8591), .ZN(n8654) );
  AOI211_X1 U9994 ( .C1(n8652), .C2(n8445), .A(n9900), .B(n4647), .ZN(n8651)
         );
  NAND2_X1 U9995 ( .A1(n8651), .A2(n6227), .ZN(n8437) );
  OAI211_X1 U9996 ( .C1(n8469), .C2(n8438), .A(n8654), .B(n8437), .ZN(n8439)
         );
  NAND2_X1 U9997 ( .A1(n8439), .A2(n9817), .ZN(n8440) );
  OAI211_X1 U9998 ( .C1(n8655), .C2(n8606), .A(n8441), .B(n8440), .ZN(P2_U3270) );
  OAI21_X1 U9999 ( .B1(n8443), .B2(n8451), .A(n8442), .ZN(n8444) );
  INV_X1 U10000 ( .A(n8444), .ZN(n8660) );
  INV_X1 U10001 ( .A(n8468), .ZN(n8447) );
  INV_X1 U10002 ( .A(n8445), .ZN(n8446) );
  AOI211_X1 U10003 ( .C1(n8657), .C2(n8447), .A(n9900), .B(n8446), .ZN(n8656)
         );
  NOR2_X1 U10004 ( .A1(n8600), .A2(n9812), .ZN(n8598) );
  AOI22_X1 U10005 ( .A1(n8600), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8448), .B2(
        n9810), .ZN(n8449) );
  OAI21_X1 U10006 ( .B1(n8450), .B2(n8626), .A(n8449), .ZN(n8456) );
  XNOR2_X1 U10007 ( .A(n8452), .B(n8451), .ZN(n8454) );
  AOI21_X1 U10008 ( .B1(n8454), .B2(n8585), .A(n8453), .ZN(n8659) );
  NOR2_X1 U10009 ( .A1(n8659), .A2(n8600), .ZN(n8455) );
  AOI211_X1 U10010 ( .C1(n8656), .C2(n8598), .A(n8456), .B(n8455), .ZN(n8457)
         );
  OAI21_X1 U10011 ( .B1(n8660), .B2(n8606), .A(n8457), .ZN(P2_U3271) );
  OAI21_X1 U10012 ( .B1(n8459), .B2(n8460), .A(n8458), .ZN(n8661) );
  INV_X1 U10013 ( .A(n8661), .ZN(n8478) );
  NAND2_X1 U10014 ( .A1(n8461), .A2(n8460), .ZN(n8462) );
  NAND3_X1 U10015 ( .A1(n8463), .A2(n8585), .A3(n8462), .ZN(n8466) );
  INV_X1 U10016 ( .A(n8464), .ZN(n8465) );
  NAND2_X1 U10017 ( .A1(n8466), .A2(n8465), .ZN(n8666) );
  AND2_X1 U10018 ( .A1(n8662), .A2(n8480), .ZN(n8467) );
  OR2_X1 U10019 ( .A1(n8468), .A2(n8467), .ZN(n8664) );
  INV_X1 U10020 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8471) );
  OAI22_X1 U10021 ( .A1(n9817), .A2(n8471), .B1(n8470), .B2(n8469), .ZN(n8472)
         );
  AOI21_X1 U10022 ( .B1(n8662), .B2(n8473), .A(n8472), .ZN(n8474) );
  OAI21_X1 U10023 ( .B1(n8664), .B2(n8475), .A(n8474), .ZN(n8476) );
  AOI21_X1 U10024 ( .B1(n8666), .B2(n9817), .A(n8476), .ZN(n8477) );
  OAI21_X1 U10025 ( .B1(n8478), .B2(n8606), .A(n8477), .ZN(P2_U3272) );
  OAI21_X1 U10026 ( .B1(n4419), .B2(n8488), .A(n8479), .ZN(n8673) );
  INV_X1 U10027 ( .A(n8499), .ZN(n8482) );
  INV_X1 U10028 ( .A(n8480), .ZN(n8481) );
  AOI21_X1 U10029 ( .B1(n8669), .B2(n8482), .A(n8481), .ZN(n8670) );
  INV_X1 U10030 ( .A(n8483), .ZN(n8484) );
  AOI22_X1 U10031 ( .A1(n8600), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8484), .B2(
        n9810), .ZN(n8485) );
  OAI21_X1 U10032 ( .B1(n8486), .B2(n8626), .A(n8485), .ZN(n8495) );
  INV_X1 U10033 ( .A(n8487), .ZN(n8506) );
  OAI21_X1 U10034 ( .B1(n8506), .B2(n8489), .A(n8488), .ZN(n8491) );
  NAND2_X1 U10035 ( .A1(n8491), .A2(n8490), .ZN(n8493) );
  AOI222_X1 U10036 ( .A1(n8585), .A2(n8493), .B1(n8525), .B2(n8591), .C1(n8492), .C2(n8590), .ZN(n8672) );
  NOR2_X1 U10037 ( .A1(n8672), .A2(n8600), .ZN(n8494) );
  AOI211_X1 U10038 ( .C1(n8670), .C2(n8632), .A(n8495), .B(n8494), .ZN(n8496)
         );
  OAI21_X1 U10039 ( .B1(n8606), .B2(n8673), .A(n8496), .ZN(P2_U3273) );
  XNOR2_X1 U10040 ( .A(n8497), .B(n8498), .ZN(n8678) );
  AOI21_X1 U10041 ( .B1(n8674), .B2(n8515), .A(n8499), .ZN(n8675) );
  INV_X1 U10042 ( .A(n8674), .ZN(n8502) );
  AOI22_X1 U10043 ( .A1(n8600), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8500), .B2(
        n9810), .ZN(n8501) );
  OAI21_X1 U10044 ( .B1(n8502), .B2(n8626), .A(n8501), .ZN(n8512) );
  AOI21_X1 U10045 ( .B1(n8522), .B2(n8504), .A(n8503), .ZN(n8505) );
  NOR3_X1 U10046 ( .A1(n8506), .A2(n8505), .A3(n8612), .ZN(n8510) );
  OAI22_X1 U10047 ( .A1(n8508), .A2(n8617), .B1(n8507), .B2(n8615), .ZN(n8509)
         );
  NOR2_X1 U10048 ( .A1(n8510), .A2(n8509), .ZN(n8677) );
  NOR2_X1 U10049 ( .A1(n8677), .A2(n8600), .ZN(n8511) );
  AOI211_X1 U10050 ( .C1(n8675), .C2(n8632), .A(n8512), .B(n8511), .ZN(n8513)
         );
  OAI21_X1 U10051 ( .B1(n8606), .B2(n8678), .A(n8513), .ZN(P2_U3274) );
  XOR2_X1 U10052 ( .A(n8514), .B(n8523), .Z(n8683) );
  INV_X1 U10053 ( .A(n8542), .ZN(n8517) );
  INV_X1 U10054 ( .A(n8515), .ZN(n8516) );
  AOI21_X1 U10055 ( .B1(n8679), .B2(n8517), .A(n8516), .ZN(n8680) );
  INV_X1 U10056 ( .A(n8518), .ZN(n8519) );
  AOI22_X1 U10057 ( .A1(n8600), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8519), .B2(
        n9810), .ZN(n8520) );
  OAI21_X1 U10058 ( .B1(n8521), .B2(n8626), .A(n8520), .ZN(n8529) );
  OAI21_X1 U10059 ( .B1(n8524), .B2(n8523), .A(n8522), .ZN(n8527) );
  AOI222_X1 U10060 ( .A1(n8585), .A2(n8527), .B1(n8526), .B2(n8591), .C1(n8525), .C2(n8590), .ZN(n8682) );
  NOR2_X1 U10061 ( .A1(n8682), .A2(n8600), .ZN(n8528) );
  AOI211_X1 U10062 ( .C1(n8680), .C2(n8632), .A(n8529), .B(n8528), .ZN(n8530)
         );
  OAI21_X1 U10063 ( .B1(n8683), .B2(n8606), .A(n8530), .ZN(P2_U3275) );
  NAND2_X1 U10064 ( .A1(n8549), .A2(n8531), .ZN(n8532) );
  XNOR2_X1 U10065 ( .A(n8532), .B(n8539), .ZN(n8534) );
  AOI222_X1 U10066 ( .A1(n8585), .A2(n8534), .B1(n8533), .B2(n8590), .C1(n8575), .C2(n8591), .ZN(n8689) );
  OR2_X1 U10067 ( .A1(n8548), .A2(n8535), .ZN(n8538) );
  NAND2_X1 U10068 ( .A1(n8538), .A2(n8536), .ZN(n8685) );
  NAND2_X1 U10069 ( .A1(n8538), .A2(n8537), .ZN(n8540) );
  NAND2_X1 U10070 ( .A1(n8540), .A2(n8539), .ZN(n8684) );
  NAND3_X1 U10071 ( .A1(n8685), .A2(n8684), .A3(n8541), .ZN(n8547) );
  AOI21_X1 U10072 ( .B1(n8686), .B2(n8556), .A(n8542), .ZN(n8687) );
  AOI22_X1 U10073 ( .A1(n8600), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8543), .B2(
        n9810), .ZN(n8544) );
  OAI21_X1 U10074 ( .B1(n4648), .B2(n8626), .A(n8544), .ZN(n8545) );
  AOI21_X1 U10075 ( .B1(n8687), .B2(n8632), .A(n8545), .ZN(n8546) );
  OAI211_X1 U10076 ( .C1(n8600), .C2(n8689), .A(n8547), .B(n8546), .ZN(
        P2_U3276) );
  XNOR2_X1 U10077 ( .A(n8548), .B(n8551), .ZN(n8695) );
  INV_X1 U10078 ( .A(n8549), .ZN(n8550) );
  AOI21_X1 U10079 ( .B1(n8552), .B2(n8551), .A(n8550), .ZN(n8553) );
  OAI222_X1 U10080 ( .A1(n8617), .A2(n8555), .B1(n8615), .B2(n8554), .C1(n8612), .C2(n8553), .ZN(n8691) );
  INV_X1 U10081 ( .A(n8556), .ZN(n8557) );
  AOI211_X1 U10082 ( .C1(n8693), .C2(n8566), .A(n9900), .B(n8557), .ZN(n8692)
         );
  NAND2_X1 U10083 ( .A1(n8692), .A2(n8598), .ZN(n8560) );
  AOI22_X1 U10084 ( .A1(n8600), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8558), .B2(
        n9810), .ZN(n8559) );
  OAI211_X1 U10085 ( .C1(n8561), .C2(n8626), .A(n8560), .B(n8559), .ZN(n8562)
         );
  AOI21_X1 U10086 ( .B1(n8691), .B2(n9817), .A(n8562), .ZN(n8563) );
  OAI21_X1 U10087 ( .B1(n8695), .B2(n8606), .A(n8563), .ZN(P2_U3277) );
  XNOR2_X1 U10088 ( .A(n8565), .B(n8564), .ZN(n8700) );
  INV_X1 U10089 ( .A(n8596), .ZN(n8568) );
  INV_X1 U10090 ( .A(n8566), .ZN(n8567) );
  AOI21_X1 U10091 ( .B1(n8696), .B2(n8568), .A(n8567), .ZN(n8697) );
  AOI22_X1 U10092 ( .A1(n8600), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8569), .B2(
        n9810), .ZN(n8570) );
  OAI21_X1 U10093 ( .B1(n8571), .B2(n8626), .A(n8570), .ZN(n8578) );
  XNOR2_X1 U10094 ( .A(n8572), .B(n8573), .ZN(n8576) );
  AOI222_X1 U10095 ( .A1(n8585), .A2(n8576), .B1(n8575), .B2(n8590), .C1(n8574), .C2(n8591), .ZN(n8699) );
  NOR2_X1 U10096 ( .A1(n8699), .A2(n8600), .ZN(n8577) );
  AOI211_X1 U10097 ( .C1(n8697), .C2(n8632), .A(n8578), .B(n8577), .ZN(n8579)
         );
  OAI21_X1 U10098 ( .B1(n8606), .B2(n8700), .A(n8579), .ZN(P2_U3278) );
  NAND2_X1 U10099 ( .A1(n8580), .A2(n8581), .ZN(n8584) );
  INV_X1 U10100 ( .A(n8582), .ZN(n8583) );
  AOI21_X1 U10101 ( .B1(n8587), .B2(n8584), .A(n8583), .ZN(n8705) );
  NAND2_X1 U10102 ( .A1(n8586), .A2(n8585), .ZN(n8595) );
  AOI21_X1 U10103 ( .B1(n8614), .B2(n8588), .A(n8587), .ZN(n8594) );
  AOI22_X1 U10104 ( .A1(n8592), .A2(n8591), .B1(n8590), .B2(n8589), .ZN(n8593)
         );
  OAI21_X1 U10105 ( .B1(n8595), .B2(n8594), .A(n8593), .ZN(n8701) );
  INV_X1 U10106 ( .A(n8622), .ZN(n8597) );
  AOI211_X1 U10107 ( .C1(n8703), .C2(n8597), .A(n9900), .B(n8596), .ZN(n8702)
         );
  NAND2_X1 U10108 ( .A1(n8702), .A2(n8598), .ZN(n8602) );
  AOI22_X1 U10109 ( .A1(n8600), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8599), .B2(
        n9810), .ZN(n8601) );
  OAI211_X1 U10110 ( .C1(n8603), .C2(n8626), .A(n8602), .B(n8601), .ZN(n8604)
         );
  AOI21_X1 U10111 ( .B1(n8701), .B2(n9817), .A(n8604), .ZN(n8605) );
  OAI21_X1 U10112 ( .B1(n8705), .B2(n8606), .A(n8605), .ZN(P2_U3279) );
  INV_X1 U10113 ( .A(n8580), .ZN(n8607) );
  AOI21_X1 U10114 ( .B1(n8609), .B2(n8608), .A(n8607), .ZN(n8628) );
  NAND2_X1 U10115 ( .A1(n8611), .A2(n8610), .ZN(n8613) );
  AOI21_X1 U10116 ( .B1(n8614), .B2(n8613), .A(n8612), .ZN(n8620) );
  OAI22_X1 U10117 ( .A1(n8618), .A2(n8617), .B1(n8616), .B2(n8615), .ZN(n8619)
         );
  AOI211_X1 U10118 ( .C1(n8628), .C2(n8621), .A(n8620), .B(n8619), .ZN(n8709)
         );
  AOI21_X1 U10119 ( .B1(n8706), .B2(n8623), .A(n8622), .ZN(n8707) );
  AOI22_X1 U10120 ( .A1(n8600), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8624), .B2(
        n9810), .ZN(n8625) );
  OAI21_X1 U10121 ( .B1(n8627), .B2(n8626), .A(n8625), .ZN(n8631) );
  INV_X1 U10122 ( .A(n8628), .ZN(n8710) );
  NOR2_X1 U10123 ( .A1(n8710), .A2(n8629), .ZN(n8630) );
  AOI211_X1 U10124 ( .C1(n8707), .C2(n8632), .A(n8631), .B(n8630), .ZN(n8633)
         );
  OAI21_X1 U10125 ( .B1(n8600), .B2(n8709), .A(n8633), .ZN(P2_U3280) );
  INV_X1 U10126 ( .A(n9868), .ZN(n9898) );
  NAND2_X1 U10127 ( .A1(n8634), .A2(n9869), .ZN(n8635) );
  OAI211_X1 U10128 ( .C1(n6359), .C2(n9898), .A(n8635), .B(n9553), .ZN(n8727)
         );
  MUX2_X1 U10129 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8727), .S(n9914), .Z(
        P2_U3551) );
  AOI22_X1 U10130 ( .A1(n8637), .A2(n9869), .B1(n9868), .B2(n8636), .ZN(n8638)
         );
  OAI211_X1 U10131 ( .C1(n8640), .C2(n8720), .A(n8639), .B(n8638), .ZN(n8728)
         );
  MUX2_X1 U10132 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8728), .S(n9914), .Z(
        P2_U3549) );
  AOI22_X1 U10133 ( .A1(n8642), .A2(n9869), .B1(n9868), .B2(n8641), .ZN(n8643)
         );
  OAI211_X1 U10134 ( .C1(n8645), .C2(n8720), .A(n8644), .B(n8643), .ZN(n8729)
         );
  MUX2_X1 U10135 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8729), .S(n9914), .Z(
        P2_U3548) );
  AOI22_X1 U10136 ( .A1(n8647), .A2(n9869), .B1(n9868), .B2(n8646), .ZN(n8648)
         );
  OAI211_X1 U10137 ( .C1(n8650), .C2(n8720), .A(n8649), .B(n8648), .ZN(n8730)
         );
  MUX2_X1 U10138 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8730), .S(n9914), .Z(
        P2_U3547) );
  AOI21_X1 U10139 ( .B1(n9868), .B2(n8652), .A(n8651), .ZN(n8653) );
  OAI211_X1 U10140 ( .C1(n8655), .C2(n8720), .A(n8654), .B(n8653), .ZN(n8731)
         );
  MUX2_X1 U10141 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8731), .S(n9914), .Z(
        P2_U3546) );
  AOI21_X1 U10142 ( .B1(n9868), .B2(n8657), .A(n8656), .ZN(n8658) );
  OAI211_X1 U10143 ( .C1(n8660), .C2(n8720), .A(n8659), .B(n8658), .ZN(n8732)
         );
  MUX2_X1 U10144 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8732), .S(n9922), .Z(
        P2_U3545) );
  NAND2_X1 U10145 ( .A1(n8661), .A2(n9904), .ZN(n8668) );
  INV_X1 U10146 ( .A(n8662), .ZN(n8663) );
  OAI22_X1 U10147 ( .A1(n8664), .A2(n9900), .B1(n8663), .B2(n9898), .ZN(n8665)
         );
  NOR2_X1 U10148 ( .A1(n8666), .A2(n8665), .ZN(n8667) );
  NAND2_X1 U10149 ( .A1(n8668), .A2(n8667), .ZN(n8733) );
  MUX2_X1 U10150 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8733), .S(n9922), .Z(
        P2_U3544) );
  AOI22_X1 U10151 ( .A1(n8670), .A2(n9869), .B1(n9868), .B2(n8669), .ZN(n8671)
         );
  OAI211_X1 U10152 ( .C1(n8673), .C2(n8720), .A(n8672), .B(n8671), .ZN(n8734)
         );
  MUX2_X1 U10153 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8734), .S(n9922), .Z(
        P2_U3543) );
  AOI22_X1 U10154 ( .A1(n8675), .A2(n9869), .B1(n9868), .B2(n8674), .ZN(n8676)
         );
  OAI211_X1 U10155 ( .C1(n8678), .C2(n8720), .A(n8677), .B(n8676), .ZN(n8735)
         );
  MUX2_X1 U10156 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8735), .S(n9922), .Z(
        P2_U3542) );
  AOI22_X1 U10157 ( .A1(n8680), .A2(n9869), .B1(n9868), .B2(n8679), .ZN(n8681)
         );
  OAI211_X1 U10158 ( .C1(n8683), .C2(n8720), .A(n8682), .B(n8681), .ZN(n8736)
         );
  MUX2_X1 U10159 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8736), .S(n9922), .Z(
        P2_U3541) );
  NAND3_X1 U10160 ( .A1(n8685), .A2(n9904), .A3(n8684), .ZN(n8690) );
  AOI22_X1 U10161 ( .A1(n8687), .A2(n9869), .B1(n9868), .B2(n8686), .ZN(n8688)
         );
  NAND3_X1 U10162 ( .A1(n8690), .A2(n8689), .A3(n8688), .ZN(n8737) );
  MUX2_X1 U10163 ( .A(n8737), .B(P2_REG1_REG_20__SCAN_IN), .S(n9919), .Z(
        P2_U3540) );
  AOI211_X1 U10164 ( .C1(n9868), .C2(n8693), .A(n8692), .B(n8691), .ZN(n8694)
         );
  OAI21_X1 U10165 ( .B1(n8720), .B2(n8695), .A(n8694), .ZN(n8738) );
  MUX2_X1 U10166 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8738), .S(n9914), .Z(
        P2_U3539) );
  AOI22_X1 U10167 ( .A1(n8697), .A2(n9869), .B1(n9868), .B2(n8696), .ZN(n8698)
         );
  OAI211_X1 U10168 ( .C1(n8700), .C2(n8720), .A(n8699), .B(n8698), .ZN(n8739)
         );
  MUX2_X1 U10169 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8739), .S(n9914), .Z(
        P2_U3538) );
  AOI211_X1 U10170 ( .C1(n9868), .C2(n8703), .A(n8702), .B(n8701), .ZN(n8704)
         );
  OAI21_X1 U10171 ( .B1(n8705), .B2(n8720), .A(n8704), .ZN(n8740) );
  MUX2_X1 U10172 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8740), .S(n9914), .Z(
        P2_U3537) );
  AOI22_X1 U10173 ( .A1(n8707), .A2(n9869), .B1(n9868), .B2(n8706), .ZN(n8708)
         );
  OAI211_X1 U10174 ( .C1(n9883), .C2(n8710), .A(n8709), .B(n8708), .ZN(n8741)
         );
  MUX2_X1 U10175 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8741), .S(n9914), .Z(
        P2_U3536) );
  AOI22_X1 U10176 ( .A1(n8712), .A2(n9869), .B1(n9868), .B2(n8711), .ZN(n8713)
         );
  OAI211_X1 U10177 ( .C1(n8715), .C2(n8720), .A(n8714), .B(n8713), .ZN(n8742)
         );
  MUX2_X1 U10178 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8742), .S(n9914), .Z(
        P2_U3535) );
  AOI22_X1 U10179 ( .A1(n8717), .A2(n9869), .B1(n9868), .B2(n8716), .ZN(n8718)
         );
  OAI211_X1 U10180 ( .C1(n8721), .C2(n8720), .A(n8719), .B(n8718), .ZN(n8743)
         );
  MUX2_X1 U10181 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8743), .S(n9914), .Z(
        P2_U3534) );
  AOI22_X1 U10182 ( .A1(n8723), .A2(n9869), .B1(n9868), .B2(n8722), .ZN(n8724)
         );
  OAI211_X1 U10183 ( .C1(n9883), .C2(n8726), .A(n8725), .B(n8724), .ZN(n8744)
         );
  MUX2_X1 U10184 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8744), .S(n9914), .Z(
        P2_U3533) );
  MUX2_X1 U10185 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8727), .S(n9908), .Z(
        P2_U3519) );
  MUX2_X1 U10186 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8728), .S(n9908), .Z(
        P2_U3517) );
  MUX2_X1 U10187 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8729), .S(n9908), .Z(
        P2_U3516) );
  MUX2_X1 U10188 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8730), .S(n9908), .Z(
        P2_U3515) );
  MUX2_X1 U10189 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8731), .S(n9908), .Z(
        P2_U3514) );
  MUX2_X1 U10190 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8732), .S(n9908), .Z(
        P2_U3513) );
  MUX2_X1 U10191 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8733), .S(n9908), .Z(
        P2_U3512) );
  MUX2_X1 U10192 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8734), .S(n9908), .Z(
        P2_U3511) );
  MUX2_X1 U10193 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8735), .S(n9908), .Z(
        P2_U3510) );
  MUX2_X1 U10194 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8736), .S(n9908), .Z(
        P2_U3509) );
  MUX2_X1 U10195 ( .A(n8737), .B(P2_REG0_REG_20__SCAN_IN), .S(n9906), .Z(
        P2_U3508) );
  MUX2_X1 U10196 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8738), .S(n9908), .Z(
        P2_U3507) );
  MUX2_X1 U10197 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8739), .S(n9908), .Z(
        P2_U3505) );
  MUX2_X1 U10198 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8740), .S(n9908), .Z(
        P2_U3502) );
  MUX2_X1 U10199 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8741), .S(n9908), .Z(
        P2_U3499) );
  MUX2_X1 U10200 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8742), .S(n9908), .Z(
        P2_U3496) );
  MUX2_X1 U10201 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8743), .S(n9908), .Z(
        P2_U3493) );
  MUX2_X1 U10202 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8744), .S(n9908), .Z(
        P2_U3490) );
  OAI222_X1 U10203 ( .A1(n8749), .A2(P2_U3152), .B1(n8747), .B2(n8746), .C1(
        n8745), .C2(n7728), .ZN(P2_U3329) );
  MUX2_X1 U10204 ( .A(n8750), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NAND2_X1 U10205 ( .A1(n8752), .A2(n8751), .ZN(n8753) );
  XNOR2_X1 U10206 ( .A(n8754), .B(n8753), .ZN(n8760) );
  AOI22_X1 U10207 ( .A1(n9299), .A2(n8868), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n8757) );
  NAND2_X1 U10208 ( .A1(n8755), .A2(n8819), .ZN(n8756) );
  OAI211_X1 U10209 ( .C1(n9242), .C2(n8865), .A(n8757), .B(n8756), .ZN(n8758)
         );
  AOI21_X1 U10210 ( .B1(n9460), .B2(n8872), .A(n8758), .ZN(n8759) );
  OAI21_X1 U10211 ( .B1(n8760), .B2(n8874), .A(n8759), .ZN(P1_U3212) );
  INV_X1 U10212 ( .A(n8761), .ZN(n8763) );
  NOR2_X1 U10213 ( .A1(n8763), .A2(n8762), .ZN(n8765) );
  XNOR2_X1 U10214 ( .A(n8765), .B(n8764), .ZN(n8771) );
  NOR2_X1 U10215 ( .A1(n9330), .A2(n8870), .ZN(n8769) );
  AOI22_X1 U10216 ( .A1(n9337), .A2(n8868), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8766) );
  OAI21_X1 U10217 ( .B1(n8767), .B2(n8865), .A(n8766), .ZN(n8768) );
  AOI211_X1 U10218 ( .C1(n9481), .C2(n8872), .A(n8769), .B(n8768), .ZN(n8770)
         );
  OAI21_X1 U10219 ( .B1(n8771), .B2(n8874), .A(n8770), .ZN(P1_U3214) );
  INV_X1 U10220 ( .A(n8773), .ZN(n8774) );
  AOI21_X1 U10221 ( .B1(n8775), .B2(n8772), .A(n8774), .ZN(n8780) );
  NAND2_X1 U10222 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9213) );
  OAI21_X1 U10223 ( .B1(n9368), .B2(n8865), .A(n9213), .ZN(n8776) );
  AOI21_X1 U10224 ( .B1(n8868), .B2(n9410), .A(n8776), .ZN(n8777) );
  OAI21_X1 U10225 ( .B1(n8870), .B2(n9401), .A(n8777), .ZN(n8778) );
  AOI21_X1 U10226 ( .B1(n9501), .B2(n8872), .A(n8778), .ZN(n8779) );
  OAI21_X1 U10227 ( .B1(n8780), .B2(n8874), .A(n8779), .ZN(P1_U3217) );
  NAND2_X1 U10228 ( .A1(n8781), .A2(n8783), .ZN(n8782) );
  OAI21_X1 U10229 ( .B1(n8783), .B2(n8781), .A(n8782), .ZN(n8784) );
  NAND2_X1 U10230 ( .A1(n8784), .A2(n8850), .ZN(n8789) );
  NOR2_X1 U10231 ( .A1(n8870), .A2(n9373), .ZN(n8787) );
  OAI22_X1 U10232 ( .A1(n9370), .A2(n8865), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8785), .ZN(n8786) );
  AOI211_X1 U10233 ( .C1(n8868), .C2(n9409), .A(n8787), .B(n8786), .ZN(n8788)
         );
  OAI211_X1 U10234 ( .C1(n9377), .C2(n8860), .A(n8789), .B(n8788), .ZN(
        P1_U3221) );
  XOR2_X1 U10235 ( .A(n8791), .B(n8790), .Z(n8797) );
  AOI22_X1 U10236 ( .A1(n9338), .A2(n8868), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8793) );
  NAND2_X1 U10237 ( .A1(n9303), .A2(n8819), .ZN(n8792) );
  OAI211_X1 U10238 ( .C1(n8794), .C2(n8865), .A(n8793), .B(n8792), .ZN(n8795)
         );
  AOI21_X1 U10239 ( .B1(n9472), .B2(n8872), .A(n8795), .ZN(n8796) );
  OAI21_X1 U10240 ( .B1(n8797), .B2(n8874), .A(n8796), .ZN(P1_U3223) );
  XOR2_X1 U10241 ( .A(n8800), .B(n8799), .Z(n8801) );
  XNOR2_X1 U10242 ( .A(n8798), .B(n8801), .ZN(n8809) );
  NOR2_X1 U10243 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8802), .ZN(n9713) );
  NOR2_X1 U10244 ( .A1(n8865), .A2(n8803), .ZN(n8804) );
  AOI211_X1 U10245 ( .C1(n8868), .C2(n9159), .A(n9713), .B(n8804), .ZN(n8805)
         );
  OAI21_X1 U10246 ( .B1(n8870), .B2(n8806), .A(n8805), .ZN(n8807) );
  AOI21_X1 U10247 ( .B1(n9519), .B2(n8872), .A(n8807), .ZN(n8808) );
  OAI21_X1 U10248 ( .B1(n8809), .B2(n8874), .A(n8808), .ZN(P1_U3224) );
  INV_X1 U10249 ( .A(n8811), .ZN(n8812) );
  AOI21_X1 U10250 ( .B1(n8813), .B2(n8810), .A(n8812), .ZN(n8822) );
  NAND2_X1 U10251 ( .A1(n8868), .A2(n9158), .ZN(n8814) );
  NAND2_X1 U10252 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9726) );
  OAI211_X1 U10253 ( .C1(n8815), .C2(n8865), .A(n8814), .B(n9726), .ZN(n8818)
         );
  NOR2_X1 U10254 ( .A1(n8816), .A2(n8860), .ZN(n8817) );
  AOI211_X1 U10255 ( .C1(n8820), .C2(n8819), .A(n8818), .B(n8817), .ZN(n8821)
         );
  OAI21_X1 U10256 ( .B1(n8822), .B2(n8874), .A(n8821), .ZN(P1_U3226) );
  XOR2_X1 U10257 ( .A(n8824), .B(n8823), .Z(n8829) );
  NOR2_X1 U10258 ( .A1(n9315), .A2(n8865), .ZN(n8827) );
  AOI22_X1 U10259 ( .A1(n9354), .A2(n8868), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8825) );
  OAI21_X1 U10260 ( .B1(n8870), .B2(n9310), .A(n8825), .ZN(n8826) );
  AOI211_X1 U10261 ( .C1(n9478), .C2(n8872), .A(n8827), .B(n8826), .ZN(n8828)
         );
  OAI21_X1 U10262 ( .B1(n8829), .B2(n8874), .A(n8828), .ZN(P1_U3227) );
  INV_X1 U10263 ( .A(n8830), .ZN(n8835) );
  AOI21_X1 U10264 ( .B1(n8834), .B2(n8832), .A(n8831), .ZN(n8833) );
  AOI21_X1 U10265 ( .B1(n8835), .B2(n8834), .A(n8833), .ZN(n8840) );
  AOI22_X1 U10266 ( .A1(n9388), .A2(n8857), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8837) );
  NAND2_X1 U10267 ( .A1(n8868), .A2(n9439), .ZN(n8836) );
  OAI211_X1 U10268 ( .C1(n8870), .C2(n9384), .A(n8837), .B(n8836), .ZN(n8838)
         );
  AOI21_X1 U10269 ( .B1(n9496), .B2(n8872), .A(n8838), .ZN(n8839) );
  OAI21_X1 U10270 ( .B1(n8840), .B2(n8874), .A(n8839), .ZN(P1_U3231) );
  AND2_X1 U10271 ( .A1(n8842), .A2(n8841), .ZN(n8843) );
  AOI21_X1 U10272 ( .B1(n8846), .B2(n8843), .A(n8845), .ZN(n8849) );
  INV_X1 U10273 ( .A(n8844), .ZN(n8848) );
  INV_X1 U10274 ( .A(n8845), .ZN(n8847) );
  OAI22_X1 U10275 ( .A1(n8849), .A2(n8848), .B1(n8847), .B2(n8846), .ZN(n8851)
         );
  NAND2_X1 U10276 ( .A1(n8851), .A2(n8850), .ZN(n8859) );
  NOR2_X1 U10277 ( .A1(n8870), .A2(n9347), .ZN(n8856) );
  OAI22_X1 U10278 ( .A1(n8854), .A2(n8853), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8852), .ZN(n8855) );
  AOI211_X1 U10279 ( .C1(n8857), .C2(n9354), .A(n8856), .B(n8855), .ZN(n8858)
         );
  OAI211_X1 U10280 ( .C1(n9350), .C2(n8860), .A(n8859), .B(n8858), .ZN(
        P1_U3233) );
  NAND2_X1 U10281 ( .A1(n8862), .A2(n8861), .ZN(n8863) );
  XOR2_X1 U10282 ( .A(n8864), .B(n8863), .Z(n8875) );
  NAND2_X1 U10283 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9742) );
  OAI21_X1 U10284 ( .B1(n8866), .B2(n8865), .A(n9742), .ZN(n8867) );
  AOI21_X1 U10285 ( .B1(n8868), .B2(n9436), .A(n8867), .ZN(n8869) );
  OAI21_X1 U10286 ( .B1(n8870), .B2(n9426), .A(n8869), .ZN(n8871) );
  AOI21_X1 U10287 ( .B1(n9509), .B2(n8872), .A(n8871), .ZN(n8873) );
  OAI21_X1 U10288 ( .B1(n8875), .B2(n8874), .A(n8873), .ZN(P1_U3236) );
  NAND2_X1 U10289 ( .A1(n8876), .A2(n8882), .ZN(n8878) );
  NAND2_X1 U10290 ( .A1(n5614), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8877) );
  NOR2_X1 U10291 ( .A1(n9563), .A2(n9240), .ZN(n8956) );
  INV_X1 U10292 ( .A(n8956), .ZN(n8881) );
  NAND2_X1 U10293 ( .A1(n5614), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8879) );
  NAND2_X1 U10294 ( .A1(n8881), .A2(n9066), .ZN(n9107) );
  INV_X1 U10295 ( .A(n9107), .ZN(n8954) );
  NAND2_X1 U10296 ( .A1(n8883), .A2(n8882), .ZN(n8885) );
  NAND2_X1 U10297 ( .A1(n5614), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8884) );
  NOR2_X1 U10298 ( .A1(n9450), .A2(n9156), .ZN(n9056) );
  INV_X1 U10299 ( .A(n9074), .ZN(n8886) );
  OR2_X1 U10300 ( .A1(n9056), .A2(n8886), .ZN(n8947) );
  NAND2_X1 U10301 ( .A1(n9042), .A2(n8887), .ZN(n9130) );
  INV_X1 U10302 ( .A(n9130), .ZN(n8942) );
  INV_X1 U10303 ( .A(n9035), .ZN(n8896) );
  NAND2_X1 U10304 ( .A1(n9023), .A2(n8888), .ZN(n8965) );
  INV_X1 U10305 ( .A(n8965), .ZN(n8890) );
  AND2_X1 U10306 ( .A1(n9025), .A2(n8964), .ZN(n9027) );
  INV_X1 U10307 ( .A(n9027), .ZN(n8889) );
  AND2_X1 U10308 ( .A1(n9362), .A2(n9022), .ZN(n9029) );
  OAI211_X1 U10309 ( .C1(n8890), .C2(n8889), .A(n9034), .B(n9029), .ZN(n8895)
         );
  INV_X1 U10310 ( .A(n9024), .ZN(n8891) );
  NAND2_X1 U10311 ( .A1(n9034), .A2(n8891), .ZN(n8893) );
  AND2_X1 U10312 ( .A1(n8893), .A2(n8892), .ZN(n8894) );
  NAND2_X1 U10313 ( .A1(n9036), .A2(n8894), .ZN(n8900) );
  NAND2_X1 U10314 ( .A1(n8900), .A2(n9035), .ZN(n9037) );
  OAI21_X1 U10315 ( .B1(n8896), .B2(n8895), .A(n9037), .ZN(n8898) );
  NAND2_X1 U10316 ( .A1(n8898), .A2(n8897), .ZN(n9128) );
  INV_X1 U10317 ( .A(n9025), .ZN(n8899) );
  OR2_X1 U10318 ( .A1(n8900), .A2(n8899), .ZN(n9124) );
  INV_X1 U10319 ( .A(n9017), .ZN(n8901) );
  NOR2_X1 U10320 ( .A1(n8902), .A2(n8901), .ZN(n8903) );
  NAND2_X1 U10321 ( .A1(n8903), .A2(n8964), .ZN(n8934) );
  NAND2_X1 U10322 ( .A1(n9524), .A2(n8904), .ZN(n8995) );
  NAND2_X1 U10323 ( .A1(n8995), .A2(n8999), .ZN(n9005) );
  INV_X1 U10324 ( .A(n9005), .ZN(n8929) );
  NAND2_X1 U10325 ( .A1(n8989), .A2(n8905), .ZN(n8997) );
  NAND2_X1 U10326 ( .A1(n8981), .A2(n8975), .ZN(n8906) );
  NOR2_X1 U10327 ( .A1(n8997), .A2(n8906), .ZN(n8907) );
  NAND3_X1 U10328 ( .A1(n9014), .A2(n8929), .A3(n8907), .ZN(n8908) );
  NOR2_X1 U10329 ( .A1(n8934), .A2(n8908), .ZN(n9121) );
  INV_X1 U10330 ( .A(n9121), .ZN(n8936) );
  INV_X1 U10331 ( .A(n8909), .ZN(n8911) );
  NAND2_X1 U10332 ( .A1(n6974), .A2(n6975), .ZN(n8910) );
  NAND3_X1 U10333 ( .A1(n8911), .A2(n9140), .A3(n8910), .ZN(n8912) );
  NAND2_X1 U10334 ( .A1(n8913), .A2(n8912), .ZN(n8915) );
  OAI21_X1 U10335 ( .B1(n7163), .B2(n8915), .A(n8914), .ZN(n8917) );
  NAND2_X1 U10336 ( .A1(n8917), .A2(n8916), .ZN(n8918) );
  NAND2_X1 U10337 ( .A1(n8918), .A2(n9120), .ZN(n8920) );
  INV_X1 U10338 ( .A(n8972), .ZN(n9123) );
  AOI21_X1 U10339 ( .B1(n8920), .B2(n8919), .A(n9123), .ZN(n8935) );
  NAND2_X1 U10340 ( .A1(n8996), .A2(n8921), .ZN(n8922) );
  NAND2_X1 U10341 ( .A1(n8922), .A2(n8989), .ZN(n8923) );
  AND2_X1 U10342 ( .A1(n9003), .A2(n8923), .ZN(n9000) );
  INV_X1 U10343 ( .A(n8924), .ZN(n8985) );
  NOR2_X1 U10344 ( .A1(n8987), .A2(n8985), .ZN(n8979) );
  INV_X1 U10345 ( .A(n8981), .ZN(n8925) );
  OR3_X1 U10346 ( .A1(n8997), .A2(n8979), .A3(n8925), .ZN(n8926) );
  NAND2_X1 U10347 ( .A1(n9000), .A2(n8926), .ZN(n8928) );
  INV_X1 U10348 ( .A(n9004), .ZN(n8927) );
  AOI21_X1 U10349 ( .B1(n8929), .B2(n8928), .A(n8927), .ZN(n8931) );
  INV_X1 U10350 ( .A(n9014), .ZN(n8930) );
  OAI211_X1 U10351 ( .C1(n8931), .C2(n8930), .A(n9018), .B(n9013), .ZN(n8932)
         );
  INV_X1 U10352 ( .A(n8932), .ZN(n8933) );
  OR2_X1 U10353 ( .A1(n8934), .A2(n8933), .ZN(n9126) );
  OAI21_X1 U10354 ( .B1(n8936), .B2(n8935), .A(n9126), .ZN(n8937) );
  INV_X1 U10355 ( .A(n8937), .ZN(n8938) );
  NOR2_X1 U10356 ( .A1(n9124), .A2(n8938), .ZN(n8939) );
  OAI21_X1 U10357 ( .B1(n9128), .B2(n8939), .A(n9127), .ZN(n8940) );
  NAND2_X1 U10358 ( .A1(n8940), .A2(n9132), .ZN(n8941) );
  NAND2_X1 U10359 ( .A1(n8942), .A2(n8941), .ZN(n8943) );
  NAND2_X1 U10360 ( .A1(n9228), .A2(n8943), .ZN(n8951) );
  NAND2_X1 U10361 ( .A1(n9455), .A2(n9242), .ZN(n9236) );
  NAND2_X1 U10362 ( .A1(n9236), .A2(n9049), .ZN(n9054) );
  INV_X1 U10363 ( .A(n9048), .ZN(n8944) );
  AND2_X1 U10364 ( .A1(n9109), .A2(n8944), .ZN(n8945) );
  NOR2_X1 U10365 ( .A1(n9054), .A2(n8945), .ZN(n8946) );
  OR2_X1 U10366 ( .A1(n8947), .A2(n8946), .ZN(n8949) );
  INV_X1 U10367 ( .A(n9060), .ZN(n8948) );
  NAND2_X1 U10368 ( .A1(n8949), .A2(n8948), .ZN(n9135) );
  INV_X1 U10369 ( .A(n9135), .ZN(n8950) );
  NAND2_X1 U10370 ( .A1(n9563), .A2(n9240), .ZN(n9104) );
  OAI211_X1 U10371 ( .C1(n9134), .C2(n8951), .A(n8950), .B(n9104), .ZN(n8953)
         );
  INV_X1 U10372 ( .A(n9139), .ZN(n8952) );
  AOI21_X1 U10373 ( .B1(n8954), .B2(n8953), .A(n8952), .ZN(n8955) );
  XNOR2_X1 U10374 ( .A(n8955), .B(n9317), .ZN(n9150) );
  NAND2_X1 U10375 ( .A1(n8956), .A2(n9445), .ZN(n8957) );
  MUX2_X1 U10376 ( .A(n9354), .B(n9481), .S(n9070), .Z(n8958) );
  NOR2_X1 U10377 ( .A1(n8958), .A2(n9318), .ZN(n9041) );
  AOI21_X1 U10378 ( .B1(n9041), .B2(n9481), .A(n9130), .ZN(n8961) );
  INV_X1 U10379 ( .A(n9132), .ZN(n8959) );
  AOI211_X1 U10380 ( .C1(n9041), .C2(n9354), .A(n8959), .B(n9044), .ZN(n8960)
         );
  MUX2_X1 U10381 ( .A(n8961), .B(n8960), .S(n9070), .Z(n9047) );
  NOR2_X1 U10382 ( .A1(n9318), .A2(n8962), .ZN(n9040) );
  NAND2_X1 U10383 ( .A1(n8964), .A2(n8963), .ZN(n8966) );
  MUX2_X1 U10384 ( .A(n8966), .B(n8965), .S(n9070), .Z(n8967) );
  INV_X1 U10385 ( .A(n8967), .ZN(n9021) );
  INV_X1 U10386 ( .A(n8973), .ZN(n9083) );
  NAND2_X1 U10387 ( .A1(n8974), .A2(n9083), .ZN(n8970) );
  NAND3_X1 U10388 ( .A1(n8970), .A2(n8969), .A3(n8968), .ZN(n8971) );
  NAND2_X1 U10389 ( .A1(n8971), .A2(n8972), .ZN(n8978) );
  OAI211_X1 U10390 ( .C1(n8974), .C2(n8973), .A(n8972), .B(n9117), .ZN(n8976)
         );
  NAND2_X1 U10391 ( .A1(n8976), .A2(n8975), .ZN(n8977) );
  INV_X1 U10392 ( .A(n9070), .ZN(n8994) );
  NAND2_X1 U10393 ( .A1(n8986), .A2(n8979), .ZN(n8982) );
  AOI21_X1 U10394 ( .B1(n8982), .B2(n8981), .A(n8980), .ZN(n8992) );
  INV_X1 U10395 ( .A(n8987), .ZN(n8991) );
  NAND2_X1 U10396 ( .A1(n8989), .A2(n8988), .ZN(n8990) );
  NAND2_X1 U10397 ( .A1(n8993), .A2(n9091), .ZN(n9012) );
  NAND2_X1 U10398 ( .A1(n8995), .A2(n8994), .ZN(n9008) );
  NAND2_X1 U10399 ( .A1(n8997), .A2(n8996), .ZN(n8998) );
  NAND2_X1 U10400 ( .A1(n8999), .A2(n8998), .ZN(n9002) );
  NAND3_X1 U10401 ( .A1(n9004), .A2(n9000), .A3(n9070), .ZN(n9001) );
  OAI21_X1 U10402 ( .B1(n9008), .B2(n9002), .A(n9001), .ZN(n9011) );
  AND2_X1 U10403 ( .A1(n9004), .A2(n9003), .ZN(n9009) );
  NAND3_X1 U10404 ( .A1(n9005), .A2(n9004), .A3(n9070), .ZN(n9006) );
  OAI211_X1 U10405 ( .C1(n9009), .C2(n9008), .A(n9007), .B(n9006), .ZN(n9010)
         );
  INV_X1 U10406 ( .A(n9096), .ZN(n9016) );
  MUX2_X1 U10407 ( .A(n9014), .B(n9013), .S(n9070), .Z(n9015) );
  NAND2_X1 U10408 ( .A1(n9016), .A2(n9015), .ZN(n9020) );
  MUX2_X1 U10409 ( .A(n9018), .B(n9017), .S(n9070), .Z(n9019) );
  NAND3_X1 U10410 ( .A1(n9026), .A2(n9025), .A3(n9024), .ZN(n9032) );
  NAND2_X1 U10411 ( .A1(n9028), .A2(n9027), .ZN(n9030) );
  NAND2_X1 U10412 ( .A1(n9030), .A2(n9029), .ZN(n9031) );
  MUX2_X1 U10413 ( .A(n9032), .B(n9031), .S(n9070), .Z(n9039) );
  NAND2_X1 U10414 ( .A1(n9035), .A2(n9034), .ZN(n9038) );
  INV_X1 U10415 ( .A(n9042), .ZN(n9043) );
  MUX2_X1 U10416 ( .A(n9044), .B(n9043), .S(n9070), .Z(n9045) );
  AOI211_X1 U10417 ( .C1(n9047), .C2(n9046), .A(n9045), .B(n9284), .ZN(n9053)
         );
  NAND2_X1 U10418 ( .A1(n9049), .A2(n9048), .ZN(n9051) );
  MUX2_X1 U10419 ( .A(n9051), .B(n9050), .S(n9070), .Z(n9052) );
  NOR2_X1 U10420 ( .A1(n9053), .A2(n9052), .ZN(n9059) );
  OAI21_X1 U10421 ( .B1(n9055), .B2(n9054), .A(n9074), .ZN(n9057) );
  AOI21_X1 U10422 ( .B1(n9057), .B2(n9237), .A(n9056), .ZN(n9065) );
  NAND2_X1 U10423 ( .A1(n9074), .A2(n9109), .ZN(n9058) );
  OAI21_X1 U10424 ( .B1(n9059), .B2(n9058), .A(n9236), .ZN(n9061) );
  AOI21_X1 U10425 ( .B1(n9061), .B2(n9237), .A(n9060), .ZN(n9062) );
  OAI211_X1 U10426 ( .C1(n9065), .C2(n8994), .A(n9138), .B(n9064), .ZN(n9069)
         );
  NAND2_X1 U10427 ( .A1(n9066), .A2(n9070), .ZN(n9068) );
  NAND2_X1 U10428 ( .A1(n9563), .A2(n9219), .ZN(n9067) );
  NAND2_X1 U10429 ( .A1(n9104), .A2(n9067), .ZN(n9136) );
  INV_X1 U10430 ( .A(n9264), .ZN(n9231) );
  INV_X1 U10431 ( .A(n9296), .ZN(n9295) );
  INV_X1 U10432 ( .A(n9318), .ZN(n9101) );
  NAND2_X1 U10433 ( .A1(n9076), .A2(n9075), .ZN(n9080) );
  NOR4_X1 U10434 ( .A1(n9080), .A2(n9079), .A3(n9078), .A4(n9077), .ZN(n9084)
         );
  NAND4_X1 U10435 ( .A1(n9084), .A2(n9083), .A3(n9082), .A4(n9081), .ZN(n9088)
         );
  NOR4_X1 U10436 ( .A1(n9088), .A2(n9087), .A3(n9086), .A4(n7331), .ZN(n9089)
         );
  NAND4_X1 U10437 ( .A1(n9092), .A2(n9091), .A3(n9090), .A4(n9089), .ZN(n9093)
         );
  NOR4_X1 U10438 ( .A1(n9096), .A2(n9095), .A3(n9094), .A4(n9093), .ZN(n9097)
         );
  NAND4_X1 U10439 ( .A1(n4803), .A2(n9098), .A3(n9418), .A4(n9097), .ZN(n9099)
         );
  NOR4_X1 U10440 ( .A1(n9325), .A2(n9366), .A3(n9391), .A4(n9099), .ZN(n9100)
         );
  NAND4_X1 U10441 ( .A1(n9295), .A2(n9101), .A3(n9352), .A4(n9100), .ZN(n9102)
         );
  NOR4_X1 U10442 ( .A1(n9231), .A2(n9284), .A3(n9103), .A4(n9102), .ZN(n9105)
         );
  NAND4_X1 U10443 ( .A1(n9139), .A2(n9237), .A3(n9105), .A4(n9104), .ZN(n9108)
         );
  INV_X1 U10444 ( .A(n9109), .ZN(n9235) );
  OAI211_X1 U10445 ( .C1(n9113), .C2(n9112), .A(n9111), .B(n9110), .ZN(n9116)
         );
  INV_X1 U10446 ( .A(n9114), .ZN(n9115) );
  NAND2_X1 U10447 ( .A1(n9116), .A2(n9115), .ZN(n9118) );
  AOI22_X1 U10448 ( .A1(n9120), .A2(n9119), .B1(n9118), .B2(n9117), .ZN(n9122)
         );
  OAI21_X1 U10449 ( .B1(n9123), .B2(n9122), .A(n9121), .ZN(n9125) );
  AOI21_X1 U10450 ( .B1(n9126), .B2(n9125), .A(n9124), .ZN(n9129) );
  OAI21_X1 U10451 ( .B1(n9129), .B2(n9128), .A(n9127), .ZN(n9131) );
  AOI21_X1 U10452 ( .B1(n9132), .B2(n9131), .A(n9130), .ZN(n9133) );
  NOR3_X1 U10453 ( .A1(n9134), .A2(n9235), .A3(n9133), .ZN(n9137) );
  NOR3_X1 U10454 ( .A1(n9137), .A2(n9136), .A3(n9135), .ZN(n9142) );
  INV_X1 U10455 ( .A(n9138), .ZN(n9141) );
  OAI211_X1 U10456 ( .C1(n9142), .C2(n9141), .A(n9140), .B(n9139), .ZN(n9143)
         );
  NAND2_X1 U10457 ( .A1(n9143), .A2(n9145), .ZN(n9144) );
  MUX2_X1 U10458 ( .A(n9145), .B(n9144), .S(n9317), .Z(n9146) );
  NAND2_X1 U10459 ( .A1(n9151), .A2(n9217), .ZN(n9152) );
  OAI211_X1 U10460 ( .C1(n5778), .C2(n9154), .A(n9152), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9153) );
  OAI21_X1 U10461 ( .B1(n9155), .B2(n9154), .A(n9153), .ZN(P1_U3240) );
  INV_X1 U10462 ( .A(n9156), .ZN(n9257) );
  MUX2_X1 U10463 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9257), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10464 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9157), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10465 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9299), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10466 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9288), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10467 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9338), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10468 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9354), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10469 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9337), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10470 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9388), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10471 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9409), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10472 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9439), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10473 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9410), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10474 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9436), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10475 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9158), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10476 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9159), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10477 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9160), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10478 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9161), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10479 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9162), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10480 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9163), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10481 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9164), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10482 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9165), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10483 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9166), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10484 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9167), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10485 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9168), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10486 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9169), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10487 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9170), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10488 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n7157), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10489 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n6719), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10490 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6974), .S(P1_U4006), .Z(
        P1_U3556) );
  INV_X1 U10491 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9182) );
  XNOR2_X1 U10492 ( .A(n9205), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9749) );
  INV_X1 U10493 ( .A(n9202), .ZN(n9728) );
  INV_X1 U10494 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10202) );
  XNOR2_X1 U10495 ( .A(n9728), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9733) );
  INV_X1 U10496 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9180) );
  NOR2_X1 U10497 ( .A1(n9715), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9171) );
  AOI21_X1 U10498 ( .B1(n9715), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9171), .ZN(
        n9717) );
  INV_X1 U10499 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9177) );
  INV_X1 U10500 ( .A(n9191), .ZN(n9675) );
  INV_X1 U10501 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10011) );
  AOI21_X1 U10502 ( .B1(n6795), .B2(n9173), .A(n9172), .ZN(n9664) );
  MUX2_X1 U10503 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9174), .S(n9189), .Z(n9663) );
  NOR2_X1 U10504 ( .A1(n9664), .A2(n9663), .ZN(n9662) );
  AOI21_X1 U10505 ( .B1(n9174), .B2(n9189), .A(n9662), .ZN(n9679) );
  NOR2_X1 U10506 ( .A1(n9191), .A2(n10011), .ZN(n9175) );
  AOI21_X1 U10507 ( .B1(n9191), .B2(n10011), .A(n9175), .ZN(n9678) );
  NOR2_X1 U10508 ( .A1(n9679), .A2(n9678), .ZN(n9677) );
  AOI21_X1 U10509 ( .B1(n9675), .B2(n10011), .A(n9677), .ZN(n9693) );
  NOR2_X1 U10510 ( .A1(n9690), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9176) );
  AOI21_X1 U10511 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9690), .A(n9176), .ZN(
        n9694) );
  NOR2_X1 U10512 ( .A1(n9693), .A2(n9694), .ZN(n9692) );
  AOI21_X1 U10513 ( .B1(n9690), .B2(n9177), .A(n9692), .ZN(n9178) );
  NAND2_X1 U10514 ( .A1(n9704), .A2(n9178), .ZN(n9179) );
  XNOR2_X1 U10515 ( .A(n9194), .B(n9178), .ZN(n9706) );
  NAND2_X1 U10516 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9706), .ZN(n9705) );
  NAND2_X1 U10517 ( .A1(n9179), .A2(n9705), .ZN(n9718) );
  NAND2_X1 U10518 ( .A1(n9717), .A2(n9718), .ZN(n9716) );
  OAI21_X1 U10519 ( .B1(n9181), .B2(n9180), .A(n9716), .ZN(n9732) );
  NAND2_X1 U10520 ( .A1(n9733), .A2(n9732), .ZN(n9730) );
  OAI21_X1 U10521 ( .B1(n9728), .B2(n10202), .A(n9730), .ZN(n9748) );
  NOR2_X1 U10522 ( .A1(n9749), .A2(n9748), .ZN(n9747) );
  AOI21_X1 U10523 ( .B1(n9182), .B2(n9744), .A(n9747), .ZN(n9183) );
  XOR2_X1 U10524 ( .A(n9183), .B(P1_REG1_REG_19__SCAN_IN), .Z(n9209) );
  INV_X1 U10525 ( .A(n9184), .ZN(n9188) );
  NOR2_X1 U10526 ( .A1(n9185), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9186) );
  AOI21_X1 U10527 ( .B1(n9188), .B2(n9187), .A(n9186), .ZN(n9656) );
  MUX2_X1 U10528 ( .A(n7609), .B(P1_REG2_REG_12__SCAN_IN), .S(n9189), .Z(n9657) );
  MUX2_X1 U10529 ( .A(n9190), .B(P1_REG2_REG_13__SCAN_IN), .S(n9191), .Z(n9668) );
  NOR2_X1 U10530 ( .A1(n9192), .A2(n9690), .ZN(n9193) );
  XNOR2_X1 U10531 ( .A(n9690), .B(n9192), .ZN(n9684) );
  NOR2_X1 U10532 ( .A1(n7801), .A2(n9684), .ZN(n9686) );
  NOR2_X1 U10533 ( .A1(n9193), .A2(n9686), .ZN(n9195) );
  NOR2_X1 U10534 ( .A1(n9195), .A2(n9194), .ZN(n9196) );
  INV_X1 U10535 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9700) );
  NOR2_X1 U10536 ( .A1(n9715), .A2(n9197), .ZN(n9198) );
  AOI21_X1 U10537 ( .B1(n9715), .B2(n9197), .A(n9198), .ZN(n9711) );
  AOI21_X1 U10538 ( .B1(n9715), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9710), .ZN(
        n9722) );
  OR2_X1 U10539 ( .A1(n9202), .A2(n9199), .ZN(n9201) );
  NAND2_X1 U10540 ( .A1(n9202), .A2(n9199), .ZN(n9200) );
  AND2_X1 U10541 ( .A1(n9201), .A2(n9200), .ZN(n9723) );
  NOR2_X1 U10542 ( .A1(n9722), .A2(n9723), .ZN(n9725) );
  AOI21_X1 U10543 ( .B1(n9202), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9725), .ZN(
        n9737) );
  OR2_X1 U10544 ( .A1(n9205), .A2(n9427), .ZN(n9204) );
  NAND2_X1 U10545 ( .A1(n9205), .A2(n9427), .ZN(n9203) );
  AND2_X1 U10546 ( .A1(n9204), .A2(n9203), .ZN(n9738) );
  NOR2_X1 U10547 ( .A1(n9737), .A2(n9738), .ZN(n9740) );
  NAND3_X1 U10548 ( .A1(n9211), .A2(n9207), .A3(n9206), .ZN(n9208) );
  OAI211_X1 U10549 ( .C1(n9209), .C2(n9751), .A(n9208), .B(n9745), .ZN(n9212)
         );
  INV_X1 U10550 ( .A(n9209), .ZN(n9210) );
  OAI21_X1 U10551 ( .B1(n9754), .B2(n9214), .A(n9213), .ZN(n9215) );
  NAND2_X1 U10552 ( .A1(n9217), .A2(P1_B_REG_SCAN_IN), .ZN(n9218) );
  NAND2_X1 U10553 ( .A1(n9438), .A2(n9218), .ZN(n9241) );
  NOR2_X1 U10554 ( .A1(n9241), .A2(n9219), .ZN(n9562) );
  NAND2_X1 U10555 ( .A1(n9562), .A2(n9379), .ZN(n9223) );
  OAI21_X1 U10556 ( .B1(n9379), .B2(n9220), .A(n9223), .ZN(n9221) );
  AOI21_X1 U10557 ( .B1(n9445), .B2(n9321), .A(n9221), .ZN(n9222) );
  OAI21_X1 U10558 ( .B1(n9447), .B2(n9247), .A(n9222), .ZN(P1_U3261) );
  XNOR2_X1 U10559 ( .A(n9563), .B(n9246), .ZN(n9560) );
  OAI21_X1 U10560 ( .B1(n9379), .B2(n9224), .A(n9223), .ZN(n9225) );
  AOI21_X1 U10561 ( .B1(n9563), .B2(n9321), .A(n9225), .ZN(n9226) );
  OAI21_X1 U10562 ( .B1(n9560), .B2(n9247), .A(n9226), .ZN(P1_U3262) );
  NAND2_X1 U10563 ( .A1(n9230), .A2(n9229), .ZN(n9262) );
  AND2_X1 U10564 ( .A1(n9231), .A2(n9262), .ZN(n9232) );
  NAND2_X1 U10565 ( .A1(n9263), .A2(n9232), .ZN(n9267) );
  INV_X1 U10566 ( .A(n9455), .ZN(n9272) );
  NAND2_X1 U10567 ( .A1(n9267), .A2(n9233), .ZN(n9234) );
  XNOR2_X1 U10568 ( .A(n9234), .B(n9237), .ZN(n9448) );
  INV_X1 U10569 ( .A(n9448), .ZN(n9254) );
  INV_X1 U10570 ( .A(n9237), .ZN(n9238) );
  XNOR2_X1 U10571 ( .A(n9239), .B(n9238), .ZN(n9245) );
  OAI22_X1 U10572 ( .A1(n9242), .A2(n9369), .B1(n9241), .B2(n9240), .ZN(n9243)
         );
  INV_X1 U10573 ( .A(n9243), .ZN(n9244) );
  OAI21_X1 U10574 ( .B1(n9245), .B2(n9389), .A(n9244), .ZN(n9451) );
  OAI21_X1 U10575 ( .B1(n9250), .B2(n9268), .A(n9246), .ZN(n9449) );
  NOR2_X1 U10576 ( .A1(n9449), .A2(n9247), .ZN(n9252) );
  AOI22_X1 U10577 ( .A1(n9248), .A2(n9402), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9404), .ZN(n9249) );
  OAI21_X1 U10578 ( .B1(n9250), .B2(n9423), .A(n9249), .ZN(n9251) );
  AOI211_X1 U10579 ( .C1(n9451), .C2(n9379), .A(n9252), .B(n9251), .ZN(n9253)
         );
  OAI21_X1 U10580 ( .B1(n9254), .B2(n9444), .A(n9253), .ZN(P1_U3355) );
  NAND2_X1 U10581 ( .A1(n9257), .A2(n9438), .ZN(n9259) );
  NAND2_X1 U10582 ( .A1(n9282), .A2(n9437), .ZN(n9258) );
  NAND2_X1 U10583 ( .A1(n9259), .A2(n9258), .ZN(n9260) );
  NAND2_X1 U10584 ( .A1(n9263), .A2(n9262), .ZN(n9265) );
  NAND2_X1 U10585 ( .A1(n9265), .A2(n9264), .ZN(n9266) );
  NAND2_X1 U10586 ( .A1(n9454), .A2(n7325), .ZN(n9275) );
  AOI21_X1 U10587 ( .B1(n9455), .B2(n9269), .A(n9268), .ZN(n9456) );
  AOI22_X1 U10588 ( .A1(n9270), .A2(n9402), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9404), .ZN(n9271) );
  OAI21_X1 U10589 ( .B1(n9272), .B2(n9423), .A(n9271), .ZN(n9273) );
  AOI21_X1 U10590 ( .B1(n9456), .B2(n9414), .A(n9273), .ZN(n9274) );
  OAI211_X1 U10591 ( .C1(n9404), .C2(n9458), .A(n9275), .B(n9274), .ZN(
        P1_U3263) );
  XOR2_X1 U10592 ( .A(n9284), .B(n9276), .Z(n9469) );
  INV_X1 U10593 ( .A(n9277), .ZN(n9278) );
  AOI21_X1 U10594 ( .B1(n9465), .B2(n4616), .A(n9278), .ZN(n9466) );
  AOI22_X1 U10595 ( .A1(n9279), .A2(n9402), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9404), .ZN(n9280) );
  OAI21_X1 U10596 ( .B1(n9281), .B2(n9423), .A(n9280), .ZN(n9290) );
  AND2_X1 U10597 ( .A1(n9282), .A2(n9438), .ZN(n9287) );
  AOI211_X1 U10598 ( .C1(n9285), .C2(n9284), .A(n9389), .B(n9283), .ZN(n9286)
         );
  AOI211_X1 U10599 ( .C1(n9437), .C2(n9288), .A(n9287), .B(n9286), .ZN(n9468)
         );
  NOR2_X1 U10600 ( .A1(n9468), .A2(n9404), .ZN(n9289) );
  AOI211_X1 U10601 ( .C1(n9466), .C2(n9414), .A(n9290), .B(n9289), .ZN(n9291)
         );
  OAI21_X1 U10602 ( .B1(n9469), .B2(n9444), .A(n9291), .ZN(P1_U3265) );
  INV_X1 U10603 ( .A(n9292), .ZN(n9293) );
  AOI21_X1 U10604 ( .B1(n9295), .B2(n9294), .A(n9293), .ZN(n9474) );
  OAI21_X1 U10605 ( .B1(n9311), .B2(n9297), .A(n9296), .ZN(n9298) );
  NAND3_X1 U10606 ( .A1(n4428), .A2(n9433), .A3(n9298), .ZN(n9301) );
  AOI22_X1 U10607 ( .A1(n9299), .A2(n9438), .B1(n9437), .B2(n9338), .ZN(n9300)
         );
  NAND2_X1 U10608 ( .A1(n9301), .A2(n9300), .ZN(n9470) );
  AOI211_X1 U10609 ( .C1(n9472), .C2(n9308), .A(n9776), .B(n9302), .ZN(n9471)
         );
  NAND2_X1 U10610 ( .A1(n9471), .A2(n9430), .ZN(n9305) );
  AOI22_X1 U10611 ( .A1(n9303), .A2(n9402), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9404), .ZN(n9304) );
  OAI211_X1 U10612 ( .C1(n4614), .C2(n9423), .A(n9305), .B(n9304), .ZN(n9306)
         );
  AOI21_X1 U10613 ( .B1(n9470), .B2(n9379), .A(n9306), .ZN(n9307) );
  OAI21_X1 U10614 ( .B1(n9474), .B2(n9444), .A(n9307), .ZN(P1_U3266) );
  INV_X1 U10615 ( .A(n9308), .ZN(n9309) );
  AOI211_X1 U10616 ( .C1(n9478), .C2(n9327), .A(n9776), .B(n9309), .ZN(n9477)
         );
  NOR2_X1 U10617 ( .A1(n9310), .A2(n9425), .ZN(n9316) );
  AOI21_X1 U10618 ( .B1(n9318), .B2(n9312), .A(n9311), .ZN(n9313) );
  OAI222_X1 U10619 ( .A1(n9371), .A2(n9315), .B1(n9369), .B2(n9314), .C1(n9389), .C2(n9313), .ZN(n9476) );
  AOI211_X1 U10620 ( .C1(n9477), .C2(n9317), .A(n9316), .B(n9476), .ZN(n9324)
         );
  OR2_X1 U10621 ( .A1(n9319), .A2(n9318), .ZN(n9475) );
  NAND3_X1 U10622 ( .A1(n9475), .A2(n9320), .A3(n7325), .ZN(n9323) );
  AOI22_X1 U10623 ( .A1(n9478), .A2(n9321), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9404), .ZN(n9322) );
  OAI211_X1 U10624 ( .C1(n9404), .C2(n9324), .A(n9323), .B(n9322), .ZN(
        P1_U3267) );
  XNOR2_X1 U10625 ( .A(n9326), .B(n9325), .ZN(n9485) );
  INV_X1 U10626 ( .A(n9345), .ZN(n9329) );
  INV_X1 U10627 ( .A(n9327), .ZN(n9328) );
  AOI21_X1 U10628 ( .B1(n9481), .B2(n9329), .A(n9328), .ZN(n9482) );
  INV_X1 U10629 ( .A(n9330), .ZN(n9331) );
  AOI22_X1 U10630 ( .A1(n9331), .A2(n9402), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9404), .ZN(n9332) );
  OAI21_X1 U10631 ( .B1(n9333), .B2(n9423), .A(n9332), .ZN(n9342) );
  OAI211_X1 U10632 ( .C1(n9336), .C2(n9335), .A(n9334), .B(n9433), .ZN(n9340)
         );
  AOI22_X1 U10633 ( .A1(n9338), .A2(n9438), .B1(n9437), .B2(n9337), .ZN(n9339)
         );
  NOR2_X1 U10634 ( .A1(n9484), .A2(n9404), .ZN(n9341) );
  AOI211_X1 U10635 ( .C1(n9482), .C2(n9414), .A(n9342), .B(n9341), .ZN(n9343)
         );
  OAI21_X1 U10636 ( .B1(n9485), .B2(n9444), .A(n9343), .ZN(P1_U3268) );
  XOR2_X1 U10637 ( .A(n9352), .B(n9344), .Z(n9490) );
  INV_X1 U10638 ( .A(n9372), .ZN(n9346) );
  AOI21_X1 U10639 ( .B1(n9486), .B2(n9346), .A(n9345), .ZN(n9487) );
  INV_X1 U10640 ( .A(n9347), .ZN(n9348) );
  AOI22_X1 U10641 ( .A1(n9348), .A2(n9402), .B1(n9404), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9349) );
  OAI21_X1 U10642 ( .B1(n9350), .B2(n9423), .A(n9349), .ZN(n9358) );
  OAI211_X1 U10643 ( .C1(n9353), .C2(n9352), .A(n9351), .B(n9433), .ZN(n9356)
         );
  AOI22_X1 U10644 ( .A1(n9354), .A2(n9438), .B1(n9437), .B2(n9388), .ZN(n9355)
         );
  NOR2_X1 U10645 ( .A1(n9489), .A2(n9404), .ZN(n9357) );
  AOI211_X1 U10646 ( .C1(n9487), .C2(n9414), .A(n9358), .B(n9357), .ZN(n9359)
         );
  OAI21_X1 U10647 ( .B1(n9490), .B2(n9444), .A(n9359), .ZN(P1_U3269) );
  OAI21_X1 U10648 ( .B1(n4398), .B2(n9366), .A(n9360), .ZN(n9495) );
  INV_X1 U10649 ( .A(n9361), .ZN(n9363) );
  NAND2_X1 U10650 ( .A1(n9363), .A2(n9362), .ZN(n9365) );
  AOI21_X1 U10651 ( .B1(n9366), .B2(n9365), .A(n9364), .ZN(n9367) );
  OAI222_X1 U10652 ( .A1(n9371), .A2(n9370), .B1(n9369), .B2(n9368), .C1(n9389), .C2(n9367), .ZN(n9491) );
  AOI211_X1 U10653 ( .C1(n9493), .C2(n9382), .A(n9776), .B(n9372), .ZN(n9492)
         );
  NAND2_X1 U10654 ( .A1(n9492), .A2(n9430), .ZN(n9376) );
  INV_X1 U10655 ( .A(n9373), .ZN(n9374) );
  AOI22_X1 U10656 ( .A1(n9404), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9374), .B2(
        n9402), .ZN(n9375) );
  OAI211_X1 U10657 ( .C1(n9377), .C2(n9423), .A(n9376), .B(n9375), .ZN(n9378)
         );
  AOI21_X1 U10658 ( .B1(n9491), .B2(n9379), .A(n9378), .ZN(n9380) );
  OAI21_X1 U10659 ( .B1(n9495), .B2(n9444), .A(n9380), .ZN(P1_U3270) );
  XNOR2_X1 U10660 ( .A(n9381), .B(n9391), .ZN(n9500) );
  INV_X1 U10661 ( .A(n9382), .ZN(n9383) );
  AOI21_X1 U10662 ( .B1(n9496), .B2(n9398), .A(n9383), .ZN(n9497) );
  INV_X1 U10663 ( .A(n9384), .ZN(n9385) );
  AOI22_X1 U10664 ( .A1(n9404), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9385), .B2(
        n9402), .ZN(n9386) );
  OAI21_X1 U10665 ( .B1(n9387), .B2(n9423), .A(n9386), .ZN(n9395) );
  AND2_X1 U10666 ( .A1(n9388), .A2(n9438), .ZN(n9393) );
  AOI211_X1 U10667 ( .C1(n9391), .C2(n9390), .A(n9389), .B(n9361), .ZN(n9392)
         );
  AOI211_X1 U10668 ( .C1(n9437), .C2(n9439), .A(n9393), .B(n9392), .ZN(n9499)
         );
  NOR2_X1 U10669 ( .A1(n9499), .A2(n9404), .ZN(n9394) );
  AOI211_X1 U10670 ( .C1(n9497), .C2(n9414), .A(n9395), .B(n9394), .ZN(n9396)
         );
  OAI21_X1 U10671 ( .B1(n9500), .B2(n9444), .A(n9396), .ZN(P1_U3271) );
  XNOR2_X1 U10672 ( .A(n9397), .B(n4803), .ZN(n9506) );
  INV_X1 U10673 ( .A(n9421), .ZN(n9400) );
  INV_X1 U10674 ( .A(n9398), .ZN(n9399) );
  AOI21_X1 U10675 ( .B1(n9501), .B2(n9400), .A(n9399), .ZN(n9503) );
  INV_X1 U10676 ( .A(n9401), .ZN(n9403) );
  AOI22_X1 U10677 ( .A1(n9404), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9403), .B2(
        n9402), .ZN(n9405) );
  OAI21_X1 U10678 ( .B1(n9406), .B2(n9423), .A(n9405), .ZN(n9413) );
  XNOR2_X1 U10679 ( .A(n9407), .B(n9408), .ZN(n9411) );
  AOI222_X1 U10680 ( .A1(n9433), .A2(n9411), .B1(n9410), .B2(n9437), .C1(n9409), .C2(n9438), .ZN(n9505) );
  NOR2_X1 U10681 ( .A1(n9505), .A2(n9404), .ZN(n9412) );
  AOI211_X1 U10682 ( .C1(n9503), .C2(n9414), .A(n9413), .B(n9412), .ZN(n9415)
         );
  OAI21_X1 U10683 ( .B1(n9506), .B2(n9444), .A(n9415), .ZN(P1_U3272) );
  AOI21_X1 U10684 ( .B1(n9418), .B2(n9417), .A(n9416), .ZN(n9419) );
  INV_X1 U10685 ( .A(n9419), .ZN(n9511) );
  INV_X1 U10686 ( .A(n9420), .ZN(n9422) );
  AOI211_X1 U10687 ( .C1(n9509), .C2(n9422), .A(n9776), .B(n9421), .ZN(n9508)
         );
  NOR2_X1 U10688 ( .A1(n9424), .A2(n9423), .ZN(n9429) );
  OAI22_X1 U10689 ( .A1(n9379), .A2(n9427), .B1(n9426), .B2(n9425), .ZN(n9428)
         );
  AOI211_X1 U10690 ( .C1(n9508), .C2(n9430), .A(n9429), .B(n9428), .ZN(n9443)
         );
  AND2_X1 U10691 ( .A1(n9432), .A2(n9431), .ZN(n9434) );
  OAI21_X1 U10692 ( .B1(n9435), .B2(n9434), .A(n9433), .ZN(n9441) );
  AOI22_X1 U10693 ( .A1(n9439), .A2(n9438), .B1(n9437), .B2(n9436), .ZN(n9440)
         );
  NAND2_X1 U10694 ( .A1(n9441), .A2(n9440), .ZN(n9507) );
  NAND2_X1 U10695 ( .A1(n9507), .A2(n9379), .ZN(n9442) );
  OAI211_X1 U10696 ( .C1(n9511), .C2(n9444), .A(n9443), .B(n9442), .ZN(
        P1_U3273) );
  AOI21_X1 U10697 ( .B1(n9445), .B2(n9564), .A(n9562), .ZN(n9446) );
  OAI21_X1 U10698 ( .B1(n9447), .B2(n9776), .A(n9446), .ZN(n9529) );
  MUX2_X1 U10699 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9529), .S(n9528), .Z(
        P1_U3554) );
  NAND2_X1 U10700 ( .A1(n9448), .A2(n9771), .ZN(n9453) );
  NAND2_X1 U10701 ( .A1(n9453), .A2(n9452), .ZN(n9530) );
  MUX2_X1 U10702 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9530), .S(n9786), .Z(
        P1_U3552) );
  NAND2_X1 U10703 ( .A1(n9454), .A2(n9771), .ZN(n9459) );
  AOI22_X1 U10704 ( .A1(n9456), .A2(n9502), .B1(n9564), .B2(n9455), .ZN(n9457)
         );
  NAND3_X1 U10705 ( .A1(n9459), .A2(n9458), .A3(n9457), .ZN(n9531) );
  MUX2_X1 U10706 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9531), .S(n9786), .Z(
        P1_U3551) );
  AOI22_X1 U10707 ( .A1(n9461), .A2(n9502), .B1(n9564), .B2(n9460), .ZN(n9462)
         );
  OAI211_X1 U10708 ( .C1(n9464), .C2(n9526), .A(n9463), .B(n9462), .ZN(n9532)
         );
  MUX2_X1 U10709 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9532), .S(n9786), .Z(
        P1_U3550) );
  AOI22_X1 U10710 ( .A1(n9466), .A2(n9502), .B1(n9564), .B2(n9465), .ZN(n9467)
         );
  OAI211_X1 U10711 ( .C1(n9469), .C2(n9526), .A(n9468), .B(n9467), .ZN(n9533)
         );
  MUX2_X1 U10712 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9533), .S(n9786), .Z(
        P1_U3549) );
  AOI211_X1 U10713 ( .C1(n9564), .C2(n9472), .A(n9471), .B(n9470), .ZN(n9473)
         );
  OAI21_X1 U10714 ( .B1(n9474), .B2(n9526), .A(n9473), .ZN(n9534) );
  MUX2_X1 U10715 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9534), .S(n9786), .Z(
        P1_U3548) );
  NAND3_X1 U10716 ( .A1(n9475), .A2(n9320), .A3(n9771), .ZN(n9480) );
  AOI211_X1 U10717 ( .C1(n9564), .C2(n9478), .A(n9477), .B(n9476), .ZN(n9479)
         );
  NAND2_X1 U10718 ( .A1(n9480), .A2(n9479), .ZN(n9535) );
  MUX2_X1 U10719 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9535), .S(n9786), .Z(
        P1_U3547) );
  AOI22_X1 U10720 ( .A1(n9482), .A2(n9502), .B1(n9564), .B2(n9481), .ZN(n9483)
         );
  OAI211_X1 U10721 ( .C1(n9485), .C2(n9526), .A(n9484), .B(n9483), .ZN(n9536)
         );
  MUX2_X1 U10722 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9536), .S(n9786), .Z(
        P1_U3546) );
  AOI22_X1 U10723 ( .A1(n9487), .A2(n9502), .B1(n9564), .B2(n9486), .ZN(n9488)
         );
  OAI211_X1 U10724 ( .C1(n9490), .C2(n9526), .A(n9489), .B(n9488), .ZN(n9537)
         );
  MUX2_X1 U10725 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9537), .S(n9786), .Z(
        P1_U3545) );
  AOI211_X1 U10726 ( .C1(n9564), .C2(n9493), .A(n9492), .B(n9491), .ZN(n9494)
         );
  OAI21_X1 U10727 ( .B1(n9495), .B2(n9526), .A(n9494), .ZN(n9538) );
  MUX2_X1 U10728 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9538), .S(n9786), .Z(
        P1_U3544) );
  AOI22_X1 U10729 ( .A1(n9497), .A2(n9502), .B1(n9564), .B2(n9496), .ZN(n9498)
         );
  OAI211_X1 U10730 ( .C1(n9500), .C2(n9526), .A(n9499), .B(n9498), .ZN(n9539)
         );
  MUX2_X1 U10731 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9539), .S(n9786), .Z(
        P1_U3543) );
  AOI22_X1 U10732 ( .A1(n9503), .A2(n9502), .B1(n9564), .B2(n9501), .ZN(n9504)
         );
  OAI211_X1 U10733 ( .C1(n9506), .C2(n9526), .A(n9505), .B(n9504), .ZN(n9540)
         );
  MUX2_X1 U10734 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9540), .S(n9786), .Z(
        P1_U3542) );
  AOI211_X1 U10735 ( .C1(n9564), .C2(n9509), .A(n9508), .B(n9507), .ZN(n9510)
         );
  OAI21_X1 U10736 ( .B1(n9511), .B2(n9526), .A(n9510), .ZN(n9541) );
  MUX2_X1 U10737 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9541), .S(n9786), .Z(
        P1_U3541) );
  AOI211_X1 U10738 ( .C1(n9564), .C2(n9514), .A(n9513), .B(n9512), .ZN(n9515)
         );
  OAI21_X1 U10739 ( .B1(n9516), .B2(n9526), .A(n9515), .ZN(n9542) );
  MUX2_X1 U10740 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9542), .S(n9786), .Z(
        P1_U3540) );
  AOI211_X1 U10741 ( .C1(n9564), .C2(n9519), .A(n9518), .B(n9517), .ZN(n9520)
         );
  OAI21_X1 U10742 ( .B1(n9521), .B2(n9526), .A(n9520), .ZN(n9543) );
  MUX2_X1 U10743 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9543), .S(n9528), .Z(
        P1_U3539) );
  AOI211_X1 U10744 ( .C1(n9564), .C2(n9524), .A(n9523), .B(n9522), .ZN(n9525)
         );
  OAI21_X1 U10745 ( .B1(n9527), .B2(n9526), .A(n9525), .ZN(n9544) );
  MUX2_X1 U10746 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9544), .S(n9528), .Z(
        P1_U3537) );
  MUX2_X1 U10747 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9529), .S(n9772), .Z(
        P1_U3522) );
  MUX2_X1 U10748 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9530), .S(n9783), .Z(
        P1_U3520) );
  MUX2_X1 U10749 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9531), .S(n9783), .Z(
        P1_U3519) );
  MUX2_X1 U10750 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9532), .S(n9783), .Z(
        P1_U3518) );
  MUX2_X1 U10751 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9533), .S(n9783), .Z(
        P1_U3517) );
  MUX2_X1 U10752 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9534), .S(n9783), .Z(
        P1_U3516) );
  MUX2_X1 U10753 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9535), .S(n9783), .Z(
        P1_U3515) );
  MUX2_X1 U10754 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9536), .S(n9783), .Z(
        P1_U3514) );
  MUX2_X1 U10755 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9537), .S(n9783), .Z(
        P1_U3513) );
  MUX2_X1 U10756 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9538), .S(n9783), .Z(
        P1_U3512) );
  MUX2_X1 U10757 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9539), .S(n9783), .Z(
        P1_U3511) );
  MUX2_X1 U10758 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9540), .S(n9783), .Z(
        P1_U3510) );
  MUX2_X1 U10759 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9541), .S(n9783), .Z(
        P1_U3508) );
  MUX2_X1 U10760 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9542), .S(n9783), .Z(
        P1_U3505) );
  MUX2_X1 U10761 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9543), .S(n9772), .Z(
        P1_U3502) );
  MUX2_X1 U10762 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9544), .S(n9772), .Z(
        P1_U3496) );
  INV_X1 U10763 ( .A(n9545), .ZN(n9551) );
  NOR4_X1 U10764 ( .A1(n4958), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9546), .A4(
        P1_U3084), .ZN(n9547) );
  AOI21_X1 U10765 ( .B1(n9548), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9547), .ZN(
        n9549) );
  OAI21_X1 U10766 ( .B1(n9551), .B2(n9550), .A(n9549), .ZN(P1_U3322) );
  MUX2_X1 U10767 ( .A(n9552), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U10768 ( .A(n9553), .ZN(n9556) );
  NOR2_X1 U10769 ( .A1(n9554), .A2(n9900), .ZN(n9555) );
  AOI22_X1 U10770 ( .A1(n9914), .A2(n9559), .B1(n5840), .B2(n9919), .ZN(
        P2_U3550) );
  INV_X1 U10771 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9558) );
  AOI22_X1 U10772 ( .A1(n9908), .A2(n9559), .B1(n9558), .B2(n9906), .ZN(
        P2_U3518) );
  NOR2_X1 U10773 ( .A1(n9560), .A2(n9776), .ZN(n9561) );
  INV_X1 U10774 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9565) );
  AOI22_X1 U10775 ( .A1(n9786), .A2(n9584), .B1(n9565), .B2(n9787), .ZN(
        P1_U3553) );
  OAI22_X1 U10776 ( .A1(n9566), .A2(n9776), .B1(n7855), .B2(n9774), .ZN(n9567)
         );
  AOI211_X1 U10777 ( .C1(n9569), .C2(n9771), .A(n9568), .B(n9567), .ZN(n9585)
         );
  INV_X1 U10778 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9570) );
  AOI22_X1 U10779 ( .A1(n9786), .A2(n9585), .B1(n9570), .B2(n9787), .ZN(
        P1_U3538) );
  INV_X1 U10780 ( .A(n9571), .ZN(n9781) );
  INV_X1 U10781 ( .A(n9572), .ZN(n9577) );
  OAI22_X1 U10782 ( .A1(n9574), .A2(n9776), .B1(n9573), .B2(n9774), .ZN(n9576)
         );
  AOI211_X1 U10783 ( .C1(n9781), .C2(n9577), .A(n9576), .B(n9575), .ZN(n9587)
         );
  AOI22_X1 U10784 ( .A1(n9786), .A2(n9587), .B1(n10011), .B2(n9787), .ZN(
        P1_U3536) );
  INV_X1 U10785 ( .A(n9578), .ZN(n9583) );
  OAI22_X1 U10786 ( .A1(n9580), .A2(n9776), .B1(n9579), .B2(n9774), .ZN(n9582)
         );
  AOI211_X1 U10787 ( .C1(n9781), .C2(n9583), .A(n9582), .B(n9581), .ZN(n9589)
         );
  AOI22_X1 U10788 ( .A1(n9786), .A2(n9589), .B1(n6795), .B2(n9787), .ZN(
        P1_U3534) );
  AOI22_X1 U10789 ( .A1(n9772), .A2(n9584), .B1(n6529), .B2(n9782), .ZN(
        P1_U3521) );
  AOI22_X1 U10790 ( .A1(n9772), .A2(n9585), .B1(n5398), .B2(n9782), .ZN(
        P1_U3499) );
  INV_X1 U10791 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9586) );
  AOI22_X1 U10792 ( .A1(n9772), .A2(n9587), .B1(n9586), .B2(n9782), .ZN(
        P1_U3493) );
  INV_X1 U10793 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9588) );
  AOI22_X1 U10794 ( .A1(n9772), .A2(n9589), .B1(n9588), .B2(n9782), .ZN(
        P1_U3487) );
  XNOR2_X1 U10795 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10796 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10797 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9598) );
  NAND2_X1 U10798 ( .A1(n4999), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9591) );
  AOI21_X1 U10799 ( .B1(n9592), .B2(n9591), .A(n9590), .ZN(n9594) );
  AOI22_X1 U10800 ( .A1(n9623), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(n9594), .B2(
        n9593), .ZN(n9597) );
  NAND3_X1 U10801 ( .A1(n9731), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9595), .ZN(
        n9596) );
  OAI211_X1 U10802 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n9598), .A(n9597), .B(
        n9596), .ZN(P1_U3241) );
  OAI21_X1 U10803 ( .B1(n9601), .B2(n9600), .A(n9599), .ZN(n9602) );
  AOI22_X1 U10804 ( .A1(n9603), .A2(n9714), .B1(n9655), .B2(n9602), .ZN(n9611)
         );
  AOI21_X1 U10805 ( .B1(n9606), .B2(n9605), .A(n9604), .ZN(n9608) );
  OAI211_X1 U10806 ( .C1(n9608), .C2(n9751), .A(n9607), .B(n4935), .ZN(n9609)
         );
  INV_X1 U10807 ( .A(n9609), .ZN(n9610) );
  OAI211_X1 U10808 ( .C1(n9754), .C2(n9612), .A(n9611), .B(n9610), .ZN(
        P1_U3245) );
  AOI211_X1 U10809 ( .C1(n9615), .C2(n9614), .A(n9613), .B(n9751), .ZN(n9616)
         );
  AOI211_X1 U10810 ( .C1(n9714), .C2(n9618), .A(n9617), .B(n9616), .ZN(n9625)
         );
  OAI21_X1 U10811 ( .B1(n9621), .B2(n9620), .A(n9619), .ZN(n9622) );
  AOI22_X1 U10812 ( .A1(n9623), .A2(P1_ADDR_REG_5__SCAN_IN), .B1(n9655), .B2(
        n9622), .ZN(n9624) );
  NAND2_X1 U10813 ( .A1(n9625), .A2(n9624), .ZN(P1_U3246) );
  OAI21_X1 U10814 ( .B1(n9628), .B2(n9627), .A(n9626), .ZN(n9634) );
  AOI211_X1 U10815 ( .C1(n9631), .C2(n9630), .A(n9629), .B(n9741), .ZN(n9632)
         );
  AOI211_X1 U10816 ( .C1(n9731), .C2(n9634), .A(n9633), .B(n9632), .ZN(n9639)
         );
  INV_X1 U10817 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9636) );
  OAI22_X1 U10818 ( .A1(n9754), .A2(n9636), .B1(n9635), .B2(n9745), .ZN(n9637)
         );
  INV_X1 U10819 ( .A(n9637), .ZN(n9638) );
  NAND2_X1 U10820 ( .A1(n9639), .A2(n9638), .ZN(P1_U3247) );
  OAI21_X1 U10821 ( .B1(n9642), .B2(n9641), .A(n9640), .ZN(n9647) );
  AOI211_X1 U10822 ( .C1(n9644), .C2(n9648), .A(n9643), .B(n9751), .ZN(n9645)
         );
  AOI211_X1 U10823 ( .C1(n9655), .C2(n9647), .A(n9646), .B(n9645), .ZN(n9653)
         );
  NOR3_X1 U10824 ( .A1(n9751), .A2(n9649), .A3(n9648), .ZN(n9651) );
  OAI21_X1 U10825 ( .B1(n9651), .B2(n9714), .A(n9650), .ZN(n9652) );
  OAI211_X1 U10826 ( .C1(n9754), .C2(n10269), .A(n9653), .B(n9652), .ZN(
        P1_U3249) );
  OAI211_X1 U10827 ( .C1(n9657), .C2(n9656), .A(n9655), .B(n9654), .ZN(n9658)
         );
  INV_X1 U10828 ( .A(n9658), .ZN(n9659) );
  AOI211_X1 U10829 ( .C1(n9714), .C2(n9661), .A(n9660), .B(n9659), .ZN(n9667)
         );
  AOI21_X1 U10830 ( .B1(n9664), .B2(n9663), .A(n9662), .ZN(n9665) );
  OR2_X1 U10831 ( .A1(n9665), .A2(n9751), .ZN(n9666) );
  OAI211_X1 U10832 ( .C1(n9754), .C2(n10038), .A(n9667), .B(n9666), .ZN(
        P1_U3253) );
  INV_X1 U10833 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9683) );
  NAND2_X1 U10834 ( .A1(n9669), .A2(n9668), .ZN(n9670) );
  NAND2_X1 U10835 ( .A1(n9670), .A2(n4458), .ZN(n9671) );
  OR2_X1 U10836 ( .A1(n9741), .A2(n9671), .ZN(n9674) );
  INV_X1 U10837 ( .A(n9672), .ZN(n9673) );
  OAI211_X1 U10838 ( .C1(n9745), .C2(n9675), .A(n9674), .B(n9673), .ZN(n9676)
         );
  INV_X1 U10839 ( .A(n9676), .ZN(n9682) );
  AOI21_X1 U10840 ( .B1(n9679), .B2(n9678), .A(n9677), .ZN(n9680) );
  OR2_X1 U10841 ( .A1(n9680), .A2(n9751), .ZN(n9681) );
  OAI211_X1 U10842 ( .C1(n9683), .C2(n9754), .A(n9682), .B(n9681), .ZN(
        P1_U3254) );
  INV_X1 U10843 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9698) );
  AND2_X1 U10844 ( .A1(n9684), .A2(n7801), .ZN(n9685) );
  OR3_X1 U10845 ( .A1(n9741), .A2(n9686), .A3(n9685), .ZN(n9689) );
  INV_X1 U10846 ( .A(n9687), .ZN(n9688) );
  OAI211_X1 U10847 ( .C1(n9745), .C2(n9690), .A(n9689), .B(n9688), .ZN(n9691)
         );
  INV_X1 U10848 ( .A(n9691), .ZN(n9697) );
  AOI21_X1 U10849 ( .B1(n9694), .B2(n9693), .A(n9692), .ZN(n9695) );
  OR2_X1 U10850 ( .A1(n9751), .A2(n9695), .ZN(n9696) );
  OAI211_X1 U10851 ( .C1(n9698), .C2(n9754), .A(n9697), .B(n9696), .ZN(
        P1_U3255) );
  INV_X1 U10852 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9709) );
  AOI211_X1 U10853 ( .C1(n9701), .C2(n9700), .A(n9699), .B(n9741), .ZN(n9702)
         );
  AOI211_X1 U10854 ( .C1(n9714), .C2(n9704), .A(n9703), .B(n9702), .ZN(n9708)
         );
  OAI211_X1 U10855 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n9706), .A(n9731), .B(
        n9705), .ZN(n9707) );
  OAI211_X1 U10856 ( .C1(n9709), .C2(n9754), .A(n9708), .B(n9707), .ZN(
        P1_U3256) );
  INV_X1 U10857 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9721) );
  AOI211_X1 U10858 ( .C1(n4449), .C2(n9711), .A(n9710), .B(n9741), .ZN(n9712)
         );
  AOI211_X1 U10859 ( .C1(n9715), .C2(n9714), .A(n9713), .B(n9712), .ZN(n9720)
         );
  OAI211_X1 U10860 ( .C1(n9718), .C2(n9717), .A(n9731), .B(n9716), .ZN(n9719)
         );
  OAI211_X1 U10861 ( .C1(n9721), .C2(n9754), .A(n9720), .B(n9719), .ZN(
        P1_U3257) );
  INV_X1 U10862 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9736) );
  AND2_X1 U10863 ( .A1(n9723), .A2(n9722), .ZN(n9724) );
  OR3_X1 U10864 ( .A1(n9741), .A2(n9725), .A3(n9724), .ZN(n9727) );
  OAI211_X1 U10865 ( .C1(n9745), .C2(n9728), .A(n9727), .B(n9726), .ZN(n9729)
         );
  INV_X1 U10866 ( .A(n9729), .ZN(n9735) );
  OAI211_X1 U10867 ( .C1(n9733), .C2(n9732), .A(n9731), .B(n9730), .ZN(n9734)
         );
  OAI211_X1 U10868 ( .C1(n9736), .C2(n9754), .A(n9735), .B(n9734), .ZN(
        P1_U3258) );
  INV_X1 U10869 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10259) );
  AND2_X1 U10870 ( .A1(n9738), .A2(n9737), .ZN(n9739) );
  OAI211_X1 U10871 ( .C1(n9745), .C2(n9744), .A(n9743), .B(n9742), .ZN(n9746)
         );
  INV_X1 U10872 ( .A(n9746), .ZN(n9753) );
  AOI21_X1 U10873 ( .B1(n9749), .B2(n9748), .A(n9747), .ZN(n9750) );
  OR2_X1 U10874 ( .A1(n9751), .A2(n9750), .ZN(n9752) );
  OAI211_X1 U10875 ( .C1(n10259), .C2(n9754), .A(n9753), .B(n9752), .ZN(
        P1_U3259) );
  AND2_X1 U10876 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9757), .ZN(P1_U3292) );
  INV_X1 U10877 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10054) );
  NOR2_X1 U10878 ( .A1(n9758), .A2(n10054), .ZN(P1_U3293) );
  INV_X1 U10879 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10221) );
  NOR2_X1 U10880 ( .A1(n9758), .A2(n10221), .ZN(P1_U3294) );
  AND2_X1 U10881 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9757), .ZN(P1_U3295) );
  AND2_X1 U10882 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9757), .ZN(P1_U3296) );
  AND2_X1 U10883 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9757), .ZN(P1_U3297) );
  AND2_X1 U10884 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9757), .ZN(P1_U3298) );
  AND2_X1 U10885 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9757), .ZN(P1_U3299) );
  INV_X1 U10886 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10163) );
  NOR2_X1 U10887 ( .A1(n9758), .A2(n10163), .ZN(P1_U3300) );
  AND2_X1 U10888 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9757), .ZN(P1_U3301) );
  INV_X1 U10889 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10224) );
  NOR2_X1 U10890 ( .A1(n9758), .A2(n10224), .ZN(P1_U3302) );
  AND2_X1 U10891 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9757), .ZN(P1_U3303) );
  AND2_X1 U10892 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9757), .ZN(P1_U3304) );
  AND2_X1 U10893 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9757), .ZN(P1_U3305) );
  NOR2_X1 U10894 ( .A1(n9758), .A2(n10096), .ZN(P1_U3306) );
  AND2_X1 U10895 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9757), .ZN(P1_U3307) );
  AND2_X1 U10896 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9757), .ZN(P1_U3308) );
  AND2_X1 U10897 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9757), .ZN(P1_U3309) );
  AND2_X1 U10898 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9757), .ZN(P1_U3310) );
  NOR2_X1 U10899 ( .A1(n9758), .A2(n10132), .ZN(P1_U3311) );
  INV_X1 U10900 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n9990) );
  NOR2_X1 U10901 ( .A1(n9758), .A2(n9990), .ZN(P1_U3312) );
  AND2_X1 U10902 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9757), .ZN(P1_U3313) );
  AND2_X1 U10903 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9757), .ZN(P1_U3314) );
  AND2_X1 U10904 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9757), .ZN(P1_U3315) );
  AND2_X1 U10905 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9757), .ZN(P1_U3316) );
  NOR2_X1 U10906 ( .A1(n9758), .A2(n9996), .ZN(P1_U3317) );
  INV_X1 U10907 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10139) );
  NOR2_X1 U10908 ( .A1(n9758), .A2(n10139), .ZN(P1_U3318) );
  AND2_X1 U10909 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9757), .ZN(P1_U3319) );
  AND2_X1 U10910 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9757), .ZN(P1_U3320) );
  NOR2_X1 U10911 ( .A1(n9758), .A2(n10081), .ZN(P1_U3321) );
  OAI22_X1 U10912 ( .A1(n9760), .A2(n9776), .B1(n9759), .B2(n9774), .ZN(n9762)
         );
  AOI211_X1 U10913 ( .C1(n9781), .C2(n9763), .A(n9762), .B(n9761), .ZN(n9784)
         );
  INV_X1 U10914 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9764) );
  AOI22_X1 U10915 ( .A1(n9772), .A2(n9784), .B1(n9764), .B2(n9782), .ZN(
        P1_U3463) );
  INV_X1 U10916 ( .A(n9765), .ZN(n9766) );
  NAND2_X1 U10917 ( .A1(n9767), .A2(n9766), .ZN(n9769) );
  AOI211_X1 U10918 ( .C1(n9771), .C2(n9770), .A(n9769), .B(n9768), .ZN(n9785)
         );
  AOI22_X1 U10919 ( .A1(n9772), .A2(n9785), .B1(n5143), .B2(n9782), .ZN(
        P1_U3472) );
  INV_X1 U10920 ( .A(n9773), .ZN(n9780) );
  OAI22_X1 U10921 ( .A1(n9777), .A2(n9776), .B1(n9775), .B2(n9774), .ZN(n9779)
         );
  AOI211_X1 U10922 ( .C1(n9781), .C2(n9780), .A(n9779), .B(n9778), .ZN(n9789)
         );
  AOI22_X1 U10923 ( .A1(n9783), .A2(n9789), .B1(n5237), .B2(n9782), .ZN(
        P1_U3481) );
  AOI22_X1 U10924 ( .A1(n9786), .A2(n9784), .B1(n6446), .B2(n9787), .ZN(
        P1_U3526) );
  AOI22_X1 U10925 ( .A1(n9786), .A2(n9785), .B1(n6443), .B2(n9787), .ZN(
        P1_U3529) );
  AOI22_X1 U10926 ( .A1(n9786), .A2(n9789), .B1(n9788), .B2(n9787), .ZN(
        P1_U3532) );
  AOI22_X1 U10927 ( .A1(n9791), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9790), .ZN(n9801) );
  OR2_X1 U10928 ( .A1(n9792), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9793) );
  OAI211_X1 U10929 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n9795), .A(n9794), .B(
        n9793), .ZN(n9796) );
  INV_X1 U10930 ( .A(n9796), .ZN(n9799) );
  AOI22_X1 U10931 ( .A1(n9797), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9798) );
  OAI221_X1 U10932 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9801), .C1(n9800), .C2(
        n9799), .A(n9798), .ZN(P2_U3245) );
  INV_X1 U10933 ( .A(n9802), .ZN(n9804) );
  AOI21_X1 U10934 ( .B1(n9805), .B2(n9804), .A(n9803), .ZN(n9816) );
  INV_X1 U10935 ( .A(n9806), .ZN(n9813) );
  AOI22_X1 U10936 ( .A1(n9810), .A2(n9809), .B1(n9808), .B2(n9807), .ZN(n9811)
         );
  OAI21_X1 U10937 ( .B1(n9813), .B2(n9812), .A(n9811), .ZN(n9814) );
  NOR3_X1 U10938 ( .A1(n9816), .A2(n9815), .A3(n9814), .ZN(n9818) );
  AOI22_X1 U10939 ( .A1(n8600), .A2(n6570), .B1(n9818), .B2(n9817), .ZN(
        P2_U3291) );
  INV_X1 U10940 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n9821) );
  NOR2_X1 U10941 ( .A1(n9845), .A2(n9821), .ZN(P2_U3297) );
  INV_X1 U10942 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n9822) );
  NOR2_X1 U10943 ( .A1(n9845), .A2(n9822), .ZN(P2_U3298) );
  NOR2_X1 U10944 ( .A1(n9845), .A2(n9973), .ZN(P2_U3299) );
  INV_X1 U10945 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n9823) );
  NOR2_X1 U10946 ( .A1(n9845), .A2(n9823), .ZN(P2_U3300) );
  INV_X1 U10947 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n9824) );
  NOR2_X1 U10948 ( .A1(n9831), .A2(n9824), .ZN(P2_U3301) );
  INV_X1 U10949 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n9825) );
  NOR2_X1 U10950 ( .A1(n9831), .A2(n9825), .ZN(P2_U3302) );
  INV_X1 U10951 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n9826) );
  NOR2_X1 U10952 ( .A1(n9831), .A2(n9826), .ZN(P2_U3303) );
  INV_X1 U10953 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n9827) );
  NOR2_X1 U10954 ( .A1(n9831), .A2(n9827), .ZN(P2_U3304) );
  INV_X1 U10955 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n9828) );
  NOR2_X1 U10956 ( .A1(n9831), .A2(n9828), .ZN(P2_U3305) );
  NOR2_X1 U10957 ( .A1(n9831), .A2(n9987), .ZN(P2_U3306) );
  NOR2_X1 U10958 ( .A1(n9831), .A2(n9971), .ZN(P2_U3307) );
  INV_X1 U10959 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n10170) );
  NOR2_X1 U10960 ( .A1(n9831), .A2(n10170), .ZN(P2_U3308) );
  INV_X1 U10961 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n9829) );
  NOR2_X1 U10962 ( .A1(n9831), .A2(n9829), .ZN(P2_U3309) );
  INV_X1 U10963 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n9830) );
  NOR2_X1 U10964 ( .A1(n9831), .A2(n9830), .ZN(P2_U3310) );
  INV_X1 U10965 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n10016) );
  NOR2_X1 U10966 ( .A1(n9845), .A2(n10016), .ZN(P2_U3311) );
  INV_X1 U10967 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n9832) );
  NOR2_X1 U10968 ( .A1(n9845), .A2(n9832), .ZN(P2_U3312) );
  INV_X1 U10969 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n9833) );
  NOR2_X1 U10970 ( .A1(n9845), .A2(n9833), .ZN(P2_U3313) );
  INV_X1 U10971 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n9834) );
  NOR2_X1 U10972 ( .A1(n9845), .A2(n9834), .ZN(P2_U3314) );
  INV_X1 U10973 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n9835) );
  NOR2_X1 U10974 ( .A1(n9845), .A2(n9835), .ZN(P2_U3315) );
  INV_X1 U10975 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n10049) );
  NOR2_X1 U10976 ( .A1(n9845), .A2(n10049), .ZN(P2_U3316) );
  INV_X1 U10977 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n9836) );
  NOR2_X1 U10978 ( .A1(n9845), .A2(n9836), .ZN(P2_U3317) );
  INV_X1 U10979 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10028) );
  NOR2_X1 U10980 ( .A1(n9845), .A2(n10028), .ZN(P2_U3318) );
  NOR2_X1 U10981 ( .A1(n9845), .A2(n10105), .ZN(P2_U3319) );
  INV_X1 U10982 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n9837) );
  NOR2_X1 U10983 ( .A1(n9845), .A2(n9837), .ZN(P2_U3320) );
  INV_X1 U10984 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n9838) );
  NOR2_X1 U10985 ( .A1(n9845), .A2(n9838), .ZN(P2_U3321) );
  INV_X1 U10986 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n9839) );
  NOR2_X1 U10987 ( .A1(n9845), .A2(n9839), .ZN(P2_U3322) );
  INV_X1 U10988 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n9840) );
  NOR2_X1 U10989 ( .A1(n9845), .A2(n9840), .ZN(P2_U3323) );
  INV_X1 U10990 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n10085) );
  NOR2_X1 U10991 ( .A1(n9845), .A2(n10085), .ZN(P2_U3324) );
  INV_X1 U10992 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10050) );
  NOR2_X1 U10993 ( .A1(n9845), .A2(n10050), .ZN(P2_U3325) );
  INV_X1 U10994 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n9984) );
  NOR2_X1 U10995 ( .A1(n9845), .A2(n9984), .ZN(P2_U3326) );
  OAI22_X1 U10996 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n9845), .B1(n9844), .B2(
        n9841), .ZN(n9842) );
  INV_X1 U10997 ( .A(n9842), .ZN(P2_U3437) );
  OAI22_X1 U10998 ( .A1(P2_D_REG_1__SCAN_IN), .A2(n9845), .B1(n9844), .B2(
        n9843), .ZN(n9846) );
  INV_X1 U10999 ( .A(n9846), .ZN(P2_U3438) );
  AOI22_X1 U11000 ( .A1(n9848), .A2(n9904), .B1(n4489), .B2(n9847), .ZN(n9849)
         );
  AND2_X1 U11001 ( .A1(n9850), .A2(n9849), .ZN(n9910) );
  INV_X1 U11002 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10025) );
  AOI22_X1 U11003 ( .A1(n9908), .A2(n9910), .B1(n10025), .B2(n9906), .ZN(
        P2_U3451) );
  INV_X1 U11004 ( .A(n9851), .ZN(n9856) );
  OAI22_X1 U11005 ( .A1(n9853), .A2(n9900), .B1(n9852), .B2(n9898), .ZN(n9855)
         );
  AOI211_X1 U11006 ( .C1(n9856), .C2(n9904), .A(n9855), .B(n9854), .ZN(n9911)
         );
  INV_X1 U11007 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9857) );
  AOI22_X1 U11008 ( .A1(n9908), .A2(n9911), .B1(n9857), .B2(n9906), .ZN(
        P2_U3454) );
  INV_X1 U11009 ( .A(n9858), .ZN(n9864) );
  OAI22_X1 U11010 ( .A1(n9860), .A2(n9900), .B1(n9859), .B2(n9898), .ZN(n9863)
         );
  INV_X1 U11011 ( .A(n9861), .ZN(n9862) );
  AOI211_X1 U11012 ( .C1(n9864), .C2(n9904), .A(n9863), .B(n9862), .ZN(n9912)
         );
  INV_X1 U11013 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9865) );
  AOI22_X1 U11014 ( .A1(n9908), .A2(n9912), .B1(n9865), .B2(n9906), .ZN(
        P2_U3457) );
  NAND2_X1 U11015 ( .A1(n9866), .A2(n9904), .ZN(n9872) );
  AOI22_X1 U11016 ( .A1(n9870), .A2(n9869), .B1(n9868), .B2(n9867), .ZN(n9871)
         );
  AND3_X1 U11017 ( .A1(n9873), .A2(n9872), .A3(n9871), .ZN(n9913) );
  INV_X1 U11018 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9874) );
  AOI22_X1 U11019 ( .A1(n9908), .A2(n9913), .B1(n9874), .B2(n9906), .ZN(
        P2_U3463) );
  INV_X1 U11020 ( .A(n9875), .ZN(n9881) );
  OAI22_X1 U11021 ( .A1(n9877), .A2(n9900), .B1(n9876), .B2(n9898), .ZN(n9880)
         );
  INV_X1 U11022 ( .A(n9878), .ZN(n9879) );
  AOI211_X1 U11023 ( .C1(n9881), .C2(n9904), .A(n9880), .B(n9879), .ZN(n9916)
         );
  INV_X1 U11024 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9882) );
  AOI22_X1 U11025 ( .A1(n9908), .A2(n9916), .B1(n9882), .B2(n9906), .ZN(
        P2_U3469) );
  INV_X1 U11026 ( .A(n9883), .ZN(n9897) );
  INV_X1 U11027 ( .A(n9884), .ZN(n9889) );
  OAI22_X1 U11028 ( .A1(n9886), .A2(n9900), .B1(n9885), .B2(n9898), .ZN(n9888)
         );
  AOI211_X1 U11029 ( .C1(n9897), .C2(n9889), .A(n9888), .B(n9887), .ZN(n9917)
         );
  INV_X1 U11030 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9890) );
  AOI22_X1 U11031 ( .A1(n9908), .A2(n9917), .B1(n9890), .B2(n9906), .ZN(
        P2_U3475) );
  INV_X1 U11032 ( .A(n9891), .ZN(n9896) );
  OAI22_X1 U11033 ( .A1(n9893), .A2(n9900), .B1(n9892), .B2(n9898), .ZN(n9895)
         );
  AOI211_X1 U11034 ( .C1(n9897), .C2(n9896), .A(n9895), .B(n9894), .ZN(n9918)
         );
  INV_X1 U11035 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10123) );
  AOI22_X1 U11036 ( .A1(n9908), .A2(n9918), .B1(n10123), .B2(n9906), .ZN(
        P2_U3481) );
  OAI22_X1 U11037 ( .A1(n9901), .A2(n9900), .B1(n9899), .B2(n9898), .ZN(n9903)
         );
  AOI211_X1 U11038 ( .C1(n9905), .C2(n9904), .A(n9903), .B(n9902), .ZN(n9921)
         );
  INV_X1 U11039 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9907) );
  AOI22_X1 U11040 ( .A1(n9908), .A2(n9921), .B1(n9907), .B2(n9906), .ZN(
        P2_U3487) );
  INV_X1 U11041 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9909) );
  AOI22_X1 U11042 ( .A1(n9914), .A2(n9910), .B1(n9909), .B2(n9919), .ZN(
        P2_U3520) );
  AOI22_X1 U11043 ( .A1(n9914), .A2(n9911), .B1(n6556), .B2(n9919), .ZN(
        P2_U3521) );
  INV_X1 U11044 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10126) );
  AOI22_X1 U11045 ( .A1(n9914), .A2(n9912), .B1(n10126), .B2(n9919), .ZN(
        P2_U3522) );
  AOI22_X1 U11046 ( .A1(n9914), .A2(n9913), .B1(n6588), .B2(n9919), .ZN(
        P2_U3524) );
  AOI22_X1 U11047 ( .A1(n9922), .A2(n9916), .B1(n9915), .B2(n9919), .ZN(
        P2_U3526) );
  AOI22_X1 U11048 ( .A1(n9922), .A2(n9917), .B1(n10141), .B2(n9919), .ZN(
        P2_U3528) );
  AOI22_X1 U11049 ( .A1(n9922), .A2(n9918), .B1(n9981), .B2(n9919), .ZN(
        P2_U3530) );
  AOI22_X1 U11050 ( .A1(n9922), .A2(n9921), .B1(n9920), .B2(n9919), .ZN(
        P2_U3532) );
  INV_X1 U11051 ( .A(n9923), .ZN(n9924) );
  NAND2_X1 U11052 ( .A1(n9925), .A2(n9924), .ZN(n9926) );
  XOR2_X1 U11053 ( .A(n9927), .B(n9926), .Z(ADD_1071_U5) );
  XOR2_X1 U11054 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11055 ( .B1(n9930), .B2(n9929), .A(n9928), .ZN(ADD_1071_U56) );
  OAI21_X1 U11056 ( .B1(n9933), .B2(n9932), .A(n9931), .ZN(ADD_1071_U57) );
  OAI21_X1 U11057 ( .B1(n9936), .B2(n9935), .A(n9934), .ZN(ADD_1071_U58) );
  OAI21_X1 U11058 ( .B1(n9939), .B2(n9938), .A(n9937), .ZN(ADD_1071_U59) );
  OAI21_X1 U11059 ( .B1(n9942), .B2(n9941), .A(n9940), .ZN(ADD_1071_U60) );
  OAI21_X1 U11060 ( .B1(n9945), .B2(n9944), .A(n9943), .ZN(ADD_1071_U61) );
  AOI21_X1 U11061 ( .B1(n9948), .B2(n9947), .A(n9946), .ZN(ADD_1071_U62) );
  AOI21_X1 U11062 ( .B1(n9951), .B2(n9950), .A(n9949), .ZN(ADD_1071_U63) );
  AOI222_X1 U11063 ( .A1(n9955), .A2(n9954), .B1(n9953), .B2(
        P2_STATE_REG_SCAN_IN), .C1(P1_DATAO_REG_20__SCAN_IN), .C2(n9952), .ZN(
        n10186) );
  INV_X1 U11064 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9957) );
  AOI22_X1 U11065 ( .A1(n9957), .A2(keyinput125), .B1(keyinput84), .B2(n10264), 
        .ZN(n9956) );
  OAI221_X1 U11066 ( .B1(n9957), .B2(keyinput125), .C1(n10264), .C2(keyinput84), .A(n9956), .ZN(n9967) );
  INV_X1 U11067 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9959) );
  INV_X1 U11068 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n10187) );
  AOI22_X1 U11069 ( .A1(n9959), .A2(keyinput123), .B1(keyinput73), .B2(n10187), 
        .ZN(n9958) );
  OAI221_X1 U11070 ( .B1(n9959), .B2(keyinput123), .C1(n10187), .C2(keyinput73), .A(n9958), .ZN(n9966) );
  AOI22_X1 U11071 ( .A1(n9961), .A2(keyinput55), .B1(n10209), .B2(keyinput98), 
        .ZN(n9960) );
  OAI221_X1 U11072 ( .B1(n9961), .B2(keyinput55), .C1(n10209), .C2(keyinput98), 
        .A(n9960), .ZN(n9965) );
  XOR2_X1 U11073 ( .A(n7431), .B(keyinput116), .Z(n9963) );
  XNOR2_X1 U11074 ( .A(P2_REG2_REG_1__SCAN_IN), .B(keyinput29), .ZN(n9962) );
  NAND2_X1 U11075 ( .A1(n9963), .A2(n9962), .ZN(n9964) );
  NOR4_X1 U11076 ( .A1(n9967), .A2(n9966), .A3(n9965), .A4(n9964), .ZN(n10009)
         );
  AOI22_X1 U11077 ( .A1(n5237), .A2(keyinput82), .B1(n5722), .B2(keyinput41), 
        .ZN(n9968) );
  OAI221_X1 U11078 ( .B1(n5237), .B2(keyinput82), .C1(n5722), .C2(keyinput41), 
        .A(n9968), .ZN(n9979) );
  AOI22_X1 U11079 ( .A1(n9971), .A2(keyinput1), .B1(n9970), .B2(keyinput63), 
        .ZN(n9969) );
  OAI221_X1 U11080 ( .B1(n9971), .B2(keyinput1), .C1(n9970), .C2(keyinput63), 
        .A(n9969), .ZN(n9978) );
  INV_X1 U11081 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9974) );
  AOI22_X1 U11082 ( .A1(n9974), .A2(keyinput108), .B1(keyinput13), .B2(n9973), 
        .ZN(n9972) );
  OAI221_X1 U11083 ( .B1(n9974), .B2(keyinput108), .C1(n9973), .C2(keyinput13), 
        .A(n9972), .ZN(n9977) );
  AOI22_X1 U11084 ( .A1(n7339), .A2(keyinput81), .B1(n10221), .B2(keyinput126), 
        .ZN(n9975) );
  OAI221_X1 U11085 ( .B1(n7339), .B2(keyinput81), .C1(n10221), .C2(keyinput126), .A(n9975), .ZN(n9976) );
  NOR4_X1 U11086 ( .A1(n9979), .A2(n9978), .A3(n9977), .A4(n9976), .ZN(n10008)
         );
  AOI22_X1 U11087 ( .A1(n9982), .A2(keyinput71), .B1(keyinput118), .B2(n9981), 
        .ZN(n9980) );
  OAI221_X1 U11088 ( .B1(n9982), .B2(keyinput71), .C1(n9981), .C2(keyinput118), 
        .A(n9980), .ZN(n9994) );
  AOI22_X1 U11089 ( .A1(n9984), .A2(keyinput110), .B1(n7609), .B2(keyinput25), 
        .ZN(n9983) );
  OAI221_X1 U11090 ( .B1(n9984), .B2(keyinput110), .C1(n7609), .C2(keyinput25), 
        .A(n9983), .ZN(n9993) );
  AOI22_X1 U11091 ( .A1(n9987), .A2(keyinput3), .B1(n9986), .B2(keyinput87), 
        .ZN(n9985) );
  OAI221_X1 U11092 ( .B1(n9987), .B2(keyinput3), .C1(n9986), .C2(keyinput87), 
        .A(n9985), .ZN(n9992) );
  INV_X1 U11093 ( .A(SI_6_), .ZN(n9989) );
  AOI22_X1 U11094 ( .A1(n9990), .A2(keyinput88), .B1(keyinput127), .B2(n9989), 
        .ZN(n9988) );
  OAI221_X1 U11095 ( .B1(n9990), .B2(keyinput88), .C1(n9989), .C2(keyinput127), 
        .A(n9988), .ZN(n9991) );
  NOR4_X1 U11096 ( .A1(n9994), .A2(n9993), .A3(n9992), .A4(n9991), .ZN(n10007)
         );
  AOI22_X1 U11097 ( .A1(n9996), .A2(keyinput49), .B1(keyinput12), .B2(n5886), 
        .ZN(n9995) );
  OAI221_X1 U11098 ( .B1(n9996), .B2(keyinput49), .C1(n5886), .C2(keyinput12), 
        .A(n9995), .ZN(n10005) );
  AOI22_X1 U11099 ( .A1(P1_U3084), .A2(keyinput114), .B1(keyinput106), .B2(
        n10270), .ZN(n9997) );
  OAI221_X1 U11100 ( .B1(P1_U3084), .B2(keyinput114), .C1(n10270), .C2(
        keyinput106), .A(n9997), .ZN(n10004) );
  AOI22_X1 U11101 ( .A1(n5143), .A2(keyinput72), .B1(n9999), .B2(keyinput62), 
        .ZN(n9998) );
  OAI221_X1 U11102 ( .B1(n5143), .B2(keyinput72), .C1(n9999), .C2(keyinput62), 
        .A(n9998), .ZN(n10003) );
  XNOR2_X1 U11103 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput7), .ZN(n10001) );
  XNOR2_X1 U11104 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput83), .ZN(n10000) );
  NAND2_X1 U11105 ( .A1(n10001), .A2(n10000), .ZN(n10002) );
  NOR4_X1 U11106 ( .A1(n10005), .A2(n10004), .A3(n10003), .A4(n10002), .ZN(
        n10006) );
  NAND4_X1 U11107 ( .A1(n10009), .A2(n10008), .A3(n10007), .A4(n10006), .ZN(
        n10184) );
  AOI22_X1 U11108 ( .A1(n10012), .A2(keyinput78), .B1(keyinput20), .B2(n10011), 
        .ZN(n10010) );
  OAI221_X1 U11109 ( .B1(n10012), .B2(keyinput78), .C1(n10011), .C2(keyinput20), .A(n10010), .ZN(n10023) );
  AOI22_X1 U11110 ( .A1(n10015), .A2(keyinput115), .B1(keyinput22), .B2(n10014), .ZN(n10013) );
  OAI221_X1 U11111 ( .B1(n10015), .B2(keyinput115), .C1(n10014), .C2(
        keyinput22), .A(n10013), .ZN(n10022) );
  XNOR2_X1 U11112 ( .A(n10016), .B(keyinput124), .ZN(n10021) );
  XNOR2_X1 U11113 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput86), .ZN(n10019) );
  XNOR2_X1 U11114 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput2), .ZN(n10018) );
  XNOR2_X1 U11115 ( .A(keyinput102), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n10017)
         );
  NAND3_X1 U11116 ( .A1(n10019), .A2(n10018), .A3(n10017), .ZN(n10020) );
  NOR4_X1 U11117 ( .A1(n10023), .A2(n10022), .A3(n10021), .A4(n10020), .ZN(
        n10064) );
  AOI22_X1 U11118 ( .A1(n5828), .A2(keyinput90), .B1(keyinput111), .B2(n10025), 
        .ZN(n10024) );
  OAI221_X1 U11119 ( .B1(n5828), .B2(keyinput90), .C1(n10025), .C2(keyinput111), .A(n10024), .ZN(n10035) );
  AOI22_X1 U11120 ( .A1(n5166), .A2(keyinput99), .B1(keyinput32), .B2(n6443), 
        .ZN(n10026) );
  OAI221_X1 U11121 ( .B1(n5166), .B2(keyinput99), .C1(n6443), .C2(keyinput32), 
        .A(n10026), .ZN(n10034) );
  INV_X1 U11122 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10029) );
  AOI22_X1 U11123 ( .A1(n10029), .A2(keyinput112), .B1(n10028), .B2(
        keyinput109), .ZN(n10027) );
  OAI221_X1 U11124 ( .B1(n10029), .B2(keyinput112), .C1(n10028), .C2(
        keyinput109), .A(n10027), .ZN(n10033) );
  XNOR2_X1 U11125 ( .A(P2_IR_REG_28__SCAN_IN), .B(keyinput19), .ZN(n10031) );
  XNOR2_X1 U11126 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput85), .ZN(n10030)
         );
  NAND2_X1 U11127 ( .A1(n10031), .A2(n10030), .ZN(n10032) );
  NOR4_X1 U11128 ( .A1(n10035), .A2(n10034), .A3(n10033), .A4(n10032), .ZN(
        n10063) );
  AOI22_X1 U11129 ( .A1(n10193), .A2(keyinput107), .B1(keyinput51), .B2(n6104), 
        .ZN(n10036) );
  OAI221_X1 U11130 ( .B1(n10193), .B2(keyinput107), .C1(n6104), .C2(keyinput51), .A(n10036), .ZN(n10047) );
  AOI22_X1 U11131 ( .A1(n10038), .A2(keyinput38), .B1(n6146), .B2(keyinput121), 
        .ZN(n10037) );
  OAI221_X1 U11132 ( .B1(n10038), .B2(keyinput38), .C1(n6146), .C2(keyinput121), .A(n10037), .ZN(n10046) );
  INV_X1 U11133 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n10040) );
  AOI22_X1 U11134 ( .A1(n9197), .A2(keyinput43), .B1(keyinput56), .B2(n10040), 
        .ZN(n10039) );
  OAI221_X1 U11135 ( .B1(n9197), .B2(keyinput43), .C1(n10040), .C2(keyinput56), 
        .A(n10039), .ZN(n10045) );
  XOR2_X1 U11136 ( .A(n10041), .B(keyinput117), .Z(n10043) );
  XNOR2_X1 U11137 ( .A(SI_1_), .B(keyinput96), .ZN(n10042) );
  NAND2_X1 U11138 ( .A1(n10043), .A2(n10042), .ZN(n10044) );
  NOR4_X1 U11139 ( .A1(n10047), .A2(n10046), .A3(n10045), .A4(n10044), .ZN(
        n10062) );
  AOI22_X1 U11140 ( .A1(n10050), .A2(keyinput80), .B1(keyinput21), .B2(n10049), 
        .ZN(n10048) );
  OAI221_X1 U11141 ( .B1(n10050), .B2(keyinput80), .C1(n10049), .C2(keyinput21), .A(n10048), .ZN(n10060) );
  AOI22_X1 U11142 ( .A1(n10190), .A2(keyinput42), .B1(n10052), .B2(keyinput65), 
        .ZN(n10051) );
  OAI221_X1 U11143 ( .B1(n10190), .B2(keyinput42), .C1(n10052), .C2(keyinput65), .A(n10051), .ZN(n10059) );
  AOI22_X1 U11144 ( .A1(n10055), .A2(keyinput91), .B1(n10054), .B2(keyinput66), 
        .ZN(n10053) );
  OAI221_X1 U11145 ( .B1(n10055), .B2(keyinput91), .C1(n10054), .C2(keyinput66), .A(n10053), .ZN(n10058) );
  INV_X1 U11146 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10220) );
  AOI22_X1 U11147 ( .A1(n5209), .A2(keyinput103), .B1(n10220), .B2(keyinput97), 
        .ZN(n10056) );
  OAI221_X1 U11148 ( .B1(n5209), .B2(keyinput103), .C1(n10220), .C2(keyinput97), .A(n10056), .ZN(n10057) );
  NOR4_X1 U11149 ( .A1(n10060), .A2(n10059), .A3(n10058), .A4(n10057), .ZN(
        n10061) );
  NAND4_X1 U11150 ( .A1(n10064), .A2(n10063), .A3(n10062), .A4(n10061), .ZN(
        n10183) );
  AOI22_X1 U11151 ( .A1(n10066), .A2(keyinput53), .B1(keyinput58), .B2(n10228), 
        .ZN(n10065) );
  OAI221_X1 U11152 ( .B1(n10066), .B2(keyinput53), .C1(n10228), .C2(keyinput58), .A(n10065), .ZN(n10079) );
  AOI22_X1 U11153 ( .A1(n10069), .A2(keyinput60), .B1(keyinput100), .B2(n10068), .ZN(n10067) );
  OAI221_X1 U11154 ( .B1(n10069), .B2(keyinput60), .C1(n10068), .C2(
        keyinput100), .A(n10067), .ZN(n10078) );
  AOI22_X1 U11155 ( .A1(n10072), .A2(keyinput36), .B1(n10071), .B2(keyinput48), 
        .ZN(n10070) );
  OAI221_X1 U11156 ( .B1(n10072), .B2(keyinput36), .C1(n10071), .C2(keyinput48), .A(n10070), .ZN(n10077) );
  AOI22_X1 U11157 ( .A1(n10075), .A2(keyinput119), .B1(n10074), .B2(keyinput6), 
        .ZN(n10073) );
  OAI221_X1 U11158 ( .B1(n10075), .B2(keyinput119), .C1(n10074), .C2(keyinput6), .A(n10073), .ZN(n10076) );
  NOR4_X1 U11159 ( .A1(n10079), .A2(n10078), .A3(n10077), .A4(n10076), .ZN(
        n10121) );
  AOI22_X1 U11160 ( .A1(n10082), .A2(keyinput67), .B1(keyinput37), .B2(n10081), 
        .ZN(n10080) );
  OAI221_X1 U11161 ( .B1(n10082), .B2(keyinput67), .C1(n10081), .C2(keyinput37), .A(n10080), .ZN(n10093) );
  AOI22_X1 U11162 ( .A1(n10188), .A2(keyinput35), .B1(keyinput15), .B2(n6176), 
        .ZN(n10083) );
  OAI221_X1 U11163 ( .B1(n10188), .B2(keyinput35), .C1(n6176), .C2(keyinput15), 
        .A(n10083), .ZN(n10092) );
  AOI22_X1 U11164 ( .A1(n10086), .A2(keyinput39), .B1(keyinput68), .B2(n10085), 
        .ZN(n10084) );
  OAI221_X1 U11165 ( .B1(n10086), .B2(keyinput39), .C1(n10085), .C2(keyinput68), .A(n10084), .ZN(n10091) );
  AOI22_X1 U11166 ( .A1(n10089), .A2(keyinput120), .B1(keyinput45), .B2(n10088), .ZN(n10087) );
  OAI221_X1 U11167 ( .B1(n10089), .B2(keyinput120), .C1(n10088), .C2(
        keyinput45), .A(n10087), .ZN(n10090) );
  NOR4_X1 U11168 ( .A1(n10093), .A2(n10092), .A3(n10091), .A4(n10090), .ZN(
        n10120) );
  AOI22_X1 U11169 ( .A1(n10203), .A2(keyinput89), .B1(keyinput14), .B2(n5169), 
        .ZN(n10094) );
  OAI221_X1 U11170 ( .B1(n10203), .B2(keyinput89), .C1(n5169), .C2(keyinput14), 
        .A(n10094), .ZN(n10103) );
  AOI22_X1 U11171 ( .A1(n10225), .A2(keyinput46), .B1(keyinput33), .B2(n10096), 
        .ZN(n10095) );
  OAI221_X1 U11172 ( .B1(n10225), .B2(keyinput46), .C1(n10096), .C2(keyinput33), .A(n10095), .ZN(n10102) );
  AOI22_X1 U11173 ( .A1(n10269), .A2(keyinput93), .B1(n10230), .B2(keyinput47), 
        .ZN(n10097) );
  OAI221_X1 U11174 ( .B1(n10269), .B2(keyinput93), .C1(n10230), .C2(keyinput47), .A(n10097), .ZN(n10101) );
  XNOR2_X1 U11175 ( .A(P1_REG3_REG_8__SCAN_IN), .B(keyinput61), .ZN(n10099) );
  XNOR2_X1 U11176 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput8), .ZN(n10098) );
  NAND2_X1 U11177 ( .A1(n10099), .A2(n10098), .ZN(n10100) );
  NOR4_X1 U11178 ( .A1(n10103), .A2(n10102), .A3(n10101), .A4(n10100), .ZN(
        n10119) );
  AOI22_X1 U11179 ( .A1(n10106), .A2(keyinput54), .B1(keyinput95), .B2(n10105), 
        .ZN(n10104) );
  OAI221_X1 U11180 ( .B1(n10106), .B2(keyinput54), .C1(n10105), .C2(keyinput95), .A(n10104), .ZN(n10108) );
  XNOR2_X1 U11181 ( .A(n10224), .B(keyinput79), .ZN(n10107) );
  NOR2_X1 U11182 ( .A1(n10108), .A2(n10107), .ZN(n10117) );
  AOI22_X1 U11183 ( .A1(n4960), .A2(keyinput30), .B1(n5870), .B2(keyinput113), 
        .ZN(n10109) );
  OAI221_X1 U11184 ( .B1(n4960), .B2(keyinput30), .C1(n5870), .C2(keyinput113), 
        .A(n10109), .ZN(n10110) );
  INV_X1 U11185 ( .A(n10110), .ZN(n10116) );
  INV_X1 U11186 ( .A(SI_14_), .ZN(n10112) );
  AOI22_X1 U11187 ( .A1(n10223), .A2(keyinput34), .B1(keyinput70), .B2(n10112), 
        .ZN(n10111) );
  OAI221_X1 U11188 ( .B1(n10223), .B2(keyinput34), .C1(n10112), .C2(keyinput70), .A(n10111), .ZN(n10113) );
  INV_X1 U11189 ( .A(n10113), .ZN(n10115) );
  XNOR2_X1 U11190 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput64), .ZN(n10114) );
  AND4_X1 U11191 ( .A1(n10117), .A2(n10116), .A3(n10115), .A4(n10114), .ZN(
        n10118) );
  NAND4_X1 U11192 ( .A1(n10121), .A2(n10120), .A3(n10119), .A4(n10118), .ZN(
        n10182) );
  AOI22_X1 U11193 ( .A1(n10202), .A2(keyinput24), .B1(keyinput27), .B2(n10123), 
        .ZN(n10122) );
  OAI221_X1 U11194 ( .B1(n10202), .B2(keyinput24), .C1(n10123), .C2(keyinput27), .A(n10122), .ZN(n10136) );
  AOI22_X1 U11195 ( .A1(n10126), .A2(keyinput122), .B1(n10125), .B2(
        keyinput104), .ZN(n10124) );
  OAI221_X1 U11196 ( .B1(n10126), .B2(keyinput122), .C1(n10125), .C2(
        keyinput104), .A(n10124), .ZN(n10135) );
  AOI22_X1 U11197 ( .A1(n10129), .A2(keyinput28), .B1(keyinput4), .B2(n10128), 
        .ZN(n10127) );
  OAI221_X1 U11198 ( .B1(n10129), .B2(keyinput28), .C1(n10128), .C2(keyinput4), 
        .A(n10127), .ZN(n10134) );
  AOI22_X1 U11199 ( .A1(n10132), .A2(keyinput59), .B1(keyinput16), .B2(n10131), 
        .ZN(n10130) );
  OAI221_X1 U11200 ( .B1(n10132), .B2(keyinput59), .C1(n10131), .C2(keyinput16), .A(n10130), .ZN(n10133) );
  NOR4_X1 U11201 ( .A1(n10136), .A2(n10135), .A3(n10134), .A4(n10133), .ZN(
        n10180) );
  AOI22_X1 U11202 ( .A1(n10139), .A2(keyinput44), .B1(n10138), .B2(keyinput52), 
        .ZN(n10137) );
  OAI221_X1 U11203 ( .B1(n10139), .B2(keyinput44), .C1(n10138), .C2(keyinput52), .A(n10137), .ZN(n10150) );
  AOI22_X1 U11204 ( .A1(n10141), .A2(keyinput50), .B1(keyinput10), .B2(n6586), 
        .ZN(n10140) );
  OAI221_X1 U11205 ( .B1(n10141), .B2(keyinput50), .C1(n6586), .C2(keyinput10), 
        .A(n10140), .ZN(n10149) );
  AOI22_X1 U11206 ( .A1(n10144), .A2(keyinput69), .B1(keyinput5), .B2(n10143), 
        .ZN(n10142) );
  OAI221_X1 U11207 ( .B1(n10144), .B2(keyinput69), .C1(n10143), .C2(keyinput5), 
        .A(n10142), .ZN(n10148) );
  INV_X1 U11208 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n10146) );
  AOI22_X1 U11209 ( .A1(n10146), .A2(keyinput0), .B1(n6592), .B2(keyinput101), 
        .ZN(n10145) );
  OAI221_X1 U11210 ( .B1(n10146), .B2(keyinput0), .C1(n6592), .C2(keyinput101), 
        .A(n10145), .ZN(n10147) );
  NOR4_X1 U11211 ( .A1(n10150), .A2(n10149), .A3(n10148), .A4(n10147), .ZN(
        n10179) );
  AOI22_X1 U11212 ( .A1(n10222), .A2(keyinput11), .B1(keyinput75), .B2(n10152), 
        .ZN(n10151) );
  OAI221_X1 U11213 ( .B1(n10222), .B2(keyinput11), .C1(n10152), .C2(keyinput75), .A(n10151), .ZN(n10161) );
  AOI22_X1 U11214 ( .A1(n5398), .A2(keyinput40), .B1(keyinput74), .B2(n6187), 
        .ZN(n10153) );
  OAI221_X1 U11215 ( .B1(n5398), .B2(keyinput40), .C1(n6187), .C2(keyinput74), 
        .A(n10153), .ZN(n10160) );
  INV_X1 U11216 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n10204) );
  AOI22_X1 U11217 ( .A1(n10204), .A2(keyinput31), .B1(n5347), .B2(keyinput105), 
        .ZN(n10154) );
  OAI221_X1 U11218 ( .B1(n10204), .B2(keyinput31), .C1(n5347), .C2(keyinput105), .A(n10154), .ZN(n10159) );
  XOR2_X1 U11219 ( .A(n10155), .B(keyinput76), .Z(n10157) );
  XNOR2_X1 U11220 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput23), .ZN(n10156) );
  NAND2_X1 U11221 ( .A1(n10157), .A2(n10156), .ZN(n10158) );
  NOR4_X1 U11222 ( .A1(n10161), .A2(n10160), .A3(n10159), .A4(n10158), .ZN(
        n10178) );
  INV_X1 U11223 ( .A(SI_7_), .ZN(n10164) );
  AOI22_X1 U11224 ( .A1(n10164), .A2(keyinput92), .B1(n10163), .B2(keyinput18), 
        .ZN(n10162) );
  OAI221_X1 U11225 ( .B1(n10164), .B2(keyinput92), .C1(n10163), .C2(keyinput18), .A(n10162), .ZN(n10176) );
  INV_X1 U11226 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10167) );
  AOI22_X1 U11227 ( .A1(n10167), .A2(keyinput17), .B1(keyinput26), .B2(n10166), 
        .ZN(n10165) );
  OAI221_X1 U11228 ( .B1(n10167), .B2(keyinput17), .C1(n10166), .C2(keyinput26), .A(n10165), .ZN(n10175) );
  AOI22_X1 U11229 ( .A1(n10170), .A2(keyinput77), .B1(keyinput9), .B2(n10169), 
        .ZN(n10168) );
  OAI221_X1 U11230 ( .B1(n10170), .B2(keyinput77), .C1(n10169), .C2(keyinput9), 
        .A(n10168), .ZN(n10174) );
  INV_X1 U11231 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n10172) );
  AOI22_X1 U11232 ( .A1(n10172), .A2(keyinput57), .B1(keyinput94), .B2(n6570), 
        .ZN(n10171) );
  OAI221_X1 U11233 ( .B1(n10172), .B2(keyinput57), .C1(n6570), .C2(keyinput94), 
        .A(n10171), .ZN(n10173) );
  NOR4_X1 U11234 ( .A1(n10176), .A2(n10175), .A3(n10174), .A4(n10173), .ZN(
        n10177) );
  NAND4_X1 U11235 ( .A1(n10180), .A2(n10179), .A3(n10178), .A4(n10177), .ZN(
        n10181) );
  NOR4_X1 U11236 ( .A1(n10184), .A2(n10183), .A3(n10182), .A4(n10181), .ZN(
        n10185) );
  XNOR2_X1 U11237 ( .A(n10186), .B(n10185), .ZN(n10250) );
  NAND4_X1 U11238 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(P2_ADDR_REG_17__SCAN_IN), .A3(n10188), .A4(n10187), .ZN(n10189) );
  NOR3_X1 U11239 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n10264), .A3(n10189), .ZN(
        n10199) );
  NAND4_X1 U11240 ( .A1(n10192), .A2(n10191), .A3(P2_ADDR_REG_8__SCAN_IN), 
        .A4(n10190), .ZN(n10197) );
  NOR4_X1 U11241 ( .A1(SI_13_), .A2(SI_9_), .A3(n10194), .A4(n10193), .ZN(
        n10195) );
  NAND3_X1 U11242 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(SI_7_), .A3(n10195), 
        .ZN(n10196) );
  NOR4_X1 U11243 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(SI_14_), .A3(n10197), 
        .A4(n10196), .ZN(n10198) );
  NAND4_X1 U11244 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), .A3(n10199), .A4(n10198), .ZN(n10200) );
  NOR4_X1 U11245 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_REG0_REG_15__SCAN_IN), 
        .A3(n10201), .A4(n10200), .ZN(n10248) );
  NAND4_X1 U11246 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG2_REG_27__SCAN_IN), 
        .A3(P2_REG2_REG_27__SCAN_IN), .A4(SI_29_), .ZN(n10208) );
  NAND4_X1 U11247 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_DATAO_REG_28__SCAN_IN), .A4(P1_REG0_REG_6__SCAN_IN), .ZN(n10207) );
  NAND4_X1 U11248 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(P1_REG2_REG_16__SCAN_IN), 
        .A3(P1_REG2_REG_12__SCAN_IN), .A4(n10202), .ZN(n10206) );
  NAND4_X1 U11249 ( .A1(n10204), .A2(n10203), .A3(P1_REG1_REG_21__SCAN_IN), 
        .A4(P1_REG0_REG_20__SCAN_IN), .ZN(n10205) );
  NOR4_X1 U11250 ( .A1(n10208), .A2(n10207), .A3(n10206), .A4(n10205), .ZN(
        n10247) );
  NAND4_X1 U11251 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_REG2_REG_24__SCAN_IN), .A4(P2_REG3_REG_4__SCAN_IN), .ZN(n10214) );
  NAND4_X1 U11252 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_REG0_REG_28__SCAN_IN), .ZN(n10213) );
  NAND4_X1 U11253 ( .A1(P1_REG0_REG_26__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), 
        .A3(P2_REG2_REG_1__SCAN_IN), .A4(P2_REG0_REG_0__SCAN_IN), .ZN(n10212)
         );
  NAND4_X1 U11254 ( .A1(n10210), .A2(n10209), .A3(P1_DATAO_REG_0__SCAN_IN), 
        .A4(SI_6_), .ZN(n10211) );
  NOR4_X1 U11255 ( .A1(n10214), .A2(n10213), .A3(n10212), .A4(n10211), .ZN(
        n10246) );
  NOR4_X1 U11256 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_DATAO_REG_25__SCAN_IN), 
        .A3(P1_REG3_REG_10__SCAN_IN), .A4(P1_REG3_REG_6__SCAN_IN), .ZN(n10218)
         );
  NOR4_X1 U11257 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .A3(
        P1_DATAO_REG_21__SCAN_IN), .A4(P2_IR_REG_28__SCAN_IN), .ZN(n10217) );
  NOR4_X1 U11258 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG0_REG_19__SCAN_IN), 
        .A3(P2_REG1_REG_22__SCAN_IN), .A4(P2_REG1_REG_23__SCAN_IN), .ZN(n10216) );
  NOR4_X1 U11259 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), 
        .A3(P2_REG3_REG_28__SCAN_IN), .A4(P2_REG0_REG_27__SCAN_IN), .ZN(n10215) );
  NAND4_X1 U11260 ( .A1(n10218), .A2(n10217), .A3(n10216), .A4(n10215), .ZN(
        n10244) );
  NOR4_X1 U11261 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(n10221), .A3(n10220), .A4(
        n10219), .ZN(n10232) );
  NOR4_X1 U11262 ( .A1(n10225), .A2(n10224), .A3(n10223), .A4(n10222), .ZN(
        n10227) );
  NOR4_X1 U11263 ( .A1(P1_STATE_REG_SCAN_IN), .A2(P2_REG3_REG_26__SCAN_IN), 
        .A3(P2_REG2_REG_21__SCAN_IN), .A4(P2_REG0_REG_16__SCAN_IN), .ZN(n10226) );
  NAND4_X1 U11264 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P2_REG3_REG_15__SCAN_IN), 
        .A3(n10227), .A4(n10226), .ZN(n10229) );
  NOR3_X1 U11265 ( .A1(n10230), .A2(n10229), .A3(n10228), .ZN(n10231) );
  NAND2_X1 U11266 ( .A1(n10232), .A2(n10231), .ZN(n10243) );
  NOR4_X1 U11267 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(P1_REG2_REG_7__SCAN_IN), 
        .A3(P1_REG1_REG_6__SCAN_IN), .A4(P1_REG2_REG_2__SCAN_IN), .ZN(n10235)
         );
  NOR4_X1 U11268 ( .A1(P1_REG0_REG_9__SCAN_IN), .A2(P1_REG1_REG_4__SCAN_IN), 
        .A3(P1_REG1_REG_2__SCAN_IN), .A4(P1_REG1_REG_1__SCAN_IN), .ZN(n10234)
         );
  NOR4_X1 U11269 ( .A1(SI_27_), .A2(P1_REG1_REG_13__SCAN_IN), .A3(
        P1_REG2_REG_0__SCAN_IN), .A4(P2_DATAO_REG_30__SCAN_IN), .ZN(n10233) );
  NAND4_X1 U11270 ( .A1(n10236), .A2(n10235), .A3(n10234), .A4(n10233), .ZN(
        n10242) );
  NOR4_X1 U11271 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(P2_REG1_REG_8__SCAN_IN), 
        .A3(P2_REG1_REG_7__SCAN_IN), .A4(P2_REG2_REG_5__SCAN_IN), .ZN(n10240)
         );
  NOR4_X1 U11272 ( .A1(P2_REG0_REG_13__SCAN_IN), .A2(P2_REG0_REG_10__SCAN_IN), 
        .A3(P2_REG1_REG_3__SCAN_IN), .A4(P2_REG1_REG_2__SCAN_IN), .ZN(n10239)
         );
  NOR4_X1 U11273 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_REG0_REG_23__SCAN_IN), 
        .A3(P1_REG1_REG_22__SCAN_IN), .A4(P1_REG0_REG_8__SCAN_IN), .ZN(n10238)
         );
  NOR4_X1 U11274 ( .A1(P1_REG1_REG_25__SCAN_IN), .A2(P1_REG1_REG_23__SCAN_IN), 
        .A3(P2_REG3_REG_6__SCAN_IN), .A4(P2_REG3_REG_3__SCAN_IN), .ZN(n10237)
         );
  NAND4_X1 U11275 ( .A1(n10240), .A2(n10239), .A3(n10238), .A4(n10237), .ZN(
        n10241) );
  NOR4_X1 U11276 ( .A1(n10244), .A2(n10243), .A3(n10242), .A4(n10241), .ZN(
        n10245) );
  NAND4_X1 U11277 ( .A1(n10248), .A2(n10247), .A3(n10246), .A4(n10245), .ZN(
        n10249) );
  XNOR2_X1 U11278 ( .A(n10250), .B(n10249), .ZN(P2_U3338) );
  XOR2_X1 U11279 ( .A(n10251), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U11280 ( .A(n10252), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11281 ( .A1(n10254), .A2(n10253), .ZN(n10255) );
  XOR2_X1 U11282 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10255), .Z(ADD_1071_U51) );
  OAI21_X1 U11283 ( .B1(n10258), .B2(n10257), .A(n10256), .ZN(n10260) );
  XOR2_X1 U11284 ( .A(n10260), .B(n10259), .Z(ADD_1071_U55) );
  OAI21_X1 U11285 ( .B1(n10263), .B2(n10262), .A(n10261), .ZN(n10265) );
  XOR2_X1 U11286 ( .A(n10265), .B(n10264), .Z(ADD_1071_U47) );
  XOR2_X1 U11287 ( .A(n10267), .B(n10266), .Z(ADD_1071_U54) );
  AOI21_X1 U11288 ( .B1(n10270), .B2(n10269), .A(n10268), .ZN(n10272) );
  XOR2_X1 U11289 ( .A(n10272), .B(n10271), .Z(ADD_1071_U48) );
  XOR2_X1 U11290 ( .A(n10274), .B(n10273), .Z(ADD_1071_U53) );
  XNOR2_X1 U11291 ( .A(n10276), .B(n10275), .ZN(ADD_1071_U52) );
  NAND2_X1 U6419 ( .A1(n8220), .A2(n8047), .ZN(n5057) );
  INV_X4 U4912 ( .A(n10279), .ZN(n4378) );
  AND2_X2 U4906 ( .A1(n8220), .A2(n4962), .ZN(n5058) );
  CLKBUF_X1 U4885 ( .A(n7213), .Z(n4379) );
  NAND2_X1 U4902 ( .A1(n5837), .A2(n8749), .ZN(n10279) );
endmodule

