

module b22_C_AntiSAT_k_128_7 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, 
        SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, 
        SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, 
        SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, 
        U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, 
        P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, 
        P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, 
        P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, 
        P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, 
        P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, 
        P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, 
        P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, 
        P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, 
        P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, 
        P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, 
        P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, 
        P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, 
        P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, 
        P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, 
        P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, 
        P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, 
        P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, 
        P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, 
        P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, 
        P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, 
        P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, 
        P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, 
        P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, 
        P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, 
        P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, 
        P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, 
        P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, 
        P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, 
        P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, 
        P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, 
        P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, 
        P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, 
        P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, 
        P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, 
        P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, 
        P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, 
        P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, 
        P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9852, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348;

  INV_X1 U7212 ( .A(n15002), .ZN(n6478) );
  INV_X4 U7213 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X4 U7214 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  OAI22_X1 U7215 ( .A1(n13309), .A2(n13311), .B1(n9525), .B2(n13647), .ZN(
        n13293) );
  AND2_X1 U7216 ( .A1(n12238), .A2(n12237), .ZN(n14134) );
  NAND2_X1 U7217 ( .A1(n7431), .A2(n7429), .ZN(n7979) );
  INV_X1 U7218 ( .A(n9769), .ZN(n9727) );
  CLKBUF_X1 U7219 ( .A(n11944), .Z(n12039) );
  INV_X2 U7220 ( .A(n12331), .ZN(n12028) );
  INV_X1 U7221 ( .A(n6544), .ZN(n9354) );
  CLKBUF_X2 U7222 ( .A(n9134), .Z(n6544) );
  INV_X1 U7223 ( .A(n7643), .ZN(n8065) );
  NAND4_X2 U7224 ( .A1(n9119), .A2(n9118), .A3(n9117), .A4(n9116), .ZN(n9559)
         );
  INV_X2 U7225 ( .A(n7662), .ZN(n12242) );
  AND2_X1 U7226 ( .A1(n9072), .A2(n7494), .ZN(n9073) );
  NAND2_X1 U7227 ( .A1(n8173), .A2(n13018), .ZN(n8569) );
  BUF_X1 U7229 ( .A(P3_IR_REG_0__SCAN_IN), .Z(n10764) );
  INV_X1 U7230 ( .A(n7655), .ZN(n7376) );
  INV_X1 U7231 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7566) );
  CLKBUF_X1 U7232 ( .A(n15003), .Z(n6464) );
  INV_X1 U7233 ( .A(n10781), .ZN(n6465) );
  XNOR2_X1 U7234 ( .A(n8210), .B(P3_IR_REG_1__SCAN_IN), .ZN(n10448) );
  XNOR2_X1 U7235 ( .A(n6466), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8172) );
  NOR2_X1 U7236 ( .A1(n6972), .A2(n13011), .ZN(n6466) );
  XNOR2_X1 U7237 ( .A(n9821), .B(n13283), .ZN(n9809) );
  OR2_X1 U7238 ( .A1(n12704), .A2(n8970), .ZN(n8974) );
  AND2_X1 U7239 ( .A1(n12703), .A2(n12702), .ZN(n12704) );
  NAND2_X1 U7240 ( .A1(n6473), .A2(n9854), .ZN(n9134) );
  CLKBUF_X3 U7241 ( .A(n9134), .Z(n6545) );
  INV_X1 U7242 ( .A(n10091), .ZN(n9353) );
  AND3_X2 U7243 ( .A1(n9043), .A2(n9041), .A3(n9042), .ZN(n9048) );
  INV_X1 U7244 ( .A(n12332), .ZN(n12025) );
  NAND2_X1 U7245 ( .A1(n7979), .A2(SI_24_), .ZN(n7980) );
  INV_X1 U7246 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n7775) );
  OR2_X1 U7247 ( .A1(n15163), .A2(n6671), .ZN(n6956) );
  NAND2_X1 U7248 ( .A1(n6789), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8188) );
  INV_X1 U7249 ( .A(n9534), .ZN(n9749) );
  NAND2_X1 U7250 ( .A1(n10896), .A2(n11552), .ZN(n11116) );
  NOR2_X2 U7251 ( .A1(n13429), .A2(n13590), .ZN(n13401) );
  NAND2_X1 U7252 ( .A1(n13401), .A2(n6557), .ZN(n13358) );
  INV_X1 U7253 ( .A(n10927), .ZN(n11223) );
  NAND2_X1 U7254 ( .A1(n8115), .A2(n12248), .ZN(n14792) );
  XNOR2_X1 U7256 ( .A(n7979), .B(SI_24_), .ZN(n7977) );
  MUX2_X1 U7257 ( .A(n12929), .B(P3_REG2_REG_28__SCAN_IN), .S(n12719), .Z(
        n12709) );
  NAND2_X1 U7258 ( .A1(n9387), .A2(n9386), .ZN(n13567) );
  CLKBUF_X2 U7259 ( .A(n9125), .Z(n9534) );
  INV_X2 U7260 ( .A(n11269), .ZN(n13490) );
  INV_X1 U7261 ( .A(n11116), .ZN(n11269) );
  OR2_X2 U7262 ( .A1(n7218), .A2(n7217), .ZN(n11166) );
  OAI21_X1 U7263 ( .B1(n14219), .B2(n9133), .A(n9758), .ZN(n13281) );
  INV_X1 U7264 ( .A(n14177), .ZN(n14058) );
  INV_X1 U7265 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n10344) );
  NAND2_X1 U7266 ( .A1(n7376), .A2(n7566), .ZN(n7684) );
  AOI211_X1 U7267 ( .C1(n12818), .C2(n12869), .A(n12710), .B(n12709), .ZN(
        n12711) );
  NAND2_X1 U7268 ( .A1(n13114), .A2(n13055), .ZN(n13179) );
  XNOR2_X1 U7269 ( .A(n7580), .B(n7579), .ZN(n14609) );
  XOR2_X1 U7270 ( .A(n12303), .B(n13915), .Z(n6467) );
  NOR2_X2 U7271 ( .A1(n13294), .A2(n13542), .ZN(n13288) );
  INV_X8 U7272 ( .A(n12104), .ZN(n12239) );
  NAND3_X2 U7273 ( .A1(n7277), .A2(n10659), .A3(n10667), .ZN(n14602) );
  NAND2_X2 U7274 ( .A1(n10655), .A2(n10654), .ZN(n7277) );
  NAND2_X2 U7275 ( .A1(n7718), .A2(n7516), .ZN(n7733) );
  INV_X1 U7276 ( .A(n13044), .ZN(n6468) );
  INV_X2 U7277 ( .A(n13044), .ZN(n6469) );
  XNOR2_X2 U7278 ( .A(n13510), .B(n13044), .ZN(n11701) );
  NAND2_X1 U7279 ( .A1(n10064), .A2(n10906), .ZN(n6470) );
  NAND2_X1 U7280 ( .A1(n10064), .A2(n10906), .ZN(n6471) );
  OAI222_X1 U7281 ( .A1(P2_U3088), .A2(n13701), .B1(n13708), .B2(n14221), .C1(
        n13700), .C2(n13705), .ZN(P2_U3300) );
  NAND2_X1 U7282 ( .A1(n9530), .A2(n13701), .ZN(n9142) );
  INV_X2 U7283 ( .A(n6534), .ZN(n7620) );
  OAI21_X2 U7284 ( .B1(n12762), .B2(n7340), .A(n7337), .ZN(n12736) );
  OAI21_X2 U7285 ( .B1(n12775), .B2(n8960), .A(n8959), .ZN(n12762) );
  NAND2_X2 U7286 ( .A1(n13861), .A2(n7639), .ZN(n10150) );
  NAND4_X4 U7287 ( .A1(n7635), .A2(n7634), .A3(n7633), .A4(n7632), .ZN(n13861)
         );
  AND2_X2 U7288 ( .A1(n11141), .A2(n10408), .ZN(n10928) );
  OAI21_X2 U7289 ( .B1(n6509), .B2(n6508), .A(n7168), .ZN(n12320) );
  NAND2_X1 U7290 ( .A1(n9530), .A2(n13701), .ZN(n6472) );
  NAND2_X1 U7291 ( .A1(n9530), .A2(n13701), .ZN(n6473) );
  BUF_X2 U7292 ( .A(n9142), .Z(n10091) );
  INV_X2 U7293 ( .A(n12331), .ZN(n6542) );
  INV_X2 U7294 ( .A(n10664), .ZN(n12331) );
  AND2_X2 U7295 ( .A1(n8133), .A2(n9905), .ZN(n8129) );
  NAND4_X4 U7296 ( .A1(n9048), .A2(n9047), .A3(n7447), .A4(n9046), .ZN(n6839)
         );
  NAND4_X2 U7297 ( .A1(n9155), .A2(n9154), .A3(n9153), .A4(n9152), .ZN(n13205)
         );
  OAI22_X2 U7298 ( .A1(n9585), .A2(n7449), .B1(n9586), .B2(n7448), .ZN(n9592)
         );
  OR2_X1 U7299 ( .A1(n9580), .A2(n9579), .ZN(n9585) );
  XNOR2_X2 U7300 ( .A(n8695), .B(n8694), .ZN(n10964) );
  OR2_X2 U7301 ( .A1(n9162), .A2(n9161), .ZN(n10927) );
  NOR2_X2 U7302 ( .A1(n14286), .A2(n15346), .ZN(n14342) );
  NAND4_X4 U7303 ( .A1(n7647), .A2(n7646), .A3(n7645), .A4(n7644), .ZN(n12090)
         );
  OR2_X2 U7304 ( .A1(n6534), .A2(n10910), .ZN(n7646) );
  OR2_X2 U7305 ( .A1(n6541), .A2(n7641), .ZN(n7645) );
  NOR4_X2 U7306 ( .A1(n8853), .A2(n8854), .A3(n8712), .A4(n8711), .ZN(n8713)
         );
  AND2_X4 U7307 ( .A1(n7591), .A2(n11930), .ZN(n7662) );
  NAND2_X1 U7308 ( .A1(n10896), .A2(n11552), .ZN(n6474) );
  NOR2_X2 U7309 ( .A1(n12580), .A2(n14381), .ZN(n14410) );
  NAND2_X4 U7310 ( .A1(n6578), .A2(n7621), .ZN(n13860) );
  AND3_X1 U7311 ( .A1(n7619), .A2(n7618), .A3(n7617), .ZN(n6578) );
  OAI22_X2 U7312 ( .A1(n9599), .A2(n7451), .B1(n7450), .B2(n9600), .ZN(n9606)
         );
  OR2_X1 U7313 ( .A1(n9594), .A2(n9593), .ZN(n9599) );
  NAND2_X1 U7314 ( .A1(n12416), .A2(n13018), .ZN(n6475) );
  XNOR2_X2 U7315 ( .A(n7545), .B(SI_18_), .ZN(n7919) );
  NAND2_X2 U7316 ( .A1(n6893), .A2(n6892), .ZN(n7545) );
  INV_X2 U7317 ( .A(n11146), .ZN(n10897) );
  OAI21_X2 U7318 ( .B1(n10185), .B2(n10183), .A(n12095), .ZN(n14715) );
  CLKBUF_X1 U7319 ( .A(n8569), .Z(n6476) );
  AND2_X2 U7321 ( .A1(n6963), .A2(n6584), .ZN(n14442) );
  XNOR2_X2 U7323 ( .A(n8124), .B(n8123), .ZN(n11911) );
  XNOR2_X2 U7324 ( .A(n9745), .B(n9744), .ZN(n13683) );
  XNOR2_X2 U7325 ( .A(n8188), .B(n8225), .ZN(n10464) );
  OAI21_X2 U7326 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n14287), .A(n14341), .ZN(
        n15343) );
  XNOR2_X2 U7327 ( .A(n13567), .B(n13186), .ZN(n13357) );
  OAI21_X1 U7328 ( .B1(n6505), .B2(n6504), .A(n8862), .ZN(n6503) );
  OAI21_X1 U7329 ( .B1(n9724), .B2(n6822), .A(n6821), .ZN(n9732) );
  XNOR2_X1 U7330 ( .A(n13038), .B(n6567), .ZN(n13149) );
  NAND2_X1 U7331 ( .A1(n8852), .A2(n8848), .ZN(n12702) );
  NOR2_X1 U7332 ( .A1(n14365), .A2(n14366), .ZN(n14364) );
  AND2_X1 U7333 ( .A1(n8841), .A2(n8840), .ZN(n12726) );
  NAND2_X1 U7334 ( .A1(n14583), .A2(n14585), .ZN(n14589) );
  NAND2_X1 U7335 ( .A1(n8832), .A2(n8830), .ZN(n12754) );
  CLKBUF_X1 U7336 ( .A(n14369), .Z(n6717) );
  NAND2_X1 U7337 ( .A1(n14226), .A2(n7676), .ZN(n14025) );
  NOR2_X1 U7338 ( .A1(n12293), .A2(n7405), .ZN(n7404) );
  NAND2_X1 U7339 ( .A1(n7070), .A2(n7069), .ZN(n14121) );
  NAND2_X1 U7340 ( .A1(n7554), .A2(n7553), .ZN(n7956) );
  NAND2_X1 U7341 ( .A1(n12359), .A2(n7239), .ZN(n11186) );
  NAND2_X1 U7342 ( .A1(n9277), .A2(n9276), .ZN(n14830) );
  INV_X1 U7343 ( .A(n12738), .ZN(n12763) );
  INV_X1 U7344 ( .A(n12110), .ZN(n14749) );
  INV_X2 U7345 ( .A(n10430), .ZN(n8978) );
  NAND2_X2 U7346 ( .A1(n10755), .A2(n12676), .ZN(n10626) );
  NAND2_X2 U7347 ( .A1(n11013), .A2(n10966), .ZN(n10430) );
  NAND2_X2 U7348 ( .A1(n15230), .A2(n8723), .ZN(n15261) );
  CLKBUF_X2 U7349 ( .A(n12104), .Z(n12227) );
  INV_X4 U7350 ( .A(n9819), .ZN(n9761) );
  CLKBUF_X1 U7351 ( .A(n8066), .Z(n6534) );
  INV_X1 U7352 ( .A(n11911), .ZN(n8130) );
  BUF_X2 U7353 ( .A(n7642), .Z(n6540) );
  CLKBUF_X2 U7354 ( .A(n7642), .Z(n6541) );
  NAND2_X1 U7355 ( .A1(n14218), .A2(n11930), .ZN(n7642) );
  NAND2_X2 U7356 ( .A1(n9559), .A2(n10897), .ZN(n10573) );
  INV_X4 U7357 ( .A(n8661), .ZN(n8284) );
  NAND2_X2 U7358 ( .A1(n12328), .A2(n12670), .ZN(n10431) );
  INV_X2 U7359 ( .A(n9798), .ZN(n11552) );
  CLKBUF_X2 U7360 ( .A(n9124), .Z(n9422) );
  BUF_X1 U7361 ( .A(n8179), .Z(n8184) );
  NAND2_X1 U7362 ( .A1(n6718), .A2(n9073), .ZN(n13701) );
  CLKBUF_X1 U7363 ( .A(n10464), .Z(n6709) );
  NOR2_X1 U7364 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n7570) );
  OAI21_X1 U7365 ( .B1(n12229), .B2(n12230), .A(n6644), .ZN(n6508) );
  XNOR2_X1 U7366 ( .A(n8888), .B(n8887), .ZN(n8917) );
  AOI21_X1 U7367 ( .B1(n12229), .B2(n12230), .A(n6510), .ZN(n6509) );
  AND2_X1 U7368 ( .A1(n8859), .A2(n8858), .ZN(n6506) );
  AOI21_X1 U7369 ( .B1(n8076), .B2(n14716), .A(n8075), .ZN(n12060) );
  AND2_X1 U7370 ( .A1(n7169), .A2(n12259), .ZN(n7168) );
  OAI21_X1 U7371 ( .B1(n6481), .B2(n6480), .A(n6479), .ZN(n8857) );
  NAND2_X1 U7372 ( .A1(n13072), .A2(n7228), .ZN(n13126) );
  NAND2_X1 U7373 ( .A1(n6481), .A2(n15237), .ZN(n6479) );
  AOI21_X1 U7374 ( .B1(n13934), .B2(n14716), .A(n13933), .ZN(n14139) );
  NAND2_X1 U7375 ( .A1(n6490), .A2(n7125), .ZN(n12221) );
  OR2_X1 U7376 ( .A1(n13546), .A2(n6750), .ZN(n13643) );
  NAND2_X1 U7377 ( .A1(n6483), .A2(n6482), .ZN(n6481) );
  OAI21_X1 U7378 ( .B1(n13043), .B2(n6629), .A(n13047), .ZN(n7222) );
  AND2_X1 U7379 ( .A1(n8983), .A2(n7369), .ZN(n9029) );
  MUX2_X1 U7380 ( .A(n12871), .B(n12870), .S(n15331), .Z(n12874) );
  NAND2_X1 U7381 ( .A1(n6484), .A2(n8856), .ZN(n6483) );
  AND2_X1 U7382 ( .A1(n9811), .A2(n9773), .ZN(n9832) );
  OR2_X1 U7383 ( .A1(n13282), .A2(n13490), .ZN(n13535) );
  OAI211_X1 U7384 ( .C1(n8850), .C2(n6488), .A(n6486), .B(n6485), .ZN(n6484)
         );
  NAND2_X1 U7385 ( .A1(n12708), .A2(n12707), .ZN(n12929) );
  NAND2_X1 U7386 ( .A1(n6528), .A2(n7133), .ZN(n12212) );
  XNOR2_X1 U7387 ( .A(n8974), .B(n8973), .ZN(n8976) );
  NAND2_X1 U7388 ( .A1(n13149), .A2(n13037), .ZN(n13150) );
  INV_X1 U7389 ( .A(n13547), .ZN(n6752) );
  INV_X1 U7390 ( .A(n13923), .ZN(n14131) );
  NAND2_X1 U7391 ( .A1(n6487), .A2(n6488), .ZN(n6486) );
  INV_X1 U7392 ( .A(n8851), .ZN(n6487) );
  INV_X1 U7393 ( .A(n14134), .ZN(n12299) );
  OR3_X1 U7394 ( .A1(n12705), .A2(n12704), .A3(n15249), .ZN(n12708) );
  NAND2_X1 U7395 ( .A1(n13797), .A2(n12004), .ZN(n13723) );
  NAND2_X1 U7396 ( .A1(n7316), .A2(n7315), .ZN(n7314) );
  OR2_X1 U7397 ( .A1(n14219), .A2(n12236), .ZN(n12238) );
  INV_X1 U7398 ( .A(n12702), .ZN(n12699) );
  OAI21_X1 U7399 ( .B1(n7089), .B2(n12297), .A(n6621), .ZN(n7085) );
  AND2_X1 U7400 ( .A1(n8972), .A2(n8852), .ZN(n6485) );
  NAND2_X1 U7401 ( .A1(n12298), .A2(n8109), .ZN(n7089) );
  NAND2_X1 U7402 ( .A1(n9757), .A2(n9742), .ZN(n9745) );
  NAND2_X1 U7403 ( .A1(n9757), .A2(n9756), .ZN(n14219) );
  OR2_X1 U7404 ( .A1(n9755), .A2(n9754), .ZN(n9757) );
  INV_X1 U7405 ( .A(n12228), .ZN(n6510) );
  OAI21_X1 U7406 ( .B1(n6566), .B2(n7401), .A(n7397), .ZN(n14003) );
  NAND2_X1 U7407 ( .A1(n8844), .A2(n8847), .ZN(n8969) );
  NAND2_X1 U7408 ( .A1(n9421), .A2(n9420), .ZN(n13542) );
  NAND2_X1 U7409 ( .A1(n8635), .A2(n8634), .ZN(n12872) );
  OR2_X1 U7410 ( .A1(n12433), .A2(n12406), .ZN(n8844) );
  XNOR2_X1 U7411 ( .A(n9737), .B(n9736), .ZN(n11928) );
  NAND2_X2 U7412 ( .A1(n9409), .A2(n9408), .ZN(n13548) );
  NAND2_X1 U7413 ( .A1(n6916), .A2(n14588), .ZN(n14365) );
  NAND2_X1 U7414 ( .A1(n8622), .A2(n8621), .ZN(n12433) );
  OAI22_X1 U7415 ( .A1(n13372), .A2(n9385), .B1(n13375), .B2(n13187), .ZN(
        n13356) );
  NAND2_X1 U7416 ( .A1(n6520), .A2(n7153), .ZN(n7151) );
  OR2_X1 U7417 ( .A1(n12880), .A2(n8966), .ZN(n8840) );
  NAND2_X1 U7418 ( .A1(n14495), .A2(n7898), .ZN(n14096) );
  AND2_X1 U7419 ( .A1(n9775), .A2(n9774), .ZN(n13335) );
  NOR2_X1 U7420 ( .A1(n13344), .A2(n7104), .ZN(n7103) );
  NOR2_X1 U7421 ( .A1(n13375), .A2(n6907), .ZN(n6906) );
  NAND2_X1 U7422 ( .A1(n6516), .A2(n8608), .ZN(n12880) );
  XNOR2_X1 U7423 ( .A(n8881), .B(n8880), .ZN(n13695) );
  AOI21_X1 U7424 ( .B1(n7402), .B2(n7399), .A(n7398), .ZN(n7397) );
  OAI21_X1 U7425 ( .B1(n12191), .B2(n12189), .A(n12188), .ZN(n6521) );
  NAND2_X1 U7426 ( .A1(n7402), .A2(n7403), .ZN(n7401) );
  NAND2_X1 U7427 ( .A1(n8619), .A2(n7047), .ZN(n7046) );
  NAND2_X1 U7428 ( .A1(n9075), .A2(n9074), .ZN(n13557) );
  INV_X1 U7429 ( .A(n14027), .ZN(n7402) );
  OR2_X1 U7430 ( .A1(n8617), .A2(n8616), .ZN(n8619) );
  NAND2_X1 U7431 ( .A1(n8595), .A2(n8594), .ZN(n12944) );
  XNOR2_X1 U7432 ( .A(n7606), .B(n7605), .ZN(n11855) );
  INV_X1 U7433 ( .A(n14025), .ZN(n14165) );
  NAND2_X1 U7434 ( .A1(n9082), .A2(n9081), .ZN(n13562) );
  NAND2_X1 U7435 ( .A1(n8583), .A2(n8582), .ZN(n12887) );
  AOI21_X1 U7436 ( .B1(n6859), .B2(n6862), .A(n6856), .ZN(n6855) );
  AOI21_X1 U7437 ( .B1(n7404), .B2(n7406), .A(n6624), .ZN(n7403) );
  AND2_X1 U7438 ( .A1(n7249), .A2(n6860), .ZN(n6859) );
  OAI21_X1 U7439 ( .B1(n6512), .B2(n6511), .A(n7157), .ZN(n7155) );
  AOI21_X1 U7440 ( .B1(n12149), .B2(n12150), .A(n6513), .ZN(n6512) );
  OAI21_X1 U7441 ( .B1(n8592), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n6514), .ZN(
        n8604) );
  NOR2_X1 U7442 ( .A1(n12149), .A2(n12150), .ZN(n6511) );
  XNOR2_X1 U7443 ( .A(n7999), .B(n7998), .ZN(n11909) );
  AND2_X1 U7444 ( .A1(n6702), .A2(n6701), .ZN(n14580) );
  OAI21_X1 U7445 ( .B1(n13473), .B2(n6773), .A(n6617), .ZN(n13446) );
  XNOR2_X1 U7446 ( .A(n6905), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14226) );
  NAND2_X1 U7447 ( .A1(n14517), .A2(n7820), .ZN(n11624) );
  OAI21_X1 U7448 ( .B1(n7473), .B2(n9632), .A(n7474), .ZN(n9646) );
  NAND2_X1 U7449 ( .A1(n6514), .A2(n8581), .ZN(n8592) );
  NAND2_X1 U7450 ( .A1(n6515), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6514) );
  NAND2_X1 U7451 ( .A1(n7958), .A2(n7957), .ZN(n14044) );
  NAND2_X1 U7452 ( .A1(n14514), .A2(n7819), .ZN(n14517) );
  NAND2_X1 U7453 ( .A1(n6526), .A2(n12140), .ZN(n12146) );
  XNOR2_X1 U7454 ( .A(n7601), .B(SI_22_), .ZN(n9092) );
  AOI21_X1 U7455 ( .B1(n11820), .B2(n11819), .A(n7480), .ZN(n12361) );
  NAND2_X1 U7456 ( .A1(n7432), .A2(n7557), .ZN(n7601) );
  AND2_X1 U7457 ( .A1(n7947), .A2(n7946), .ZN(n14177) );
  NAND2_X1 U7458 ( .A1(n9096), .A2(n9095), .ZN(n13590) );
  NAND2_X1 U7459 ( .A1(n6527), .A2(n7121), .ZN(n12141) );
  OR3_X1 U7460 ( .A1(n7462), .A2(n7465), .A3(n6845), .ZN(n6842) );
  NAND2_X1 U7461 ( .A1(n8545), .A2(n8544), .ZN(n12966) );
  NAND2_X1 U7462 ( .A1(n7939), .A2(n7938), .ZN(n14181) );
  NAND2_X1 U7463 ( .A1(n6494), .A2(n8566), .ZN(n8577) );
  NOR2_X1 U7464 ( .A1(n15110), .A2(n12575), .ZN(n15129) );
  NOR2_X1 U7465 ( .A1(n11686), .A2(n7271), .ZN(n7270) );
  NAND2_X1 U7466 ( .A1(n6493), .A2(n6491), .ZN(n6494) );
  NAND2_X1 U7467 ( .A1(n11188), .A2(n11045), .ZN(n11260) );
  NAND2_X1 U7468 ( .A1(n6493), .A2(n8556), .ZN(n8565) );
  NAND2_X2 U7469 ( .A1(n9302), .A2(n9301), .ZN(n13672) );
  NAND2_X1 U7470 ( .A1(n9332), .A2(n9331), .ZN(n12073) );
  NAND2_X1 U7471 ( .A1(n8555), .A2(n8554), .ZN(n6493) );
  NAND2_X2 U7472 ( .A1(n9289), .A2(n9288), .ZN(n13510) );
  OAI21_X1 U7473 ( .B1(n7933), .B2(n7932), .A(n7550), .ZN(n7552) );
  AND2_X1 U7474 ( .A1(n11198), .A2(n7767), .ZN(n14656) );
  NAND2_X1 U7475 ( .A1(n7854), .A2(n7853), .ZN(n14545) );
  NAND2_X1 U7476 ( .A1(n11186), .A2(n11037), .ZN(n11043) );
  NAND2_X1 U7477 ( .A1(n9316), .A2(n9315), .ZN(n13477) );
  OAI21_X1 U7478 ( .B1(n7919), .B2(n7446), .A(n7546), .ZN(n7933) );
  OR2_X1 U7479 ( .A1(n8530), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8542) );
  INV_X1 U7480 ( .A(n12148), .ZN(n6513) );
  NAND2_X1 U7481 ( .A1(n8541), .A2(n6518), .ZN(n8530) );
  NAND2_X1 U7482 ( .A1(n6522), .A2(n7129), .ZN(n12121) );
  OR2_X1 U7483 ( .A1(n6519), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6518) );
  NAND2_X2 U7484 ( .A1(n6710), .A2(n9249), .ZN(n13526) );
  NAND2_X1 U7485 ( .A1(n7811), .A2(n7810), .ZN(n14521) );
  NAND2_X1 U7486 ( .A1(n7835), .A2(n7443), .ZN(n7439) );
  AND4_X1 U7487 ( .A1(n8601), .A2(n8600), .A3(n8599), .A4(n8598), .ZN(n12393)
         );
  NAND2_X1 U7488 ( .A1(n9265), .A2(n9264), .ZN(n11741) );
  NAND2_X1 U7489 ( .A1(n7825), .A2(n7824), .ZN(n12147) );
  NAND2_X1 U7490 ( .A1(n7795), .A2(n7794), .ZN(n14478) );
  NAND2_X1 U7491 ( .A1(n6889), .A2(n7532), .ZN(n7835) );
  NAND2_X1 U7492 ( .A1(n9221), .A2(n9220), .ZN(n11363) );
  NAND2_X1 U7493 ( .A1(n6687), .A2(n6651), .ZN(n12572) );
  NAND2_X1 U7494 ( .A1(n7757), .A2(n7756), .ZN(n12127) );
  OAI22_X1 U7495 ( .A1(n12112), .A2(n7117), .B1(n12113), .B2(n7118), .ZN(
        n12115) );
  AND2_X1 U7496 ( .A1(n10675), .A2(n10674), .ZN(n10867) );
  NAND2_X1 U7497 ( .A1(n7771), .A2(n7525), .ZN(n7789) );
  AND2_X1 U7498 ( .A1(n6497), .A2(n6496), .ZN(n6495) );
  NAND2_X1 U7499 ( .A1(n10637), .A2(n7476), .ZN(n10710) );
  NAND2_X2 U7500 ( .A1(n13519), .A2(n10403), .ZN(n13461) );
  INV_X1 U7501 ( .A(n7021), .ZN(n7020) );
  NAND2_X1 U7502 ( .A1(n7021), .A2(n8446), .ZN(n6496) );
  OR2_X1 U7503 ( .A1(n8406), .A2(n10423), .ZN(n8424) );
  OR2_X1 U7504 ( .A1(n8406), .A2(n6498), .ZN(n6497) );
  AND2_X1 U7505 ( .A1(n10709), .A2(n10633), .ZN(n10637) );
  NAND2_X1 U7506 ( .A1(n9181), .A2(n9180), .ZN(n10959) );
  NAND2_X2 U7507 ( .A1(n8901), .A2(n14719), .ZN(n14721) );
  NAND2_X1 U7508 ( .A1(n15335), .A2(n14293), .ZN(n14294) );
  AND2_X2 U7509 ( .A1(n13521), .A2(n9476), .ZN(n13517) );
  INV_X1 U7510 ( .A(n8978), .ZN(n6488) );
  INV_X1 U7511 ( .A(n10620), .ZN(n6480) );
  NAND2_X1 U7512 ( .A1(n8389), .A2(n8388), .ZN(n8402) );
  NAND2_X1 U7513 ( .A1(n8731), .A2(n8730), .ZN(n11018) );
  AND2_X2 U7515 ( .A1(n10063), .A2(n14792), .ZN(n11944) );
  NAND4_X1 U7516 ( .A1(n8237), .A2(n8236), .A3(n8235), .A4(n8234), .ZN(n15217)
         );
  OR2_X1 U7517 ( .A1(n11016), .A2(n15224), .ZN(n8740) );
  NAND2_X1 U7518 ( .A1(n8353), .A2(n8352), .ZN(n8356) );
  INV_X1 U7519 ( .A(n10627), .ZN(n10755) );
  NAND2_X1 U7520 ( .A1(n15332), .A2(n14290), .ZN(n14292) );
  NAND2_X1 U7521 ( .A1(n6888), .A2(n7507), .ZN(n7671) );
  NAND4_X1 U7522 ( .A1(n8197), .A2(n8196), .A3(n8195), .A4(n8194), .ZN(n15257)
         );
  INV_X2 U7523 ( .A(n8345), .ZN(n8674) );
  AND3_X1 U7524 ( .A1(n8213), .A2(n8212), .A3(n8211), .ZN(n15254) );
  CLKBUF_X2 U7525 ( .A(n9611), .Z(n9819) );
  AND3_X1 U7526 ( .A1(n8176), .A2(n8177), .A3(n8175), .ZN(n6986) );
  OR2_X1 U7527 ( .A1(n8483), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8501) );
  CLKBUF_X3 U7528 ( .A(n8066), .Z(n6535) );
  NAND2_X1 U7529 ( .A1(n7651), .A2(n7506), .ZN(n6888) );
  NAND2_X2 U7530 ( .A1(n10406), .A2(n10405), .ZN(n10932) );
  CLKBUF_X1 U7531 ( .A(n7643), .Z(n12241) );
  INV_X1 U7532 ( .A(n6477), .ZN(n8636) );
  OAI21_X1 U7533 ( .B1(n8696), .B2(P3_IR_REG_20__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8695) );
  NAND2_X2 U7534 ( .A1(n7276), .A2(n10906), .ZN(n12332) );
  XNOR2_X1 U7535 ( .A(n8126), .B(P1_IR_REG_24__SCAN_IN), .ZN(n8133) );
  NAND2_X1 U7536 ( .A1(n8294), .A2(n8293), .ZN(n8297) );
  NAND4_X1 U7537 ( .A1(n9141), .A2(n9140), .A3(n9139), .A4(n9138), .ZN(n13206)
         );
  NAND2_X2 U7538 ( .A1(n12416), .A2(n13018), .ZN(n8679) );
  NAND2_X1 U7539 ( .A1(n7591), .A2(n7594), .ZN(n8066) );
  INV_X1 U7540 ( .A(n7589), .ZN(n14218) );
  XNOR2_X1 U7541 ( .A(n8865), .B(n8864), .ZN(n8985) );
  NAND4_X1 U7542 ( .A1(n9108), .A2(n9107), .A3(n9106), .A4(n9105), .ZN(n9552)
         );
  INV_X1 U7543 ( .A(n13915), .ZN(n14511) );
  INV_X1 U7544 ( .A(n10906), .ZN(n12086) );
  INV_X1 U7545 ( .A(n8171), .ZN(n13018) );
  NAND2_X1 U7546 ( .A1(n8870), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8865) );
  XNOR2_X1 U7547 ( .A(n7585), .B(P1_IR_REG_30__SCAN_IN), .ZN(n7589) );
  NAND2_X1 U7548 ( .A1(n6517), .A2(n8278), .ZN(n8292) );
  NOR2_X1 U7549 ( .A1(n8495), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n6681) );
  MUX2_X1 U7550 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8183), .S(
        P3_IR_REG_27__SCAN_IN), .Z(n8185) );
  NOR2_X1 U7551 ( .A1(n8395), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8416) );
  NAND2_X1 U7552 ( .A1(n12255), .A2(n8114), .ZN(n10906) );
  INV_X1 U7553 ( .A(n11930), .ZN(n7594) );
  INV_X1 U7554 ( .A(n9136), .ZN(n9753) );
  INV_X1 U7555 ( .A(n8114), .ZN(n12248) );
  NAND2_X1 U7556 ( .A1(n14212), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7585) );
  AND2_X1 U7557 ( .A1(n9448), .A2(n9447), .ZN(n9449) );
  CLKBUF_X1 U7558 ( .A(n8450), .Z(n8717) );
  OR2_X1 U7559 ( .A1(n9450), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n9453) );
  XNOR2_X1 U7560 ( .A(n7588), .B(n7587), .ZN(n11930) );
  NAND2_X1 U7561 ( .A1(n7578), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7580) );
  NAND2_X1 U7562 ( .A1(n7511), .A2(SI_5_), .ZN(n7513) );
  NAND2_X1 U7563 ( .A1(n8430), .A2(n6678), .ZN(n8179) );
  OR3_X1 U7564 ( .A1(n9446), .A2(n9454), .A3(n9431), .ZN(n9448) );
  AND2_X1 U7565 ( .A1(n7906), .A2(n7905), .ZN(n7923) );
  XNOR2_X1 U7566 ( .A(n8245), .B(n8244), .ZN(n12626) );
  NAND2_X2 U7567 ( .A1(n9874), .A2(P1_U3086), .ZN(n14216) );
  NOR2_X1 U7568 ( .A1(n9339), .A2(n7244), .ZN(n9446) );
  NAND2_X1 U7569 ( .A1(n6500), .A2(n8223), .ZN(n8240) );
  NAND2_X1 U7570 ( .A1(n13684), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9056) );
  NAND2_X1 U7571 ( .A1(n9072), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9070) );
  INV_X2 U7572 ( .A(n9854), .ZN(n9874) );
  INV_X2 U7573 ( .A(n9854), .ZN(n6533) );
  NAND2_X1 U7574 ( .A1(n6788), .A2(n6600), .ZN(n14853) );
  XNOR2_X1 U7575 ( .A(n8227), .B(n8226), .ZN(n10490) );
  NAND2_X1 U7576 ( .A1(n8222), .A2(n6501), .ZN(n6500) );
  INV_X2 U7577 ( .A(n7503), .ZN(n9854) );
  NAND2_X1 U7578 ( .A1(n6502), .A2(n8186), .ZN(n8222) );
  NOR2_X1 U7579 ( .A1(n8564), .A2(n6492), .ZN(n6491) );
  AND2_X1 U7580 ( .A1(n9434), .A2(n6591), .ZN(n6547) );
  AND2_X1 U7581 ( .A1(n6645), .A2(n7575), .ZN(n7407) );
  INV_X1 U7582 ( .A(n8556), .ZN(n6492) );
  NAND2_X1 U7583 ( .A1(n8223), .A2(n8187), .ZN(n8221) );
  AND3_X1 U7584 ( .A1(n7177), .A2(n7176), .A3(n7175), .ZN(n9434) );
  AND2_X2 U7585 ( .A1(n6969), .A2(n6970), .ZN(n10435) );
  AND4_X1 U7586 ( .A1(n9052), .A2(n9051), .A3(n9050), .A4(n9049), .ZN(n9053)
         );
  AND2_X1 U7587 ( .A1(n7571), .A2(n7570), .ZN(n7378) );
  AND2_X1 U7589 ( .A1(n9120), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8208) );
  NOR2_X1 U7590 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n7176) );
  INV_X1 U7591 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8341) );
  INV_X1 U7592 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n14332) );
  INV_X1 U7593 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n6970) );
  INV_X1 U7594 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n6969) );
  INV_X1 U7595 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8302) );
  INV_X1 U7596 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9120) );
  NOR2_X1 U7597 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n8155) );
  NOR2_X1 U7598 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n7177) );
  INV_X1 U7599 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8131) );
  INV_X4 U7600 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U7601 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n8159) );
  NOR2_X1 U7602 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n8158) );
  INV_X1 U7603 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7447) );
  NOR2_X1 U7604 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n7175) );
  INV_X1 U7605 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9437) );
  NOR2_X1 U7606 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n7571) );
  INV_X1 U7607 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n7567) );
  NAND2_X1 U7608 ( .A1(n8854), .A2(n8855), .ZN(n6482) );
  NAND2_X1 U7609 ( .A1(n8689), .A2(n8688), .ZN(n8854) );
  NAND2_X1 U7610 ( .A1(n6489), .A2(n12220), .ZN(n12226) );
  NAND2_X1 U7611 ( .A1(n12221), .A2(n12222), .ZN(n6489) );
  NAND3_X1 U7612 ( .A1(n12217), .A2(n12216), .A3(n7123), .ZN(n6490) );
  NAND2_X1 U7613 ( .A1(n8577), .A2(n8576), .ZN(n8579) );
  NAND3_X1 U7614 ( .A1(n6497), .A2(n6496), .A3(n8460), .ZN(n8463) );
  NAND3_X1 U7615 ( .A1(n8426), .A2(n8446), .A3(P1_DATAO_REG_13__SCAN_IN), .ZN(
        n6498) );
  INV_X1 U7616 ( .A(n8221), .ZN(n6501) );
  NAND2_X1 U7617 ( .A1(n8208), .A2(n8209), .ZN(n6502) );
  NAND2_X1 U7618 ( .A1(n6503), .A2(n8877), .ZN(P3_U3296) );
  NOR2_X1 U7619 ( .A1(n8691), .A2(n7003), .ZN(n6504) );
  NAND2_X1 U7620 ( .A1(n6507), .A2(n6506), .ZN(n6505) );
  NAND3_X1 U7621 ( .A1(n8691), .A2(n9020), .A3(n7004), .ZN(n6507) );
  INV_X1 U7622 ( .A(n8580), .ZN(n6515) );
  NAND2_X1 U7623 ( .A1(n11694), .A2(n8673), .ZN(n6516) );
  NAND2_X1 U7624 ( .A1(n8292), .A2(n8291), .ZN(n8294) );
  NAND2_X1 U7625 ( .A1(n8277), .A2(n8276), .ZN(n6517) );
  NAND2_X1 U7626 ( .A1(n7019), .A2(n8259), .ZN(n8277) );
  NAND2_X1 U7627 ( .A1(n8404), .A2(n8403), .ZN(n8423) );
  NAND2_X1 U7628 ( .A1(n8402), .A2(n8401), .ZN(n8404) );
  NAND2_X1 U7629 ( .A1(n7027), .A2(n7028), .ZN(n8389) );
  NAND2_X1 U7630 ( .A1(n6519), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8541) );
  OAI21_X1 U7631 ( .B1(n8511), .B2(n7026), .A(n7023), .ZN(n6519) );
  NAND3_X1 U7632 ( .A1(n6521), .A2(n14074), .A3(n12192), .ZN(n6520) );
  NAND2_X1 U7633 ( .A1(n12186), .A2(n12185), .ZN(n12191) );
  NAND3_X1 U7634 ( .A1(n6524), .A2(n7127), .A3(n6523), .ZN(n6522) );
  OR2_X1 U7635 ( .A1(n12115), .A2(n12116), .ZN(n6523) );
  NAND2_X1 U7636 ( .A1(n6525), .A2(n12114), .ZN(n6524) );
  NAND2_X1 U7637 ( .A1(n12115), .A2(n12116), .ZN(n6525) );
  NAND2_X1 U7638 ( .A1(n12141), .A2(n12142), .ZN(n6526) );
  NAND3_X1 U7639 ( .A1(n12136), .A2(n12137), .A3(n7119), .ZN(n6527) );
  NAND3_X1 U7640 ( .A1(n6530), .A2(n7131), .A3(n6529), .ZN(n6528) );
  OR2_X1 U7641 ( .A1(n12206), .A2(n12207), .ZN(n6529) );
  NAND2_X1 U7642 ( .A1(n6531), .A2(n12205), .ZN(n6530) );
  NAND2_X1 U7643 ( .A1(n12206), .A2(n12207), .ZN(n6531) );
  NOR2_X2 U7644 ( .A1(n7684), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n7905) );
  NOR2_X2 U7645 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n7627) );
  NAND2_X4 U7646 ( .A1(n10064), .A2(n10906), .ZN(n10660) );
  NAND2_X4 U7647 ( .A1(n8130), .A2(n8129), .ZN(n10064) );
  NAND2_X1 U7648 ( .A1(n6857), .A2(n6855), .ZN(n13788) );
  OAI21_X2 U7649 ( .B1(n13028), .B2(n13027), .A(n13026), .ZN(n13163) );
  OAI21_X2 U7650 ( .B1(n11806), .B2(n6570), .A(n7229), .ZN(n13026) );
  NOR2_X2 U7651 ( .A1(n15165), .A2(n15164), .ZN(n15163) );
  INV_X1 U7652 ( .A(n9854), .ZN(n6532) );
  AND2_X2 U7653 ( .A1(n6851), .A2(n6849), .ZN(n7503) );
  NOR2_X2 U7654 ( .A1(n10562), .A2(n14818), .ZN(n10553) );
  NAND2_X2 U7655 ( .A1(n8089), .A2(n8088), .ZN(n11532) );
  OAI22_X2 U7656 ( .A1(n11942), .A2(n11941), .B1(n11940), .B2(n11939), .ZN(
        n13714) );
  NOR2_X2 U7657 ( .A1(n11768), .A2(n7479), .ZN(n11942) );
  AND2_X1 U7658 ( .A1(n10063), .A2(n14792), .ZN(n6536) );
  AND2_X1 U7659 ( .A1(n10063), .A2(n14792), .ZN(n6537) );
  NAND2_X1 U7660 ( .A1(n11953), .A2(n11952), .ZN(n7263) );
  NOR2_X2 U7661 ( .A1(n14125), .A2(n14545), .ZN(n11843) );
  OR2_X1 U7662 ( .A1(n10172), .A2(n12025), .ZN(n10174) );
  NAND2_X1 U7663 ( .A1(n10071), .A2(n10172), .ZN(n10173) );
  NAND2_X2 U7664 ( .A1(n14602), .A2(n10670), .ZN(n10866) );
  NAND2_X2 U7665 ( .A1(n13723), .A2(n13724), .ZN(n13722) );
  NAND2_X1 U7666 ( .A1(n13747), .A2(n12034), .ZN(n13819) );
  NAND2_X2 U7667 ( .A1(n13819), .A2(n13820), .ZN(n13818) );
  CLKBUF_X1 U7668 ( .A(n14609), .Z(n6538) );
  NAND2_X1 U7669 ( .A1(n14218), .A2(n7594), .ZN(n6539) );
  NOR2_X2 U7670 ( .A1(n8501), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8522) );
  NOR2_X2 U7671 ( .A1(n14410), .A2(n14409), .ZN(n14411) );
  AOI21_X2 U7672 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(n14321), .A(n14364), .ZN(
        n14336) );
  NOR2_X2 U7673 ( .A1(n13509), .A2(n13510), .ZN(n13489) );
  OR2_X2 U7674 ( .A1(n11667), .A2(n14830), .ZN(n13509) );
  OAI21_X2 U7675 ( .B1(n13748), .B2(n13750), .A(n13749), .ZN(n13747) );
  AOI21_X2 U7676 ( .B1(n13722), .B2(n13780), .A(n13779), .ZN(n13748) );
  AND2_X2 U7677 ( .A1(n10064), .A2(n12086), .ZN(n10664) );
  INV_X2 U7678 ( .A(n12331), .ZN(n10693) );
  NOR2_X2 U7679 ( .A1(n13329), .A2(n13317), .ZN(n6913) );
  NOR2_X2 U7680 ( .A1(n13460), .A2(n13601), .ZN(n6911) );
  NAND2_X1 U7681 ( .A1(n6633), .A2(n7166), .ZN(n7164) );
  INV_X1 U7682 ( .A(n7535), .ZN(n7445) );
  OR2_X1 U7683 ( .A1(n14192), .A2(n14497), .ZN(n12272) );
  AOI21_X1 U7684 ( .B1(n7093), .B2(n7097), .A(n9786), .ZN(n7092) );
  NAND2_X1 U7685 ( .A1(n6749), .A2(n6598), .ZN(n11425) );
  XOR2_X1 U7686 ( .A(n13842), .B(n12232), .Z(n12301) );
  NAND2_X1 U7687 ( .A1(n6946), .A2(n6945), .ZN(n13956) );
  INV_X1 U7688 ( .A(n13960), .ZN(n6945) );
  INV_X1 U7689 ( .A(n7081), .ZN(n7080) );
  OAI21_X1 U7690 ( .B1(n7083), .B2(n7082), .A(n13946), .ZN(n7081) );
  INV_X1 U7691 ( .A(n8107), .ZN(n7082) );
  INV_X1 U7692 ( .A(n12236), .ZN(n12260) );
  OAI211_X1 U7693 ( .C1(n12098), .C2(n12099), .A(n12097), .B(n7140), .ZN(
        n12100) );
  NAND2_X1 U7694 ( .A1(n6819), .A2(n6818), .ZN(n9578) );
  NAND2_X1 U7695 ( .A1(n6820), .A2(n6574), .ZN(n6819) );
  AND2_X1 U7696 ( .A1(n7167), .A2(n7161), .ZN(n7160) );
  INV_X1 U7697 ( .A(n12162), .ZN(n7167) );
  NAND2_X1 U7698 ( .A1(n7162), .A2(n7165), .ZN(n7161) );
  INV_X1 U7699 ( .A(n6846), .ZN(n6845) );
  NAND2_X1 U7700 ( .A1(n9677), .A2(n6604), .ZN(n7460) );
  OR2_X1 U7701 ( .A1(n7457), .A2(n7456), .ZN(n7455) );
  INV_X1 U7702 ( .A(n7557), .ZN(n7435) );
  INV_X1 U7703 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n9045) );
  INV_X1 U7704 ( .A(n7444), .ZN(n7443) );
  OAI21_X1 U7705 ( .B1(n7834), .B2(n7445), .A(n7537), .ZN(n7444) );
  AND2_X1 U7706 ( .A1(n7536), .A2(n7539), .ZN(n7537) );
  NAND2_X1 U7707 ( .A1(n12512), .A2(n12385), .ZN(n12388) );
  INV_X1 U7708 ( .A(n12449), .ZN(n7285) );
  INV_X1 U7709 ( .A(n10625), .ZN(n8714) );
  NAND2_X1 U7710 ( .A1(n8855), .A2(n8685), .ZN(n8853) );
  NOR2_X1 U7711 ( .A1(n8939), .A2(n7362), .ZN(n7361) );
  NAND2_X1 U7712 ( .A1(n8364), .A2(n8365), .ZN(n7012) );
  NAND2_X1 U7713 ( .A1(n11017), .A2(n7353), .ZN(n7352) );
  NOR2_X1 U7714 ( .A1(n15202), .A2(n7354), .ZN(n7353) );
  OR2_X1 U7715 ( .A1(n12694), .A2(n12405), .ZN(n8972) );
  NAND2_X1 U7716 ( .A1(n12761), .A2(n8962), .ZN(n7341) );
  NAND2_X1 U7717 ( .A1(n11387), .A2(n11386), .ZN(n11385) );
  AND2_X1 U7718 ( .A1(n8168), .A2(n6679), .ZN(n6678) );
  AND2_X1 U7719 ( .A1(n7365), .A2(n7366), .ZN(n6679) );
  NOR2_X1 U7720 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_27__SCAN_IN), .ZN(
        n7365) );
  AND2_X1 U7721 ( .A1(n8716), .A2(n8165), .ZN(n7323) );
  INV_X1 U7722 ( .A(n8167), .ZN(n8716) );
  NAND2_X1 U7723 ( .A1(n8717), .A2(n7323), .ZN(n8863) );
  NAND2_X1 U7724 ( .A1(n9867), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8223) );
  OR2_X1 U7725 ( .A1(n13548), .A2(n9418), .ZN(n9526) );
  NAND2_X1 U7726 ( .A1(n7103), .A2(n6728), .ZN(n6727) );
  NAND2_X1 U7727 ( .A1(n9521), .A2(n9522), .ZN(n6728) );
  NOR2_X1 U7728 ( .A1(n9513), .A2(n6735), .ZN(n6734) );
  INV_X1 U7729 ( .A(n9511), .ZN(n6735) );
  NAND2_X1 U7730 ( .A1(n12073), .A2(n13193), .ZN(n7199) );
  INV_X1 U7731 ( .A(n9509), .ZN(n6739) );
  AND2_X1 U7732 ( .A1(n9243), .A2(n9242), .ZN(n9783) );
  NAND2_X1 U7733 ( .A1(n7205), .A2(n6772), .ZN(n9312) );
  NOR2_X1 U7734 ( .A1(n13486), .A2(n9777), .ZN(n6772) );
  INV_X1 U7735 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n9041) );
  INV_X1 U7736 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n7569) );
  INV_X1 U7737 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n7568) );
  NAND2_X1 U7738 ( .A1(n7917), .A2(n7916), .ZN(n7390) );
  OR2_X1 U7739 ( .A1(n11950), .A2(n14113), .ZN(n12159) );
  OR2_X1 U7740 ( .A1(n14545), .A2(n11772), .ZN(n12156) );
  NAND2_X1 U7741 ( .A1(n8885), .A2(n8884), .ZN(n12231) );
  NAND2_X1 U7742 ( .A1(n6944), .A2(n12336), .ZN(n8893) );
  INV_X1 U7743 ( .A(n13847), .ZN(n7371) );
  NAND2_X1 U7744 ( .A1(n7053), .A2(n7052), .ZN(n14057) );
  AOI21_X1 U7745 ( .B1(n6549), .B2(n7057), .A(n6614), .ZN(n7052) );
  XNOR2_X1 U7746 ( .A(n7542), .B(SI_16_), .ZN(n7882) );
  NAND2_X1 U7747 ( .A1(n6890), .A2(n7423), .ZN(n6889) );
  AOI21_X1 U7748 ( .B1(n7425), .B2(n7426), .A(n7424), .ZN(n7423) );
  XNOR2_X1 U7749 ( .A(n14237), .B(n6934), .ZN(n14276) );
  XNOR2_X1 U7750 ( .A(n14239), .B(n6932), .ZN(n14275) );
  INV_X1 U7751 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n6932) );
  NAND2_X1 U7752 ( .A1(n7314), .A2(n8961), .ZN(n7313) );
  XNOR2_X1 U7753 ( .A(n10969), .B(n7322), .ZN(n11320) );
  NOR2_X1 U7754 ( .A1(n12540), .A2(n6606), .ZN(n7301) );
  AND4_X1 U7755 ( .A1(n8488), .A2(n8487), .A3(n8486), .A4(n8485), .ZN(n12371)
         );
  NAND2_X1 U7756 ( .A1(n10777), .A2(n10427), .ZN(n6795) );
  NAND2_X1 U7757 ( .A1(n15138), .A2(n6808), .ZN(n15154) );
  NOR2_X1 U7758 ( .A1(n15157), .A2(n6809), .ZN(n6808) );
  INV_X1 U7759 ( .A(n12655), .ZN(n6809) );
  NOR2_X1 U7760 ( .A1(n8956), .A2(n6976), .ZN(n6975) );
  AND2_X1 U7761 ( .A1(n6979), .A2(n6978), .ZN(n6976) );
  INV_X1 U7762 ( .A(n8358), .ZN(n8532) );
  INV_X1 U7763 ( .A(n8532), .ZN(n8673) );
  NAND2_X1 U7764 ( .A1(n8648), .A2(n8647), .ZN(n8657) );
  NAND2_X1 U7765 ( .A1(n7046), .A2(n6565), .ZN(n8648) );
  INV_X1 U7766 ( .A(n7031), .ZN(n7030) );
  OAI21_X1 U7767 ( .B1(n8355), .B2(n7032), .A(n8380), .ZN(n7031) );
  NAND2_X1 U7768 ( .A1(n8356), .A2(n8355), .ZN(n8378) );
  OR2_X1 U7769 ( .A1(n8297), .A2(n8296), .ZN(n8317) );
  NAND2_X1 U7770 ( .A1(n11699), .A2(n11702), .ZN(n11713) );
  AND2_X1 U7771 ( .A1(n14864), .A2(n14865), .ZN(n14861) );
  NAND2_X1 U7772 ( .A1(n6913), .A2(n6912), .ZN(n13294) );
  NAND3_X1 U7773 ( .A1(n13310), .A2(n13300), .A3(n13301), .ZN(n13302) );
  OR2_X1 U7774 ( .A1(n13434), .A2(n13141), .ZN(n7483) );
  NAND2_X1 U7775 ( .A1(n6568), .A2(n9506), .ZN(n7098) );
  NAND2_X1 U7776 ( .A1(n6747), .A2(n6555), .ZN(n6749) );
  NOR2_X1 U7777 ( .A1(n9460), .A2(n13704), .ZN(n14947) );
  AND2_X1 U7778 ( .A1(n6547), .A2(n9054), .ZN(n6720) );
  NAND2_X1 U7779 ( .A1(n6566), .A2(n7404), .ZN(n7396) );
  NAND2_X1 U7780 ( .A1(n14055), .A2(n7079), .ZN(n14040) );
  AND2_X1 U7781 ( .A1(n12293), .A2(n8101), .ZN(n7079) );
  NAND2_X1 U7782 ( .A1(n7086), .A2(n7084), .ZN(n8888) );
  INV_X1 U7783 ( .A(n7085), .ZN(n7084) );
  NAND2_X1 U7784 ( .A1(n7985), .A2(n7984), .ZN(n14147) );
  NAND2_X1 U7785 ( .A1(n6764), .A2(n7717), .ZN(n7718) );
  NAND2_X1 U7786 ( .A1(n6869), .A2(SI_4_), .ZN(n7510) );
  MUX2_X1 U7787 ( .A(n10446), .B(n12563), .S(n10441), .Z(n15170) );
  AND2_X1 U7788 ( .A1(n13034), .A2(n13033), .ZN(n6707) );
  NAND2_X1 U7789 ( .A1(n6467), .A2(n8117), .ZN(n6695) );
  NAND2_X1 U7790 ( .A1(n12092), .A2(n12090), .ZN(n7141) );
  INV_X1 U7791 ( .A(n12111), .ZN(n7118) );
  NAND2_X1 U7792 ( .A1(n12118), .A2(n7128), .ZN(n7127) );
  INV_X1 U7793 ( .A(n12117), .ZN(n7128) );
  AOI21_X1 U7794 ( .B1(n6551), .B2(n7146), .A(n7145), .ZN(n7144) );
  NAND2_X1 U7795 ( .A1(n12139), .A2(n7120), .ZN(n7119) );
  INV_X1 U7796 ( .A(n12138), .ZN(n7120) );
  NAND2_X1 U7797 ( .A1(n9551), .A2(n9550), .ZN(n9566) );
  NOR2_X1 U7798 ( .A1(n9587), .A2(n9584), .ZN(n7449) );
  INV_X1 U7799 ( .A(n9584), .ZN(n7448) );
  AOI21_X1 U7800 ( .B1(n7157), .B2(n7159), .A(n6585), .ZN(n7156) );
  INV_X1 U7801 ( .A(n7160), .ZN(n7159) );
  AOI21_X1 U7802 ( .B1(n9623), .B2(n9624), .A(n6630), .ZN(n6848) );
  OR2_X1 U7803 ( .A1(n9617), .A2(n7463), .ZN(n7462) );
  NOR2_X1 U7804 ( .A1(n6596), .A2(n7464), .ZN(n7463) );
  AND2_X1 U7805 ( .A1(n6558), .A2(n6847), .ZN(n6846) );
  OR2_X1 U7806 ( .A1(n9623), .A2(n9624), .ZN(n6847) );
  INV_X1 U7807 ( .A(n6640), .ZN(n7467) );
  INV_X1 U7808 ( .A(n7152), .ZN(n7148) );
  NOR2_X1 U7809 ( .A1(n7152), .A2(n7150), .ZN(n7149) );
  NAND2_X1 U7810 ( .A1(n12204), .A2(n7137), .ZN(n7136) );
  INV_X1 U7811 ( .A(n12203), .ZN(n7137) );
  NOR3_X1 U7812 ( .A1(n8772), .A2(n8771), .A3(n14451), .ZN(n8781) );
  NAND2_X1 U7813 ( .A1(n9640), .A2(n6548), .ZN(n7474) );
  OR2_X1 U7814 ( .A1(n9635), .A2(n7475), .ZN(n7473) );
  OR2_X1 U7815 ( .A1(n7460), .A2(n9681), .ZN(n7458) );
  AND2_X1 U7816 ( .A1(n7460), .A2(n9681), .ZN(n7456) );
  OR2_X1 U7817 ( .A1(n7461), .A2(n9681), .ZN(n7459) );
  NAND2_X1 U7818 ( .A1(n12209), .A2(n7132), .ZN(n7131) );
  INV_X1 U7819 ( .A(n12208), .ZN(n7132) );
  NAND2_X1 U7820 ( .A1(n12219), .A2(n7124), .ZN(n7123) );
  INV_X1 U7821 ( .A(n12218), .ZN(n7124) );
  NAND2_X1 U7822 ( .A1(n9695), .A2(n6575), .ZN(n9700) );
  NOR2_X1 U7823 ( .A1(n6832), .A2(n6831), .ZN(n6830) );
  NOR2_X1 U7824 ( .A1(n9699), .A2(n9698), .ZN(n6831) );
  AND2_X1 U7825 ( .A1(n6834), .A2(n6833), .ZN(n6832) );
  INV_X1 U7826 ( .A(n6641), .ZN(n6834) );
  AND2_X1 U7827 ( .A1(n6636), .A2(n6825), .ZN(n6824) );
  NAND2_X1 U7828 ( .A1(n9719), .A2(n9718), .ZN(n7472) );
  INV_X1 U7829 ( .A(n12235), .ZN(n7170) );
  NAND2_X1 U7830 ( .A1(n7173), .A2(n7172), .ZN(n7171) );
  INV_X1 U7831 ( .A(n12257), .ZN(n7172) );
  INV_X1 U7832 ( .A(n12258), .ZN(n7173) );
  NAND2_X1 U7833 ( .A1(n7640), .A2(n7639), .ZN(n12084) );
  AOI21_X1 U7834 ( .B1(n7433), .B2(n7435), .A(n7430), .ZN(n7429) );
  INV_X1 U7835 ( .A(n7434), .ZN(n7433) );
  AOI21_X1 U7836 ( .B1(n6550), .B2(n6897), .A(n6659), .ZN(n6892) );
  NAND2_X1 U7837 ( .A1(n7789), .A2(n7425), .ZN(n6890) );
  NOR2_X1 U7838 ( .A1(n7804), .A2(n7428), .ZN(n7427) );
  INV_X1 U7839 ( .A(n7528), .ZN(n7428) );
  AND2_X1 U7840 ( .A1(n8854), .A2(n12681), .ZN(n8690) );
  INV_X1 U7841 ( .A(n12628), .ZN(n6801) );
  INV_X1 U7842 ( .A(n12662), .ZN(n6959) );
  OR2_X1 U7843 ( .A1(n12558), .A2(n14455), .ZN(n8773) );
  OR2_X1 U7844 ( .A1(n15190), .A2(n11391), .ZN(n8756) );
  OR2_X1 U7845 ( .A1(n12562), .A2(n15196), .ZN(n8755) );
  INV_X1 U7846 ( .A(n6985), .ZN(n6984) );
  AND2_X1 U7847 ( .A1(n10431), .A2(n6533), .ZN(n8274) );
  NAND2_X1 U7848 ( .A1(n13010), .A2(n8673), .ZN(n7015) );
  NAND2_X1 U7849 ( .A1(n8819), .A2(n6992), .ZN(n6991) );
  INV_X1 U7850 ( .A(n8820), .ZN(n6992) );
  INV_X1 U7851 ( .A(n8823), .ZN(n6989) );
  INV_X1 U7852 ( .A(n7335), .ZN(n7334) );
  OAI21_X1 U7853 ( .B1(n8956), .B2(n7336), .A(n8958), .ZN(n7335) );
  INV_X1 U7854 ( .A(n8957), .ZN(n7336) );
  INV_X1 U7855 ( .A(n7000), .ZN(n6997) );
  NAND2_X1 U7856 ( .A1(n15191), .A2(n8931), .ZN(n11387) );
  NAND2_X1 U7857 ( .A1(n8989), .A2(n8987), .ZN(n7304) );
  INV_X1 U7858 ( .A(n8316), .ZN(n7042) );
  NAND2_X1 U7859 ( .A1(n9878), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8259) );
  INV_X1 U7860 ( .A(n13125), .ZN(n7227) );
  INV_X1 U7861 ( .A(n13183), .ZN(n9525) );
  INV_X1 U7862 ( .A(n9522), .ZN(n6724) );
  NOR2_X1 U7863 ( .A1(n13357), .A2(n7105), .ZN(n7104) );
  INV_X1 U7864 ( .A(n9523), .ZN(n7105) );
  INV_X1 U7865 ( .A(n9397), .ZN(n7211) );
  INV_X1 U7866 ( .A(n13357), .ZN(n7212) );
  NOR2_X1 U7867 ( .A1(n13580), .A2(n13404), .ZN(n6908) );
  NOR2_X1 U7868 ( .A1(n13404), .A2(n13189), .ZN(n7178) );
  INV_X1 U7869 ( .A(n6761), .ZN(n6760) );
  NAND2_X1 U7870 ( .A1(n6762), .A2(n13399), .ZN(n6756) );
  INV_X1 U7871 ( .A(n7178), .ZN(n6757) );
  NOR2_X1 U7872 ( .A1(n7493), .A2(n7189), .ZN(n7188) );
  INV_X1 U7873 ( .A(n9243), .ZN(n7189) );
  NOR2_X1 U7874 ( .A1(n11288), .A2(n6745), .ZN(n6746) );
  INV_X1 U7875 ( .A(n9491), .ZN(n6745) );
  INV_X1 U7876 ( .A(n7113), .ZN(n7112) );
  AOI21_X1 U7877 ( .B1(n7113), .B2(n7111), .A(n6615), .ZN(n7110) );
  NOR2_X1 U7878 ( .A1(n13385), .A2(n7114), .ZN(n7113) );
  INV_X1 U7879 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n9055) );
  INV_X1 U7880 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9456) );
  NAND2_X1 U7881 ( .A1(n9340), .A2(n7248), .ZN(n7247) );
  INV_X1 U7882 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n7248) );
  NAND2_X1 U7883 ( .A1(n7775), .A2(n6935), .ZN(n7806) );
  INV_X1 U7884 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6935) );
  NAND2_X1 U7885 ( .A1(n8878), .A2(n8052), .ZN(n12298) );
  INV_X1 U7886 ( .A(n7954), .ZN(n7406) );
  INV_X1 U7887 ( .A(n7077), .ZN(n7076) );
  OAI21_X1 U7888 ( .B1(n12290), .B2(n7078), .A(n14503), .ZN(n7077) );
  INV_X1 U7889 ( .A(n8096), .ZN(n7078) );
  INV_X1 U7890 ( .A(n11842), .ZN(n8095) );
  INV_X1 U7891 ( .A(n7064), .ZN(n7063) );
  OAI21_X1 U7892 ( .B1(n12284), .B2(n7065), .A(n14523), .ZN(n7064) );
  INV_X1 U7893 ( .A(n8090), .ZN(n7065) );
  INV_X1 U7894 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7779) );
  OR2_X1 U7895 ( .A1(n12090), .A2(n12092), .ZN(n12095) );
  INV_X1 U7896 ( .A(n12090), .ZN(n7660) );
  NAND2_X1 U7897 ( .A1(n6899), .A2(n6602), .ZN(n13963) );
  NAND2_X1 U7898 ( .A1(n11624), .A2(n12285), .ZN(n11629) );
  NAND2_X1 U7899 ( .A1(n14227), .A2(n14511), .ZN(n12249) );
  NAND2_X1 U7900 ( .A1(n8883), .A2(n8882), .ZN(n9737) );
  AND4_X1 U7901 ( .A1(n7573), .A2(n7572), .A3(n10344), .A4(n8131), .ZN(n7574)
         );
  NAND2_X1 U7902 ( .A1(n7935), .A2(n7142), .ZN(n8057) );
  NOR2_X1 U7903 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n7142) );
  AOI21_X1 U7904 ( .B1(n7443), .B2(n7445), .A(n7441), .ZN(n7440) );
  INV_X1 U7905 ( .A(n7541), .ZN(n7441) );
  NAND2_X1 U7906 ( .A1(n7526), .A2(SI_10_), .ZN(n7528) );
  XNOR2_X1 U7907 ( .A(n7529), .B(SI_11_), .ZN(n7804) );
  NAND2_X1 U7908 ( .A1(n7520), .A2(SI_8_), .ZN(n7522) );
  OR2_X1 U7909 ( .A1(n7754), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n7772) );
  INV_X1 U7910 ( .A(n14282), .ZN(n14281) );
  XNOR2_X1 U7911 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n14280) );
  NAND2_X1 U7912 ( .A1(n6925), .A2(n6923), .ZN(n14233) );
  NAND2_X1 U7913 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n6924), .ZN(n6923) );
  INV_X1 U7914 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6924) );
  NAND2_X1 U7915 ( .A1(n6933), .A2(n14238), .ZN(n14239) );
  NAND2_X1 U7916 ( .A1(n14276), .A2(n14639), .ZN(n6933) );
  INV_X1 U7917 ( .A(n12387), .ZN(n7315) );
  INV_X1 U7918 ( .A(n12388), .ZN(n7316) );
  AOI21_X1 U7919 ( .B1(n7301), .B2(n6569), .A(n6561), .ZN(n7300) );
  INV_X1 U7920 ( .A(n12367), .ZN(n7303) );
  OR2_X1 U7921 ( .A1(n7296), .A2(n6588), .ZN(n7293) );
  AOI21_X1 U7922 ( .B1(n7298), .B2(n7300), .A(n7297), .ZN(n7296) );
  INV_X1 U7923 ( .A(n12474), .ZN(n7297) );
  INV_X1 U7924 ( .A(n7301), .ZN(n7298) );
  NAND2_X1 U7925 ( .A1(n12388), .A2(n12387), .ZN(n12491) );
  NAND2_X1 U7926 ( .A1(n8328), .A2(n11328), .ZN(n8346) );
  INV_X1 U7927 ( .A(n11467), .ZN(n11317) );
  OR2_X1 U7928 ( .A1(n11325), .A2(n11326), .ZN(n7321) );
  AOI21_X1 U7929 ( .B1(n6546), .B2(n7280), .A(n12379), .ZN(n7279) );
  INV_X1 U7930 ( .A(n6572), .ZN(n7280) );
  NAND2_X1 U7931 ( .A1(n7319), .A2(n6573), .ZN(n7318) );
  NAND2_X1 U7932 ( .A1(n11410), .A2(n6573), .ZN(n7317) );
  AND2_X1 U7933 ( .A1(n8384), .A2(n8383), .ZN(n11641) );
  AND2_X1 U7934 ( .A1(n7293), .A2(n7291), .ZN(n7290) );
  INV_X1 U7935 ( .A(n12482), .ZN(n7291) );
  OR2_X1 U7936 ( .A1(n7299), .A2(n6588), .ZN(n7294) );
  INV_X1 U7937 ( .A(n7300), .ZN(n7299) );
  NAND2_X1 U7938 ( .A1(n8715), .A2(n8714), .ZN(n8859) );
  OR2_X1 U7939 ( .A1(n8690), .A2(n12676), .ZN(n7005) );
  AOI21_X1 U7940 ( .B1(n8690), .B2(n12676), .A(n8975), .ZN(n7004) );
  AOI211_X1 U7941 ( .C1(n9015), .C2(n8972), .A(n8686), .B(n8853), .ZN(n8691)
         );
  AND4_X1 U7942 ( .A1(n8315), .A2(n8314), .A3(n8313), .A4(n8312), .ZN(n11452)
         );
  NOR2_X1 U7943 ( .A1(n6954), .A2(n10490), .ZN(n6953) );
  INV_X1 U7944 ( .A(n10438), .ZN(n6954) );
  NAND2_X1 U7945 ( .A1(n10479), .A2(n10480), .ZN(n6804) );
  NAND2_X1 U7946 ( .A1(n6952), .A2(n10490), .ZN(n10486) );
  NAND2_X1 U7947 ( .A1(n10461), .A2(n10438), .ZN(n6952) );
  NAND2_X1 U7948 ( .A1(n10486), .A2(n6950), .ZN(n10488) );
  AND2_X1 U7949 ( .A1(n6951), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n6950) );
  NAND2_X1 U7950 ( .A1(n6967), .A2(n6966), .ZN(n6965) );
  INV_X1 U7951 ( .A(n15026), .ZN(n6966) );
  OR2_X1 U7952 ( .A1(n15069), .A2(n15068), .ZN(n6687) );
  OR2_X1 U7953 ( .A1(n15127), .A2(n6662), .ZN(n6964) );
  NAND2_X1 U7954 ( .A1(n6957), .A2(n12662), .ZN(n12579) );
  INV_X1 U7955 ( .A(n15163), .ZN(n6957) );
  INV_X1 U7956 ( .A(n7358), .ZN(n7357) );
  AOI21_X1 U7957 ( .B1(n7358), .B2(n7356), .A(n6608), .ZN(n7355) );
  NAND2_X1 U7958 ( .A1(n7360), .A2(n8938), .ZN(n11611) );
  NOR2_X1 U7959 ( .A1(n11615), .A2(n7359), .ZN(n7358) );
  INV_X1 U7960 ( .A(n8938), .ZN(n7359) );
  NAND2_X1 U7961 ( .A1(n8937), .A2(n7361), .ZN(n7360) );
  AND4_X1 U7962 ( .A1(n8422), .A2(n8421), .A3(n8420), .A4(n8419), .ZN(n12363)
         );
  INV_X1 U7963 ( .A(n12559), .ZN(n14453) );
  AOI21_X1 U7964 ( .B1(n7327), .B2(n7330), .A(n6590), .ZN(n7325) );
  INV_X1 U7965 ( .A(n15192), .ZN(n15187) );
  AOI21_X1 U7966 ( .B1(n7339), .B2(n7338), .A(n6601), .ZN(n7337) );
  INV_X1 U7967 ( .A(n8962), .ZN(n7338) );
  OR2_X1 U7968 ( .A1(n12954), .A2(n8961), .ZN(n12747) );
  NAND2_X1 U7969 ( .A1(n7342), .A2(n8698), .ZN(n12766) );
  AND2_X1 U7970 ( .A1(n8823), .A2(n8824), .ZN(n12774) );
  NAND2_X1 U7971 ( .A1(n8810), .A2(n12821), .ZN(n6979) );
  NAND2_X1 U7972 ( .A1(n6634), .A2(n8810), .ZN(n6978) );
  INV_X1 U7973 ( .A(n8803), .ZN(n6980) );
  AND2_X1 U7974 ( .A1(n8540), .A2(n8539), .ZN(n12808) );
  INV_X1 U7975 ( .A(n7347), .ZN(n7346) );
  AND2_X1 U7976 ( .A1(n8954), .A2(n7344), .ZN(n7343) );
  NAND2_X1 U7977 ( .A1(n7347), .A2(n7345), .ZN(n7344) );
  OR2_X1 U7978 ( .A1(n10430), .A2(n8977), .ZN(n15243) );
  OR2_X1 U7979 ( .A1(n12986), .A2(n12807), .ZN(n8803) );
  NAND2_X1 U7980 ( .A1(n8489), .A2(n8807), .ZN(n12822) );
  INV_X1 U7981 ( .A(n8785), .ZN(n6999) );
  NAND2_X1 U7982 ( .A1(n8400), .A2(n8778), .ZN(n11829) );
  NOR2_X1 U7983 ( .A1(n8943), .A2(n7001), .ZN(n7000) );
  INV_X1 U7984 ( .A(n15259), .ZN(n15241) );
  NAND2_X1 U7985 ( .A1(n8992), .A2(n8991), .ZN(n10505) );
  NAND2_X1 U7986 ( .A1(n8169), .A2(n8180), .ZN(n6973) );
  OAI22_X1 U7987 ( .A1(n8657), .A2(n8656), .B1(P2_DATAO_REG_29__SCAN_IN), .B2(
        n13691), .ZN(n8668) );
  NOR2_X1 U7988 ( .A1(n8630), .A2(n7048), .ZN(n7047) );
  INV_X1 U7989 ( .A(n8618), .ZN(n7048) );
  NOR2_X1 U7990 ( .A1(n8167), .A2(n8166), .ZN(n8168) );
  NAND2_X1 U7991 ( .A1(n8717), .A2(n8716), .ZN(n8719) );
  NAND2_X1 U7992 ( .A1(n8696), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8697) );
  AOI21_X1 U7993 ( .B1(n7036), .B2(n7038), .A(n7035), .ZN(n7034) );
  INV_X1 U7994 ( .A(n8493), .ZN(n7035) );
  NAND2_X1 U7995 ( .A1(n8463), .A2(n8462), .ZN(n8477) );
  OAI21_X1 U7996 ( .B1(n8423), .B2(n7022), .A(n8443), .ZN(n7021) );
  INV_X1 U7997 ( .A(n8426), .ZN(n7022) );
  NAND2_X1 U7998 ( .A1(n8423), .A2(n8405), .ZN(n8406) );
  OR2_X1 U7999 ( .A1(n8404), .A2(n8403), .ZN(n8405) );
  INV_X1 U8000 ( .A(n8377), .ZN(n7032) );
  AND2_X1 U8001 ( .A1(n8377), .A2(n8354), .ZN(n8355) );
  NAND2_X1 U8002 ( .A1(n9899), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8316) );
  AND2_X1 U8003 ( .A1(n8334), .A2(n8319), .ZN(n8320) );
  INV_X1 U8004 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n8318) );
  NAND2_X1 U8005 ( .A1(n8317), .A2(n8316), .ZN(n8321) );
  AND2_X1 U8006 ( .A1(n7045), .A2(n8320), .ZN(n7044) );
  NAND2_X1 U8007 ( .A1(n8296), .A2(n8316), .ZN(n7045) );
  NAND2_X1 U8008 ( .A1(n9868), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8241) );
  OR3_X1 U8009 ( .A1(n11864), .A2(n13710), .A3(n13704), .ZN(n9848) );
  OR2_X1 U8010 ( .A1(n12420), .A2(n11053), .ZN(n11054) );
  NOR2_X1 U8011 ( .A1(n7227), .A2(n7225), .ZN(n7224) );
  INV_X1 U8012 ( .A(n13041), .ZN(n7225) );
  AND2_X1 U8013 ( .A1(n13053), .A2(n13051), .ZN(n13111) );
  INV_X1 U8014 ( .A(n7485), .ZN(n7232) );
  INV_X1 U8015 ( .A(n11809), .ZN(n7233) );
  NAND2_X1 U8016 ( .A1(n9037), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n9388) );
  INV_X1 U8017 ( .A(n13201), .ZN(n11256) );
  NAND2_X1 U8018 ( .A1(n11708), .A2(n11698), .ZN(n11712) );
  INV_X1 U8019 ( .A(n9832), .ZN(n9833) );
  NAND2_X1 U8020 ( .A1(n7437), .A2(n7436), .ZN(n6684) );
  NAND2_X1 U8021 ( .A1(n9831), .A2(n6840), .ZN(n7436) );
  INV_X1 U8022 ( .A(n9732), .ZN(n9735) );
  OR2_X1 U8023 ( .A1(n9123), .A2(n11135), .ZN(n9107) );
  NOR2_X1 U8024 ( .A1(n14861), .A2(n6620), .ZN(n10120) );
  OR2_X1 U8025 ( .A1(n10120), .A2(n10119), .ZN(n6783) );
  NOR2_X1 U8026 ( .A1(n11915), .A2(n6784), .ZN(n14892) );
  AND2_X1 U8027 ( .A1(n10103), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6784) );
  NOR2_X1 U8028 ( .A1(n14892), .A2(n14891), .ZN(n14890) );
  NOR2_X1 U8029 ( .A1(n14906), .A2(n6652), .ZN(n10748) );
  NOR2_X1 U8030 ( .A1(n10747), .A2(n10748), .ZN(n10848) );
  OR2_X1 U8031 ( .A1(n11103), .A2(n11104), .ZN(n6781) );
  AND2_X1 U8032 ( .A1(n6781), .A2(n6780), .ZN(n11484) );
  NAND2_X1 U8033 ( .A1(n11482), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6780) );
  OR2_X1 U8034 ( .A1(n11484), .A2(n11483), .ZN(n6779) );
  AND2_X1 U8035 ( .A1(n9053), .A2(n9054), .ZN(n6835) );
  NAND2_X1 U8036 ( .A1(n9526), .A2(n9419), .ZN(n13292) );
  INV_X1 U8037 ( .A(n13308), .ZN(n13311) );
  NAND2_X1 U8038 ( .A1(n13312), .A2(n13311), .ZN(n13310) );
  AND2_X1 U8039 ( .A1(n13567), .A2(n13186), .ZN(n9397) );
  NAND2_X1 U8040 ( .A1(n7213), .A2(n7212), .ZN(n7209) );
  INV_X1 U8041 ( .A(n13356), .ZN(n7213) );
  NAND2_X1 U8042 ( .A1(n13352), .A2(n13357), .ZN(n7102) );
  INV_X1 U8043 ( .A(n7209), .ZN(n13355) );
  NAND2_X1 U8044 ( .A1(n6725), .A2(n9522), .ZN(n13352) );
  OR2_X1 U8045 ( .A1(n13366), .A2(n9521), .ZN(n6725) );
  AND2_X1 U8046 ( .A1(n7180), .A2(n9362), .ZN(n6761) );
  NAND2_X1 U8047 ( .A1(n13418), .A2(n9516), .ZN(n7180) );
  OR2_X1 U8048 ( .A1(n13596), .A2(n13191), .ZN(n9362) );
  NAND2_X1 U8049 ( .A1(n6911), .A2(n13434), .ZN(n13429) );
  INV_X1 U8050 ( .A(n6734), .ZN(n6733) );
  AOI21_X1 U8051 ( .B1(n6734), .B2(n6738), .A(n6556), .ZN(n6732) );
  NAND2_X1 U8052 ( .A1(n13446), .A2(n9351), .ZN(n13424) );
  NAND2_X1 U8053 ( .A1(n9326), .A2(n7199), .ZN(n7197) );
  NAND2_X1 U8054 ( .A1(n6632), .A2(n7199), .ZN(n7196) );
  NAND2_X1 U8055 ( .A1(n13474), .A2(n9326), .ZN(n7198) );
  INV_X1 U8056 ( .A(n13473), .ZN(n9325) );
  NAND2_X1 U8057 ( .A1(n9325), .A2(n9786), .ZN(n13476) );
  AOI21_X1 U8058 ( .B1(n7096), .B2(n7094), .A(n6619), .ZN(n7093) );
  INV_X1 U8059 ( .A(n6568), .ZN(n7094) );
  NAND2_X1 U8060 ( .A1(n6771), .A2(n6769), .ZN(n7205) );
  NOR2_X1 U8061 ( .A1(n9776), .A2(n6770), .ZN(n6769) );
  INV_X1 U8062 ( .A(n9286), .ZN(n6770) );
  NAND2_X1 U8063 ( .A1(n6721), .A2(n9504), .ZN(n13502) );
  NAND2_X1 U8064 ( .A1(n11664), .A2(n9503), .ZN(n6721) );
  AOI21_X1 U8065 ( .B1(n7184), .B2(n7186), .A(n6611), .ZN(n7182) );
  NAND2_X1 U8066 ( .A1(n7190), .A2(n6592), .ZN(n7187) );
  NAND2_X1 U8067 ( .A1(n9244), .A2(n7188), .ZN(n7183) );
  AOI21_X1 U8068 ( .B1(n7185), .B2(n7187), .A(n11578), .ZN(n7184) );
  INV_X1 U8069 ( .A(n7188), .ZN(n7185) );
  INV_X1 U8070 ( .A(n7187), .ZN(n7186) );
  NAND2_X1 U8071 ( .A1(n9500), .A2(n11596), .ZN(n11601) );
  INV_X1 U8072 ( .A(n11603), .ZN(n9500) );
  AND2_X1 U8073 ( .A1(n11598), .A2(n11606), .ZN(n11599) );
  NAND2_X1 U8074 ( .A1(n7200), .A2(n7201), .ZN(n11342) );
  AOI21_X1 U8075 ( .B1(n9782), .B2(n7203), .A(n7202), .ZN(n7201) );
  INV_X1 U8076 ( .A(n9231), .ZN(n7202) );
  NOR2_X2 U8077 ( .A1(n11357), .A2(n11493), .ZN(n11598) );
  AOI21_X1 U8078 ( .B1(n9493), .B2(n7100), .A(n6586), .ZN(n7099) );
  INV_X1 U8079 ( .A(n9492), .ZN(n7100) );
  AOI21_X1 U8080 ( .B1(n11288), .B2(n7193), .A(n6609), .ZN(n7191) );
  INV_X1 U8081 ( .A(n11121), .ZN(n6748) );
  NAND2_X1 U8082 ( .A1(n6747), .A2(n6746), .ZN(n11282) );
  OAI22_X1 U8083 ( .A1(n10575), .A2(n10576), .B1(n11131), .B2(n9552), .ZN(
        n10565) );
  XNOR2_X1 U8084 ( .A(n9552), .B(n11131), .ZN(n10575) );
  NAND2_X1 U8085 ( .A1(n10575), .A2(n10573), .ZN(n10572) );
  NAND2_X1 U8086 ( .A1(n9399), .A2(n9398), .ZN(n13317) );
  INV_X1 U8087 ( .A(n9133), .ZN(n9746) );
  AND2_X1 U8088 ( .A1(n6547), .A2(n7470), .ZN(n7469) );
  NOR2_X1 U8089 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n7470) );
  INV_X1 U8090 ( .A(n9053), .ZN(n6838) );
  INV_X1 U8091 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n9071) );
  NAND2_X1 U8092 ( .A1(n7469), .A2(n9327), .ZN(n9072) );
  NOR2_X1 U8093 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n9130) );
  NAND2_X1 U8094 ( .A1(n9454), .A2(n9042), .ZN(n6787) );
  OR2_X1 U8095 ( .A1(n7759), .A2(n7758), .ZN(n7780) );
  NAND2_X1 U8096 ( .A1(n10070), .A2(n10069), .ZN(n10172) );
  NAND2_X1 U8097 ( .A1(n7826), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7842) );
  NAND2_X1 U8098 ( .A1(n6577), .A2(n7269), .ZN(n7268) );
  INV_X1 U8099 ( .A(n7270), .ZN(n7269) );
  NOR2_X1 U8100 ( .A1(n7780), .A2(n7779), .ZN(n7812) );
  NAND2_X1 U8101 ( .A1(n12307), .A2(n12268), .ZN(n12269) );
  AND4_X1 U8102 ( .A1(n7881), .A2(n7880), .A3(n7879), .A4(n7878), .ZN(n14113)
         );
  OR2_X1 U8103 ( .A1(n11887), .A2(n11886), .ZN(n6880) );
  NAND2_X1 U8104 ( .A1(n14160), .A2(n6901), .ZN(n6900) );
  INV_X1 U8105 ( .A(n13848), .ZN(n6901) );
  NOR2_X1 U8106 ( .A1(n14002), .A2(n7072), .ZN(n7071) );
  INV_X1 U8107 ( .A(n8103), .ZN(n7072) );
  NAND2_X1 U8108 ( .A1(n14020), .A2(n14025), .ZN(n14021) );
  NAND2_X1 U8109 ( .A1(n14099), .A2(n6940), .ZN(n14054) );
  AOI21_X1 U8110 ( .B1(n7382), .B2(n7389), .A(n7381), .ZN(n7380) );
  INV_X1 U8111 ( .A(n12194), .ZN(n7381) );
  NOR2_X1 U8112 ( .A1(n12190), .A2(n7059), .ZN(n7058) );
  INV_X1 U8113 ( .A(n12271), .ZN(n7059) );
  AND2_X1 U8114 ( .A1(n12193), .A2(n12194), .ZN(n14074) );
  INV_X1 U8115 ( .A(n14096), .ZN(n7385) );
  AOI21_X1 U8116 ( .B1(n7388), .B2(n7387), .A(n6582), .ZN(n7386) );
  INV_X1 U8117 ( .A(n7916), .ZN(n7387) );
  NAND2_X1 U8118 ( .A1(n8095), .A2(n12290), .ZN(n11840) );
  NAND2_X1 U8119 ( .A1(n7871), .A2(n7870), .ZN(n11950) );
  AND2_X1 U8120 ( .A1(n12286), .A2(n7394), .ZN(n7393) );
  OR2_X1 U8121 ( .A1(n12285), .A2(n7395), .ZN(n7394) );
  INV_X1 U8122 ( .A(n7833), .ZN(n7395) );
  NAND2_X1 U8123 ( .A1(n11629), .A2(n7833), .ZN(n11650) );
  NAND2_X1 U8124 ( .A1(n14655), .A2(n7787), .ZN(n11535) );
  AND2_X1 U8125 ( .A1(n12281), .A2(n7749), .ZN(n7408) );
  INV_X1 U8126 ( .A(n14689), .ZN(n7714) );
  INV_X1 U8127 ( .A(n14690), .ZN(n7715) );
  AND3_X2 U8128 ( .A1(n7631), .A2(n7630), .A3(n7629), .ZN(n11902) );
  AOI21_X1 U8129 ( .B1(n12231), .B2(n14761), .A(n8894), .ZN(n6949) );
  NAND2_X1 U8130 ( .A1(n8021), .A2(n8020), .ZN(n14137) );
  INV_X1 U8131 ( .A(n14056), .ZN(n8099) );
  INV_X1 U8132 ( .A(n14104), .ZN(n14192) );
  INV_X1 U8133 ( .A(n14761), .ZN(n14781) );
  INV_X1 U8134 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n6853) );
  NAND2_X1 U8135 ( .A1(n6894), .A2(n6895), .ZN(n7901) );
  OR2_X1 U8136 ( .A1(n7439), .A2(n6897), .ZN(n6894) );
  NAND2_X1 U8137 ( .A1(n7789), .A2(n7788), .ZN(n7791) );
  INV_X1 U8138 ( .A(n7414), .ZN(n7413) );
  OAI21_X1 U8139 ( .B1(n7732), .B2(n7415), .A(n7751), .ZN(n7414) );
  NAND2_X1 U8140 ( .A1(n7733), .A2(n7732), .ZN(n7735) );
  OR2_X1 U8141 ( .A1(n6891), .A2(n7679), .ZN(n6763) );
  NOR2_X1 U8142 ( .A1(n6891), .A2(n6866), .ZN(n6864) );
  NAND2_X1 U8143 ( .A1(n7671), .A2(n7508), .ZN(n7680) );
  NAND2_X1 U8144 ( .A1(n7626), .A2(n7502), .ZN(n7648) );
  CLKBUF_X1 U8145 ( .A(n7627), .Z(n7628) );
  NOR2_X1 U8146 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6875) );
  XNOR2_X1 U8147 ( .A(n14281), .B(n6682), .ZN(n14284) );
  INV_X1 U8148 ( .A(n14280), .ZN(n6682) );
  XNOR2_X1 U8149 ( .A(n14233), .B(n6922), .ZN(n14277) );
  INV_X1 U8150 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n6922) );
  NOR2_X1 U8151 ( .A1(n15339), .A2(n14301), .ZN(n14304) );
  OAI21_X1 U8152 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n14255), .A(n14254), .ZN(
        n14270) );
  AND2_X1 U8153 ( .A1(n6914), .A2(n14579), .ZN(n14320) );
  OAI21_X1 U8154 ( .B1(n14580), .B2(n14581), .A(n6915), .ZN(n6914) );
  INV_X1 U8155 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6915) );
  NAND2_X1 U8156 ( .A1(n8874), .A2(n8873), .ZN(n10607) );
  XNOR2_X1 U8157 ( .A(n11386), .B(n12386), .ZN(n11465) );
  XNOR2_X1 U8158 ( .A(n11320), .B(n11452), .ZN(n11467) );
  INV_X1 U8159 ( .A(n12557), .ZN(n14454) );
  INV_X1 U8160 ( .A(n12393), .ZN(n12553) );
  INV_X1 U8161 ( .A(n12363), .ZN(n12556) );
  NAND2_X1 U8162 ( .A1(n10463), .A2(n10462), .ZN(n10461) );
  AND2_X1 U8163 ( .A1(n10481), .A2(n6796), .ZN(n6802) );
  NAND2_X1 U8164 ( .A1(n6631), .A2(n6795), .ZN(n6803) );
  NOR2_X1 U8165 ( .A1(n10446), .A2(n10433), .ZN(n15054) );
  NOR2_X1 U8166 ( .A1(n15129), .A2(n15128), .ZN(n15127) );
  NAND2_X1 U8167 ( .A1(n15120), .A2(n6664), .ZN(n15138) );
  XNOR2_X1 U8168 ( .A(n6964), .B(n15151), .ZN(n15145) );
  NOR2_X1 U8169 ( .A1(n15145), .A2(n11835), .ZN(n15144) );
  NOR2_X1 U8170 ( .A1(n14435), .A2(n6816), .ZN(n6815) );
  INV_X1 U8171 ( .A(n12673), .ZN(n6814) );
  NAND2_X1 U8172 ( .A1(n6812), .A2(n6811), .ZN(n6810) );
  INV_X1 U8173 ( .A(n12677), .ZN(n6811) );
  NAND2_X1 U8174 ( .A1(n12678), .A2(n15176), .ZN(n6812) );
  OR2_X1 U8175 ( .A1(n10627), .A2(n12676), .ZN(n15267) );
  NOR2_X1 U8176 ( .A1(n8984), .A2(n8981), .ZN(n7369) );
  NAND2_X1 U8177 ( .A1(n8520), .A2(n8519), .ZN(n12982) );
  NAND2_X1 U8178 ( .A1(n8482), .A2(n8481), .ZN(n12992) );
  NAND2_X1 U8179 ( .A1(n8454), .A2(n8453), .ZN(n13004) );
  OR2_X1 U8180 ( .A1(n10030), .A2(n8532), .ZN(n8454) );
  NAND2_X1 U8181 ( .A1(n8434), .A2(n8433), .ZN(n14374) );
  NOR2_X1 U8182 ( .A1(n13063), .A2(n7235), .ZN(n7234) );
  INV_X1 U8183 ( .A(n13059), .ZN(n7235) );
  NAND2_X1 U8184 ( .A1(n13179), .A2(n13059), .ZN(n13062) );
  NAND2_X1 U8185 ( .A1(n13071), .A2(n13041), .ZN(n13072) );
  NAND2_X1 U8186 ( .A1(n13126), .A2(n13125), .ZN(n13124) );
  NAND2_X1 U8187 ( .A1(n13142), .A2(n13032), .ZN(n7236) );
  NAND2_X1 U8188 ( .A1(n10933), .A2(n11157), .ZN(n11169) );
  INV_X2 U8189 ( .A(n13148), .ZN(n14824) );
  XNOR2_X1 U8190 ( .A(n13287), .B(n9821), .ZN(n13282) );
  NAND2_X1 U8191 ( .A1(n9538), .A2(n9537), .ZN(n9539) );
  NAND2_X1 U8192 ( .A1(n14954), .A2(n9458), .ZN(n13521) );
  AND2_X1 U8193 ( .A1(n13519), .A2(n13276), .ZN(n13529) );
  NOR2_X1 U8194 ( .A1(n9875), .A2(n9133), .ZN(n7218) );
  OAI22_X1 U8195 ( .A1(n6545), .A2(n9867), .B1(n10091), .B2(n14853), .ZN(n7217) );
  NAND2_X1 U8196 ( .A1(n9462), .A2(n9461), .ZN(n14953) );
  INV_X1 U8197 ( .A(n9799), .ZN(n13276) );
  NAND2_X1 U8198 ( .A1(n7889), .A2(n7888), .ZN(n14531) );
  INV_X1 U8199 ( .A(n14593), .ZN(n14488) );
  AND2_X1 U8200 ( .A1(n12313), .A2(n12312), .ZN(n6694) );
  OR2_X1 U8201 ( .A1(n7915), .A2(n7914), .ZN(n14497) );
  AND4_X1 U8202 ( .A1(n7861), .A2(n7860), .A3(n7859), .A4(n7858), .ZN(n11772)
         );
  INV_X1 U8203 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7498) );
  OAI21_X1 U8204 ( .B1(n13913), .B2(n13911), .A(n6873), .ZN(n6872) );
  AOI21_X1 U8205 ( .B1(n13912), .B2(n14649), .A(n14645), .ZN(n6873) );
  INV_X1 U8206 ( .A(n13911), .ZN(n14648) );
  OAI21_X1 U8207 ( .B1(n8917), .B2(n14107), .A(n8916), .ZN(n8918) );
  XNOR2_X1 U8208 ( .A(n8886), .B(n12301), .ZN(n6904) );
  NAND2_X1 U8209 ( .A1(n8002), .A2(n8001), .ZN(n13960) );
  NAND2_X1 U8210 ( .A1(n14150), .A2(n8107), .ZN(n13947) );
  NAND2_X1 U8211 ( .A1(n7934), .A2(n6594), .ZN(n7267) );
  NAND2_X1 U8212 ( .A1(n7719), .A2(n7266), .ZN(n7265) );
  XNOR2_X1 U8213 ( .A(n14284), .B(n14285), .ZN(n15347) );
  NOR2_X1 U8214 ( .A1(n14309), .A2(n14350), .ZN(n14355) );
  NAND2_X1 U8215 ( .A1(n6700), .A2(n6699), .ZN(n14585) );
  INV_X1 U8216 ( .A(n14319), .ZN(n6699) );
  INV_X1 U8217 ( .A(n14320), .ZN(n6700) );
  OAI21_X1 U8218 ( .B1(n14336), .B2(n14337), .A(n13254), .ZN(n6931) );
  AND2_X1 U8219 ( .A1(n12113), .A2(n7118), .ZN(n7117) );
  NAND2_X1 U8220 ( .A1(n7130), .A2(n12117), .ZN(n7129) );
  INV_X1 U8221 ( .A(n12128), .ZN(n7147) );
  OR2_X1 U8222 ( .A1(n7147), .A2(n12130), .ZN(n7146) );
  NAND2_X1 U8223 ( .A1(n7122), .A2(n12138), .ZN(n7121) );
  NAND2_X1 U8224 ( .A1(n12153), .A2(n12154), .ZN(n7166) );
  AOI21_X1 U8225 ( .B1(n9578), .B2(n9577), .A(n9576), .ZN(n9580) );
  INV_X1 U8226 ( .A(n7166), .ZN(n7165) );
  INV_X1 U8227 ( .A(n12161), .ZN(n7158) );
  AOI211_X1 U8228 ( .C1(n8728), .C2(n8727), .A(n15231), .B(n8726), .ZN(n8738)
         );
  INV_X1 U8229 ( .A(n9598), .ZN(n7450) );
  NOR2_X1 U8230 ( .A1(n9598), .A2(n9601), .ZN(n7451) );
  INV_X1 U8231 ( .A(n9620), .ZN(n7464) );
  INV_X1 U8232 ( .A(n9628), .ZN(n7466) );
  NOR2_X1 U8233 ( .A1(n12196), .A2(n12197), .ZN(n7152) );
  AOI21_X1 U8234 ( .B1(n12196), .B2(n12197), .A(n7154), .ZN(n7153) );
  INV_X1 U8235 ( .A(n12195), .ZN(n7154) );
  NOR2_X1 U8236 ( .A1(n9640), .A2(n6548), .ZN(n7475) );
  AOI21_X1 U8237 ( .B1(n6846), .B2(n6844), .A(n6553), .ZN(n6843) );
  INV_X1 U8238 ( .A(n6848), .ZN(n6844) );
  NAND2_X1 U8239 ( .A1(n7139), .A2(n12203), .ZN(n7138) );
  AOI22_X1 U8240 ( .A1(n7457), .A2(n7459), .B1(n7456), .B2(n7461), .ZN(n7452)
         );
  NAND2_X1 U8241 ( .A1(n7134), .A2(n12208), .ZN(n7133) );
  NAND2_X1 U8242 ( .A1(n7126), .A2(n12218), .ZN(n7125) );
  NOR2_X1 U8243 ( .A1(n6576), .A2(n6827), .ZN(n6826) );
  NAND2_X1 U8244 ( .A1(n6829), .A2(n6828), .ZN(n9710) );
  AOI21_X1 U8245 ( .B1(n6830), .B2(n7468), .A(n6562), .ZN(n6828) );
  AND2_X1 U8246 ( .A1(n9698), .A2(n9699), .ZN(n7468) );
  NAND2_X1 U8247 ( .A1(n6576), .A2(n6827), .ZN(n6825) );
  OAI21_X1 U8248 ( .B1(n7555), .B2(n7435), .A(n7559), .ZN(n7434) );
  INV_X1 U8249 ( .A(n7564), .ZN(n7430) );
  NAND2_X1 U8250 ( .A1(n7015), .A2(n7013), .ZN(n8855) );
  NOR2_X1 U8251 ( .A1(n8687), .A2(n7014), .ZN(n7013) );
  INV_X1 U8252 ( .A(n8675), .ZN(n7014) );
  INV_X1 U8253 ( .A(n8510), .ZN(n7025) );
  AND2_X1 U8254 ( .A1(n9519), .A2(n9520), .ZN(n7114) );
  INV_X1 U8255 ( .A(n9520), .ZN(n7111) );
  INV_X1 U8256 ( .A(n7403), .ZN(n7400) );
  NOR2_X1 U8257 ( .A1(n14025), .A2(n14032), .ZN(n7398) );
  NAND2_X1 U8258 ( .A1(n7056), .A2(n12189), .ZN(n7055) );
  INV_X1 U8259 ( .A(n7058), .ZN(n7056) );
  INV_X1 U8260 ( .A(n12189), .ZN(n7057) );
  NOR2_X1 U8261 ( .A1(n7998), .A2(n7978), .ZN(n7420) );
  INV_X1 U8262 ( .A(n7997), .ZN(n7419) );
  INV_X1 U8263 ( .A(n7998), .ZN(n7421) );
  NAND2_X1 U8264 ( .A1(n7547), .A2(n10422), .ZN(n7550) );
  NAND2_X1 U8265 ( .A1(n7538), .A2(SI_15_), .ZN(n7539) );
  INV_X1 U8266 ( .A(n7821), .ZN(n7424) );
  NAND2_X1 U8267 ( .A1(n14235), .A2(n14236), .ZN(n14237) );
  INV_X1 U8268 ( .A(n11326), .ZN(n7319) );
  OR2_X1 U8269 ( .A1(n12362), .A2(n12556), .ZN(n12360) );
  NAND2_X1 U8270 ( .A1(n6965), .A2(n6580), .ZN(n12569) );
  AND2_X1 U8271 ( .A1(n15179), .A2(n12663), .ZN(n6793) );
  AND2_X1 U8272 ( .A1(n6793), .A2(n8452), .ZN(n12664) );
  INV_X1 U8273 ( .A(n7361), .ZN(n7356) );
  AND2_X1 U8274 ( .A1(n7328), .A2(n8935), .ZN(n7327) );
  NAND2_X1 U8275 ( .A1(n8934), .A2(n7329), .ZN(n7328) );
  INV_X1 U8276 ( .A(n8933), .ZN(n7329) );
  INV_X1 U8277 ( .A(n8934), .ZN(n7330) );
  INV_X1 U8278 ( .A(n10964), .ZN(n11013) );
  OR2_X1 U8279 ( .A1(n12872), .A2(n8980), .ZN(n8852) );
  NOR2_X1 U8280 ( .A1(n12821), .A2(n7348), .ZN(n7347) );
  INV_X1 U8281 ( .A(n8953), .ZN(n7348) );
  OR2_X1 U8282 ( .A1(n14374), .A2(n12856), .ZN(n8785) );
  INV_X1 U8283 ( .A(n8513), .ZN(n7026) );
  AOI21_X1 U8284 ( .B1(n8513), .B2(n7025), .A(n7024), .ZN(n7023) );
  INV_X1 U8285 ( .A(n8528), .ZN(n7024) );
  INV_X1 U8286 ( .A(n7037), .ZN(n7036) );
  OAI21_X1 U8287 ( .B1(n8462), .B2(n7038), .A(n8491), .ZN(n7037) );
  INV_X1 U8288 ( .A(n8476), .ZN(n7038) );
  NAND2_X1 U8289 ( .A1(n9887), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8278) );
  INV_X1 U8290 ( .A(n10932), .ZN(n13044) );
  NAND2_X1 U8291 ( .A1(n9723), .A2(n6597), .ZN(n6821) );
  NOR2_X1 U8292 ( .A1(n9723), .A2(n6597), .ZN(n6822) );
  AND2_X1 U8293 ( .A1(n6779), .A2(n6778), .ZN(n13239) );
  NAND2_X1 U8294 ( .A1(n13238), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6778) );
  NAND2_X1 U8295 ( .A1(n7215), .A2(n13128), .ZN(n7214) );
  OR2_X1 U8296 ( .A1(n13557), .A2(n13118), .ZN(n9775) );
  INV_X1 U8297 ( .A(n6908), .ZN(n6907) );
  NAND2_X1 U8298 ( .A1(n9036), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n9378) );
  NAND2_X1 U8299 ( .A1(n6732), .A2(n6733), .ZN(n6731) );
  OR2_X1 U8300 ( .A1(n9290), .A2(n11567), .ZN(n9305) );
  INV_X1 U8301 ( .A(n9218), .ZN(n7203) );
  INV_X1 U8302 ( .A(n9178), .ZN(n7193) );
  NAND2_X1 U8303 ( .A1(n13401), .A2(n9542), .ZN(n13402) );
  INV_X1 U8304 ( .A(n9133), .ZN(n6744) );
  INV_X1 U8305 ( .A(n9898), .ZN(n6743) );
  NOR2_X1 U8306 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n6837) );
  OR2_X1 U8307 ( .A1(n9274), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n9297) );
  INV_X1 U8308 ( .A(n7609), .ZN(n7593) );
  INV_X1 U8309 ( .A(n7960), .ZN(n7971) );
  NAND2_X1 U8310 ( .A1(n7971), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n7970) );
  NAND2_X1 U8311 ( .A1(n11684), .A2(n7275), .ZN(n7274) );
  INV_X1 U8312 ( .A(n14484), .ZN(n7275) );
  NAND2_X1 U8313 ( .A1(n7171), .A2(n6603), .ZN(n7169) );
  INV_X1 U8314 ( .A(n13843), .ZN(n12335) );
  NOR2_X1 U8315 ( .A1(n14058), .A2(n6941), .ZN(n6940) );
  INV_X1 U8316 ( .A(n6942), .ZN(n6941) );
  INV_X1 U8317 ( .A(n7386), .ZN(n7383) );
  NOR2_X1 U8318 ( .A1(n14181), .A2(n14091), .ZN(n6942) );
  INV_X1 U8320 ( .A(n13852), .ZN(n11676) );
  NAND2_X1 U8321 ( .A1(n11902), .A2(n13860), .ZN(n12094) );
  NAND2_X1 U8322 ( .A1(n13940), .A2(n7087), .ZN(n7086) );
  INV_X1 U8323 ( .A(n7089), .ZN(n7087) );
  NAND2_X1 U8324 ( .A1(n13963), .A2(n7996), .ZN(n13949) );
  AOI21_X1 U8325 ( .B1(n7393), .B2(n7395), .A(n6616), .ZN(n7391) );
  AND2_X1 U8326 ( .A1(n9919), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9850) );
  INV_X1 U8327 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n7583) );
  INV_X1 U8328 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7575) );
  INV_X1 U8329 ( .A(n8127), .ZN(n7576) );
  INV_X1 U8330 ( .A(P2_RD_REG_SCAN_IN), .ZN(n6850) );
  INV_X1 U8331 ( .A(P1_RD_REG_SCAN_IN), .ZN(n6852) );
  INV_X1 U8332 ( .A(n7918), .ZN(n7446) );
  INV_X1 U8333 ( .A(n6896), .ZN(n6895) );
  OAI21_X1 U8334 ( .B1(n7440), .B2(n6897), .A(n7543), .ZN(n6896) );
  INV_X1 U8335 ( .A(n7882), .ZN(n6897) );
  NAND2_X1 U8336 ( .A1(n7442), .A2(n7535), .ZN(n7862) );
  XNOR2_X1 U8337 ( .A(n7531), .B(SI_12_), .ZN(n7821) );
  AOI21_X1 U8338 ( .B1(n7527), .B2(n7427), .A(n6627), .ZN(n7425) );
  INV_X1 U8339 ( .A(n7427), .ZN(n7426) );
  NAND2_X1 U8340 ( .A1(n7523), .A2(SI_9_), .ZN(n7525) );
  INV_X1 U8341 ( .A(n7508), .ZN(n6866) );
  INV_X1 U8342 ( .A(n7510), .ZN(n6891) );
  OAI21_X1 U8343 ( .B1(n9854), .B2(n9868), .A(n6775), .ZN(n7409) );
  NAND2_X1 U8344 ( .A1(n9854), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6775) );
  NAND2_X1 U8345 ( .A1(n7409), .A2(SI_3_), .ZN(n7508) );
  NAND2_X1 U8346 ( .A1(n7503), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6714) );
  OAI21_X1 U8347 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n14249), .A(n14248), .ZN(
        n14274) );
  AOI21_X1 U8348 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n14251), .A(n14250), .ZN(
        n14252) );
  NOR2_X1 U8349 ( .A1(n14274), .A2(n14273), .ZN(n14250) );
  AOI21_X1 U8350 ( .B1(n12435), .B2(n12400), .A(n12403), .ZN(n7311) );
  INV_X1 U8351 ( .A(n7311), .ZN(n7308) );
  AND2_X1 U8352 ( .A1(n7284), .A2(n6637), .ZN(n7283) );
  NAND2_X1 U8353 ( .A1(n12504), .A2(n7287), .ZN(n7284) );
  NAND2_X1 U8354 ( .A1(n7282), .A2(n6572), .ZN(n7281) );
  AND2_X1 U8355 ( .A1(n8394), .A2(n8393), .ZN(n11724) );
  AND2_X1 U8356 ( .A1(n12398), .A2(n12396), .ZN(n12465) );
  NAND2_X1 U8357 ( .A1(n8470), .A2(n8469), .ZN(n8483) );
  NAND2_X1 U8358 ( .A1(n12392), .A2(n12492), .ZN(n12494) );
  AND2_X1 U8359 ( .A1(n8309), .A2(n8308), .ZN(n8328) );
  AND4_X1 U8360 ( .A1(n8629), .A2(n8628), .A3(n8627), .A4(n8626), .ZN(n12406)
         );
  AND4_X1 U8361 ( .A1(n8614), .A2(n8613), .A3(n8612), .A4(n8611), .ZN(n8966)
         );
  AND4_X1 U8362 ( .A1(n8475), .A2(n8474), .A3(n8473), .A4(n8472), .ZN(n12485)
         );
  NAND2_X1 U8363 ( .A1(n10426), .A2(n6465), .ZN(n6794) );
  NAND2_X1 U8364 ( .A1(n6800), .A2(n6798), .ZN(n15011) );
  INV_X1 U8365 ( .A(n6799), .ZN(n6798) );
  OAI22_X1 U8366 ( .A1(n12628), .A2(n6804), .B1(n12626), .B2(n12627), .ZN(
        n6799) );
  NAND2_X1 U8367 ( .A1(n15006), .A2(n6968), .ZN(n6967) );
  INV_X1 U8368 ( .A(n6805), .ZN(n15105) );
  INV_X1 U8369 ( .A(n15081), .ZN(n6807) );
  OAI21_X1 U8370 ( .B1(n15081), .B2(n12639), .A(n6660), .ZN(n6806) );
  NOR2_X1 U8371 ( .A1(n15092), .A2(n6708), .ZN(n12574) );
  AND2_X1 U8372 ( .A1(n15100), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6708) );
  NAND2_X1 U8373 ( .A1(n14389), .A2(n6959), .ZN(n6958) );
  NAND2_X1 U8374 ( .A1(n6792), .A2(n6790), .ZN(n14393) );
  NAND2_X1 U8375 ( .A1(n6791), .A2(n14389), .ZN(n6790) );
  INV_X1 U8376 ( .A(n12664), .ZN(n6792) );
  INV_X1 U8377 ( .A(n6793), .ZN(n6791) );
  NOR2_X1 U8378 ( .A1(n14393), .A2(n14394), .ZN(n14392) );
  OR2_X1 U8379 ( .A1(n14411), .A2(n6673), .ZN(n6961) );
  NAND2_X1 U8380 ( .A1(n14411), .A2(n12666), .ZN(n6960) );
  NAND2_X1 U8381 ( .A1(n6668), .A2(n12666), .ZN(n6962) );
  INV_X1 U8382 ( .A(n8969), .ZN(n12716) );
  INV_X1 U8383 ( .A(n8609), .ZN(n8610) );
  NAND2_X1 U8384 ( .A1(n8965), .A2(n8964), .ZN(n12725) );
  INV_X1 U8385 ( .A(n8596), .ZN(n8597) );
  NOR2_X1 U8386 ( .A1(n8597), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8609) );
  INV_X1 U8387 ( .A(n8584), .ZN(n8585) );
  INV_X1 U8388 ( .A(n8570), .ZN(n8571) );
  NOR2_X1 U8389 ( .A1(n8571), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8584) );
  NOR2_X1 U8390 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(n7478), .ZN(n8570) );
  NAND2_X1 U8391 ( .A1(n8536), .A2(n8535), .ZN(n8546) );
  AOI21_X1 U8392 ( .B1(n7010), .B2(n7009), .A(n7008), .ZN(n7007) );
  INV_X1 U8393 ( .A(n8365), .ZN(n7009) );
  INV_X1 U8394 ( .A(n8773), .ZN(n7008) );
  OR2_X1 U8395 ( .A1(n8367), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8395) );
  INV_X1 U8396 ( .A(n11641), .ZN(n14455) );
  NAND2_X1 U8397 ( .A1(n11396), .A2(n8933), .ZN(n7326) );
  NAND2_X1 U8398 ( .A1(n8756), .A2(n8757), .ZN(n11386) );
  NOR2_X1 U8399 ( .A1(n8285), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8309) );
  OR2_X1 U8400 ( .A1(n8532), .A2(n8299), .ZN(n8306) );
  OR2_X1 U8401 ( .A1(n8267), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8285) );
  NOR2_X1 U8402 ( .A1(n15187), .A2(n7351), .ZN(n7350) );
  INV_X1 U8403 ( .A(n8930), .ZN(n7351) );
  AND3_X1 U8404 ( .A1(n8283), .A2(n8282), .A3(n8281), .ZN(n15196) );
  INV_X1 U8405 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n10975) );
  NOR2_X1 U8406 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8250) );
  NAND2_X1 U8407 ( .A1(n6984), .A2(n8190), .ZN(n15235) );
  OR2_X1 U8408 ( .A1(n9021), .A2(n9020), .ZN(n15266) );
  NAND2_X1 U8409 ( .A1(n7015), .A2(n8675), .ZN(n12681) );
  AOI21_X1 U8410 ( .B1(n6583), .B2(n6993), .A(n6989), .ZN(n6988) );
  INV_X1 U8411 ( .A(n8819), .ZN(n6993) );
  NAND2_X1 U8412 ( .A1(n12760), .A2(n12761), .ZN(n12746) );
  AOI21_X1 U8413 ( .B1(n7334), .B2(n7336), .A(n6581), .ZN(n7332) );
  NAND2_X1 U8414 ( .A1(n12832), .A2(n8952), .ZN(n7349) );
  AOI21_X1 U8415 ( .B1(n6998), .B2(n6997), .A(n8946), .ZN(n6996) );
  NAND2_X1 U8416 ( .A1(n6680), .A2(n6998), .ZN(n6994) );
  INV_X1 U8417 ( .A(n8949), .ZN(n12843) );
  AND2_X1 U8418 ( .A1(n8978), .A2(n8977), .ZN(n15259) );
  INV_X1 U8419 ( .A(n15243), .ZN(n15256) );
  INV_X1 U8420 ( .A(n15253), .ZN(n12888) );
  AND2_X1 U8421 ( .A1(n8168), .A2(n7364), .ZN(n7363) );
  AND2_X1 U8422 ( .A1(n7366), .A2(n8161), .ZN(n7364) );
  INV_X1 U8423 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8871) );
  INV_X1 U8424 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8864) );
  NAND2_X1 U8425 ( .A1(n8717), .A2(n6607), .ZN(n8870) );
  NAND2_X1 U8426 ( .A1(n8542), .A2(n8541), .ZN(n8555) );
  INV_X1 U8427 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n6817) );
  NOR2_X1 U8428 ( .A1(n8160), .A2(n8374), .ZN(n8391) );
  AOI21_X1 U8429 ( .B1(n7030), .B2(n7032), .A(n7029), .ZN(n7028) );
  INV_X1 U8430 ( .A(n8385), .ZN(n7029) );
  AND2_X1 U8431 ( .A1(n8401), .A2(n8387), .ZN(n8388) );
  AOI21_X1 U8432 ( .B1(n7044), .B2(n7042), .A(n7041), .ZN(n7040) );
  INV_X1 U8433 ( .A(n7044), .ZN(n7043) );
  INV_X1 U8434 ( .A(n8334), .ZN(n7041) );
  AND2_X1 U8435 ( .A1(n8352), .A2(n8336), .ZN(n8337) );
  OR2_X1 U8436 ( .A1(n8340), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8359) );
  OAI21_X1 U8437 ( .B1(n8240), .B2(n7018), .A(n7017), .ZN(n7019) );
  INV_X1 U8438 ( .A(n8241), .ZN(n7018) );
  AOI21_X1 U8439 ( .B1(n8238), .B2(n8241), .A(n8257), .ZN(n7017) );
  OR2_X1 U8440 ( .A1(n8243), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n8261) );
  INV_X1 U8441 ( .A(n10435), .ZN(n6789) );
  OR2_X1 U8442 ( .A1(n13058), .A2(n13057), .ZN(n13059) );
  XNOR2_X1 U8443 ( .A(n10932), .B(n11166), .ZN(n10934) );
  NOR2_X1 U8444 ( .A1(n9193), .A2(n9033), .ZN(n9210) );
  INV_X1 U8445 ( .A(n9359), .ZN(n9035) );
  OR2_X1 U8446 ( .A1(n9366), .A2(n13107), .ZN(n9368) );
  AND2_X1 U8447 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n9171) );
  NAND2_X1 U8448 ( .A1(n9266), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9278) );
  OR2_X1 U8449 ( .A1(n9278), .A2(n14820), .ZN(n9290) );
  INV_X1 U8450 ( .A(n14826), .ZN(n7219) );
  NAND2_X1 U8451 ( .A1(n13035), .A2(n6706), .ZN(n6705) );
  INV_X1 U8452 ( .A(n13036), .ZN(n6706) );
  NOR2_X1 U8453 ( .A1(n9235), .A2(n14905), .ZN(n9251) );
  XNOR2_X1 U8454 ( .A(n10932), .B(n11131), .ZN(n11155) );
  INV_X1 U8455 ( .A(n10956), .ZN(n10953) );
  AND2_X1 U8456 ( .A1(n6783), .A2(n6782), .ZN(n14880) );
  NAND2_X1 U8457 ( .A1(n10102), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6782) );
  AND2_X1 U8458 ( .A1(n13257), .A2(n13256), .ZN(n13270) );
  NAND2_X1 U8459 ( .A1(n13288), .A2(n13641), .ZN(n13287) );
  INV_X1 U8460 ( .A(n9794), .ZN(n9527) );
  XNOR2_X1 U8461 ( .A(n13317), .B(n9525), .ZN(n13308) );
  INV_X1 U8462 ( .A(n6765), .ZN(n13309) );
  OAI21_X1 U8463 ( .B1(n13336), .B2(n6767), .A(n6766), .ZN(n6765) );
  NAND2_X1 U8464 ( .A1(n13557), .A2(n13184), .ZN(n6766) );
  NOR2_X1 U8465 ( .A1(n13557), .A2(n13184), .ZN(n6767) );
  AND2_X1 U8466 ( .A1(n9040), .A2(n9401), .ZN(n13331) );
  NAND2_X1 U8467 ( .A1(n6768), .A2(n7207), .ZN(n13336) );
  INV_X1 U8468 ( .A(n7208), .ZN(n7207) );
  NAND2_X1 U8469 ( .A1(n13356), .A2(n7206), .ZN(n6768) );
  OAI21_X1 U8470 ( .B1(n7210), .B2(n7212), .A(n7214), .ZN(n7208) );
  AOI21_X1 U8471 ( .B1(n7103), .B2(n7105), .A(n6595), .ZN(n7101) );
  NAND2_X1 U8472 ( .A1(n13401), .A2(n6908), .ZN(n13387) );
  NAND2_X1 U8473 ( .A1(n6758), .A2(n6755), .ZN(n13386) );
  NAND2_X1 U8474 ( .A1(n6757), .A2(n6756), .ZN(n6755) );
  NOR2_X1 U8475 ( .A1(n7178), .A2(n6760), .ZN(n6759) );
  INV_X1 U8476 ( .A(n9790), .ZN(n13420) );
  OR2_X1 U8477 ( .A1(n9334), .A2(n12070), .ZN(n9345) );
  NAND2_X1 U8478 ( .A1(n9034), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9357) );
  INV_X1 U8479 ( .A(n9345), .ZN(n9034) );
  INV_X1 U8480 ( .A(n7196), .ZN(n6773) );
  NAND2_X1 U8481 ( .A1(n7196), .A2(n7197), .ZN(n7195) );
  INV_X1 U8482 ( .A(n13135), .ZN(n13172) );
  INV_X1 U8483 ( .A(n13136), .ZN(n13173) );
  NAND2_X1 U8484 ( .A1(n6722), .A2(n7108), .ZN(n11664) );
  AOI21_X1 U8485 ( .B1(n11604), .B2(n7109), .A(n6560), .ZN(n7108) );
  NAND2_X1 U8486 ( .A1(n11603), .A2(n7109), .ZN(n6722) );
  NAND2_X1 U8487 ( .A1(n11599), .A2(n11738), .ZN(n11667) );
  INV_X1 U8488 ( .A(n9783), .ZN(n11344) );
  AND2_X1 U8489 ( .A1(n9492), .A2(n6774), .ZN(n11283) );
  INV_X1 U8490 ( .A(n11283), .ZN(n11288) );
  XNOR2_X1 U8491 ( .A(n13205), .B(n11223), .ZN(n10533) );
  XNOR2_X1 U8492 ( .A(n13206), .B(n9145), .ZN(n10554) );
  XNOR2_X1 U8493 ( .A(n13207), .B(n6909), .ZN(n10564) );
  NAND2_X1 U8494 ( .A1(n6910), .A2(n6909), .ZN(n10562) );
  OR2_X1 U8495 ( .A1(n13549), .A2(n13622), .ZN(n6753) );
  AND2_X1 U8496 ( .A1(n13330), .A2(n13329), .ZN(n13556) );
  CLKBUF_X1 U8497 ( .A(n10406), .Z(n14986) );
  AND3_X1 U8498 ( .A1(n6742), .A2(n6741), .A3(n6740), .ZN(n9145) );
  OR2_X1 U8499 ( .A1(n9142), .A2(n10100), .ZN(n6740) );
  OR2_X1 U8500 ( .A1(n6545), .A2(n9868), .ZN(n6741) );
  NAND2_X1 U8501 ( .A1(n6744), .A2(n6743), .ZN(n6742) );
  NAND2_X1 U8502 ( .A1(n7245), .A2(n9456), .ZN(n7244) );
  INV_X1 U8503 ( .A(n7247), .ZN(n7245) );
  XNOR2_X1 U8504 ( .A(n9352), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9799) );
  NAND2_X1 U8505 ( .A1(n9430), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9352) );
  OR2_X1 U8506 ( .A1(n9132), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n9157) );
  INV_X1 U8507 ( .A(n7970), .ZN(n7610) );
  NAND2_X1 U8508 ( .A1(n7610), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n7609) );
  AOI21_X1 U8509 ( .B1(n12046), .B2(n12044), .A(n12329), .ZN(n7260) );
  INV_X1 U8510 ( .A(n7260), .ZN(n7258) );
  INV_X1 U8511 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7758) );
  NAND2_X1 U8512 ( .A1(n10989), .A2(n6605), .ZN(n11440) );
  INV_X1 U8513 ( .A(n10992), .ZN(n6868) );
  NOR2_X1 U8514 ( .A1(n7873), .A2(n7872), .ZN(n7890) );
  NAND2_X1 U8515 ( .A1(n6858), .A2(n6861), .ZN(n13768) );
  NAND2_X1 U8516 ( .A1(n6676), .A2(n11961), .ZN(n6858) );
  AND2_X1 U8517 ( .A1(n7940), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n7948) );
  NAND2_X1 U8518 ( .A1(n11961), .A2(n13759), .ZN(n6863) );
  NOR2_X1 U8519 ( .A1(n7253), .A2(n7250), .ZN(n7249) );
  INV_X1 U8520 ( .A(n11970), .ZN(n7250) );
  INV_X1 U8521 ( .A(n7491), .ZN(n7253) );
  NAND2_X1 U8522 ( .A1(n6861), .A2(n13770), .ZN(n6860) );
  INV_X1 U8523 ( .A(n7251), .ZN(n6856) );
  AOI21_X1 U8524 ( .B1(n7491), .B2(n7252), .A(n6628), .ZN(n7251) );
  INV_X1 U8525 ( .A(n13807), .ZN(n7252) );
  OR2_X1 U8526 ( .A1(n7842), .A2(n7841), .ZN(n7856) );
  AND2_X1 U8527 ( .A1(n7812), .A2(n7592), .ZN(n7826) );
  INV_X1 U8528 ( .A(n7273), .ZN(n7271) );
  NAND2_X1 U8529 ( .A1(n14484), .A2(n14483), .ZN(n7273) );
  NAND2_X1 U8530 ( .A1(n14482), .A2(n7274), .ZN(n7272) );
  OR2_X1 U8531 ( .A1(n6470), .A2(n11902), .ZN(n10169) );
  OR2_X1 U8532 ( .A1(n7910), .A2(n11881), .ZN(n7928) );
  NOR2_X1 U8533 ( .A1(n7928), .A2(n7927), .ZN(n7940) );
  NAND2_X1 U8534 ( .A1(n13768), .A2(n11970), .ZN(n13808) );
  NAND2_X1 U8535 ( .A1(n13808), .A2(n13807), .ZN(n13806) );
  NAND2_X1 U8536 ( .A1(n8114), .A2(n14227), .ZN(n12264) );
  INV_X1 U8537 ( .A(n13831), .ZN(n7262) );
  INV_X1 U8538 ( .A(n11954), .ZN(n7264) );
  INV_X1 U8539 ( .A(n12264), .ZN(n9920) );
  OR2_X1 U8540 ( .A1(n7642), .A2(n7616), .ZN(n7617) );
  AOI21_X1 U8541 ( .B1(n14628), .B2(n14629), .A(n6885), .ZN(n14626) );
  NOR2_X1 U8542 ( .A1(n14626), .A2(n6883), .ZN(n10004) );
  NOR2_X1 U8543 ( .A1(n6884), .A2(n14801), .ZN(n6883) );
  NOR2_X1 U8544 ( .A1(n10035), .A2(n6881), .ZN(n10039) );
  AND2_X1 U8545 ( .A1(n10036), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6881) );
  NAND2_X1 U8546 ( .A1(n10039), .A2(n10038), .ZN(n10197) );
  NOR2_X1 U8547 ( .A1(n11374), .A2(n6887), .ZN(n11376) );
  AND2_X1 U8548 ( .A1(n11375), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6887) );
  NAND2_X1 U8549 ( .A1(n11376), .A2(n11377), .ZN(n11780) );
  INV_X1 U8550 ( .A(n7806), .ZN(n7373) );
  NAND2_X1 U8551 ( .A1(n11780), .A2(n6886), .ZN(n11782) );
  OR2_X1 U8552 ( .A1(n11781), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6886) );
  NAND2_X1 U8553 ( .A1(n6880), .A2(n6879), .ZN(n6878) );
  NAND2_X1 U8554 ( .A1(n13890), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6879) );
  AND2_X1 U8555 ( .A1(n6878), .A2(n13903), .ZN(n13908) );
  INV_X1 U8556 ( .A(n12231), .ZN(n12232) );
  AND2_X1 U8557 ( .A1(n12294), .A2(n8106), .ZN(n7083) );
  AND2_X1 U8558 ( .A1(n7948), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n7959) );
  NAND2_X1 U8559 ( .A1(n7959), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n7960) );
  AND2_X1 U8560 ( .A1(n14049), .A2(n7954), .ZN(n14031) );
  NAND2_X1 U8561 ( .A1(n6566), .A2(n14056), .ZN(n14049) );
  NAND2_X1 U8562 ( .A1(n14099), .A2(n14188), .ZN(n14087) );
  OAI21_X1 U8563 ( .B1(n14096), .B2(n7917), .A(n7916), .ZN(n14080) );
  AOI21_X1 U8564 ( .B1(n7076), .B2(n7078), .A(n6612), .ZN(n7075) );
  INV_X1 U8565 ( .A(n7276), .ZN(n8111) );
  NAND2_X1 U8567 ( .A1(n11847), .A2(n12159), .ZN(n14493) );
  NAND2_X1 U8568 ( .A1(n11849), .A2(n11848), .ZN(n11847) );
  NAND2_X1 U8569 ( .A1(n11843), .A2(n13832), .ZN(n14505) );
  NAND2_X1 U8570 ( .A1(n6943), .A2(n14552), .ZN(n14125) );
  INV_X1 U8571 ( .A(n6943), .ZN(n11653) );
  AOI21_X1 U8572 ( .B1(n7063), .B2(n7065), .A(n6613), .ZN(n7061) );
  NAND2_X1 U8573 ( .A1(n7370), .A2(n7802), .ZN(n11533) );
  INV_X1 U8574 ( .A(n12279), .ZN(n14674) );
  NOR2_X1 U8575 ( .A1(n14749), .A2(n14697), .ZN(n7066) );
  INV_X1 U8576 ( .A(n7068), .ZN(n7067) );
  OAI21_X1 U8577 ( .B1(n12110), .B2(n14598), .A(n8078), .ZN(n7068) );
  NAND2_X1 U8578 ( .A1(n7678), .A2(n7677), .ZN(n11076) );
  AND2_X1 U8579 ( .A1(n6898), .A2(n6554), .ZN(n13964) );
  INV_X1 U8580 ( .A(n14521), .ZN(n14558) );
  NAND2_X1 U8581 ( .A1(n10061), .A2(n8905), .ZN(n14761) );
  INV_X1 U8582 ( .A(n14792), .ZN(n14726) );
  INV_X1 U8583 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7587) );
  AND2_X1 U8584 ( .A1(n8882), .A2(n8040), .ZN(n8880) );
  XNOR2_X1 U8585 ( .A(n8035), .B(n8019), .ZN(n13699) );
  OAI21_X1 U8586 ( .B1(n7977), .B2(n7422), .A(n7980), .ZN(n7999) );
  NAND2_X1 U8587 ( .A1(n8125), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8126) );
  XNOR2_X1 U8588 ( .A(n7977), .B(n7978), .ZN(n11859) );
  NAND2_X1 U8589 ( .A1(n8059), .A2(n8121), .ZN(n7116) );
  MUX2_X1 U8590 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8058), .S(
        P1_IR_REG_22__SCAN_IN), .Z(n8059) );
  NAND2_X1 U8591 ( .A1(n7923), .A2(n7922), .ZN(n7934) );
  INV_X1 U8592 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7922) );
  NAND2_X1 U8593 ( .A1(n7439), .A2(n7440), .ZN(n7883) );
  XNOR2_X1 U8594 ( .A(n7805), .B(n7804), .ZN(n10045) );
  AOI21_X1 U8595 ( .B1(n7413), .B2(n7415), .A(n7411), .ZN(n7410) );
  INV_X1 U8596 ( .A(n7522), .ZN(n7411) );
  OR2_X1 U8597 ( .A1(n7772), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n7773) );
  NAND2_X1 U8598 ( .A1(n7702), .A2(n7513), .ZN(n6764) );
  AND2_X1 U8599 ( .A1(n7905), .A2(n7704), .ZN(n7737) );
  OAI21_X1 U8600 ( .B1(SI_3_), .B2(n7409), .A(n7508), .ZN(n7669) );
  INV_X1 U8601 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n7565) );
  INV_X1 U8602 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n14283) );
  NAND2_X1 U8603 ( .A1(n14231), .A2(n6926), .ZN(n14279) );
  NAND2_X1 U8604 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n6927), .ZN(n6926) );
  INV_X1 U8605 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6927) );
  NAND2_X1 U8606 ( .A1(n14242), .A2(n14241), .ZN(n14296) );
  NOR2_X1 U8607 ( .A1(n14345), .A2(n14297), .ZN(n14299) );
  NAND2_X1 U8608 ( .A1(n14348), .A2(n14306), .ZN(n14308) );
  NOR2_X1 U8609 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14252), .ZN(n14310) );
  NOR2_X1 U8610 ( .A1(n14310), .A2(n14253), .ZN(n14272) );
  AND2_X1 U8611 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(n14312), .ZN(n14253) );
  AOI21_X1 U8612 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n14257), .A(n14256), .ZN(
        n14315) );
  OR2_X1 U8613 ( .A1(n10642), .A2(n10621), .ZN(n12533) );
  INV_X1 U8614 ( .A(n7313), .ZN(n7312) );
  NAND2_X1 U8615 ( .A1(n7314), .A2(n12491), .ZN(n12443) );
  INV_X1 U8616 ( .A(n11410), .ZN(n7320) );
  NAND2_X1 U8617 ( .A1(n12435), .A2(n12404), .ZN(n7310) );
  NAND2_X1 U8618 ( .A1(n6717), .A2(n7301), .ZN(n7295) );
  NAND2_X1 U8619 ( .A1(n7292), .A2(n7293), .ZN(n12483) );
  OR2_X1 U8620 ( .A1(n6717), .A2(n7294), .ZN(n7292) );
  AND2_X1 U8621 ( .A1(n11322), .A2(n7481), .ZN(n11323) );
  OR2_X1 U8622 ( .A1(n11321), .A2(n11452), .ZN(n7481) );
  INV_X1 U8623 ( .A(n7321), .ZN(n11411) );
  NAND2_X1 U8624 ( .A1(n7289), .A2(n7288), .ZN(n12521) );
  AOI21_X1 U8625 ( .B1(n7290), .B2(n7294), .A(n6623), .ZN(n7288) );
  NAND2_X1 U8626 ( .A1(n10645), .A2(n10644), .ZN(n14376) );
  AOI21_X1 U8627 ( .B1(n6717), .B2(n14368), .A(n6569), .ZN(n12541) );
  INV_X1 U8628 ( .A(n14376), .ZN(n12550) );
  NAND2_X1 U8629 ( .A1(n7005), .A2(n7004), .ZN(n7003) );
  AND4_X1 U8630 ( .A1(n8683), .A2(n8682), .A3(n8681), .A4(n8680), .ZN(n11149)
         );
  AND4_X1 U8631 ( .A1(n8683), .A2(n8654), .A3(n8653), .A4(n8652), .ZN(n12405)
         );
  INV_X1 U8632 ( .A(n12406), .ZN(n12552) );
  INV_X1 U8633 ( .A(n8966), .ZN(n12739) );
  INV_X1 U8634 ( .A(n12807), .ZN(n12833) );
  OR2_X1 U8635 ( .A1(n6477), .A2(n11618), .ZN(n8396) );
  NAND4_X1 U8636 ( .A1(n8351), .A2(n8350), .A3(n8349), .A4(n8348), .ZN(n12559)
         );
  NAND4_X1 U8637 ( .A1(n8333), .A2(n8332), .A3(n8331), .A4(n8330), .ZN(n12560)
         );
  INV_X1 U8638 ( .A(n11452), .ZN(n12561) );
  INV_X1 U8639 ( .A(P3_U3897), .ZN(n12563) );
  NAND2_X1 U8640 ( .A1(n6951), .A2(n10486), .ZN(n10439) );
  INV_X1 U8641 ( .A(n6804), .ZN(n6797) );
  INV_X1 U8642 ( .A(n6687), .ZN(n15067) );
  NOR2_X1 U8643 ( .A1(n15080), .A2(n15081), .ZN(n15079) );
  NOR2_X1 U8644 ( .A1(n15062), .A2(n12642), .ZN(n15080) );
  NOR2_X1 U8645 ( .A1(n15094), .A2(n15093), .ZN(n15092) );
  XNOR2_X1 U8646 ( .A(n12574), .B(n12650), .ZN(n15111) );
  NOR2_X1 U8647 ( .A1(n15111), .A2(n8366), .ZN(n15110) );
  AND2_X1 U8648 ( .A1(n15120), .A2(n12652), .ZN(n15140) );
  NAND2_X1 U8649 ( .A1(n15138), .A2(n12655), .ZN(n15156) );
  NOR2_X1 U8650 ( .A1(n15144), .A2(n12578), .ZN(n15165) );
  INV_X1 U8651 ( .A(n6964), .ZN(n12577) );
  AND2_X1 U8652 ( .A1(n15154), .A2(n12659), .ZN(n15181) );
  NAND2_X1 U8653 ( .A1(n8650), .A2(n8649), .ZN(n12694) );
  AND2_X1 U8654 ( .A1(n12685), .A2(n8640), .ZN(n12701) );
  NAND2_X1 U8655 ( .A1(n12766), .A2(n8962), .ZN(n12755) );
  NAND2_X1 U8656 ( .A1(n7360), .A2(n7358), .ZN(n11613) );
  NAND2_X1 U8657 ( .A1(n10508), .A2(n10619), .ZN(n15268) );
  AND2_X1 U8658 ( .A1(n15227), .A2(n12888), .ZN(n12860) );
  INV_X1 U8659 ( .A(n15268), .ZN(n15226) );
  OAI21_X1 U8660 ( .B1(n7369), .B2(n15329), .A(n6663), .ZN(n7368) );
  INV_X1 U8661 ( .A(n12681), .ZN(n12924) );
  NAND2_X1 U8662 ( .A1(n8660), .A2(n8659), .ZN(n12925) );
  NAND2_X1 U8663 ( .A1(n8568), .A2(n8567), .ZN(n12954) );
  NAND2_X1 U8664 ( .A1(n8559), .A2(n8558), .ZN(n12960) );
  NAND2_X1 U8665 ( .A1(n6990), .A2(n8819), .ZN(n12773) );
  NAND2_X1 U8666 ( .A1(n12783), .A2(n8820), .ZN(n6990) );
  NAND2_X1 U8667 ( .A1(n7333), .A2(n8957), .ZN(n12784) );
  NAND2_X1 U8668 ( .A1(n12795), .A2(n8956), .ZN(n7333) );
  NAND2_X1 U8669 ( .A1(n8534), .A2(n8533), .ZN(n12972) );
  OR2_X1 U8670 ( .A1(n10753), .A2(n8532), .ZN(n8534) );
  NAND2_X1 U8671 ( .A1(n6974), .A2(n6978), .ZN(n12793) );
  OR2_X1 U8672 ( .A1(n12822), .A2(n6979), .ZN(n6974) );
  NAND2_X1 U8673 ( .A1(n6981), .A2(n8803), .ZN(n12813) );
  OR2_X1 U8674 ( .A1(n12822), .A2(n12823), .ZN(n6981) );
  NAND2_X1 U8675 ( .A1(n8500), .A2(n8499), .ZN(n12986) );
  NAND2_X1 U8676 ( .A1(n8467), .A2(n8466), .ZN(n12998) );
  OR2_X1 U8677 ( .A1(n10054), .A2(n8532), .ZN(n8467) );
  NAND2_X1 U8678 ( .A1(n6995), .A2(n6998), .ZN(n12852) );
  NAND2_X1 U8679 ( .A1(n11829), .A2(n7000), .ZN(n6995) );
  INV_X1 U8680 ( .A(n12983), .ZN(n13005) );
  NAND2_X1 U8681 ( .A1(n7002), .A2(n7000), .ZN(n11867) );
  OR2_X1 U8682 ( .A1(n11829), .A2(n8782), .ZN(n7002) );
  INV_X2 U8683 ( .A(n15316), .ZN(n15318) );
  XNOR2_X1 U8684 ( .A(n8672), .B(n8671), .ZN(n13010) );
  BUF_X1 U8685 ( .A(n8172), .Z(n12416) );
  NAND2_X1 U8686 ( .A1(n7046), .A2(n8632), .ZN(n8646) );
  NAND2_X1 U8687 ( .A1(n8717), .A2(n8168), .ZN(n8866) );
  XNOR2_X1 U8688 ( .A(n8872), .B(n8871), .ZN(n11593) );
  OAI21_X1 U8689 ( .B1(n8870), .B2(P3_IR_REG_24__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8872) );
  NAND2_X1 U8690 ( .A1(n8514), .A2(n8513), .ZN(n8529) );
  NAND2_X1 U8691 ( .A1(n8511), .A2(n8510), .ZN(n8514) );
  NAND2_X1 U8692 ( .A1(n8477), .A2(n8476), .ZN(n8492) );
  OAI21_X1 U8693 ( .B1(n8424), .B2(n7022), .A(n7020), .ZN(n8447) );
  NAND2_X1 U8694 ( .A1(n8427), .A2(n8426), .ZN(n8444) );
  NAND2_X1 U8695 ( .A1(n8424), .A2(n8423), .ZN(n8427) );
  OAI21_X1 U8696 ( .B1(n8356), .B2(n7032), .A(n7030), .ZN(n8386) );
  NAND2_X1 U8697 ( .A1(n8378), .A2(n8377), .ZN(n8381) );
  NAND2_X1 U8698 ( .A1(n7039), .A2(n7044), .ZN(n8335) );
  NAND2_X1 U8699 ( .A1(n8297), .A2(n8316), .ZN(n7039) );
  NAND2_X1 U8700 ( .A1(n7016), .A2(n8241), .ZN(n8258) );
  NAND2_X1 U8701 ( .A1(n8240), .A2(n8239), .ZN(n7016) );
  NAND2_X1 U8702 ( .A1(n11263), .A2(n11059), .ZN(n12422) );
  INV_X1 U8703 ( .A(n7222), .ZN(n7221) );
  NAND2_X1 U8704 ( .A1(n11807), .A2(n11806), .ZN(n11808) );
  NOR2_X1 U8705 ( .A1(n6570), .A2(n7232), .ZN(n7231) );
  OAI21_X1 U8706 ( .B1(n7233), .B2(n6570), .A(n12075), .ZN(n7230) );
  AND3_X1 U8707 ( .A1(n11806), .A2(n7233), .A3(n11807), .ZN(n12077) );
  NAND2_X1 U8708 ( .A1(n13042), .A2(n7226), .ZN(n7228) );
  AND2_X1 U8709 ( .A1(n10404), .A2(n13521), .ZN(n13133) );
  OR2_X1 U8710 ( .A1(n13086), .A2(n13031), .ZN(n7238) );
  NAND2_X1 U8711 ( .A1(n12422), .A2(n11265), .ZN(n12432) );
  NAND2_X1 U8712 ( .A1(n9344), .A2(n9343), .ZN(n13601) );
  NAND2_X1 U8713 ( .A1(n12359), .A2(n10952), .ZN(n10955) );
  NAND2_X1 U8714 ( .A1(n10919), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14832) );
  INV_X1 U8715 ( .A(n13159), .ZN(n14822) );
  NAND2_X1 U8716 ( .A1(n6716), .A2(n7485), .ZN(n11807) );
  CLKBUF_X1 U8717 ( .A(n11714), .Z(n6716) );
  NOR2_X1 U8718 ( .A1(n14824), .A2(n11269), .ZN(n13167) );
  AND2_X1 U8719 ( .A1(n10415), .A2(n10412), .ZN(n13148) );
  INV_X1 U8720 ( .A(n12065), .ZN(n9843) );
  OR2_X1 U8721 ( .A1(n9829), .A2(n9834), .ZN(n7438) );
  AND3_X1 U8722 ( .A1(n9837), .A2(n9835), .A3(n9832), .ZN(n9818) );
  INV_X1 U8723 ( .A(n9816), .ZN(n9817) );
  AOI21_X1 U8724 ( .B1(n9824), .B2(n9830), .A(n9825), .ZN(n9816) );
  NAND2_X1 U8725 ( .A1(n9417), .A2(n9416), .ZN(n13182) );
  OR2_X1 U8726 ( .A1(n13297), .A2(n9422), .ZN(n9417) );
  NAND2_X1 U8727 ( .A1(n9407), .A2(n9406), .ZN(n13183) );
  OR2_X1 U8728 ( .A1(n9124), .A2(n11130), .ZN(n9105) );
  OR2_X1 U8729 ( .A1(n9125), .A2(n10078), .ZN(n9106) );
  INV_X1 U8730 ( .A(n6783), .ZN(n10118) );
  NOR2_X1 U8731 ( .A1(n14890), .A2(n6653), .ZN(n10089) );
  NAND2_X1 U8732 ( .A1(n10089), .A2(n10088), .ZN(n10743) );
  NOR2_X1 U8733 ( .A1(n10848), .A2(n6654), .ZN(n10852) );
  NAND2_X1 U8734 ( .A1(n10852), .A2(n10851), .ZN(n11101) );
  INV_X1 U8735 ( .A(n6781), .ZN(n11481) );
  INV_X1 U8736 ( .A(n6779), .ZN(n13237) );
  AOI21_X1 U8737 ( .B1(n6786), .B2(n14863), .A(n6785), .ZN(n13278) );
  INV_X1 U8738 ( .A(n13274), .ZN(n6786) );
  OAI21_X1 U8739 ( .B1(n13275), .B2(n14913), .A(n14930), .ZN(n6785) );
  OAI21_X1 U8740 ( .B1(n13305), .B2(n6754), .A(n13304), .ZN(n13546) );
  NAND2_X1 U8741 ( .A1(n7209), .A2(n7206), .ZN(n13343) );
  NAND2_X1 U8742 ( .A1(n7102), .A2(n9523), .ZN(n13340) );
  AOI21_X1 U8743 ( .B1(n9363), .B2(n6761), .A(n7179), .ZN(n13400) );
  NAND2_X1 U8744 ( .A1(n6730), .A2(n6732), .ZN(n13425) );
  OR2_X1 U8745 ( .A1(n9510), .A2(n6733), .ZN(n6730) );
  NAND2_X1 U8746 ( .A1(n6736), .A2(n9511), .ZN(n13438) );
  NAND2_X1 U8747 ( .A1(n9510), .A2(n6737), .ZN(n6736) );
  NAND2_X1 U8748 ( .A1(n9510), .A2(n9509), .ZN(n13454) );
  NAND2_X1 U8749 ( .A1(n13476), .A2(n9326), .ZN(n13452) );
  NAND2_X1 U8750 ( .A1(n7091), .A2(n7093), .ZN(n13469) );
  OR2_X1 U8751 ( .A1(n13502), .A2(n7097), .ZN(n7091) );
  NAND2_X1 U8752 ( .A1(n7095), .A2(n6568), .ZN(n13483) );
  OR2_X1 U8753 ( .A1(n13502), .A2(n9506), .ZN(n7095) );
  NAND2_X1 U8754 ( .A1(n7205), .A2(n9296), .ZN(n13488) );
  NAND2_X1 U8755 ( .A1(n6771), .A2(n9286), .ZN(n13507) );
  NAND2_X1 U8756 ( .A1(n11601), .A2(n7109), .ZN(n11577) );
  OAI21_X1 U8757 ( .B1(n9244), .B2(n7186), .A(n7184), .ZN(n11575) );
  NAND2_X1 U8758 ( .A1(n7183), .A2(n7187), .ZN(n11576) );
  NAND2_X1 U8759 ( .A1(n9244), .A2(n9243), .ZN(n11597) );
  NAND2_X1 U8760 ( .A1(n11420), .A2(n9218), .ZN(n11355) );
  NAND2_X1 U8761 ( .A1(n6749), .A2(n7099), .ZN(n11423) );
  NAND2_X1 U8762 ( .A1(n11282), .A2(n9492), .ZN(n11298) );
  INV_X1 U8763 ( .A(n13529), .ZN(n13498) );
  INV_X1 U8764 ( .A(n13467), .ZN(n13527) );
  INV_X1 U8765 ( .A(n11131), .ZN(n10582) );
  INV_X1 U8766 ( .A(n13281), .ZN(n13641) );
  AND2_X1 U8767 ( .A1(n13538), .A2(n13537), .ZN(n13639) );
  NAND2_X1 U8768 ( .A1(n6777), .A2(n14982), .ZN(n6776) );
  INV_X1 U8769 ( .A(n13545), .ZN(n6777) );
  INV_X1 U8770 ( .A(n12073), .ZN(n13665) );
  INV_X1 U8771 ( .A(n13510), .ZN(n13678) );
  OR2_X1 U8772 ( .A1(n9967), .A2(n9133), .ZN(n9234) );
  INV_X2 U8773 ( .A(n9145), .ZN(n14818) );
  INV_X1 U8774 ( .A(n14995), .ZN(n14994) );
  AND2_X1 U8775 ( .A1(n10916), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14954) );
  NOR2_X1 U8776 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n7115) );
  NAND2_X1 U8777 ( .A1(n9057), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9059) );
  NAND2_X1 U8778 ( .A1(n9442), .A2(n6719), .ZN(n6718) );
  NOR2_X1 U8779 ( .A1(n9071), .A2(n9454), .ZN(n6719) );
  XNOR2_X1 U8780 ( .A(n9433), .B(n9432), .ZN(n11864) );
  OAI21_X1 U8781 ( .B1(n9453), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9433) );
  INV_X1 U8782 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11247) );
  INV_X1 U8783 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10761) );
  INV_X1 U8784 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10732) );
  INV_X1 U8785 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10046) );
  INV_X1 U8786 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9966) );
  INV_X1 U8787 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9926) );
  INV_X1 U8788 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9900) );
  INV_X1 U8789 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9892) );
  INV_X1 U8790 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9887) );
  INV_X1 U8791 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9878) );
  NAND2_X1 U8792 ( .A1(n9131), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n6788) );
  NAND2_X1 U8793 ( .A1(n10824), .A2(n10823), .ZN(n10989) );
  NAND2_X1 U8794 ( .A1(n7277), .A2(n10659), .ZN(n14595) );
  NAND2_X1 U8795 ( .A1(n13806), .A2(n7491), .ZN(n13732) );
  NAND2_X1 U8796 ( .A1(n10989), .A2(n10988), .ZN(n10991) );
  OR2_X1 U8798 ( .A1(n10074), .A2(n12321), .ZN(n13836) );
  AND2_X1 U8799 ( .A1(n7264), .A2(n7261), .ZN(n13829) );
  NAND2_X1 U8800 ( .A1(n7263), .A2(n7264), .ZN(n13830) );
  OR3_X1 U8801 ( .A1(n12246), .A2(n12245), .A3(n12244), .ZN(n13920) );
  OR2_X1 U8802 ( .A1(n6535), .A2(n10879), .ZN(n7633) );
  OR2_X1 U8803 ( .A1(n12242), .A2(n10880), .ZN(n7634) );
  NAND2_X1 U8804 ( .A1(n13864), .A2(n13863), .ZN(n13862) );
  NAND2_X1 U8805 ( .A1(n13876), .A2(n13877), .ZN(n14628) );
  NOR2_X1 U8806 ( .A1(n9979), .A2(n9978), .ZN(n10035) );
  NOR2_X1 U8807 ( .A1(n10015), .A2(n6882), .ZN(n9979) );
  AND2_X1 U8808 ( .A1(n9990), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6882) );
  XNOR2_X1 U8809 ( .A(n11782), .B(n14646), .ZN(n14644) );
  INV_X1 U8810 ( .A(n6880), .ZN(n13889) );
  NOR2_X1 U8811 ( .A1(n13908), .A2(n6877), .ZN(n13892) );
  NOR2_X1 U8812 ( .A1(n6878), .A2(n13903), .ZN(n6877) );
  OR2_X1 U8813 ( .A1(n13939), .A2(n8110), .ZN(n7088) );
  OR2_X1 U8814 ( .A1(n13939), .A2(n7089), .ZN(n12057) );
  NAND2_X1 U8815 ( .A1(n8074), .A2(n8073), .ZN(n8075) );
  NAND2_X1 U8816 ( .A1(n13991), .A2(n7083), .ZN(n14150) );
  NAND2_X1 U8817 ( .A1(n13991), .A2(n8106), .ZN(n13976) );
  NAND2_X1 U8818 ( .A1(n14001), .A2(n6900), .ZN(n13981) );
  NAND2_X1 U8819 ( .A1(n7073), .A2(n8103), .ZN(n13998) );
  NAND2_X1 U8820 ( .A1(n7396), .A2(n7403), .ZN(n14016) );
  NAND2_X1 U8821 ( .A1(n14055), .A2(n8101), .ZN(n14038) );
  NAND2_X1 U8822 ( .A1(n8098), .A2(n7058), .ZN(n7054) );
  NAND2_X1 U8823 ( .A1(n7384), .A2(n7386), .ZN(n14065) );
  NAND2_X1 U8824 ( .A1(n7385), .A2(n7388), .ZN(n7384) );
  NAND2_X1 U8825 ( .A1(n8098), .A2(n12271), .ZN(n14078) );
  AND2_X1 U8826 ( .A1(n7909), .A2(n7908), .ZN(n14104) );
  NAND2_X1 U8827 ( .A1(n11840), .A2(n8096), .ZN(n14502) );
  AND2_X1 U8828 ( .A1(n12288), .A2(n8093), .ZN(n7069) );
  NAND2_X1 U8829 ( .A1(n7070), .A2(n8093), .ZN(n14123) );
  OAI21_X1 U8830 ( .B1(n11624), .B2(n7395), .A(n7393), .ZN(n11649) );
  NAND2_X1 U8831 ( .A1(n11532), .A2(n12284), .ZN(n7062) );
  NAND2_X1 U8832 ( .A1(n7778), .A2(n7777), .ZN(n14665) );
  NAND2_X1 U8833 ( .A1(n7750), .A2(n7749), .ZN(n11200) );
  INV_X1 U8834 ( .A(n14731), .ZN(n14088) );
  NAND2_X1 U8835 ( .A1(n14711), .A2(n8078), .ZN(n11071) );
  AND2_X1 U8836 ( .A1(n14721), .A2(n13915), .ZN(n14731) );
  NAND2_X1 U8837 ( .A1(n8903), .A2(n6947), .ZN(n8921) );
  NOR2_X1 U8838 ( .A1(n8915), .A2(n6948), .ZN(n6947) );
  OAI21_X1 U8839 ( .B1(n8917), .B2(n14537), .A(n6949), .ZN(n6948) );
  AND4_X1 U8840 ( .A1(n14144), .A2(n14143), .A3(n14142), .A4(n14141), .ZN(
        n14145) );
  OR2_X1 U8841 ( .A1(n14179), .A2(n14178), .ZN(n14206) );
  NAND2_X1 U8842 ( .A1(n7603), .A2(n7602), .ZN(n7606) );
  OR2_X1 U8843 ( .A1(n9092), .A2(n6533), .ZN(n6905) );
  INV_X1 U8844 ( .A(n7116), .ZN(n14227) );
  INV_X1 U8845 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10757) );
  INV_X1 U8846 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10603) );
  INV_X1 U8847 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10056) );
  INV_X1 U8848 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9965) );
  INV_X1 U8849 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9924) );
  INV_X1 U8850 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9913) );
  NAND2_X1 U8851 ( .A1(n7735), .A2(n6867), .ZN(n7752) );
  NOR2_X1 U8852 ( .A1(n7751), .A2(n7415), .ZN(n6867) );
  INV_X1 U8853 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9899) );
  INV_X1 U8854 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9891) );
  OAI21_X1 U8855 ( .B1(n6764), .B2(n7717), .A(n7718), .ZN(n9893) );
  INV_X1 U8856 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9881) );
  NAND2_X1 U8857 ( .A1(n7682), .A2(n7510), .ZN(n7700) );
  INV_X1 U8858 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9879) );
  INV_X1 U8859 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9876) );
  INV_X1 U8860 ( .A(n7648), .ZN(n7650) );
  NAND2_X1 U8861 ( .A1(n6876), .A2(n6874), .ZN(n13868) );
  NAND2_X1 U8862 ( .A1(n6589), .A2(P1_IR_REG_1__SCAN_IN), .ZN(n6876) );
  NOR2_X1 U8863 ( .A1(n7628), .A2(n6875), .ZN(n6874) );
  AOI21_X1 U8864 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n14288), .A(n15342), .ZN(
        n15334) );
  XNOR2_X1 U8865 ( .A(n6683), .B(n14292), .ZN(n15337) );
  INV_X1 U8866 ( .A(n14291), .ZN(n6683) );
  XNOR2_X1 U8867 ( .A(n14294), .B(n14889), .ZN(n14347) );
  XNOR2_X1 U8868 ( .A(n14299), .B(n14300), .ZN(n15340) );
  INV_X1 U8869 ( .A(n14305), .ZN(n6928) );
  NAND2_X1 U8870 ( .A1(n14349), .A2(n14904), .ZN(n14348) );
  XNOR2_X1 U8871 ( .A(n14308), .B(n14307), .ZN(n14351) );
  OAI21_X1 U8872 ( .B1(n14355), .B2(n14354), .A(n6704), .ZN(n6703) );
  NAND2_X1 U8873 ( .A1(n6920), .A2(n14567), .ZN(n14573) );
  OAI21_X1 U8874 ( .B1(n14568), .B2(n14569), .A(n6921), .ZN(n6920) );
  INV_X1 U8875 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n6921) );
  NAND2_X1 U8876 ( .A1(n6918), .A2(n14571), .ZN(n14577) );
  OAI21_X1 U8877 ( .B1(n14573), .B2(n14572), .A(n6919), .ZN(n6918) );
  INV_X1 U8878 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6919) );
  NOR2_X1 U8879 ( .A1(n14577), .A2(n14576), .ZN(n14575) );
  NAND2_X1 U8880 ( .A1(n14589), .A2(n14590), .ZN(n14588) );
  OAI21_X1 U8881 ( .B1(n14589), .B2(n14590), .A(n6917), .ZN(n6916) );
  AOI21_X1 U8882 ( .B1(n6802), .B2(n6803), .A(n6797), .ZN(n12629) );
  AOI21_X1 U8883 ( .B1(n6813), .B2(n15178), .A(n6810), .ZN(n12679) );
  XNOR2_X1 U8884 ( .A(n6815), .B(n6814), .ZN(n6813) );
  OAI21_X1 U8885 ( .B1(n12697), .B2(n12903), .A(n6688), .ZN(P3_U3488) );
  INV_X1 U8886 ( .A(n6689), .ZN(n6688) );
  OAI21_X1 U8887 ( .B1(n8983), .B2(n15329), .A(n7367), .ZN(n6689) );
  INV_X1 U8888 ( .A(n7368), .ZN(n7367) );
  OR2_X1 U8889 ( .A1(n12697), .A2(n12975), .ZN(n9031) );
  NAND2_X1 U8890 ( .A1(n9549), .A2(n6599), .ZN(P2_U3236) );
  AND2_X1 U8891 ( .A1(n9821), .A2(n13634), .ZN(n6690) );
  NAND2_X1 U8892 ( .A1(n7107), .A2(n7106), .ZN(P2_U3528) );
  NAND2_X1 U8893 ( .A1(n6478), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n7106) );
  NAND2_X1 U8894 ( .A1(n13642), .A2(n15002), .ZN(n7107) );
  AND2_X1 U8895 ( .A1(n9821), .A2(n13680), .ZN(n6691) );
  INV_X1 U8896 ( .A(n6697), .ZN(n6696) );
  OAI21_X1 U8897 ( .B1(n13938), .B2(n13817), .A(n12051), .ZN(n6697) );
  OAI21_X1 U8898 ( .B1(n13916), .B2(n14511), .A(n6870), .ZN(P1_U3262) );
  AOI21_X1 U8899 ( .B1(n6872), .B2(n14511), .A(n6871), .ZN(n6870) );
  OAI21_X1 U8900 ( .B1(n14653), .B2(n7498), .A(n13917), .ZN(n6871) );
  INV_X1 U8901 ( .A(n8918), .ZN(n8919) );
  INV_X1 U8902 ( .A(n8902), .ZN(n6903) );
  INV_X1 U8903 ( .A(n14585), .ZN(n14584) );
  XNOR2_X1 U8904 ( .A(n14331), .B(n14334), .ZN(n6929) );
  NAND2_X1 U8905 ( .A1(n14079), .A2(n7390), .ZN(n7389) );
  NAND2_X1 U8906 ( .A1(n7840), .A2(n7839), .ZN(n12151) );
  INV_X2 U8907 ( .A(n10719), .ZN(n10969) );
  AND2_X1 U8908 ( .A1(n7283), .A2(n12457), .ZN(n6546) );
  NAND2_X1 U8909 ( .A1(n7349), .A2(n7347), .ZN(n12803) );
  AND2_X1 U8910 ( .A1(n9637), .A2(n9636), .ZN(n6548) );
  OR2_X1 U8911 ( .A1(n12982), .A2(n12824), .ZN(n8810) );
  NAND2_X1 U8912 ( .A1(n9365), .A2(n9364), .ZN(n13404) );
  INV_X1 U8913 ( .A(n8952), .ZN(n7345) );
  AND2_X1 U8914 ( .A1(n14064), .A2(n7055), .ZN(n6549) );
  AND2_X1 U8915 ( .A1(n6895), .A2(n6610), .ZN(n6550) );
  AND2_X1 U8916 ( .A1(n12130), .A2(n7147), .ZN(n6551) );
  OR2_X1 U8917 ( .A1(n10428), .A2(n6709), .ZN(n6552) );
  NAND2_X1 U8918 ( .A1(n8042), .A2(n8041), .ZN(n12344) );
  AND2_X1 U8919 ( .A1(n9628), .A2(n6640), .ZN(n6553) );
  OR2_X1 U8920 ( .A1(n14155), .A2(n7371), .ZN(n6554) );
  INV_X1 U8921 ( .A(n12200), .ZN(n7150) );
  AND2_X1 U8922 ( .A1(n6746), .A2(n9493), .ZN(n6555) );
  NAND2_X1 U8923 ( .A1(n7267), .A2(n6559), .ZN(n13915) );
  AND2_X1 U8924 ( .A1(n13601), .A2(n9350), .ZN(n6556) );
  AND2_X1 U8925 ( .A1(n6906), .A2(n13359), .ZN(n6557) );
  NAND2_X1 U8926 ( .A1(n7467), .A2(n7466), .ZN(n6558) );
  AND2_X1 U8927 ( .A1(n8062), .A2(n7265), .ZN(n6559) );
  AND2_X1 U8928 ( .A1(n11578), .A2(n9501), .ZN(n7109) );
  INV_X1 U8929 ( .A(n9611), .ZN(n9641) );
  NAND3_X1 U8930 ( .A1(n6840), .A2(n6841), .A3(n12065), .ZN(n9611) );
  NOR2_X1 U8931 ( .A1(n11741), .A2(n9502), .ZN(n6560) );
  INV_X1 U8932 ( .A(n12297), .ZN(n13941) );
  INV_X1 U8933 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n9069) );
  INV_X1 U8934 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8161) );
  INV_X1 U8935 ( .A(n9705), .ZN(n6833) );
  AND2_X1 U8936 ( .A1(n7303), .A2(n7302), .ZN(n6561) );
  AND2_X1 U8937 ( .A1(n9705), .A2(n6641), .ZN(n6562) );
  AND2_X1 U8938 ( .A1(n6939), .A2(n6940), .ZN(n6563) );
  AND2_X1 U8939 ( .A1(n7272), .A2(n7270), .ZN(n6564) );
  INV_X1 U8940 ( .A(n7389), .ZN(n7388) );
  AND2_X1 U8941 ( .A1(n13590), .A2(n13190), .ZN(n7179) );
  NAND2_X1 U8942 ( .A1(n7281), .A2(n6546), .ZN(n12456) );
  NOR2_X1 U8943 ( .A1(n6836), .A2(n6839), .ZN(n7246) );
  INV_X2 U8944 ( .A(n15329), .ZN(n15331) );
  AND2_X1 U8945 ( .A1(n9501), .A2(n9499), .ZN(n11596) );
  NAND2_X1 U8946 ( .A1(n9449), .A2(n9450), .ZN(n12419) );
  INV_X1 U8947 ( .A(n12419), .ZN(n6841) );
  AND2_X1 U8948 ( .A1(n6672), .A2(n8632), .ZN(n6565) );
  AND2_X1 U8949 ( .A1(n7379), .A2(n7380), .ZN(n6566) );
  INV_X1 U8950 ( .A(n9048), .ZN(n9132) );
  INV_X1 U8951 ( .A(n12290), .ZN(n11848) );
  XOR2_X1 U8952 ( .A(n13580), .B(n6469), .Z(n6567) );
  INV_X1 U8953 ( .A(n9677), .ZN(n7461) );
  OR2_X1 U8954 ( .A1(n13678), .A2(n13196), .ZN(n6568) );
  INV_X1 U8955 ( .A(n6839), .ZN(n9205) );
  AND2_X1 U8956 ( .A1(n12366), .A2(n12856), .ZN(n6569) );
  NOR2_X1 U8957 ( .A1(n12074), .A2(n12069), .ZN(n6570) );
  NOR2_X1 U8958 ( .A1(n6676), .A2(n13759), .ZN(n13758) );
  AND2_X1 U8959 ( .A1(n7312), .A2(n12491), .ZN(n6571) );
  AND2_X1 U8960 ( .A1(n12504), .A2(n7285), .ZN(n6572) );
  NAND2_X1 U8961 ( .A1(n11640), .A2(n12559), .ZN(n6573) );
  AND2_X1 U8962 ( .A1(n9569), .A2(n9568), .ZN(n6574) );
  OR2_X1 U8963 ( .A1(n9694), .A2(n9693), .ZN(n6575) );
  INV_X1 U8964 ( .A(n13344), .ZN(n7216) );
  AND2_X1 U8965 ( .A1(n9714), .A2(n9713), .ZN(n6576) );
  NOR2_X1 U8966 ( .A1(n11750), .A2(n11751), .ZN(n6577) );
  AND2_X1 U8967 ( .A1(n6906), .A2(n13401), .ZN(n6579) );
  OR2_X1 U8968 ( .A1(n12632), .A2(n15200), .ZN(n6580) );
  INV_X1 U8969 ( .A(n7097), .ZN(n7096) );
  NAND2_X1 U8970 ( .A1(n13486), .A2(n7098), .ZN(n7097) );
  AND2_X1 U8971 ( .A1(n12966), .A2(n12796), .ZN(n6581) );
  AND2_X1 U8972 ( .A1(n14188), .A2(n14066), .ZN(n6582) );
  AND2_X1 U8973 ( .A1(n8824), .A2(n6991), .ZN(n6583) );
  NAND2_X1 U8974 ( .A1(n9356), .A2(n9355), .ZN(n13596) );
  INV_X1 U8975 ( .A(n8956), .ZN(n12794) );
  OR2_X1 U8976 ( .A1(n14416), .A2(n12583), .ZN(n6584) );
  AND3_X1 U8977 ( .A1(n8326), .A2(n8325), .A3(n8324), .ZN(n11402) );
  INV_X1 U8978 ( .A(n11402), .ZN(n7322) );
  INV_X1 U8979 ( .A(n7487), .ZN(n7226) );
  NOR3_X1 U8980 ( .A1(n12171), .A2(n12170), .A3(n12179), .ZN(n6585) );
  AND2_X1 U8981 ( .A1(n11038), .A2(n11170), .ZN(n6586) );
  AND2_X1 U8982 ( .A1(n7926), .A2(n7925), .ZN(n14188) );
  INV_X1 U8983 ( .A(n14188), .ZN(n14091) );
  AND4_X1 U8984 ( .A1(n6695), .A2(n6694), .A3(n12319), .A4(n6692), .ZN(n6587)
         );
  NAND4_X1 U8985 ( .A1(n7050), .A2(n7049), .A3(n7376), .A4(n7574), .ZN(n8127)
         );
  AND2_X1 U8986 ( .A1(n12369), .A2(n12855), .ZN(n6588) );
  INV_X1 U8987 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9166) );
  AND2_X1 U8988 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6589) );
  AND2_X1 U8989 ( .A1(n12560), .A2(n11327), .ZN(n6590) );
  INV_X1 U8990 ( .A(n13548), .ZN(n6912) );
  AND3_X1 U8991 ( .A1(n9340), .A2(n9437), .A3(n9055), .ZN(n6591) );
  NOR2_X1 U8992 ( .A1(n13526), .A2(n13198), .ZN(n6592) );
  AOI21_X1 U8993 ( .B1(n7000), .B2(n8782), .A(n6999), .ZN(n6998) );
  NAND2_X1 U8994 ( .A1(n7582), .A2(n7581), .ZN(n14155) );
  NOR2_X1 U8995 ( .A1(n13355), .A2(n9397), .ZN(n6593) );
  AND2_X1 U8996 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n6594) );
  AND2_X1 U8997 ( .A1(n13562), .A2(n13128), .ZN(n6595) );
  AND2_X1 U8998 ( .A1(n9619), .A2(n9618), .ZN(n6596) );
  AND2_X1 U8999 ( .A1(n8803), .A2(n8806), .ZN(n12821) );
  AND2_X1 U9000 ( .A1(n9721), .A2(n9720), .ZN(n6597) );
  NAND2_X1 U9001 ( .A1(n13344), .A2(n7211), .ZN(n7210) );
  INV_X1 U9002 ( .A(n7210), .ZN(n7206) );
  INV_X1 U9003 ( .A(n6944), .ZN(n13935) );
  INV_X1 U9004 ( .A(n6913), .ZN(n13316) );
  INV_X1 U9005 ( .A(n12134), .ZN(n7145) );
  INV_X1 U9006 ( .A(n7287), .ZN(n7286) );
  AND2_X1 U9007 ( .A1(n9216), .A2(n7099), .ZN(n6598) );
  AND2_X1 U9008 ( .A1(n7490), .A2(n9548), .ZN(n6599) );
  AND2_X1 U9009 ( .A1(n9132), .A2(n6787), .ZN(n6600) );
  INV_X1 U9010 ( .A(n6862), .ZN(n6861) );
  NAND2_X1 U9011 ( .A1(n13769), .A2(n6863), .ZN(n6862) );
  NAND2_X1 U9012 ( .A1(n7517), .A2(SI_7_), .ZN(n7519) );
  INV_X1 U9013 ( .A(n7519), .ZN(n7415) );
  AND2_X1 U9014 ( .A1(n12887), .A2(n12738), .ZN(n6601) );
  AND2_X1 U9015 ( .A1(n13975), .A2(n6554), .ZN(n6602) );
  AND2_X1 U9016 ( .A1(n7174), .A2(n7170), .ZN(n6603) );
  NAND2_X1 U9017 ( .A1(n9659), .A2(n9656), .ZN(n6604) );
  AND2_X1 U9018 ( .A1(n6868), .A2(n10988), .ZN(n6605) );
  INV_X1 U9019 ( .A(n7163), .ZN(n7162) );
  NAND2_X1 U9020 ( .A1(n14122), .A2(n7164), .ZN(n7163) );
  NOR2_X1 U9021 ( .A1(n14368), .A2(n6569), .ZN(n6606) );
  INV_X1 U9022 ( .A(n6946), .ZN(n13970) );
  INV_X1 U9023 ( .A(n6738), .ZN(n6737) );
  OR2_X1 U9024 ( .A1(n9512), .A2(n6739), .ZN(n6738) );
  NAND4_X2 U9025 ( .A1(n7696), .A2(n7695), .A3(n7694), .A4(n7693), .ZN(n14598)
         );
  AND2_X1 U9026 ( .A1(n7323), .A2(n8860), .ZN(n6607) );
  INV_X1 U9027 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8860) );
  INV_X1 U9028 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7579) );
  AND2_X1 U9029 ( .A1(n11731), .A2(n12557), .ZN(n6608) );
  AND2_X1 U9030 ( .A1(n14975), .A2(n11191), .ZN(n6609) );
  NAND2_X1 U9031 ( .A1(n9446), .A2(n9431), .ZN(n9450) );
  OR2_X1 U9032 ( .A1(n7544), .A2(SI_17_), .ZN(n6610) );
  INV_X1 U9033 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n7719) );
  NOR2_X1 U9034 ( .A1(n11741), .A2(n13197), .ZN(n6611) );
  NOR2_X1 U9035 ( .A1(n14531), .A2(n13850), .ZN(n6612) );
  NOR2_X1 U9036 ( .A1(n14521), .A2(n13852), .ZN(n6613) );
  NOR2_X1 U9037 ( .A1(n14181), .A2(n14081), .ZN(n6614) );
  INV_X1 U9038 ( .A(n8109), .ZN(n8110) );
  NOR2_X1 U9039 ( .A1(n13580), .A2(n9704), .ZN(n6615) );
  NOR2_X1 U9040 ( .A1(n12151), .A2(n12152), .ZN(n6616) );
  INV_X1 U9041 ( .A(n7493), .ZN(n7190) );
  INV_X1 U9042 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9897) );
  AND2_X1 U9043 ( .A1(n13447), .A2(n7195), .ZN(n6617) );
  OR2_X1 U9044 ( .A1(n7174), .A2(n7170), .ZN(n6618) );
  AND2_X1 U9045 ( .A1(n13672), .A2(n9507), .ZN(n6619) );
  AND2_X1 U9046 ( .A1(n10083), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6620) );
  OR2_X1 U9047 ( .A1(n12336), .A2(n12335), .ZN(n6621) );
  NAND2_X1 U9048 ( .A1(n7151), .A2(n7148), .ZN(n6622) );
  NOR2_X1 U9049 ( .A1(n12370), .A2(n12371), .ZN(n6623) );
  NOR2_X1 U9050 ( .A1(n14044), .A2(n7968), .ZN(n6624) );
  INV_X1 U9051 ( .A(n12139), .ZN(n7122) );
  OR2_X1 U9052 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), .ZN(
        n6625) );
  AND3_X1 U9053 ( .A1(n9793), .A2(n9795), .A3(n9794), .ZN(n6626) );
  INV_X1 U9054 ( .A(n8946), .ZN(n12854) );
  AND2_X1 U9055 ( .A1(n7530), .A2(n9889), .ZN(n6627) );
  INV_X1 U9056 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9868) );
  INV_X1 U9057 ( .A(n7011), .ZN(n7010) );
  AND2_X1 U9058 ( .A1(n11983), .A2(n11982), .ZN(n6628) );
  INV_X1 U9059 ( .A(n12293), .ZN(n14037) );
  OR2_X1 U9060 ( .A1(n7227), .A2(n7487), .ZN(n6629) );
  AND2_X1 U9061 ( .A1(n9326), .A2(n9324), .ZN(n9786) );
  INV_X1 U9062 ( .A(n9786), .ZN(n13474) );
  AND2_X1 U9063 ( .A1(n7464), .A2(n6596), .ZN(n6630) );
  AND2_X1 U9064 ( .A1(n6552), .A2(n6794), .ZN(n6631) );
  NAND2_X1 U9065 ( .A1(n13451), .A2(n7198), .ZN(n6632) );
  NOR2_X1 U9066 ( .A1(n12153), .A2(n12154), .ZN(n6633) );
  OR2_X1 U9067 ( .A1(n8804), .A2(n6980), .ZN(n6634) );
  INV_X1 U9068 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n14232) );
  INV_X1 U9069 ( .A(n7179), .ZN(n6762) );
  INV_X1 U9070 ( .A(n12219), .ZN(n7126) );
  INV_X1 U9071 ( .A(n12118), .ZN(n7130) );
  INV_X1 U9072 ( .A(n12209), .ZN(n7134) );
  INV_X1 U9073 ( .A(n12204), .ZN(n7139) );
  AND2_X1 U9074 ( .A1(n6731), .A2(n13426), .ZN(n6635) );
  OR2_X1 U9075 ( .A1(n9718), .A2(n9719), .ZN(n6636) );
  OR2_X1 U9076 ( .A1(n12377), .A2(n12808), .ZN(n6637) );
  INV_X1 U9077 ( .A(n12288), .ZN(n14122) );
  INV_X1 U9078 ( .A(n12294), .ZN(n13975) );
  AND2_X1 U9079 ( .A1(n12159), .A2(n7897), .ZN(n6638) );
  NOR2_X1 U9080 ( .A1(n7383), .A2(n14064), .ZN(n7382) );
  NAND2_X1 U9081 ( .A1(n9490), .A2(n14964), .ZN(n6639) );
  AND2_X1 U9082 ( .A1(n9626), .A2(n9625), .ZN(n6640) );
  AND2_X1 U9083 ( .A1(n9702), .A2(n9701), .ZN(n6641) );
  OR2_X1 U9084 ( .A1(n9831), .A2(n9830), .ZN(n6642) );
  AND2_X1 U9085 ( .A1(n6900), .A2(n13994), .ZN(n6643) );
  INV_X1 U9086 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n9054) );
  AND2_X1 U9087 ( .A1(n7171), .A2(n6618), .ZN(n6644) );
  AND2_X1 U9088 ( .A1(n7583), .A2(n7579), .ZN(n6645) );
  AND2_X1 U9089 ( .A1(n6577), .A2(n7274), .ZN(n6646) );
  AND2_X1 U9090 ( .A1(n12270), .A2(n12269), .ZN(n6647) );
  AND2_X1 U9091 ( .A1(n9231), .A2(n9230), .ZN(n9782) );
  INV_X1 U9092 ( .A(n9782), .ZN(n7204) );
  INV_X1 U9093 ( .A(n11268), .ZN(n7243) );
  INV_X1 U9094 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7266) );
  INV_X1 U9095 ( .A(n7340), .ZN(n7339) );
  OR2_X1 U9096 ( .A1(n13637), .A2(n6691), .ZN(P2_U3498) );
  OR2_X1 U9097 ( .A1(n13536), .A2(n6690), .ZN(P2_U3530) );
  NAND2_X1 U9098 ( .A1(n9799), .A2(n11552), .ZN(n9478) );
  INV_X1 U9099 ( .A(n12476), .ZN(n7302) );
  INV_X1 U9100 ( .A(n13562), .ZN(n7215) );
  INV_X1 U9101 ( .A(n14044), .ZN(n6939) );
  NAND2_X1 U9102 ( .A1(n9205), .A2(n6835), .ZN(n9339) );
  NAND2_X1 U9103 ( .A1(n6983), .A2(n6982), .ZN(n8411) );
  AND2_X1 U9104 ( .A1(n14099), .A2(n6942), .ZN(n6650) );
  INV_X1 U9105 ( .A(n8699), .ZN(n7001) );
  INV_X1 U9106 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6715) );
  OR2_X1 U9107 ( .A1(n12640), .A2(n12622), .ZN(n6651) );
  AND2_X1 U9108 ( .A1(n14911), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6652) );
  OAI21_X1 U9109 ( .B1(n12450), .B2(n12449), .A(n7286), .ZN(n12503) );
  AND2_X1 U9110 ( .A1(n10105), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6653) );
  NAND2_X1 U9111 ( .A1(n7295), .A2(n7300), .ZN(n12473) );
  NAND2_X1 U9112 ( .A1(n9363), .A2(n9362), .ZN(n13419) );
  INV_X1 U9113 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7366) );
  AND2_X1 U9114 ( .A1(n10849), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6654) );
  NAND2_X1 U9115 ( .A1(n7272), .A2(n7273), .ZN(n11685) );
  INV_X1 U9116 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n7704) );
  AND3_X1 U9117 ( .A1(n7378), .A2(n7375), .A3(n7373), .ZN(n6655) );
  INV_X1 U9118 ( .A(n13184), .ZN(n13118) );
  INV_X1 U9119 ( .A(n8961), .ZN(n12776) );
  AND2_X1 U9120 ( .A1(n12747), .A2(n8829), .ZN(n12761) );
  INV_X1 U9121 ( .A(n6911), .ZN(n7495) );
  AND2_X1 U9122 ( .A1(n7002), .A2(n8699), .ZN(n6656) );
  AND2_X1 U9123 ( .A1(n7686), .A2(n7685), .ZN(n14620) );
  INV_X1 U9124 ( .A(n14620), .ZN(n6884) );
  AND2_X1 U9125 ( .A1(n7349), .A2(n8953), .ZN(n6657) );
  AND2_X1 U9126 ( .A1(n11601), .A2(n9501), .ZN(n6658) );
  AND2_X1 U9127 ( .A1(n7544), .A2(SI_17_), .ZN(n6659) );
  NAND2_X1 U9128 ( .A1(n12644), .A2(n12643), .ZN(n6660) );
  NAND2_X1 U9129 ( .A1(n7054), .A2(n12189), .ZN(n14073) );
  INV_X1 U9130 ( .A(n7246), .ZN(n9430) );
  INV_X1 U9131 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9043) );
  AND2_X1 U9132 ( .A1(n7281), .A2(n7283), .ZN(n6661) );
  NAND2_X1 U9133 ( .A1(n6748), .A2(n6639), .ZN(n6747) );
  NAND2_X1 U9134 ( .A1(n7326), .A2(n8934), .ZN(n11454) );
  NAND2_X1 U9135 ( .A1(n7194), .A2(n9178), .ZN(n11287) );
  NAND2_X1 U9136 ( .A1(n7062), .A2(n8090), .ZN(n14522) );
  AND2_X1 U9137 ( .A1(n15135), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n6662) );
  NAND2_X1 U9138 ( .A1(n7304), .A2(n8988), .ZN(n10624) );
  OR2_X1 U9139 ( .A1(n15331), .A2(n9014), .ZN(n6663) );
  AND2_X1 U9140 ( .A1(n15139), .A2(n12652), .ZN(n6664) );
  AND2_X1 U9141 ( .A1(n6747), .A2(n9491), .ZN(n6665) );
  INV_X1 U9142 ( .A(n7978), .ZN(n7422) );
  AND2_X1 U9143 ( .A1(n7352), .A2(n8930), .ZN(n6666) );
  NAND2_X1 U9144 ( .A1(n7321), .A2(n7320), .ZN(n6667) );
  AND2_X1 U9145 ( .A1(n12613), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n6668) );
  OR2_X1 U9146 ( .A1(n9478), .A2(n12419), .ZN(n6669) );
  AND2_X1 U9147 ( .A1(n6795), .A2(n6794), .ZN(n6670) );
  NAND2_X1 U9148 ( .A1(n11131), .A2(n11146), .ZN(n10574) );
  INV_X1 U9149 ( .A(n10574), .ZN(n6910) );
  INV_X1 U9150 ( .A(n9473), .ZN(n9798) );
  AND2_X1 U9151 ( .A1(n14986), .A2(n14987), .ZN(n13622) );
  OR2_X1 U9152 ( .A1(n14389), .A2(n6959), .ZN(n6671) );
  NAND2_X1 U9153 ( .A1(n12061), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6672) );
  OR2_X1 U9155 ( .A1(n6668), .A2(n12666), .ZN(n6673) );
  NAND2_X1 U9156 ( .A1(n12249), .A2(n8064), .ZN(n14716) );
  INV_X1 U9157 ( .A(n14627), .ZN(n6885) );
  INV_X1 U9158 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n6934) );
  INV_X1 U9159 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n6704) );
  INV_X1 U9160 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n6917) );
  NAND2_X1 U9161 ( .A1(n10072), .A2(n9904), .ZN(n6674) );
  AND2_X1 U9162 ( .A1(n10064), .A2(n9850), .ZN(n10072) );
  NAND2_X1 U9163 ( .A1(n6675), .A2(n9529), .ZN(n13484) );
  NAND2_X1 U9164 ( .A1(n9798), .A2(n6841), .ZN(n6675) );
  NAND2_X1 U9165 ( .A1(n13302), .A2(n13484), .ZN(n6754) );
  INV_X1 U9166 ( .A(n13484), .ZN(n13504) );
  NAND2_X1 U9167 ( .A1(n10723), .A2(n10722), .ZN(n10799) );
  NAND2_X1 U9168 ( .A1(n10971), .A2(n10970), .ZN(n10972) );
  NAND2_X1 U9169 ( .A1(n12469), .A2(n12398), .ZN(n12529) );
  OAI21_X1 U9170 ( .B1(n11325), .B2(n7318), .A(n7317), .ZN(n7489) );
  XNOR2_X1 U9171 ( .A(n12434), .B(n12435), .ZN(n12436) );
  XNOR2_X1 U9172 ( .A(n7489), .B(n11722), .ZN(n11723) );
  NAND2_X1 U9173 ( .A1(n8156), .A2(n8157), .ZN(n8160) );
  OR2_X2 U9174 ( .A1(n12514), .A2(n12554), .ZN(n12512) );
  NAND2_X1 U9175 ( .A1(n12384), .A2(n12385), .ZN(n12514) );
  NAND2_X1 U9176 ( .A1(n10804), .A2(n10803), .ZN(n10971) );
  NAND2_X1 U9177 ( .A1(n11324), .A2(n11323), .ZN(n11325) );
  NAND2_X1 U9178 ( .A1(n10972), .A2(n10973), .ZN(n11313) );
  NAND2_X1 U9179 ( .A1(n12365), .A2(n7484), .ZN(n14369) );
  NAND2_X1 U9180 ( .A1(n13104), .A2(n6705), .ZN(n13038) );
  AOI21_X2 U9181 ( .B1(n7237), .B2(n7236), .A(n13144), .ZN(n13134) );
  OAI21_X1 U9182 ( .B1(n6869), .B2(SI_4_), .A(n7510), .ZN(n7509) );
  NAND2_X2 U9183 ( .A1(n10948), .A2(n12352), .ZN(n12359) );
  NAND2_X1 U9184 ( .A1(n7220), .A2(n7219), .ZN(n11699) );
  NAND2_X1 U9185 ( .A1(n6677), .A2(n7268), .ZN(n11768) );
  NAND2_X1 U9186 ( .A1(n13741), .A2(n13740), .ZN(n13739) );
  NAND2_X1 U9187 ( .A1(n11680), .A2(n11679), .ZN(n14482) );
  NOR2_X1 U9188 ( .A1(n11713), .A2(n11571), .ZN(n11804) );
  NAND2_X1 U9189 ( .A1(n11260), .A2(n11048), .ZN(n11049) );
  NAND2_X1 U9190 ( .A1(n14482), .A2(n6646), .ZN(n6677) );
  NAND2_X1 U9191 ( .A1(n10378), .A2(n10377), .ZN(n10383) );
  NAND2_X1 U9192 ( .A1(n10173), .A2(n10174), .ZN(n10377) );
  NOR2_X2 U9193 ( .A1(n13714), .A2(n13715), .ZN(n13713) );
  NAND2_X1 U9194 ( .A1(n11444), .A2(n11443), .ZN(n11680) );
  AOI21_X1 U9195 ( .B1(n9540), .B2(n13484), .A(n9539), .ZN(n13544) );
  INV_X1 U9196 ( .A(n6727), .ZN(n6726) );
  NAND2_X1 U9197 ( .A1(n6726), .A2(n6724), .ZN(n6723) );
  NAND2_X1 U9198 ( .A1(n7682), .A2(n7681), .ZN(n9880) );
  XNOR2_X1 U9199 ( .A(n10932), .B(n10927), .ZN(n12351) );
  NAND2_X1 U9200 ( .A1(n11000), .A2(n7731), .ZN(n14675) );
  NAND2_X1 U9201 ( .A1(n7715), .A2(n7714), .ZN(n14693) );
  INV_X1 U9203 ( .A(n7241), .ZN(n7240) );
  NAND2_X1 U9204 ( .A1(n7392), .A2(n7391), .ZN(n14112) );
  OAI21_X2 U9205 ( .B1(n7417), .B2(n7418), .A(n7416), .ZN(n8016) );
  OAI21_X1 U9206 ( .B1(n8035), .B2(n11762), .A(n8034), .ZN(n8037) );
  INV_X1 U9207 ( .A(n12320), .ZN(n6693) );
  NAND2_X1 U9208 ( .A1(n6693), .A2(n6647), .ZN(n6692) );
  NAND2_X1 U9209 ( .A1(n12257), .A2(n12258), .ZN(n12259) );
  NAND2_X1 U9210 ( .A1(n8037), .A2(n8036), .ZN(n8881) );
  NAND2_X1 U9211 ( .A1(n9740), .A2(n9739), .ZN(n9755) );
  NOR2_X1 U9212 ( .A1(n7400), .A2(n7404), .ZN(n7399) );
  NAND2_X1 U9213 ( .A1(n8018), .A2(n8017), .ZN(n8035) );
  NOR2_X1 U9214 ( .A1(n14056), .A2(n7406), .ZN(n7405) );
  NOR2_X1 U9215 ( .A1(n9834), .A2(n9833), .ZN(n9836) );
  NAND2_X1 U9216 ( .A1(n14573), .A2(n14572), .ZN(n14571) );
  NAND2_X1 U9217 ( .A1(n12792), .A2(n8815), .ZN(n12783) );
  NAND2_X1 U9218 ( .A1(n15337), .A2(n15336), .ZN(n15335) );
  AND3_X2 U9219 ( .A1(n6982), .A2(n6983), .A3(n6817), .ZN(n8430) );
  NAND2_X1 U9220 ( .A1(n14568), .A2(n14569), .ZN(n14567) );
  XNOR2_X1 U9221 ( .A(n14304), .B(n6928), .ZN(n14349) );
  NAND2_X1 U9222 ( .A1(n14316), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6701) );
  NAND2_X1 U9223 ( .A1(n14279), .A2(n14278), .ZN(n6925) );
  INV_X1 U9224 ( .A(n11829), .ZN(n6680) );
  OAI21_X2 U9225 ( .B1(n11514), .B2(n7011), .A(n7007), .ZN(n11616) );
  NAND2_X1 U9226 ( .A1(n14586), .A2(n14587), .ZN(n14583) );
  NOR2_X1 U9227 ( .A1(n14347), .A2(n14346), .ZN(n14345) );
  NOR2_X1 U9228 ( .A1(n15341), .A2(n15340), .ZN(n15339) );
  NAND2_X1 U9229 ( .A1(n8214), .A2(n15239), .ZN(n15234) );
  NAND2_X1 U9230 ( .A1(n14336), .A2(n14337), .ZN(n14335) );
  NAND3_X1 U9231 ( .A1(n8163), .A2(n8164), .A3(n8162), .ZN(n8167) );
  OAI21_X2 U9232 ( .B1(n8179), .B2(P3_IR_REG_28__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8170) );
  NAND2_X1 U9233 ( .A1(n11049), .A2(n11255), .ZN(n11263) );
  INV_X1 U9234 ( .A(n6681), .ZN(n8497) );
  NOR2_X4 U9235 ( .A1(n6838), .A2(n6839), .ZN(n9327) );
  NAND2_X1 U9236 ( .A1(n14353), .A2(n6703), .ZN(n14568) );
  NAND2_X1 U9237 ( .A1(n6931), .A2(n14335), .ZN(n6930) );
  XNOR2_X1 U9238 ( .A(n6930), .B(n6929), .ZN(SUB_1596_U4) );
  NAND4_X1 U9239 ( .A1(n6684), .A2(n9838), .A3(n6642), .A4(n7438), .ZN(n9840)
         );
  NAND2_X1 U9240 ( .A1(n9809), .A2(n6626), .ZN(n9796) );
  NAND2_X2 U9241 ( .A1(n8097), .A2(n12272), .ZN(n8098) );
  NAND3_X1 U9242 ( .A1(n6865), .A2(n7699), .A3(n6763), .ZN(n7702) );
  NAND2_X1 U9243 ( .A1(n14026), .A2(n14027), .ZN(n7073) );
  NAND2_X1 U9244 ( .A1(n11647), .A2(n11648), .ZN(n7070) );
  INV_X1 U9245 ( .A(n9824), .ZN(n7437) );
  OAI21_X1 U9246 ( .B1(n7503), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n6685), .ZN(
        n7500) );
  NAND2_X1 U9247 ( .A1(n7503), .A2(n9120), .ZN(n6685) );
  NAND2_X1 U9248 ( .A1(n6686), .A2(n10941), .ZN(n14814) );
  NAND2_X1 U9249 ( .A1(n11213), .A2(n10940), .ZN(n6686) );
  NAND2_X1 U9250 ( .A1(n10407), .A2(n6474), .ZN(n11141) );
  NAND2_X1 U9251 ( .A1(n13052), .A2(n13111), .ZN(n13114) );
  NAND2_X1 U9252 ( .A1(n9327), .A2(n6720), .ZN(n9442) );
  NAND2_X1 U9253 ( .A1(n11169), .A2(n10937), .ZN(n14815) );
  NAND2_X1 U9254 ( .A1(n10943), .A2(n10942), .ZN(n11212) );
  NOR2_X1 U9255 ( .A1(n9339), .A2(n7247), .ZN(n9455) );
  INV_X1 U9256 ( .A(n11699), .ZN(n14823) );
  NAND2_X1 U9257 ( .A1(n8509), .A2(n8508), .ZN(n8511) );
  NOR2_X1 U9258 ( .A1(n13134), .A2(n6707), .ZN(n13106) );
  OAI211_X1 U9259 ( .C1(n11713), .C2(n11712), .A(n11711), .B(n11710), .ZN(
        n11714) );
  NAND2_X1 U9260 ( .A1(n8338), .A2(n8337), .ZN(n8353) );
  NOR2_X1 U9261 ( .A1(n14442), .A2(n14441), .ZN(n14443) );
  NOR2_X1 U9262 ( .A1(n12573), .A2(n15077), .ZN(n15094) );
  AOI21_X2 U9263 ( .B1(n10689), .B2(n10688), .A(n10687), .ZN(n10696) );
  XNOR2_X2 U9264 ( .A(n8181), .B(n8180), .ZN(n12328) );
  NAND2_X1 U9265 ( .A1(n12841), .A2(n12843), .ZN(n12840) );
  NAND2_X1 U9266 ( .A1(n12717), .A2(n12716), .ZN(n12715) );
  NAND2_X1 U9267 ( .A1(n15188), .A2(n15187), .ZN(n15186) );
  INV_X1 U9268 ( .A(n15239), .ZN(n15231) );
  AND2_X1 U9269 ( .A1(n8729), .A2(n8739), .ZN(n15239) );
  INV_X2 U9270 ( .A(n8274), .ZN(n8345) );
  XNOR2_X1 U9271 ( .A(n11678), .B(n11441), .ZN(n11444) );
  NAND2_X1 U9272 ( .A1(n13818), .A2(n12045), .ZN(n6854) );
  NOR2_X2 U9273 ( .A1(n7261), .A2(n11954), .ZN(n13760) );
  NAND3_X2 U9274 ( .A1(n10435), .A2(n8159), .A3(n8158), .ZN(n8374) );
  NAND2_X1 U9275 ( .A1(n8327), .A2(n8762), .ZN(n11450) );
  NAND2_X1 U9276 ( .A1(n8231), .A2(n8740), .ZN(n6971) );
  NAND2_X1 U9277 ( .A1(n6977), .A2(n6975), .ZN(n12792) );
  NAND2_X1 U9278 ( .A1(n13328), .A2(n13334), .ZN(n13329) );
  NAND2_X1 U9279 ( .A1(n13458), .A2(n13665), .ZN(n13460) );
  AOI22_X1 U9280 ( .A1(n13788), .A2(n13787), .B1(n11986), .B2(n11985), .ZN(
        n13741) );
  NOR2_X2 U9281 ( .A1(n13713), .A2(n11949), .ZN(n11953) );
  NAND2_X1 U9282 ( .A1(n6698), .A2(n6696), .ZN(P1_U3214) );
  NAND2_X1 U9283 ( .A1(n12047), .A2(n14488), .ZN(n6698) );
  INV_X1 U9284 ( .A(n14594), .ZN(n10667) );
  NAND2_X1 U9285 ( .A1(n12262), .A2(n12261), .ZN(n13923) );
  NAND2_X1 U9286 ( .A1(n11440), .A2(n11439), .ZN(n11678) );
  INV_X1 U9287 ( .A(n7499), .ZN(n6713) );
  INV_X1 U9288 ( .A(n6888), .ZN(n7670) );
  NAND2_X1 U9290 ( .A1(n7502), .A2(n6711), .ZN(n7624) );
  AND2_X2 U9291 ( .A1(n7375), .A2(n7378), .ZN(n7050) );
  AND4_X2 U9292 ( .A1(n7704), .A2(n7569), .A3(n7568), .A4(n7567), .ZN(n7375)
         );
  NAND2_X1 U9293 ( .A1(n10818), .A2(n10817), .ZN(n10824) );
  NAND2_X1 U9294 ( .A1(n7935), .A2(n10344), .ZN(n8060) );
  NOR2_X2 U9295 ( .A1(n7377), .A2(n7051), .ZN(n7935) );
  NAND2_X1 U9296 ( .A1(n10696), .A2(n10695), .ZN(n10818) );
  XNOR2_X1 U9297 ( .A(n6854), .B(n12046), .ZN(n12047) );
  NAND2_X1 U9298 ( .A1(n8122), .A2(n8131), .ZN(n8125) );
  NAND2_X1 U9299 ( .A1(n14580), .A2(n14581), .ZN(n14579) );
  INV_X1 U9300 ( .A(n14575), .ZN(n6702) );
  NOR2_X2 U9301 ( .A1(n11953), .A2(n11952), .ZN(n11954) );
  NAND3_X1 U9302 ( .A1(n11263), .A2(n11059), .A3(n11268), .ZN(n7242) );
  NAND2_X1 U9303 ( .A1(n10045), .A2(n9746), .ZN(n6710) );
  NAND2_X1 U9304 ( .A1(n6713), .A2(n6712), .ZN(n6711) );
  INV_X1 U9305 ( .A(SI_1_), .ZN(n6712) );
  OAI21_X1 U9306 ( .B1(n7503), .B2(n6715), .A(n6714), .ZN(n7499) );
  NAND2_X1 U9307 ( .A1(n7648), .A2(n7505), .ZN(n7651) );
  OAI21_X1 U9308 ( .B1(n11265), .B2(n7243), .A(n11275), .ZN(n7241) );
  INV_X1 U9309 ( .A(n14825), .ZN(n7220) );
  NAND2_X1 U9310 ( .A1(n7791), .A2(n7528), .ZN(n7805) );
  NAND2_X1 U9311 ( .A1(n7412), .A2(n7410), .ZN(n7769) );
  NAND2_X1 U9312 ( .A1(n7278), .A2(n7279), .ZN(n12380) );
  NOR2_X2 U9313 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n9046) );
  OAI211_X1 U9314 ( .C1(n13366), .C2(n6727), .A(n6723), .B(n7101), .ZN(n13325)
         );
  NAND2_X1 U9315 ( .A1(n6729), .A2(n6635), .ZN(n9515) );
  NAND2_X1 U9316 ( .A1(n9510), .A2(n6732), .ZN(n6729) );
  NAND3_X1 U9317 ( .A1(n6753), .A2(n6752), .A3(n6751), .ZN(n6750) );
  NAND2_X1 U9318 ( .A1(n13548), .A2(n14972), .ZN(n6751) );
  NAND2_X1 U9319 ( .A1(n9363), .A2(n6759), .ZN(n6758) );
  NAND2_X1 U9320 ( .A1(n11661), .A2(n9285), .ZN(n6771) );
  INV_X1 U9321 ( .A(n13486), .ZN(n13487) );
  INV_X1 U9322 ( .A(n10959), .ZN(n14975) );
  NAND2_X1 U9323 ( .A1(n14975), .A2(n13203), .ZN(n6774) );
  NAND3_X1 U9324 ( .A1(n13544), .A2(n6776), .A3(n13543), .ZN(n13642) );
  MUX2_X1 U9325 ( .A(n10079), .B(P2_REG1_REG_2__SCAN_IN), .S(n14853), .Z(
        n14851) );
  MUX2_X1 U9326 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9110), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n9112) );
  NAND2_X1 U9327 ( .A1(n10460), .A2(n6552), .ZN(n6796) );
  NAND3_X1 U9328 ( .A1(n6803), .A2(n6802), .A3(n6801), .ZN(n6800) );
  OAI21_X1 U9329 ( .B1(n6670), .B2(n10460), .A(n6552), .ZN(n10482) );
  AOI21_X1 U9330 ( .B1(n15062), .B2(n6807), .A(n6806), .ZN(n6805) );
  AND2_X1 U9331 ( .A1(n12668), .A2(n14431), .ZN(n6816) );
  NAND2_X1 U9332 ( .A1(n8430), .A2(n7363), .ZN(n8182) );
  NAND2_X1 U9333 ( .A1(n9573), .A2(n9572), .ZN(n6820) );
  OR2_X1 U9334 ( .A1(n9572), .A2(n9573), .ZN(n6818) );
  NAND3_X1 U9335 ( .A1(n9551), .A2(n9550), .A3(n9565), .ZN(n9564) );
  OAI21_X1 U9336 ( .B1(n6823), .B2(n9712), .A(n6824), .ZN(n7471) );
  OR2_X1 U9337 ( .A1(n9711), .A2(n6826), .ZN(n6823) );
  INV_X1 U9338 ( .A(n9715), .ZN(n6827) );
  NAND2_X1 U9339 ( .A1(n9700), .A2(n6830), .ZN(n6829) );
  NAND2_X1 U9340 ( .A1(n9053), .A2(n6837), .ZN(n6836) );
  INV_X1 U9341 ( .A(n9478), .ZN(n6840) );
  NAND2_X1 U9342 ( .A1(n6842), .A2(n6843), .ZN(n9634) );
  NAND4_X1 U9343 ( .A1(n14332), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(n6850), .A4(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n6849) );
  NAND4_X1 U9344 ( .A1(n7498), .A2(n6853), .A3(P3_ADDR_REG_19__SCAN_IN), .A4(
        n6852), .ZN(n6851) );
  NAND2_X1 U9345 ( .A1(n13760), .A2(n6859), .ZN(n6857) );
  NAND2_X1 U9346 ( .A1(n7671), .A2(n6864), .ZN(n6865) );
  MUX2_X1 U9347 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n9854), .Z(n6869) );
  MUX2_X1 U9348 ( .A(n9969), .B(P1_REG1_REG_1__SCAN_IN), .S(n13868), .Z(n13864) );
  NAND2_X1 U9349 ( .A1(n7680), .A2(n7679), .ZN(n7682) );
  NAND2_X1 U9350 ( .A1(n7439), .A2(n6550), .ZN(n6893) );
  NAND2_X1 U9351 ( .A1(n14001), .A2(n6643), .ZN(n6899) );
  CLKBUF_X1 U9352 ( .A(n6899), .Z(n6898) );
  INV_X1 U9353 ( .A(n6898), .ZN(n13980) );
  NAND2_X1 U9354 ( .A1(n6904), .A2(n14716), .ZN(n8903) );
  OAI21_X1 U9355 ( .B1(n6904), .B2(n6903), .A(n6902), .ZN(n8920) );
  AOI21_X1 U9356 ( .B1(n8902), .B2(n14691), .A(n14701), .ZN(n6902) );
  INV_X1 U9357 ( .A(n11166), .ZN(n6909) );
  AND3_X2 U9358 ( .A1(n9113), .A2(n9114), .A3(n7486), .ZN(n11131) );
  NOR2_X2 U9359 ( .A1(n13492), .A2(n13477), .ZN(n13458) );
  NOR2_X2 U9360 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n6936) );
  AND3_X2 U9361 ( .A1(n6937), .A2(n6936), .A3(n7775), .ZN(n7374) );
  NOR2_X2 U9362 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n6937) );
  AND2_X2 U9363 ( .A1(n7374), .A2(n7372), .ZN(n7049) );
  AND3_X2 U9364 ( .A1(n6938), .A2(n7566), .A3(n7266), .ZN(n7372) );
  NOR2_X2 U9365 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n6938) );
  NOR2_X2 U9367 ( .A1(n13956), .A2(n14137), .ZN(n6944) );
  NOR2_X2 U9368 ( .A1(n13986), .A2(n14147), .ZN(n6946) );
  NAND2_X1 U9369 ( .A1(n10461), .A2(n6953), .ZN(n6951) );
  NAND2_X1 U9370 ( .A1(n15163), .A2(n14389), .ZN(n6955) );
  NAND3_X1 U9371 ( .A1(n6956), .A2(n6958), .A3(n6955), .ZN(n14382) );
  AND4_X2 U9372 ( .A1(n6956), .A2(n6958), .A3(n6955), .A4(
        P3_REG2_REG_15__SCAN_IN), .ZN(n14381) );
  NOR2_X1 U9373 ( .A1(n14411), .A2(n6668), .ZN(n12583) );
  NAND3_X1 U9374 ( .A1(n6961), .A2(n6962), .A3(n6960), .ZN(n14424) );
  NAND4_X1 U9375 ( .A1(n6961), .A2(n6962), .A3(n6960), .A4(
        P3_REG2_REG_17__SCAN_IN), .ZN(n6963) );
  INV_X1 U9376 ( .A(n6963), .ZN(n14426) );
  INV_X1 U9377 ( .A(n6967), .ZN(n15027) );
  INV_X1 U9378 ( .A(n6965), .ZN(n15025) );
  NAND2_X1 U9379 ( .A1(n12567), .A2(n15014), .ZN(n6968) );
  NAND2_X1 U9380 ( .A1(n6971), .A2(n8248), .ZN(n8249) );
  XNOR2_X1 U9381 ( .A(n6971), .B(n11018), .ZN(n11022) );
  INV_X1 U9382 ( .A(n6972), .ZN(n13012) );
  NOR2_X2 U9383 ( .A1(n8179), .A2(n6973), .ZN(n6972) );
  NAND2_X1 U9384 ( .A1(n12822), .A2(n6978), .ZN(n6977) );
  INV_X1 U9385 ( .A(n8160), .ZN(n6983) );
  NOR2_X2 U9386 ( .A1(n8374), .A2(n6625), .ZN(n6982) );
  OAI21_X1 U9387 ( .B1(SI_2_), .B2(n8345), .A(n8189), .ZN(n6985) );
  NAND2_X2 U9388 ( .A1(n6986), .A2(n8178), .ZN(n15258) );
  NAND4_X1 U9389 ( .A1(n6984), .A2(n6986), .A3(n8190), .A4(n8178), .ZN(n8739)
         );
  NAND2_X1 U9390 ( .A1(n15258), .A2(n15235), .ZN(n8729) );
  NAND2_X1 U9391 ( .A1(n12783), .A2(n6583), .ZN(n6987) );
  NAND2_X1 U9392 ( .A1(n6987), .A2(n6988), .ZN(n12760) );
  NAND2_X1 U9393 ( .A1(n6994), .A2(n6996), .ZN(n8459) );
  OAI21_X1 U9394 ( .B1(n11514), .B2(n8364), .A(n8365), .ZN(n14449) );
  NAND2_X1 U9395 ( .A1(n14448), .A2(n7012), .ZN(n7011) );
  NAND2_X1 U9396 ( .A1(n8356), .A2(n7030), .ZN(n7027) );
  NAND2_X1 U9397 ( .A1(n8463), .A2(n7036), .ZN(n7033) );
  NAND2_X1 U9398 ( .A1(n7033), .A2(n7034), .ZN(n8509) );
  OAI21_X1 U9399 ( .B1(n8297), .B2(n7043), .A(n7040), .ZN(n8338) );
  NAND2_X1 U9400 ( .A1(n8619), .A2(n8618), .ZN(n8631) );
  NAND2_X1 U9401 ( .A1(n7376), .A2(n7372), .ZN(n7051) );
  NAND2_X1 U9402 ( .A1(n7050), .A2(n7374), .ZN(n7377) );
  NAND2_X1 U9403 ( .A1(n8098), .A2(n6549), .ZN(n7053) );
  NAND2_X1 U9404 ( .A1(n11532), .A2(n7063), .ZN(n7060) );
  NAND2_X1 U9405 ( .A1(n7060), .A2(n7061), .ZN(n11623) );
  AOI21_X2 U9406 ( .B1(n14711), .B2(n7067), .A(n7066), .ZN(n14688) );
  NAND2_X1 U9407 ( .A1(n14713), .A2(n14712), .ZN(n14711) );
  NAND2_X1 U9408 ( .A1(n7073), .A2(n7071), .ZN(n14000) );
  NAND2_X1 U9409 ( .A1(n7074), .A2(n7075), .ZN(n14105) );
  NAND2_X1 U9410 ( .A1(n8095), .A2(n7076), .ZN(n7074) );
  NAND2_X2 U9411 ( .A1(n8100), .A2(n8099), .ZN(n14055) );
  OAI21_X2 U9412 ( .B1(n13991), .B2(n7082), .A(n7080), .ZN(n13945) );
  NOR2_X2 U9413 ( .A1(n13940), .A2(n13941), .ZN(n13939) );
  NAND2_X1 U9414 ( .A1(n7090), .A2(n7092), .ZN(n9510) );
  NAND2_X1 U9415 ( .A1(n13502), .A2(n7093), .ZN(n7090) );
  OAI21_X1 U9416 ( .B1(n13396), .B2(n7112), .A(n7110), .ZN(n13366) );
  OAI21_X1 U9417 ( .B1(n13396), .B2(n9519), .A(n9520), .ZN(n13380) );
  NAND3_X1 U9418 ( .A1(n7469), .A2(n9327), .A3(n9069), .ZN(n9057) );
  NAND3_X1 U9419 ( .A1(n7469), .A2(n9327), .A3(n7115), .ZN(n13684) );
  NAND2_X1 U9420 ( .A1(n9485), .A2(n9484), .ZN(n10534) );
  NAND2_X1 U9421 ( .A1(n9518), .A2(n9517), .ZN(n13396) );
  NAND2_X1 U9422 ( .A1(n9515), .A2(n9514), .ZN(n13411) );
  NAND2_X1 U9423 ( .A1(n11360), .A2(n7204), .ZN(n11359) );
  NAND2_X1 U9424 ( .A1(n9524), .A2(n9774), .ZN(n13312) );
  NAND2_X1 U9425 ( .A1(n9483), .A2(n9482), .ZN(n10555) );
  INV_X1 U9426 ( .A(n8857), .ZN(n8858) );
  NAND2_X1 U9427 ( .A1(n8606), .A2(n8605), .ZN(n8617) );
  NAND2_X1 U9428 ( .A1(n8579), .A2(n8578), .ZN(n8580) );
  NAND2_X1 U9429 ( .A1(n8105), .A2(n13982), .ZN(n13991) );
  NAND2_X4 U9430 ( .A1(n7676), .A2(n6533), .ZN(n7673) );
  XNOR2_X1 U9431 ( .A(n13859), .B(n14724), .ZN(n14714) );
  NAND2_X1 U9432 ( .A1(n8604), .A2(n8603), .ZN(n8606) );
  XNOR2_X1 U9433 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8209) );
  NAND2_X1 U9434 ( .A1(n11425), .A2(n9494), .ZN(n11360) );
  INV_X1 U9435 ( .A(n10554), .ZN(n9778) );
  NAND2_X1 U9436 ( .A1(n7116), .A2(n13915), .ZN(n12247) );
  NAND2_X1 U9437 ( .A1(n7116), .A2(n12255), .ZN(n12263) );
  NAND2_X1 U9438 ( .A1(n13915), .A2(n14227), .ZN(n7276) );
  NAND2_X1 U9439 ( .A1(n12248), .A2(n7116), .ZN(n10048) );
  NAND2_X1 U9440 ( .A1(n8117), .A2(n7116), .ZN(n8905) );
  NAND2_X1 U9441 ( .A1(n7135), .A2(n7138), .ZN(n12206) );
  NAND3_X1 U9442 ( .A1(n12202), .A2(n7136), .A3(n12201), .ZN(n7135) );
  NAND3_X1 U9443 ( .A1(n12093), .A2(n12227), .A3(n7141), .ZN(n7140) );
  NAND2_X1 U9444 ( .A1(n8057), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8058) );
  NAND2_X1 U9445 ( .A1(n12129), .A2(n7146), .ZN(n7143) );
  OAI21_X1 U9446 ( .B1(n12129), .B2(n6551), .A(n7146), .ZN(n12133) );
  NAND2_X1 U9447 ( .A1(n7143), .A2(n7144), .ZN(n12132) );
  NAND2_X1 U9448 ( .A1(n7151), .A2(n7149), .ZN(n12199) );
  NAND2_X1 U9449 ( .A1(n7155), .A2(n7156), .ZN(n12186) );
  AOI21_X1 U9450 ( .B1(n7160), .B2(n7163), .A(n7158), .ZN(n7157) );
  INV_X1 U9451 ( .A(n12234), .ZN(n7174) );
  NAND2_X1 U9452 ( .A1(n9244), .A2(n7184), .ZN(n7181) );
  NAND2_X1 U9453 ( .A1(n7181), .A2(n7182), .ZN(n11661) );
  NAND2_X1 U9454 ( .A1(n7192), .A2(n7191), .ZN(n11302) );
  NAND3_X1 U9455 ( .A1(n11114), .A2(n9177), .A3(n11288), .ZN(n7192) );
  NAND2_X1 U9456 ( .A1(n11114), .A2(n9177), .ZN(n7194) );
  OAI21_X1 U9457 ( .B1(n9325), .B2(n7197), .A(n7196), .ZN(n13448) );
  INV_X1 U9458 ( .A(n9217), .ZN(n11420) );
  NAND2_X1 U9459 ( .A1(n9217), .A2(n9782), .ZN(n7200) );
  NAND2_X2 U9460 ( .A1(n9142), .A2(n9874), .ZN(n9133) );
  NAND2_X1 U9461 ( .A1(n7651), .A2(n7652), .ZN(n9875) );
  NAND2_X1 U9462 ( .A1(n13071), .A2(n7224), .ZN(n7223) );
  NAND2_X1 U9463 ( .A1(n7223), .A2(n7221), .ZN(n13052) );
  AOI21_X1 U9464 ( .B1(n11714), .B2(n7231), .A(n7230), .ZN(n7229) );
  NAND2_X1 U9465 ( .A1(n13179), .A2(n7234), .ZN(n13091) );
  OR2_X2 U9466 ( .A1(n13161), .A2(n7238), .ZN(n7237) );
  NOR2_X2 U9467 ( .A1(n13163), .A2(n13162), .ZN(n13161) );
  AND2_X1 U9468 ( .A1(n10953), .A2(n10952), .ZN(n7239) );
  NAND2_X1 U9469 ( .A1(n7242), .A2(n7240), .ZN(n11557) );
  NAND2_X1 U9470 ( .A1(n9477), .A2(n13276), .ZN(n10406) );
  OAI211_X1 U9471 ( .C1(n13818), .C2(n7259), .A(n7256), .B(n7254), .ZN(n12346)
         );
  OAI22_X1 U9472 ( .A1(n7258), .A2(n7255), .B1(n12339), .B2(n7260), .ZN(n7254)
         );
  NOR2_X1 U9473 ( .A1(n12339), .A2(n12046), .ZN(n7255) );
  NAND2_X1 U9474 ( .A1(n13818), .A2(n7257), .ZN(n7256) );
  NOR2_X1 U9475 ( .A1(n7258), .A2(n12339), .ZN(n7257) );
  NAND2_X1 U9476 ( .A1(n12046), .A2(n12339), .ZN(n7259) );
  AND2_X2 U9477 ( .A1(n7263), .A2(n7262), .ZN(n7261) );
  NAND2_X1 U9478 ( .A1(n12450), .A2(n6546), .ZN(n7278) );
  INV_X1 U9479 ( .A(n12450), .ZN(n7282) );
  NOR2_X1 U9480 ( .A1(n12375), .A2(n12376), .ZN(n7287) );
  NAND2_X1 U9481 ( .A1(n14369), .A2(n7290), .ZN(n7289) );
  NAND3_X1 U9482 ( .A1(n7304), .A2(n8988), .A3(n8714), .ZN(n10630) );
  NAND2_X1 U9483 ( .A1(n12528), .A2(n12401), .ZN(n12434) );
  OAI211_X1 U9484 ( .C1(n12528), .C2(n7310), .A(n7307), .B(n7305), .ZN(n12412)
         );
  NAND2_X1 U9485 ( .A1(n12528), .A2(n7306), .ZN(n7305) );
  NOR2_X1 U9486 ( .A1(n7308), .A2(n12404), .ZN(n7306) );
  OAI22_X1 U9487 ( .A1(n7309), .A2(n7308), .B1(n12404), .B2(n7311), .ZN(n7307)
         );
  NOR2_X1 U9488 ( .A1(n12404), .A2(n12435), .ZN(n7309) );
  NAND2_X1 U9489 ( .A1(n7313), .A2(n12491), .ZN(n12392) );
  AOI21_X2 U9490 ( .B1(n12712), .B2(n8969), .A(n8968), .ZN(n12703) );
  OAI21_X2 U9491 ( .B1(n12725), .B2(n12726), .A(n8967), .ZN(n12712) );
  NAND2_X1 U9492 ( .A1(n11396), .A2(n7327), .ZN(n7324) );
  NAND2_X1 U9493 ( .A1(n7324), .A2(n7325), .ZN(n11518) );
  NAND2_X1 U9494 ( .A1(n12795), .A2(n7334), .ZN(n7331) );
  NAND2_X1 U9495 ( .A1(n7331), .A2(n7332), .ZN(n12775) );
  NAND2_X1 U9496 ( .A1(n8963), .A2(n7341), .ZN(n7340) );
  INV_X1 U9497 ( .A(n12762), .ZN(n7342) );
  OAI21_X1 U9498 ( .B1(n12832), .B2(n7346), .A(n7343), .ZN(n12802) );
  NAND2_X1 U9499 ( .A1(n7352), .A2(n7350), .ZN(n15191) );
  NAND2_X1 U9500 ( .A1(n11017), .A2(n8929), .ZN(n15204) );
  INV_X1 U9501 ( .A(n8929), .ZN(n7354) );
  OAI21_X2 U9502 ( .B1(n8937), .B2(n7357), .A(n7355), .ZN(n11831) );
  NAND2_X1 U9503 ( .A1(n8937), .A2(n8936), .ZN(n14450) );
  INV_X1 U9504 ( .A(n8936), .ZN(n7362) );
  AND2_X1 U9505 ( .A1(n8430), .A2(n8161), .ZN(n8450) );
  NAND2_X1 U9506 ( .A1(n8983), .A2(n8982), .ZN(n12690) );
  NAND2_X1 U9507 ( .A1(n11533), .A2(n7803), .ZN(n14514) );
  INV_X1 U9508 ( .A(n11535), .ZN(n7370) );
  INV_X1 U9509 ( .A(n7377), .ZN(n7906) );
  NAND2_X1 U9510 ( .A1(n14096), .A2(n7382), .ZN(n7379) );
  NAND2_X1 U9511 ( .A1(n11624), .A2(n7393), .ZN(n7392) );
  NAND2_X1 U9512 ( .A1(n11847), .A2(n6638), .ZN(n14495) );
  OAI21_X1 U9513 ( .B1(n11076), .B2(n7697), .A(n7698), .ZN(n14690) );
  NAND2_X1 U9514 ( .A1(n7576), .A2(n7407), .ZN(n7586) );
  NAND2_X1 U9515 ( .A1(n7576), .A2(n7575), .ZN(n7578) );
  INV_X1 U9516 ( .A(n7586), .ZN(n7584) );
  NAND2_X1 U9517 ( .A1(n7750), .A2(n7408), .ZN(n11198) );
  OAI21_X1 U9518 ( .B1(n7733), .B2(n7415), .A(n7413), .ZN(n7753) );
  NAND2_X1 U9519 ( .A1(n7733), .A2(n7413), .ZN(n7412) );
  INV_X1 U9520 ( .A(n7977), .ZN(n7417) );
  AOI21_X2 U9521 ( .B1(n7980), .B2(n7420), .A(n7419), .ZN(n7416) );
  NAND2_X1 U9522 ( .A1(n7980), .A2(n7421), .ZN(n7418) );
  OAI21_X1 U9523 ( .B1(n7789), .B2(n7426), .A(n7425), .ZN(n7822) );
  NAND2_X1 U9524 ( .A1(n7956), .A2(n7433), .ZN(n7431) );
  NAND2_X1 U9525 ( .A1(n7956), .A2(n7555), .ZN(n7432) );
  NAND2_X1 U9526 ( .A1(n7835), .A2(n7834), .ZN(n7442) );
  NAND3_X1 U9527 ( .A1(n9048), .A2(n9047), .A3(n9046), .ZN(n9202) );
  AOI21_X1 U9528 ( .B1(n9592), .B2(n9591), .A(n9590), .ZN(n9594) );
  NOR2_X1 U9529 ( .A1(n9606), .A2(n9605), .ZN(n9607) );
  NAND2_X1 U9530 ( .A1(n9657), .A2(n7455), .ZN(n7453) );
  NAND2_X1 U9531 ( .A1(n9658), .A2(n7455), .ZN(n7454) );
  NAND3_X1 U9532 ( .A1(n7454), .A2(n7453), .A3(n7452), .ZN(n9686) );
  AND2_X1 U9533 ( .A1(n7458), .A2(n9680), .ZN(n7457) );
  AND2_X1 U9534 ( .A1(n9614), .A2(n9613), .ZN(n7465) );
  NAND2_X1 U9535 ( .A1(n7471), .A2(n7472), .ZN(n9724) );
  OR2_X1 U9536 ( .A1(n11709), .A2(n11802), .ZN(n11710) );
  NAND2_X2 U9537 ( .A1(n8740), .A2(n8743), .ZN(n15219) );
  AND2_X1 U9538 ( .A1(n10067), .A2(n10066), .ZN(n10071) );
  INV_X4 U9539 ( .A(n10660), .ZN(n12035) );
  INV_X1 U9540 ( .A(n13861), .ZN(n7640) );
  OR2_X1 U9541 ( .A1(n9455), .A2(n9454), .ZN(n9457) );
  CLKBUF_X1 U9542 ( .A(n8072), .Z(n12062) );
  XNOR2_X1 U9543 ( .A(n9015), .B(n9016), .ZN(n12697) );
  NAND2_X1 U9544 ( .A1(n12361), .A2(n12360), .ZN(n12365) );
  NAND2_X1 U9545 ( .A1(n12320), .A2(n12318), .ZN(n12319) );
  NAND2_X1 U9546 ( .A1(n11343), .A2(n9498), .ZN(n11603) );
  XNOR2_X1 U9547 ( .A(n9528), .B(n9527), .ZN(n9540) );
  AOI22_X2 U9548 ( .A1(n12521), .A2(n12520), .B1(n12373), .B2(n12833), .ZN(
        n12450) );
  AND2_X2 U9549 ( .A1(n12083), .A2(n12082), .ZN(n12104) );
  XNOR2_X1 U9550 ( .A(n7552), .B(SI_20_), .ZN(n7945) );
  NAND2_X1 U9551 ( .A1(n7945), .A2(n7551), .ZN(n7554) );
  NAND2_X1 U9552 ( .A1(n7545), .A2(SI_18_), .ZN(n7546) );
  OR2_X1 U9553 ( .A1(n8053), .A2(n8113), .ZN(n8054) );
  OR2_X1 U9554 ( .A1(n13544), .A2(n13517), .ZN(n9549) );
  INV_X1 U9555 ( .A(n13693), .ZN(n9060) );
  AND2_X1 U9556 ( .A1(n12419), .A2(n12065), .ZN(n10896) );
  NAND2_X1 U9557 ( .A1(n9136), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n9108) );
  NAND2_X1 U9558 ( .A1(n7586), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7588) );
  NAND2_X1 U9559 ( .A1(n8976), .A2(n15262), .ZN(n8983) );
  MUX2_X2 U9560 ( .A(n9030), .B(n9029), .S(n15318), .Z(n9032) );
  OAI211_X1 U9561 ( .C1(n8679), .C2(n12965), .A(n8552), .B(n8551), .ZN(n12796)
         );
  NAND2_X1 U9562 ( .A1(n8016), .A2(n11696), .ZN(n8017) );
  OAI21_X1 U9563 ( .B1(n8016), .B2(n11696), .A(n8015), .ZN(n8018) );
  XNOR2_X1 U9564 ( .A(n8016), .B(n8000), .ZN(n13702) );
  NOR2_X1 U9565 ( .A1(n9818), .A2(n9817), .ZN(n9841) );
  INV_X1 U9566 ( .A(n12273), .ZN(n10183) );
  OR2_X1 U9567 ( .A1(n12564), .A2(n15254), .ZN(n15230) );
  INV_X1 U9568 ( .A(n8172), .ZN(n8173) );
  OR2_X1 U9569 ( .A1(n8651), .A2(n12437), .ZN(n8627) );
  NAND2_X1 U9570 ( .A1(n15232), .A2(n10634), .ZN(n7476) );
  AND2_X1 U9571 ( .A1(n8395), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7477) );
  OR2_X1 U9572 ( .A1(n8546), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n7478) );
  INV_X1 U9573 ( .A(n11578), .ZN(n9272) );
  INV_X1 U9574 ( .A(n13489), .ZN(n13508) );
  INV_X1 U9575 ( .A(n11843), .ZN(n14124) );
  AND2_X1 U9576 ( .A1(n11767), .A2(n11766), .ZN(n7479) );
  AND2_X1 U9577 ( .A1(n11818), .A2(n14454), .ZN(n7480) );
  OR4_X1 U9578 ( .A1(n15243), .A2(n10641), .A3(n12328), .A4(n10626), .ZN(n7482) );
  OR2_X1 U9579 ( .A1(n12364), .A2(n12363), .ZN(n7484) );
  AND2_X1 U9580 ( .A1(n13195), .A2(n13490), .ZN(n7485) );
  INV_X1 U9581 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n13011) );
  AND2_X1 U9582 ( .A1(n8975), .A2(n9023), .ZN(n15249) );
  INV_X1 U9583 ( .A(n10154), .ZN(n7639) );
  INV_X1 U9584 ( .A(n11152), .ZN(n8862) );
  OR2_X1 U9585 ( .A1(n9142), .A2(n10097), .ZN(n7486) );
  XOR2_X1 U9586 ( .A(n13375), .B(n6468), .Z(n7487) );
  INV_X1 U9587 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7723) );
  INV_X1 U9588 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n8403) );
  AND3_X1 U9589 ( .A1(n11312), .A2(n11311), .A3(n11467), .ZN(n7488) );
  OR2_X1 U9590 ( .A1(n13545), .A2(n13467), .ZN(n7490) );
  AND2_X1 U9591 ( .A1(n13733), .A2(n13731), .ZN(n7491) );
  AND2_X1 U9592 ( .A1(n8120), .A2(n8119), .ZN(n7492) );
  INV_X1 U9593 ( .A(n13401), .ZN(n13414) );
  AND2_X1 U9594 ( .A1(n13526), .A2(n13198), .ZN(n7493) );
  OR2_X1 U9595 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n7494) );
  NOR3_X1 U9596 ( .A1(n14536), .A2(n14535), .A3(n14534), .ZN(n7496) );
  NOR3_X1 U9597 ( .A1(n14536), .A2(n14513), .A3(n14512), .ZN(n7497) );
  INV_X1 U9598 ( .A(n12094), .ZN(n12096) );
  INV_X1 U9599 ( .A(n12088), .ZN(n12099) );
  MUX2_X1 U9600 ( .A(n12085), .B(n12084), .S(n12227), .Z(n12103) );
  OAI21_X1 U9601 ( .B1(n11256), .B2(n9819), .A(n9612), .ZN(n9613) );
  INV_X1 U9602 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9044) );
  AND2_X1 U9603 ( .A1(n12872), .A2(n12438), .ZN(n8970) );
  INV_X1 U9604 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8165) );
  INV_X1 U9605 ( .A(n13404), .ZN(n9542) );
  INV_X1 U9606 ( .A(n7899), .ZN(n7544) );
  INV_X1 U9607 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n8308) );
  INV_X1 U9608 ( .A(n9016), .ZN(n8973) );
  INV_X1 U9609 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8154) );
  OR2_X1 U9610 ( .A1(n14953), .A2(n10401), .ZN(n10416) );
  INV_X1 U9611 ( .A(n9368), .ZN(n9036) );
  INV_X1 U9612 ( .A(n9378), .ZN(n9037) );
  NOR2_X1 U9613 ( .A1(n9305), .A2(n9304), .ZN(n9303) );
  NAND2_X1 U9614 ( .A1(n12091), .A2(n12094), .ZN(n10149) );
  OR2_X1 U9615 ( .A1(n11412), .A2(n11413), .ZN(n11410) );
  INV_X1 U9616 ( .A(n10806), .ZN(n10803) );
  OR2_X1 U9617 ( .A1(n8651), .A2(n12701), .ZN(n8643) );
  OAI22_X1 U9618 ( .A1(n8980), .A2(n15243), .B1(n12682), .B2(n11149), .ZN(
        n8981) );
  NOR2_X1 U9619 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(n8585), .ZN(n8596) );
  INV_X1 U9620 ( .A(n12821), .ZN(n12823) );
  NAND2_X1 U9621 ( .A1(n9913), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8334) );
  OR2_X1 U9622 ( .A1(n13039), .A2(n6567), .ZN(n13040) );
  INV_X1 U9623 ( .A(n14814), .ZN(n10942) );
  OR2_X1 U9624 ( .A1(n10932), .A2(n10897), .ZN(n10408) );
  OR2_X1 U9626 ( .A1(n11701), .A2(n11703), .ZN(n11698) );
  OR2_X1 U9627 ( .A1(n9390), .A2(n9039), .ZN(n9401) );
  OR2_X1 U9628 ( .A1(n9388), .A2(n13129), .ZN(n9390) );
  NAND2_X1 U9629 ( .A1(n9035), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n9366) );
  OR2_X1 U9630 ( .A1(n13225), .A2(n13224), .ZN(n13226) );
  AND2_X1 U9631 ( .A1(n6841), .A2(n9843), .ZN(n10411) );
  INV_X1 U9632 ( .A(n13192), .ZN(n9350) );
  NAND2_X1 U9633 ( .A1(n13489), .A2(n9541), .ZN(n13492) );
  AND2_X1 U9634 ( .A1(n9251), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n9266) );
  OR2_X1 U9635 ( .A1(n9223), .A2(n9222), .ZN(n9235) );
  NAND2_X1 U9636 ( .A1(n9171), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9193) );
  INV_X1 U9637 ( .A(n11980), .ZN(n11983) );
  NAND2_X1 U9638 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n7593), .ZN(n7987) );
  INV_X1 U9639 ( .A(n12301), .ZN(n8887) );
  OR2_X1 U9640 ( .A1(n7856), .A2(n7855), .ZN(n7873) );
  NOR2_X1 U9641 ( .A1(n7724), .A2(n7723), .ZN(n7741) );
  INV_X1 U9642 ( .A(n10149), .ZN(n12275) );
  INV_X1 U9643 ( .A(n8121), .ZN(n8122) );
  OR2_X1 U9644 ( .A1(n7552), .A2(n10754), .ZN(n7553) );
  NOR2_X1 U9645 ( .A1(n14270), .A2(n14269), .ZN(n14256) );
  AND2_X1 U9646 ( .A1(n8522), .A2(n8521), .ZN(n8536) );
  AND2_X1 U9647 ( .A1(n12467), .A2(n12391), .ZN(n12492) );
  AND2_X1 U9648 ( .A1(n8416), .A2(n8415), .ZN(n8436) );
  INV_X1 U9649 ( .A(n12545), .ZN(n12507) );
  AND4_X1 U9650 ( .A1(n8645), .A2(n8644), .A3(n8643), .A4(n8642), .ZN(n8980)
         );
  AND4_X1 U9651 ( .A1(n8458), .A2(n8457), .A3(n8456), .A4(n8455), .ZN(n12476)
         );
  OR2_X1 U9652 ( .A1(n8679), .A2(n8191), .ZN(n8197) );
  INV_X1 U9653 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n11328) );
  INV_X1 U9654 ( .A(n8981), .ZN(n8982) );
  AND2_X1 U9655 ( .A1(n8436), .A2(n8435), .ZN(n8470) );
  AND2_X1 U9656 ( .A1(n10607), .A2(n9910), .ZN(n10619) );
  AND2_X1 U9657 ( .A1(n12694), .A2(n12888), .ZN(n8984) );
  INV_X1 U9658 ( .A(n15249), .ZN(n15262) );
  AND2_X1 U9659 ( .A1(n8777), .A2(n8778), .ZN(n11615) );
  INV_X1 U9660 ( .A(n15205), .ZN(n15202) );
  NAND2_X1 U9661 ( .A1(n10964), .A2(n9022), .ZN(n15253) );
  AND2_X1 U9662 ( .A1(n8443), .A2(n8425), .ZN(n8426) );
  AND2_X1 U9663 ( .A1(n8385), .A2(n8379), .ZN(n8380) );
  AND2_X1 U9664 ( .A1(n13187), .A2(n13490), .ZN(n13041) );
  INV_X1 U9665 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n14820) );
  AND2_X1 U9666 ( .A1(n14954), .A2(n10402), .ZN(n10415) );
  OR2_X1 U9667 ( .A1(n9357), .A2(n13080), .ZN(n9359) );
  INV_X1 U9668 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n14905) );
  NAND2_X1 U9669 ( .A1(n13441), .A2(n9350), .ZN(n9351) );
  INV_X1 U9670 ( .A(n9787), .ZN(n13447) );
  XNOR2_X1 U9671 ( .A(n13542), .B(n13181), .ZN(n9794) );
  AND2_X1 U9672 ( .A1(n12034), .A2(n12033), .ZN(n13749) );
  AND2_X1 U9673 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n7708) );
  INV_X1 U9674 ( .A(n10681), .ZN(n10688) );
  INV_X1 U9675 ( .A(n12298), .ZN(n8113) );
  INV_X1 U9676 ( .A(n14074), .ZN(n14064) );
  INV_X1 U9677 ( .A(n14498), .ZN(n14694) );
  NAND2_X2 U9678 ( .A1(n8072), .A2(n14609), .ZN(n7676) );
  XNOR2_X1 U9679 ( .A(n14025), .B(n14032), .ZN(n14027) );
  INV_X1 U9680 ( .A(n12281), .ZN(n11201) );
  OR2_X1 U9681 ( .A1(n9904), .A2(n8148), .ZN(n10058) );
  XNOR2_X1 U9682 ( .A(n7533), .B(n9915), .ZN(n7834) );
  AOI22_X1 U9683 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14244), .B1(n14296), .B2(
        n14243), .ZN(n14245) );
  AND2_X1 U9684 ( .A1(n8869), .A2(n8868), .ZN(n8874) );
  OR2_X1 U9685 ( .A1(n8346), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8367) );
  INV_X1 U9686 ( .A(n11724), .ZN(n11731) );
  NAND2_X1 U9687 ( .A1(n10799), .A2(n10798), .ZN(n10807) );
  NAND2_X1 U9688 ( .A1(n10618), .A2(n15268), .ZN(n12548) );
  OR2_X1 U9689 ( .A1(n8651), .A2(n12685), .ZN(n8683) );
  AND4_X1 U9690 ( .A1(n8575), .A2(n8574), .A3(n8573), .A4(n8572), .ZN(n8961)
         );
  AND4_X1 U9691 ( .A1(n8506), .A2(n8505), .A3(n8504), .A4(n8503), .ZN(n12807)
         );
  OR2_X1 U9692 ( .A1(n8651), .A2(n11525), .ZN(n8348) );
  OR2_X1 U9693 ( .A1(n10443), .A2(n10442), .ZN(n10446) );
  NOR2_X1 U9694 ( .A1(n10510), .A2(n15237), .ZN(n15227) );
  INV_X1 U9695 ( .A(n12907), .ZN(n12918) );
  OR2_X1 U9696 ( .A1(n9004), .A2(n9003), .ZN(n10507) );
  OR2_X1 U9697 ( .A1(n10642), .A2(n9026), .ZN(n9027) );
  INV_X1 U9698 ( .A(n15275), .ZN(n15312) );
  INV_X1 U9699 ( .A(n9022), .ZN(n10966) );
  INV_X1 U9700 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8692) );
  INV_X1 U9701 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8225) );
  INV_X1 U9702 ( .A(n14832), .ZN(n13174) );
  AND2_X1 U9703 ( .A1(n10415), .A2(n10414), .ZN(n13159) );
  OR2_X1 U9704 ( .A1(n10918), .A2(n10917), .ZN(n10919) );
  INV_X1 U9705 ( .A(n13133), .ZN(n14829) );
  INV_X1 U9706 ( .A(n14863), .ZN(n14932) );
  AND2_X1 U9707 ( .A1(n10109), .A2(n13701), .ZN(n14863) );
  AOI21_X1 U9708 ( .B1(n13541), .B2(n13529), .A(n9547), .ZN(n9548) );
  INV_X1 U9709 ( .A(n13630), .ZN(n13634) );
  NOR2_X1 U9710 ( .A1(n14955), .A2(n10542), .ZN(n10546) );
  INV_X1 U9711 ( .A(n13622), .ZN(n14982) );
  AND2_X1 U9712 ( .A1(n9848), .A2(n10090), .ZN(n10916) );
  AND2_X1 U9713 ( .A1(n9168), .A2(n9189), .ZN(n10102) );
  AND2_X1 U9714 ( .A1(n14592), .A2(n14761), .ZN(n13794) );
  AND2_X1 U9715 ( .A1(n10698), .A2(n10072), .ZN(n14592) );
  OR2_X1 U9716 ( .A1(n14618), .A2(n9977), .ZN(n13911) );
  INV_X1 U9717 ( .A(n13899), .ZN(n14649) );
  NAND2_X1 U9718 ( .A1(n8014), .A2(n8013), .ZN(n13946) );
  NAND2_X1 U9719 ( .A1(n10072), .A2(n8900), .ZN(n14719) );
  INV_X1 U9720 ( .A(n14103), .ZN(n14723) );
  AND2_X1 U9721 ( .A1(n9920), .A2(n12062), .ZN(n14498) );
  INV_X1 U9722 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n8897) );
  INV_X1 U9723 ( .A(n14797), .ZN(n14537) );
  NOR2_X1 U9724 ( .A1(n12263), .A2(n13915), .ZN(n14787) );
  AND3_X1 U9725 ( .A1(n10062), .A2(n10057), .A3(n10058), .ZN(n8907) );
  AND2_X1 U9726 ( .A1(n7776), .A2(n7792), .ZN(n10518) );
  INV_X1 U9727 ( .A(n9910), .ZN(n9931) );
  AND2_X1 U9728 ( .A1(n10617), .A2(n10616), .ZN(n14379) );
  NAND2_X1 U9729 ( .A1(n7482), .A2(n8876), .ZN(n8877) );
  INV_X1 U9730 ( .A(n12485), .ZN(n12855) );
  INV_X1 U9731 ( .A(n15054), .ZN(n15184) );
  NAND2_X1 U9732 ( .A1(n15273), .A2(n15209), .ZN(n12863) );
  AND2_X1 U9733 ( .A1(n11523), .A2(n11522), .ZN(n15315) );
  NAND2_X2 U9734 ( .A1(n10510), .A2(n15268), .ZN(n15273) );
  OR2_X1 U9735 ( .A1(n10507), .A2(n9013), .ZN(n15329) );
  INV_X1 U9736 ( .A(n12433), .ZN(n12937) );
  AND2_X1 U9737 ( .A1(n15315), .A2(n15314), .ZN(n15330) );
  AND2_X1 U9738 ( .A1(n9028), .A2(n9027), .ZN(n15316) );
  AND2_X1 U9739 ( .A1(n10606), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9910) );
  XNOR2_X1 U9740 ( .A(n8867), .B(n7366), .ZN(n11697) );
  INV_X1 U9741 ( .A(SI_13_), .ZN(n9915) );
  INV_X1 U9742 ( .A(SI_11_), .ZN(n9889) );
  INV_X1 U9743 ( .A(n13014), .ZN(n11761) );
  OR2_X1 U9744 ( .A1(n9845), .A2(n9844), .ZN(n9846) );
  OR2_X1 U9745 ( .A1(n9338), .A2(n9337), .ZN(n13193) );
  OR2_X1 U9746 ( .A1(n14895), .A2(P2_U3088), .ZN(n14930) );
  OR2_X1 U9747 ( .A1(n10111), .A2(P2_U3088), .ZN(n14946) );
  NAND2_X1 U9748 ( .A1(n13519), .A2(n9479), .ZN(n13467) );
  AND2_X2 U9749 ( .A1(n10546), .A2(n10545), .ZN(n15002) );
  INV_X1 U9750 ( .A(n13317), .ZN(n13647) );
  AND2_X2 U9751 ( .A1(n10546), .A2(n14953), .ZN(n14995) );
  INV_X1 U9752 ( .A(n14950), .ZN(n14951) );
  INV_X1 U9753 ( .A(n14954), .ZN(n14957) );
  INV_X1 U9754 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10181) );
  AND2_X1 U9755 ( .A1(n9976), .A2(n9923), .ZN(n14615) );
  AND2_X1 U9756 ( .A1(n10700), .A2(n12324), .ZN(n14606) );
  OR2_X1 U9757 ( .A1(n10074), .A2(n10073), .ZN(n14593) );
  OR2_X1 U9758 ( .A1(n10064), .A2(n9906), .ZN(n13849) );
  OR2_X1 U9759 ( .A1(n14618), .A2(n9996), .ZN(n14634) );
  OR2_X1 U9760 ( .A1(n14618), .A2(n9980), .ZN(n13899) );
  NAND2_X1 U9761 ( .A1(n14721), .A2(n14504), .ZN(n14107) );
  INV_X1 U9762 ( .A(n14721), .ZN(n14736) );
  OR2_X1 U9763 ( .A1(n14811), .A2(n8897), .ZN(n8898) );
  AND2_X2 U9764 ( .A1(n8896), .A2(n8895), .ZN(n14811) );
  OR2_X1 U9765 ( .A1(n14799), .A2(n8067), .ZN(n8922) );
  AND3_X1 U9766 ( .A1(n14549), .A2(n14548), .A3(n14547), .ZN(n14563) );
  INV_X1 U9767 ( .A(n14799), .ZN(n14798) );
  AND2_X2 U9768 ( .A1(n8907), .A2(n8151), .ZN(n14799) );
  INV_X1 U9769 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11249) );
  INV_X1 U9770 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10376) );
  NOR2_X1 U9771 ( .A1(n14352), .A2(n14351), .ZN(n14350) );
  NOR2_X1 U9772 ( .A1(P2_U3088), .A2(n10094), .ZN(P2_U3947) );
  NAND2_X1 U9773 ( .A1(n8153), .A2(n8152), .ZN(P1_U3524) );
  NAND2_X1 U9774 ( .A1(n7499), .A2(SI_1_), .ZN(n7502) );
  INV_X1 U9775 ( .A(n7624), .ZN(n7501) );
  INV_X1 U9776 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8198) );
  INV_X1 U9777 ( .A(SI_0_), .ZN(n7636) );
  NOR2_X1 U9778 ( .A1(n7500), .A2(n7636), .ZN(n7622) );
  NAND2_X1 U9779 ( .A1(n7501), .A2(n7622), .ZN(n7626) );
  MUX2_X1 U9780 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n7503), .Z(n7504) );
  NAND2_X1 U9781 ( .A1(n7504), .A2(SI_2_), .ZN(n7506) );
  OAI21_X1 U9782 ( .B1(n7504), .B2(SI_2_), .A(n7506), .ZN(n7649) );
  INV_X1 U9783 ( .A(n7649), .ZN(n7505) );
  INV_X1 U9784 ( .A(n7669), .ZN(n7507) );
  INV_X1 U9785 ( .A(n7509), .ZN(n7679) );
  MUX2_X1 U9786 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n6532), .Z(n7511) );
  OAI21_X1 U9787 ( .B1(n7511), .B2(SI_5_), .A(n7513), .ZN(n7512) );
  INV_X1 U9788 ( .A(n7512), .ZN(n7699) );
  MUX2_X1 U9789 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n6533), .Z(n7514) );
  NAND2_X1 U9790 ( .A1(n7514), .A2(SI_6_), .ZN(n7516) );
  OAI21_X1 U9791 ( .B1(n7514), .B2(SI_6_), .A(n7516), .ZN(n7515) );
  INV_X1 U9792 ( .A(n7515), .ZN(n7717) );
  MUX2_X1 U9793 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9874), .Z(n7517) );
  OAI21_X1 U9794 ( .B1(n7517), .B2(SI_7_), .A(n7519), .ZN(n7518) );
  INV_X1 U9795 ( .A(n7518), .ZN(n7732) );
  MUX2_X1 U9796 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9874), .Z(n7520) );
  OAI21_X1 U9797 ( .B1(n7520), .B2(SI_8_), .A(n7522), .ZN(n7521) );
  INV_X1 U9798 ( .A(n7521), .ZN(n7751) );
  MUX2_X1 U9799 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n6533), .Z(n7523) );
  OAI21_X1 U9800 ( .B1(n7523), .B2(SI_9_), .A(n7525), .ZN(n7524) );
  INV_X1 U9801 ( .A(n7524), .ZN(n7768) );
  NAND2_X1 U9802 ( .A1(n7769), .A2(n7768), .ZN(n7771) );
  MUX2_X1 U9803 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n6533), .Z(n7526) );
  OAI21_X1 U9804 ( .B1(n7526), .B2(SI_10_), .A(n7528), .ZN(n7527) );
  INV_X1 U9805 ( .A(n7527), .ZN(n7788) );
  MUX2_X1 U9806 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n9874), .Z(n7529) );
  INV_X1 U9807 ( .A(n7529), .ZN(n7530) );
  MUX2_X1 U9808 ( .A(n10376), .B(n10181), .S(n9874), .Z(n7531) );
  INV_X1 U9809 ( .A(SI_12_), .ZN(n9895) );
  NAND2_X1 U9810 ( .A1(n7531), .A2(n9895), .ZN(n7532) );
  MUX2_X1 U9811 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n6533), .Z(n7533) );
  INV_X1 U9812 ( .A(n7533), .ZN(n7534) );
  NAND2_X1 U9813 ( .A1(n7534), .A2(n9915), .ZN(n7535) );
  MUX2_X1 U9814 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n9874), .Z(n7864) );
  NAND2_X1 U9815 ( .A1(n7864), .A2(SI_14_), .ZN(n7536) );
  MUX2_X1 U9816 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n9874), .Z(n7538) );
  NOR2_X1 U9817 ( .A1(n7864), .A2(SI_14_), .ZN(n7540) );
  INV_X1 U9818 ( .A(n7538), .ZN(n7866) );
  INV_X1 U9819 ( .A(SI_15_), .ZN(n10029) );
  AOI22_X1 U9820 ( .A1(n7540), .A2(n7539), .B1(n7866), .B2(n10029), .ZN(n7541)
         );
  MUX2_X1 U9821 ( .A(n10603), .B(n10732), .S(n9874), .Z(n7542) );
  INV_X1 U9822 ( .A(SI_16_), .ZN(n10053) );
  NAND2_X1 U9823 ( .A1(n7542), .A2(n10053), .ZN(n7543) );
  MUX2_X1 U9824 ( .A(n10757), .B(n10761), .S(n9874), .Z(n7899) );
  MUX2_X1 U9825 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n9874), .Z(n7918) );
  MUX2_X1 U9826 ( .A(n11249), .B(n11247), .S(n6533), .Z(n7547) );
  INV_X1 U9827 ( .A(SI_19_), .ZN(n10422) );
  INV_X1 U9828 ( .A(n7547), .ZN(n7548) );
  NAND2_X1 U9829 ( .A1(n7548), .A2(SI_19_), .ZN(n7549) );
  NAND2_X1 U9830 ( .A1(n7550), .A2(n7549), .ZN(n7932) );
  INV_X1 U9831 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11546) );
  INV_X1 U9832 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11550) );
  MUX2_X1 U9833 ( .A(n11546), .B(n11550), .S(n9874), .Z(n7944) );
  INV_X1 U9834 ( .A(n7944), .ZN(n7551) );
  INV_X1 U9835 ( .A(SI_20_), .ZN(n10754) );
  MUX2_X1 U9836 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n6533), .Z(n7556) );
  XNOR2_X1 U9837 ( .A(n7556), .B(SI_21_), .ZN(n7955) );
  INV_X1 U9838 ( .A(n7955), .ZN(n7555) );
  NAND2_X1 U9839 ( .A1(n7556), .A2(SI_21_), .ZN(n7557) );
  INV_X1 U9840 ( .A(SI_22_), .ZN(n7560) );
  MUX2_X1 U9841 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n6533), .Z(n9091) );
  INV_X1 U9842 ( .A(n9091), .ZN(n7561) );
  MUX2_X1 U9843 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n6533), .Z(n7604) );
  INV_X1 U9844 ( .A(n7604), .ZN(n7558) );
  INV_X1 U9845 ( .A(SI_23_), .ZN(n11154) );
  AOI22_X1 U9846 ( .A1(n7560), .A2(n7561), .B1(n7558), .B2(n11154), .ZN(n7559)
         );
  OAI21_X1 U9847 ( .B1(n7561), .B2(n7560), .A(n11154), .ZN(n7563) );
  AND2_X1 U9848 ( .A1(SI_22_), .A2(SI_23_), .ZN(n7562) );
  AOI22_X1 U9849 ( .A1(n7563), .A2(n7604), .B1(n9091), .B2(n7562), .ZN(n7564)
         );
  MUX2_X1 U9850 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9874), .Z(n7978) );
  NAND2_X1 U9851 ( .A1(n7627), .A2(n7565), .ZN(n7655) );
  NOR2_X1 U9852 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n7573) );
  NOR2_X1 U9853 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n7572) );
  XNOR2_X1 U9854 ( .A(n7577), .B(n7583), .ZN(n8072) );
  NAND2_X1 U9856 ( .A1(n11859), .A2(n12260), .ZN(n7582) );
  INV_X1 U9857 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11861) );
  OR2_X1 U9858 ( .A1(n7673), .A2(n11861), .ZN(n7581) );
  INV_X1 U9859 ( .A(n14155), .ZN(n13990) );
  NAND2_X1 U9860 ( .A1(n7584), .A2(n7587), .ZN(n14212) );
  BUF_X2 U9861 ( .A(n7589), .Z(n7591) );
  NAND2_X1 U9862 ( .A1(n7662), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n7599) );
  INV_X1 U9863 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n7590) );
  OR2_X1 U9864 ( .A1(n6541), .A2(n7590), .ZN(n7598) );
  NAND2_X1 U9865 ( .A1(n7708), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7724) );
  NAND2_X1 U9866 ( .A1(n7741), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7759) );
  AND2_X1 U9867 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n7592) );
  INV_X1 U9868 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7841) );
  INV_X1 U9869 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7855) );
  INV_X1 U9870 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7872) );
  NAND2_X1 U9871 ( .A1(n7890), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7910) );
  INV_X1 U9872 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n11881) );
  INV_X1 U9873 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n7927) );
  OAI21_X1 U9874 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n7593), .A(n7987), .ZN(
        n13782) );
  OR2_X1 U9875 ( .A1(n6535), .A2(n13782), .ZN(n7597) );
  NAND2_X1 U9876 ( .A1(n14218), .A2(n7594), .ZN(n7643) );
  INV_X1 U9877 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n7595) );
  OR2_X1 U9878 ( .A1(n12241), .A2(n7595), .ZN(n7596) );
  NAND4_X1 U9879 ( .A1(n7599), .A2(n7598), .A3(n7597), .A4(n7596), .ZN(n13847)
         );
  INV_X1 U9880 ( .A(n9092), .ZN(n7600) );
  NAND2_X1 U9881 ( .A1(n7600), .A2(n9091), .ZN(n7603) );
  NAND2_X1 U9882 ( .A1(n7601), .A2(SI_22_), .ZN(n7602) );
  XNOR2_X1 U9883 ( .A(n7604), .B(SI_23_), .ZN(n7605) );
  NAND2_X1 U9884 ( .A1(n11855), .A2(n12260), .ZN(n7608) );
  INV_X1 U9885 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11854) );
  OR2_X1 U9886 ( .A1(n7673), .A2(n11854), .ZN(n7607) );
  NAND2_X2 U9887 ( .A1(n7608), .A2(n7607), .ZN(n14160) );
  INV_X1 U9888 ( .A(n14160), .ZN(n14012) );
  NAND2_X1 U9889 ( .A1(n8065), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n7615) );
  INV_X1 U9890 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n14011) );
  OR2_X1 U9891 ( .A1(n12242), .A2(n14011), .ZN(n7614) );
  OAI21_X1 U9892 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n7610), .A(n7609), .ZN(
        n14007) );
  OR2_X1 U9893 ( .A1(n6535), .A2(n14007), .ZN(n7613) );
  INV_X1 U9894 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n7611) );
  OR2_X1 U9895 ( .A1(n6541), .A2(n7611), .ZN(n7612) );
  NAND4_X1 U9896 ( .A1(n7615), .A2(n7614), .A3(n7613), .A4(n7612), .ZN(n13848)
         );
  NAND2_X1 U9897 ( .A1(n7662), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7619) );
  INV_X1 U9898 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9969) );
  OR2_X1 U9899 ( .A1(n6539), .A2(n9969), .ZN(n7618) );
  INV_X1 U9900 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7616) );
  NAND2_X1 U9901 ( .A1(n7620), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n7621) );
  OR2_X1 U9902 ( .A1(n7673), .A2(n6715), .ZN(n7631) );
  INV_X1 U9903 ( .A(n7622), .ZN(n7623) );
  NAND2_X1 U9904 ( .A1(n7624), .A2(n7623), .ZN(n7625) );
  NAND2_X1 U9905 ( .A1(n7626), .A2(n7625), .ZN(n9877) );
  OR2_X1 U9906 ( .A1(n12236), .A2(n9877), .ZN(n7630) );
  OR2_X1 U9907 ( .A1(n7676), .A2(n13868), .ZN(n7629) );
  INV_X2 U9908 ( .A(n6540), .ZN(n8889) );
  NAND2_X1 U9909 ( .A1(n8889), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n7635) );
  INV_X1 U9910 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10880) );
  INV_X1 U9911 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10879) );
  INV_X1 U9912 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n14608) );
  OR2_X1 U9913 ( .A1(n7643), .A2(n14608), .ZN(n7632) );
  INV_X1 U9914 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7638) );
  NOR2_X1 U9915 ( .A1(n9874), .A2(n7636), .ZN(n7637) );
  XNOR2_X1 U9916 ( .A(n7637), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n14228) );
  MUX2_X1 U9917 ( .A(n7638), .B(n14228), .S(n7676), .Z(n10154) );
  OR2_X2 U9918 ( .A1(n13860), .A2(n11902), .ZN(n12091) );
  NAND2_X1 U9919 ( .A1(n12084), .A2(n12091), .ZN(n12085) );
  NAND2_X1 U9920 ( .A1(n12094), .A2(n12085), .ZN(n10185) );
  NAND2_X1 U9921 ( .A1(n7662), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7647) );
  INV_X1 U9922 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10910) );
  INV_X1 U9923 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7641) );
  INV_X1 U9924 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9970) );
  OR2_X1 U9925 ( .A1(n7643), .A2(n9970), .ZN(n7644) );
  NAND2_X1 U9927 ( .A1(n7650), .A2(n7649), .ZN(n7652) );
  OR2_X1 U9928 ( .A1(n12236), .A2(n9875), .ZN(n7658) );
  NOR2_X1 U9929 ( .A1(n7628), .A2(n7719), .ZN(n7653) );
  MUX2_X1 U9930 ( .A(n7719), .B(n7653), .S(P1_IR_REG_2__SCAN_IN), .Z(n7654) );
  INV_X1 U9931 ( .A(n7654), .ZN(n7656) );
  NAND2_X1 U9932 ( .A1(n7656), .A2(n7655), .ZN(n10139) );
  OR2_X1 U9933 ( .A1(n7676), .A2(n10139), .ZN(n7657) );
  AND3_X2 U9934 ( .A1(n7659), .A2(n7658), .A3(n7657), .ZN(n12092) );
  NAND2_X1 U9936 ( .A1(n7660), .A2(n12092), .ZN(n12088) );
  NAND2_X1 U9937 ( .A1(n12090), .A2(n12089), .ZN(n7661) );
  NAND2_X1 U9938 ( .A1(n12088), .A2(n7661), .ZN(n12273) );
  NAND2_X1 U9939 ( .A1(n8889), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n7666) );
  OR2_X1 U9940 ( .A1(n6535), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7665) );
  INV_X1 U9941 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n14720) );
  OR2_X1 U9942 ( .A1(n12242), .A2(n14720), .ZN(n7664) );
  INV_X1 U9943 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9972) );
  OR2_X1 U9944 ( .A1(n7643), .A2(n9972), .ZN(n7663) );
  NAND4_X2 U9945 ( .A1(n7666), .A2(n7665), .A3(n7664), .A4(n7663), .ZN(n13859)
         );
  NAND2_X1 U9946 ( .A1(n7655), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7667) );
  MUX2_X1 U9947 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7667), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n7668) );
  NAND2_X1 U9948 ( .A1(n7668), .A2(n7684), .ZN(n13878) );
  NAND2_X1 U9949 ( .A1(n7670), .A2(n7669), .ZN(n7672) );
  NAND2_X1 U9950 ( .A1(n7672), .A2(n7671), .ZN(n9898) );
  OR2_X1 U9951 ( .A1(n9898), .A2(n12236), .ZN(n7675) );
  OR2_X1 U9952 ( .A1(n7673), .A2(n9897), .ZN(n7674) );
  NAND2_X1 U9953 ( .A1(n14715), .A2(n14714), .ZN(n7678) );
  INV_X1 U9954 ( .A(n14724), .ZN(n12105) );
  OR2_X1 U9955 ( .A1(n13859), .A2(n12105), .ZN(n7677) );
  OR2_X1 U9956 ( .A1(n7680), .A2(n7679), .ZN(n7681) );
  INV_X2 U9957 ( .A(n7673), .ZN(n7937) );
  NAND2_X1 U9959 ( .A1(n7684), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7683) );
  MUX2_X1 U9960 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7683), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n7686) );
  INV_X1 U9961 ( .A(n7905), .ZN(n7685) );
  AOI22_X1 U9962 ( .A1(n7937), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n7936), .B2(
        n14620), .ZN(n7687) );
  OAI21_X1 U9963 ( .B1(n9880), .B2(n12236), .A(n7687), .ZN(n12110) );
  NAND2_X1 U9964 ( .A1(n8065), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7696) );
  INV_X1 U9965 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9981) );
  OR2_X1 U9966 ( .A1(n12242), .A2(n9981), .ZN(n7695) );
  INV_X1 U9967 ( .A(n7708), .ZN(n7691) );
  INV_X1 U9968 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7689) );
  INV_X1 U9969 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n7688) );
  NAND2_X1 U9970 ( .A1(n7689), .A2(n7688), .ZN(n7690) );
  NAND2_X1 U9971 ( .A1(n7691), .A2(n7690), .ZN(n11072) );
  OR2_X1 U9972 ( .A1(n6535), .A2(n11072), .ZN(n7694) );
  INV_X1 U9973 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7692) );
  OR2_X1 U9974 ( .A1(n6540), .A2(n7692), .ZN(n7693) );
  NOR2_X1 U9975 ( .A1(n14749), .A2(n14598), .ZN(n7697) );
  NAND2_X1 U9976 ( .A1(n14749), .A2(n14598), .ZN(n7698) );
  OR2_X1 U9977 ( .A1(n7700), .A2(n7699), .ZN(n7701) );
  NAND2_X1 U9978 ( .A1(n7702), .A2(n7701), .ZN(n9888) );
  OR2_X1 U9979 ( .A1(n9888), .A2(n12236), .ZN(n7707) );
  NOR2_X1 U9980 ( .A1(n7905), .A2(n7719), .ZN(n7703) );
  MUX2_X1 U9981 ( .A(n7719), .B(n7703), .S(P1_IR_REG_5__SCAN_IN), .Z(n7705) );
  OR2_X1 U9982 ( .A1(n7705), .A2(n7737), .ZN(n10014) );
  INV_X1 U9983 ( .A(n10014), .ZN(n9989) );
  AOI22_X1 U9984 ( .A1(n7937), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n7936), .B2(
        n9989), .ZN(n7706) );
  NAND2_X1 U9985 ( .A1(n7707), .A2(n7706), .ZN(n14704) );
  INV_X1 U9986 ( .A(n14704), .ZN(n14754) );
  NAND2_X1 U9987 ( .A1(n8889), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n7712) );
  INV_X1 U9988 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9973) );
  OR2_X1 U9989 ( .A1(n7643), .A2(n9973), .ZN(n7711) );
  INV_X1 U9990 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9988) );
  OR2_X1 U9991 ( .A1(n12242), .A2(n9988), .ZN(n7710) );
  OAI21_X1 U9992 ( .B1(n7708), .B2(P1_REG3_REG_5__SCAN_IN), .A(n7724), .ZN(
        n14700) );
  OR2_X1 U9993 ( .A1(n6535), .A2(n14700), .ZN(n7709) );
  NAND4_X1 U9994 ( .A1(n7712), .A2(n7711), .A3(n7710), .A4(n7709), .ZN(n13858)
         );
  NAND2_X1 U9995 ( .A1(n14754), .A2(n13858), .ZN(n7713) );
  INV_X1 U9996 ( .A(n13858), .ZN(n11003) );
  NAND2_X1 U9997 ( .A1(n11003), .A2(n14704), .ZN(n7716) );
  NAND2_X1 U9998 ( .A1(n7713), .A2(n7716), .ZN(n14689) );
  NAND2_X1 U9999 ( .A1(n14693), .A2(n7716), .ZN(n11001) );
  OR2_X1 U10000 ( .A1(n9893), .A2(n12236), .ZN(n7722) );
  OR2_X1 U10001 ( .A1(n7737), .A2(n7719), .ZN(n7720) );
  XNOR2_X1 U10002 ( .A(n7720), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9990) );
  AOI22_X1 U10003 ( .A1(n7937), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7936), .B2(
        n9990), .ZN(n7721) );
  NAND2_X1 U10004 ( .A1(n7722), .A2(n7721), .ZN(n14762) );
  NAND2_X1 U10005 ( .A1(n8065), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7730) );
  INV_X1 U10006 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11007) );
  OR2_X1 U10007 ( .A1(n12242), .A2(n11007), .ZN(n7729) );
  AND2_X1 U10008 ( .A1(n7724), .A2(n7723), .ZN(n7725) );
  OR2_X1 U10009 ( .A1(n7725), .A2(n7741), .ZN(n11008) );
  OR2_X1 U10010 ( .A1(n6535), .A2(n11008), .ZN(n7728) );
  INV_X1 U10011 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7726) );
  OR2_X1 U10012 ( .A1(n6540), .A2(n7726), .ZN(n7727) );
  NAND4_X1 U10013 ( .A1(n7730), .A2(n7729), .A3(n7728), .A4(n7727), .ZN(n13857) );
  XNOR2_X1 U10014 ( .A(n14762), .B(n13857), .ZN(n12278) );
  NAND2_X1 U10015 ( .A1(n11001), .A2(n12278), .ZN(n11000) );
  INV_X1 U10016 ( .A(n13857), .ZN(n14695) );
  NAND2_X1 U10017 ( .A1(n14762), .A2(n14695), .ZN(n7731) );
  OR2_X1 U10018 ( .A1(n7733), .A2(n7732), .ZN(n7734) );
  NAND2_X1 U10019 ( .A1(n7735), .A2(n7734), .ZN(n9901) );
  OR2_X1 U10020 ( .A1(n9901), .A2(n12236), .ZN(n7740) );
  INV_X1 U10021 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n7736) );
  NAND2_X1 U10022 ( .A1(n7737), .A2(n7736), .ZN(n7754) );
  NAND2_X1 U10023 ( .A1(n7754), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7738) );
  XNOR2_X1 U10024 ( .A(n7738), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10036) );
  AOI22_X1 U10025 ( .A1(n7937), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7936), .B2(
        n10036), .ZN(n7739) );
  NAND2_X1 U10026 ( .A1(n7740), .A2(n7739), .ZN(n14681) );
  NAND2_X1 U10027 ( .A1(n8065), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7747) );
  INV_X1 U10028 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9991) );
  OR2_X1 U10029 ( .A1(n12242), .A2(n9991), .ZN(n7746) );
  OR2_X1 U10030 ( .A1(n7741), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7742) );
  NAND2_X1 U10031 ( .A1(n7759), .A2(n7742), .ZN(n14679) );
  OR2_X1 U10032 ( .A1(n6535), .A2(n14679), .ZN(n7745) );
  INV_X1 U10033 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7743) );
  OR2_X1 U10034 ( .A1(n6540), .A2(n7743), .ZN(n7744) );
  NAND4_X1 U10035 ( .A1(n7747), .A2(n7746), .A3(n7745), .A4(n7744), .ZN(n13856) );
  INV_X1 U10036 ( .A(n13856), .ZN(n11002) );
  OR2_X1 U10037 ( .A1(n14681), .A2(n11002), .ZN(n7748) );
  NAND2_X1 U10038 ( .A1(n14675), .A2(n7748), .ZN(n7750) );
  NAND2_X1 U10039 ( .A1(n14681), .A2(n11002), .ZN(n7749) );
  NAND2_X1 U10040 ( .A1(n7753), .A2(n7752), .ZN(n9914) );
  OR2_X1 U10041 ( .A1(n9914), .A2(n12236), .ZN(n7757) );
  NAND2_X1 U10042 ( .A1(n7772), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7755) );
  XNOR2_X1 U10043 ( .A(n7755), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10198) );
  AOI22_X1 U10044 ( .A1(n7937), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7936), .B2(
        n10198), .ZN(n7756) );
  NAND2_X1 U10045 ( .A1(n7662), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7765) );
  INV_X1 U10046 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10037) );
  OR2_X1 U10047 ( .A1(n7643), .A2(n10037), .ZN(n7764) );
  NAND2_X1 U10048 ( .A1(n7759), .A2(n7758), .ZN(n7760) );
  NAND2_X1 U10049 ( .A1(n7780), .A2(n7760), .ZN(n11205) );
  OR2_X1 U10050 ( .A1(n6535), .A2(n11205), .ZN(n7763) );
  INV_X1 U10051 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7761) );
  OR2_X1 U10052 ( .A1(n6541), .A2(n7761), .ZN(n7762) );
  NAND4_X1 U10053 ( .A1(n7765), .A2(n7764), .A3(n7763), .A4(n7762), .ZN(n13855) );
  XNOR2_X1 U10054 ( .A(n12127), .B(n13855), .ZN(n12281) );
  INV_X1 U10055 ( .A(n13855), .ZN(n7766) );
  OR2_X1 U10056 ( .A1(n12127), .A2(n7766), .ZN(n7767) );
  OR2_X1 U10057 ( .A1(n7769), .A2(n7768), .ZN(n7770) );
  NAND2_X1 U10058 ( .A1(n7771), .A2(n7770), .ZN(n9927) );
  OR2_X1 U10059 ( .A1(n9927), .A2(n12236), .ZN(n7778) );
  NAND2_X1 U10060 ( .A1(n7773), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7808) );
  INV_X1 U10061 ( .A(n7808), .ZN(n7774) );
  NAND2_X1 U10062 ( .A1(n7774), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n7776) );
  NAND2_X1 U10063 ( .A1(n7808), .A2(n7775), .ZN(n7792) );
  AOI22_X1 U10064 ( .A1(n7937), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7936), .B2(
        n10518), .ZN(n7777) );
  NAND2_X1 U10065 ( .A1(n8889), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7785) );
  INV_X1 U10066 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10196) );
  OR2_X1 U10067 ( .A1(n12241), .A2(n10196), .ZN(n7784) );
  INV_X1 U10068 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10202) );
  OR2_X1 U10069 ( .A1(n12242), .A2(n10202), .ZN(n7783) );
  AND2_X1 U10070 ( .A1(n7780), .A2(n7779), .ZN(n7781) );
  OR2_X1 U10071 ( .A1(n7781), .A2(n7812), .ZN(n11445) );
  OR2_X1 U10072 ( .A1(n6535), .A2(n11445), .ZN(n7782) );
  NAND4_X1 U10073 ( .A1(n7785), .A2(n7784), .A3(n7783), .A4(n7782), .ZN(n13854) );
  INV_X1 U10074 ( .A(n13854), .ZN(n7786) );
  XNOR2_X1 U10075 ( .A(n14665), .B(n7786), .ZN(n12283) );
  INV_X1 U10076 ( .A(n12283), .ZN(n14659) );
  NAND2_X1 U10077 ( .A1(n14656), .A2(n14659), .ZN(n14655) );
  NAND2_X1 U10078 ( .A1(n14665), .A2(n7786), .ZN(n7787) );
  OR2_X1 U10079 ( .A1(n7789), .A2(n7788), .ZN(n7790) );
  NAND2_X1 U10080 ( .A1(n7791), .A2(n7790), .ZN(n9967) );
  OR2_X1 U10081 ( .A1(n9967), .A2(n12236), .ZN(n7795) );
  NAND2_X1 U10082 ( .A1(n7792), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7793) );
  XNOR2_X1 U10083 ( .A(n7793), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10586) );
  AOI22_X1 U10084 ( .A1(n7937), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7936), 
        .B2(n10586), .ZN(n7794) );
  NAND2_X1 U10085 ( .A1(n8065), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7800) );
  INV_X1 U10086 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10590) );
  OR2_X1 U10087 ( .A1(n12242), .A2(n10590), .ZN(n7799) );
  INV_X1 U10088 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7796) );
  OR2_X1 U10089 ( .A1(n6541), .A2(n7796), .ZN(n7798) );
  XNOR2_X1 U10090 ( .A(n7812), .B(P1_REG3_REG_10__SCAN_IN), .ZN(n14492) );
  OR2_X1 U10091 ( .A1(n6535), .A2(n14492), .ZN(n7797) );
  NAND4_X1 U10092 ( .A1(n7800), .A2(n7799), .A3(n7798), .A4(n7797), .ZN(n13853) );
  INV_X1 U10093 ( .A(n13853), .ZN(n11681) );
  OR2_X1 U10094 ( .A1(n14478), .A2(n11681), .ZN(n7803) );
  NAND2_X1 U10095 ( .A1(n14478), .A2(n11681), .ZN(n7801) );
  NAND2_X1 U10096 ( .A1(n7803), .A2(n7801), .ZN(n12284) );
  INV_X1 U10097 ( .A(n12284), .ZN(n7802) );
  NAND2_X1 U10098 ( .A1(n10045), .A2(n12260), .ZN(n7811) );
  NAND2_X1 U10099 ( .A1(n7806), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7807) );
  NAND2_X1 U10100 ( .A1(n7808), .A2(n7807), .ZN(n7823) );
  INV_X1 U10101 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n7809) );
  XNOR2_X1 U10102 ( .A(n7823), .B(n7809), .ZN(n10833) );
  AOI22_X1 U10103 ( .A1(n7937), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7936), 
        .B2(n10833), .ZN(n7810) );
  NAND2_X1 U10104 ( .A1(n8889), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7817) );
  AOI21_X1 U10105 ( .B1(n7812), .B2(P1_REG3_REG_10__SCAN_IN), .A(
        P1_REG3_REG_11__SCAN_IN), .ZN(n7813) );
  OR2_X1 U10106 ( .A1(n7826), .A2(n7813), .ZN(n14519) );
  OR2_X1 U10107 ( .A1(n6535), .A2(n14519), .ZN(n7816) );
  INV_X1 U10108 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10837) );
  OR2_X1 U10109 ( .A1(n12242), .A2(n10837), .ZN(n7815) );
  INV_X1 U10110 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10587) );
  OR2_X1 U10111 ( .A1(n7643), .A2(n10587), .ZN(n7814) );
  NAND4_X1 U10112 ( .A1(n7817), .A2(n7816), .A3(n7815), .A4(n7814), .ZN(n13852) );
  OR2_X1 U10113 ( .A1(n14521), .A2(n11676), .ZN(n7820) );
  NAND2_X1 U10114 ( .A1(n14521), .A2(n11676), .ZN(n7818) );
  NAND2_X1 U10115 ( .A1(n7820), .A2(n7818), .ZN(n14523) );
  INV_X1 U10116 ( .A(n14523), .ZN(n7819) );
  XNOR2_X1 U10117 ( .A(n7822), .B(n7821), .ZN(n10180) );
  NAND2_X1 U10118 ( .A1(n10180), .A2(n12260), .ZN(n7825) );
  OAI21_X1 U10119 ( .B1(n7823), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7837) );
  XNOR2_X1 U10120 ( .A(n7837), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11236) );
  AOI22_X1 U10121 ( .A1(n11236), .A2(n7936), .B1(n7937), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n7824) );
  NAND2_X1 U10122 ( .A1(n8889), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7831) );
  INV_X1 U10123 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11632) );
  OR2_X1 U10124 ( .A1(n12242), .A2(n11632), .ZN(n7830) );
  OR2_X1 U10125 ( .A1(n7826), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7827) );
  NAND2_X1 U10126 ( .A1(n7842), .A2(n7827), .ZN(n11754) );
  OR2_X1 U10127 ( .A1(n6535), .A2(n11754), .ZN(n7829) );
  INV_X1 U10128 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10831) );
  OR2_X1 U10129 ( .A1(n12241), .A2(n10831), .ZN(n7828) );
  NAND4_X1 U10130 ( .A1(n7831), .A2(n7830), .A3(n7829), .A4(n7828), .ZN(n13851) );
  XNOR2_X1 U10131 ( .A(n12147), .B(n13851), .ZN(n12285) );
  INV_X1 U10132 ( .A(n13851), .ZN(n7832) );
  OR2_X1 U10133 ( .A1(n12147), .A2(n7832), .ZN(n7833) );
  XNOR2_X1 U10134 ( .A(n7835), .B(n7834), .ZN(n10399) );
  NAND2_X1 U10135 ( .A1(n10399), .A2(n12260), .ZN(n7840) );
  INV_X1 U10136 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n7836) );
  NAND2_X1 U10137 ( .A1(n7837), .A2(n7836), .ZN(n7838) );
  NAND2_X1 U10138 ( .A1(n7838), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7850) );
  XNOR2_X1 U10139 ( .A(n7850), .B(P1_IR_REG_13__SCAN_IN), .ZN(n11375) );
  AOI22_X1 U10140 ( .A1(n11375), .A2(n7936), .B1(n7937), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n7839) );
  NAND2_X1 U10141 ( .A1(n8065), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7848) );
  INV_X1 U10142 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11655) );
  OR2_X1 U10143 ( .A1(n12242), .A2(n11655), .ZN(n7847) );
  NAND2_X1 U10144 ( .A1(n7842), .A2(n7841), .ZN(n7843) );
  NAND2_X1 U10145 ( .A1(n7856), .A2(n7843), .ZN(n11775) );
  OR2_X1 U10146 ( .A1(n6535), .A2(n11775), .ZN(n7846) );
  INV_X1 U10147 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7844) );
  OR2_X1 U10148 ( .A1(n6541), .A2(n7844), .ZN(n7845) );
  NAND4_X1 U10149 ( .A1(n7848), .A2(n7847), .A3(n7846), .A4(n7845), .ZN(n14114) );
  XNOR2_X1 U10150 ( .A(n12151), .B(n14114), .ZN(n12286) );
  INV_X1 U10151 ( .A(n14114), .ZN(n12152) );
  INV_X1 U10152 ( .A(SI_14_), .ZN(n9929) );
  XNOR2_X1 U10153 ( .A(n7862), .B(n9929), .ZN(n7865) );
  XNOR2_X1 U10154 ( .A(n7865), .B(n7864), .ZN(n10730) );
  NAND2_X1 U10155 ( .A1(n10730), .A2(n12260), .ZN(n7854) );
  INV_X1 U10156 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n7849) );
  NAND2_X1 U10157 ( .A1(n7850), .A2(n7849), .ZN(n7851) );
  NAND2_X1 U10158 ( .A1(n7851), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7852) );
  XNOR2_X1 U10159 ( .A(n7852), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11781) );
  AOI22_X1 U10160 ( .A1(n11781), .A2(n7936), .B1(n7937), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n7853) );
  NAND2_X1 U10161 ( .A1(n8889), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7861) );
  INV_X1 U10162 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11373) );
  OR2_X1 U10163 ( .A1(n12241), .A2(n11373), .ZN(n7860) );
  INV_X1 U10164 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n14119) );
  OR2_X1 U10165 ( .A1(n12242), .A2(n14119), .ZN(n7859) );
  NAND2_X1 U10166 ( .A1(n7856), .A2(n7855), .ZN(n7857) );
  NAND2_X1 U10167 ( .A1(n7873), .A2(n7857), .ZN(n14118) );
  OR2_X1 U10168 ( .A1(n6535), .A2(n14118), .ZN(n7858) );
  NAND2_X1 U10169 ( .A1(n14545), .A2(n11772), .ZN(n12155) );
  NAND2_X1 U10170 ( .A1(n12156), .A2(n12155), .ZN(n12288) );
  NAND2_X1 U10171 ( .A1(n14112), .A2(n14122), .ZN(n14111) );
  NAND2_X1 U10172 ( .A1(n14111), .A2(n12156), .ZN(n11849) );
  INV_X1 U10173 ( .A(n7862), .ZN(n7863) );
  OAI22_X1 U10174 ( .A1(n7865), .A2(n7864), .B1(n7863), .B2(SI_14_), .ZN(n7868) );
  XNOR2_X1 U10175 ( .A(n7866), .B(SI_15_), .ZN(n7867) );
  XNOR2_X1 U10176 ( .A(n7868), .B(n7867), .ZN(n10758) );
  NAND2_X1 U10177 ( .A1(n10758), .A2(n12260), .ZN(n7871) );
  NAND2_X1 U10178 ( .A1(n7905), .A2(n6655), .ZN(n7884) );
  NAND2_X1 U10179 ( .A1(n7884), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7869) );
  XNOR2_X1 U10180 ( .A(n7869), .B(P1_IR_REG_15__SCAN_IN), .ZN(n14646) );
  AOI22_X1 U10181 ( .A1(n7937), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7936), 
        .B2(n14646), .ZN(n7870) );
  AND2_X1 U10182 ( .A1(n7873), .A2(n7872), .ZN(n7874) );
  NOR2_X1 U10183 ( .A1(n7890), .A2(n7874), .ZN(n13833) );
  NAND2_X1 U10184 ( .A1(n7620), .A2(n13833), .ZN(n7881) );
  INV_X1 U10185 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7875) );
  OR2_X1 U10186 ( .A1(n12241), .A2(n7875), .ZN(n7880) );
  INV_X1 U10187 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7876) );
  OR2_X1 U10188 ( .A1(n12242), .A2(n7876), .ZN(n7879) );
  INV_X1 U10189 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n7877) );
  OR2_X1 U10190 ( .A1(n6541), .A2(n7877), .ZN(n7878) );
  NAND2_X1 U10191 ( .A1(n11950), .A2(n14113), .ZN(n12160) );
  NAND2_X1 U10192 ( .A1(n12159), .A2(n12160), .ZN(n12290) );
  XNOR2_X1 U10193 ( .A(n7883), .B(n7882), .ZN(n10602) );
  NAND2_X1 U10194 ( .A1(n10602), .A2(n12260), .ZN(n7889) );
  OR2_X1 U10195 ( .A1(n7884), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n7886) );
  NAND2_X1 U10196 ( .A1(n7886), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7885) );
  MUX2_X1 U10197 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7885), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n7887) );
  OR2_X1 U10198 ( .A1(n7886), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n7902) );
  AND2_X1 U10199 ( .A1(n7887), .A2(n7902), .ZN(n11885) );
  AOI22_X1 U10200 ( .A1(n7937), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7936), 
        .B2(n11885), .ZN(n7888) );
  OR2_X1 U10201 ( .A1(n7890), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7891) );
  AND2_X1 U10202 ( .A1(n7910), .A2(n7891), .ZN(n14508) );
  NAND2_X1 U10203 ( .A1(n7620), .A2(n14508), .ZN(n7896) );
  INV_X1 U10204 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11795) );
  OR2_X1 U10205 ( .A1(n12242), .A2(n11795), .ZN(n7895) );
  INV_X1 U10206 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n7892) );
  OR2_X1 U10207 ( .A1(n6540), .A2(n7892), .ZN(n7894) );
  INV_X1 U10208 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n11784) );
  OR2_X1 U10209 ( .A1(n12241), .A2(n11784), .ZN(n7893) );
  NAND4_X1 U10210 ( .A1(n7896), .A2(n7895), .A3(n7894), .A4(n7893), .ZN(n13850) );
  INV_X1 U10211 ( .A(n13850), .ZN(n12163) );
  XNOR2_X1 U10212 ( .A(n14531), .B(n12163), .ZN(n14503) );
  INV_X1 U10213 ( .A(n14503), .ZN(n7897) );
  NAND2_X1 U10214 ( .A1(n14531), .A2(n12163), .ZN(n7898) );
  XNOR2_X1 U10215 ( .A(n7899), .B(SI_17_), .ZN(n7900) );
  XNOR2_X1 U10216 ( .A(n7901), .B(n7900), .ZN(n10756) );
  NAND2_X1 U10217 ( .A1(n10756), .A2(n12260), .ZN(n7909) );
  NAND2_X1 U10218 ( .A1(n7902), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7903) );
  MUX2_X1 U10219 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7903), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n7904) );
  INV_X1 U10220 ( .A(n7904), .ZN(n7907) );
  NOR2_X1 U10221 ( .A1(n7907), .A2(n7923), .ZN(n13890) );
  AOI22_X1 U10222 ( .A1(n7937), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7936), 
        .B2(n13890), .ZN(n7908) );
  NAND2_X1 U10223 ( .A1(n7910), .A2(n11881), .ZN(n7911) );
  NAND2_X1 U10224 ( .A1(n7928), .A2(n7911), .ZN(n14100) );
  INV_X1 U10225 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n10336) );
  OAI22_X1 U10226 ( .A1(n14100), .A2(n6535), .B1(n6540), .B2(n10336), .ZN(
        n7915) );
  INV_X1 U10227 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n7913) );
  NAND2_X1 U10228 ( .A1(n7662), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7912) );
  OAI21_X1 U10229 ( .B1(n7913), .B2(n12241), .A(n7912), .ZN(n7914) );
  NOR2_X1 U10230 ( .A1(n14104), .A2(n14497), .ZN(n7917) );
  NAND2_X1 U10231 ( .A1(n14104), .A2(n14497), .ZN(n7916) );
  XNOR2_X1 U10232 ( .A(n7919), .B(n7918), .ZN(n11067) );
  NAND2_X1 U10233 ( .A1(n11067), .A2(n12260), .ZN(n7926) );
  INV_X1 U10234 ( .A(n7923), .ZN(n7920) );
  NAND2_X1 U10235 ( .A1(n7920), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7921) );
  MUX2_X1 U10236 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7921), .S(
        P1_IR_REG_18__SCAN_IN), .Z(n7924) );
  NAND2_X1 U10237 ( .A1(n7924), .A2(n7934), .ZN(n13895) );
  INV_X1 U10238 ( .A(n13895), .ZN(n13903) );
  AOI22_X1 U10239 ( .A1(n7937), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7936), 
        .B2(n13903), .ZN(n7925) );
  AND2_X1 U10240 ( .A1(n7928), .A2(n7927), .ZN(n7929) );
  OR2_X1 U10241 ( .A1(n7929), .A2(n7940), .ZN(n14085) );
  AOI22_X1 U10242 ( .A1(n8065), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n7662), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n7931) );
  NAND2_X1 U10243 ( .A1(n8889), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n7930) );
  OAI211_X1 U10244 ( .C1(n14085), .C2(n6535), .A(n7931), .B(n7930), .ZN(n14066) );
  XNOR2_X1 U10245 ( .A(n14091), .B(n14066), .ZN(n14079) );
  XNOR2_X1 U10246 ( .A(n7933), .B(n7932), .ZN(n11246) );
  NAND2_X1 U10247 ( .A1(n11246), .A2(n12260), .ZN(n7939) );
  INV_X1 U10248 ( .A(n7935), .ZN(n8062) );
  AOI22_X1 U10249 ( .A1(n7937), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14511), 
        .B2(n7936), .ZN(n7938) );
  NOR2_X1 U10250 ( .A1(n7940), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n7941) );
  OR2_X1 U10251 ( .A1(n7948), .A2(n7941), .ZN(n14069) );
  AOI22_X1 U10252 ( .A1(n7662), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n8889), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n7943) );
  NAND2_X1 U10253 ( .A1(n8065), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n7942) );
  OAI211_X1 U10254 ( .C1(n14069), .C2(n6535), .A(n7943), .B(n7942), .ZN(n14081) );
  INV_X1 U10255 ( .A(n14081), .ZN(n13810) );
  OR2_X1 U10256 ( .A1(n14181), .A2(n13810), .ZN(n12193) );
  NAND2_X1 U10257 ( .A1(n14181), .A2(n13810), .ZN(n12194) );
  XNOR2_X1 U10258 ( .A(n7945), .B(n7944), .ZN(n11545) );
  NAND2_X1 U10259 ( .A1(n11545), .A2(n12260), .ZN(n7947) );
  OR2_X1 U10260 ( .A1(n7673), .A2(n11546), .ZN(n7946) );
  NOR2_X1 U10261 ( .A1(n7948), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n7949) );
  OR2_X1 U10262 ( .A1(n7959), .A2(n7949), .ZN(n13792) );
  INV_X1 U10263 ( .A(n13792), .ZN(n14053) );
  INV_X1 U10264 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n7952) );
  NAND2_X1 U10265 ( .A1(n7662), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n7951) );
  NAND2_X1 U10266 ( .A1(n8889), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n7950) );
  OAI211_X1 U10267 ( .C1(n12241), .C2(n7952), .A(n7951), .B(n7950), .ZN(n7953)
         );
  AOI21_X1 U10268 ( .B1(n14053), .B2(n7620), .A(n7953), .ZN(n14034) );
  INV_X1 U10269 ( .A(n14034), .ZN(n14067) );
  XNOR2_X1 U10270 ( .A(n14058), .B(n14067), .ZN(n14056) );
  NAND2_X1 U10271 ( .A1(n14177), .A2(n14067), .ZN(n7954) );
  XNOR2_X1 U10272 ( .A(n7956), .B(n7955), .ZN(n11594) );
  NAND2_X1 U10273 ( .A1(n11594), .A2(n12260), .ZN(n7958) );
  INV_X1 U10274 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11595) );
  OR2_X1 U10275 ( .A1(n7673), .A2(n11595), .ZN(n7957) );
  OR2_X1 U10276 ( .A1(n7959), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n7961) );
  AND2_X1 U10277 ( .A1(n7961), .A2(n7960), .ZN(n14043) );
  NAND2_X1 U10278 ( .A1(n14043), .A2(n7620), .ZN(n7967) );
  INV_X1 U10279 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n7964) );
  NAND2_X1 U10280 ( .A1(n8889), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n7963) );
  NAND2_X1 U10281 ( .A1(n8065), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n7962) );
  OAI211_X1 U10282 ( .C1(n12242), .C2(n7964), .A(n7963), .B(n7962), .ZN(n7965)
         );
  INV_X1 U10283 ( .A(n7965), .ZN(n7966) );
  NAND2_X1 U10284 ( .A1(n7967), .A2(n7966), .ZN(n14050) );
  INV_X1 U10285 ( .A(n14050), .ZN(n7968) );
  XNOR2_X1 U10286 ( .A(n14044), .B(n7968), .ZN(n12293) );
  NAND2_X1 U10287 ( .A1(n8065), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n7976) );
  INV_X1 U10288 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n7969) );
  OR2_X1 U10289 ( .A1(n12242), .A2(n7969), .ZN(n7975) );
  OAI21_X1 U10290 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n7971), .A(n7970), .ZN(
        n13801) );
  OR2_X1 U10291 ( .A1(n6535), .A2(n13801), .ZN(n7974) );
  INV_X1 U10292 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n7972) );
  OR2_X1 U10293 ( .A1(n6540), .A2(n7972), .ZN(n7973) );
  NAND4_X1 U10294 ( .A1(n7976), .A2(n7975), .A3(n7974), .A4(n7973), .ZN(n14032) );
  XNOR2_X1 U10295 ( .A(n14160), .B(n13848), .ZN(n14002) );
  NAND2_X1 U10296 ( .A1(n14003), .A2(n14002), .ZN(n14001) );
  XNOR2_X1 U10297 ( .A(n14155), .B(n13847), .ZN(n13994) );
  INV_X1 U10298 ( .A(n13994), .ZN(n13982) );
  INV_X1 U10299 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11910) );
  INV_X1 U10300 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13706) );
  MUX2_X1 U10301 ( .A(n11910), .B(n13706), .S(n6533), .Z(n7981) );
  INV_X1 U10302 ( .A(SI_25_), .ZN(n11592) );
  NAND2_X1 U10303 ( .A1(n7981), .A2(n11592), .ZN(n7997) );
  INV_X1 U10304 ( .A(n7981), .ZN(n7982) );
  NAND2_X1 U10305 ( .A1(n7982), .A2(SI_25_), .ZN(n7983) );
  NAND2_X1 U10306 ( .A1(n7997), .A2(n7983), .ZN(n7998) );
  NAND2_X1 U10307 ( .A1(n11909), .A2(n12260), .ZN(n7985) );
  OR2_X1 U10308 ( .A1(n7673), .A2(n11910), .ZN(n7984) );
  NAND2_X1 U10309 ( .A1(n8065), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n7993) );
  INV_X1 U10310 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n13971) );
  OR2_X1 U10311 ( .A1(n12242), .A2(n13971), .ZN(n7992) );
  INV_X1 U10312 ( .A(n7987), .ZN(n7986) );
  NAND2_X1 U10313 ( .A1(n7986), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8005) );
  INV_X1 U10314 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n13754) );
  NAND2_X1 U10315 ( .A1(n13754), .A2(n7987), .ZN(n7988) );
  NAND2_X1 U10316 ( .A1(n8005), .A2(n7988), .ZN(n13753) );
  OR2_X1 U10317 ( .A1(n6535), .A2(n13753), .ZN(n7991) );
  INV_X1 U10318 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n7989) );
  OR2_X1 U10319 ( .A1(n6540), .A2(n7989), .ZN(n7990) );
  NAND4_X1 U10320 ( .A1(n7993), .A2(n7992), .A3(n7991), .A4(n7990), .ZN(n13846) );
  INV_X1 U10321 ( .A(n13846), .ZN(n7994) );
  NAND2_X1 U10322 ( .A1(n14147), .A2(n7994), .ZN(n7996) );
  OR2_X1 U10323 ( .A1(n14147), .A2(n7994), .ZN(n7995) );
  NAND2_X1 U10324 ( .A1(n7996), .A2(n7995), .ZN(n12294) );
  INV_X1 U10325 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14222) );
  INV_X1 U10326 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13703) );
  MUX2_X1 U10327 ( .A(n14222), .B(n13703), .S(n9874), .Z(n8015) );
  XNOR2_X1 U10328 ( .A(n8015), .B(SI_26_), .ZN(n8000) );
  NAND2_X1 U10329 ( .A1(n13702), .A2(n12260), .ZN(n8002) );
  OR2_X1 U10330 ( .A1(n7673), .A2(n14222), .ZN(n8001) );
  NAND2_X1 U10331 ( .A1(n7662), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8011) );
  INV_X1 U10332 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n8003) );
  OR2_X1 U10333 ( .A1(n12241), .A2(n8003), .ZN(n8010) );
  INV_X1 U10334 ( .A(n8005), .ZN(n8004) );
  NAND2_X1 U10335 ( .A1(n8004), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8024) );
  INV_X1 U10336 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n13824) );
  NAND2_X1 U10337 ( .A1(n8005), .A2(n13824), .ZN(n8006) );
  NAND2_X1 U10338 ( .A1(n8024), .A2(n8006), .ZN(n13954) );
  OR2_X1 U10339 ( .A1(n6535), .A2(n13954), .ZN(n8009) );
  INV_X1 U10340 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n8007) );
  OR2_X1 U10341 ( .A1(n6540), .A2(n8007), .ZN(n8008) );
  NAND4_X1 U10342 ( .A1(n8011), .A2(n8010), .A3(n8009), .A4(n8008), .ZN(n13845) );
  INV_X1 U10343 ( .A(n13845), .ZN(n8012) );
  NAND2_X1 U10344 ( .A1(n13960), .A2(n8012), .ZN(n8014) );
  OR2_X1 U10345 ( .A1(n13960), .A2(n8012), .ZN(n8013) );
  INV_X1 U10346 ( .A(n13946), .ZN(n13950) );
  NAND2_X1 U10347 ( .A1(n13949), .A2(n13950), .ZN(n13948) );
  NAND2_X1 U10348 ( .A1(n13948), .A2(n8014), .ZN(n13931) );
  INV_X1 U10349 ( .A(SI_26_), .ZN(n11696) );
  INV_X1 U10350 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14220) );
  INV_X1 U10351 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13700) );
  MUX2_X1 U10352 ( .A(n14220), .B(n13700), .S(n9874), .Z(n8034) );
  XNOR2_X1 U10353 ( .A(n8034), .B(SI_27_), .ZN(n8019) );
  NAND2_X1 U10354 ( .A1(n13699), .A2(n12260), .ZN(n8021) );
  OR2_X1 U10355 ( .A1(n7673), .A2(n14220), .ZN(n8020) );
  NAND2_X1 U10356 ( .A1(n8065), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8030) );
  INV_X1 U10357 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n8022) );
  OR2_X1 U10358 ( .A1(n12242), .A2(n8022), .ZN(n8029) );
  INV_X1 U10359 ( .A(n8024), .ZN(n8023) );
  NAND2_X1 U10360 ( .A1(n8023), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8045) );
  INV_X1 U10361 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n12049) );
  NAND2_X1 U10362 ( .A1(n8024), .A2(n12049), .ZN(n8025) );
  NAND2_X1 U10363 ( .A1(n8045), .A2(n8025), .ZN(n12048) );
  OR2_X1 U10364 ( .A1(n6535), .A2(n12048), .ZN(n8028) );
  INV_X1 U10365 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n8026) );
  OR2_X1 U10366 ( .A1(n6541), .A2(n8026), .ZN(n8027) );
  NAND4_X1 U10367 ( .A1(n8030), .A2(n8029), .A3(n8028), .A4(n8027), .ZN(n13844) );
  INV_X1 U10368 ( .A(n13844), .ZN(n8031) );
  NAND2_X1 U10369 ( .A1(n14137), .A2(n8031), .ZN(n8033) );
  OR2_X1 U10370 ( .A1(n14137), .A2(n8031), .ZN(n8032) );
  NAND2_X1 U10371 ( .A1(n8033), .A2(n8032), .ZN(n12297) );
  NAND2_X1 U10372 ( .A1(n13931), .A2(n13941), .ZN(n13930) );
  NAND2_X1 U10373 ( .A1(n13930), .A2(n8033), .ZN(n8053) );
  INV_X1 U10374 ( .A(SI_27_), .ZN(n11762) );
  NAND2_X1 U10375 ( .A1(n8035), .A2(n11762), .ZN(n8036) );
  INV_X1 U10376 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12061) );
  INV_X1 U10377 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13698) );
  MUX2_X1 U10378 ( .A(n12061), .B(n13698), .S(n6533), .Z(n8038) );
  INV_X1 U10379 ( .A(SI_28_), .ZN(n12327) );
  NAND2_X1 U10380 ( .A1(n8038), .A2(n12327), .ZN(n8882) );
  INV_X1 U10381 ( .A(n8038), .ZN(n8039) );
  NAND2_X1 U10382 ( .A1(n8039), .A2(SI_28_), .ZN(n8040) );
  NAND2_X1 U10383 ( .A1(n13695), .A2(n12260), .ZN(n8042) );
  OR2_X1 U10384 ( .A1(n7673), .A2(n12061), .ZN(n8041) );
  NAND2_X1 U10385 ( .A1(n8065), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8051) );
  INV_X1 U10386 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n12052) );
  OR2_X1 U10387 ( .A1(n12242), .A2(n12052), .ZN(n8050) );
  INV_X1 U10388 ( .A(n8045), .ZN(n8043) );
  NAND2_X1 U10389 ( .A1(n8043), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8906) );
  INV_X1 U10390 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8044) );
  NAND2_X1 U10391 ( .A1(n8045), .A2(n8044), .ZN(n8046) );
  NAND2_X1 U10392 ( .A1(n8906), .A2(n8046), .ZN(n12342) );
  OR2_X1 U10393 ( .A1(n6535), .A2(n12342), .ZN(n8049) );
  INV_X1 U10394 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n8047) );
  OR2_X1 U10395 ( .A1(n6540), .A2(n8047), .ZN(n8048) );
  NAND4_X1 U10396 ( .A1(n8051), .A2(n8050), .A3(n8049), .A4(n8048), .ZN(n13843) );
  NAND2_X1 U10397 ( .A1(n12344), .A2(n12335), .ZN(n8878) );
  OR2_X1 U10398 ( .A1(n12344), .A2(n12335), .ZN(n8052) );
  NAND2_X1 U10399 ( .A1(n8053), .A2(n8113), .ZN(n8879) );
  NAND2_X1 U10400 ( .A1(n8879), .A2(n8054), .ZN(n8076) );
  INV_X1 U10401 ( .A(n8057), .ZN(n8056) );
  INV_X1 U10402 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8055) );
  NAND2_X1 U10403 ( .A1(n8056), .A2(n8055), .ZN(n8121) );
  NAND2_X1 U10404 ( .A1(n8060), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8061) );
  XNOR2_X1 U10405 ( .A(n8061), .B(P1_IR_REG_21__SCAN_IN), .ZN(n8114) );
  NAND2_X1 U10406 ( .A1(n8062), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8063) );
  XNOR2_X1 U10407 ( .A(n8063), .B(n10344), .ZN(n12255) );
  INV_X1 U10408 ( .A(n12255), .ZN(n10878) );
  NAND2_X1 U10409 ( .A1(n8114), .A2(n10878), .ZN(n8064) );
  NAND2_X1 U10410 ( .A1(n8065), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8071) );
  NAND2_X1 U10411 ( .A1(n7662), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8070) );
  OR2_X1 U10412 ( .A1(n6535), .A2(n8906), .ZN(n8069) );
  INV_X1 U10413 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8067) );
  OR2_X1 U10414 ( .A1(n6540), .A2(n8067), .ZN(n8068) );
  NAND4_X1 U10415 ( .A1(n8071), .A2(n8070), .A3(n8069), .A4(n8068), .ZN(n13842) );
  NAND2_X1 U10416 ( .A1(n13842), .A2(n14498), .ZN(n8074) );
  INV_X1 U10417 ( .A(n12062), .ZN(n9996) );
  NAND2_X1 U10418 ( .A1(n9920), .A2(n9996), .ZN(n14696) );
  INV_X2 U10419 ( .A(n14696), .ZN(n14596) );
  NAND2_X1 U10420 ( .A1(n13844), .A2(n14596), .ZN(n8073) );
  NAND2_X1 U10421 ( .A1(n10149), .A2(n10150), .ZN(n10153) );
  INV_X1 U10422 ( .A(n11902), .ZN(n10177) );
  OR2_X1 U10423 ( .A1(n13860), .A2(n10177), .ZN(n8077) );
  NAND2_X1 U10424 ( .A1(n10153), .A2(n8077), .ZN(n10184) );
  NAND2_X1 U10425 ( .A1(n10184), .A2(n10183), .ZN(n10182) );
  NAND2_X1 U10426 ( .A1(n10182), .A2(n12088), .ZN(n14713) );
  INV_X1 U10427 ( .A(n14714), .ZN(n14712) );
  OR2_X1 U10428 ( .A1(n13859), .A2(n14724), .ZN(n8078) );
  INV_X1 U10429 ( .A(n14598), .ZN(n14697) );
  NAND2_X1 U10430 ( .A1(n14688), .A2(n14689), .ZN(n8080) );
  NAND2_X1 U10431 ( .A1(n14754), .A2(n11003), .ZN(n8079) );
  NAND2_X1 U10432 ( .A1(n8080), .A2(n8079), .ZN(n10999) );
  INV_X1 U10433 ( .A(n12278), .ZN(n8081) );
  NAND2_X1 U10434 ( .A1(n10999), .A2(n8081), .ZN(n8083) );
  INV_X1 U10435 ( .A(n14762), .ZN(n11009) );
  NAND2_X1 U10436 ( .A1(n11009), .A2(n14695), .ZN(n8082) );
  NAND2_X1 U10437 ( .A1(n8083), .A2(n8082), .ZN(n14673) );
  XNOR2_X1 U10438 ( .A(n14681), .B(n13856), .ZN(n12279) );
  NAND2_X1 U10439 ( .A1(n14673), .A2(n14674), .ZN(n8085) );
  OR2_X1 U10440 ( .A1(n14681), .A2(n13856), .ZN(n8084) );
  NAND2_X1 U10441 ( .A1(n8085), .A2(n8084), .ZN(n11197) );
  NAND2_X1 U10442 ( .A1(n11197), .A2(n11201), .ZN(n8087) );
  OR2_X1 U10443 ( .A1(n12127), .A2(n13855), .ZN(n8086) );
  NAND2_X1 U10444 ( .A1(n8087), .A2(n8086), .ZN(n14658) );
  NAND2_X1 U10445 ( .A1(n14658), .A2(n12283), .ZN(n8089) );
  OR2_X1 U10446 ( .A1(n14665), .A2(n13854), .ZN(n8088) );
  OR2_X1 U10447 ( .A1(n14478), .A2(n13853), .ZN(n8090) );
  INV_X1 U10448 ( .A(n12285), .ZN(n11625) );
  NAND2_X1 U10449 ( .A1(n11623), .A2(n11625), .ZN(n8092) );
  OR2_X1 U10450 ( .A1(n12147), .A2(n13851), .ZN(n8091) );
  NAND2_X1 U10451 ( .A1(n8092), .A2(n8091), .ZN(n11647) );
  INV_X1 U10452 ( .A(n12286), .ZN(n11648) );
  OR2_X1 U10453 ( .A1(n12151), .A2(n14114), .ZN(n8093) );
  INV_X1 U10454 ( .A(n11772), .ZN(n11945) );
  NAND2_X1 U10455 ( .A1(n14545), .A2(n11945), .ZN(n8094) );
  NAND2_X1 U10456 ( .A1(n14121), .A2(n8094), .ZN(n11842) );
  INV_X1 U10457 ( .A(n14113), .ZN(n14499) );
  OR2_X1 U10458 ( .A1(n11950), .A2(n14499), .ZN(n8096) );
  INV_X1 U10459 ( .A(n14105), .ZN(n8097) );
  NAND2_X1 U10460 ( .A1(n14192), .A2(n14497), .ZN(n12271) );
  AND2_X1 U10461 ( .A1(n14091), .A2(n14066), .ZN(n12190) );
  OR2_X1 U10462 ( .A1(n14091), .A2(n14066), .ZN(n12189) );
  INV_X1 U10463 ( .A(n14057), .ZN(n8100) );
  OR2_X1 U10464 ( .A1(n14177), .A2(n14034), .ZN(n8101) );
  OR2_X1 U10465 ( .A1(n14044), .A2(n14050), .ZN(n8102) );
  NAND2_X1 U10466 ( .A1(n14040), .A2(n8102), .ZN(n14026) );
  OR2_X1 U10467 ( .A1(n14165), .A2(n14032), .ZN(n8103) );
  NAND2_X1 U10468 ( .A1(n14160), .A2(n13848), .ZN(n8104) );
  NAND2_X1 U10469 ( .A1(n14000), .A2(n8104), .ZN(n13993) );
  INV_X1 U10470 ( .A(n13993), .ZN(n8105) );
  OR2_X1 U10471 ( .A1(n14155), .A2(n13847), .ZN(n8106) );
  NAND2_X1 U10472 ( .A1(n14147), .A2(n13846), .ZN(n8107) );
  NAND2_X1 U10473 ( .A1(n13960), .A2(n13845), .ZN(n8108) );
  NAND2_X1 U10474 ( .A1(n13945), .A2(n8108), .ZN(n13940) );
  OR2_X1 U10475 ( .A1(n14137), .A2(n13844), .ZN(n8109) );
  NAND2_X1 U10476 ( .A1(n8111), .A2(n12086), .ZN(n8112) );
  NAND2_X1 U10477 ( .A1(n8112), .A2(n12332), .ZN(n8904) );
  OR2_X1 U10478 ( .A1(n8904), .A2(n14511), .ZN(n14660) );
  INV_X1 U10479 ( .A(n14787), .ZN(n14766) );
  NAND2_X1 U10480 ( .A1(n14660), .A2(n14766), .ZN(n14797) );
  NAND2_X1 U10481 ( .A1(n7088), .A2(n8113), .ZN(n12056) );
  NAND3_X1 U10482 ( .A1(n12057), .A2(n14797), .A3(n12056), .ZN(n8120) );
  NAND2_X1 U10483 ( .A1(n11902), .A2(n10154), .ZN(n10191) );
  NOR2_X1 U10485 ( .A1(n14725), .A2(n14724), .ZN(n14728) );
  NAND2_X1 U10486 ( .A1(n14728), .A2(n14749), .ZN(n14705) );
  NOR2_X2 U10488 ( .A1(n14706), .A2(n14762), .ZN(n14684) );
  INV_X1 U10489 ( .A(n14681), .ZN(n14769) );
  INV_X1 U10491 ( .A(n12127), .ZN(n14776) );
  NAND2_X1 U10492 ( .A1(n14682), .A2(n14776), .ZN(n14667) );
  OR2_X2 U10493 ( .A1(n14667), .A2(n14665), .ZN(n14668) );
  NOR2_X2 U10494 ( .A1(n14668), .A2(n14478), .ZN(n14525) );
  NAND2_X1 U10495 ( .A1(n14558), .A2(n14525), .ZN(n14524) );
  NOR2_X4 U10496 ( .A1(n14506), .A2(n14192), .ZN(n14099) );
  OR2_X2 U10497 ( .A1(n14021), .A2(n14160), .ZN(n14009) );
  OR2_X2 U10498 ( .A1(n14009), .A2(n14155), .ZN(n13986) );
  INV_X1 U10499 ( .A(n12263), .ZN(n8115) );
  AOI21_X1 U10500 ( .B1(n12344), .B2(n13935), .A(n14792), .ZN(n8116) );
  NAND2_X1 U10501 ( .A1(n8116), .A2(n8893), .ZN(n12053) );
  NAND2_X1 U10502 ( .A1(n14787), .A2(n12248), .ZN(n10061) );
  NAND2_X1 U10503 ( .A1(n12248), .A2(n10878), .ZN(n12314) );
  INV_X1 U10504 ( .A(n12314), .ZN(n8117) );
  NAND2_X1 U10505 ( .A1(n12344), .A2(n14761), .ZN(n8118) );
  AND2_X1 U10506 ( .A1(n12053), .A2(n8118), .ZN(n8119) );
  NAND2_X1 U10507 ( .A1(n12060), .A2(n7492), .ZN(n14135) );
  OAI21_X2 U10508 ( .B1(n8125), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8124) );
  INV_X1 U10509 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8123) );
  NAND2_X1 U10510 ( .A1(n8127), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8128) );
  XNOR2_X1 U10511 ( .A(n8128), .B(P1_IR_REG_26__SCAN_IN), .ZN(n9905) );
  NAND2_X1 U10512 ( .A1(n8121), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8132) );
  XNOR2_X1 U10513 ( .A(n8132), .B(n8131), .ZN(n9919) );
  NAND2_X1 U10514 ( .A1(n14716), .A2(n9920), .ZN(n10697) );
  NAND2_X1 U10515 ( .A1(n10072), .A2(n10697), .ZN(n12321) );
  INV_X1 U10516 ( .A(n12321), .ZN(n10062) );
  INV_X1 U10517 ( .A(n8133), .ZN(n11860) );
  NAND3_X1 U10518 ( .A1(n11860), .A2(n11911), .A3(P1_B_REG_SCAN_IN), .ZN(n8136) );
  INV_X1 U10519 ( .A(P1_B_REG_SCAN_IN), .ZN(n8134) );
  INV_X1 U10520 ( .A(n9905), .ZN(n14223) );
  AOI21_X1 U10521 ( .B1(n8133), .B2(n8134), .A(n14223), .ZN(n8135) );
  NAND2_X1 U10522 ( .A1(n8136), .A2(n8135), .ZN(n9904) );
  OR2_X1 U10523 ( .A1(n9904), .A2(P1_D_REG_0__SCAN_IN), .ZN(n8138) );
  OR2_X1 U10524 ( .A1(n8133), .A2(n9905), .ZN(n8137) );
  NAND2_X1 U10525 ( .A1(n8138), .A2(n8137), .ZN(n10057) );
  NOR4_X1 U10526 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n8147) );
  NOR4_X1 U10527 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n8146) );
  OR4_X1 U10528 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n8144) );
  NOR4_X1 U10529 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n8142) );
  NOR4_X1 U10530 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n8141) );
  NOR4_X1 U10531 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n8140) );
  NOR4_X1 U10532 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n8139) );
  NAND4_X1 U10533 ( .A1(n8142), .A2(n8141), .A3(n8140), .A4(n8139), .ZN(n8143)
         );
  NOR4_X1 U10534 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n8144), .A4(n8143), .ZN(n8145) );
  AND3_X1 U10535 ( .A1(n8147), .A2(n8146), .A3(n8145), .ZN(n8148) );
  OR2_X1 U10536 ( .A1(n9904), .A2(P1_D_REG_1__SCAN_IN), .ZN(n8150) );
  NAND2_X1 U10537 ( .A1(n11911), .A2(n14223), .ZN(n8149) );
  NAND2_X1 U10538 ( .A1(n8150), .A2(n8149), .ZN(n8908) );
  AND2_X1 U10539 ( .A1(n8908), .A2(n10061), .ZN(n8151) );
  NAND2_X1 U10540 ( .A1(n14135), .A2(n14799), .ZN(n8153) );
  NAND2_X1 U10541 ( .A1(n14798), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8152) );
  INV_X1 U10542 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8157) );
  NAND4_X1 U10543 ( .A1(n8155), .A2(n8154), .A3(n8341), .A4(n8302), .ZN(n8373)
         );
  INV_X1 U10544 ( .A(n8373), .ZN(n8156) );
  NOR2_X1 U10545 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), 
        .ZN(n8164) );
  NOR2_X1 U10546 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), 
        .ZN(n8163) );
  NOR2_X1 U10547 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), 
        .ZN(n8162) );
  NAND4_X1 U10548 ( .A1(n8864), .A2(n8860), .A3(n8165), .A4(n8871), .ZN(n8166)
         );
  INV_X1 U10549 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8169) );
  XNOR2_X2 U10550 ( .A(n8170), .B(P3_IR_REG_29__SCAN_IN), .ZN(n8171) );
  INV_X2 U10551 ( .A(n8679), .ZN(n8538) );
  NAND2_X1 U10552 ( .A1(n8538), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8178) );
  NAND2_X4 U10553 ( .A1(n8173), .A2(n8171), .ZN(n8651) );
  INV_X1 U10554 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15236) );
  OR2_X1 U10555 ( .A1(n8651), .A2(n15236), .ZN(n8177) );
  AND2_X2 U10556 ( .A1(n8172), .A2(n8171), .ZN(n8661) );
  INV_X1 U10557 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10447) );
  OR2_X1 U10558 ( .A1(n8284), .A2(n10447), .ZN(n8176) );
  INV_X1 U10559 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n8174) );
  OR2_X1 U10560 ( .A1(n6476), .A2(n8174), .ZN(n8175) );
  NAND2_X1 U10561 ( .A1(n8184), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8181) );
  INV_X1 U10562 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8180) );
  NAND2_X1 U10563 ( .A1(n8182), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8183) );
  NAND2_X4 U10564 ( .A1(n8185), .A2(n8184), .ZN(n12670) );
  AND2_X2 U10565 ( .A1(n10431), .A2(n9854), .ZN(n8358) );
  INV_X1 U10566 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9109) );
  NAND2_X1 U10567 ( .A1(n9109), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8186) );
  INV_X1 U10568 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9867) );
  NAND2_X1 U10569 ( .A1(n9876), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8187) );
  XNOR2_X1 U10570 ( .A(n8222), .B(n8221), .ZN(n9858) );
  NAND2_X1 U10571 ( .A1(n8358), .A2(n9858), .ZN(n8190) );
  INV_X4 U10572 ( .A(n10431), .ZN(n8518) );
  NAND2_X1 U10573 ( .A1(n8518), .A2(n6709), .ZN(n8189) );
  INV_X1 U10574 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n8191) );
  INV_X1 U10575 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10653) );
  OR2_X1 U10576 ( .A1(n8651), .A2(n10653), .ZN(n8196) );
  INV_X1 U10577 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n8192) );
  OR2_X1 U10578 ( .A1(n8284), .A2(n8192), .ZN(n8195) );
  INV_X1 U10579 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n8193) );
  OR2_X1 U10580 ( .A1(n6476), .A2(n8193), .ZN(n8194) );
  INV_X1 U10581 ( .A(n8208), .ZN(n8200) );
  NAND2_X1 U10582 ( .A1(n8198), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8199) );
  AND2_X1 U10583 ( .A1(n8200), .A2(n8199), .ZN(n8201) );
  NAND2_X1 U10584 ( .A1(n6533), .A2(SI_0_), .ZN(n9121) );
  OAI21_X1 U10585 ( .B1(n9874), .B2(n8201), .A(n9121), .ZN(n13024) );
  MUX2_X1 U10586 ( .A(n10764), .B(n13024), .S(n10431), .Z(n10511) );
  INV_X1 U10587 ( .A(n10511), .ZN(n10649) );
  NOR2_X2 U10588 ( .A1(n15257), .A2(n10649), .ZN(n15255) );
  NAND2_X1 U10589 ( .A1(n8661), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8207) );
  INV_X1 U10590 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n15269) );
  OR2_X1 U10591 ( .A1(n8651), .A2(n15269), .ZN(n8206) );
  INV_X1 U10592 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n8202) );
  OR2_X1 U10593 ( .A1(n6475), .A2(n8202), .ZN(n8205) );
  INV_X1 U10594 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n8203) );
  OR2_X1 U10595 ( .A1(n6476), .A2(n8203), .ZN(n8204) );
  NAND4_X1 U10596 ( .A1(n8207), .A2(n8206), .A3(n8205), .A4(n8204), .ZN(n12564) );
  NAND2_X1 U10597 ( .A1(n8274), .A2(SI_1_), .ZN(n8213) );
  XNOR2_X1 U10598 ( .A(n8209), .B(n8208), .ZN(n9865) );
  NAND2_X1 U10599 ( .A1(n8358), .A2(n9865), .ZN(n8212) );
  NAND2_X1 U10600 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n10764), .ZN(n8210) );
  NAND2_X1 U10601 ( .A1(n8518), .A2(n6465), .ZN(n8211) );
  NAND2_X1 U10602 ( .A1(n12564), .A2(n15254), .ZN(n8723) );
  NAND2_X1 U10603 ( .A1(n15255), .A2(n8723), .ZN(n15232) );
  NAND2_X1 U10604 ( .A1(n15232), .A2(n15230), .ZN(n8214) );
  NAND2_X1 U10605 ( .A1(n15234), .A2(n8739), .ZN(n15216) );
  NAND2_X1 U10606 ( .A1(n8661), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8220) );
  OR2_X1 U10607 ( .A1(n8651), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8219) );
  INV_X1 U10608 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n8215) );
  OR2_X1 U10609 ( .A1(n8679), .A2(n8215), .ZN(n8218) );
  INV_X1 U10610 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n8216) );
  OR2_X1 U10611 ( .A1(n6477), .A2(n8216), .ZN(n8217) );
  NAND4_X1 U10612 ( .A1(n8220), .A2(n8219), .A3(n8218), .A4(n8217), .ZN(n11016) );
  NAND2_X1 U10613 ( .A1(n9897), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8224) );
  NAND2_X1 U10614 ( .A1(n8241), .A2(n8224), .ZN(n8238) );
  XNOR2_X1 U10615 ( .A(n8240), .B(n8238), .ZN(n9860) );
  NAND2_X1 U10616 ( .A1(n8358), .A2(n9860), .ZN(n8229) );
  NAND2_X1 U10617 ( .A1(n10435), .A2(n8225), .ZN(n8243) );
  NAND2_X1 U10618 ( .A1(n8243), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8227) );
  INV_X1 U10619 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8226) );
  NAND2_X1 U10620 ( .A1(n8518), .A2(n10490), .ZN(n8228) );
  OAI211_X1 U10621 ( .C1(n8345), .C2(SI_3_), .A(n8229), .B(n8228), .ZN(n15224)
         );
  NAND2_X1 U10622 ( .A1(n11016), .A2(n15224), .ZN(n8743) );
  INV_X1 U10623 ( .A(n15219), .ZN(n8230) );
  NAND2_X1 U10624 ( .A1(n15216), .A2(n8230), .ZN(n8231) );
  NAND2_X1 U10625 ( .A1(n8636), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8237) );
  INV_X1 U10626 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n12590) );
  OR2_X1 U10627 ( .A1(n8284), .A2(n12590), .ZN(n8236) );
  AND2_X1 U10628 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8232) );
  NOR2_X1 U10629 ( .A1(n8250), .A2(n8232), .ZN(n11015) );
  OR2_X1 U10630 ( .A1(n8651), .A2(n11015), .ZN(n8235) );
  INV_X1 U10631 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n8233) );
  OR2_X1 U10632 ( .A1(n8679), .A2(n8233), .ZN(n8234) );
  INV_X1 U10633 ( .A(n8238), .ZN(n8239) );
  NAND2_X1 U10634 ( .A1(n9879), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8242) );
  NAND2_X1 U10635 ( .A1(n8259), .A2(n8242), .ZN(n8257) );
  XNOR2_X1 U10636 ( .A(n8258), .B(n8257), .ZN(n9862) );
  NAND2_X1 U10637 ( .A1(n8358), .A2(n9862), .ZN(n8247) );
  NAND2_X1 U10638 ( .A1(n8261), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8245) );
  INV_X1 U10639 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8244) );
  NAND2_X1 U10640 ( .A1(n8518), .A2(n12626), .ZN(n8246) );
  OAI211_X1 U10641 ( .C1(n8345), .C2(SI_4_), .A(n8247), .B(n8246), .ZN(n8928)
         );
  OR2_X1 U10642 ( .A1(n15217), .A2(n8928), .ZN(n8731) );
  NAND2_X1 U10643 ( .A1(n15217), .A2(n8928), .ZN(n8730) );
  INV_X1 U10644 ( .A(n11018), .ZN(n8248) );
  NAND2_X1 U10645 ( .A1(n8249), .A2(n8731), .ZN(n15203) );
  NAND2_X1 U10646 ( .A1(n8636), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8256) );
  INV_X1 U10647 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n12597) );
  OR2_X1 U10648 ( .A1(n8284), .A2(n12597), .ZN(n8255) );
  NAND2_X1 U10649 ( .A1(n8250), .A2(n10975), .ZN(n8267) );
  OR2_X1 U10650 ( .A1(n8250), .A2(n10975), .ZN(n8251) );
  AND2_X1 U10651 ( .A1(n8267), .A2(n8251), .ZN(n15211) );
  OR2_X1 U10652 ( .A1(n8651), .A2(n15211), .ZN(n8254) );
  INV_X1 U10653 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n8252) );
  OR2_X1 U10654 ( .A1(n8679), .A2(n8252), .ZN(n8253) );
  NAND4_X1 U10655 ( .A1(n8256), .A2(n8255), .A3(n8254), .A4(n8253), .ZN(n15189) );
  NAND2_X1 U10656 ( .A1(n9881), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8260) );
  NAND2_X1 U10657 ( .A1(n8278), .A2(n8260), .ZN(n8275) );
  XNOR2_X1 U10658 ( .A(n8277), .B(n8275), .ZN(n9856) );
  NAND2_X1 U10659 ( .A1(n8358), .A2(n9856), .ZN(n8265) );
  OAI21_X1 U10660 ( .B1(n8261), .B2(P3_IR_REG_4__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8262) );
  MUX2_X1 U10661 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8262), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n8263) );
  NAND2_X1 U10662 ( .A1(n8263), .A2(n8374), .ZN(n15014) );
  NAND2_X1 U10663 ( .A1(n8518), .A2(n15014), .ZN(n8264) );
  OAI211_X1 U10664 ( .C1(n8345), .C2(SI_5_), .A(n8265), .B(n8264), .ZN(n15210)
         );
  OR2_X1 U10665 ( .A1(n15189), .A2(n15210), .ZN(n8734) );
  NAND2_X1 U10666 ( .A1(n15189), .A2(n15210), .ZN(n8750) );
  NAND2_X1 U10667 ( .A1(n8734), .A2(n8750), .ZN(n15205) );
  NAND2_X1 U10668 ( .A1(n15203), .A2(n15202), .ZN(n8266) );
  NAND2_X1 U10669 ( .A1(n8266), .A2(n8734), .ZN(n15188) );
  NAND2_X1 U10670 ( .A1(n8636), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8273) );
  INV_X1 U10671 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n12625) );
  OR2_X1 U10672 ( .A1(n8284), .A2(n12625), .ZN(n8272) );
  NAND2_X1 U10673 ( .A1(n8267), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8268) );
  AND2_X1 U10674 ( .A1(n8285), .A2(n8268), .ZN(n15197) );
  OR2_X1 U10675 ( .A1(n8651), .A2(n15197), .ZN(n8271) );
  INV_X1 U10676 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n8269) );
  OR2_X1 U10677 ( .A1(n8679), .A2(n8269), .ZN(n8270) );
  NAND4_X1 U10678 ( .A1(n8273), .A2(n8272), .A3(n8271), .A4(n8270), .ZN(n12562) );
  NAND2_X1 U10679 ( .A1(n8674), .A2(SI_6_), .ZN(n8283) );
  INV_X1 U10680 ( .A(n8275), .ZN(n8276) );
  XNOR2_X1 U10681 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n8279) );
  XNOR2_X1 U10682 ( .A(n8292), .B(n8279), .ZN(n9884) );
  NAND2_X1 U10683 ( .A1(n8358), .A2(n9884), .ZN(n8282) );
  NAND2_X1 U10684 ( .A1(n8374), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8280) );
  XNOR2_X1 U10685 ( .A(n8280), .B(P3_IR_REG_6__SCAN_IN), .ZN(n12632) );
  NAND2_X1 U10686 ( .A1(n8518), .A2(n12632), .ZN(n8281) );
  NAND2_X1 U10687 ( .A1(n12562), .A2(n15196), .ZN(n8752) );
  NAND2_X1 U10688 ( .A1(n8755), .A2(n8752), .ZN(n15192) );
  NAND2_X1 U10689 ( .A1(n15186), .A2(n8755), .ZN(n11384) );
  NAND2_X1 U10690 ( .A1(n8538), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8290) );
  INV_X1 U10691 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n12623) );
  OR2_X1 U10692 ( .A1(n8284), .A2(n12623), .ZN(n8289) );
  AND2_X1 U10693 ( .A1(n8285), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8286) );
  NOR2_X1 U10694 ( .A1(n8309), .A2(n8286), .ZN(n11392) );
  OR2_X1 U10695 ( .A1(n8651), .A2(n11392), .ZN(n8288) );
  INV_X1 U10696 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n12624) );
  OR2_X1 U10697 ( .A1(n6477), .A2(n12624), .ZN(n8287) );
  NAND4_X1 U10698 ( .A1(n8290), .A2(n8289), .A3(n8288), .A4(n8287), .ZN(n15190) );
  NAND2_X1 U10699 ( .A1(n9891), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8291) );
  NAND2_X1 U10700 ( .A1(n9892), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8293) );
  NAND2_X1 U10701 ( .A1(n9900), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8295) );
  NAND2_X1 U10702 ( .A1(n8316), .A2(n8295), .ZN(n8296) );
  NAND2_X1 U10703 ( .A1(n8297), .A2(n8296), .ZN(n8298) );
  NAND2_X1 U10704 ( .A1(n8317), .A2(n8298), .ZN(n9864) );
  INV_X1 U10705 ( .A(n9864), .ZN(n8299) );
  OR2_X1 U10706 ( .A1(n8374), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n8301) );
  NAND2_X1 U10707 ( .A1(n8301), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8300) );
  MUX2_X1 U10708 ( .A(n8300), .B(P3_IR_REG_31__SCAN_IN), .S(n8302), .Z(n8304)
         );
  INV_X1 U10709 ( .A(n8301), .ZN(n8303) );
  NAND2_X1 U10710 ( .A1(n8303), .A2(n8302), .ZN(n8340) );
  NAND2_X1 U10711 ( .A1(n8304), .A2(n8340), .ZN(n15052) );
  NAND2_X1 U10712 ( .A1(n8518), .A2(n15052), .ZN(n8305) );
  OAI211_X1 U10713 ( .C1(n8345), .C2(SI_7_), .A(n8306), .B(n8305), .ZN(n11391)
         );
  NAND2_X1 U10714 ( .A1(n15190), .A2(n11391), .ZN(n8757) );
  INV_X1 U10715 ( .A(n11386), .ZN(n8754) );
  NAND2_X1 U10716 ( .A1(n11384), .A2(n8754), .ZN(n8307) );
  NAND2_X1 U10717 ( .A1(n8307), .A2(n8756), .ZN(n11398) );
  NAND2_X1 U10718 ( .A1(n8636), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8315) );
  INV_X1 U10719 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n12621) );
  OR2_X1 U10720 ( .A1(n8284), .A2(n12621), .ZN(n8314) );
  NOR2_X1 U10721 ( .A1(n8309), .A2(n8308), .ZN(n8310) );
  OR2_X1 U10722 ( .A1(n8328), .A2(n8310), .ZN(n11403) );
  INV_X1 U10723 ( .A(n11403), .ZN(n11472) );
  OR2_X1 U10724 ( .A1(n8651), .A2(n11472), .ZN(n8313) );
  INV_X1 U10725 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n8311) );
  OR2_X1 U10726 ( .A1(n8679), .A2(n8311), .ZN(n8312) );
  NAND2_X1 U10727 ( .A1(n8674), .A2(SI_8_), .ZN(n8326) );
  NAND2_X1 U10728 ( .A1(n8318), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8319) );
  OR2_X1 U10729 ( .A1(n8321), .A2(n8320), .ZN(n8322) );
  AND2_X1 U10730 ( .A1(n8335), .A2(n8322), .ZN(n9869) );
  NAND2_X1 U10731 ( .A1(n8358), .A2(n9869), .ZN(n8325) );
  NAND2_X1 U10732 ( .A1(n8340), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8323) );
  XNOR2_X1 U10733 ( .A(n8323), .B(P3_IR_REG_8__SCAN_IN), .ZN(n12640) );
  NAND2_X1 U10734 ( .A1(n8518), .A2(n12640), .ZN(n8324) );
  XNOR2_X1 U10735 ( .A(n12561), .B(n7322), .ZN(n11397) );
  NAND2_X1 U10736 ( .A1(n11398), .A2(n11397), .ZN(n8327) );
  NAND2_X1 U10737 ( .A1(n11452), .A2(n7322), .ZN(n8762) );
  NAND2_X1 U10738 ( .A1(n8538), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8333) );
  INV_X1 U10739 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n12620) );
  OR2_X1 U10740 ( .A1(n6477), .A2(n12620), .ZN(n8332) );
  INV_X1 U10741 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n12619) );
  OR2_X1 U10742 ( .A1(n8284), .A2(n12619), .ZN(n8331) );
  OR2_X1 U10743 ( .A1(n8328), .A2(n11328), .ZN(n8329) );
  AND2_X1 U10744 ( .A1(n8346), .A2(n8329), .ZN(n11460) );
  OR2_X1 U10745 ( .A1(n8651), .A2(n11460), .ZN(n8330) );
  NAND2_X1 U10746 ( .A1(n9924), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8352) );
  NAND2_X1 U10747 ( .A1(n9926), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8336) );
  OR2_X1 U10748 ( .A1(n8338), .A2(n8337), .ZN(n8339) );
  NAND2_X1 U10749 ( .A1(n8353), .A2(n8339), .ZN(n9873) );
  NAND2_X1 U10750 ( .A1(n8358), .A2(n9873), .ZN(n8344) );
  NAND2_X1 U10751 ( .A1(n8359), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8342) );
  XNOR2_X1 U10752 ( .A(n8342), .B(n8341), .ZN(n15083) );
  NAND2_X1 U10753 ( .A1(n8518), .A2(n15083), .ZN(n8343) );
  OAI211_X1 U10754 ( .C1(n8345), .C2(SI_9_), .A(n8344), .B(n8343), .ZN(n11459)
         );
  NOR2_X1 U10755 ( .A1(n12560), .A2(n11459), .ZN(n8765) );
  NAND2_X1 U10756 ( .A1(n12560), .A2(n11459), .ZN(n8767) );
  OAI21_X2 U10757 ( .B1(n11450), .B2(n8765), .A(n8767), .ZN(n11514) );
  NAND2_X1 U10758 ( .A1(n8538), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8351) );
  INV_X1 U10759 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11528) );
  OR2_X1 U10760 ( .A1(n6477), .A2(n11528), .ZN(n8350) );
  INV_X1 U10761 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n12589) );
  OR2_X1 U10762 ( .A1(n8284), .A2(n12589), .ZN(n8349) );
  NAND2_X1 U10763 ( .A1(n8346), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8347) );
  AND2_X1 U10764 ( .A1(n8367), .A2(n8347), .ZN(n11525) );
  NAND2_X1 U10765 ( .A1(n9965), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8377) );
  NAND2_X1 U10766 ( .A1(n9966), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8354) );
  OR2_X1 U10767 ( .A1(n8356), .A2(n8355), .ZN(n8357) );
  NAND2_X1 U10768 ( .A1(n8378), .A2(n8357), .ZN(n9883) );
  NAND2_X1 U10769 ( .A1(n8358), .A2(n9883), .ZN(n8363) );
  OAI21_X1 U10770 ( .B1(n8359), .B2(P3_IR_REG_9__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8361) );
  INV_X1 U10771 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8360) );
  XNOR2_X1 U10772 ( .A(n8361), .B(n8360), .ZN(n15100) );
  NAND2_X1 U10773 ( .A1(n8518), .A2(n15100), .ZN(n8362) );
  OAI211_X1 U10774 ( .C1(n8345), .C2(SI_10_), .A(n8363), .B(n8362), .ZN(n11524) );
  AND2_X1 U10775 ( .A1(n12559), .A2(n11524), .ZN(n8364) );
  INV_X1 U10776 ( .A(n11524), .ZN(n11408) );
  NAND2_X1 U10777 ( .A1(n14453), .A2(n11408), .ZN(n8365) );
  NAND2_X1 U10778 ( .A1(n8538), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8372) );
  INV_X1 U10779 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n8366) );
  OR2_X1 U10780 ( .A1(n6477), .A2(n8366), .ZN(n8371) );
  OR2_X1 U10781 ( .A1(n8284), .A2(n14471), .ZN(n8370) );
  NAND2_X1 U10782 ( .A1(n8367), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8368) );
  AND2_X1 U10783 ( .A1(n8395), .A2(n8368), .ZN(n14456) );
  OR2_X1 U10784 ( .A1(n8651), .A2(n14456), .ZN(n8369) );
  NAND4_X1 U10785 ( .A1(n8372), .A2(n8371), .A3(n8370), .A4(n8369), .ZN(n12558) );
  OR2_X1 U10786 ( .A1(n8374), .A2(n8373), .ZN(n8375) );
  NAND2_X1 U10787 ( .A1(n8375), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8376) );
  XNOR2_X1 U10788 ( .A(n8376), .B(n8157), .ZN(n15117) );
  AOI22_X1 U10789 ( .A1(n8674), .A2(n9889), .B1(n8518), .B2(n15117), .ZN(n8384) );
  NAND2_X1 U10790 ( .A1(n10056), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8385) );
  NAND2_X1 U10791 ( .A1(n10046), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8379) );
  OR2_X1 U10792 ( .A1(n8381), .A2(n8380), .ZN(n8382) );
  NAND2_X1 U10793 ( .A1(n8386), .A2(n8382), .ZN(n9890) );
  NAND2_X1 U10794 ( .A1(n9890), .A2(n8673), .ZN(n8383) );
  NAND2_X1 U10795 ( .A1(n12558), .A2(n14455), .ZN(n8774) );
  NAND2_X1 U10796 ( .A1(n8773), .A2(n8774), .ZN(n14451) );
  INV_X1 U10797 ( .A(n14451), .ZN(n14448) );
  NAND2_X1 U10798 ( .A1(n10376), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8401) );
  NAND2_X1 U10799 ( .A1(n10181), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8387) );
  OR2_X1 U10800 ( .A1(n8389), .A2(n8388), .ZN(n8390) );
  NAND2_X1 U10801 ( .A1(n8402), .A2(n8390), .ZN(n9896) );
  OR2_X1 U10802 ( .A1(n9896), .A2(n8532), .ZN(n8394) );
  OR2_X1 U10803 ( .A1(n8391), .A2(n13011), .ZN(n8392) );
  INV_X1 U10804 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8408) );
  XNOR2_X1 U10805 ( .A(n8392), .B(n8408), .ZN(n15135) );
  INV_X1 U10806 ( .A(n15135), .ZN(n12653) );
  AOI22_X1 U10807 ( .A1(n8674), .A2(SI_12_), .B1(n8518), .B2(n12653), .ZN(
        n8393) );
  NAND2_X1 U10808 ( .A1(n8538), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8399) );
  INV_X1 U10809 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n12588) );
  OR2_X1 U10810 ( .A1(n8284), .A2(n12588), .ZN(n8398) );
  NOR2_X1 U10811 ( .A1(n8416), .A2(n7477), .ZN(n11728) );
  OR2_X1 U10812 ( .A1(n8651), .A2(n11728), .ZN(n8397) );
  INV_X1 U10813 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11618) );
  NAND4_X1 U10814 ( .A1(n8399), .A2(n8398), .A3(n8397), .A4(n8396), .ZN(n12557) );
  NAND2_X1 U10815 ( .A1(n11724), .A2(n12557), .ZN(n8777) );
  NAND2_X1 U10816 ( .A1(n14454), .A2(n11731), .ZN(n8778) );
  NAND2_X1 U10817 ( .A1(n11616), .A2(n11615), .ZN(n8400) );
  INV_X1 U10818 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10423) );
  NAND2_X1 U10819 ( .A1(n8406), .A2(n10423), .ZN(n8407) );
  NAND2_X1 U10820 ( .A1(n8424), .A2(n8407), .ZN(n9916) );
  NAND2_X1 U10821 ( .A1(n9916), .A2(n8673), .ZN(n8414) );
  NAND2_X1 U10822 ( .A1(n8391), .A2(n8408), .ZN(n8409) );
  NAND2_X1 U10823 ( .A1(n8409), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8410) );
  MUX2_X1 U10824 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8410), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n8412) );
  NAND2_X1 U10825 ( .A1(n8412), .A2(n8411), .ZN(n15151) );
  AOI22_X1 U10826 ( .A1(n8674), .A2(n9915), .B1(n8518), .B2(n15151), .ZN(n8413) );
  NAND2_X1 U10827 ( .A1(n8414), .A2(n8413), .ZN(n11833) );
  NAND2_X1 U10828 ( .A1(n8538), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8422) );
  INV_X1 U10829 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8415) );
  NOR2_X1 U10830 ( .A1(n8416), .A2(n8415), .ZN(n8417) );
  OR2_X1 U10831 ( .A1(n8436), .A2(n8417), .ZN(n11825) );
  INV_X1 U10832 ( .A(n11825), .ZN(n11834) );
  OR2_X1 U10833 ( .A1(n8651), .A2(n11834), .ZN(n8421) );
  INV_X1 U10834 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n8418) );
  OR2_X1 U10835 ( .A1(n8284), .A2(n8418), .ZN(n8420) );
  INV_X1 U10836 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n11835) );
  OR2_X1 U10837 ( .A1(n6477), .A2(n11835), .ZN(n8419) );
  NOR2_X1 U10838 ( .A1(n11833), .A2(n12556), .ZN(n8782) );
  NAND2_X1 U10839 ( .A1(n11833), .A2(n12556), .ZN(n8699) );
  INV_X1 U10840 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10731) );
  NAND2_X1 U10841 ( .A1(n10731), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8443) );
  INV_X1 U10842 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10735) );
  NAND2_X1 U10843 ( .A1(n10735), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8425) );
  OR2_X1 U10844 ( .A1(n8427), .A2(n8426), .ZN(n8428) );
  NAND2_X1 U10845 ( .A1(n8444), .A2(n8428), .ZN(n9930) );
  NAND2_X1 U10846 ( .A1(n9930), .A2(n8673), .ZN(n8434) );
  NAND2_X1 U10847 ( .A1(n8411), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8429) );
  MUX2_X1 U10848 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8429), .S(
        P3_IR_REG_14__SCAN_IN), .Z(n8432) );
  INV_X1 U10849 ( .A(n8430), .ZN(n8431) );
  NAND2_X1 U10850 ( .A1(n8432), .A2(n8431), .ZN(n15169) );
  AOI22_X1 U10851 ( .A1(n8674), .A2(n9929), .B1(n8518), .B2(n15169), .ZN(n8433) );
  NAND2_X1 U10852 ( .A1(n8661), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8442) );
  INV_X1 U10853 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n8435) );
  NOR2_X1 U10854 ( .A1(n8436), .A2(n8435), .ZN(n8437) );
  OR2_X1 U10855 ( .A1(n8470), .A2(n8437), .ZN(n11876) );
  INV_X1 U10856 ( .A(n11876), .ZN(n14380) );
  OR2_X1 U10857 ( .A1(n8651), .A2(n14380), .ZN(n8441) );
  INV_X1 U10858 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n11871) );
  OR2_X1 U10859 ( .A1(n8679), .A2(n11871), .ZN(n8440) );
  INV_X1 U10860 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n8438) );
  OR2_X1 U10861 ( .A1(n6477), .A2(n8438), .ZN(n8439) );
  NAND4_X1 U10862 ( .A1(n8442), .A2(n8441), .A3(n8440), .A4(n8439), .ZN(n12856) );
  NAND2_X1 U10863 ( .A1(n14374), .A2(n12856), .ZN(n8786) );
  NAND2_X1 U10864 ( .A1(n8785), .A2(n8786), .ZN(n8943) );
  INV_X1 U10865 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10759) );
  NAND2_X1 U10866 ( .A1(n10759), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8460) );
  INV_X1 U10867 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10794) );
  NAND2_X1 U10868 ( .A1(n10794), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8445) );
  AND2_X1 U10869 ( .A1(n8460), .A2(n8445), .ZN(n8446) );
  OR2_X1 U10870 ( .A1(n8447), .A2(n8446), .ZN(n8448) );
  NAND2_X1 U10871 ( .A1(n6495), .A2(n8448), .ZN(n10030) );
  NOR2_X1 U10872 ( .A1(n8430), .A2(n13011), .ZN(n8449) );
  MUX2_X1 U10873 ( .A(n13011), .B(n8449), .S(P3_IR_REG_15__SCAN_IN), .Z(n8451)
         );
  OR2_X1 U10874 ( .A1(n8451), .A2(n8717), .ZN(n14389) );
  INV_X1 U10875 ( .A(n14389), .ZN(n8452) );
  AOI22_X1 U10876 ( .A1(n8674), .A2(SI_15_), .B1(n8518), .B2(n8452), .ZN(n8453) );
  INV_X1 U10877 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14383) );
  OR2_X1 U10878 ( .A1(n6477), .A2(n14383), .ZN(n8458) );
  INV_X1 U10879 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12917) );
  OR2_X1 U10880 ( .A1(n8284), .A2(n12917), .ZN(n8457) );
  XNOR2_X1 U10881 ( .A(n8470), .B(P3_REG3_REG_15__SCAN_IN), .ZN(n12858) );
  OR2_X1 U10882 ( .A1(n8651), .A2(n12858), .ZN(n8456) );
  INV_X1 U10883 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13003) );
  OR2_X1 U10884 ( .A1(n8679), .A2(n13003), .ZN(n8455) );
  OR2_X1 U10885 ( .A1(n13004), .A2(n12476), .ZN(n8789) );
  NAND2_X1 U10886 ( .A1(n13004), .A2(n12476), .ZN(n8793) );
  NAND2_X1 U10887 ( .A1(n8789), .A2(n8793), .ZN(n8946) );
  NAND2_X1 U10888 ( .A1(n8459), .A2(n8793), .ZN(n12841) );
  NAND2_X1 U10889 ( .A1(n10603), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8476) );
  NAND2_X1 U10890 ( .A1(n10732), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8461) );
  AND2_X1 U10891 ( .A1(n8476), .A2(n8461), .ZN(n8462) );
  OR2_X1 U10892 ( .A1(n8463), .A2(n8462), .ZN(n8464) );
  NAND2_X1 U10893 ( .A1(n8477), .A2(n8464), .ZN(n10054) );
  OR2_X1 U10894 ( .A1(n8717), .A2(n13011), .ZN(n8465) );
  XNOR2_X1 U10895 ( .A(n8465), .B(P3_IR_REG_16__SCAN_IN), .ZN(n14399) );
  AOI22_X1 U10896 ( .A1(n8674), .A2(SI_16_), .B1(n8518), .B2(n14399), .ZN(
        n8466) );
  NAND2_X1 U10897 ( .A1(n8538), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8475) );
  INV_X1 U10898 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12846) );
  OR2_X1 U10899 ( .A1(n6477), .A2(n12846), .ZN(n8474) );
  INV_X1 U10900 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12914) );
  OR2_X1 U10901 ( .A1(n8284), .A2(n12914), .ZN(n8473) );
  INV_X1 U10902 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n14386) );
  NAND2_X1 U10903 ( .A1(n8470), .A2(n14386), .ZN(n8468) );
  NAND2_X1 U10904 ( .A1(n8468), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8471) );
  NOR2_X1 U10905 ( .A1(P3_REG3_REG_15__SCAN_IN), .A2(P3_REG3_REG_16__SCAN_IN), 
        .ZN(n8469) );
  AND2_X1 U10906 ( .A1(n8471), .A2(n8483), .ZN(n12847) );
  OR2_X1 U10907 ( .A1(n8651), .A2(n12847), .ZN(n8472) );
  OR2_X1 U10908 ( .A1(n12998), .A2(n12485), .ZN(n8790) );
  NAND2_X1 U10909 ( .A1(n12998), .A2(n12485), .ZN(n8794) );
  NAND2_X1 U10910 ( .A1(n8790), .A2(n8794), .ZN(n8949) );
  NAND2_X1 U10911 ( .A1(n12840), .A2(n8794), .ZN(n12831) );
  NAND2_X1 U10912 ( .A1(n10757), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8493) );
  NAND2_X1 U10913 ( .A1(n10761), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8478) );
  NAND2_X1 U10914 ( .A1(n8493), .A2(n8478), .ZN(n8490) );
  XNOR2_X1 U10915 ( .A(n8492), .B(n8490), .ZN(n10146) );
  NAND2_X1 U10916 ( .A1(n10146), .A2(n8673), .ZN(n8482) );
  INV_X1 U10917 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8479) );
  NAND2_X1 U10918 ( .A1(n8450), .A2(n8479), .ZN(n8495) );
  NAND2_X1 U10919 ( .A1(n8495), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8480) );
  XNOR2_X1 U10920 ( .A(n8480), .B(P3_IR_REG_17__SCAN_IN), .ZN(n14416) );
  AOI22_X1 U10921 ( .A1(n8674), .A2(SI_17_), .B1(n8518), .B2(n14416), .ZN(
        n8481) );
  NAND2_X1 U10922 ( .A1(n8538), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8488) );
  INV_X1 U10923 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14425) );
  OR2_X1 U10924 ( .A1(n6477), .A2(n14425), .ZN(n8487) );
  INV_X1 U10925 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12911) );
  OR2_X1 U10926 ( .A1(n8284), .A2(n12911), .ZN(n8486) );
  NAND2_X1 U10927 ( .A1(n8483), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8484) );
  AND2_X1 U10928 ( .A1(n8501), .A2(n8484), .ZN(n12835) );
  OR2_X1 U10929 ( .A1(n8651), .A2(n12835), .ZN(n8485) );
  OR2_X1 U10930 ( .A1(n12992), .A2(n12371), .ZN(n8802) );
  NAND2_X1 U10931 ( .A1(n12992), .A2(n12371), .ZN(n8807) );
  NAND2_X1 U10932 ( .A1(n8802), .A2(n8807), .ZN(n8952) );
  NAND2_X1 U10933 ( .A1(n12831), .A2(n7345), .ZN(n8489) );
  INV_X1 U10934 ( .A(n8490), .ZN(n8491) );
  INV_X1 U10935 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11068) );
  NAND2_X1 U10936 ( .A1(n11068), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8510) );
  INV_X1 U10937 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11069) );
  NAND2_X1 U10938 ( .A1(n11069), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8494) );
  NAND2_X1 U10939 ( .A1(n8510), .A2(n8494), .ZN(n8507) );
  XNOR2_X1 U10940 ( .A(n8509), .B(n8507), .ZN(n10393) );
  NAND2_X1 U10941 ( .A1(n10393), .A2(n8673), .ZN(n8500) );
  NAND2_X1 U10942 ( .A1(n8497), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8496) );
  MUX2_X1 U10943 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8496), .S(
        P3_IR_REG_18__SCAN_IN), .Z(n8498) );
  NOR2_X2 U10944 ( .A1(n8497), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n8693) );
  INV_X1 U10945 ( .A(n8693), .ZN(n8516) );
  NAND2_X1 U10946 ( .A1(n8498), .A2(n8516), .ZN(n12617) );
  INV_X1 U10947 ( .A(n12617), .ZN(n14431) );
  AOI22_X1 U10948 ( .A1(n8674), .A2(SI_18_), .B1(n8518), .B2(n14431), .ZN(
        n8499) );
  NAND2_X1 U10949 ( .A1(n8636), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8506) );
  INV_X1 U10950 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12908) );
  OR2_X1 U10951 ( .A1(n8284), .A2(n12908), .ZN(n8505) );
  AND2_X1 U10952 ( .A1(n8501), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8502) );
  NOR2_X1 U10953 ( .A1(n8522), .A2(n8502), .ZN(n12826) );
  OR2_X1 U10954 ( .A1(n8651), .A2(n12826), .ZN(n8504) );
  INV_X1 U10955 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12985) );
  OR2_X1 U10956 ( .A1(n8679), .A2(n12985), .ZN(n8503) );
  NAND2_X1 U10957 ( .A1(n12986), .A2(n12807), .ZN(n8806) );
  INV_X1 U10958 ( .A(n8507), .ZN(n8508) );
  NAND2_X1 U10959 ( .A1(n11249), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8528) );
  NAND2_X1 U10960 ( .A1(n11247), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8512) );
  AND2_X1 U10961 ( .A1(n8528), .A2(n8512), .ZN(n8513) );
  OR2_X1 U10962 ( .A1(n8514), .A2(n8513), .ZN(n8515) );
  NAND2_X1 U10963 ( .A1(n8529), .A2(n8515), .ZN(n10421) );
  NAND2_X1 U10964 ( .A1(n10421), .A2(n8673), .ZN(n8520) );
  NAND2_X1 U10965 ( .A1(n8516), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8517) );
  XNOR2_X2 U10966 ( .A(n8517), .B(n8692), .ZN(n12676) );
  AOI22_X1 U10967 ( .A1(n8674), .A2(n10422), .B1(n8518), .B2(n12676), .ZN(
        n8519) );
  INV_X1 U10968 ( .A(n8651), .ZN(n8548) );
  INV_X1 U10969 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n8521) );
  NOR2_X1 U10970 ( .A1(n8522), .A2(n8521), .ZN(n8523) );
  OR2_X1 U10971 ( .A1(n8536), .A2(n8523), .ZN(n12814) );
  NAND2_X1 U10972 ( .A1(n8548), .A2(n12814), .ZN(n8527) );
  INV_X1 U10973 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12811) );
  OR2_X1 U10974 ( .A1(n6477), .A2(n12811), .ZN(n8526) );
  INV_X1 U10975 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12904) );
  OR2_X1 U10976 ( .A1(n8284), .A2(n12904), .ZN(n8525) );
  INV_X1 U10977 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12978) );
  OR2_X1 U10978 ( .A1(n8679), .A2(n12978), .ZN(n8524) );
  NAND4_X1 U10979 ( .A1(n8527), .A2(n8526), .A3(n8525), .A4(n8524), .ZN(n12824) );
  NAND2_X1 U10980 ( .A1(n12982), .A2(n12824), .ZN(n8811) );
  INV_X1 U10981 ( .A(n8811), .ZN(n8804) );
  NAND2_X1 U10982 ( .A1(n8530), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8531) );
  NAND2_X1 U10983 ( .A1(n8542), .A2(n8531), .ZN(n10753) );
  NAND2_X1 U10984 ( .A1(n8674), .A2(SI_20_), .ZN(n8533) );
  INV_X1 U10985 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n8535) );
  OR2_X1 U10986 ( .A1(n8536), .A2(n8535), .ZN(n8537) );
  NAND2_X1 U10987 ( .A1(n8546), .A2(n8537), .ZN(n12799) );
  AOI22_X1 U10988 ( .A1(n12799), .A2(n8548), .B1(n8538), .B2(
        P3_REG0_REG_20__SCAN_IN), .ZN(n8540) );
  AOI22_X1 U10989 ( .A1(n8636), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n8661), .B2(
        P3_REG1_REG_20__SCAN_IN), .ZN(n8539) );
  XNOR2_X1 U10990 ( .A(n12972), .B(n12808), .ZN(n8956) );
  OR2_X1 U10991 ( .A1(n12972), .A2(n12808), .ZN(n8815) );
  NAND2_X1 U10992 ( .A1(n11595), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8556) );
  INV_X1 U10993 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n12417) );
  NAND2_X1 U10994 ( .A1(n12417), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8543) );
  NAND2_X1 U10995 ( .A1(n8556), .A2(n8543), .ZN(n8553) );
  XNOR2_X1 U10996 ( .A(n8555), .B(n8553), .ZN(n10961) );
  NAND2_X1 U10997 ( .A1(n10961), .A2(n8673), .ZN(n8545) );
  NAND2_X1 U10998 ( .A1(n8674), .A2(SI_21_), .ZN(n8544) );
  INV_X1 U10999 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12965) );
  NAND2_X1 U11000 ( .A1(n8546), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8547) );
  NAND2_X1 U11001 ( .A1(n8547), .A2(n7478), .ZN(n12789) );
  NAND2_X1 U11002 ( .A1(n12789), .A2(n8548), .ZN(n8552) );
  INV_X1 U11003 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n12788) );
  OR2_X1 U11004 ( .A1(n6477), .A2(n12788), .ZN(n8550) );
  INV_X1 U11005 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12897) );
  OR2_X1 U11006 ( .A1(n8284), .A2(n12897), .ZN(n8549) );
  AND2_X1 U11007 ( .A1(n8550), .A2(n8549), .ZN(n8551) );
  INV_X1 U11008 ( .A(n12796), .ZN(n12508) );
  NAND2_X1 U11009 ( .A1(n12966), .A2(n12508), .ZN(n8820) );
  OR2_X1 U11010 ( .A1(n12966), .A2(n12508), .ZN(n8819) );
  INV_X1 U11011 ( .A(n8553), .ZN(n8554) );
  INV_X1 U11012 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8557) );
  XNOR2_X1 U11013 ( .A(n8557), .B(P1_DATAO_REG_22__SCAN_IN), .ZN(n8564) );
  XNOR2_X1 U11014 ( .A(n8565), .B(n8564), .ZN(n10965) );
  NAND2_X1 U11015 ( .A1(n10965), .A2(n8673), .ZN(n8559) );
  NAND2_X1 U11016 ( .A1(n8674), .A2(SI_22_), .ZN(n8558) );
  NAND2_X1 U11017 ( .A1(n8636), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8563) );
  INV_X1 U11018 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12894) );
  OR2_X1 U11019 ( .A1(n8284), .A2(n12894), .ZN(n8562) );
  AOI21_X1 U11020 ( .B1(P3_REG3_REG_22__SCAN_IN), .B2(n7478), .A(n8570), .ZN(
        n12779) );
  OR2_X1 U11021 ( .A1(n8651), .A2(n12779), .ZN(n8561) );
  INV_X1 U11022 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12959) );
  OR2_X1 U11023 ( .A1(n8679), .A2(n12959), .ZN(n8560) );
  NAND4_X1 U11024 ( .A1(n8563), .A2(n8562), .A3(n8561), .A4(n8560), .ZN(n12554) );
  INV_X1 U11025 ( .A(n12554), .ZN(n12764) );
  NAND2_X1 U11026 ( .A1(n12960), .A2(n12764), .ZN(n8824) );
  OR2_X1 U11027 ( .A1(n12960), .A2(n12764), .ZN(n8823) );
  INV_X1 U11028 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12067) );
  NAND2_X1 U11029 ( .A1(n12067), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8566) );
  XNOR2_X1 U11030 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8576) );
  XNOR2_X1 U11031 ( .A(n8577), .B(n8576), .ZN(n11151) );
  NAND2_X1 U11032 ( .A1(n11151), .A2(n8673), .ZN(n8568) );
  NAND2_X1 U11033 ( .A1(n8674), .A2(SI_23_), .ZN(n8567) );
  NAND2_X1 U11034 ( .A1(n8661), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8575) );
  INV_X1 U11035 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12768) );
  OR2_X1 U11036 ( .A1(n6477), .A2(n12768), .ZN(n8574) );
  AOI21_X1 U11037 ( .B1(P3_REG3_REG_23__SCAN_IN), .B2(n8571), .A(n8584), .ZN(
        n12769) );
  OR2_X1 U11038 ( .A1(n8651), .A2(n12769), .ZN(n8573) );
  INV_X1 U11039 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12953) );
  OR2_X1 U11040 ( .A1(n8679), .A2(n12953), .ZN(n8572) );
  NAND2_X1 U11041 ( .A1(n12954), .A2(n8961), .ZN(n8829) );
  INV_X1 U11042 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11858) );
  NAND2_X1 U11043 ( .A1(n11858), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8578) );
  INV_X1 U11044 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11862) );
  NAND2_X1 U11045 ( .A1(n8580), .A2(n11862), .ZN(n8581) );
  XNOR2_X1 U11046 ( .A(n8592), .B(n11861), .ZN(n11547) );
  NAND2_X1 U11047 ( .A1(n11547), .A2(n8673), .ZN(n8583) );
  NAND2_X1 U11048 ( .A1(n8674), .A2(SI_24_), .ZN(n8582) );
  NAND2_X1 U11049 ( .A1(n8636), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8589) );
  INV_X1 U11050 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12889) );
  OR2_X1 U11051 ( .A1(n8284), .A2(n12889), .ZN(n8588) );
  AOI21_X1 U11052 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(n8585), .A(n8596), .ZN(
        n12751) );
  OR2_X1 U11053 ( .A1(n8651), .A2(n12751), .ZN(n8587) );
  INV_X1 U11054 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12949) );
  OR2_X1 U11055 ( .A1(n8679), .A2(n12949), .ZN(n8586) );
  NAND4_X1 U11056 ( .A1(n8589), .A2(n8588), .A3(n8587), .A4(n8586), .ZN(n12738) );
  OR2_X1 U11057 ( .A1(n12887), .A2(n12763), .ZN(n8832) );
  NAND2_X1 U11058 ( .A1(n12887), .A2(n12763), .ZN(n8830) );
  INV_X1 U11059 ( .A(n12747), .ZN(n8590) );
  NOR2_X1 U11060 ( .A1(n12754), .A2(n8590), .ZN(n8591) );
  NAND2_X1 U11061 ( .A1(n12746), .A2(n8591), .ZN(n12748) );
  NAND2_X1 U11062 ( .A1(n12748), .A2(n8830), .ZN(n12735) );
  XNOR2_X1 U11063 ( .A(n13706), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8593) );
  XNOR2_X1 U11064 ( .A(n8604), .B(n8593), .ZN(n11590) );
  NAND2_X1 U11065 ( .A1(n11590), .A2(n8673), .ZN(n8595) );
  NAND2_X1 U11066 ( .A1(n8674), .A2(SI_25_), .ZN(n8594) );
  NAND2_X1 U11067 ( .A1(n8636), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8601) );
  INV_X1 U11068 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12883) );
  OR2_X1 U11069 ( .A1(n8284), .A2(n12883), .ZN(n8600) );
  AOI21_X1 U11070 ( .B1(P3_REG3_REG_25__SCAN_IN), .B2(n8597), .A(n8609), .ZN(
        n12742) );
  OR2_X1 U11071 ( .A1(n8651), .A2(n12742), .ZN(n8599) );
  INV_X1 U11072 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12943) );
  OR2_X1 U11073 ( .A1(n8679), .A2(n12943), .ZN(n8598) );
  OR2_X1 U11074 ( .A1(n12944), .A2(n12393), .ZN(n8835) );
  NAND2_X1 U11075 ( .A1(n12944), .A2(n12393), .ZN(n8836) );
  NAND2_X1 U11076 ( .A1(n8835), .A2(n8836), .ZN(n12734) );
  INV_X1 U11077 ( .A(n12734), .ZN(n12737) );
  NAND2_X1 U11078 ( .A1(n12735), .A2(n12737), .ZN(n8602) );
  NAND2_X1 U11079 ( .A1(n8602), .A2(n8836), .ZN(n12724) );
  NAND2_X1 U11080 ( .A1(n13706), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8603) );
  NAND2_X1 U11081 ( .A1(n11910), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8605) );
  XNOR2_X1 U11082 ( .A(n13703), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n8607) );
  XNOR2_X1 U11083 ( .A(n8617), .B(n8607), .ZN(n11694) );
  NAND2_X1 U11084 ( .A1(n8674), .A2(SI_26_), .ZN(n8608) );
  NAND2_X1 U11085 ( .A1(n8636), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8614) );
  INV_X1 U11086 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12881) );
  OR2_X1 U11087 ( .A1(n8284), .A2(n12881), .ZN(n8613) );
  NOR2_X2 U11088 ( .A1(P3_REG3_REG_26__SCAN_IN), .A2(n8610), .ZN(n8623) );
  AOI21_X1 U11089 ( .B1(P3_REG3_REG_26__SCAN_IN), .B2(n8610), .A(n8623), .ZN(
        n12729) );
  OR2_X1 U11090 ( .A1(n8651), .A2(n12729), .ZN(n8612) );
  INV_X1 U11091 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12939) );
  OR2_X1 U11092 ( .A1(n8679), .A2(n12939), .ZN(n8611) );
  NAND2_X1 U11093 ( .A1(n12724), .A2(n8840), .ZN(n8615) );
  NAND2_X1 U11094 ( .A1(n12880), .A2(n8966), .ZN(n8841) );
  NAND2_X1 U11095 ( .A1(n8615), .A2(n8841), .ZN(n12717) );
  AND2_X1 U11096 ( .A1(n14222), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8616) );
  NAND2_X1 U11097 ( .A1(n13703), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8618) );
  XNOR2_X1 U11098 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n8620) );
  XNOR2_X1 U11099 ( .A(n8631), .B(n8620), .ZN(n11760) );
  NAND2_X1 U11100 ( .A1(n11760), .A2(n8673), .ZN(n8622) );
  NAND2_X1 U11101 ( .A1(n8674), .A2(SI_27_), .ZN(n8621) );
  NAND2_X1 U11102 ( .A1(n8636), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8629) );
  INV_X1 U11103 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12877) );
  OR2_X1 U11104 ( .A1(n8284), .A2(n12877), .ZN(n8628) );
  INV_X1 U11105 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n12439) );
  NAND2_X1 U11106 ( .A1(n12439), .A2(n8623), .ZN(n8639) );
  INV_X1 U11107 ( .A(n8623), .ZN(n8624) );
  NAND2_X1 U11108 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(n8624), .ZN(n8625) );
  AND2_X1 U11109 ( .A1(n8639), .A2(n8625), .ZN(n12437) );
  INV_X1 U11110 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12935) );
  OR2_X1 U11111 ( .A1(n6475), .A2(n12935), .ZN(n8626) );
  NAND2_X1 U11112 ( .A1(n12433), .A2(n12406), .ZN(n8847) );
  NAND2_X1 U11113 ( .A1(n12715), .A2(n8847), .ZN(n12700) );
  AND2_X1 U11114 ( .A1(n13700), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8630) );
  NAND2_X1 U11115 ( .A1(n14220), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8632) );
  XNOR2_X1 U11116 ( .A(n13698), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n8633) );
  XNOR2_X1 U11117 ( .A(n8646), .B(n8633), .ZN(n12325) );
  NAND2_X1 U11118 ( .A1(n12325), .A2(n8673), .ZN(n8635) );
  NAND2_X1 U11119 ( .A1(n8674), .A2(SI_28_), .ZN(n8634) );
  NAND2_X1 U11120 ( .A1(n8636), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8645) );
  INV_X1 U11121 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12871) );
  OR2_X1 U11122 ( .A1(n8284), .A2(n12871), .ZN(n8644) );
  INV_X1 U11123 ( .A(n8639), .ZN(n8638) );
  INV_X1 U11124 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n8637) );
  NAND2_X1 U11125 ( .A1(n8638), .A2(n8637), .ZN(n12685) );
  NAND2_X1 U11126 ( .A1(n8639), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8640) );
  INV_X1 U11127 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n8641) );
  OR2_X1 U11128 ( .A1(n8679), .A2(n8641), .ZN(n8642) );
  NAND2_X1 U11129 ( .A1(n12872), .A2(n8980), .ZN(n8848) );
  NAND2_X1 U11130 ( .A1(n12700), .A2(n12699), .ZN(n12698) );
  NAND2_X1 U11131 ( .A1(n13698), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8647) );
  XNOR2_X1 U11132 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n8655) );
  XNOR2_X1 U11133 ( .A(n8657), .B(n8655), .ZN(n13017) );
  NAND2_X1 U11134 ( .A1(n13017), .A2(n8673), .ZN(n8650) );
  NAND2_X1 U11135 ( .A1(n8674), .A2(SI_29_), .ZN(n8649) );
  INV_X1 U11136 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9014) );
  OR2_X1 U11137 ( .A1(n8284), .A2(n9014), .ZN(n8654) );
  INV_X1 U11138 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9030) );
  OR2_X1 U11139 ( .A1(n8679), .A2(n9030), .ZN(n8653) );
  INV_X1 U11140 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n12692) );
  OR2_X1 U11141 ( .A1(n6477), .A2(n12692), .ZN(n8652) );
  INV_X1 U11142 ( .A(n8655), .ZN(n8656) );
  INV_X1 U11143 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13691) );
  XNOR2_X1 U11144 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n8667) );
  INV_X1 U11145 ( .A(n8667), .ZN(n8658) );
  XNOR2_X1 U11146 ( .A(n8668), .B(n8658), .ZN(n12413) );
  NAND2_X1 U11147 ( .A1(n12413), .A2(n8673), .ZN(n8660) );
  NAND2_X1 U11148 ( .A1(n8674), .A2(SI_30_), .ZN(n8659) );
  INV_X1 U11149 ( .A(n12925), .ZN(n12689) );
  NAND2_X1 U11150 ( .A1(n8661), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n8666) );
  INV_X1 U11151 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n8662) );
  OR2_X1 U11152 ( .A1(n6477), .A2(n8662), .ZN(n8665) );
  INV_X1 U11153 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n8663) );
  OR2_X1 U11154 ( .A1(n6475), .A2(n8663), .ZN(n8664) );
  NAND4_X1 U11155 ( .A1(n8683), .A2(n8666), .A3(n8665), .A4(n8664), .ZN(n12683) );
  NOR2_X1 U11156 ( .A1(n12689), .A2(n12683), .ZN(n8686) );
  NAND2_X1 U11157 ( .A1(n8668), .A2(n8667), .ZN(n8670) );
  INV_X1 U11158 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14217) );
  NAND2_X1 U11159 ( .A1(n14217), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8669) );
  NAND2_X1 U11160 ( .A1(n8670), .A2(n8669), .ZN(n8672) );
  INV_X1 U11161 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13686) );
  XNOR2_X1 U11162 ( .A(n13686), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n8671) );
  NAND2_X1 U11163 ( .A1(n8674), .A2(SI_31_), .ZN(n8675) );
  INV_X1 U11164 ( .A(n12683), .ZN(n8687) );
  INV_X1 U11165 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n8676) );
  OR2_X1 U11166 ( .A1(n6477), .A2(n8676), .ZN(n8682) );
  INV_X1 U11167 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n8677) );
  OR2_X1 U11168 ( .A1(n8284), .A2(n8677), .ZN(n8681) );
  INV_X1 U11169 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n8678) );
  OR2_X1 U11170 ( .A1(n8679), .A2(n8678), .ZN(n8680) );
  NAND2_X1 U11171 ( .A1(n12694), .A2(n12405), .ZN(n8971) );
  INV_X1 U11172 ( .A(n8971), .ZN(n8684) );
  AOI21_X1 U11173 ( .B1(n12925), .B2(n11149), .A(n8684), .ZN(n8685) );
  NAND2_X1 U11174 ( .A1(n12681), .A2(n8687), .ZN(n8689) );
  OR2_X1 U11175 ( .A1(n12925), .A2(n11149), .ZN(n8688) );
  INV_X1 U11176 ( .A(n12676), .ZN(n9020) );
  NAND2_X1 U11177 ( .A1(n8693), .A2(n8692), .ZN(n8696) );
  INV_X1 U11178 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8694) );
  XNOR2_X2 U11179 ( .A(n8697), .B(P3_IR_REG_20__SCAN_IN), .ZN(n10627) );
  NAND2_X1 U11180 ( .A1(n11013), .A2(n10627), .ZN(n8975) );
  INV_X1 U11181 ( .A(n8972), .ZN(n8712) );
  INV_X1 U11182 ( .A(n12761), .ZN(n8698) );
  NOR2_X1 U11183 ( .A1(n12754), .A2(n8698), .ZN(n8826) );
  INV_X1 U11184 ( .A(n8826), .ZN(n8709) );
  XNOR2_X1 U11185 ( .A(n12966), .B(n12796), .ZN(n12785) );
  INV_X1 U11186 ( .A(n12785), .ZN(n8708) );
  NAND2_X1 U11187 ( .A1(n8810), .A2(n8811), .ZN(n12812) );
  INV_X1 U11188 ( .A(n8943), .ZN(n11868) );
  OR2_X1 U11189 ( .A1(n8782), .A2(n7001), .ZN(n11830) );
  INV_X1 U11190 ( .A(n11830), .ZN(n11828) );
  INV_X1 U11191 ( .A(n11615), .ZN(n8703) );
  XNOR2_X1 U11192 ( .A(n12559), .B(n11524), .ZN(n11519) );
  INV_X1 U11193 ( .A(n15255), .ZN(n10635) );
  AND2_X1 U11194 ( .A1(n15257), .A2(n10649), .ZN(n8722) );
  INV_X1 U11195 ( .A(n8722), .ZN(n8721) );
  NAND2_X1 U11196 ( .A1(n10635), .A2(n8721), .ZN(n10651) );
  NOR4_X1 U11197 ( .A1(n15192), .A2(n10651), .A3(n15219), .A4(n15261), .ZN(
        n8701) );
  NOR4_X1 U11198 ( .A1(n11386), .A2(n15205), .A3(n11018), .A4(n15231), .ZN(
        n8700) );
  XNOR2_X1 U11199 ( .A(n12560), .B(n11459), .ZN(n8935) );
  INV_X1 U11200 ( .A(n8935), .ZN(n11455) );
  NAND4_X1 U11201 ( .A1(n8701), .A2(n8700), .A3(n11455), .A4(n11397), .ZN(
        n8702) );
  NOR4_X1 U11202 ( .A1(n8703), .A2(n11519), .A3(n8702), .A4(n14451), .ZN(n8704) );
  NAND4_X1 U11203 ( .A1(n12854), .A2(n11868), .A3(n11828), .A4(n8704), .ZN(
        n8705) );
  NOR4_X1 U11204 ( .A1(n12812), .A2(n8952), .A3(n8705), .A4(n8949), .ZN(n8706)
         );
  NAND4_X1 U11205 ( .A1(n12774), .A2(n12821), .A3(n8706), .A4(n12794), .ZN(
        n8707) );
  NOR4_X1 U11206 ( .A1(n8709), .A2(n12734), .A3(n8708), .A4(n8707), .ZN(n8710)
         );
  NAND4_X1 U11207 ( .A1(n12699), .A2(n12716), .A3(n12726), .A4(n8710), .ZN(
        n8711) );
  XNOR2_X1 U11208 ( .A(n8713), .B(n12676), .ZN(n8715) );
  NAND2_X1 U11209 ( .A1(n10964), .A2(n10627), .ZN(n10625) );
  INV_X1 U11210 ( .A(n15267), .ZN(n15237) );
  INV_X1 U11211 ( .A(n10626), .ZN(n10620) );
  NAND2_X1 U11212 ( .A1(n8719), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8718) );
  MUX2_X1 U11213 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8718), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n8720) );
  NAND2_X1 U11214 ( .A1(n8720), .A2(n8863), .ZN(n9022) );
  OAI211_X1 U11215 ( .C1(n15255), .C2(n11013), .A(n8721), .B(n10430), .ZN(
        n8728) );
  INV_X1 U11216 ( .A(n15230), .ZN(n8724) );
  OAI22_X1 U11217 ( .A1(n8722), .A2(n15261), .B1(n8724), .B2(n8978), .ZN(n8727) );
  INV_X1 U11218 ( .A(n8723), .ZN(n8725) );
  MUX2_X1 U11219 ( .A(n8725), .B(n8724), .S(n8978), .Z(n8726) );
  AOI21_X1 U11220 ( .B1(n8743), .B2(n8729), .A(n10430), .ZN(n8742) );
  OAI21_X1 U11221 ( .B1(n8738), .B2(n8742), .A(n8740), .ZN(n8737) );
  MUX2_X1 U11222 ( .A(n8731), .B(n8730), .S(n8978), .Z(n8732) );
  INV_X1 U11223 ( .A(n8732), .ZN(n8733) );
  NOR2_X1 U11224 ( .A1(n8733), .A2(n15205), .ZN(n8746) );
  INV_X1 U11225 ( .A(n8755), .ZN(n8736) );
  INV_X1 U11226 ( .A(n8734), .ZN(n8735) );
  AOI211_X1 U11227 ( .C1(n8737), .C2(n8746), .A(n8736), .B(n8735), .ZN(n8749)
         );
  INV_X1 U11228 ( .A(n8738), .ZN(n8741) );
  NAND3_X1 U11229 ( .A1(n8741), .A2(n8740), .A3(n8739), .ZN(n8744) );
  AOI21_X1 U11230 ( .B1(n8744), .B2(n8743), .A(n8742), .ZN(n8745) );
  NOR2_X1 U11231 ( .A1(n8745), .A2(n11018), .ZN(n8748) );
  INV_X1 U11232 ( .A(n8746), .ZN(n8747) );
  OAI22_X1 U11233 ( .A1(n8749), .A2(n10430), .B1(n8748), .B2(n8747), .ZN(n8753) );
  AOI21_X1 U11234 ( .B1(n8752), .B2(n8750), .A(n8978), .ZN(n8751) );
  AOI21_X1 U11235 ( .B1(n8753), .B2(n8752), .A(n8751), .ZN(n8760) );
  OAI21_X1 U11236 ( .B1(n8978), .B2(n8755), .A(n8754), .ZN(n8759) );
  MUX2_X1 U11237 ( .A(n8757), .B(n8756), .S(n8978), .Z(n8758) );
  OAI211_X1 U11238 ( .C1(n8760), .C2(n8759), .A(n11397), .B(n8758), .ZN(n8764)
         );
  NAND2_X1 U11239 ( .A1(n12561), .A2(n11402), .ZN(n8761) );
  MUX2_X1 U11240 ( .A(n8762), .B(n8761), .S(n8978), .Z(n8763) );
  NAND3_X1 U11241 ( .A1(n8764), .A2(n11455), .A3(n8763), .ZN(n8769) );
  INV_X1 U11242 ( .A(n8765), .ZN(n8766) );
  MUX2_X1 U11243 ( .A(n8767), .B(n8766), .S(n8978), .Z(n8768) );
  AOI21_X1 U11244 ( .B1(n8769), .B2(n8768), .A(n11519), .ZN(n8772) );
  MUX2_X1 U11245 ( .A(n8978), .B(n12559), .S(n11408), .Z(n8770) );
  AOI21_X1 U11246 ( .B1(n14453), .B2(n10430), .A(n8770), .ZN(n8771) );
  NAND2_X1 U11247 ( .A1(n8778), .A2(n8773), .ZN(n8776) );
  NAND2_X1 U11248 ( .A1(n8777), .A2(n8774), .ZN(n8775) );
  MUX2_X1 U11249 ( .A(n8776), .B(n8775), .S(n8978), .Z(n8780) );
  MUX2_X1 U11250 ( .A(n8778), .B(n8777), .S(n10430), .Z(n8779) );
  OAI21_X1 U11251 ( .B1(n8781), .B2(n8780), .A(n8779), .ZN(n8784) );
  MUX2_X1 U11252 ( .A(n8782), .B(n7001), .S(n10430), .Z(n8783) );
  AOI21_X1 U11253 ( .B1(n8784), .B2(n11828), .A(n8783), .ZN(n8788) );
  MUX2_X1 U11254 ( .A(n8786), .B(n8785), .S(n8978), .Z(n8787) );
  OAI21_X1 U11255 ( .B1(n8788), .B2(n8943), .A(n8787), .ZN(n8792) );
  AOI21_X1 U11256 ( .B1(n8790), .B2(n8789), .A(n8978), .ZN(n8791) );
  AOI21_X1 U11257 ( .B1(n8792), .B2(n12854), .A(n8791), .ZN(n8797) );
  INV_X1 U11258 ( .A(n8794), .ZN(n8796) );
  AND2_X1 U11259 ( .A1(n8794), .A2(n8793), .ZN(n8795) );
  OAI22_X1 U11260 ( .A1(n8797), .A2(n8796), .B1(n8795), .B2(n10430), .ZN(n8800) );
  INV_X1 U11261 ( .A(n12998), .ZN(n8798) );
  NAND3_X1 U11262 ( .A1(n8798), .A2(n8978), .A3(n12855), .ZN(n8799) );
  AOI211_X1 U11263 ( .C1(n8800), .C2(n8799), .A(n8952), .B(n12823), .ZN(n8814)
         );
  INV_X1 U11264 ( .A(n8806), .ZN(n8801) );
  AOI21_X1 U11265 ( .B1(n8803), .B2(n8802), .A(n8801), .ZN(n8805) );
  OR2_X1 U11266 ( .A1(n8805), .A2(n8804), .ZN(n8809) );
  OAI211_X1 U11267 ( .C1(n12823), .C2(n8807), .A(n8806), .B(n8810), .ZN(n8808)
         );
  MUX2_X1 U11268 ( .A(n8809), .B(n8808), .S(n10430), .Z(n8813) );
  MUX2_X1 U11269 ( .A(n8811), .B(n8810), .S(n8978), .Z(n8812) );
  OAI211_X1 U11270 ( .C1(n8814), .C2(n8813), .A(n12794), .B(n8812), .ZN(n8818)
         );
  NAND2_X1 U11271 ( .A1(n12972), .A2(n12808), .ZN(n8816) );
  MUX2_X1 U11272 ( .A(n8816), .B(n8815), .S(n8978), .Z(n8817) );
  NAND3_X1 U11273 ( .A1(n8818), .A2(n12785), .A3(n8817), .ZN(n8822) );
  MUX2_X1 U11274 ( .A(n8820), .B(n8819), .S(n10430), .Z(n8821) );
  NAND3_X1 U11275 ( .A1(n8822), .A2(n12774), .A3(n8821), .ZN(n8827) );
  MUX2_X1 U11276 ( .A(n8824), .B(n8823), .S(n8978), .Z(n8825) );
  NAND3_X1 U11277 ( .A1(n8827), .A2(n8826), .A3(n8825), .ZN(n8828) );
  NAND2_X1 U11278 ( .A1(n8828), .A2(n12737), .ZN(n8839) );
  OAI21_X1 U11279 ( .B1(n12754), .B2(n8829), .A(n8830), .ZN(n8834) );
  INV_X1 U11280 ( .A(n8830), .ZN(n8831) );
  AOI21_X1 U11281 ( .B1(n12747), .B2(n8832), .A(n8831), .ZN(n8833) );
  MUX2_X1 U11282 ( .A(n8834), .B(n8833), .S(n10430), .Z(n8838) );
  MUX2_X1 U11283 ( .A(n8836), .B(n8835), .S(n8978), .Z(n8837) );
  OAI211_X1 U11284 ( .C1(n8839), .C2(n8838), .A(n12726), .B(n8837), .ZN(n8843)
         );
  MUX2_X1 U11285 ( .A(n8841), .B(n8840), .S(n10430), .Z(n8842) );
  AOI21_X1 U11286 ( .B1(n8843), .B2(n8842), .A(n8969), .ZN(n8846) );
  INV_X1 U11287 ( .A(n8844), .ZN(n8845) );
  OAI21_X1 U11288 ( .B1(n8846), .B2(n8845), .A(n12699), .ZN(n8851) );
  INV_X1 U11289 ( .A(n8846), .ZN(n8849) );
  NAND3_X1 U11290 ( .A1(n8849), .A2(n8848), .A3(n8847), .ZN(n8850) );
  INV_X1 U11291 ( .A(n8853), .ZN(n8856) );
  NAND2_X1 U11292 ( .A1(n8863), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8861) );
  XNOR2_X1 U11293 ( .A(n8861), .B(n8860), .ZN(n10606) );
  OR2_X1 U11294 ( .A1(n10606), .A2(P3_U3151), .ZN(n11152) );
  INV_X1 U11295 ( .A(n12328), .ZN(n10441) );
  INV_X1 U11296 ( .A(n12670), .ZN(n10445) );
  NAND2_X1 U11297 ( .A1(n10441), .A2(n10445), .ZN(n10433) );
  NAND2_X1 U11298 ( .A1(n10433), .A2(n10431), .ZN(n8977) );
  INV_X1 U11299 ( .A(n8985), .ZN(n8869) );
  NAND2_X1 U11300 ( .A1(n8866), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8867) );
  INV_X1 U11301 ( .A(n11697), .ZN(n8868) );
  INV_X1 U11302 ( .A(n11593), .ZN(n8873) );
  INV_X1 U11303 ( .A(n10619), .ZN(n10641) );
  OAI21_X1 U11304 ( .B1(n11152), .B2(n10966), .A(P3_B_REG_SCAN_IN), .ZN(n8875)
         );
  INV_X1 U11305 ( .A(n8875), .ZN(n8876) );
  NAND2_X1 U11306 ( .A1(n8879), .A2(n8878), .ZN(n8886) );
  NAND2_X1 U11307 ( .A1(n8881), .A2(n8880), .ZN(n8883) );
  INV_X1 U11308 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n11929) );
  MUX2_X1 U11309 ( .A(n11929), .B(n13691), .S(n6533), .Z(n9738) );
  XNOR2_X1 U11310 ( .A(n9738), .B(SI_29_), .ZN(n9736) );
  NAND2_X1 U11311 ( .A1(n11928), .A2(n12260), .ZN(n8885) );
  OR2_X1 U11312 ( .A1(n7673), .A2(n11929), .ZN(n8884) );
  INV_X1 U11313 ( .A(n12344), .ZN(n12336) );
  INV_X1 U11314 ( .A(n6538), .ZN(n9977) );
  AOI21_X1 U11315 ( .B1(n9977), .B2(P1_B_REG_SCAN_IN), .A(n14694), .ZN(n13921)
         );
  INV_X1 U11316 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8892) );
  NAND2_X1 U11317 ( .A1(n7662), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8891) );
  NAND2_X1 U11318 ( .A1(n8889), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8890) );
  OAI211_X1 U11319 ( .C1(n12241), .C2(n8892), .A(n8891), .B(n8890), .ZN(n13841) );
  NAND2_X1 U11320 ( .A1(n13921), .A2(n13841), .ZN(n8909) );
  NAND2_X1 U11321 ( .A1(n13843), .A2(n14596), .ZN(n8902) );
  NAND2_X1 U11322 ( .A1(n8909), .A2(n8902), .ZN(n8894) );
  NOR2_X2 U11323 ( .A1(n8893), .A2(n12231), .ZN(n13926) );
  AOI211_X1 U11324 ( .C1(n12231), .C2(n8893), .A(n14792), .B(n13926), .ZN(
        n8915) );
  AND3_X1 U11325 ( .A1(n8908), .A2(n10061), .A3(n10058), .ZN(n8896) );
  NOR2_X1 U11326 ( .A1(n10057), .A2(n12321), .ZN(n8895) );
  NAND2_X1 U11327 ( .A1(n8921), .A2(n14811), .ZN(n8899) );
  NAND2_X1 U11328 ( .A1(n8899), .A2(n8898), .ZN(P1_U3557) );
  INV_X1 U11329 ( .A(n8908), .ZN(n10060) );
  NAND2_X1 U11330 ( .A1(n8907), .A2(n10060), .ZN(n8901) );
  INV_X1 U11331 ( .A(n10061), .ZN(n8900) );
  INV_X1 U11332 ( .A(n8904), .ZN(n14504) );
  INV_X1 U11333 ( .A(n8905), .ZN(n14509) );
  NAND2_X1 U11334 ( .A1(n14721), .A2(n14509), .ZN(n14103) );
  NOR2_X1 U11335 ( .A1(n14719), .A2(n8906), .ZN(n8912) );
  INV_X1 U11336 ( .A(n8907), .ZN(n8910) );
  NOR3_X1 U11337 ( .A1(n8910), .A2(n8909), .A3(n8908), .ZN(n8911) );
  AOI211_X1 U11338 ( .C1(n14736), .C2(P1_REG2_REG_29__SCAN_IN), .A(n8912), .B(
        n8911), .ZN(n8913) );
  OAI21_X1 U11339 ( .B1(n12232), .B2(n14103), .A(n8913), .ZN(n8914) );
  AOI21_X1 U11340 ( .B1(n8915), .B2(n14731), .A(n8914), .ZN(n8916) );
  NAND2_X1 U11341 ( .A1(n8920), .A2(n8919), .ZN(P1_U3356) );
  NAND2_X1 U11342 ( .A1(n8921), .A2(n14799), .ZN(n8923) );
  NAND2_X1 U11343 ( .A1(n8923), .A2(n8922), .ZN(P1_U3525) );
  NAND2_X1 U11344 ( .A1(n15257), .A2(n10511), .ZN(n15260) );
  NAND2_X1 U11345 ( .A1(n15261), .A2(n15260), .ZN(n8925) );
  INV_X1 U11346 ( .A(n12564), .ZN(n15244) );
  NAND2_X1 U11347 ( .A1(n15244), .A2(n15254), .ZN(n8924) );
  NAND2_X1 U11348 ( .A1(n8925), .A2(n8924), .ZN(n15240) );
  INV_X1 U11349 ( .A(n15235), .ZN(n10708) );
  NOR2_X1 U11350 ( .A1(n15258), .A2(n10708), .ZN(n8926) );
  AOI21_X1 U11351 ( .B1(n15240), .B2(n15231), .A(n8926), .ZN(n15220) );
  NAND2_X1 U11352 ( .A1(n15220), .A2(n15219), .ZN(n15218) );
  INV_X1 U11353 ( .A(n15224), .ZN(n10718) );
  NAND2_X1 U11354 ( .A1(n11016), .A2(n10718), .ZN(n8927) );
  NAND2_X1 U11355 ( .A1(n15218), .A2(n8927), .ZN(n11019) );
  NAND2_X1 U11356 ( .A1(n11019), .A2(n11018), .ZN(n11017) );
  INV_X1 U11357 ( .A(n8928), .ZN(n11014) );
  NAND2_X1 U11358 ( .A1(n15217), .A2(n11014), .ZN(n8929) );
  INV_X1 U11359 ( .A(n15189), .ZN(n11027) );
  NAND2_X1 U11360 ( .A1(n11027), .A2(n15210), .ZN(n8930) );
  INV_X1 U11361 ( .A(n15196), .ZN(n11029) );
  NAND2_X1 U11362 ( .A1(n12562), .A2(n11029), .ZN(n8931) );
  INV_X1 U11363 ( .A(n11391), .ZN(n11336) );
  NAND2_X1 U11364 ( .A1(n15190), .A2(n11336), .ZN(n8932) );
  NAND2_X2 U11365 ( .A1(n11385), .A2(n8932), .ZN(n11396) );
  NAND2_X1 U11366 ( .A1(n11452), .A2(n11402), .ZN(n8933) );
  NAND2_X1 U11367 ( .A1(n12561), .A2(n7322), .ZN(n8934) );
  INV_X1 U11368 ( .A(n11459), .ZN(n11327) );
  NAND2_X1 U11369 ( .A1(n11518), .A2(n11519), .ZN(n8937) );
  NAND2_X1 U11370 ( .A1(n12559), .A2(n11408), .ZN(n8936) );
  AND2_X1 U11371 ( .A1(n12558), .A2(n11641), .ZN(n8939) );
  INV_X1 U11372 ( .A(n12558), .ZN(n11727) );
  NAND2_X1 U11373 ( .A1(n11727), .A2(n14455), .ZN(n8938) );
  NAND2_X1 U11374 ( .A1(n11833), .A2(n12363), .ZN(n8940) );
  NAND2_X1 U11375 ( .A1(n11831), .A2(n8940), .ZN(n8942) );
  OR2_X1 U11376 ( .A1(n11833), .A2(n12363), .ZN(n8941) );
  NAND2_X1 U11377 ( .A1(n8942), .A2(n8941), .ZN(n11865) );
  NAND2_X1 U11378 ( .A1(n11865), .A2(n8943), .ZN(n8945) );
  INV_X1 U11379 ( .A(n12856), .ZN(n12542) );
  OR2_X1 U11380 ( .A1(n14374), .A2(n12542), .ZN(n8944) );
  NAND2_X1 U11381 ( .A1(n8945), .A2(n8944), .ZN(n12853) );
  NAND2_X1 U11382 ( .A1(n12853), .A2(n8946), .ZN(n8948) );
  NAND2_X1 U11383 ( .A1(n13004), .A2(n7302), .ZN(n8947) );
  NAND2_X1 U11384 ( .A1(n8948), .A2(n8947), .ZN(n12842) );
  NAND2_X1 U11385 ( .A1(n12842), .A2(n8949), .ZN(n8951) );
  NAND2_X1 U11386 ( .A1(n12998), .A2(n12855), .ZN(n8950) );
  NAND2_X1 U11387 ( .A1(n8951), .A2(n8950), .ZN(n12832) );
  INV_X1 U11388 ( .A(n12371), .ZN(n12844) );
  NAND2_X1 U11389 ( .A1(n12992), .A2(n12844), .ZN(n8953) );
  OR2_X1 U11390 ( .A1(n12986), .A2(n12833), .ZN(n12804) );
  AND2_X1 U11391 ( .A1(n12812), .A2(n12804), .ZN(n8954) );
  INV_X1 U11392 ( .A(n12824), .ZN(n12376) );
  OR2_X1 U11393 ( .A1(n12982), .A2(n12376), .ZN(n8955) );
  NAND2_X1 U11394 ( .A1(n12802), .A2(n8955), .ZN(n12795) );
  INV_X1 U11395 ( .A(n12808), .ZN(n12555) );
  NAND2_X1 U11396 ( .A1(n12972), .A2(n12555), .ZN(n8957) );
  OR2_X1 U11397 ( .A1(n12966), .A2(n12796), .ZN(n8958) );
  AND2_X1 U11398 ( .A1(n12960), .A2(n12554), .ZN(n8960) );
  OR2_X1 U11399 ( .A1(n12960), .A2(n12554), .ZN(n8959) );
  NAND2_X1 U11400 ( .A1(n12954), .A2(n12776), .ZN(n8962) );
  OR2_X1 U11401 ( .A1(n12887), .A2(n12738), .ZN(n8963) );
  NAND2_X1 U11402 ( .A1(n12736), .A2(n12734), .ZN(n8965) );
  NAND2_X1 U11403 ( .A1(n12944), .A2(n12553), .ZN(n8964) );
  OR2_X1 U11404 ( .A1(n12880), .A2(n12739), .ZN(n8967) );
  NOR2_X1 U11405 ( .A1(n12433), .A2(n12552), .ZN(n8968) );
  INV_X1 U11406 ( .A(n8980), .ZN(n12438) );
  NAND2_X1 U11407 ( .A1(n8972), .A2(n8971), .ZN(n9016) );
  NAND2_X1 U11408 ( .A1(n9020), .A2(n10966), .ZN(n9023) );
  NAND2_X1 U11409 ( .A1(n10441), .A2(P3_B_REG_SCAN_IN), .ZN(n8979) );
  NAND2_X1 U11410 ( .A1(n15259), .A2(n8979), .ZN(n12682) );
  XNOR2_X1 U11411 ( .A(n8985), .B(P3_B_REG_SCAN_IN), .ZN(n8986) );
  AOI21_X1 U11412 ( .B1(n8986), .B2(n11593), .A(n11697), .ZN(n8989) );
  INV_X1 U11413 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n8987) );
  NAND2_X1 U11414 ( .A1(n8985), .A2(n11697), .ZN(n8988) );
  INV_X1 U11415 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8990) );
  NAND2_X1 U11416 ( .A1(n8989), .A2(n8990), .ZN(n8992) );
  NAND2_X1 U11417 ( .A1(n11593), .A2(n11697), .ZN(n8991) );
  XNOR2_X1 U11418 ( .A(n10624), .B(n10505), .ZN(n9004) );
  NOR2_X1 U11419 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n8996) );
  NOR4_X1 U11420 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n8995) );
  NOR4_X1 U11421 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n8994) );
  NOR4_X1 U11422 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8993) );
  NAND4_X1 U11423 ( .A1(n8996), .A2(n8995), .A3(n8994), .A4(n8993), .ZN(n9002)
         );
  NOR4_X1 U11424 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n9000) );
  NOR4_X1 U11425 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n8999) );
  NOR4_X1 U11426 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8998) );
  NOR4_X1 U11427 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8997) );
  NAND4_X1 U11428 ( .A1(n9000), .A2(n8999), .A3(n8998), .A4(n8997), .ZN(n9001)
         );
  OAI21_X1 U11429 ( .B1(n9002), .B2(n9001), .A(n8989), .ZN(n9025) );
  NAND2_X1 U11430 ( .A1(n9025), .A2(n10619), .ZN(n9003) );
  NAND2_X1 U11431 ( .A1(n12676), .A2(n10966), .ZN(n9008) );
  OAI21_X1 U11432 ( .B1(n15253), .B2(n10627), .A(n9008), .ZN(n9005) );
  NAND2_X1 U11433 ( .A1(n9005), .A2(n10626), .ZN(n9006) );
  NAND2_X1 U11434 ( .A1(n9006), .A2(n10430), .ZN(n9007) );
  NAND2_X1 U11435 ( .A1(n9007), .A2(n10505), .ZN(n9012) );
  INV_X1 U11436 ( .A(n10505), .ZN(n9908) );
  OR2_X1 U11437 ( .A1(n10430), .A2(n10620), .ZN(n10609) );
  INV_X1 U11438 ( .A(n9008), .ZN(n9009) );
  NAND2_X1 U11439 ( .A1(n10627), .A2(n9009), .ZN(n9010) );
  NAND2_X1 U11440 ( .A1(n10430), .A2(n9010), .ZN(n10501) );
  NAND2_X1 U11441 ( .A1(n10609), .A2(n10501), .ZN(n10502) );
  NAND2_X1 U11442 ( .A1(n9908), .A2(n10502), .ZN(n9011) );
  NAND2_X1 U11443 ( .A1(n9012), .A2(n9011), .ZN(n9013) );
  NAND2_X1 U11444 ( .A1(n10964), .A2(n10755), .ZN(n9017) );
  XNOR2_X1 U11445 ( .A(n9017), .B(n10966), .ZN(n9019) );
  NAND2_X1 U11446 ( .A1(n10964), .A2(n12676), .ZN(n9018) );
  NAND2_X1 U11447 ( .A1(n9019), .A2(n9018), .ZN(n10604) );
  NAND2_X1 U11448 ( .A1(n10604), .A2(n15253), .ZN(n10638) );
  MUX2_X1 U11449 ( .A(n9022), .B(n10638), .S(n10755), .Z(n9021) );
  NAND2_X1 U11450 ( .A1(n15237), .A2(n9022), .ZN(n15275) );
  NAND2_X1 U11451 ( .A1(n15266), .A2(n15275), .ZN(n15293) );
  NAND2_X1 U11452 ( .A1(n15331), .A2(n15293), .ZN(n12903) );
  INV_X1 U11453 ( .A(n10624), .ZN(n9902) );
  NAND3_X1 U11454 ( .A1(n9908), .A2(n9902), .A3(n9025), .ZN(n10605) );
  OR2_X1 U11455 ( .A1(n10605), .A2(n10641), .ZN(n10639) );
  OR2_X1 U11456 ( .A1(n10430), .A2(n10626), .ZN(n10614) );
  OR2_X1 U11457 ( .A1(n10625), .A2(n9023), .ZN(n10640) );
  AND2_X1 U11458 ( .A1(n10614), .A2(n10640), .ZN(n9024) );
  OR2_X1 U11459 ( .A1(n10639), .A2(n9024), .ZN(n9028) );
  NAND3_X1 U11460 ( .A1(n10505), .A2(n10624), .A3(n9025), .ZN(n10642) );
  NAND2_X1 U11461 ( .A1(n10604), .A2(n10619), .ZN(n9026) );
  NAND2_X1 U11462 ( .A1(n15318), .A2(n15293), .ZN(n12975) );
  NAND2_X1 U11463 ( .A1(n9032), .A2(n9031), .ZN(P3_U3456) );
  NAND2_X1 U11464 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n9033) );
  NAND2_X1 U11465 ( .A1(n9210), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n9223) );
  INV_X1 U11466 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9222) );
  INV_X1 U11467 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n11567) );
  INV_X1 U11468 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9304) );
  NAND2_X1 U11469 ( .A1(n9303), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9334) );
  INV_X1 U11470 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n12070) );
  INV_X1 U11471 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n13080) );
  INV_X1 U11472 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13107) );
  INV_X1 U11473 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13129) );
  INV_X1 U11474 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13119) );
  INV_X1 U11475 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9038) );
  OAI21_X1 U11476 ( .B1(n9390), .B2(n13119), .A(n9038), .ZN(n9040) );
  NAND2_X1 U11477 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n9039) );
  INV_X1 U11478 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9042) );
  AND3_X2 U11479 ( .A1(n9045), .A2(n9166), .A3(n9044), .ZN(n9047) );
  NOR2_X1 U11480 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), 
        .ZN(n9052) );
  NOR2_X1 U11481 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), 
        .ZN(n9051) );
  NOR2_X1 U11482 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), 
        .ZN(n9050) );
  NOR2_X1 U11483 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n9049) );
  INV_X1 U11484 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n13685) );
  XNOR2_X2 U11485 ( .A(n9056), .B(n13685), .ZN(n9062) );
  INV_X1 U11486 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n9058) );
  XNOR2_X2 U11487 ( .A(n9059), .B(n9058), .ZN(n13693) );
  OR2_X2 U11488 ( .A1(n9062), .A2(n13693), .ZN(n9124) );
  INV_X1 U11489 ( .A(n9124), .ZN(n9369) );
  NAND2_X1 U11490 ( .A1(n13331), .A2(n9369), .ZN(n9068) );
  INV_X1 U11491 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9065) );
  NAND2_X1 U11492 ( .A1(n9062), .A2(n9060), .ZN(n9125) );
  INV_X1 U11493 ( .A(n9062), .ZN(n9061) );
  NAND2_X2 U11494 ( .A1(n13693), .A2(n9061), .ZN(n9123) );
  INV_X2 U11495 ( .A(n9123), .ZN(n9750) );
  NAND2_X1 U11496 ( .A1(n9750), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n9064) );
  AND2_X4 U11497 ( .A1(n9062), .A2(n13693), .ZN(n9136) );
  NAND2_X1 U11498 ( .A1(n9136), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n9063) );
  OAI211_X1 U11499 ( .C1(n9065), .C2(n9534), .A(n9064), .B(n9063), .ZN(n9066)
         );
  INV_X1 U11500 ( .A(n9066), .ZN(n9067) );
  NAND2_X1 U11501 ( .A1(n9068), .A2(n9067), .ZN(n13184) );
  XNOR2_X2 U11502 ( .A(n9070), .B(n9069), .ZN(n9530) );
  NAND2_X1 U11503 ( .A1(n13702), .A2(n9746), .ZN(n9075) );
  OR2_X1 U11504 ( .A1(n6545), .A2(n13703), .ZN(n9074) );
  INV_X1 U11505 ( .A(n13557), .ZN(n13334) );
  XNOR2_X1 U11506 ( .A(n9390), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n13347) );
  NAND2_X1 U11507 ( .A1(n13347), .A2(n9369), .ZN(n9080) );
  INV_X1 U11508 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n10351) );
  NAND2_X1 U11509 ( .A1(n9136), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9077) );
  NAND2_X1 U11510 ( .A1(n9750), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9076) );
  OAI211_X1 U11511 ( .C1(n9534), .C2(n10351), .A(n9077), .B(n9076), .ZN(n9078)
         );
  INV_X1 U11512 ( .A(n9078), .ZN(n9079) );
  NAND2_X1 U11513 ( .A1(n9080), .A2(n9079), .ZN(n13185) );
  NAND2_X1 U11514 ( .A1(n11909), .A2(n9746), .ZN(n9082) );
  OR2_X1 U11515 ( .A1(n6544), .A2(n13706), .ZN(n9081) );
  INV_X1 U11516 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9083) );
  NAND2_X1 U11517 ( .A1(n9368), .A2(n9083), .ZN(n9084) );
  NAND2_X1 U11518 ( .A1(n9378), .A2(n9084), .ZN(n13151) );
  OR2_X1 U11519 ( .A1(n13151), .A2(n9124), .ZN(n9090) );
  INV_X1 U11520 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9087) );
  NAND2_X1 U11521 ( .A1(n9136), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9086) );
  NAND2_X1 U11522 ( .A1(n9750), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n9085) );
  OAI211_X1 U11523 ( .C1(n9534), .C2(n9087), .A(n9086), .B(n9085), .ZN(n9088)
         );
  INV_X1 U11524 ( .A(n9088), .ZN(n9089) );
  NAND2_X1 U11525 ( .A1(n9090), .A2(n9089), .ZN(n13188) );
  INV_X1 U11526 ( .A(n13188), .ZN(n9704) );
  XNOR2_X1 U11527 ( .A(n9092), .B(n9091), .ZN(n12064) );
  NAND2_X1 U11528 ( .A1(n12064), .A2(n9746), .ZN(n9094) );
  OR2_X1 U11529 ( .A1(n6545), .A2(n12067), .ZN(n9093) );
  NAND2_X2 U11530 ( .A1(n9094), .A2(n9093), .ZN(n13580) );
  INV_X1 U11531 ( .A(n13580), .ZN(n13392) );
  NAND2_X1 U11532 ( .A1(n11545), .A2(n9746), .ZN(n9096) );
  OR2_X1 U11533 ( .A1(n6545), .A2(n11550), .ZN(n9095) );
  INV_X1 U11534 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9097) );
  NAND2_X1 U11535 ( .A1(n9359), .A2(n9097), .ZN(n9098) );
  NAND2_X1 U11536 ( .A1(n9366), .A2(n9098), .ZN(n13415) );
  OR2_X1 U11537 ( .A1(n13415), .A2(n9124), .ZN(n9104) );
  INV_X1 U11538 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9101) );
  NAND2_X1 U11539 ( .A1(n9136), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n9100) );
  NAND2_X1 U11540 ( .A1(n9750), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n9099) );
  OAI211_X1 U11541 ( .C1(n9534), .C2(n9101), .A(n9100), .B(n9099), .ZN(n9102)
         );
  INV_X1 U11542 ( .A(n9102), .ZN(n9103) );
  NAND2_X1 U11543 ( .A1(n9104), .A2(n9103), .ZN(n13190) );
  INV_X1 U11544 ( .A(n13590), .ZN(n13418) );
  INV_X1 U11545 ( .A(n13190), .ZN(n9516) );
  INV_X1 U11546 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n11135) );
  INV_X1 U11547 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10078) );
  INV_X1 U11548 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n11130) );
  OR2_X1 U11549 ( .A1(n6544), .A2(n9109), .ZN(n9114) );
  NAND2_X1 U11550 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9110) );
  INV_X1 U11551 ( .A(n9130), .ZN(n9111) );
  NAND2_X1 U11552 ( .A1(n9112), .A2(n9111), .ZN(n10097) );
  OR2_X1 U11553 ( .A1(n9133), .A2(n9877), .ZN(n9113) );
  INV_X1 U11554 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10901) );
  OR2_X1 U11555 ( .A1(n9123), .A2(n10901), .ZN(n9119) );
  INV_X1 U11556 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10900) );
  OR2_X1 U11557 ( .A1(n9124), .A2(n10900), .ZN(n9118) );
  NAND2_X1 U11558 ( .A1(n9136), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n9117) );
  INV_X1 U11559 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9115) );
  OR2_X1 U11560 ( .A1(n9125), .A2(n9115), .ZN(n9116) );
  XNOR2_X1 U11561 ( .A(n9121), .B(n9120), .ZN(n13711) );
  MUX2_X1 U11562 ( .A(n9043), .B(n13711), .S(n6472), .Z(n11146) );
  INV_X1 U11563 ( .A(n9552), .ZN(n11156) );
  NAND2_X1 U11564 ( .A1(n11156), .A2(n11131), .ZN(n9122) );
  NAND2_X1 U11565 ( .A1(n10572), .A2(n9122), .ZN(n10561) );
  INV_X1 U11566 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10098) );
  OR2_X1 U11567 ( .A1(n9123), .A2(n10098), .ZN(n9129) );
  NAND2_X1 U11568 ( .A1(n9136), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n9128) );
  INV_X1 U11569 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11162) );
  OR2_X1 U11570 ( .A1(n9124), .A2(n11162), .ZN(n9127) );
  INV_X1 U11571 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10079) );
  OR2_X1 U11572 ( .A1(n9125), .A2(n10079), .ZN(n9126) );
  NAND4_X1 U11573 ( .A1(n9129), .A2(n9128), .A3(n9127), .A4(n9126), .ZN(n13207) );
  NOR2_X1 U11574 ( .A1(n9130), .A2(n9454), .ZN(n9131) );
  NAND2_X1 U11575 ( .A1(n10561), .A2(n10564), .ZN(n10560) );
  INV_X1 U11576 ( .A(n13207), .ZN(n9481) );
  NAND2_X1 U11577 ( .A1(n9481), .A2(n6909), .ZN(n9135) );
  NAND2_X1 U11578 ( .A1(n10560), .A2(n9135), .ZN(n10552) );
  NAND2_X1 U11579 ( .A1(n9750), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9141) );
  OR2_X1 U11580 ( .A1(n9422), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n9140) );
  INV_X1 U11581 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9137) );
  OR2_X1 U11582 ( .A1(n9753), .A2(n9137), .ZN(n9139) );
  INV_X1 U11583 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10081) );
  OR2_X1 U11584 ( .A1(n9125), .A2(n10081), .ZN(n9138) );
  NAND2_X1 U11585 ( .A1(n9132), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9143) );
  MUX2_X1 U11586 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9143), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n9144) );
  NAND2_X1 U11587 ( .A1(n9144), .A2(n9157), .ZN(n10100) );
  NAND2_X1 U11588 ( .A1(n10552), .A2(n10554), .ZN(n10551) );
  INV_X1 U11589 ( .A(n13206), .ZN(n11214) );
  NAND2_X1 U11590 ( .A1(n11214), .A2(n9145), .ZN(n9146) );
  NAND2_X1 U11591 ( .A1(n10551), .A2(n9146), .ZN(n10530) );
  NAND2_X1 U11592 ( .A1(n9749), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9155) );
  INV_X1 U11593 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11094) );
  OR2_X1 U11594 ( .A1(n9123), .A2(n11094), .ZN(n9154) );
  INV_X1 U11595 ( .A(n9171), .ZN(n9150) );
  INV_X1 U11596 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9148) );
  INV_X1 U11597 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9147) );
  NAND2_X1 U11598 ( .A1(n9148), .A2(n9147), .ZN(n9149) );
  NAND2_X1 U11599 ( .A1(n9150), .A2(n9149), .ZN(n11219) );
  OR2_X1 U11600 ( .A1(n9422), .A2(n11219), .ZN(n9153) );
  INV_X1 U11601 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9151) );
  OR2_X1 U11602 ( .A1(n9753), .A2(n9151), .ZN(n9152) );
  NOR2_X1 U11603 ( .A1(n9880), .A2(n9133), .ZN(n9162) );
  NAND2_X1 U11604 ( .A1(n9157), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9156) );
  MUX2_X1 U11605 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9156), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n9160) );
  INV_X1 U11606 ( .A(n9157), .ZN(n9159) );
  INV_X1 U11607 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n9158) );
  NAND2_X1 U11608 ( .A1(n9159), .A2(n9158), .ZN(n9165) );
  NAND2_X1 U11609 ( .A1(n9160), .A2(n9165), .ZN(n14868) );
  OAI22_X1 U11610 ( .A1(n6545), .A2(n9878), .B1(n10091), .B2(n14868), .ZN(
        n9161) );
  NAND2_X1 U11611 ( .A1(n10530), .A2(n10533), .ZN(n10529) );
  INV_X1 U11612 ( .A(n13205), .ZN(n9487) );
  NAND2_X1 U11613 ( .A1(n9487), .A2(n11223), .ZN(n9163) );
  NAND2_X1 U11614 ( .A1(n10529), .A2(n9163), .ZN(n11114) );
  OR2_X1 U11615 ( .A1(n9888), .A2(n9133), .ZN(n9170) );
  NAND2_X1 U11616 ( .A1(n9165), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9164) );
  MUX2_X1 U11617 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9164), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n9168) );
  INV_X1 U11618 ( .A(n9165), .ZN(n9167) );
  NAND2_X1 U11619 ( .A1(n9167), .A2(n9166), .ZN(n9189) );
  AOI22_X1 U11620 ( .A1(n9354), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9353), .B2(
        n10102), .ZN(n9169) );
  NAND2_X1 U11621 ( .A1(n9170), .A2(n9169), .ZN(n14964) );
  NAND2_X1 U11622 ( .A1(n9749), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9176) );
  INV_X1 U11623 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11125) );
  OR2_X1 U11624 ( .A1(n9123), .A2(n11125), .ZN(n9175) );
  OAI21_X1 U11625 ( .B1(n9171), .B2(P2_REG3_REG_5__SCAN_IN), .A(n9193), .ZN(
        n12347) );
  OR2_X1 U11626 ( .A1(n9422), .A2(n12347), .ZN(n9174) );
  INV_X1 U11627 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9172) );
  OR2_X1 U11628 ( .A1(n9753), .A2(n9172), .ZN(n9173) );
  NAND4_X1 U11629 ( .A1(n9176), .A2(n9175), .A3(n9174), .A4(n9173), .ZN(n13204) );
  NAND2_X1 U11630 ( .A1(n14964), .A2(n13204), .ZN(n9177) );
  INV_X1 U11631 ( .A(n14964), .ZN(n12350) );
  INV_X1 U11632 ( .A(n13204), .ZN(n9490) );
  NAND2_X1 U11633 ( .A1(n12350), .A2(n9490), .ZN(n9178) );
  OR2_X1 U11634 ( .A1(n9893), .A2(n9133), .ZN(n9181) );
  NAND2_X1 U11635 ( .A1(n9189), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9179) );
  XNOR2_X1 U11636 ( .A(n9179), .B(P2_IR_REG_6__SCAN_IN), .ZN(n14883) );
  AOI22_X1 U11637 ( .A1(n9354), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9353), .B2(
        n14883), .ZN(n9180) );
  NAND2_X1 U11638 ( .A1(n9750), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9188) );
  INV_X1 U11639 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9182) );
  OR2_X1 U11640 ( .A1(n9534), .A2(n9182), .ZN(n9187) );
  INV_X1 U11641 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9183) );
  XNOR2_X1 U11642 ( .A(n9193), .B(n9183), .ZN(n11292) );
  OR2_X1 U11643 ( .A1(n9422), .A2(n11292), .ZN(n9186) );
  INV_X1 U11644 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9184) );
  OR2_X1 U11645 ( .A1(n9753), .A2(n9184), .ZN(n9185) );
  NAND4_X1 U11646 ( .A1(n9188), .A2(n9187), .A3(n9186), .A4(n9185), .ZN(n13203) );
  INV_X1 U11647 ( .A(n13203), .ZN(n11191) );
  NAND2_X1 U11648 ( .A1(n10959), .A2(n11191), .ZN(n9492) );
  OR2_X1 U11649 ( .A1(n9901), .A2(n9133), .ZN(n9192) );
  OAI21_X1 U11650 ( .B1(n9189), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9190) );
  XNOR2_X1 U11651 ( .A(n9190), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10103) );
  AOI22_X1 U11652 ( .A1(n9354), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n9353), .B2(
        n10103), .ZN(n9191) );
  NAND2_X1 U11653 ( .A1(n9192), .A2(n9191), .ZN(n11038) );
  NAND2_X1 U11654 ( .A1(n9136), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n9199) );
  INV_X1 U11655 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11301) );
  OR2_X1 U11656 ( .A1(n9123), .A2(n11301), .ZN(n9198) );
  INV_X1 U11657 ( .A(n9193), .ZN(n9194) );
  AOI21_X1 U11658 ( .B1(n9194), .B2(P2_REG3_REG_6__SCAN_IN), .A(
        P2_REG3_REG_7__SCAN_IN), .ZN(n9195) );
  OR2_X1 U11659 ( .A1(n9195), .A2(n9210), .ZN(n11306) );
  OR2_X1 U11660 ( .A1(n9422), .A2(n11306), .ZN(n9197) );
  INV_X1 U11661 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10085) );
  OR2_X1 U11662 ( .A1(n9534), .A2(n10085), .ZN(n9196) );
  NAND4_X1 U11663 ( .A1(n9199), .A2(n9198), .A3(n9197), .A4(n9196), .ZN(n13202) );
  XNOR2_X1 U11664 ( .A(n11038), .B(n13202), .ZN(n11297) );
  INV_X1 U11665 ( .A(n11297), .ZN(n11303) );
  NAND2_X1 U11666 ( .A1(n11302), .A2(n11303), .ZN(n9201) );
  OR2_X1 U11667 ( .A1(n11038), .A2(n13202), .ZN(n9200) );
  NAND2_X1 U11668 ( .A1(n9201), .A2(n9200), .ZN(n11419) );
  OR2_X1 U11669 ( .A1(n9914), .A2(n9133), .ZN(n9208) );
  NAND2_X1 U11670 ( .A1(n9202), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9203) );
  MUX2_X1 U11671 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9203), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n9204) );
  INV_X1 U11672 ( .A(n9204), .ZN(n9206) );
  NOR2_X1 U11673 ( .A1(n9206), .A2(n9205), .ZN(n10105) );
  AOI22_X1 U11674 ( .A1(n9354), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n9353), .B2(
        n10105), .ZN(n9207) );
  NAND2_X1 U11675 ( .A1(n9208), .A2(n9207), .ZN(n11180) );
  NAND2_X1 U11676 ( .A1(n9750), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9215) );
  INV_X1 U11677 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9209) );
  OR2_X1 U11678 ( .A1(n9753), .A2(n9209), .ZN(n9214) );
  OR2_X1 U11679 ( .A1(n9210), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n9211) );
  NAND2_X1 U11680 ( .A1(n9223), .A2(n9211), .ZN(n11430) );
  OR2_X1 U11681 ( .A1(n9422), .A2(n11430), .ZN(n9213) );
  INV_X1 U11682 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10086) );
  OR2_X1 U11683 ( .A1(n9534), .A2(n10086), .ZN(n9212) );
  NAND4_X1 U11684 ( .A1(n9215), .A2(n9214), .A3(n9213), .A4(n9212), .ZN(n13201) );
  XNOR2_X1 U11685 ( .A(n11180), .B(n11256), .ZN(n11422) );
  INV_X1 U11686 ( .A(n11422), .ZN(n9216) );
  NOR2_X1 U11687 ( .A1(n11419), .A2(n9216), .ZN(n9217) );
  NAND2_X1 U11688 ( .A1(n11180), .A2(n13201), .ZN(n9218) );
  OR2_X1 U11689 ( .A1(n9927), .A2(n9133), .ZN(n9221) );
  OR2_X1 U11690 ( .A1(n9205), .A2(n9454), .ZN(n9219) );
  XNOR2_X1 U11691 ( .A(n9219), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10744) );
  AOI22_X1 U11692 ( .A1(n9354), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n9353), .B2(
        n10744), .ZN(n9220) );
  NAND2_X1 U11693 ( .A1(n9750), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n9229) );
  INV_X1 U11694 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10087) );
  OR2_X1 U11695 ( .A1(n9534), .A2(n10087), .ZN(n9228) );
  NAND2_X1 U11696 ( .A1(n9223), .A2(n9222), .ZN(n9224) );
  NAND2_X1 U11697 ( .A1(n9235), .A2(n9224), .ZN(n11507) );
  OR2_X1 U11698 ( .A1(n9422), .A2(n11507), .ZN(n9227) );
  INV_X1 U11699 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9225) );
  OR2_X1 U11700 ( .A1(n9753), .A2(n9225), .ZN(n9226) );
  NAND4_X1 U11701 ( .A1(n9229), .A2(n9228), .A3(n9227), .A4(n9226), .ZN(n13200) );
  NAND2_X1 U11702 ( .A1(n11363), .A2(n13200), .ZN(n9231) );
  OR2_X1 U11703 ( .A1(n11363), .A2(n13200), .ZN(n9230) );
  INV_X1 U11704 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9232) );
  AND2_X1 U11705 ( .A1(n9205), .A2(n9232), .ZN(n9258) );
  OR2_X1 U11706 ( .A1(n9258), .A2(n9454), .ZN(n9246) );
  XNOR2_X1 U11707 ( .A(n9246), .B(P2_IR_REG_10__SCAN_IN), .ZN(n14911) );
  AOI22_X1 U11708 ( .A1(n9354), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n9353), 
        .B2(n14911), .ZN(n9233) );
  NAND2_X2 U11709 ( .A1(n9234), .A2(n9233), .ZN(n11493) );
  NAND2_X1 U11710 ( .A1(n9750), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9241) );
  INV_X1 U11711 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10745) );
  OR2_X1 U11712 ( .A1(n9534), .A2(n10745), .ZN(n9240) );
  AND2_X1 U11713 ( .A1(n9235), .A2(n14905), .ZN(n9236) );
  OR2_X1 U11714 ( .A1(n9236), .A2(n9251), .ZN(n11349) );
  OR2_X1 U11715 ( .A1(n9422), .A2(n11349), .ZN(n9239) );
  INV_X1 U11716 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9237) );
  OR2_X1 U11717 ( .A1(n9753), .A2(n9237), .ZN(n9238) );
  NAND4_X1 U11718 ( .A1(n9241), .A2(n9240), .A3(n9239), .A4(n9238), .ZN(n13199) );
  NAND2_X1 U11719 ( .A1(n11493), .A2(n13199), .ZN(n9243) );
  OR2_X1 U11720 ( .A1(n11493), .A2(n13199), .ZN(n9242) );
  NAND2_X1 U11721 ( .A1(n11342), .A2(n9783), .ZN(n9244) );
  INV_X1 U11722 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n9245) );
  NAND2_X1 U11723 ( .A1(n9246), .A2(n9245), .ZN(n9247) );
  NAND2_X1 U11724 ( .A1(n9247), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9248) );
  XNOR2_X1 U11725 ( .A(n9248), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10849) );
  AOI22_X1 U11726 ( .A1(n9354), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n9353), 
        .B2(n10849), .ZN(n9249) );
  NAND2_X1 U11727 ( .A1(n9750), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n9256) );
  INV_X1 U11728 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9250) );
  OR2_X1 U11729 ( .A1(n9753), .A2(n9250), .ZN(n9255) );
  NOR2_X1 U11730 ( .A1(n9251), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n9252) );
  OR2_X1 U11731 ( .A1(n9266), .A2(n9252), .ZN(n13522) );
  OR2_X1 U11732 ( .A1(n9422), .A2(n13522), .ZN(n9254) );
  INV_X1 U11733 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10746) );
  OR2_X1 U11734 ( .A1(n9534), .A2(n10746), .ZN(n9253) );
  NAND4_X1 U11735 ( .A1(n9256), .A2(n9255), .A3(n9254), .A4(n9253), .ZN(n13198) );
  NAND2_X1 U11736 ( .A1(n10180), .A2(n9746), .ZN(n9265) );
  NOR2_X1 U11737 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), 
        .ZN(n9257) );
  AND2_X1 U11738 ( .A1(n9258), .A2(n9257), .ZN(n9261) );
  NOR2_X1 U11739 ( .A1(n9261), .A2(n9454), .ZN(n9259) );
  MUX2_X1 U11740 ( .A(n9454), .B(n9259), .S(P2_IR_REG_12__SCAN_IN), .Z(n9263)
         );
  INV_X1 U11741 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n9260) );
  NAND2_X1 U11742 ( .A1(n9261), .A2(n9260), .ZN(n9274) );
  INV_X1 U11743 ( .A(n9274), .ZN(n9262) );
  NOR2_X1 U11744 ( .A1(n9263), .A2(n9262), .ZN(n11102) );
  AOI22_X1 U11745 ( .A1(n9354), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n9353), 
        .B2(n11102), .ZN(n9264) );
  NAND2_X1 U11746 ( .A1(n9136), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9271) );
  INV_X1 U11747 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10850) );
  OR2_X1 U11748 ( .A1(n9534), .A2(n10850), .ZN(n9270) );
  INV_X1 U11749 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11584) );
  OR2_X1 U11750 ( .A1(n9123), .A2(n11584), .ZN(n9269) );
  OR2_X1 U11751 ( .A1(n9266), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9267) );
  NAND2_X1 U11752 ( .A1(n9278), .A2(n9267), .ZN(n11583) );
  OR2_X1 U11753 ( .A1(n9124), .A2(n11583), .ZN(n9268) );
  NAND4_X1 U11754 ( .A1(n9271), .A2(n9270), .A3(n9269), .A4(n9268), .ZN(n13197) );
  XNOR2_X1 U11755 ( .A(n11741), .B(n13197), .ZN(n11578) );
  NAND2_X1 U11756 ( .A1(n10399), .A2(n9746), .ZN(n9277) );
  NAND2_X1 U11757 ( .A1(n9274), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9273) );
  MUX2_X1 U11758 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9273), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n9275) );
  AND2_X1 U11759 ( .A1(n9275), .A2(n9297), .ZN(n11482) );
  AOI22_X1 U11760 ( .A1(n9354), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n9353), 
        .B2(n11482), .ZN(n9276) );
  NAND2_X1 U11761 ( .A1(n9749), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9284) );
  INV_X1 U11762 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11669) );
  OR2_X1 U11763 ( .A1(n9123), .A2(n11669), .ZN(n9283) );
  NAND2_X1 U11764 ( .A1(n9278), .A2(n14820), .ZN(n9279) );
  NAND2_X1 U11765 ( .A1(n9290), .A2(n9279), .ZN(n14833) );
  OR2_X1 U11766 ( .A1(n9422), .A2(n14833), .ZN(n9282) );
  INV_X1 U11767 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9280) );
  OR2_X1 U11768 ( .A1(n9753), .A2(n9280), .ZN(n9281) );
  NAND4_X1 U11769 ( .A1(n9284), .A2(n9283), .A3(n9282), .A4(n9281), .ZN(n11566) );
  NAND2_X1 U11770 ( .A1(n14830), .A2(n11566), .ZN(n9285) );
  OR2_X1 U11771 ( .A1(n14830), .A2(n11566), .ZN(n9286) );
  NAND2_X1 U11772 ( .A1(n10730), .A2(n9746), .ZN(n9289) );
  NAND2_X1 U11773 ( .A1(n9297), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9287) );
  XNOR2_X1 U11774 ( .A(n9287), .B(P2_IR_REG_14__SCAN_IN), .ZN(n13238) );
  AOI22_X1 U11775 ( .A1(n9354), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n9353), 
        .B2(n13238), .ZN(n9288) );
  NAND2_X1 U11776 ( .A1(n9749), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n9295) );
  INV_X1 U11777 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n13224) );
  OR2_X1 U11778 ( .A1(n9123), .A2(n13224), .ZN(n9294) );
  NAND2_X1 U11779 ( .A1(n9290), .A2(n11567), .ZN(n9291) );
  NAND2_X1 U11780 ( .A1(n9305), .A2(n9291), .ZN(n11565) );
  OR2_X1 U11781 ( .A1(n9124), .A2(n11565), .ZN(n9293) );
  INV_X1 U11782 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n13675) );
  OR2_X1 U11783 ( .A1(n9753), .A2(n13675), .ZN(n9292) );
  NAND4_X1 U11784 ( .A1(n9295), .A2(n9294), .A3(n9293), .A4(n9292), .ZN(n13196) );
  NOR2_X1 U11785 ( .A1(n13510), .A2(n13196), .ZN(n9776) );
  AND2_X1 U11786 ( .A1(n13510), .A2(n13196), .ZN(n9777) );
  INV_X1 U11787 ( .A(n9777), .ZN(n9296) );
  NAND2_X1 U11788 ( .A1(n10758), .A2(n9746), .ZN(n9302) );
  OAI21_X1 U11789 ( .B1(n9297), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9299) );
  INV_X1 U11790 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n9298) );
  NAND2_X1 U11791 ( .A1(n9299), .A2(n9298), .ZN(n9313) );
  OR2_X1 U11792 ( .A1(n9299), .A2(n9298), .ZN(n9300) );
  AND2_X1 U11793 ( .A1(n9313), .A2(n9300), .ZN(n13228) );
  AOI22_X1 U11794 ( .A1(n9354), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n9353), 
        .B2(n13228), .ZN(n9301) );
  INV_X1 U11795 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14920) );
  OR2_X1 U11796 ( .A1(n9534), .A2(n14920), .ZN(n9310) );
  INV_X1 U11797 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n13495) );
  OR2_X1 U11798 ( .A1(n9123), .A2(n13495), .ZN(n9309) );
  INV_X1 U11799 ( .A(n9303), .ZN(n9318) );
  NAND2_X1 U11800 ( .A1(n9305), .A2(n9304), .ZN(n9306) );
  NAND2_X1 U11801 ( .A1(n9318), .A2(n9306), .ZN(n13494) );
  OR2_X1 U11802 ( .A1(n9124), .A2(n13494), .ZN(n9308) );
  INV_X1 U11803 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n10223) );
  OR2_X1 U11804 ( .A1(n9753), .A2(n10223), .ZN(n9307) );
  NAND4_X1 U11805 ( .A1(n9310), .A2(n9309), .A3(n9308), .A4(n9307), .ZN(n13195) );
  XNOR2_X1 U11806 ( .A(n13672), .B(n13195), .ZN(n13486) );
  OR2_X1 U11807 ( .A1(n13672), .A2(n13195), .ZN(n9311) );
  NAND2_X1 U11808 ( .A1(n9312), .A2(n9311), .ZN(n13473) );
  NAND2_X1 U11809 ( .A1(n10602), .A2(n9746), .ZN(n9316) );
  NAND2_X1 U11810 ( .A1(n9313), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9314) );
  XNOR2_X1 U11811 ( .A(n9314), .B(P2_IR_REG_16__SCAN_IN), .ZN(n14938) );
  AOI22_X1 U11812 ( .A1(n14938), .A2(n9353), .B1(n9354), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n9315) );
  NAND2_X1 U11813 ( .A1(n9749), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n9323) );
  INV_X1 U11814 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9317) );
  OR2_X1 U11815 ( .A1(n9123), .A2(n9317), .ZN(n9322) );
  INV_X1 U11816 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n14931) );
  NAND2_X1 U11817 ( .A1(n9318), .A2(n14931), .ZN(n9319) );
  NAND2_X1 U11818 ( .A1(n9334), .A2(n9319), .ZN(n13471) );
  OR2_X1 U11819 ( .A1(n9422), .A2(n13471), .ZN(n9321) );
  INV_X1 U11820 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n13667) );
  OR2_X1 U11821 ( .A1(n9753), .A2(n13667), .ZN(n9320) );
  NAND4_X1 U11822 ( .A1(n9323), .A2(n9322), .A3(n9321), .A4(n9320), .ZN(n13194) );
  NAND2_X1 U11823 ( .A1(n13477), .A2(n13194), .ZN(n9326) );
  OR2_X1 U11824 ( .A1(n13477), .A2(n13194), .ZN(n9324) );
  NAND2_X1 U11825 ( .A1(n10756), .A2(n9746), .ZN(n9332) );
  NOR2_X1 U11826 ( .A1(n9327), .A2(n9454), .ZN(n9328) );
  MUX2_X1 U11827 ( .A(n9454), .B(n9328), .S(P2_IR_REG_17__SCAN_IN), .Z(n9330)
         );
  INV_X1 U11828 ( .A(n9339), .ZN(n9329) );
  NOR2_X1 U11829 ( .A1(n9330), .A2(n9329), .ZN(n13255) );
  AOI22_X1 U11830 ( .A1(n9354), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n9353), 
        .B2(n13255), .ZN(n9331) );
  INV_X1 U11831 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13609) );
  NAND2_X1 U11832 ( .A1(n9750), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n9333) );
  OAI21_X1 U11833 ( .B1(n13609), .B2(n9534), .A(n9333), .ZN(n9338) );
  NAND2_X1 U11834 ( .A1(n9334), .A2(n12070), .ZN(n9335) );
  NAND2_X1 U11835 ( .A1(n9345), .A2(n9335), .ZN(n13462) );
  NAND2_X1 U11836 ( .A1(n9136), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n9336) );
  OAI21_X1 U11837 ( .B1(n13462), .B2(n9124), .A(n9336), .ZN(n9337) );
  INV_X1 U11838 ( .A(n13193), .ZN(n9667) );
  XNOR2_X1 U11839 ( .A(n12073), .B(n9667), .ZN(n13451) );
  NAND2_X1 U11840 ( .A1(n11067), .A2(n9746), .ZN(n9344) );
  INV_X1 U11841 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n9340) );
  NAND2_X1 U11842 ( .A1(n9339), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9341) );
  MUX2_X1 U11843 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9341), .S(
        P2_IR_REG_18__SCAN_IN), .Z(n9342) );
  AND2_X1 U11844 ( .A1(n9430), .A2(n9342), .ZN(n13265) );
  AOI22_X1 U11845 ( .A1(n9354), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n9353), 
        .B2(n13265), .ZN(n9343) );
  INV_X1 U11846 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9349) );
  INV_X1 U11847 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10324) );
  NAND2_X1 U11848 ( .A1(n9345), .A2(n10324), .ZN(n9346) );
  NAND2_X1 U11849 ( .A1(n9357), .A2(n9346), .ZN(n13442) );
  OR2_X1 U11850 ( .A1(n13442), .A2(n9124), .ZN(n9348) );
  AOI22_X1 U11851 ( .A1(n9749), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n9750), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n9347) );
  OAI211_X1 U11852 ( .C1(n9753), .C2(n9349), .A(n9348), .B(n9347), .ZN(n13192)
         );
  XNOR2_X1 U11853 ( .A(n13601), .B(n13192), .ZN(n9787) );
  NAND2_X1 U11854 ( .A1(n11246), .A2(n9746), .ZN(n9356) );
  AOI22_X1 U11855 ( .A1(n9354), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9799), 
        .B2(n9353), .ZN(n9355) );
  INV_X1 U11856 ( .A(n13596), .ZN(n13434) );
  NAND2_X1 U11857 ( .A1(n9357), .A2(n13080), .ZN(n9358) );
  NAND2_X1 U11858 ( .A1(n9359), .A2(n9358), .ZN(n13431) );
  AOI22_X1 U11859 ( .A1(n9749), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n9750), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n9361) );
  NAND2_X1 U11860 ( .A1(n9136), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n9360) );
  OAI211_X1 U11861 ( .C1(n13431), .C2(n9422), .A(n9361), .B(n9360), .ZN(n13191) );
  INV_X1 U11862 ( .A(n13191), .ZN(n13141) );
  NAND2_X1 U11863 ( .A1(n13424), .A2(n7483), .ZN(n9363) );
  NAND2_X1 U11864 ( .A1(n11594), .A2(n9746), .ZN(n9365) );
  OR2_X1 U11865 ( .A1(n6544), .A2(n12417), .ZN(n9364) );
  NAND2_X1 U11866 ( .A1(n9366), .A2(n13107), .ZN(n9367) );
  AND2_X1 U11867 ( .A1(n9368), .A2(n9367), .ZN(n13405) );
  NAND2_X1 U11868 ( .A1(n13405), .A2(n9369), .ZN(n9374) );
  INV_X1 U11869 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n13587) );
  NAND2_X1 U11870 ( .A1(n9750), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n9371) );
  NAND2_X1 U11871 ( .A1(n9136), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n9370) );
  OAI211_X1 U11872 ( .C1(n9534), .C2(n13587), .A(n9371), .B(n9370), .ZN(n9372)
         );
  INV_X1 U11873 ( .A(n9372), .ZN(n9373) );
  NAND2_X1 U11874 ( .A1(n9374), .A2(n9373), .ZN(n13189) );
  INV_X1 U11875 ( .A(n13189), .ZN(n13137) );
  XNOR2_X1 U11876 ( .A(n13404), .B(n13137), .ZN(n13399) );
  XNOR2_X1 U11877 ( .A(n13580), .B(n9704), .ZN(n13385) );
  NAND2_X1 U11878 ( .A1(n13386), .A2(n13385), .ZN(n13384) );
  OAI21_X1 U11879 ( .B1(n9704), .B2(n13392), .A(n13384), .ZN(n13372) );
  NAND2_X1 U11880 ( .A1(n11855), .A2(n9746), .ZN(n9376) );
  OR2_X1 U11881 ( .A1(n6545), .A2(n11858), .ZN(n9375) );
  NAND2_X2 U11882 ( .A1(n9376), .A2(n9375), .ZN(n13375) );
  INV_X1 U11883 ( .A(n13375), .ZN(n13654) );
  INV_X1 U11884 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9377) );
  NAND2_X1 U11885 ( .A1(n9378), .A2(n9377), .ZN(n9379) );
  NAND2_X1 U11886 ( .A1(n9388), .A2(n9379), .ZN(n13074) );
  OR2_X1 U11887 ( .A1(n13074), .A2(n9422), .ZN(n9384) );
  INV_X1 U11888 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n13652) );
  NAND2_X1 U11889 ( .A1(n9749), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n9381) );
  NAND2_X1 U11890 ( .A1(n9750), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n9380) );
  OAI211_X1 U11891 ( .C1(n13652), .C2(n9753), .A(n9381), .B(n9380), .ZN(n9382)
         );
  INV_X1 U11892 ( .A(n9382), .ZN(n9383) );
  NAND2_X1 U11893 ( .A1(n9384), .A2(n9383), .ZN(n13187) );
  INV_X1 U11894 ( .A(n13187), .ZN(n13127) );
  NOR2_X1 U11895 ( .A1(n13654), .A2(n13127), .ZN(n9385) );
  NAND2_X1 U11896 ( .A1(n11859), .A2(n9746), .ZN(n9387) );
  OR2_X1 U11897 ( .A1(n6544), .A2(n11862), .ZN(n9386) );
  NAND2_X1 U11898 ( .A1(n9388), .A2(n13129), .ZN(n9389) );
  NAND2_X1 U11899 ( .A1(n9390), .A2(n9389), .ZN(n13361) );
  OR2_X1 U11900 ( .A1(n13361), .A2(n9124), .ZN(n9396) );
  INV_X1 U11901 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9393) );
  NAND2_X1 U11902 ( .A1(n9136), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9392) );
  NAND2_X1 U11903 ( .A1(n9750), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9391) );
  OAI211_X1 U11904 ( .C1(n9534), .C2(n9393), .A(n9392), .B(n9391), .ZN(n9394)
         );
  INV_X1 U11905 ( .A(n9394), .ZN(n9395) );
  NAND2_X1 U11906 ( .A1(n9396), .A2(n9395), .ZN(n13186) );
  INV_X1 U11907 ( .A(n13185), .ZN(n13128) );
  XNOR2_X1 U11908 ( .A(n13562), .B(n13128), .ZN(n13344) );
  NAND2_X1 U11909 ( .A1(n13699), .A2(n9746), .ZN(n9399) );
  OR2_X1 U11910 ( .A1(n6544), .A2(n13700), .ZN(n9398) );
  INV_X1 U11911 ( .A(n9401), .ZN(n9400) );
  NAND2_X1 U11912 ( .A1(n9400), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n9411) );
  INV_X1 U11913 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13066) );
  NAND2_X1 U11914 ( .A1(n9401), .A2(n13066), .ZN(n9402) );
  NAND2_X1 U11915 ( .A1(n9411), .A2(n9402), .ZN(n13318) );
  OR2_X1 U11916 ( .A1(n13318), .A2(n9124), .ZN(n9407) );
  INV_X1 U11917 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n13553) );
  NAND2_X1 U11918 ( .A1(n9750), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9404) );
  NAND2_X1 U11919 ( .A1(n9136), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9403) );
  OAI211_X1 U11920 ( .C1(n9534), .C2(n13553), .A(n9404), .B(n9403), .ZN(n9405)
         );
  INV_X1 U11921 ( .A(n9405), .ZN(n9406) );
  NAND2_X1 U11922 ( .A1(n13695), .A2(n9746), .ZN(n9409) );
  OR2_X1 U11923 ( .A1(n6545), .A2(n13698), .ZN(n9408) );
  INV_X1 U11924 ( .A(n9411), .ZN(n9410) );
  NAND2_X1 U11925 ( .A1(n9410), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n9543) );
  INV_X1 U11926 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n13099) );
  NAND2_X1 U11927 ( .A1(n9411), .A2(n13099), .ZN(n9412) );
  NAND2_X1 U11928 ( .A1(n9543), .A2(n9412), .ZN(n13297) );
  INV_X1 U11929 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13296) );
  NAND2_X1 U11930 ( .A1(n9749), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n9414) );
  NAND2_X1 U11931 ( .A1(n9136), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9413) );
  OAI211_X1 U11932 ( .C1(n9123), .C2(n13296), .A(n9414), .B(n9413), .ZN(n9415)
         );
  INV_X1 U11933 ( .A(n9415), .ZN(n9416) );
  INV_X1 U11934 ( .A(n13182), .ZN(n9418) );
  NAND2_X1 U11935 ( .A1(n13548), .A2(n9418), .ZN(n9419) );
  AOI22_X1 U11936 ( .A1(n13293), .A2(n13292), .B1(n13548), .B2(n13182), .ZN(
        n9429) );
  NAND2_X1 U11937 ( .A1(n11928), .A2(n9746), .ZN(n9421) );
  OR2_X1 U11938 ( .A1(n6544), .A2(n13691), .ZN(n9420) );
  OR2_X1 U11939 ( .A1(n9543), .A2(n9422), .ZN(n9428) );
  INV_X1 U11940 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9425) );
  NAND2_X1 U11941 ( .A1(n9750), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9424) );
  NAND2_X1 U11942 ( .A1(n9136), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9423) );
  OAI211_X1 U11943 ( .C1(n9425), .C2(n9534), .A(n9424), .B(n9423), .ZN(n9426)
         );
  INV_X1 U11944 ( .A(n9426), .ZN(n9427) );
  NAND2_X1 U11945 ( .A1(n9428), .A2(n9427), .ZN(n13181) );
  XNOR2_X1 U11946 ( .A(n9429), .B(n9794), .ZN(n13545) );
  INV_X1 U11947 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n9431) );
  INV_X1 U11948 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9432) );
  NAND2_X1 U11949 ( .A1(n7246), .A2(n9434), .ZN(n9436) );
  NAND2_X1 U11950 ( .A1(n9436), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9435) );
  MUX2_X1 U11951 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9435), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n9439) );
  INV_X1 U11952 ( .A(n9436), .ZN(n9438) );
  NAND2_X1 U11953 ( .A1(n9438), .A2(n9437), .ZN(n9440) );
  NAND2_X1 U11954 ( .A1(n9439), .A2(n9440), .ZN(n13710) );
  NAND2_X1 U11955 ( .A1(n9440), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9441) );
  MUX2_X1 U11956 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9441), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n9443) );
  NAND2_X1 U11957 ( .A1(n9443), .A2(n9442), .ZN(n13704) );
  NAND2_X1 U11958 ( .A1(n9453), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9445) );
  INV_X1 U11959 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9444) );
  XNOR2_X1 U11960 ( .A(n9445), .B(n9444), .ZN(n10090) );
  NAND2_X1 U11961 ( .A1(n9454), .A2(n9431), .ZN(n9447) );
  NAND2_X1 U11962 ( .A1(n9450), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9451) );
  MUX2_X1 U11963 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9451), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n9452) );
  NAND2_X2 U11964 ( .A1(n9453), .A2(n9452), .ZN(n12065) );
  XNOR2_X1 U11965 ( .A(n9457), .B(n9456), .ZN(n9473) );
  NAND2_X1 U11966 ( .A1(n10896), .A2(n6840), .ZN(n10540) );
  INV_X1 U11967 ( .A(n10540), .ZN(n9458) );
  NAND2_X1 U11968 ( .A1(n11864), .A2(n13704), .ZN(n9462) );
  XNOR2_X1 U11969 ( .A(n11864), .B(P2_B_REG_SCAN_IN), .ZN(n9459) );
  AND2_X1 U11970 ( .A1(n13710), .A2(n9459), .ZN(n9460) );
  INV_X1 U11971 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14952) );
  NAND2_X1 U11972 ( .A1(n14947), .A2(n14952), .ZN(n9461) );
  INV_X1 U11973 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14958) );
  AOI22_X1 U11974 ( .A1(n14947), .A2(n14958), .B1(n13704), .B2(n13710), .ZN(
        n10538) );
  NOR4_X1 U11975 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n9466) );
  NOR4_X1 U11976 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n9465) );
  NOR4_X1 U11977 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9464) );
  NOR4_X1 U11978 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n9463) );
  NAND4_X1 U11979 ( .A1(n9466), .A2(n9465), .A3(n9464), .A4(n9463), .ZN(n9472)
         );
  NOR2_X1 U11980 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .ZN(
        n9470) );
  NOR4_X1 U11981 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n9469) );
  NOR4_X1 U11982 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n9468) );
  NOR4_X1 U11983 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n9467) );
  NAND4_X1 U11984 ( .A1(n9470), .A2(n9469), .A3(n9468), .A4(n9467), .ZN(n9471)
         );
  OAI21_X1 U11985 ( .B1(n9472), .B2(n9471), .A(n14947), .ZN(n10541) );
  NAND2_X1 U11986 ( .A1(n10538), .A2(n10541), .ZN(n10401) );
  INV_X1 U11987 ( .A(n10401), .ZN(n9474) );
  NAND2_X1 U11988 ( .A1(n11552), .A2(n13276), .ZN(n9842) );
  NAND2_X1 U11989 ( .A1(n10411), .A2(n9842), .ZN(n10539) );
  AND3_X1 U11990 ( .A1(n14953), .A2(n9474), .A3(n10539), .ZN(n9475) );
  NAND2_X1 U11991 ( .A1(n14954), .A2(n9475), .ZN(n9476) );
  NOR2_X2 U11992 ( .A1(n12419), .A2(n9798), .ZN(n9826) );
  XNOR2_X1 U11993 ( .A(n9826), .B(n12065), .ZN(n9477) );
  NAND2_X1 U11994 ( .A1(n14986), .A2(n6669), .ZN(n9479) );
  INV_X1 U11995 ( .A(n9559), .ZN(n11140) );
  NAND2_X1 U11996 ( .A1(n11140), .A2(n10897), .ZN(n10576) );
  INV_X1 U11997 ( .A(n10564), .ZN(n9480) );
  NAND2_X1 U11998 ( .A1(n10565), .A2(n9480), .ZN(n9483) );
  NAND2_X1 U11999 ( .A1(n9481), .A2(n11166), .ZN(n9482) );
  NAND2_X1 U12000 ( .A1(n10555), .A2(n9778), .ZN(n9485) );
  NAND2_X1 U12001 ( .A1(n11214), .A2(n14818), .ZN(n9484) );
  INV_X1 U12002 ( .A(n10533), .ZN(n9486) );
  NAND2_X1 U12003 ( .A1(n10534), .A2(n9486), .ZN(n9489) );
  NAND2_X1 U12004 ( .A1(n9487), .A2(n10927), .ZN(n9488) );
  NAND2_X1 U12005 ( .A1(n9489), .A2(n9488), .ZN(n11121) );
  NAND2_X1 U12006 ( .A1(n12350), .A2(n13204), .ZN(n9491) );
  INV_X1 U12007 ( .A(n13202), .ZN(n11170) );
  OR2_X1 U12008 ( .A1(n11038), .A2(n11170), .ZN(n9493) );
  OR2_X1 U12009 ( .A1(n11180), .A2(n11256), .ZN(n9494) );
  INV_X1 U12010 ( .A(n13200), .ZN(n9495) );
  OR2_X1 U12011 ( .A1(n11363), .A2(n9495), .ZN(n9496) );
  NAND2_X1 U12012 ( .A1(n11359), .A2(n9496), .ZN(n11345) );
  NAND2_X1 U12013 ( .A1(n11345), .A2(n11344), .ZN(n11343) );
  INV_X1 U12014 ( .A(n13199), .ZN(n9497) );
  OR2_X1 U12015 ( .A1(n11493), .A2(n9497), .ZN(n9498) );
  INV_X1 U12016 ( .A(n13198), .ZN(n11276) );
  NAND2_X1 U12017 ( .A1(n13526), .A2(n11276), .ZN(n9501) );
  OR2_X1 U12018 ( .A1(n13526), .A2(n11276), .ZN(n9499) );
  INV_X1 U12019 ( .A(n11596), .ZN(n11604) );
  INV_X1 U12020 ( .A(n13197), .ZN(n9502) );
  INV_X1 U12021 ( .A(n11566), .ZN(n9639) );
  NAND2_X1 U12022 ( .A1(n14830), .A2(n9639), .ZN(n9503) );
  OR2_X1 U12023 ( .A1(n14830), .A2(n9639), .ZN(n9504) );
  INV_X1 U12024 ( .A(n13196), .ZN(n9505) );
  NOR2_X1 U12025 ( .A1(n13510), .A2(n9505), .ZN(n9506) );
  INV_X1 U12026 ( .A(n13195), .ZN(n9507) );
  INV_X1 U12027 ( .A(n13194), .ZN(n9508) );
  NAND2_X1 U12028 ( .A1(n13477), .A2(n9508), .ZN(n9509) );
  AND2_X1 U12029 ( .A1(n12073), .A2(n9667), .ZN(n9512) );
  OR2_X1 U12030 ( .A1(n12073), .A2(n9667), .ZN(n9511) );
  NOR2_X1 U12031 ( .A1(n13601), .A2(n9350), .ZN(n9513) );
  XNOR2_X1 U12032 ( .A(n13596), .B(n13191), .ZN(n13426) );
  NAND2_X1 U12033 ( .A1(n13596), .A2(n13141), .ZN(n9514) );
  XNOR2_X1 U12034 ( .A(n13590), .B(n9516), .ZN(n9790) );
  NAND2_X1 U12035 ( .A1(n13411), .A2(n13420), .ZN(n9518) );
  NAND2_X1 U12036 ( .A1(n13590), .A2(n9516), .ZN(n9517) );
  AND2_X1 U12037 ( .A1(n13404), .A2(n13137), .ZN(n9519) );
  OR2_X1 U12038 ( .A1(n13404), .A2(n13137), .ZN(n9520) );
  NOR2_X1 U12039 ( .A1(n13375), .A2(n13127), .ZN(n9521) );
  NAND2_X1 U12040 ( .A1(n13375), .A2(n13127), .ZN(n9522) );
  INV_X1 U12041 ( .A(n13186), .ZN(n13117) );
  NAND2_X1 U12042 ( .A1(n13567), .A2(n13117), .ZN(n9523) );
  NAND2_X1 U12043 ( .A1(n13325), .A2(n9775), .ZN(n9524) );
  NAND2_X1 U12044 ( .A1(n13557), .A2(n13118), .ZN(n9774) );
  INV_X1 U12045 ( .A(n13292), .ZN(n13300) );
  NAND2_X1 U12046 ( .A1(n13317), .A2(n9525), .ZN(n13301) );
  NAND2_X1 U12047 ( .A1(n13302), .A2(n9526), .ZN(n9528) );
  OR2_X1 U12048 ( .A1(n12065), .A2(n13276), .ZN(n9529) );
  INV_X1 U12049 ( .A(n9530), .ZN(n9531) );
  NAND2_X1 U12050 ( .A1(n10411), .A2(n9531), .ZN(n13135) );
  NAND2_X1 U12051 ( .A1(n13182), .A2(n13172), .ZN(n9538) );
  INV_X1 U12052 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13539) );
  NAND2_X1 U12053 ( .A1(n9750), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9533) );
  NAND2_X1 U12054 ( .A1(n9136), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9532) );
  OAI211_X1 U12055 ( .C1(n9534), .C2(n13539), .A(n9533), .B(n9532), .ZN(n13180) );
  NAND2_X1 U12056 ( .A1(n10411), .A2(n9530), .ZN(n13136) );
  INV_X1 U12057 ( .A(P2_B_REG_SCAN_IN), .ZN(n9535) );
  NOR2_X1 U12058 ( .A1(n13701), .A2(n9535), .ZN(n9536) );
  NOR2_X1 U12059 ( .A1(n13136), .A2(n9536), .ZN(n13284) );
  NAND2_X1 U12060 ( .A1(n13180), .A2(n13284), .ZN(n9537) );
  INV_X1 U12061 ( .A(n11741), .ZN(n11738) );
  INV_X1 U12062 ( .A(n13526), .ZN(n11606) );
  NAND2_X1 U12063 ( .A1(n10553), .A2(n11223), .ZN(n11115) );
  OR2_X1 U12064 ( .A1(n11115), .A2(n14964), .ZN(n11289) );
  NOR2_X2 U12065 ( .A1(n11289), .A2(n10959), .ZN(n11305) );
  INV_X1 U12066 ( .A(n11038), .ZN(n14980) );
  AND2_X2 U12067 ( .A1(n11305), .A2(n14980), .ZN(n11429) );
  INV_X1 U12068 ( .A(n11180), .ZN(n14990) );
  NAND2_X1 U12069 ( .A1(n11429), .A2(n14990), .ZN(n11356) );
  OR2_X2 U12070 ( .A1(n11356), .A2(n11363), .ZN(n11357) );
  INV_X1 U12071 ( .A(n13672), .ZN(n9541) );
  INV_X1 U12072 ( .A(n13567), .ZN(n13359) );
  NOR2_X2 U12073 ( .A1(n13358), .A2(n13562), .ZN(n13328) );
  AOI211_X1 U12074 ( .C1(n13542), .C2(n13294), .A(n13490), .B(n13288), .ZN(
        n13541) );
  INV_X1 U12075 ( .A(n13542), .ZN(n9546) );
  AND2_X1 U12076 ( .A1(n10896), .A2(n9798), .ZN(n10403) );
  INV_X1 U12077 ( .A(n9543), .ZN(n9544) );
  INV_X1 U12078 ( .A(n13521), .ZN(n13511) );
  AOI22_X1 U12079 ( .A1(n9544), .A2(n13511), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n13517), .ZN(n9545) );
  OAI21_X1 U12080 ( .B1(n9546), .B2(n13461), .A(n9545), .ZN(n9547) );
  NAND2_X1 U12081 ( .A1(n9641), .A2(n10582), .ZN(n9551) );
  NAND2_X1 U12082 ( .A1(n9552), .A2(n9611), .ZN(n9550) );
  NAND2_X1 U12083 ( .A1(n9552), .A2(n9641), .ZN(n9554) );
  NAND2_X1 U12084 ( .A1(n9819), .A2(n10582), .ZN(n9553) );
  NAND2_X1 U12085 ( .A1(n9554), .A2(n9553), .ZN(n9565) );
  NAND2_X1 U12086 ( .A1(n12065), .A2(n9799), .ZN(n9555) );
  NAND2_X1 U12087 ( .A1(n9826), .A2(n9555), .ZN(n9560) );
  NAND2_X1 U12088 ( .A1(n9560), .A2(n11146), .ZN(n9557) );
  NAND2_X1 U12089 ( .A1(n10897), .A2(n9641), .ZN(n9556) );
  OAI21_X1 U12090 ( .B1(n9559), .B2(n9557), .A(n9556), .ZN(n9558) );
  INV_X1 U12091 ( .A(n9558), .ZN(n9562) );
  OAI211_X1 U12092 ( .C1(n9560), .C2(n11146), .A(n9559), .B(n9819), .ZN(n9561)
         );
  NAND2_X1 U12093 ( .A1(n9562), .A2(n9561), .ZN(n9563) );
  NAND2_X1 U12094 ( .A1(n9564), .A2(n9563), .ZN(n9569) );
  INV_X1 U12095 ( .A(n9565), .ZN(n9567) );
  NAND2_X1 U12096 ( .A1(n9567), .A2(n9566), .ZN(n9568) );
  NAND2_X1 U12097 ( .A1(n13207), .A2(n9819), .ZN(n9571) );
  NAND2_X1 U12098 ( .A1(n9761), .A2(n11166), .ZN(n9570) );
  NAND2_X1 U12099 ( .A1(n9571), .A2(n9570), .ZN(n9573) );
  AOI22_X1 U12100 ( .A1(n13207), .A2(n9641), .B1(n9819), .B2(n11166), .ZN(
        n9572) );
  NAND2_X1 U12101 ( .A1(n13206), .A2(n9761), .ZN(n9575) );
  INV_X2 U12102 ( .A(n9641), .ZN(n9769) );
  NAND2_X1 U12103 ( .A1(n9769), .A2(n14818), .ZN(n9574) );
  NAND2_X1 U12104 ( .A1(n9575), .A2(n9574), .ZN(n9577) );
  INV_X1 U12105 ( .A(n9641), .ZN(n9770) );
  AOI22_X1 U12106 ( .A1(n13206), .A2(n9770), .B1(n9761), .B2(n14818), .ZN(
        n9576) );
  NOR2_X1 U12107 ( .A1(n9578), .A2(n9577), .ZN(n9579) );
  NAND2_X1 U12108 ( .A1(n13205), .A2(n9770), .ZN(n9582) );
  NAND2_X1 U12109 ( .A1(n9761), .A2(n10927), .ZN(n9581) );
  NAND2_X1 U12110 ( .A1(n9582), .A2(n9581), .ZN(n9586) );
  NAND2_X1 U12111 ( .A1(n13205), .A2(n9761), .ZN(n9583) );
  OAI21_X1 U12112 ( .B1(n11223), .B2(n9761), .A(n9583), .ZN(n9584) );
  INV_X1 U12113 ( .A(n9586), .ZN(n9587) );
  NAND2_X1 U12114 ( .A1(n14964), .A2(n9769), .ZN(n9589) );
  NAND2_X1 U12115 ( .A1(n13204), .A2(n9761), .ZN(n9588) );
  NAND2_X1 U12116 ( .A1(n9589), .A2(n9588), .ZN(n9591) );
  AOI22_X1 U12117 ( .A1(n14964), .A2(n9727), .B1(n13204), .B2(n9769), .ZN(
        n9590) );
  NOR2_X1 U12118 ( .A1(n9592), .A2(n9591), .ZN(n9593) );
  NAND2_X1 U12119 ( .A1(n10959), .A2(n9761), .ZN(n9596) );
  NAND2_X1 U12120 ( .A1(n13203), .A2(n9769), .ZN(n9595) );
  NAND2_X1 U12121 ( .A1(n9596), .A2(n9595), .ZN(n9600) );
  NAND2_X1 U12122 ( .A1(n10959), .A2(n9769), .ZN(n9597) );
  OAI21_X1 U12123 ( .B1(n11191), .B2(n9769), .A(n9597), .ZN(n9598) );
  INV_X1 U12124 ( .A(n9600), .ZN(n9601) );
  NAND2_X1 U12125 ( .A1(n11038), .A2(n9769), .ZN(n9603) );
  NAND2_X1 U12126 ( .A1(n13202), .A2(n9727), .ZN(n9602) );
  NAND2_X1 U12127 ( .A1(n9603), .A2(n9602), .ZN(n9605) );
  AOI22_X1 U12128 ( .A1(n11038), .A2(n9761), .B1(n13202), .B2(n9769), .ZN(
        n9604) );
  AOI21_X1 U12129 ( .B1(n9606), .B2(n9605), .A(n9604), .ZN(n9608) );
  OR2_X1 U12130 ( .A1(n9608), .A2(n9607), .ZN(n9616) );
  NAND2_X1 U12131 ( .A1(n11180), .A2(n9761), .ZN(n9610) );
  NAND2_X1 U12132 ( .A1(n13201), .A2(n9770), .ZN(n9609) );
  NAND2_X1 U12133 ( .A1(n9610), .A2(n9609), .ZN(n9615) );
  NAND2_X1 U12134 ( .A1(n9616), .A2(n9615), .ZN(n9614) );
  NAND2_X1 U12135 ( .A1(n11180), .A2(n9770), .ZN(n9612) );
  NOR2_X1 U12136 ( .A1(n9616), .A2(n9615), .ZN(n9617) );
  NAND2_X1 U12137 ( .A1(n11363), .A2(n9769), .ZN(n9619) );
  NAND2_X1 U12138 ( .A1(n13200), .A2(n9761), .ZN(n9618) );
  AOI22_X1 U12139 ( .A1(n11363), .A2(n9761), .B1(n13200), .B2(n9769), .ZN(
        n9620) );
  NAND2_X1 U12140 ( .A1(n11493), .A2(n9727), .ZN(n9622) );
  NAND2_X1 U12141 ( .A1(n13199), .A2(n9769), .ZN(n9621) );
  NAND2_X1 U12142 ( .A1(n9622), .A2(n9621), .ZN(n9624) );
  AOI22_X1 U12143 ( .A1(n11493), .A2(n9770), .B1(n9761), .B2(n13199), .ZN(
        n9623) );
  NAND2_X1 U12144 ( .A1(n13526), .A2(n9769), .ZN(n9626) );
  NAND2_X1 U12145 ( .A1(n13198), .A2(n9761), .ZN(n9625) );
  NAND2_X1 U12146 ( .A1(n13526), .A2(n9761), .ZN(n9627) );
  OAI21_X1 U12147 ( .B1(n11276), .B2(n9727), .A(n9627), .ZN(n9628) );
  NAND2_X1 U12148 ( .A1(n11741), .A2(n9761), .ZN(n9630) );
  NAND2_X1 U12149 ( .A1(n13197), .A2(n9769), .ZN(n9629) );
  NAND2_X1 U12150 ( .A1(n9630), .A2(n9629), .ZN(n9633) );
  AOI22_X1 U12151 ( .A1(n11741), .A2(n9770), .B1(n9761), .B2(n13197), .ZN(
        n9631) );
  AOI21_X1 U12152 ( .B1(n9634), .B2(n9633), .A(n9631), .ZN(n9632) );
  NOR2_X1 U12153 ( .A1(n9634), .A2(n9633), .ZN(n9635) );
  NAND2_X1 U12154 ( .A1(n14830), .A2(n9770), .ZN(n9637) );
  NAND2_X1 U12155 ( .A1(n11566), .A2(n9727), .ZN(n9636) );
  NAND2_X1 U12156 ( .A1(n14830), .A2(n9727), .ZN(n9638) );
  OAI21_X1 U12157 ( .B1(n9639), .B2(n9761), .A(n9638), .ZN(n9640) );
  NAND2_X1 U12158 ( .A1(n13510), .A2(n9641), .ZN(n9643) );
  NAND2_X1 U12159 ( .A1(n13196), .A2(n9769), .ZN(n9642) );
  NAND2_X1 U12160 ( .A1(n9643), .A2(n9642), .ZN(n9645) );
  AOI22_X1 U12161 ( .A1(n13510), .A2(n9770), .B1(n9727), .B2(n13196), .ZN(
        n9644) );
  AOI21_X1 U12162 ( .B1(n9646), .B2(n9645), .A(n9644), .ZN(n9658) );
  NOR2_X1 U12163 ( .A1(n9646), .A2(n9645), .ZN(n9657) );
  AND2_X1 U12164 ( .A1(n13193), .A2(n9727), .ZN(n9647) );
  AOI21_X1 U12165 ( .B1(n12073), .B2(n9769), .A(n9647), .ZN(n9670) );
  NAND2_X1 U12166 ( .A1(n12073), .A2(n9727), .ZN(n9649) );
  NAND2_X1 U12167 ( .A1(n13193), .A2(n9769), .ZN(n9648) );
  NAND2_X1 U12168 ( .A1(n9649), .A2(n9648), .ZN(n9668) );
  AND2_X1 U12169 ( .A1(n13194), .A2(n9727), .ZN(n9650) );
  AOI21_X1 U12170 ( .B1(n13477), .B2(n9769), .A(n9650), .ZN(n9664) );
  NAND2_X1 U12171 ( .A1(n13477), .A2(n9727), .ZN(n9652) );
  NAND2_X1 U12172 ( .A1(n13194), .A2(n9769), .ZN(n9651) );
  NAND2_X1 U12173 ( .A1(n9652), .A2(n9651), .ZN(n9663) );
  AOI22_X1 U12174 ( .A1(n9670), .A2(n9668), .B1(n9664), .B2(n9663), .ZN(n9659)
         );
  AND2_X1 U12175 ( .A1(n13195), .A2(n9727), .ZN(n9653) );
  AOI21_X1 U12176 ( .B1(n13672), .B2(n9769), .A(n9653), .ZN(n9661) );
  NAND2_X1 U12177 ( .A1(n13672), .A2(n9761), .ZN(n9655) );
  NAND2_X1 U12178 ( .A1(n13195), .A2(n9769), .ZN(n9654) );
  NAND2_X1 U12179 ( .A1(n9655), .A2(n9654), .ZN(n9660) );
  NAND2_X1 U12180 ( .A1(n9661), .A2(n9660), .ZN(n9656) );
  INV_X1 U12181 ( .A(n9659), .ZN(n9662) );
  OR3_X1 U12182 ( .A1(n9662), .A2(n9661), .A3(n9660), .ZN(n9676) );
  INV_X1 U12183 ( .A(n9663), .ZN(n9666) );
  INV_X1 U12184 ( .A(n9664), .ZN(n9665) );
  NAND2_X1 U12185 ( .A1(n9666), .A2(n9665), .ZN(n9669) );
  NAND3_X1 U12186 ( .A1(n9669), .A2(n9667), .A3(n13665), .ZN(n9674) );
  INV_X1 U12187 ( .A(n9668), .ZN(n9673) );
  INV_X1 U12188 ( .A(n9669), .ZN(n9672) );
  INV_X1 U12189 ( .A(n9670), .ZN(n9671) );
  AOI22_X1 U12190 ( .A1(n9674), .A2(n9673), .B1(n9672), .B2(n9671), .ZN(n9675)
         );
  AND2_X1 U12191 ( .A1(n9676), .A2(n9675), .ZN(n9677) );
  AND2_X1 U12192 ( .A1(n13192), .A2(n9769), .ZN(n9678) );
  AOI21_X1 U12193 ( .B1(n13601), .B2(n9727), .A(n9678), .ZN(n9681) );
  NAND2_X1 U12194 ( .A1(n13601), .A2(n9770), .ZN(n9679) );
  OAI21_X1 U12195 ( .B1(n9350), .B2(n9770), .A(n9679), .ZN(n9680) );
  NAND2_X1 U12196 ( .A1(n13596), .A2(n9770), .ZN(n9683) );
  NAND2_X1 U12197 ( .A1(n13191), .A2(n9761), .ZN(n9682) );
  NAND2_X1 U12198 ( .A1(n9683), .A2(n9682), .ZN(n9685) );
  AOI22_X1 U12199 ( .A1(n13596), .A2(n9727), .B1(n13191), .B2(n9769), .ZN(
        n9684) );
  AOI21_X1 U12200 ( .B1(n9686), .B2(n9685), .A(n9684), .ZN(n9688) );
  NOR2_X1 U12201 ( .A1(n9686), .A2(n9685), .ZN(n9687) );
  OR2_X1 U12202 ( .A1(n9688), .A2(n9687), .ZN(n9694) );
  NAND2_X1 U12203 ( .A1(n13590), .A2(n9727), .ZN(n9690) );
  NAND2_X1 U12204 ( .A1(n13190), .A2(n9769), .ZN(n9689) );
  NAND2_X1 U12205 ( .A1(n9690), .A2(n9689), .ZN(n9693) );
  AOI22_X1 U12206 ( .A1(n13590), .A2(n9770), .B1(n9761), .B2(n13190), .ZN(
        n9691) );
  AOI21_X1 U12207 ( .B1(n9694), .B2(n9693), .A(n9691), .ZN(n9692) );
  INV_X1 U12208 ( .A(n9692), .ZN(n9695) );
  NAND2_X1 U12209 ( .A1(n13404), .A2(n9769), .ZN(n9697) );
  NAND2_X1 U12210 ( .A1(n13189), .A2(n9727), .ZN(n9696) );
  NAND2_X1 U12211 ( .A1(n9697), .A2(n9696), .ZN(n9699) );
  AOI22_X1 U12212 ( .A1(n13404), .A2(n9727), .B1(n13189), .B2(n9769), .ZN(
        n9698) );
  NAND2_X1 U12213 ( .A1(n13580), .A2(n9727), .ZN(n9702) );
  NAND2_X1 U12214 ( .A1(n13188), .A2(n9770), .ZN(n9701) );
  NAND2_X1 U12215 ( .A1(n13580), .A2(n9769), .ZN(n9703) );
  OAI21_X1 U12216 ( .B1(n9704), .B2(n9769), .A(n9703), .ZN(n9705) );
  NAND2_X1 U12217 ( .A1(n13375), .A2(n9769), .ZN(n9707) );
  NAND2_X1 U12218 ( .A1(n13187), .A2(n9727), .ZN(n9706) );
  NAND2_X1 U12219 ( .A1(n9707), .A2(n9706), .ZN(n9709) );
  AOI22_X1 U12220 ( .A1(n13375), .A2(n9761), .B1(n13187), .B2(n9769), .ZN(
        n9708) );
  AOI21_X1 U12221 ( .B1(n9710), .B2(n9709), .A(n9708), .ZN(n9712) );
  NOR2_X1 U12222 ( .A1(n9710), .A2(n9709), .ZN(n9711) );
  NAND2_X1 U12223 ( .A1(n13567), .A2(n9761), .ZN(n9714) );
  NAND2_X1 U12224 ( .A1(n13186), .A2(n9769), .ZN(n9713) );
  AOI22_X1 U12225 ( .A1(n13567), .A2(n9769), .B1(n9761), .B2(n13186), .ZN(
        n9715) );
  AND2_X1 U12226 ( .A1(n13185), .A2(n9761), .ZN(n9716) );
  AOI21_X1 U12227 ( .B1(n13562), .B2(n9769), .A(n9716), .ZN(n9719) );
  NAND2_X1 U12228 ( .A1(n13562), .A2(n9761), .ZN(n9717) );
  OAI21_X1 U12229 ( .B1(n13128), .B2(n9727), .A(n9717), .ZN(n9718) );
  NAND2_X1 U12230 ( .A1(n13557), .A2(n9761), .ZN(n9721) );
  NAND2_X1 U12231 ( .A1(n13184), .A2(n9769), .ZN(n9720) );
  NAND2_X1 U12232 ( .A1(n13557), .A2(n9769), .ZN(n9722) );
  OAI21_X1 U12233 ( .B1(n13118), .B2(n9769), .A(n9722), .ZN(n9723) );
  NAND2_X1 U12234 ( .A1(n13317), .A2(n9769), .ZN(n9726) );
  NAND2_X1 U12235 ( .A1(n13183), .A2(n9727), .ZN(n9725) );
  NAND2_X1 U12236 ( .A1(n9726), .A2(n9725), .ZN(n9733) );
  NAND2_X1 U12237 ( .A1(n9732), .A2(n9733), .ZN(n9731) );
  NAND2_X1 U12238 ( .A1(n13317), .A2(n9727), .ZN(n9729) );
  NAND2_X1 U12239 ( .A1(n13183), .A2(n9769), .ZN(n9728) );
  NAND2_X1 U12240 ( .A1(n9729), .A2(n9728), .ZN(n9730) );
  NAND2_X1 U12241 ( .A1(n9731), .A2(n9730), .ZN(n9837) );
  INV_X1 U12242 ( .A(n9733), .ZN(n9734) );
  NAND2_X1 U12243 ( .A1(n9735), .A2(n9734), .ZN(n9835) );
  NAND2_X1 U12244 ( .A1(n9737), .A2(n9736), .ZN(n9740) );
  INV_X1 U12245 ( .A(SI_29_), .ZN(n13022) );
  NAND2_X1 U12246 ( .A1(n9738), .A2(n13022), .ZN(n9739) );
  MUX2_X1 U12247 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9874), .Z(n9741) );
  NAND2_X1 U12248 ( .A1(n9741), .A2(SI_30_), .ZN(n9742) );
  OAI21_X1 U12249 ( .B1(SI_30_), .B2(n9741), .A(n9742), .ZN(n9754) );
  MUX2_X1 U12250 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6533), .Z(n9743) );
  XNOR2_X1 U12251 ( .A(n9743), .B(SI_31_), .ZN(n9744) );
  NAND2_X1 U12252 ( .A1(n13683), .A2(n9746), .ZN(n9748) );
  OR2_X1 U12253 ( .A1(n6544), .A2(n13686), .ZN(n9747) );
  NAND2_X2 U12254 ( .A1(n9748), .A2(n9747), .ZN(n9821) );
  INV_X1 U12255 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n10333) );
  NAND2_X1 U12256 ( .A1(n9749), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9752) );
  NAND2_X1 U12257 ( .A1(n9750), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9751) );
  OAI211_X1 U12258 ( .C1(n9753), .C2(n10333), .A(n9752), .B(n9751), .ZN(n13283) );
  NAND2_X1 U12259 ( .A1(n9755), .A2(n9754), .ZN(n9756) );
  INV_X1 U12260 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13690) );
  OR2_X1 U12261 ( .A1(n6545), .A2(n13690), .ZN(n9758) );
  NAND2_X1 U12262 ( .A1(n13283), .A2(n9819), .ZN(n9820) );
  NAND2_X1 U12263 ( .A1(n9843), .A2(n6840), .ZN(n9801) );
  NAND4_X1 U12264 ( .A1(n9820), .A2(n6841), .A3(n9801), .A4(n9842), .ZN(n9759)
         );
  AND2_X1 U12265 ( .A1(n9759), .A2(n13180), .ZN(n9760) );
  AOI21_X1 U12266 ( .B1(n13281), .B2(n9761), .A(n9760), .ZN(n9813) );
  NAND2_X1 U12267 ( .A1(n13281), .A2(n9769), .ZN(n9763) );
  NAND2_X1 U12268 ( .A1(n13180), .A2(n9761), .ZN(n9762) );
  NAND2_X1 U12269 ( .A1(n9763), .A2(n9762), .ZN(n9812) );
  AND2_X1 U12270 ( .A1(n13181), .A2(n9769), .ZN(n9764) );
  AOI21_X1 U12271 ( .B1(n13542), .B2(n9761), .A(n9764), .ZN(n9807) );
  NAND2_X1 U12272 ( .A1(n13542), .A2(n9769), .ZN(n9766) );
  NAND2_X1 U12273 ( .A1(n13181), .A2(n9727), .ZN(n9765) );
  NAND2_X1 U12274 ( .A1(n9766), .A2(n9765), .ZN(n9806) );
  OAI22_X1 U12275 ( .A1(n9813), .A2(n9812), .B1(n9807), .B2(n9806), .ZN(n9767)
         );
  NAND2_X1 U12276 ( .A1(n9809), .A2(n9767), .ZN(n9811) );
  AND2_X1 U12277 ( .A1(n13182), .A2(n9761), .ZN(n9768) );
  AOI21_X1 U12278 ( .B1(n13548), .B2(n9769), .A(n9768), .ZN(n9803) );
  NAND2_X1 U12279 ( .A1(n13548), .A2(n9727), .ZN(n9772) );
  NAND2_X1 U12280 ( .A1(n13182), .A2(n9770), .ZN(n9771) );
  NAND2_X1 U12281 ( .A1(n9772), .A2(n9771), .ZN(n9802) );
  NAND2_X1 U12282 ( .A1(n9803), .A2(n9802), .ZN(n9773) );
  NOR2_X1 U12283 ( .A1(n9777), .A2(n9776), .ZN(n13506) );
  OAI21_X1 U12284 ( .B1(n9559), .B2(n10897), .A(n10573), .ZN(n14961) );
  NAND3_X1 U12285 ( .A1(n9778), .A2(n9798), .A3(n14961), .ZN(n9779) );
  NOR4_X1 U12286 ( .A1(n10533), .A2(n10575), .A3(n9779), .A4(n10564), .ZN(
        n9780) );
  XNOR2_X1 U12287 ( .A(n14964), .B(n13204), .ZN(n11120) );
  NAND4_X1 U12288 ( .A1(n11297), .A2(n11283), .A3(n9780), .A4(n11120), .ZN(
        n9781) );
  NOR4_X1 U12289 ( .A1(n9783), .A2(n11422), .A3(n9782), .A4(n9781), .ZN(n9784)
         );
  XNOR2_X1 U12290 ( .A(n14830), .B(n11566), .ZN(n11663) );
  NAND4_X1 U12291 ( .A1(n9784), .A2(n11596), .A3(n11663), .A4(n11578), .ZN(
        n9785) );
  NOR4_X1 U12292 ( .A1(n9786), .A2(n13506), .A3(n13451), .A4(n9785), .ZN(n9788) );
  NAND4_X1 U12293 ( .A1(n13426), .A2(n9788), .A3(n9787), .A4(n13486), .ZN(
        n9789) );
  NOR4_X1 U12294 ( .A1(n13385), .A2(n13399), .A3(n9790), .A4(n9789), .ZN(n9791) );
  XNOR2_X1 U12295 ( .A(n13375), .B(n13187), .ZN(n13371) );
  NAND4_X1 U12296 ( .A1(n13335), .A2(n9791), .A3(n13371), .A4(n13357), .ZN(
        n9792) );
  NOR4_X1 U12297 ( .A1(n13292), .A2(n13308), .A3(n13344), .A4(n9792), .ZN(
        n9795) );
  XNOR2_X1 U12298 ( .A(n13281), .B(n13180), .ZN(n9793) );
  XNOR2_X1 U12299 ( .A(n9796), .B(n9799), .ZN(n9797) );
  NAND2_X1 U12300 ( .A1(n9797), .A2(n12419), .ZN(n9824) );
  NAND3_X1 U12301 ( .A1(n6841), .A2(n9799), .A3(n9798), .ZN(n9800) );
  AND2_X1 U12302 ( .A1(n9801), .A2(n9800), .ZN(n9830) );
  INV_X1 U12303 ( .A(n9802), .ZN(n9805) );
  INV_X1 U12304 ( .A(n9803), .ZN(n9804) );
  AOI22_X1 U12305 ( .A1(n9807), .A2(n9806), .B1(n9805), .B2(n9804), .ZN(n9808)
         );
  NAND2_X1 U12306 ( .A1(n9809), .A2(n9808), .ZN(n9810) );
  NAND2_X1 U12307 ( .A1(n9811), .A2(n9810), .ZN(n9815) );
  NAND2_X1 U12308 ( .A1(n9813), .A2(n9812), .ZN(n9814) );
  NAND2_X1 U12309 ( .A1(n9815), .A2(n9814), .ZN(n9825) );
  NAND2_X1 U12310 ( .A1(n13283), .A2(n9761), .ZN(n9823) );
  NAND2_X1 U12311 ( .A1(n9820), .A2(n9819), .ZN(n9822) );
  MUX2_X1 U12312 ( .A(n9823), .B(n9822), .S(n9821), .Z(n9831) );
  INV_X1 U12313 ( .A(n9825), .ZN(n9829) );
  INV_X1 U12314 ( .A(n9826), .ZN(n10405) );
  INV_X1 U12315 ( .A(n9842), .ZN(n10414) );
  AOI21_X1 U12316 ( .B1(n6841), .B2(n13276), .A(n10414), .ZN(n9827) );
  OAI21_X1 U12317 ( .B1(n10405), .B2(n9843), .A(n9827), .ZN(n9828) );
  NAND2_X1 U12318 ( .A1(n9831), .A2(n9828), .ZN(n9834) );
  NAND3_X1 U12319 ( .A1(n9837), .A2(n9836), .A3(n9835), .ZN(n9838) );
  OR2_X1 U12320 ( .A1(n10090), .A2(P2_U3088), .ZN(n11856) );
  INV_X1 U12321 ( .A(n11856), .ZN(n9839) );
  OAI21_X1 U12322 ( .B1(n9841), .B2(n9840), .A(n9839), .ZN(n9847) );
  NOR4_X1 U12323 ( .A1(n14957), .A2(n13135), .A3(n9842), .A4(n13701), .ZN(
        n9845) );
  OAI21_X1 U12324 ( .B1(n11856), .B2(n9843), .A(P2_B_REG_SCAN_IN), .ZN(n9844)
         );
  NAND2_X1 U12325 ( .A1(n9847), .A2(n9846), .ZN(P2_U3328) );
  INV_X1 U12326 ( .A(n9848), .ZN(n9849) );
  NAND2_X1 U12327 ( .A1(n9849), .A2(n10090), .ZN(n10094) );
  NOR2_X4 U12328 ( .A1(n10607), .A2(n9931), .ZN(P3_U3897) );
  INV_X1 U12329 ( .A(n9850), .ZN(n9906) );
  INV_X2 U12330 ( .A(n13849), .ZN(P1_U4016) );
  AND2_X1 U12331 ( .A1(n9874), .A2(P2_U3088), .ZN(n13694) );
  INV_X2 U12332 ( .A(n13694), .ZN(n13708) );
  AND2_X1 U12333 ( .A1(n9854), .A2(P2_U3088), .ZN(n9911) );
  NOR2_X1 U12334 ( .A1(n10097), .A2(P2_U3088), .ZN(n14840) );
  AOI21_X1 U12335 ( .B1(n9911), .B2(P1_DATAO_REG_1__SCAN_IN), .A(n14840), .ZN(
        n9852) );
  OAI21_X1 U12336 ( .B1(n9877), .B2(n13708), .A(n9852), .ZN(P2_U3326) );
  AND2_X1 U12337 ( .A1(n9854), .A2(P3_U3151), .ZN(n11150) );
  INV_X2 U12338 ( .A(n11150), .ZN(n13021) );
  NAND2_X1 U12339 ( .A1(n6532), .A2(P3_U3151), .ZN(n13023) );
  INV_X1 U12340 ( .A(SI_5_), .ZN(n9855) );
  OAI222_X1 U12341 ( .A1(n13021), .A2(n9856), .B1(n13023), .B2(n9855), .C1(
        n15014), .C2(P3_U3151), .ZN(P3_U3290) );
  INV_X1 U12342 ( .A(SI_2_), .ZN(n9857) );
  OAI222_X1 U12343 ( .A1(n13021), .A2(n9858), .B1(n13023), .B2(n9857), .C1(
        n6709), .C2(P3_U3151), .ZN(P3_U3293) );
  INV_X1 U12344 ( .A(SI_3_), .ZN(n9859) );
  OAI222_X1 U12345 ( .A1(n13021), .A2(n9860), .B1(n13023), .B2(n9859), .C1(
        n10490), .C2(P3_U3151), .ZN(P3_U3292) );
  INV_X1 U12346 ( .A(SI_4_), .ZN(n9861) );
  OAI222_X1 U12347 ( .A1(n13021), .A2(n9862), .B1(n13023), .B2(n9861), .C1(
        n12626), .C2(P3_U3151), .ZN(P3_U3291) );
  INV_X1 U12348 ( .A(SI_7_), .ZN(n9863) );
  OAI222_X1 U12349 ( .A1(n13021), .A2(n9864), .B1(n13023), .B2(n9863), .C1(
        n15052), .C2(P3_U3151), .ZN(P3_U3288) );
  INV_X1 U12350 ( .A(n10448), .ZN(n10781) );
  INV_X1 U12351 ( .A(n9865), .ZN(n9866) );
  OAI222_X1 U12352 ( .A1(P3_U3151), .A2(n10781), .B1(n13023), .B2(n6712), .C1(
        n13021), .C2(n9866), .ZN(P3_U3294) );
  INV_X2 U12353 ( .A(n9911), .ZN(n13705) );
  OAI222_X1 U12354 ( .A1(n13705), .A2(n9867), .B1(n13708), .B2(n9875), .C1(
        P2_U3088), .C2(n14853), .ZN(P2_U3325) );
  OAI222_X1 U12355 ( .A1(P2_U3088), .A2(n10100), .B1(n13708), .B2(n9898), .C1(
        n9868), .C2(n13705), .ZN(P2_U3324) );
  INV_X1 U12356 ( .A(n12640), .ZN(n15066) );
  INV_X1 U12357 ( .A(SI_8_), .ZN(n9871) );
  INV_X1 U12358 ( .A(n9869), .ZN(n9870) );
  OAI222_X1 U12359 ( .A1(P3_U3151), .A2(n15066), .B1(n13023), .B2(n9871), .C1(
        n13021), .C2(n9870), .ZN(P3_U3287) );
  INV_X1 U12360 ( .A(SI_9_), .ZN(n9872) );
  OAI222_X1 U12361 ( .A1(n13021), .A2(n9873), .B1(n13023), .B2(n9872), .C1(
        n15083), .C2(P3_U3151), .ZN(P3_U3286) );
  NOR2_X1 U12362 ( .A1(n6533), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14210) );
  INV_X2 U12363 ( .A(n14210), .ZN(n14225) );
  OAI222_X1 U12364 ( .A1(n14216), .A2(n9876), .B1(n10139), .B2(P1_U3086), .C1(
        n14225), .C2(n9875), .ZN(P1_U3353) );
  OAI222_X1 U12365 ( .A1(n14216), .A2(n6715), .B1(n13868), .B2(P1_U3086), .C1(
        n14225), .C2(n9877), .ZN(P1_U3354) );
  OAI222_X1 U12366 ( .A1(P2_U3088), .A2(n14868), .B1(n13708), .B2(n9880), .C1(
        n9878), .C2(n13705), .ZN(P2_U3323) );
  OAI222_X1 U12367 ( .A1(n14225), .A2(n9880), .B1(n6884), .B2(P1_U3086), .C1(
        n9879), .C2(n14216), .ZN(P1_U3351) );
  OAI222_X1 U12368 ( .A1(n14225), .A2(n9888), .B1(n10014), .B2(P1_U3086), .C1(
        n9881), .C2(n14216), .ZN(P1_U3350) );
  INV_X1 U12369 ( .A(n13023), .ZN(n13014) );
  INV_X1 U12370 ( .A(SI_10_), .ZN(n9882) );
  OAI222_X1 U12371 ( .A1(n13021), .A2(n9883), .B1(n11761), .B2(n9882), .C1(
        n15100), .C2(P3_U3151), .ZN(P3_U3285) );
  INV_X1 U12372 ( .A(n12632), .ZN(n15028) );
  INV_X1 U12373 ( .A(n9884), .ZN(n9886) );
  INV_X1 U12374 ( .A(SI_6_), .ZN(n9885) );
  OAI222_X1 U12375 ( .A1(n15028), .A2(P3_U3151), .B1(n13021), .B2(n9886), .C1(
        n9885), .C2(n11761), .ZN(P3_U3289) );
  INV_X1 U12376 ( .A(n10102), .ZN(n10129) );
  OAI222_X1 U12377 ( .A1(P2_U3088), .A2(n10129), .B1(n13708), .B2(n9888), .C1(
        n9887), .C2(n13705), .ZN(P2_U3322) );
  OAI222_X1 U12378 ( .A1(n13021), .A2(n9890), .B1(n13023), .B2(n9889), .C1(
        n15117), .C2(P3_U3151), .ZN(P3_U3284) );
  INV_X1 U12379 ( .A(n9990), .ZN(n10027) );
  OAI222_X1 U12380 ( .A1(n14225), .A2(n9893), .B1(n10027), .B2(P1_U3086), .C1(
        n9891), .C2(n14216), .ZN(P1_U3349) );
  INV_X1 U12381 ( .A(n14883), .ZN(n9894) );
  OAI222_X1 U12382 ( .A1(P2_U3088), .A2(n9894), .B1(n13708), .B2(n9893), .C1(
        n9892), .C2(n13705), .ZN(P2_U3321) );
  OAI222_X1 U12383 ( .A1(n13021), .A2(n9896), .B1(n15135), .B2(P3_U3151), .C1(
        n9895), .C2(n11761), .ZN(P3_U3283) );
  OAI222_X1 U12384 ( .A1(n14225), .A2(n9898), .B1(n13878), .B2(P1_U3086), .C1(
        n9897), .C2(n14216), .ZN(P1_U3352) );
  INV_X1 U12385 ( .A(n10036), .ZN(n9998) );
  OAI222_X1 U12386 ( .A1(n14225), .A2(n9901), .B1(n9998), .B2(P1_U3086), .C1(
        n9899), .C2(n14216), .ZN(P1_U3348) );
  INV_X1 U12387 ( .A(n10103), .ZN(n11927) );
  OAI222_X1 U12388 ( .A1(P2_U3088), .A2(n11927), .B1(n13708), .B2(n9901), .C1(
        n9900), .C2(n13705), .ZN(P2_U3320) );
  NAND2_X1 U12389 ( .A1(n9902), .A2(n9910), .ZN(n9903) );
  OAI21_X1 U12390 ( .B1(n9910), .B2(n8987), .A(n9903), .ZN(P3_U3376) );
  NAND2_X1 U12391 ( .A1(n10072), .A2(n9904), .ZN(n14739) );
  INV_X1 U12392 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9907) );
  NOR2_X1 U12393 ( .A1(n9906), .A2(n9905), .ZN(n11912) );
  AOI22_X1 U12394 ( .A1(n6674), .A2(n9907), .B1(n11912), .B2(n11860), .ZN(
        P1_U3445) );
  NAND2_X1 U12395 ( .A1(n9908), .A2(n9910), .ZN(n9909) );
  OAI21_X1 U12396 ( .B1(n9910), .B2(n8990), .A(n9909), .ZN(P3_U3377) );
  NAND2_X1 U12397 ( .A1(n10105), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14894) );
  NAND2_X1 U12398 ( .A1(n9911), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n9912) );
  OAI211_X1 U12399 ( .C1(n9914), .C2(n13708), .A(n14894), .B(n9912), .ZN(
        P2_U3319) );
  INV_X1 U12400 ( .A(n10198), .ZN(n10201) );
  OAI222_X1 U12401 ( .A1(n14225), .A2(n9914), .B1(n10201), .B2(P1_U3086), .C1(
        n9913), .C2(n14216), .ZN(P1_U3347) );
  OAI222_X1 U12402 ( .A1(n13021), .A2(n9916), .B1(n11761), .B2(n9915), .C1(
        n15151), .C2(P3_U3151), .ZN(P3_U3282) );
  INV_X1 U12403 ( .A(n10072), .ZN(n9918) );
  INV_X1 U12404 ( .A(n9919), .ZN(n9917) );
  NAND2_X1 U12405 ( .A1(n9917), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12324) );
  NAND2_X1 U12406 ( .A1(n9918), .A2(n12324), .ZN(n9976) );
  NAND2_X1 U12407 ( .A1(n9920), .A2(n9919), .ZN(n9922) );
  AND2_X1 U12408 ( .A1(n9922), .A2(n7676), .ZN(n9975) );
  INV_X1 U12409 ( .A(n9975), .ZN(n9923) );
  NOR2_X1 U12410 ( .A1(n14615), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12411 ( .A(n10518), .ZN(n9925) );
  OAI222_X1 U12412 ( .A1(n14225), .A2(n9927), .B1(n9925), .B2(P1_U3086), .C1(
        n9924), .C2(n14216), .ZN(P1_U3346) );
  INV_X1 U12413 ( .A(n10744), .ZN(n10113) );
  OAI222_X1 U12414 ( .A1(P2_U3088), .A2(n10113), .B1(n13708), .B2(n9927), .C1(
        n9926), .C2(n13705), .ZN(P2_U3318) );
  INV_X1 U12415 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n10356) );
  NAND2_X1 U12416 ( .A1(n11016), .A2(P3_U3897), .ZN(n9928) );
  OAI21_X1 U12417 ( .B1(P3_U3897), .B2(n10356), .A(n9928), .ZN(P3_U3494) );
  OAI222_X1 U12418 ( .A1(n13021), .A2(n9930), .B1(n13023), .B2(n9929), .C1(
        n15169), .C2(P3_U3151), .ZN(P3_U3281) );
  NOR2_X1 U12419 ( .A1(n8989), .A2(n9931), .ZN(n9934) );
  INV_X1 U12420 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n9932) );
  NOR2_X1 U12421 ( .A1(n9963), .A2(n9932), .ZN(P3_U3236) );
  INV_X1 U12422 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n9933) );
  NOR2_X1 U12423 ( .A1(n9934), .A2(n9933), .ZN(P3_U3238) );
  CLKBUF_X1 U12424 ( .A(n9934), .Z(n9963) );
  INV_X1 U12425 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n9935) );
  NOR2_X1 U12426 ( .A1(n9963), .A2(n9935), .ZN(P3_U3251) );
  INV_X1 U12427 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n9936) );
  NOR2_X1 U12428 ( .A1(n9963), .A2(n9936), .ZN(P3_U3250) );
  INV_X1 U12429 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n9937) );
  NOR2_X1 U12430 ( .A1(n9934), .A2(n9937), .ZN(P3_U3237) );
  INV_X1 U12431 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n9938) );
  NOR2_X1 U12432 ( .A1(n9934), .A2(n9938), .ZN(P3_U3235) );
  INV_X1 U12433 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n9939) );
  NOR2_X1 U12434 ( .A1(n9934), .A2(n9939), .ZN(P3_U3240) );
  INV_X1 U12435 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n9940) );
  NOR2_X1 U12436 ( .A1(n9934), .A2(n9940), .ZN(P3_U3239) );
  INV_X1 U12437 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9941) );
  NOR2_X1 U12438 ( .A1(n9934), .A2(n9941), .ZN(P3_U3262) );
  INV_X1 U12439 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n9942) );
  NOR2_X1 U12440 ( .A1(n9963), .A2(n9942), .ZN(P3_U3252) );
  INV_X1 U12441 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n9943) );
  NOR2_X1 U12442 ( .A1(n9934), .A2(n9943), .ZN(P3_U3260) );
  INV_X1 U12443 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n9944) );
  NOR2_X1 U12444 ( .A1(n9963), .A2(n9944), .ZN(P3_U3259) );
  INV_X1 U12445 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n9945) );
  NOR2_X1 U12446 ( .A1(n9934), .A2(n9945), .ZN(P3_U3258) );
  INV_X1 U12447 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n9946) );
  NOR2_X1 U12448 ( .A1(n9963), .A2(n9946), .ZN(P3_U3257) );
  INV_X1 U12449 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n9947) );
  NOR2_X1 U12450 ( .A1(n9963), .A2(n9947), .ZN(P3_U3256) );
  INV_X1 U12451 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n9948) );
  NOR2_X1 U12452 ( .A1(n9963), .A2(n9948), .ZN(P3_U3263) );
  INV_X1 U12453 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n9949) );
  NOR2_X1 U12454 ( .A1(n9963), .A2(n9949), .ZN(P3_U3254) );
  INV_X1 U12455 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n9950) );
  NOR2_X1 U12456 ( .A1(n9963), .A2(n9950), .ZN(P3_U3261) );
  INV_X1 U12457 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n9951) );
  NOR2_X1 U12458 ( .A1(n9963), .A2(n9951), .ZN(P3_U3246) );
  INV_X1 U12459 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n9952) );
  NOR2_X1 U12460 ( .A1(n9934), .A2(n9952), .ZN(P3_U3245) );
  INV_X1 U12461 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n9953) );
  NOR2_X1 U12462 ( .A1(n9934), .A2(n9953), .ZN(P3_U3244) );
  INV_X1 U12463 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n9954) );
  NOR2_X1 U12464 ( .A1(n9934), .A2(n9954), .ZN(P3_U3234) );
  INV_X1 U12465 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n9955) );
  NOR2_X1 U12466 ( .A1(n9963), .A2(n9955), .ZN(P3_U3242) );
  INV_X1 U12467 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n9956) );
  NOR2_X1 U12468 ( .A1(n9963), .A2(n9956), .ZN(P3_U3255) );
  INV_X1 U12469 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n9957) );
  NOR2_X1 U12470 ( .A1(n9963), .A2(n9957), .ZN(P3_U3248) );
  INV_X1 U12471 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9958) );
  NOR2_X1 U12472 ( .A1(n9963), .A2(n9958), .ZN(P3_U3247) );
  INV_X1 U12473 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n9959) );
  NOR2_X1 U12474 ( .A1(n9963), .A2(n9959), .ZN(P3_U3243) );
  INV_X1 U12475 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n9960) );
  NOR2_X1 U12476 ( .A1(n9963), .A2(n9960), .ZN(P3_U3249) );
  INV_X1 U12477 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n9961) );
  NOR2_X1 U12478 ( .A1(n9963), .A2(n9961), .ZN(P3_U3241) );
  INV_X1 U12479 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n9962) );
  NOR2_X1 U12480 ( .A1(n9963), .A2(n9962), .ZN(P3_U3253) );
  INV_X1 U12481 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n10349) );
  NAND2_X1 U12482 ( .A1(n15257), .A2(P3_U3897), .ZN(n9964) );
  OAI21_X1 U12483 ( .B1(P3_U3897), .B2(n10349), .A(n9964), .ZN(P3_U3491) );
  INV_X1 U12484 ( .A(n10586), .ZN(n10591) );
  OAI222_X1 U12485 ( .A1(n14225), .A2(n9967), .B1(n10591), .B2(P1_U3086), .C1(
        n9965), .C2(n14216), .ZN(P1_U3345) );
  INV_X1 U12486 ( .A(n14911), .ZN(n9968) );
  OAI222_X1 U12487 ( .A1(P2_U3088), .A2(n9968), .B1(n13708), .B2(n9967), .C1(
        n9966), .C2(n13705), .ZN(P2_U3317) );
  MUX2_X1 U12488 ( .A(n9970), .B(P1_REG1_REG_2__SCAN_IN), .S(n10139), .Z(
        n10136) );
  AND2_X1 U12489 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n13863) );
  OAI21_X1 U12490 ( .B1(n13868), .B2(n9969), .A(n13862), .ZN(n10135) );
  NAND2_X1 U12491 ( .A1(n10136), .A2(n10135), .ZN(n10134) );
  OR2_X1 U12492 ( .A1(n10139), .A2(n9970), .ZN(n9971) );
  NAND2_X1 U12493 ( .A1(n10134), .A2(n9971), .ZN(n13876) );
  MUX2_X1 U12494 ( .A(n9972), .B(P1_REG1_REG_3__SCAN_IN), .S(n13878), .Z(
        n13877) );
  OR2_X1 U12495 ( .A1(n13878), .A2(n9972), .ZN(n14629) );
  INV_X1 U12496 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n14801) );
  MUX2_X1 U12497 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n14801), .S(n14620), .Z(
        n14627) );
  MUX2_X1 U12498 ( .A(n9973), .B(P1_REG1_REG_5__SCAN_IN), .S(n10014), .Z(
        n10003) );
  NAND2_X1 U12499 ( .A1(n10004), .A2(n10003), .ZN(n10002) );
  OAI21_X1 U12500 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n9989), .A(n10002), .ZN(
        n10016) );
  XNOR2_X1 U12501 ( .A(n9990), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n10017) );
  NOR2_X1 U12502 ( .A1(n10016), .A2(n10017), .ZN(n10015) );
  INV_X1 U12503 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9974) );
  MUX2_X1 U12504 ( .A(n9974), .B(P1_REG1_REG_7__SCAN_IN), .S(n10036), .Z(n9978) );
  NAND2_X1 U12505 ( .A1(n9976), .A2(n9975), .ZN(n14618) );
  AOI211_X1 U12506 ( .C1(n9979), .C2(n9978), .A(n13911), .B(n10035), .ZN(
        n10001) );
  OR2_X1 U12507 ( .A1(n12062), .A2(n6538), .ZN(n9980) );
  MUX2_X1 U12508 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n9981), .S(n14620), .Z(n9987) );
  INV_X1 U12509 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10909) );
  MUX2_X1 U12510 ( .A(n10909), .B(P1_REG2_REG_2__SCAN_IN), .S(n10139), .Z(
        n10138) );
  INV_X1 U12511 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9983) );
  MUX2_X1 U12512 ( .A(n9983), .B(P1_REG2_REG_1__SCAN_IN), .S(n13868), .Z(
        n13867) );
  AND2_X1 U12513 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9982) );
  NAND2_X1 U12514 ( .A1(n13867), .A2(n9982), .ZN(n13866) );
  OAI21_X1 U12515 ( .B1(n9983), .B2(n13868), .A(n13866), .ZN(n10137) );
  NAND2_X1 U12516 ( .A1(n10138), .A2(n10137), .ZN(n13881) );
  OR2_X1 U12517 ( .A1(n10139), .A2(n10909), .ZN(n13880) );
  NAND2_X1 U12518 ( .A1(n13881), .A2(n13880), .ZN(n9985) );
  MUX2_X1 U12519 ( .A(n14720), .B(P1_REG2_REG_3__SCAN_IN), .S(n13878), .Z(
        n9984) );
  NAND2_X1 U12520 ( .A1(n9985), .A2(n9984), .ZN(n14622) );
  OR2_X1 U12521 ( .A1(n13878), .A2(n14720), .ZN(n14621) );
  NAND2_X1 U12522 ( .A1(n14622), .A2(n14621), .ZN(n9986) );
  AND2_X1 U12523 ( .A1(n9987), .A2(n9986), .ZN(n14619) );
  NOR2_X1 U12524 ( .A1(n6884), .A2(n9981), .ZN(n10006) );
  MUX2_X1 U12525 ( .A(n9988), .B(P1_REG2_REG_5__SCAN_IN), .S(n10014), .Z(
        n10005) );
  OAI21_X1 U12526 ( .B1(n14619), .B2(n10006), .A(n10005), .ZN(n10020) );
  NAND2_X1 U12527 ( .A1(n9989), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10019) );
  MUX2_X1 U12528 ( .A(n11007), .B(P1_REG2_REG_6__SCAN_IN), .S(n9990), .Z(
        n10018) );
  AOI21_X1 U12529 ( .B1(n10020), .B2(n10019), .A(n10018), .ZN(n10022) );
  NOR2_X1 U12530 ( .A1(n10027), .A2(n11007), .ZN(n9993) );
  MUX2_X1 U12531 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n9991), .S(n10036), .Z(n9992) );
  OAI21_X1 U12532 ( .B1(n10022), .B2(n9993), .A(n9992), .ZN(n10033) );
  INV_X1 U12533 ( .A(n10033), .ZN(n9995) );
  NOR3_X1 U12534 ( .A1(n10022), .A2(n9993), .A3(n9992), .ZN(n9994) );
  NOR3_X1 U12535 ( .A1(n13899), .A2(n9995), .A3(n9994), .ZN(n10000) );
  AND2_X1 U12536 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10828) );
  AOI21_X1 U12537 ( .B1(n14615), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n10828), .ZN(
        n9997) );
  OAI21_X1 U12538 ( .B1(n14634), .B2(n9998), .A(n9997), .ZN(n9999) );
  OR3_X1 U12539 ( .A1(n10001), .A2(n10000), .A3(n9999), .ZN(P1_U3250) );
  OAI21_X1 U12540 ( .B1(n10004), .B2(n10003), .A(n10002), .ZN(n10010) );
  INV_X1 U12541 ( .A(n10020), .ZN(n10008) );
  NOR3_X1 U12542 ( .A1(n14619), .A2(n10006), .A3(n10005), .ZN(n10007) );
  NOR3_X1 U12543 ( .A1(n13899), .A2(n10008), .A3(n10007), .ZN(n10009) );
  AOI21_X1 U12544 ( .B1(n14648), .B2(n10010), .A(n10009), .ZN(n10013) );
  NAND2_X1 U12545 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n10871) );
  INV_X1 U12546 ( .A(n10871), .ZN(n10011) );
  AOI21_X1 U12547 ( .B1(n14615), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10011), .ZN(
        n10012) );
  OAI211_X1 U12548 ( .C1(n10014), .C2(n14634), .A(n10013), .B(n10012), .ZN(
        P1_U3248) );
  AOI211_X1 U12549 ( .C1(n10017), .C2(n10016), .A(n10015), .B(n13911), .ZN(
        n10024) );
  AND3_X1 U12550 ( .A1(n10020), .A2(n10019), .A3(n10018), .ZN(n10021) );
  NOR3_X1 U12551 ( .A1(n13899), .A2(n10022), .A3(n10021), .ZN(n10023) );
  NOR2_X1 U12552 ( .A1(n10024), .A2(n10023), .ZN(n10026) );
  NOR2_X1 U12553 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7723), .ZN(n10701) );
  AOI21_X1 U12554 ( .B1(n14615), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10701), .ZN(
        n10025) );
  OAI211_X1 U12555 ( .C1(n10027), .C2(n14634), .A(n10026), .B(n10025), .ZN(
        P1_U3249) );
  MUX2_X1 U12556 ( .A(n10735), .B(n11772), .S(P1_U4016), .Z(n10028) );
  INV_X1 U12557 ( .A(n10028), .ZN(P1_U3574) );
  OAI222_X1 U12558 ( .A1(n13021), .A2(n10030), .B1(n13023), .B2(n10029), .C1(
        n14389), .C2(P3_U3151), .ZN(P3_U3280) );
  NAND2_X1 U12559 ( .A1(n10036), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10032) );
  INV_X1 U12560 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n11206) );
  MUX2_X1 U12561 ( .A(n11206), .B(P1_REG2_REG_8__SCAN_IN), .S(n10198), .Z(
        n10031) );
  AOI21_X1 U12562 ( .B1(n10033), .B2(n10032), .A(n10031), .ZN(n10205) );
  NAND3_X1 U12563 ( .A1(n10033), .A2(n10032), .A3(n10031), .ZN(n10034) );
  NAND2_X1 U12564 ( .A1(n14649), .A2(n10034), .ZN(n10044) );
  MUX2_X1 U12565 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10037), .S(n10198), .Z(
        n10038) );
  OAI21_X1 U12566 ( .B1(n10039), .B2(n10038), .A(n10197), .ZN(n10040) );
  NAND2_X1 U12567 ( .A1(n10040), .A2(n14648), .ZN(n10043) );
  AND2_X1 U12568 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n10993) );
  NOR2_X1 U12569 ( .A1(n14634), .A2(n10201), .ZN(n10041) );
  AOI211_X1 U12570 ( .C1(n14615), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n10993), .B(
        n10041), .ZN(n10042) );
  OAI211_X1 U12571 ( .C1(n10205), .C2(n10044), .A(n10043), .B(n10042), .ZN(
        P1_U3251) );
  INV_X1 U12572 ( .A(n10849), .ZN(n10853) );
  INV_X1 U12573 ( .A(n10045), .ZN(n10055) );
  OAI222_X1 U12574 ( .A1(n10853), .A2(P2_U3088), .B1(n13708), .B2(n10055), 
        .C1(n10046), .C2(n13705), .ZN(P2_U3316) );
  INV_X1 U12575 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10052) );
  OR2_X1 U12576 ( .A1(n13861), .A2(n7639), .ZN(n10047) );
  NAND2_X1 U12577 ( .A1(n10150), .A2(n10047), .ZN(n12274) );
  INV_X1 U12578 ( .A(n12274), .ZN(n10882) );
  OAI21_X1 U12579 ( .B1(n14716), .B2(n14797), .A(n10882), .ZN(n10050) );
  NOR2_X1 U12580 ( .A1(n10154), .A2(n10048), .ZN(n10049) );
  AOI21_X1 U12581 ( .B1(n13860), .B2(n14498), .A(n10049), .ZN(n10885) );
  NAND2_X1 U12582 ( .A1(n10050), .A2(n10885), .ZN(n14196) );
  NAND2_X1 U12583 ( .A1(n14196), .A2(n14799), .ZN(n10051) );
  OAI21_X1 U12584 ( .B1(n14799), .B2(n10052), .A(n10051), .ZN(P1_U3459) );
  INV_X1 U12585 ( .A(n14399), .ZN(n12613) );
  OAI222_X1 U12586 ( .A1(n13021), .A2(n10054), .B1(n12613), .B2(P3_U3151), 
        .C1(n10053), .C2(n11761), .ZN(P3_U3279) );
  INV_X1 U12587 ( .A(n10833), .ZN(n10838) );
  OAI222_X1 U12588 ( .A1(n14216), .A2(n10056), .B1(P1_U3086), .B2(n10838), 
        .C1(n14225), .C2(n10055), .ZN(P1_U3344) );
  INV_X1 U12589 ( .A(n10057), .ZN(n10059) );
  NAND3_X1 U12590 ( .A1(n10060), .A2(n10059), .A3(n10058), .ZN(n10074) );
  NAND2_X1 U12591 ( .A1(n10074), .A2(n10061), .ZN(n10698) );
  INV_X1 U12592 ( .A(n13794), .ZN(n13817) );
  NOR2_X1 U12593 ( .A1(n13836), .A2(n14694), .ZN(n13789) );
  NAND2_X1 U12594 ( .A1(n10698), .A2(n10062), .ZN(n10387) );
  AOI22_X1 U12595 ( .A1(n13789), .A2(n13860), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n10387), .ZN(n10076) );
  INV_X1 U12596 ( .A(n10660), .ZN(n10063) );
  NAND2_X1 U12597 ( .A1(n13861), .A2(n6537), .ZN(n10067) );
  INV_X1 U12598 ( .A(n10064), .ZN(n10065) );
  AOI22_X1 U12599 ( .A1(n7639), .A2(n10664), .B1(n10065), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n10066) );
  NAND2_X1 U12600 ( .A1(n13861), .A2(n10664), .ZN(n10070) );
  OAI22_X1 U12601 ( .A1(n10154), .A2(n6471), .B1(n10064), .B2(n14608), .ZN(
        n10068) );
  INV_X1 U12602 ( .A(n10068), .ZN(n10069) );
  OAI21_X1 U12603 ( .B1(n10071), .B2(n10172), .A(n10173), .ZN(n10130) );
  NAND3_X1 U12604 ( .A1(n10072), .A2(n14781), .A3(n12264), .ZN(n10073) );
  NAND2_X1 U12605 ( .A1(n10130), .A2(n14488), .ZN(n10075) );
  OAI211_X1 U12606 ( .C1(n13817), .C2(n10154), .A(n10076), .B(n10075), .ZN(
        P1_U3232) );
  INV_X1 U12607 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n10343) );
  NAND2_X1 U12608 ( .A1(n7302), .A2(P3_U3897), .ZN(n10077) );
  OAI21_X1 U12609 ( .B1(P3_U3897), .B2(n10343), .A(n10077), .ZN(P3_U3506) );
  INV_X1 U12610 ( .A(n14868), .ZN(n10083) );
  MUX2_X1 U12611 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n10078), .S(n10097), .Z(
        n14838) );
  NAND2_X1 U12612 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n14839) );
  OAI22_X1 U12613 ( .A1(n14838), .A2(n14839), .B1(n10078), .B2(n10097), .ZN(
        n14850) );
  NAND2_X1 U12614 ( .A1(n14851), .A2(n14850), .ZN(n14849) );
  OR2_X1 U12615 ( .A1(n14853), .A2(n10079), .ZN(n10080) );
  NAND2_X1 U12616 ( .A1(n14849), .A2(n10080), .ZN(n13217) );
  MUX2_X1 U12617 ( .A(n10081), .B(P2_REG1_REG_3__SCAN_IN), .S(n10100), .Z(
        n13218) );
  NAND2_X1 U12618 ( .A1(n13217), .A2(n13218), .ZN(n13216) );
  OR2_X1 U12619 ( .A1(n10100), .A2(n10081), .ZN(n10082) );
  NAND2_X1 U12620 ( .A1(n13216), .A2(n10082), .ZN(n14864) );
  INV_X1 U12621 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10547) );
  MUX2_X1 U12622 ( .A(n10547), .B(P2_REG1_REG_4__SCAN_IN), .S(n14868), .Z(
        n14865) );
  INV_X1 U12623 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10084) );
  MUX2_X1 U12624 ( .A(n10084), .B(P2_REG1_REG_5__SCAN_IN), .S(n10102), .Z(
        n10119) );
  XNOR2_X1 U12625 ( .A(n14883), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n14879) );
  NOR2_X1 U12626 ( .A1(n14880), .A2(n14879), .ZN(n14878) );
  AOI21_X1 U12627 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n14883), .A(n14878), .ZN(
        n11917) );
  MUX2_X1 U12628 ( .A(n10085), .B(P2_REG1_REG_7__SCAN_IN), .S(n10103), .Z(
        n11916) );
  NOR2_X1 U12629 ( .A1(n11917), .A2(n11916), .ZN(n11915) );
  MUX2_X1 U12630 ( .A(n10086), .B(P2_REG1_REG_8__SCAN_IN), .S(n10105), .Z(
        n14891) );
  MUX2_X1 U12631 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10087), .S(n10744), .Z(
        n10088) );
  OAI21_X1 U12632 ( .B1(n10089), .B2(n10088), .A(n10743), .ZN(n10096) );
  NAND2_X1 U12633 ( .A1(n10411), .A2(n10090), .ZN(n10092) );
  NAND2_X1 U12634 ( .A1(n10092), .A2(n10091), .ZN(n10093) );
  NAND2_X1 U12635 ( .A1(n10094), .A2(n10093), .ZN(n10111) );
  OR2_X1 U12636 ( .A1(n9530), .A2(P2_U3088), .ZN(n13696) );
  INV_X1 U12637 ( .A(n13696), .ZN(n10095) );
  AND2_X1 U12638 ( .A1(n10111), .A2(n10095), .ZN(n10109) );
  NAND2_X1 U12639 ( .A1(n10096), .A2(n14863), .ZN(n10117) );
  INV_X1 U12640 ( .A(n10100), .ZN(n13214) );
  INV_X1 U12641 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10101) );
  MUX2_X1 U12642 ( .A(n11135), .B(P2_REG2_REG_1__SCAN_IN), .S(n10097), .Z(
        n14844) );
  NAND3_X1 U12643 ( .A1(n14844), .A2(P2_IR_REG_0__SCAN_IN), .A3(
        P2_REG2_REG_0__SCAN_IN), .ZN(n14843) );
  OAI21_X1 U12644 ( .B1(n11135), .B2(n10097), .A(n14843), .ZN(n14857) );
  MUX2_X1 U12645 ( .A(n10098), .B(P2_REG2_REG_2__SCAN_IN), .S(n14853), .Z(
        n14856) );
  NAND2_X1 U12646 ( .A1(n14857), .A2(n14856), .ZN(n14855) );
  INV_X1 U12647 ( .A(n14853), .ZN(n10099) );
  NAND2_X1 U12648 ( .A1(n10099), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n13210) );
  MUX2_X1 U12649 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10101), .S(n10100), .Z(
        n13209) );
  AOI21_X1 U12650 ( .B1(n14855), .B2(n13210), .A(n13209), .ZN(n13212) );
  AOI21_X1 U12651 ( .B1(n13214), .B2(P2_REG2_REG_3__SCAN_IN), .A(n13212), .ZN(
        n14872) );
  MUX2_X1 U12652 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n11094), .S(n14868), .Z(
        n14871) );
  NOR2_X1 U12653 ( .A1(n14872), .A2(n14871), .ZN(n14870) );
  NOR2_X1 U12654 ( .A1(n14868), .A2(n11094), .ZN(n10124) );
  MUX2_X1 U12655 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11125), .S(n10102), .Z(
        n10123) );
  OAI21_X1 U12656 ( .B1(n14870), .B2(n10124), .A(n10123), .ZN(n10126) );
  OAI21_X1 U12657 ( .B1(n11125), .B2(n10129), .A(n10126), .ZN(n14886) );
  INV_X1 U12658 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11286) );
  MUX2_X1 U12659 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11286), .S(n14883), .Z(
        n14885) );
  NAND2_X1 U12660 ( .A1(n14886), .A2(n14885), .ZN(n14884) );
  NAND2_X1 U12661 ( .A1(n14883), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n11922) );
  MUX2_X1 U12662 ( .A(n11301), .B(P2_REG2_REG_7__SCAN_IN), .S(n10103), .Z(
        n11921) );
  AOI21_X1 U12663 ( .B1(n14884), .B2(n11922), .A(n11921), .ZN(n11920) );
  AOI21_X1 U12664 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n10103), .A(n11920), .ZN(
        n14900) );
  INV_X1 U12665 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10104) );
  MUX2_X1 U12666 ( .A(n10104), .B(P2_REG2_REG_8__SCAN_IN), .S(n10105), .Z(
        n14899) );
  NOR2_X1 U12667 ( .A1(n14900), .A2(n14899), .ZN(n14898) );
  AOI21_X1 U12668 ( .B1(n10105), .B2(P2_REG2_REG_8__SCAN_IN), .A(n14898), .ZN(
        n10108) );
  INV_X1 U12669 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10106) );
  MUX2_X1 U12670 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n10106), .S(n10744), .Z(
        n10107) );
  NAND2_X1 U12671 ( .A1(n10108), .A2(n10107), .ZN(n10737) );
  OAI21_X1 U12672 ( .B1(n10108), .B2(n10107), .A(n10737), .ZN(n10115) );
  INV_X1 U12673 ( .A(n10109), .ZN(n10110) );
  OR2_X1 U12674 ( .A1(n10110), .A2(n13701), .ZN(n14913) );
  INV_X1 U12675 ( .A(n14913), .ZN(n14941) );
  NAND2_X1 U12676 ( .A1(n10111), .A2(n9530), .ZN(n14895) );
  INV_X1 U12677 ( .A(n14946), .ZN(n14924) );
  NAND2_X1 U12678 ( .A1(n14924), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n10112) );
  NAND2_X1 U12679 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n11252) );
  OAI211_X1 U12680 ( .C1(n14930), .C2(n10113), .A(n10112), .B(n11252), .ZN(
        n10114) );
  AOI21_X1 U12681 ( .B1(n10115), .B2(n14941), .A(n10114), .ZN(n10116) );
  NAND2_X1 U12682 ( .A1(n10117), .A2(n10116), .ZN(P2_U3223) );
  AND2_X1 U12683 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10122) );
  AOI211_X1 U12684 ( .C1(n10120), .C2(n10119), .A(n10118), .B(n14932), .ZN(
        n10121) );
  AOI211_X1 U12685 ( .C1(n14924), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n10122), .B(
        n10121), .ZN(n10128) );
  OR3_X1 U12686 ( .A1(n14870), .A2(n10124), .A3(n10123), .ZN(n10125) );
  NAND3_X1 U12687 ( .A1(n14941), .A2(n10126), .A3(n10125), .ZN(n10127) );
  OAI211_X1 U12688 ( .C1(n14930), .C2(n10129), .A(n10128), .B(n10127), .ZN(
        P2_U3219) );
  NAND2_X1 U12689 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13865) );
  MUX2_X1 U12690 ( .A(n13865), .B(n10130), .S(n6538), .Z(n10131) );
  NOR2_X1 U12691 ( .A1(n10131), .A2(n12062), .ZN(n10133) );
  NOR2_X1 U12692 ( .A1(n6538), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10132) );
  NOR2_X1 U12693 ( .A1(n12062), .A2(n10132), .ZN(n14610) );
  NOR2_X1 U12694 ( .A1(n14610), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n14607) );
  NOR3_X1 U12695 ( .A1(n10133), .A2(n14607), .A3(n13849), .ZN(n14636) );
  OAI211_X1 U12696 ( .C1(n10136), .C2(n10135), .A(n14648), .B(n10134), .ZN(
        n10144) );
  OAI211_X1 U12697 ( .C1(n10138), .C2(n10137), .A(n14649), .B(n13881), .ZN(
        n10143) );
  AOI22_X1 U12698 ( .A1(n14615), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n10142) );
  INV_X1 U12699 ( .A(n14634), .ZN(n14645) );
  INV_X1 U12700 ( .A(n10139), .ZN(n10140) );
  NAND2_X1 U12701 ( .A1(n14645), .A2(n10140), .ZN(n10141) );
  NAND4_X1 U12702 ( .A1(n10144), .A2(n10143), .A3(n10142), .A4(n10141), .ZN(
        n10145) );
  OR2_X1 U12703 ( .A1(n14636), .A2(n10145), .ZN(P1_U3245) );
  INV_X1 U12704 ( .A(n14416), .ZN(n12666) );
  INV_X1 U12705 ( .A(n10146), .ZN(n10148) );
  INV_X1 U12706 ( .A(SI_17_), .ZN(n10147) );
  OAI222_X1 U12707 ( .A1(n12666), .A2(P3_U3151), .B1(n13021), .B2(n10148), 
        .C1(n10147), .C2(n11761), .ZN(P3_U3278) );
  INV_X1 U12708 ( .A(n10150), .ZN(n10151) );
  NAND2_X1 U12709 ( .A1(n12275), .A2(n10151), .ZN(n10152) );
  NAND2_X1 U12710 ( .A1(n10153), .A2(n10152), .ZN(n10158) );
  INV_X1 U12711 ( .A(n10158), .ZN(n11906) );
  INV_X1 U12712 ( .A(n14716), .ZN(n14691) );
  INV_X1 U12713 ( .A(n13860), .ZN(n10156) );
  OR2_X1 U12714 ( .A1(n11902), .A2(n10154), .ZN(n10155) );
  NAND2_X1 U12715 ( .A1(n10191), .A2(n10155), .ZN(n10162) );
  XNOR2_X1 U12716 ( .A(n10156), .B(n10162), .ZN(n10157) );
  MUX2_X1 U12717 ( .A(n10157), .B(n12275), .S(n13861), .Z(n10161) );
  INV_X1 U12718 ( .A(n14660), .ZN(n14718) );
  NAND2_X1 U12719 ( .A1(n10158), .A2(n14718), .ZN(n10160) );
  AOI22_X1 U12720 ( .A1(n14596), .A2(n13861), .B1(n12090), .B2(n14498), .ZN(
        n10159) );
  OAI211_X1 U12721 ( .C1(n14691), .C2(n10161), .A(n10160), .B(n10159), .ZN(
        n11899) );
  INV_X1 U12722 ( .A(n11899), .ZN(n10164) );
  INV_X1 U12723 ( .A(n10162), .ZN(n11900) );
  AOI22_X1 U12724 ( .A1(n11900), .A2(n14726), .B1(n10177), .B2(n14761), .ZN(
        n10163) );
  OAI211_X1 U12725 ( .C1(n11906), .C2(n14766), .A(n10164), .B(n10163), .ZN(
        n10166) );
  NAND2_X1 U12726 ( .A1(n10166), .A2(n14811), .ZN(n10165) );
  OAI21_X1 U12727 ( .B1(n14811), .B2(n9969), .A(n10165), .ZN(P1_U3529) );
  NAND2_X1 U12728 ( .A1(n10166), .A2(n14799), .ZN(n10167) );
  OAI21_X1 U12729 ( .B1(n14799), .B2(n7616), .A(n10167), .ZN(P1_U3462) );
  CLKBUF_X2 U12730 ( .A(P2_U3947), .Z(n13208) );
  NAND2_X1 U12731 ( .A1(n11566), .A2(n13208), .ZN(n10168) );
  OAI21_X1 U12732 ( .B1(n8403), .B2(n13208), .A(n10168), .ZN(P2_U3544) );
  NAND2_X1 U12733 ( .A1(n13860), .A2(n10664), .ZN(n10170) );
  NAND2_X1 U12734 ( .A1(n10170), .A2(n10169), .ZN(n10171) );
  XNOR2_X1 U12735 ( .A(n10171), .B(n12332), .ZN(n10379) );
  AOI22_X1 U12736 ( .A1(n13860), .A2(n6536), .B1(n10177), .B2(n10664), .ZN(
        n10380) );
  XNOR2_X1 U12737 ( .A(n10379), .B(n10380), .ZN(n10378) );
  XOR2_X1 U12738 ( .A(n10378), .B(n10377), .Z(n10179) );
  NOR2_X1 U12739 ( .A1(n13836), .A2(n14696), .ZN(n13814) );
  INV_X1 U12740 ( .A(n13814), .ZN(n13763) );
  AOI22_X1 U12741 ( .A1(n13789), .A2(n12090), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n10387), .ZN(n10175) );
  OAI21_X1 U12742 ( .B1(n7640), .B2(n13763), .A(n10175), .ZN(n10176) );
  AOI21_X1 U12743 ( .B1(n13794), .B2(n10177), .A(n10176), .ZN(n10178) );
  OAI21_X1 U12744 ( .B1(n14593), .B2(n10179), .A(n10178), .ZN(P1_U3222) );
  INV_X1 U12745 ( .A(n11102), .ZN(n11106) );
  INV_X1 U12746 ( .A(n10180), .ZN(n10375) );
  OAI222_X1 U12747 ( .A1(P2_U3088), .A2(n11106), .B1(n13708), .B2(n10375), 
        .C1(n10181), .C2(n13705), .ZN(P2_U3315) );
  OAI21_X1 U12748 ( .B1(n10184), .B2(n10183), .A(n10182), .ZN(n10189) );
  INV_X1 U12749 ( .A(n10189), .ZN(n10915) );
  XNOR2_X1 U12750 ( .A(n12273), .B(n10185), .ZN(n10187) );
  INV_X1 U12751 ( .A(n14694), .ZN(n14597) );
  AOI22_X1 U12752 ( .A1(n14596), .A2(n13860), .B1(n13859), .B2(n14597), .ZN(
        n10186) );
  OAI21_X1 U12753 ( .B1(n10187), .B2(n14691), .A(n10186), .ZN(n10188) );
  AOI21_X1 U12754 ( .B1(n10189), .B2(n14718), .A(n10188), .ZN(n10908) );
  INV_X1 U12755 ( .A(n14725), .ZN(n10190) );
  AOI211_X1 U12756 ( .C1(n12089), .C2(n10191), .A(n14792), .B(n10190), .ZN(
        n10912) );
  AOI21_X1 U12757 ( .B1(n12089), .B2(n14761), .A(n10912), .ZN(n10192) );
  OAI211_X1 U12758 ( .C1(n10915), .C2(n14766), .A(n10908), .B(n10192), .ZN(
        n10194) );
  NAND2_X1 U12759 ( .A1(n10194), .A2(n14811), .ZN(n10193) );
  OAI21_X1 U12760 ( .B1(n14811), .B2(n9970), .A(n10193), .ZN(P1_U3530) );
  NAND2_X1 U12761 ( .A1(n10194), .A2(n14799), .ZN(n10195) );
  OAI21_X1 U12762 ( .B1(n14799), .B2(n7641), .A(n10195), .ZN(P1_U3465) );
  MUX2_X1 U12763 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10196), .S(n10518), .Z(
        n10200) );
  OAI21_X1 U12764 ( .B1(n10198), .B2(P1_REG1_REG_8__SCAN_IN), .A(n10197), .ZN(
        n10199) );
  NAND2_X1 U12765 ( .A1(n10199), .A2(n10200), .ZN(n10515) );
  OAI21_X1 U12766 ( .B1(n10200), .B2(n10199), .A(n10515), .ZN(n10211) );
  NOR2_X1 U12767 ( .A1(n10201), .A2(n11206), .ZN(n10204) );
  MUX2_X1 U12768 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10202), .S(n10518), .Z(
        n10203) );
  OAI21_X1 U12769 ( .B1(n10205), .B2(n10204), .A(n10203), .ZN(n10521) );
  INV_X1 U12770 ( .A(n10521), .ZN(n10207) );
  NOR3_X1 U12771 ( .A1(n10205), .A2(n10204), .A3(n10203), .ZN(n10206) );
  NOR3_X1 U12772 ( .A1(n10207), .A2(n10206), .A3(n13899), .ZN(n10210) );
  INV_X1 U12773 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14251) );
  INV_X1 U12774 ( .A(n14615), .ZN(n14653) );
  NAND2_X1 U12775 ( .A1(n14645), .A2(n10518), .ZN(n10208) );
  NAND2_X1 U12776 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n11446) );
  OAI211_X1 U12777 ( .C1(n14251), .C2(n14653), .A(n10208), .B(n11446), .ZN(
        n10209) );
  AOI211_X1 U12778 ( .C1(n10211), .C2(n14648), .A(n10210), .B(n10209), .ZN(
        n10374) );
  INV_X1 U12779 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14362) );
  AOI22_X1 U12780 ( .A1(n14362), .A2(keyinput85), .B1(n9137), .B2(keyinput112), 
        .ZN(n10212) );
  OAI221_X1 U12781 ( .B1(n14362), .B2(keyinput85), .C1(n9137), .C2(keyinput112), .A(n10212), .ZN(n10219) );
  INV_X1 U12782 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n14737) );
  AOI22_X1 U12783 ( .A1(n7875), .A2(keyinput123), .B1(n14737), .B2(keyinput106), .ZN(n10213) );
  OAI221_X1 U12784 ( .B1(n7875), .B2(keyinput123), .C1(n14737), .C2(
        keyinput106), .A(n10213), .ZN(n10218) );
  INV_X1 U12785 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n11436) );
  AOI22_X1 U12786 ( .A1(n14232), .A2(keyinput83), .B1(keyinput93), .B2(n11436), 
        .ZN(n10214) );
  OAI221_X1 U12787 ( .B1(n14232), .B2(keyinput83), .C1(n11436), .C2(keyinput93), .A(n10214), .ZN(n10217) );
  INV_X1 U12788 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14324) );
  INV_X1 U12789 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n14949) );
  AOI22_X1 U12790 ( .A1(n14324), .A2(keyinput120), .B1(n14949), .B2(keyinput99), .ZN(n10215) );
  OAI221_X1 U12791 ( .B1(n14324), .B2(keyinput120), .C1(n14949), .C2(
        keyinput99), .A(n10215), .ZN(n10216) );
  NOR4_X1 U12792 ( .A1(n10219), .A2(n10218), .A3(n10217), .A4(n10216), .ZN(
        n10250) );
  AOI22_X1 U12793 ( .A1(n13296), .A2(keyinput64), .B1(keyinput72), .B2(n13652), 
        .ZN(n10220) );
  OAI221_X1 U12794 ( .B1(n13296), .B2(keyinput64), .C1(n13652), .C2(keyinput72), .A(n10220), .ZN(n10228) );
  INV_X1 U12795 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n14948) );
  AOI22_X1 U12796 ( .A1(P3_REG2_REG_21__SCAN_IN), .A2(keyinput95), .B1(n14948), 
        .B2(keyinput78), .ZN(n10221) );
  OAI221_X1 U12797 ( .B1(P3_REG2_REG_21__SCAN_IN), .B2(keyinput95), .C1(n14948), .C2(keyinput78), .A(n10221), .ZN(n10227) );
  AOI22_X1 U12798 ( .A1(n13022), .A2(keyinput96), .B1(keyinput105), .B2(n10223), .ZN(n10222) );
  OAI221_X1 U12799 ( .B1(n13022), .B2(keyinput96), .C1(n10223), .C2(
        keyinput105), .A(n10222), .ZN(n10226) );
  INV_X1 U12800 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n12475) );
  AOI22_X1 U12801 ( .A1(n11286), .A2(keyinput91), .B1(n12475), .B2(keyinput116), .ZN(n10224) );
  OAI221_X1 U12802 ( .B1(n11286), .B2(keyinput91), .C1(n12475), .C2(
        keyinput116), .A(n10224), .ZN(n10225) );
  NOR4_X1 U12803 ( .A1(n10228), .A2(n10227), .A3(n10226), .A4(n10225), .ZN(
        n10249) );
  INV_X1 U12804 ( .A(SI_24_), .ZN(n11548) );
  AOI22_X1 U12805 ( .A1(n11548), .A2(keyinput109), .B1(keyinput110), .B2(
        n10910), .ZN(n10229) );
  OAI221_X1 U12806 ( .B1(n11548), .B2(keyinput109), .C1(n10910), .C2(
        keyinput110), .A(n10229), .ZN(n10237) );
  AOI22_X1 U12807 ( .A1(n13686), .A2(keyinput66), .B1(keyinput104), .B2(n7641), 
        .ZN(n10230) );
  OAI221_X1 U12808 ( .B1(n13686), .B2(keyinput66), .C1(n7641), .C2(keyinput104), .A(n10230), .ZN(n10236) );
  INV_X1 U12809 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14876) );
  AOI22_X1 U12810 ( .A1(n14876), .A2(keyinput68), .B1(n9182), .B2(keyinput101), 
        .ZN(n10231) );
  OAI221_X1 U12811 ( .B1(n14876), .B2(keyinput68), .C1(n9182), .C2(keyinput101), .A(n10231), .ZN(n10235) );
  XNOR2_X1 U12812 ( .A(P3_IR_REG_4__SCAN_IN), .B(keyinput117), .ZN(n10233) );
  XNOR2_X1 U12813 ( .A(P2_REG0_REG_31__SCAN_IN), .B(keyinput73), .ZN(n10232)
         );
  NAND2_X1 U12814 ( .A1(n10233), .A2(n10232), .ZN(n10234) );
  NOR4_X1 U12815 ( .A1(n10237), .A2(n10236), .A3(n10235), .A4(n10234), .ZN(
        n10248) );
  AOI22_X1 U12816 ( .A1(n11861), .A2(keyinput108), .B1(keyinput80), .B2(n10086), .ZN(n10238) );
  OAI221_X1 U12817 ( .B1(n11861), .B2(keyinput108), .C1(n10086), .C2(
        keyinput80), .A(n10238), .ZN(n10246) );
  AOI22_X1 U12818 ( .A1(n10336), .A2(keyinput81), .B1(keyinput76), .B2(n10343), 
        .ZN(n10239) );
  OAI221_X1 U12819 ( .B1(n10336), .B2(keyinput81), .C1(n10343), .C2(keyinput76), .A(n10239), .ZN(n10245) );
  AOI22_X1 U12820 ( .A1(n9237), .A2(keyinput127), .B1(n13003), .B2(keyinput89), 
        .ZN(n10240) );
  OAI221_X1 U12821 ( .B1(n9237), .B2(keyinput127), .C1(n13003), .C2(keyinput89), .A(n10240), .ZN(n10244) );
  XOR2_X1 U12822 ( .A(n12621), .B(keyinput107), .Z(n10242) );
  XNOR2_X1 U12823 ( .A(P3_IR_REG_12__SCAN_IN), .B(keyinput97), .ZN(n10241) );
  NAND2_X1 U12824 ( .A1(n10242), .A2(n10241), .ZN(n10243) );
  NOR4_X1 U12825 ( .A1(n10246), .A2(n10245), .A3(n10244), .A4(n10243), .ZN(
        n10247) );
  AND4_X1 U12826 ( .A1(n10250), .A2(n10249), .A3(n10248), .A4(n10247), .ZN(
        n10372) );
  OAI22_X1 U12827 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(keyinput102), .B1(
        P3_REG3_REG_18__SCAN_IN), .B2(keyinput114), .ZN(n10251) );
  AOI221_X1 U12828 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(keyinput102), .C1(
        keyinput114), .C2(P3_REG3_REG_18__SCAN_IN), .A(n10251), .ZN(n10258) );
  OAI22_X1 U12829 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput88), .B1(
        keyinput122), .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n10252) );
  AOI221_X1 U12830 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput88), .C1(
        P3_DATAO_REG_26__SCAN_IN), .C2(keyinput122), .A(n10252), .ZN(n10257)
         );
  OAI22_X1 U12831 ( .A1(P3_REG0_REG_4__SCAN_IN), .A2(keyinput79), .B1(
        P1_REG2_REG_21__SCAN_IN), .B2(keyinput111), .ZN(n10253) );
  AOI221_X1 U12832 ( .B1(P3_REG0_REG_4__SCAN_IN), .B2(keyinput79), .C1(
        keyinput111), .C2(P1_REG2_REG_21__SCAN_IN), .A(n10253), .ZN(n10256) );
  OAI22_X1 U12833 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(keyinput75), .B1(
        keyinput115), .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n10254) );
  AOI221_X1 U12834 ( .B1(P1_DATAO_REG_19__SCAN_IN), .B2(keyinput75), .C1(
        P3_DATAO_REG_3__SCAN_IN), .C2(keyinput115), .A(n10254), .ZN(n10255) );
  NAND4_X1 U12835 ( .A1(n10258), .A2(n10257), .A3(n10256), .A4(n10255), .ZN(
        n10286) );
  OAI22_X1 U12836 ( .A1(SI_18_), .A2(keyinput77), .B1(keyinput90), .B2(
        P3_REG2_REG_7__SCAN_IN), .ZN(n10259) );
  AOI221_X1 U12837 ( .B1(SI_18_), .B2(keyinput77), .C1(P3_REG2_REG_7__SCAN_IN), 
        .C2(keyinput90), .A(n10259), .ZN(n10266) );
  OAI22_X1 U12838 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput126), .B1(
        P2_REG1_REG_1__SCAN_IN), .B2(keyinput70), .ZN(n10260) );
  AOI221_X1 U12839 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput126), .C1(
        keyinput70), .C2(P2_REG1_REG_1__SCAN_IN), .A(n10260), .ZN(n10265) );
  OAI22_X1 U12840 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(keyinput69), .B1(
        P2_REG1_REG_25__SCAN_IN), .B2(keyinput87), .ZN(n10261) );
  AOI221_X1 U12841 ( .B1(P3_IR_REG_11__SCAN_IN), .B2(keyinput69), .C1(
        keyinput87), .C2(P2_REG1_REG_25__SCAN_IN), .A(n10261), .ZN(n10264) );
  OAI22_X1 U12842 ( .A1(P3_REG2_REG_9__SCAN_IN), .A2(keyinput121), .B1(
        keyinput113), .B2(P3_B_REG_SCAN_IN), .ZN(n10262) );
  AOI221_X1 U12843 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(keyinput121), .C1(
        P3_B_REG_SCAN_IN), .C2(keyinput113), .A(n10262), .ZN(n10263) );
  NAND4_X1 U12844 ( .A1(n10266), .A2(n10265), .A3(n10264), .A4(n10263), .ZN(
        n10285) );
  OAI22_X1 U12845 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(keyinput67), .B1(
        keyinput71), .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n10267) );
  AOI221_X1 U12846 ( .B1(P2_IR_REG_14__SCAN_IN), .B2(keyinput67), .C1(
        P3_DATAO_REG_0__SCAN_IN), .C2(keyinput71), .A(n10267), .ZN(n10274) );
  OAI22_X1 U12847 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(keyinput125), .B1(
        keyinput100), .B2(P1_ADDR_REG_8__SCAN_IN), .ZN(n10268) );
  AOI221_X1 U12848 ( .B1(P1_REG3_REG_17__SCAN_IN), .B2(keyinput125), .C1(
        P1_ADDR_REG_8__SCAN_IN), .C2(keyinput100), .A(n10268), .ZN(n10273) );
  OAI22_X1 U12849 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput103), .B1(
        P1_REG2_REG_25__SCAN_IN), .B2(keyinput84), .ZN(n10269) );
  AOI221_X1 U12850 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput103), .C1(
        keyinput84), .C2(P1_REG2_REG_25__SCAN_IN), .A(n10269), .ZN(n10272) );
  OAI22_X1 U12851 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput118), .B1(
        P3_ADDR_REG_8__SCAN_IN), .B2(keyinput119), .ZN(n10270) );
  AOI221_X1 U12852 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput118), .C1(
        keyinput119), .C2(P3_ADDR_REG_8__SCAN_IN), .A(n10270), .ZN(n10271) );
  NAND4_X1 U12853 ( .A1(n10274), .A2(n10273), .A3(n10272), .A4(n10271), .ZN(
        n10284) );
  OAI22_X1 U12854 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput74), .B1(
        keyinput98), .B2(P1_REG3_REG_25__SCAN_IN), .ZN(n10275) );
  AOI221_X1 U12855 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput74), .C1(
        P1_REG3_REG_25__SCAN_IN), .C2(keyinput98), .A(n10275), .ZN(n10282) );
  OAI22_X1 U12856 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput82), .B1(
        keyinput92), .B2(P1_REG2_REG_19__SCAN_IN), .ZN(n10276) );
  AOI221_X1 U12857 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput82), .C1(
        P1_REG2_REG_19__SCAN_IN), .C2(keyinput92), .A(n10276), .ZN(n10281) );
  OAI22_X1 U12858 ( .A1(SI_6_), .A2(keyinput124), .B1(keyinput94), .B2(
        P1_IR_REG_3__SCAN_IN), .ZN(n10277) );
  AOI221_X1 U12859 ( .B1(SI_6_), .B2(keyinput124), .C1(P1_IR_REG_3__SCAN_IN), 
        .C2(keyinput94), .A(n10277), .ZN(n10280) );
  OAI22_X1 U12860 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(keyinput65), .B1(
        P1_REG2_REG_8__SCAN_IN), .B2(keyinput86), .ZN(n10278) );
  AOI221_X1 U12861 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(keyinput65), .C1(
        keyinput86), .C2(P1_REG2_REG_8__SCAN_IN), .A(n10278), .ZN(n10279) );
  NAND4_X1 U12862 ( .A1(n10282), .A2(n10281), .A3(n10280), .A4(n10279), .ZN(
        n10283) );
  NOR4_X1 U12863 ( .A1(n10286), .A2(n10285), .A3(n10284), .A4(n10283), .ZN(
        n10371) );
  AOI22_X1 U12864 ( .A1(P2_REG2_REG_28__SCAN_IN), .A2(keyinput0), .B1(
        P3_IR_REG_12__SCAN_IN), .B2(keyinput33), .ZN(n10287) );
  OAI221_X1 U12865 ( .B1(P2_REG2_REG_28__SCAN_IN), .B2(keyinput0), .C1(
        P3_IR_REG_12__SCAN_IN), .C2(keyinput33), .A(n10287), .ZN(n10294) );
  AOI22_X1 U12866 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(keyinput61), .B1(
        P2_D_REG_5__SCAN_IN), .B2(keyinput35), .ZN(n10288) );
  OAI221_X1 U12867 ( .B1(P1_REG3_REG_17__SCAN_IN), .B2(keyinput61), .C1(
        P2_D_REG_5__SCAN_IN), .C2(keyinput35), .A(n10288), .ZN(n10293) );
  AOI22_X1 U12868 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(keyinput30), .B1(
        P3_REG2_REG_7__SCAN_IN), .B2(keyinput26), .ZN(n10289) );
  OAI221_X1 U12869 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(keyinput30), .C1(
        P3_REG2_REG_7__SCAN_IN), .C2(keyinput26), .A(n10289), .ZN(n10292) );
  AOI22_X1 U12870 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput39), .B1(SI_18_), 
        .B2(keyinput13), .ZN(n10290) );
  OAI221_X1 U12871 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput39), .C1(SI_18_), 
        .C2(keyinput13), .A(n10290), .ZN(n10291) );
  NOR4_X1 U12872 ( .A1(n10294), .A2(n10293), .A3(n10292), .A4(n10291), .ZN(
        n10322) );
  AOI22_X1 U12873 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(keyinput52), .B1(
        P3_IR_REG_4__SCAN_IN), .B2(keyinput53), .ZN(n10295) );
  OAI221_X1 U12874 ( .B1(P3_REG3_REG_16__SCAN_IN), .B2(keyinput52), .C1(
        P3_IR_REG_4__SCAN_IN), .C2(keyinput53), .A(n10295), .ZN(n10302) );
  AOI22_X1 U12875 ( .A1(P3_REG2_REG_9__SCAN_IN), .A2(keyinput57), .B1(
        P3_REG3_REG_24__SCAN_IN), .B2(keyinput38), .ZN(n10296) );
  OAI221_X1 U12876 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(keyinput57), .C1(
        P3_REG3_REG_24__SCAN_IN), .C2(keyinput38), .A(n10296), .ZN(n10301) );
  AOI22_X1 U12877 ( .A1(P1_REG3_REG_2__SCAN_IN), .A2(keyinput46), .B1(
        P3_REG0_REG_15__SCAN_IN), .B2(keyinput25), .ZN(n10297) );
  OAI221_X1 U12878 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(keyinput46), .C1(
        P3_REG0_REG_15__SCAN_IN), .C2(keyinput25), .A(n10297), .ZN(n10300) );
  AOI22_X1 U12879 ( .A1(P3_DATAO_REG_26__SCAN_IN), .A2(keyinput58), .B1(SI_6_), 
        .B2(keyinput60), .ZN(n10298) );
  OAI221_X1 U12880 ( .B1(P3_DATAO_REG_26__SCAN_IN), .B2(keyinput58), .C1(SI_6_), .C2(keyinput60), .A(n10298), .ZN(n10299) );
  NOR4_X1 U12881 ( .A1(n10302), .A2(n10301), .A3(n10300), .A4(n10299), .ZN(
        n10321) );
  AOI22_X1 U12882 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(keyinput36), .B1(
        P3_IR_REG_11__SCAN_IN), .B2(keyinput5), .ZN(n10303) );
  OAI221_X1 U12883 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(keyinput36), .C1(
        P3_IR_REG_11__SCAN_IN), .C2(keyinput5), .A(n10303), .ZN(n10310) );
  AOI22_X1 U12884 ( .A1(P2_REG0_REG_15__SCAN_IN), .A2(keyinput41), .B1(
        P2_IR_REG_14__SCAN_IN), .B2(keyinput3), .ZN(n10304) );
  OAI221_X1 U12885 ( .B1(P2_REG0_REG_15__SCAN_IN), .B2(keyinput41), .C1(
        P2_IR_REG_14__SCAN_IN), .C2(keyinput3), .A(n10304), .ZN(n10309) );
  AOI22_X1 U12886 ( .A1(P1_REG2_REG_19__SCAN_IN), .A2(keyinput28), .B1(
        P3_REG1_REG_8__SCAN_IN), .B2(keyinput43), .ZN(n10305) );
  OAI221_X1 U12887 ( .B1(P1_REG2_REG_19__SCAN_IN), .B2(keyinput28), .C1(
        P3_REG1_REG_8__SCAN_IN), .C2(keyinput43), .A(n10305), .ZN(n10308) );
  AOI22_X1 U12888 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(keyinput37), .B1(
        P3_REG2_REG_21__SCAN_IN), .B2(keyinput31), .ZN(n10306) );
  OAI221_X1 U12889 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(keyinput37), .C1(
        P3_REG2_REG_21__SCAN_IN), .C2(keyinput31), .A(n10306), .ZN(n10307) );
  NOR4_X1 U12890 ( .A1(n10310), .A2(n10309), .A3(n10308), .A4(n10307), .ZN(
        n10320) );
  AOI22_X1 U12891 ( .A1(P3_DATAO_REG_28__SCAN_IN), .A2(keyinput29), .B1(
        P3_ADDR_REG_8__SCAN_IN), .B2(keyinput55), .ZN(n10311) );
  OAI221_X1 U12892 ( .B1(P3_DATAO_REG_28__SCAN_IN), .B2(keyinput29), .C1(
        P3_ADDR_REG_8__SCAN_IN), .C2(keyinput55), .A(n10311), .ZN(n10318) );
  AOI22_X1 U12893 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(keyinput4), .B1(
        P1_REG2_REG_25__SCAN_IN), .B2(keyinput20), .ZN(n10312) );
  OAI221_X1 U12894 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(keyinput4), .C1(
        P1_REG2_REG_25__SCAN_IN), .C2(keyinput20), .A(n10312), .ZN(n10317) );
  AOI22_X1 U12895 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(keyinput59), .B1(
        P3_B_REG_SCAN_IN), .B2(keyinput49), .ZN(n10313) );
  OAI221_X1 U12896 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(keyinput59), .C1(
        P3_B_REG_SCAN_IN), .C2(keyinput49), .A(n10313), .ZN(n10316) );
  AOI22_X1 U12897 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput62), .B1(
        P2_REG3_REG_9__SCAN_IN), .B2(keyinput10), .ZN(n10314) );
  OAI221_X1 U12898 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput62), .C1(
        P2_REG3_REG_9__SCAN_IN), .C2(keyinput10), .A(n10314), .ZN(n10315) );
  NOR4_X1 U12899 ( .A1(n10318), .A2(n10317), .A3(n10316), .A4(n10315), .ZN(
        n10319) );
  NAND4_X1 U12900 ( .A1(n10322), .A2(n10321), .A3(n10320), .A4(n10319), .ZN(
        n10370) );
  AOI22_X1 U12901 ( .A1(n13652), .A2(keyinput8), .B1(n10324), .B2(keyinput24), 
        .ZN(n10323) );
  OAI221_X1 U12902 ( .B1(n13652), .B2(keyinput8), .C1(n10324), .C2(keyinput24), 
        .A(n10323), .ZN(n10331) );
  AOI22_X1 U12903 ( .A1(n11247), .A2(keyinput11), .B1(keyinput27), .B2(n11286), 
        .ZN(n10325) );
  OAI221_X1 U12904 ( .B1(n11247), .B2(keyinput11), .C1(n11286), .C2(keyinput27), .A(n10325), .ZN(n10330) );
  AOI22_X1 U12905 ( .A1(n10086), .A2(keyinput16), .B1(n13686), .B2(keyinput2), 
        .ZN(n10326) );
  OAI221_X1 U12906 ( .B1(n10086), .B2(keyinput16), .C1(n13686), .C2(keyinput2), 
        .A(n10326), .ZN(n10329) );
  AOI22_X1 U12907 ( .A1(n7641), .A2(keyinput40), .B1(n7964), .B2(keyinput47), 
        .ZN(n10327) );
  OAI221_X1 U12908 ( .B1(n7641), .B2(keyinput40), .C1(n7964), .C2(keyinput47), 
        .A(n10327), .ZN(n10328) );
  NOR4_X1 U12909 ( .A1(n10331), .A2(n10330), .A3(n10329), .A4(n10328), .ZN(
        n10368) );
  AOI22_X1 U12910 ( .A1(n14931), .A2(keyinput54), .B1(keyinput9), .B2(n10333), 
        .ZN(n10332) );
  OAI221_X1 U12911 ( .B1(n14931), .B2(keyinput54), .C1(n10333), .C2(keyinput9), 
        .A(n10332), .ZN(n10341) );
  AOI22_X1 U12912 ( .A1(n9237), .A2(keyinput63), .B1(n11861), .B2(keyinput44), 
        .ZN(n10334) );
  OAI221_X1 U12913 ( .B1(n9237), .B2(keyinput63), .C1(n11861), .C2(keyinput44), 
        .A(n10334), .ZN(n10340) );
  AOI22_X1 U12914 ( .A1(n14324), .A2(keyinput56), .B1(n10336), .B2(keyinput17), 
        .ZN(n10335) );
  OAI221_X1 U12915 ( .B1(n14324), .B2(keyinput56), .C1(n10336), .C2(keyinput17), .A(n10335), .ZN(n10339) );
  AOI22_X1 U12916 ( .A1(n11528), .A2(keyinput1), .B1(keyinput42), .B2(n14737), 
        .ZN(n10337) );
  OAI221_X1 U12917 ( .B1(n11528), .B2(keyinput1), .C1(n14737), .C2(keyinput42), 
        .A(n10337), .ZN(n10338) );
  NOR4_X1 U12918 ( .A1(n10341), .A2(n10340), .A3(n10339), .A4(n10338), .ZN(
        n10367) );
  AOI22_X1 U12919 ( .A1(n8233), .A2(keyinput15), .B1(keyinput34), .B2(n13754), 
        .ZN(n10342) );
  OAI221_X1 U12920 ( .B1(n8233), .B2(keyinput15), .C1(n13754), .C2(keyinput34), 
        .A(n10342), .ZN(n10347) );
  XNOR2_X1 U12921 ( .A(n10343), .B(keyinput12), .ZN(n10346) );
  XNOR2_X1 U12922 ( .A(n10344), .B(keyinput18), .ZN(n10345) );
  OR3_X1 U12923 ( .A1(n10347), .A2(n10346), .A3(n10345), .ZN(n10354) );
  AOI22_X1 U12924 ( .A1(n10349), .A2(keyinput7), .B1(n13022), .B2(keyinput32), 
        .ZN(n10348) );
  OAI221_X1 U12925 ( .B1(n10349), .B2(keyinput7), .C1(n13022), .C2(keyinput32), 
        .A(n10348), .ZN(n10353) );
  AOI22_X1 U12926 ( .A1(n14362), .A2(keyinput21), .B1(n10351), .B2(keyinput23), 
        .ZN(n10350) );
  OAI221_X1 U12927 ( .B1(n14362), .B2(keyinput21), .C1(n10351), .C2(keyinput23), .A(n10350), .ZN(n10352) );
  NOR3_X1 U12928 ( .A1(n10354), .A2(n10353), .A3(n10352), .ZN(n10366) );
  AOI22_X1 U12929 ( .A1(n10356), .A2(keyinput51), .B1(n11548), .B2(keyinput45), 
        .ZN(n10355) );
  OAI221_X1 U12930 ( .B1(n10356), .B2(keyinput51), .C1(n11548), .C2(keyinput45), .A(n10355), .ZN(n10364) );
  INV_X1 U12931 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n10358) );
  AOI22_X1 U12932 ( .A1(n10358), .A2(keyinput50), .B1(keyinput22), .B2(n11206), 
        .ZN(n10357) );
  OAI221_X1 U12933 ( .B1(n10358), .B2(keyinput50), .C1(n11206), .C2(keyinput22), .A(n10357), .ZN(n10363) );
  AOI22_X1 U12934 ( .A1(n14232), .A2(keyinput19), .B1(n9137), .B2(keyinput48), 
        .ZN(n10359) );
  OAI221_X1 U12935 ( .B1(n14232), .B2(keyinput19), .C1(n9137), .C2(keyinput48), 
        .A(n10359), .ZN(n10362) );
  AOI22_X1 U12936 ( .A1(n14948), .A2(keyinput14), .B1(keyinput6), .B2(n10078), 
        .ZN(n10360) );
  OAI221_X1 U12937 ( .B1(n14948), .B2(keyinput14), .C1(n10078), .C2(keyinput6), 
        .A(n10360), .ZN(n10361) );
  NOR4_X1 U12938 ( .A1(n10364), .A2(n10363), .A3(n10362), .A4(n10361), .ZN(
        n10365) );
  NAND4_X1 U12939 ( .A1(n10368), .A2(n10367), .A3(n10366), .A4(n10365), .ZN(
        n10369) );
  AOI211_X1 U12940 ( .C1(n10372), .C2(n10371), .A(n10370), .B(n10369), .ZN(
        n10373) );
  XNOR2_X1 U12941 ( .A(n10374), .B(n10373), .ZN(P1_U3252) );
  INV_X1 U12942 ( .A(n11236), .ZN(n10839) );
  OAI222_X1 U12943 ( .A1(n14216), .A2(n10376), .B1(n10839), .B2(P1_U3086), 
        .C1(n14225), .C2(n10375), .ZN(P1_U3343) );
  INV_X1 U12944 ( .A(n10379), .ZN(n10381) );
  NAND2_X1 U12945 ( .A1(n10381), .A2(n10380), .ZN(n10382) );
  NAND2_X1 U12946 ( .A1(n10383), .A2(n10382), .ZN(n10655) );
  NAND2_X1 U12947 ( .A1(n12090), .A2(n10664), .ZN(n10385) );
  OR2_X1 U12948 ( .A1(n12092), .A2(n6471), .ZN(n10384) );
  NAND2_X1 U12949 ( .A1(n10385), .A2(n10384), .ZN(n10386) );
  XNOR2_X1 U12950 ( .A(n10386), .B(n12332), .ZN(n10656) );
  AOI22_X1 U12951 ( .A1(n12090), .A2(n11944), .B1(n12089), .B2(n10664), .ZN(
        n10657) );
  XNOR2_X1 U12952 ( .A(n10656), .B(n10657), .ZN(n10654) );
  XOR2_X1 U12953 ( .A(n10655), .B(n10654), .Z(n10392) );
  INV_X1 U12954 ( .A(n13859), .ZN(n10389) );
  INV_X1 U12955 ( .A(n13789), .ZN(n13811) );
  AOI22_X1 U12956 ( .A1(n13814), .A2(n13860), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n10387), .ZN(n10388) );
  OAI21_X1 U12957 ( .B1(n10389), .B2(n13811), .A(n10388), .ZN(n10390) );
  AOI21_X1 U12958 ( .B1(n13794), .B2(n12089), .A(n10390), .ZN(n10391) );
  OAI21_X1 U12959 ( .B1(n10392), .B2(n14593), .A(n10391), .ZN(P1_U3237) );
  INV_X1 U12960 ( .A(n10393), .ZN(n10395) );
  INV_X1 U12961 ( .A(SI_18_), .ZN(n10394) );
  OAI222_X1 U12962 ( .A1(n12617), .A2(P3_U3151), .B1(n13021), .B2(n10395), 
        .C1(n10394), .C2(n11761), .ZN(P3_U3277) );
  NAND2_X1 U12963 ( .A1(n15331), .A2(n12888), .ZN(n12907) );
  NAND3_X1 U12964 ( .A1(n10651), .A2(n15253), .A3(n10614), .ZN(n10396) );
  OAI21_X1 U12965 ( .B1(n15244), .B2(n15241), .A(n10396), .ZN(n10509) );
  NOR2_X1 U12966 ( .A1(n15331), .A2(n8192), .ZN(n10397) );
  AOI21_X1 U12967 ( .B1(n10509), .B2(n15331), .A(n10397), .ZN(n10398) );
  OAI21_X1 U12968 ( .B1(n10649), .B2(n12907), .A(n10398), .ZN(P3_U3459) );
  INV_X1 U12969 ( .A(n10399), .ZN(n10424) );
  INV_X1 U12970 ( .A(n11375), .ZN(n10400) );
  OAI222_X1 U12971 ( .A1(n14225), .A2(n10424), .B1(n14216), .B2(n8403), .C1(
        P1_U3086), .C2(n10400), .ZN(P1_U3342) );
  INV_X1 U12972 ( .A(n10416), .ZN(n10402) );
  NAND2_X1 U12973 ( .A1(n10415), .A2(n10403), .ZN(n10404) );
  NAND2_X1 U12974 ( .A1(n9552), .A2(n11116), .ZN(n10929) );
  XOR2_X1 U12975 ( .A(n10929), .B(n11155), .Z(n10409) );
  INV_X1 U12976 ( .A(n10573), .ZN(n10407) );
  NAND2_X1 U12977 ( .A1(n10409), .A2(n10928), .ZN(n11158) );
  OAI21_X1 U12978 ( .B1(n10409), .B2(n10928), .A(n11158), .ZN(n10413) );
  INV_X1 U12979 ( .A(n10896), .ZN(n10410) );
  NOR2_X2 U12980 ( .A1(n10410), .A2(n10414), .ZN(n14972) );
  NOR2_X1 U12981 ( .A1(n14972), .A2(n10411), .ZN(n10412) );
  NAND2_X1 U12982 ( .A1(n10413), .A2(n13148), .ZN(n10420) );
  AOI22_X1 U12983 ( .A1(n13172), .A2(n9559), .B1(n13173), .B2(n13207), .ZN(
        n10577) );
  INV_X1 U12984 ( .A(n10577), .ZN(n10418) );
  NAND2_X1 U12985 ( .A1(n10416), .A2(n10540), .ZN(n10417) );
  NAND2_X1 U12986 ( .A1(n10417), .A2(n10539), .ZN(n10918) );
  OR2_X1 U12987 ( .A1(n14957), .A2(n10918), .ZN(n11161) );
  AOI22_X1 U12988 ( .A1(n13159), .A2(n10418), .B1(n11161), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n10419) );
  OAI211_X1 U12989 ( .C1(n11131), .C2(n13133), .A(n10420), .B(n10419), .ZN(
        P2_U3194) );
  OAI222_X1 U12990 ( .A1(P3_U3151), .A2(n12676), .B1(n11761), .B2(n10422), 
        .C1(n13021), .C2(n10421), .ZN(P3_U3276) );
  INV_X1 U12991 ( .A(n11482), .ZN(n11477) );
  OAI222_X1 U12992 ( .A1(P2_U3088), .A2(n11477), .B1(n13708), .B2(n10424), 
        .C1(n10423), .C2(n13705), .ZN(P2_U3314) );
  MUX2_X1 U12993 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12670), .Z(n10478) );
  XOR2_X1 U12994 ( .A(n10490), .B(n10478), .Z(n10481) );
  MUX2_X1 U12995 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n12670), .Z(n10425) );
  XNOR2_X1 U12996 ( .A(n10425), .B(n6465), .ZN(n10777) );
  MUX2_X1 U12997 ( .A(n8193), .B(n8192), .S(n12670), .Z(n10765) );
  INV_X1 U12998 ( .A(n10764), .ZN(n10775) );
  NAND2_X1 U12999 ( .A1(n10765), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10776) );
  INV_X1 U13000 ( .A(n10776), .ZN(n10427) );
  INV_X1 U13001 ( .A(n10425), .ZN(n10426) );
  MUX2_X1 U13002 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12670), .Z(n10428) );
  XNOR2_X1 U13003 ( .A(n10428), .B(n6709), .ZN(n10460) );
  XOR2_X1 U13004 ( .A(n10481), .B(n10482), .Z(n10459) );
  NAND2_X1 U13005 ( .A1(P3_U3897), .A2(n12328), .ZN(n15158) );
  INV_X1 U13006 ( .A(n10606), .ZN(n10429) );
  OR2_X1 U13007 ( .A1(n10430), .A2(n10429), .ZN(n10432) );
  NAND2_X1 U13008 ( .A1(n10432), .A2(n10431), .ZN(n10443) );
  NOR2_X1 U13009 ( .A1(n10619), .A2(n8862), .ZN(n10442) );
  MUX2_X1 U13010 ( .A(P3_REG2_REG_2__SCAN_IN), .B(n8174), .S(n10464), .Z(
        n10463) );
  NOR2_X1 U13011 ( .A1(n10764), .A2(n8193), .ZN(n10773) );
  INV_X1 U13012 ( .A(n10773), .ZN(n10434) );
  NAND2_X1 U13013 ( .A1(n10448), .A2(n10434), .ZN(n10436) );
  NAND2_X1 U13014 ( .A1(n10435), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10437) );
  NAND2_X1 U13015 ( .A1(n10436), .A2(n10437), .ZN(n10778) );
  OR2_X1 U13016 ( .A1(n10778), .A2(n8203), .ZN(n10780) );
  NAND2_X1 U13017 ( .A1(n10780), .A2(n10437), .ZN(n10462) );
  NAND2_X1 U13018 ( .A1(n10464), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10438) );
  NAND2_X1 U13019 ( .A1(n10439), .A2(n8216), .ZN(n10440) );
  NAND2_X1 U13020 ( .A1(n10488), .A2(n10440), .ZN(n10457) );
  NOR2_X1 U13021 ( .A1(n15170), .A2(n10490), .ZN(n10456) );
  INV_X1 U13022 ( .A(n10442), .ZN(n10444) );
  AND2_X1 U13023 ( .A1(n10444), .A2(n10443), .ZN(n15149) );
  AOI22_X1 U13024 ( .A1(n15149), .A2(P3_ADDR_REG_3__SCAN_IN), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(P3_U3151), .ZN(n10454) );
  NOR2_X2 U13025 ( .A1(n10446), .A2(n10445), .ZN(n15176) );
  MUX2_X1 U13026 ( .A(P3_REG1_REG_2__SCAN_IN), .B(n10447), .S(n10464), .Z(
        n10467) );
  NAND2_X1 U13027 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n10775), .ZN(n10762) );
  NAND2_X1 U13028 ( .A1(n10448), .A2(n10762), .ZN(n10449) );
  OR2_X1 U13029 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10762), .ZN(n10450) );
  NAND2_X1 U13030 ( .A1(n10449), .A2(n10450), .ZN(n10783) );
  INV_X1 U13031 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10782) );
  OR2_X1 U13032 ( .A1(n10783), .A2(n10782), .ZN(n10785) );
  NAND2_X1 U13033 ( .A1(n10785), .A2(n10450), .ZN(n10466) );
  NAND2_X1 U13034 ( .A1(n10467), .A2(n10466), .ZN(n10465) );
  NAND2_X1 U13035 ( .A1(n6709), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10451) );
  NAND2_X1 U13036 ( .A1(n10465), .A2(n10451), .ZN(n10491) );
  INV_X1 U13037 ( .A(n10490), .ZN(n10480) );
  XNOR2_X1 U13038 ( .A(n10491), .B(n10480), .ZN(n10493) );
  XNOR2_X1 U13039 ( .A(n10493), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n10452) );
  NAND2_X1 U13040 ( .A1(n15176), .A2(n10452), .ZN(n10453) );
  NAND2_X1 U13041 ( .A1(n10454), .A2(n10453), .ZN(n10455) );
  AOI211_X1 U13042 ( .C1(n15054), .C2(n10457), .A(n10456), .B(n10455), .ZN(
        n10458) );
  OAI21_X1 U13043 ( .B1(n10459), .B2(n15158), .A(n10458), .ZN(P3_U3185) );
  XOR2_X1 U13044 ( .A(n10460), .B(n6670), .Z(n10475) );
  OAI21_X1 U13045 ( .B1(n10463), .B2(n10462), .A(n10461), .ZN(n10473) );
  NOR2_X1 U13046 ( .A1(n15170), .A2(n6709), .ZN(n10472) );
  OAI21_X1 U13047 ( .B1(n10467), .B2(n10466), .A(n10465), .ZN(n10468) );
  NAND2_X1 U13048 ( .A1(n15176), .A2(n10468), .ZN(n10470) );
  NAND2_X1 U13049 ( .A1(n15149), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n10469) );
  OAI211_X1 U13050 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n15236), .A(n10470), .B(
        n10469), .ZN(n10471) );
  AOI211_X1 U13051 ( .C1(n15054), .C2(n10473), .A(n10472), .B(n10471), .ZN(
        n10474) );
  OAI21_X1 U13052 ( .B1(n10475), .B2(n15158), .A(n10474), .ZN(P3_U3184) );
  NAND2_X1 U13053 ( .A1(n15318), .A2(n12888), .ZN(n12983) );
  NOR2_X1 U13054 ( .A1(n15318), .A2(n8191), .ZN(n10476) );
  AOI21_X1 U13055 ( .B1(n15318), .B2(n10509), .A(n10476), .ZN(n10477) );
  OAI21_X1 U13056 ( .B1(n10649), .B2(n12983), .A(n10477), .ZN(P3_U3390) );
  MUX2_X1 U13057 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12670), .Z(n12627) );
  XNOR2_X1 U13058 ( .A(n12627), .B(n12626), .ZN(n12628) );
  INV_X1 U13059 ( .A(n10478), .ZN(n10479) );
  XOR2_X1 U13060 ( .A(n12628), .B(n12629), .Z(n10500) );
  NAND2_X1 U13061 ( .A1(n10488), .A2(n10486), .ZN(n10484) );
  INV_X1 U13062 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10483) );
  XNOR2_X1 U13063 ( .A(n12626), .B(n10483), .ZN(n10485) );
  NAND2_X1 U13064 ( .A1(n10484), .A2(n10485), .ZN(n12566) );
  INV_X1 U13065 ( .A(n10485), .ZN(n10487) );
  NAND3_X1 U13066 ( .A1(n10488), .A2(n10487), .A3(n10486), .ZN(n10489) );
  NAND2_X1 U13067 ( .A1(n12566), .A2(n10489), .ZN(n10498) );
  NOR2_X1 U13068 ( .A1(n15170), .A2(n12626), .ZN(n10497) );
  INV_X1 U13069 ( .A(n15149), .ZN(n15173) );
  NAND2_X1 U13070 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_U3151), .ZN(n10808) );
  AND2_X1 U13071 ( .A1(n10491), .A2(n10490), .ZN(n10492) );
  AOI21_X1 U13072 ( .B1(n10493), .B2(P3_REG1_REG_3__SCAN_IN), .A(n10492), .ZN(
        n12593) );
  MUX2_X1 U13073 ( .A(n12590), .B(P3_REG1_REG_4__SCAN_IN), .S(n12626), .Z(
        n12592) );
  XNOR2_X1 U13074 ( .A(n12593), .B(n12592), .ZN(n10494) );
  NAND2_X1 U13075 ( .A1(n15176), .A2(n10494), .ZN(n10495) );
  OAI211_X1 U13076 ( .C1(n15173), .C2(n6934), .A(n10808), .B(n10495), .ZN(
        n10496) );
  AOI211_X1 U13077 ( .C1(n15054), .C2(n10498), .A(n10497), .B(n10496), .ZN(
        n10499) );
  OAI21_X1 U13078 ( .B1(n10500), .B2(n15158), .A(n10499), .ZN(P3_U3186) );
  INV_X1 U13079 ( .A(n10501), .ZN(n10504) );
  NAND2_X1 U13080 ( .A1(n10502), .A2(n10505), .ZN(n10503) );
  OAI21_X1 U13081 ( .B1(n10505), .B2(n10504), .A(n10503), .ZN(n10506) );
  OR2_X1 U13082 ( .A1(n10507), .A2(n10506), .ZN(n10510) );
  NOR2_X1 U13083 ( .A1(n15253), .A2(n15267), .ZN(n10508) );
  AOI22_X1 U13084 ( .A1(n10509), .A2(n15273), .B1(P3_REG3_REG_0__SCAN_IN), 
        .B2(n15226), .ZN(n10513) );
  NAND2_X1 U13085 ( .A1(n12860), .A2(n10511), .ZN(n10512) );
  OAI211_X1 U13086 ( .C1(n8193), .C2(n15273), .A(n10513), .B(n10512), .ZN(
        P3_U3233) );
  INV_X1 U13087 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10514) );
  MUX2_X1 U13088 ( .A(n10514), .B(P1_REG1_REG_10__SCAN_IN), .S(n10586), .Z(
        n10517) );
  OAI21_X1 U13089 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n10518), .A(n10515), .ZN(
        n10516) );
  NOR2_X1 U13090 ( .A1(n10516), .A2(n10517), .ZN(n10585) );
  AOI211_X1 U13091 ( .C1(n10517), .C2(n10516), .A(n13911), .B(n10585), .ZN(
        n10528) );
  NAND2_X1 U13092 ( .A1(n10518), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10520) );
  MUX2_X1 U13093 ( .A(n10590), .B(P1_REG2_REG_10__SCAN_IN), .S(n10586), .Z(
        n10519) );
  AOI21_X1 U13094 ( .B1(n10521), .B2(n10520), .A(n10519), .ZN(n10594) );
  INV_X1 U13095 ( .A(n10594), .ZN(n10523) );
  NAND3_X1 U13096 ( .A1(n10521), .A2(n10520), .A3(n10519), .ZN(n10522) );
  NAND3_X1 U13097 ( .A1(n10523), .A2(n14649), .A3(n10522), .ZN(n10526) );
  AND2_X1 U13098 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10524) );
  AOI21_X1 U13099 ( .B1(n14615), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n10524), 
        .ZN(n10525) );
  OAI211_X1 U13100 ( .C1(n14634), .C2(n10591), .A(n10526), .B(n10525), .ZN(
        n10527) );
  OR2_X1 U13101 ( .A1(n10528), .A2(n10527), .ZN(P1_U3253) );
  AND2_X1 U13102 ( .A1(n12065), .A2(n6840), .ZN(n14963) );
  INV_X1 U13103 ( .A(n14963), .ZN(n14987) );
  OAI21_X1 U13104 ( .B1(n10530), .B2(n10533), .A(n10529), .ZN(n11091) );
  INV_X1 U13105 ( .A(n10553), .ZN(n10532) );
  INV_X1 U13106 ( .A(n11115), .ZN(n10531) );
  AOI211_X1 U13107 ( .C1(n10927), .C2(n10532), .A(n13490), .B(n10531), .ZN(
        n11096) );
  XNOR2_X1 U13108 ( .A(n10534), .B(n10533), .ZN(n10537) );
  NAND2_X1 U13109 ( .A1(n13173), .A2(n13204), .ZN(n10536) );
  NAND2_X1 U13110 ( .A1(n13172), .A2(n13206), .ZN(n10535) );
  AND2_X1 U13111 ( .A1(n10536), .A2(n10535), .ZN(n11217) );
  OAI21_X1 U13112 ( .B1(n10537), .B2(n13504), .A(n11217), .ZN(n11092) );
  AOI211_X1 U13113 ( .C1(n14982), .C2(n11091), .A(n11096), .B(n11092), .ZN(
        n10550) );
  OR2_X1 U13114 ( .A1(n10538), .A2(n14957), .ZN(n14955) );
  NAND3_X1 U13115 ( .A1(n10541), .A2(n10540), .A3(n10539), .ZN(n10542) );
  NAND2_X1 U13116 ( .A1(n14995), .A2(n14972), .ZN(n13677) );
  OAI22_X1 U13117 ( .A1(n13677), .A2(n11223), .B1(n14995), .B2(n9151), .ZN(
        n10543) );
  INV_X1 U13118 ( .A(n10543), .ZN(n10544) );
  OAI21_X1 U13119 ( .B1(n10550), .B2(n14994), .A(n10544), .ZN(P2_U3442) );
  INV_X1 U13120 ( .A(n14953), .ZN(n10545) );
  NAND2_X1 U13121 ( .A1(n15002), .A2(n14972), .ZN(n13630) );
  OAI22_X1 U13122 ( .A1(n13630), .A2(n11223), .B1(n15002), .B2(n10547), .ZN(
        n10548) );
  INV_X1 U13123 ( .A(n10548), .ZN(n10549) );
  OAI21_X1 U13124 ( .B1(n10550), .B2(n6478), .A(n10549), .ZN(P2_U3503) );
  OAI21_X1 U13125 ( .B1(n10552), .B2(n10554), .A(n10551), .ZN(n11502) );
  AOI211_X1 U13126 ( .C1(n14818), .C2(n10562), .A(n13490), .B(n10553), .ZN(
        n11496) );
  XNOR2_X1 U13127 ( .A(n10555), .B(n10554), .ZN(n10556) );
  AOI22_X1 U13128 ( .A1(n13172), .A2(n13207), .B1(n13173), .B2(n13205), .ZN(
        n14812) );
  OAI21_X1 U13129 ( .B1(n10556), .B2(n13504), .A(n14812), .ZN(n11499) );
  AOI211_X1 U13130 ( .C1(n14982), .C2(n11502), .A(n11496), .B(n11499), .ZN(
        n10559) );
  AOI22_X1 U13131 ( .A1(n13634), .A2(n14818), .B1(n6478), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n10557) );
  OAI21_X1 U13132 ( .B1(n10559), .B2(n6478), .A(n10557), .ZN(P2_U3502) );
  INV_X1 U13133 ( .A(n13677), .ZN(n13680) );
  AOI22_X1 U13134 ( .A1(n13680), .A2(n14818), .B1(n14994), .B2(
        P2_REG0_REG_3__SCAN_IN), .ZN(n10558) );
  OAI21_X1 U13135 ( .B1(n10559), .B2(n14994), .A(n10558), .ZN(P2_U3439) );
  OAI21_X1 U13136 ( .B1(n10561), .B2(n10564), .A(n10560), .ZN(n11083) );
  INV_X1 U13137 ( .A(n10562), .ZN(n10563) );
  AOI211_X1 U13138 ( .C1(n11166), .C2(n10574), .A(n13490), .B(n10563), .ZN(
        n11086) );
  XNOR2_X1 U13139 ( .A(n10565), .B(n10564), .ZN(n10566) );
  AOI22_X1 U13140 ( .A1(n13172), .A2(n9552), .B1(n13173), .B2(n13206), .ZN(
        n11164) );
  OAI21_X1 U13141 ( .B1(n10566), .B2(n13504), .A(n11164), .ZN(n11087) );
  AOI211_X1 U13142 ( .C1(n14982), .C2(n11083), .A(n11086), .B(n11087), .ZN(
        n10571) );
  INV_X1 U13143 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10567) );
  OAI22_X1 U13144 ( .A1(n13677), .A2(n6909), .B1(n14995), .B2(n10567), .ZN(
        n10568) );
  INV_X1 U13145 ( .A(n10568), .ZN(n10569) );
  OAI21_X1 U13146 ( .B1(n10571), .B2(n14994), .A(n10569), .ZN(P2_U3436) );
  AOI22_X1 U13147 ( .A1(n13634), .A2(n11166), .B1(n6478), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n10570) );
  OAI21_X1 U13148 ( .B1(n10571), .B2(n6478), .A(n10570), .ZN(P2_U3501) );
  OAI21_X1 U13149 ( .B1(n10575), .B2(n10573), .A(n10572), .ZN(n11129) );
  AOI211_X1 U13150 ( .C1(n10897), .C2(n10582), .A(n13490), .B(n6910), .ZN(
        n11133) );
  XOR2_X1 U13151 ( .A(n10576), .B(n10575), .Z(n10578) );
  OAI21_X1 U13152 ( .B1(n10578), .B2(n13504), .A(n10577), .ZN(n11134) );
  AOI211_X1 U13153 ( .C1(n14982), .C2(n11129), .A(n11133), .B(n11134), .ZN(
        n10584) );
  INV_X1 U13154 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10579) );
  OAI22_X1 U13155 ( .A1(n13677), .A2(n11131), .B1(n14995), .B2(n10579), .ZN(
        n10580) );
  INV_X1 U13156 ( .A(n10580), .ZN(n10581) );
  OAI21_X1 U13157 ( .B1(n10584), .B2(n14994), .A(n10581), .ZN(P2_U3433) );
  AOI22_X1 U13158 ( .A1(n13634), .A2(n10582), .B1(n6478), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n10583) );
  OAI21_X1 U13159 ( .B1(n10584), .B2(n6478), .A(n10583), .ZN(P2_U3500) );
  AOI21_X1 U13160 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n10586), .A(n10585), 
        .ZN(n10589) );
  MUX2_X1 U13161 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10587), .S(n10833), .Z(
        n10588) );
  NAND2_X1 U13162 ( .A1(n10589), .A2(n10588), .ZN(n10832) );
  OAI21_X1 U13163 ( .B1(n10589), .B2(n10588), .A(n10832), .ZN(n10600) );
  NOR2_X1 U13164 ( .A1(n10591), .A2(n10590), .ZN(n10593) );
  MUX2_X1 U13165 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n10837), .S(n10833), .Z(
        n10592) );
  OAI21_X1 U13166 ( .B1(n10594), .B2(n10593), .A(n10592), .ZN(n10836) );
  OR3_X1 U13167 ( .A1(n10594), .A2(n10593), .A3(n10592), .ZN(n10595) );
  NAND3_X1 U13168 ( .A1(n10836), .A2(n14649), .A3(n10595), .ZN(n10598) );
  NAND2_X1 U13169 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n11690)
         );
  INV_X1 U13170 ( .A(n11690), .ZN(n10596) );
  AOI21_X1 U13171 ( .B1(n14615), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n10596), 
        .ZN(n10597) );
  OAI211_X1 U13172 ( .C1(n10838), .C2(n14634), .A(n10598), .B(n10597), .ZN(
        n10599) );
  AOI21_X1 U13173 ( .B1(n10600), .B2(n14648), .A(n10599), .ZN(n10601) );
  INV_X1 U13174 ( .A(n10601), .ZN(P1_U3254) );
  INV_X1 U13175 ( .A(n10602), .ZN(n10733) );
  INV_X1 U13176 ( .A(n11885), .ZN(n11796) );
  OAI222_X1 U13177 ( .A1(n14225), .A2(n10733), .B1(n11796), .B2(P1_U3086), 
        .C1(n10603), .C2(n14216), .ZN(P1_U3339) );
  NAND2_X1 U13178 ( .A1(n10605), .A2(n10604), .ZN(n10612) );
  AND2_X1 U13179 ( .A1(n10607), .A2(n10606), .ZN(n10611) );
  INV_X1 U13180 ( .A(n10640), .ZN(n10608) );
  NAND2_X1 U13181 ( .A1(n10642), .A2(n10608), .ZN(n10610) );
  NAND4_X1 U13182 ( .A1(n10612), .A2(n10611), .A3(n10610), .A4(n10609), .ZN(
        n10613) );
  NAND2_X1 U13183 ( .A1(n10613), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10617) );
  INV_X1 U13184 ( .A(n10614), .ZN(n10615) );
  NAND3_X1 U13185 ( .A1(n10642), .A2(n10619), .A3(n10615), .ZN(n10616) );
  INV_X1 U13186 ( .A(n14379), .ZN(n12535) );
  NOR2_X1 U13187 ( .A1(n12535), .A2(P3_U3151), .ZN(n10716) );
  INV_X1 U13188 ( .A(n15254), .ZN(n10632) );
  OR2_X1 U13189 ( .A1(n10639), .A2(n15253), .ZN(n10618) );
  INV_X1 U13190 ( .A(n15258), .ZN(n10724) );
  NAND2_X1 U13191 ( .A1(n10620), .A2(n10619), .ZN(n10621) );
  NOR2_X2 U13192 ( .A1(n12533), .A2(n15241), .ZN(n12545) );
  NOR2_X2 U13193 ( .A1(n12533), .A2(n15243), .ZN(n12522) );
  INV_X1 U13194 ( .A(n12522), .ZN(n12543) );
  INV_X1 U13195 ( .A(n15257), .ZN(n10622) );
  OAI22_X1 U13196 ( .A1(n10724), .A2(n12507), .B1(n12543), .B2(n10622), .ZN(
        n10623) );
  AOI21_X1 U13197 ( .B1(n10632), .B2(n12548), .A(n10623), .ZN(n10648) );
  OAI21_X1 U13198 ( .B1(n10964), .B2(n10627), .A(n10626), .ZN(n10628) );
  INV_X1 U13199 ( .A(n10628), .ZN(n10629) );
  NAND2_X2 U13200 ( .A1(n10630), .A2(n10629), .ZN(n10719) );
  XNOR2_X1 U13201 ( .A(n10719), .B(n10632), .ZN(n10631) );
  NAND2_X1 U13202 ( .A1(n10631), .A2(n15244), .ZN(n10709) );
  NAND3_X1 U13203 ( .A1(n10969), .A2(n12564), .A3(n10632), .ZN(n10633) );
  NAND2_X1 U13204 ( .A1(n10969), .A2(n15260), .ZN(n10634) );
  NAND3_X1 U13205 ( .A1(n10635), .A2(n12386), .A3(n15261), .ZN(n10636) );
  OAI211_X1 U13206 ( .C1(n10637), .C2(n15260), .A(n10710), .B(n10636), .ZN(
        n10646) );
  OR2_X1 U13207 ( .A1(n10639), .A2(n10638), .ZN(n10645) );
  OR2_X1 U13208 ( .A1(n10641), .A2(n10640), .ZN(n10643) );
  OR2_X1 U13209 ( .A1(n10643), .A2(n10642), .ZN(n10644) );
  NAND2_X1 U13210 ( .A1(n10646), .A2(n14376), .ZN(n10647) );
  OAI211_X1 U13211 ( .C1(n10716), .C2(n15269), .A(n10648), .B(n10647), .ZN(
        P3_U3162) );
  INV_X1 U13212 ( .A(n12548), .ZN(n14373) );
  OAI22_X1 U13213 ( .A1(n14373), .A2(n10649), .B1(n12507), .B2(n15244), .ZN(
        n10650) );
  AOI21_X1 U13214 ( .B1(n14376), .B2(n10651), .A(n10650), .ZN(n10652) );
  OAI21_X1 U13215 ( .B1(n10716), .B2(n10653), .A(n10652), .ZN(P3_U3172) );
  INV_X1 U13216 ( .A(n10656), .ZN(n10658) );
  NAND2_X1 U13217 ( .A1(n10658), .A2(n10657), .ZN(n10659) );
  NAND2_X1 U13218 ( .A1(n13859), .A2(n10664), .ZN(n10662) );
  NAND2_X1 U13219 ( .A1(n12035), .A2(n14724), .ZN(n10661) );
  NAND2_X1 U13220 ( .A1(n10662), .A2(n10661), .ZN(n10663) );
  XNOR2_X1 U13221 ( .A(n10663), .B(n12332), .ZN(n10669) );
  NAND2_X1 U13222 ( .A1(n13859), .A2(n11944), .ZN(n10666) );
  NAND2_X1 U13223 ( .A1(n12028), .A2(n14724), .ZN(n10665) );
  NAND2_X1 U13224 ( .A1(n10666), .A2(n10665), .ZN(n10668) );
  XNOR2_X1 U13225 ( .A(n10669), .B(n10668), .ZN(n14594) );
  NAND2_X1 U13226 ( .A1(n10669), .A2(n10668), .ZN(n10670) );
  INV_X1 U13227 ( .A(n10866), .ZN(n10689) );
  NAND2_X1 U13228 ( .A1(n14704), .A2(n12035), .ZN(n10672) );
  NAND2_X1 U13229 ( .A1(n13858), .A2(n10693), .ZN(n10671) );
  NAND2_X1 U13230 ( .A1(n10672), .A2(n10671), .ZN(n10673) );
  XNOR2_X1 U13231 ( .A(n10673), .B(n12025), .ZN(n10868) );
  NAND2_X1 U13232 ( .A1(n14704), .A2(n12028), .ZN(n10675) );
  NAND2_X1 U13233 ( .A1(n13858), .A2(n11944), .ZN(n10674) );
  NAND2_X1 U13234 ( .A1(n14598), .A2(n10664), .ZN(n10677) );
  NAND2_X1 U13235 ( .A1(n12110), .A2(n12035), .ZN(n10676) );
  NAND2_X1 U13236 ( .A1(n10677), .A2(n10676), .ZN(n10678) );
  XNOR2_X1 U13237 ( .A(n10678), .B(n12025), .ZN(n10889) );
  NAND2_X1 U13238 ( .A1(n14598), .A2(n11944), .ZN(n10680) );
  NAND2_X1 U13239 ( .A1(n12110), .A2(n6542), .ZN(n10679) );
  AND2_X1 U13240 ( .A1(n10680), .A2(n10679), .ZN(n10864) );
  OAI22_X1 U13241 ( .A1(n10868), .A2(n10867), .B1(n10889), .B2(n10864), .ZN(
        n10681) );
  NAND2_X1 U13242 ( .A1(n10889), .A2(n10864), .ZN(n10683) );
  INV_X1 U13243 ( .A(n10867), .ZN(n10682) );
  NAND2_X1 U13244 ( .A1(n10683), .A2(n10682), .ZN(n10685) );
  INV_X1 U13245 ( .A(n10683), .ZN(n10684) );
  AOI22_X1 U13246 ( .A1(n10868), .A2(n10685), .B1(n10684), .B2(n10867), .ZN(
        n10686) );
  INV_X1 U13247 ( .A(n10686), .ZN(n10687) );
  NAND2_X1 U13248 ( .A1(n14762), .A2(n12035), .ZN(n10691) );
  NAND2_X1 U13249 ( .A1(n13857), .A2(n12028), .ZN(n10690) );
  NAND2_X1 U13250 ( .A1(n10691), .A2(n10690), .ZN(n10692) );
  XNOR2_X1 U13251 ( .A(n10692), .B(n12332), .ZN(n10816) );
  AND2_X1 U13252 ( .A1(n12039), .A2(n13857), .ZN(n10694) );
  AOI21_X1 U13253 ( .B1(n14762), .B2(n10693), .A(n10694), .ZN(n10814) );
  XNOR2_X1 U13254 ( .A(n10816), .B(n10814), .ZN(n10695) );
  OAI211_X1 U13255 ( .C1(n10696), .C2(n10695), .A(n10818), .B(n14488), .ZN(
        n10706) );
  NAND3_X1 U13256 ( .A1(n10698), .A2(n10697), .A3(n10064), .ZN(n10699) );
  NAND2_X1 U13257 ( .A1(n10699), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10700) );
  AOI21_X1 U13258 ( .B1(n13789), .B2(n13856), .A(n10701), .ZN(n10703) );
  NAND2_X1 U13259 ( .A1(n13814), .A2(n13858), .ZN(n10702) );
  OAI211_X1 U13260 ( .C1(n14606), .C2(n11008), .A(n10703), .B(n10702), .ZN(
        n10704) );
  AOI21_X1 U13261 ( .B1(n13794), .B2(n14762), .A(n10704), .ZN(n10705) );
  NAND2_X1 U13262 ( .A1(n10706), .A2(n10705), .ZN(P1_U3239) );
  INV_X1 U13263 ( .A(n11016), .ZN(n15242) );
  OAI22_X1 U13264 ( .A1(n15244), .A2(n12543), .B1(n12507), .B2(n15242), .ZN(
        n10707) );
  AOI21_X1 U13265 ( .B1(n10708), .B2(n12548), .A(n10707), .ZN(n10715) );
  XNOR2_X1 U13266 ( .A(n10719), .B(n10708), .ZN(n10717) );
  XNOR2_X1 U13267 ( .A(n10717), .B(n15258), .ZN(n10712) );
  NAND2_X1 U13268 ( .A1(n10710), .A2(n10709), .ZN(n10711) );
  NAND2_X1 U13269 ( .A1(n10711), .A2(n10712), .ZN(n10723) );
  OAI21_X1 U13270 ( .B1(n10712), .B2(n10711), .A(n10723), .ZN(n10713) );
  NAND2_X1 U13271 ( .A1(n10713), .A2(n14376), .ZN(n10714) );
  OAI211_X1 U13272 ( .C1(n10716), .C2(n15236), .A(n10715), .B(n10714), .ZN(
        P3_U3177) );
  NAND2_X1 U13273 ( .A1(n10717), .A2(n10724), .ZN(n10720) );
  XNOR2_X1 U13274 ( .A(n10719), .B(n10718), .ZN(n10796) );
  XNOR2_X1 U13275 ( .A(n10796), .B(n11016), .ZN(n10721) );
  AOI21_X1 U13276 ( .B1(n10723), .B2(n10720), .A(n10721), .ZN(n10729) );
  AND2_X1 U13277 ( .A1(n10721), .A2(n10720), .ZN(n10722) );
  NAND2_X1 U13278 ( .A1(n10799), .A2(n14376), .ZN(n10728) );
  INV_X1 U13279 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n15225) );
  OAI22_X1 U13280 ( .A1(n12543), .A2(n10724), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15225), .ZN(n10726) );
  INV_X1 U13281 ( .A(n15217), .ZN(n15208) );
  OAI22_X1 U13282 ( .A1(n14373), .A2(n15224), .B1(n12507), .B2(n15208), .ZN(
        n10725) );
  AOI211_X1 U13283 ( .C1(n15225), .C2(n12535), .A(n10726), .B(n10725), .ZN(
        n10727) );
  OAI21_X1 U13284 ( .B1(n10729), .B2(n10728), .A(n10727), .ZN(P3_U3158) );
  INV_X1 U13285 ( .A(n10730), .ZN(n10736) );
  INV_X1 U13286 ( .A(n11781), .ZN(n11791) );
  OAI222_X1 U13287 ( .A1(n14225), .A2(n10736), .B1(n11791), .B2(P1_U3086), 
        .C1(n10731), .C2(n14216), .ZN(P1_U3341) );
  INV_X1 U13288 ( .A(n14938), .ZN(n10734) );
  OAI222_X1 U13289 ( .A1(P2_U3088), .A2(n10734), .B1(n13708), .B2(n10733), 
        .C1(n10732), .C2(n13705), .ZN(P2_U3311) );
  INV_X1 U13290 ( .A(n13238), .ZN(n11480) );
  OAI222_X1 U13291 ( .A1(P2_U3088), .A2(n11480), .B1(n13708), .B2(n10736), 
        .C1(n10735), .C2(n13705), .ZN(P2_U3313) );
  OAI21_X1 U13292 ( .B1(n10744), .B2(P2_REG2_REG_9__SCAN_IN), .A(n10737), .ZN(
        n14914) );
  INV_X1 U13293 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10738) );
  MUX2_X1 U13294 ( .A(n10738), .B(P2_REG2_REG_10__SCAN_IN), .S(n14911), .Z(
        n14915) );
  NOR2_X1 U13295 ( .A1(n14914), .A2(n14915), .ZN(n14912) );
  AOI21_X1 U13296 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n14911), .A(n14912), 
        .ZN(n10740) );
  MUX2_X1 U13297 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n13523), .S(n10849), .Z(
        n10739) );
  NAND2_X1 U13298 ( .A1(n10740), .A2(n10739), .ZN(n10856) );
  OAI21_X1 U13299 ( .B1(n10740), .B2(n10739), .A(n10856), .ZN(n10751) );
  INV_X1 U13300 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n12426) );
  NOR2_X1 U13301 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n12426), .ZN(n10741) );
  AOI21_X1 U13302 ( .B1(n14924), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n10741), 
        .ZN(n10742) );
  OAI21_X1 U13303 ( .B1(n10853), .B2(n14930), .A(n10742), .ZN(n10750) );
  OAI21_X1 U13304 ( .B1(n10744), .B2(P2_REG1_REG_9__SCAN_IN), .A(n10743), .ZN(
        n14907) );
  MUX2_X1 U13305 ( .A(n10745), .B(P2_REG1_REG_10__SCAN_IN), .S(n14911), .Z(
        n14908) );
  NOR2_X1 U13306 ( .A1(n14907), .A2(n14908), .ZN(n14906) );
  MUX2_X1 U13307 ( .A(n10746), .B(P2_REG1_REG_11__SCAN_IN), .S(n10849), .Z(
        n10747) );
  AOI211_X1 U13308 ( .C1(n10748), .C2(n10747), .A(n14932), .B(n10848), .ZN(
        n10749) );
  AOI211_X1 U13309 ( .C1(n14941), .C2(n10751), .A(n10750), .B(n10749), .ZN(
        n10752) );
  INV_X1 U13310 ( .A(n10752), .ZN(P2_U3225) );
  OAI222_X1 U13311 ( .A1(P3_U3151), .A2(n10755), .B1(n11761), .B2(n10754), 
        .C1(n13021), .C2(n10753), .ZN(P3_U3275) );
  INV_X1 U13312 ( .A(n10756), .ZN(n10760) );
  INV_X1 U13313 ( .A(n13890), .ZN(n13887) );
  OAI222_X1 U13314 ( .A1(n14225), .A2(n10760), .B1(n13887), .B2(P1_U3086), 
        .C1(n10757), .C2(n14216), .ZN(P1_U3338) );
  INV_X1 U13315 ( .A(n10758), .ZN(n10795) );
  INV_X1 U13316 ( .A(n14646), .ZN(n11793) );
  OAI222_X1 U13317 ( .A1(n14225), .A2(n10795), .B1(n11793), .B2(P1_U3086), 
        .C1(n10759), .C2(n14216), .ZN(P1_U3340) );
  INV_X1 U13318 ( .A(n13255), .ZN(n13250) );
  OAI222_X1 U13319 ( .A1(n13705), .A2(n10761), .B1(n13708), .B2(n10760), .C1(
        P2_U3088), .C2(n13250), .ZN(P2_U3310) );
  INV_X1 U13320 ( .A(n10762), .ZN(n10763) );
  NAND2_X1 U13321 ( .A1(n15176), .A2(n10763), .ZN(n10769) );
  INV_X1 U13322 ( .A(n15158), .ZN(n15178) );
  NOR2_X1 U13323 ( .A1(n10765), .A2(n10764), .ZN(n10766) );
  AOI22_X1 U13324 ( .A1(n15178), .A2(n10766), .B1(P3_REG3_REG_0__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10768) );
  NAND2_X1 U13325 ( .A1(n15149), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n10767) );
  NAND3_X1 U13326 ( .A1(n10769), .A2(n10768), .A3(n10767), .ZN(n10772) );
  NOR3_X1 U13327 ( .A1(n15054), .A2(n15176), .A3(n15178), .ZN(n10770) );
  NOR2_X1 U13328 ( .A1(n10770), .A2(n10776), .ZN(n10771) );
  AOI211_X1 U13329 ( .C1(n10773), .C2(n15054), .A(n10772), .B(n10771), .ZN(
        n10774) );
  OAI21_X1 U13330 ( .B1(n10775), .B2(n15170), .A(n10774), .ZN(P3_U3182) );
  XNOR2_X1 U13331 ( .A(n10777), .B(n10776), .ZN(n10793) );
  NAND2_X1 U13332 ( .A1(n10778), .A2(n8203), .ZN(n10779) );
  NAND2_X1 U13333 ( .A1(n10780), .A2(n10779), .ZN(n10791) );
  NOR2_X1 U13334 ( .A1(n15170), .A2(n10781), .ZN(n10790) );
  NAND2_X1 U13335 ( .A1(n10783), .A2(n10782), .ZN(n10784) );
  NAND2_X1 U13336 ( .A1(n10785), .A2(n10784), .ZN(n10786) );
  NAND2_X1 U13337 ( .A1(n15176), .A2(n10786), .ZN(n10788) );
  NAND2_X1 U13338 ( .A1(n15149), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n10787) );
  OAI211_X1 U13339 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n15269), .A(n10788), .B(
        n10787), .ZN(n10789) );
  AOI211_X1 U13340 ( .C1(n15054), .C2(n10791), .A(n10790), .B(n10789), .ZN(
        n10792) );
  OAI21_X1 U13341 ( .B1(n15158), .B2(n10793), .A(n10792), .ZN(P3_U3183) );
  INV_X1 U13342 ( .A(n13228), .ZN(n14929) );
  OAI222_X1 U13343 ( .A1(P2_U3088), .A2(n14929), .B1(n13708), .B2(n10795), 
        .C1(n10794), .C2(n13705), .ZN(P2_U3312) );
  INV_X1 U13344 ( .A(n10796), .ZN(n10797) );
  NAND2_X1 U13345 ( .A1(n10797), .A2(n11016), .ZN(n10798) );
  XNOR2_X1 U13346 ( .A(n12386), .B(n11014), .ZN(n10800) );
  NAND2_X1 U13347 ( .A1(n10800), .A2(n15208), .ZN(n10970) );
  INV_X1 U13348 ( .A(n10800), .ZN(n10801) );
  NAND2_X1 U13349 ( .A1(n10801), .A2(n15217), .ZN(n10802) );
  NAND2_X1 U13350 ( .A1(n10970), .A2(n10802), .ZN(n10806) );
  INV_X1 U13351 ( .A(n10807), .ZN(n10804) );
  INV_X1 U13352 ( .A(n10971), .ZN(n10805) );
  AOI21_X1 U13353 ( .B1(n10807), .B2(n10806), .A(n10805), .ZN(n10813) );
  INV_X1 U13354 ( .A(n11015), .ZN(n10811) );
  AOI22_X1 U13355 ( .A1(n12548), .A2(n11014), .B1(n12545), .B2(n15189), .ZN(
        n10809) );
  OAI211_X1 U13356 ( .C1(n15242), .C2(n12543), .A(n10809), .B(n10808), .ZN(
        n10810) );
  AOI21_X1 U13357 ( .B1(n10811), .B2(n12535), .A(n10810), .ZN(n10812) );
  OAI21_X1 U13358 ( .B1(n10813), .B2(n12550), .A(n10812), .ZN(P3_U3170) );
  INV_X1 U13359 ( .A(n10814), .ZN(n10815) );
  NAND2_X1 U13360 ( .A1(n10816), .A2(n10815), .ZN(n10817) );
  NAND2_X1 U13361 ( .A1(n14681), .A2(n12035), .ZN(n10820) );
  NAND2_X1 U13362 ( .A1(n13856), .A2(n12028), .ZN(n10819) );
  NAND2_X1 U13363 ( .A1(n10820), .A2(n10819), .ZN(n10821) );
  XNOR2_X1 U13364 ( .A(n10821), .B(n12332), .ZN(n10987) );
  AND2_X1 U13365 ( .A1(n12039), .A2(n13856), .ZN(n10822) );
  AOI21_X1 U13366 ( .B1(n14681), .B2(n12028), .A(n10822), .ZN(n10985) );
  XNOR2_X1 U13367 ( .A(n10987), .B(n10985), .ZN(n10823) );
  OAI211_X1 U13368 ( .C1(n10824), .C2(n10823), .A(n10989), .B(n14488), .ZN(
        n10830) );
  INV_X1 U13369 ( .A(n13836), .ZN(n14601) );
  NAND2_X1 U13370 ( .A1(n13857), .A2(n14596), .ZN(n10826) );
  NAND2_X1 U13371 ( .A1(n13855), .A2(n14597), .ZN(n10825) );
  NAND2_X1 U13372 ( .A1(n10826), .A2(n10825), .ZN(n14678) );
  NOR2_X1 U13373 ( .A1(n14606), .A2(n14679), .ZN(n10827) );
  AOI211_X1 U13374 ( .C1(n14601), .C2(n14678), .A(n10828), .B(n10827), .ZN(
        n10829) );
  OAI211_X1 U13375 ( .C1(n14769), .C2(n13817), .A(n10830), .B(n10829), .ZN(
        P1_U3213) );
  MUX2_X1 U13376 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10831), .S(n11236), .Z(
        n10835) );
  OAI21_X1 U13377 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n10833), .A(n10832), 
        .ZN(n10834) );
  NAND2_X1 U13378 ( .A1(n10834), .A2(n10835), .ZN(n11230) );
  OAI21_X1 U13379 ( .B1(n10835), .B2(n10834), .A(n11230), .ZN(n10846) );
  OAI21_X1 U13380 ( .B1(n10838), .B2(n10837), .A(n10836), .ZN(n10841) );
  AOI22_X1 U13381 ( .A1(n11236), .A2(n11632), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n10839), .ZN(n10840) );
  NOR2_X1 U13382 ( .A1(n10840), .A2(n10841), .ZN(n11237) );
  AOI21_X1 U13383 ( .B1(n10841), .B2(n10840), .A(n11237), .ZN(n10844) );
  AND2_X1 U13384 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n11756) );
  AOI21_X1 U13385 ( .B1(n14615), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n11756), 
        .ZN(n10843) );
  NAND2_X1 U13386 ( .A1(n14645), .A2(n11236), .ZN(n10842) );
  OAI211_X1 U13387 ( .C1(n10844), .C2(n13899), .A(n10843), .B(n10842), .ZN(
        n10845) );
  AOI21_X1 U13388 ( .B1(n10846), .B2(n14648), .A(n10845), .ZN(n10847) );
  INV_X1 U13389 ( .A(n10847), .ZN(P1_U3255) );
  MUX2_X1 U13390 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n10850), .S(n11102), .Z(
        n10851) );
  OAI21_X1 U13391 ( .B1(n10852), .B2(n10851), .A(n11101), .ZN(n10862) );
  INV_X1 U13392 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n13523) );
  NAND2_X1 U13393 ( .A1(n10853), .A2(n13523), .ZN(n10854) );
  MUX2_X1 U13394 ( .A(n11584), .B(P2_REG2_REG_12__SCAN_IN), .S(n11102), .Z(
        n10855) );
  AOI21_X1 U13395 ( .B1(n10856), .B2(n10854), .A(n10855), .ZN(n11105) );
  INV_X1 U13396 ( .A(n11105), .ZN(n10858) );
  NAND3_X1 U13397 ( .A1(n10856), .A2(n10855), .A3(n10854), .ZN(n10857) );
  AOI21_X1 U13398 ( .B1(n10858), .B2(n10857), .A(n14913), .ZN(n10861) );
  NAND2_X1 U13399 ( .A1(n14924), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n10859) );
  NAND2_X1 U13400 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n11272)
         );
  OAI211_X1 U13401 ( .C1(n14930), .C2(n11106), .A(n10859), .B(n11272), .ZN(
        n10860) );
  AOI211_X1 U13402 ( .C1(n10862), .C2(n14863), .A(n10861), .B(n10860), .ZN(
        n10863) );
  INV_X1 U13403 ( .A(n10863), .ZN(P2_U3226) );
  INV_X1 U13404 ( .A(n10864), .ZN(n10865) );
  XOR2_X1 U13405 ( .A(n10866), .B(n10864), .Z(n10888) );
  NOR2_X1 U13406 ( .A1(n10888), .A2(n10889), .ZN(n10887) );
  AOI21_X1 U13407 ( .B1(n10866), .B2(n10865), .A(n10887), .ZN(n10870) );
  XNOR2_X1 U13408 ( .A(n10868), .B(n10867), .ZN(n10869) );
  XNOR2_X1 U13409 ( .A(n10870), .B(n10869), .ZN(n10877) );
  NAND2_X1 U13410 ( .A1(n13814), .A2(n14598), .ZN(n10873) );
  NAND2_X1 U13411 ( .A1(n13789), .A2(n13857), .ZN(n10872) );
  NAND3_X1 U13412 ( .A1(n10873), .A2(n10872), .A3(n10871), .ZN(n10875) );
  NOR2_X1 U13413 ( .A1(n14606), .A2(n14700), .ZN(n10874) );
  AOI211_X1 U13414 ( .C1(n13794), .C2(n14704), .A(n10875), .B(n10874), .ZN(
        n10876) );
  OAI21_X1 U13415 ( .B1(n10877), .B2(n14593), .A(n10876), .ZN(P1_U3227) );
  AOI21_X1 U13416 ( .B1(n10878), .B2(n14721), .A(n14731), .ZN(n10886) );
  OAI21_X1 U13417 ( .B1(n14736), .B2(n14691), .A(n14107), .ZN(n10883) );
  OAI22_X1 U13418 ( .A1(n14721), .A2(n10880), .B1(n10879), .B2(n14719), .ZN(
        n10881) );
  AOI21_X1 U13419 ( .B1(n10883), .B2(n10882), .A(n10881), .ZN(n10884) );
  OAI21_X1 U13420 ( .B1(n10886), .B2(n10885), .A(n10884), .ZN(P1_U3293) );
  AOI211_X1 U13421 ( .C1(n10889), .C2(n10888), .A(n14593), .B(n10887), .ZN(
        n10890) );
  INV_X1 U13422 ( .A(n10890), .ZN(n10895) );
  NAND2_X1 U13423 ( .A1(n13859), .A2(n14596), .ZN(n10892) );
  NAND2_X1 U13424 ( .A1(n13858), .A2(n14597), .ZN(n10891) );
  AND2_X1 U13425 ( .A1(n10892), .A2(n10891), .ZN(n11078) );
  NAND2_X1 U13426 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n14637) );
  OAI21_X1 U13427 ( .B1(n13836), .B2(n11078), .A(n14637), .ZN(n10893) );
  AOI21_X1 U13428 ( .B1(n13794), .B2(n12110), .A(n10893), .ZN(n10894) );
  OAI211_X1 U13429 ( .C1(n14606), .C2(n11072), .A(n10895), .B(n10894), .ZN(
        P1_U3230) );
  OR2_X1 U13430 ( .A1(n13517), .A2(n6669), .ZN(n10905) );
  INV_X2 U13431 ( .A(n13517), .ZN(n13519) );
  NAND2_X1 U13432 ( .A1(n10897), .A2(n10896), .ZN(n14959) );
  INV_X1 U13433 ( .A(n14961), .ZN(n10899) );
  NAND2_X1 U13434 ( .A1(n14986), .A2(n13504), .ZN(n10898) );
  AND2_X1 U13435 ( .A1(n13173), .A2(n9552), .ZN(n11143) );
  AOI21_X1 U13436 ( .B1(n10899), .B2(n10898), .A(n11143), .ZN(n14960) );
  OAI21_X1 U13437 ( .B1(n6840), .B2(n14959), .A(n14960), .ZN(n10903) );
  OAI22_X1 U13438 ( .A1(n13519), .A2(n10901), .B1(n10900), .B2(n13521), .ZN(
        n10902) );
  AOI21_X1 U13439 ( .B1(n13519), .B2(n10903), .A(n10902), .ZN(n10904) );
  OAI21_X1 U13440 ( .B1(n10905), .B2(n14961), .A(n10904), .ZN(P2_U3265) );
  OR2_X1 U13441 ( .A1(n10906), .A2(n13915), .ZN(n12265) );
  INV_X1 U13442 ( .A(n12265), .ZN(n10907) );
  AND2_X1 U13443 ( .A1(n14721), .A2(n10907), .ZN(n14732) );
  INV_X1 U13444 ( .A(n14732), .ZN(n14094) );
  MUX2_X1 U13445 ( .A(n10909), .B(n10908), .S(n14721), .Z(n10914) );
  OAI22_X1 U13446 ( .A1(n14103), .A2(n12092), .B1(n10910), .B2(n14719), .ZN(
        n10911) );
  AOI21_X1 U13447 ( .B1(n14731), .B2(n10912), .A(n10911), .ZN(n10913) );
  OAI211_X1 U13448 ( .C1(n10915), .C2(n14094), .A(n10914), .B(n10913), .ZN(
        P1_U3291) );
  INV_X1 U13449 ( .A(n10916), .ZN(n10917) );
  NAND2_X1 U13450 ( .A1(n13172), .A2(n13204), .ZN(n10921) );
  NAND2_X1 U13451 ( .A1(n13173), .A2(n13202), .ZN(n10920) );
  NAND2_X1 U13452 ( .A1(n10921), .A2(n10920), .ZN(n11284) );
  NAND2_X1 U13453 ( .A1(n13159), .A2(n11284), .ZN(n10922) );
  NAND2_X1 U13454 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n14877) );
  OAI211_X1 U13455 ( .C1(n14832), .C2(n11292), .A(n10922), .B(n14877), .ZN(
        n10958) );
  XNOR2_X1 U13456 ( .A(n10959), .B(n6468), .ZN(n10923) );
  AND2_X1 U13457 ( .A1(n13203), .A2(n6474), .ZN(n10924) );
  NAND2_X1 U13458 ( .A1(n10923), .A2(n10924), .ZN(n11037) );
  INV_X1 U13459 ( .A(n10923), .ZN(n11187) );
  INV_X1 U13460 ( .A(n10924), .ZN(n10925) );
  NAND2_X1 U13461 ( .A1(n11187), .A2(n10925), .ZN(n10926) );
  NAND2_X1 U13462 ( .A1(n11037), .A2(n10926), .ZN(n10956) );
  NAND2_X1 U13463 ( .A1(n13205), .A2(n11116), .ZN(n10945) );
  XNOR2_X1 U13464 ( .A(n12351), .B(n10945), .ZN(n11226) );
  XNOR2_X1 U13465 ( .A(n10932), .B(n14818), .ZN(n10938) );
  AND2_X1 U13466 ( .A1(n13206), .A2(n11116), .ZN(n10939) );
  NAND2_X1 U13467 ( .A1(n10938), .A2(n10939), .ZN(n10941) );
  AND2_X1 U13468 ( .A1(n11226), .A2(n10941), .ZN(n10944) );
  OAI21_X1 U13469 ( .B1(n11155), .B2(n10929), .A(n10928), .ZN(n10931) );
  NAND2_X1 U13470 ( .A1(n11155), .A2(n10929), .ZN(n10930) );
  NAND2_X1 U13471 ( .A1(n10931), .A2(n10930), .ZN(n10933) );
  NAND2_X1 U13472 ( .A1(n13207), .A2(n11116), .ZN(n10935) );
  XNOR2_X1 U13473 ( .A(n10934), .B(n10935), .ZN(n11157) );
  INV_X1 U13474 ( .A(n10934), .ZN(n10936) );
  NAND2_X1 U13475 ( .A1(n10936), .A2(n10935), .ZN(n10937) );
  INV_X1 U13476 ( .A(n14815), .ZN(n10943) );
  INV_X1 U13477 ( .A(n10938), .ZN(n11213) );
  INV_X1 U13478 ( .A(n10939), .ZN(n10940) );
  NAND2_X1 U13479 ( .A1(n10944), .A2(n11212), .ZN(n11216) );
  INV_X1 U13480 ( .A(n12351), .ZN(n10946) );
  NAND2_X1 U13481 ( .A1(n10946), .A2(n10945), .ZN(n10947) );
  NAND2_X1 U13482 ( .A1(n11216), .A2(n10947), .ZN(n10948) );
  XNOR2_X1 U13483 ( .A(n10932), .B(n14964), .ZN(n10949) );
  NAND2_X1 U13484 ( .A1(n13204), .A2(n6474), .ZN(n10950) );
  XNOR2_X1 U13485 ( .A(n10949), .B(n10950), .ZN(n12352) );
  INV_X1 U13486 ( .A(n10949), .ZN(n10951) );
  NAND2_X1 U13487 ( .A1(n10951), .A2(n10950), .ZN(n10952) );
  INV_X1 U13488 ( .A(n11186), .ZN(n10954) );
  AOI211_X1 U13489 ( .C1(n10956), .C2(n10955), .A(n14824), .B(n10954), .ZN(
        n10957) );
  AOI211_X1 U13490 ( .C1(n10959), .C2(n14829), .A(n10958), .B(n10957), .ZN(
        n10960) );
  INV_X1 U13491 ( .A(n10960), .ZN(P2_U3211) );
  INV_X1 U13492 ( .A(n10961), .ZN(n10963) );
  INV_X1 U13493 ( .A(SI_21_), .ZN(n10962) );
  OAI222_X1 U13494 ( .A1(n10964), .A2(P3_U3151), .B1(n13021), .B2(n10963), 
        .C1(n10962), .C2(n11761), .ZN(P3_U3274) );
  INV_X1 U13495 ( .A(n10965), .ZN(n10968) );
  OAI22_X1 U13496 ( .A1(n10966), .A2(P3_U3151), .B1(SI_22_), .B2(n13023), .ZN(
        n10967) );
  AOI21_X1 U13497 ( .B1(n10968), .B2(n11150), .A(n10967), .ZN(P3_U3273) );
  INV_X4 U13498 ( .A(n10969), .ZN(n12386) );
  XNOR2_X1 U13499 ( .A(n12386), .B(n15210), .ZN(n11026) );
  XNOR2_X1 U13500 ( .A(n11026), .B(n11027), .ZN(n10973) );
  OAI21_X1 U13501 ( .B1(n10973), .B2(n10972), .A(n11313), .ZN(n10979) );
  INV_X1 U13502 ( .A(n15210), .ZN(n10974) );
  AOI22_X1 U13503 ( .A1(n12548), .A2(n10974), .B1(n12545), .B2(n12562), .ZN(
        n10977) );
  NOR2_X1 U13504 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10975), .ZN(n15012) );
  AOI21_X1 U13505 ( .B1(n12522), .B2(n15217), .A(n15012), .ZN(n10976) );
  OAI211_X1 U13506 ( .C1(n14379), .C2(n15211), .A(n10977), .B(n10976), .ZN(
        n10978) );
  AOI21_X1 U13507 ( .B1(n10979), .B2(n14376), .A(n10978), .ZN(n10980) );
  INV_X1 U13508 ( .A(n10980), .ZN(P3_U3167) );
  NAND2_X1 U13509 ( .A1(n12127), .A2(n12035), .ZN(n10982) );
  NAND2_X1 U13510 ( .A1(n13855), .A2(n12028), .ZN(n10981) );
  NAND2_X1 U13511 ( .A1(n10982), .A2(n10981), .ZN(n10983) );
  XNOR2_X1 U13512 ( .A(n10983), .B(n12025), .ZN(n11438) );
  AND2_X1 U13513 ( .A1(n12039), .A2(n13855), .ZN(n10984) );
  AOI21_X1 U13514 ( .B1(n12127), .B2(n10693), .A(n10984), .ZN(n11437) );
  XNOR2_X1 U13515 ( .A(n11438), .B(n11437), .ZN(n10992) );
  INV_X1 U13516 ( .A(n10985), .ZN(n10986) );
  NAND2_X1 U13517 ( .A1(n10987), .A2(n10986), .ZN(n10988) );
  INV_X1 U13518 ( .A(n11440), .ZN(n10990) );
  AOI21_X1 U13519 ( .B1(n10992), .B2(n10991), .A(n10990), .ZN(n10998) );
  AOI21_X1 U13520 ( .B1(n13789), .B2(n13854), .A(n10993), .ZN(n10995) );
  NAND2_X1 U13521 ( .A1(n13814), .A2(n13856), .ZN(n10994) );
  OAI211_X1 U13522 ( .C1(n14606), .C2(n11205), .A(n10995), .B(n10994), .ZN(
        n10996) );
  AOI21_X1 U13523 ( .B1(n13794), .B2(n12127), .A(n10996), .ZN(n10997) );
  OAI21_X1 U13524 ( .B1(n10998), .B2(n14593), .A(n10997), .ZN(P1_U3221) );
  XNOR2_X1 U13525 ( .A(n10999), .B(n12278), .ZN(n14765) );
  OAI21_X1 U13526 ( .B1(n11001), .B2(n12278), .A(n11000), .ZN(n11006) );
  OAI22_X1 U13527 ( .A1(n11003), .A2(n14696), .B1(n11002), .B2(n14694), .ZN(
        n11005) );
  NOR2_X1 U13528 ( .A1(n14765), .A2(n14660), .ZN(n11004) );
  AOI211_X1 U13529 ( .C1(n14716), .C2(n11006), .A(n11005), .B(n11004), .ZN(
        n14764) );
  MUX2_X1 U13530 ( .A(n11007), .B(n14764), .S(n14721), .Z(n11012) );
  AOI211_X1 U13531 ( .C1(n14762), .C2(n14706), .A(n14792), .B(n14684), .ZN(
        n14760) );
  OAI22_X1 U13532 ( .A1(n14103), .A2(n11009), .B1(n14719), .B2(n11008), .ZN(
        n11010) );
  AOI21_X1 U13533 ( .B1(n14760), .B2(n14731), .A(n11010), .ZN(n11011) );
  OAI211_X1 U13534 ( .C1(n14765), .C2(n14094), .A(n11012), .B(n11011), .ZN(
        P1_U3287) );
  INV_X1 U13535 ( .A(n11022), .ZN(n15290) );
  NAND2_X1 U13536 ( .A1(n15237), .A2(n11013), .ZN(n11617) );
  INV_X1 U13537 ( .A(n11617), .ZN(n15251) );
  NAND2_X1 U13538 ( .A1(n15273), .A2(n15251), .ZN(n15270) );
  INV_X1 U13539 ( .A(n15270), .ZN(n11530) );
  INV_X1 U13540 ( .A(n15227), .ZN(n11619) );
  NAND2_X1 U13541 ( .A1(n11014), .A2(n12888), .ZN(n15287) );
  OAI22_X1 U13542 ( .A1(n11619), .A2(n15287), .B1(n11015), .B2(n15268), .ZN(
        n11024) );
  AOI22_X1 U13543 ( .A1(n15259), .A2(n15189), .B1(n11016), .B2(n15256), .ZN(
        n11021) );
  OAI211_X1 U13544 ( .C1(n11019), .C2(n11018), .A(n11017), .B(n15262), .ZN(
        n11020) );
  OAI211_X1 U13545 ( .C1(n11022), .C2(n15266), .A(n11021), .B(n11020), .ZN(
        n15288) );
  MUX2_X1 U13546 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n15288), .S(n15273), .Z(
        n11023) );
  AOI211_X1 U13547 ( .C1(n15290), .C2(n11530), .A(n11024), .B(n11023), .ZN(
        n11025) );
  INV_X1 U13548 ( .A(n11025), .ZN(P3_U3229) );
  INV_X1 U13549 ( .A(n11026), .ZN(n11028) );
  NAND2_X1 U13550 ( .A1(n11028), .A2(n11027), .ZN(n11311) );
  NAND2_X1 U13551 ( .A1(n11313), .A2(n11311), .ZN(n11031) );
  XNOR2_X1 U13552 ( .A(n12386), .B(n11029), .ZN(n11314) );
  INV_X1 U13553 ( .A(n12562), .ZN(n15207) );
  XNOR2_X1 U13554 ( .A(n11314), .B(n15207), .ZN(n11030) );
  AOI21_X1 U13555 ( .B1(n11031), .B2(n11030), .A(n12550), .ZN(n11032) );
  OR2_X1 U13556 ( .A1(n11031), .A2(n11030), .ZN(n11335) );
  NAND2_X1 U13557 ( .A1(n11032), .A2(n11335), .ZN(n11036) );
  NAND2_X1 U13558 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n15037) );
  INV_X1 U13559 ( .A(n15037), .ZN(n11034) );
  INV_X1 U13560 ( .A(n15190), .ZN(n11316) );
  OAI22_X1 U13561 ( .A1(n14373), .A2(n15196), .B1(n12507), .B2(n11316), .ZN(
        n11033) );
  AOI211_X1 U13562 ( .C1(n12522), .C2(n15189), .A(n11034), .B(n11033), .ZN(
        n11035) );
  OAI211_X1 U13563 ( .C1(n15197), .C2(n14379), .A(n11036), .B(n11035), .ZN(
        P3_U3179) );
  INV_X1 U13564 ( .A(n11493), .ZN(n11348) );
  XNOR2_X1 U13565 ( .A(n11038), .B(n6469), .ZN(n11039) );
  AND2_X1 U13566 ( .A1(n13202), .A2(n13490), .ZN(n11040) );
  NAND2_X1 U13567 ( .A1(n11039), .A2(n11040), .ZN(n11044) );
  INV_X1 U13568 ( .A(n11039), .ZN(n11171) );
  INV_X1 U13569 ( .A(n11040), .ZN(n11041) );
  NAND2_X1 U13570 ( .A1(n11171), .A2(n11041), .ZN(n11042) );
  AND2_X1 U13571 ( .A1(n11044), .A2(n11042), .ZN(n11184) );
  NAND2_X2 U13572 ( .A1(n11043), .A2(n11184), .ZN(n11188) );
  XNOR2_X1 U13573 ( .A(n11180), .B(n6469), .ZN(n11046) );
  NAND2_X1 U13574 ( .A1(n13201), .A2(n13490), .ZN(n11047) );
  XNOR2_X1 U13575 ( .A(n11046), .B(n11047), .ZN(n11182) );
  AND2_X1 U13576 ( .A1(n11182), .A2(n11044), .ZN(n11045) );
  INV_X1 U13577 ( .A(n11046), .ZN(n11257) );
  NAND2_X1 U13578 ( .A1(n11257), .A2(n11047), .ZN(n11048) );
  XNOR2_X1 U13579 ( .A(n11363), .B(n6469), .ZN(n11050) );
  NAND2_X1 U13580 ( .A1(n13200), .A2(n13490), .ZN(n11051) );
  XNOR2_X1 U13581 ( .A(n11050), .B(n11051), .ZN(n11255) );
  INV_X1 U13582 ( .A(n11050), .ZN(n11052) );
  NAND2_X1 U13583 ( .A1(n11052), .A2(n11051), .ZN(n11058) );
  NAND2_X1 U13584 ( .A1(n11263), .A2(n11058), .ZN(n11055) );
  XNOR2_X1 U13585 ( .A(n11493), .B(n6469), .ZN(n12420) );
  AND2_X1 U13586 ( .A1(n13199), .A2(n13490), .ZN(n11053) );
  NAND2_X1 U13587 ( .A1(n12420), .A2(n11053), .ZN(n11264) );
  NAND2_X1 U13588 ( .A1(n11264), .A2(n11054), .ZN(n11056) );
  AOI21_X1 U13589 ( .B1(n11055), .B2(n11056), .A(n14824), .ZN(n11060) );
  INV_X1 U13590 ( .A(n11056), .ZN(n11057) );
  AND2_X1 U13591 ( .A1(n11058), .A2(n11057), .ZN(n11059) );
  NAND2_X1 U13592 ( .A1(n11060), .A2(n12422), .ZN(n11066) );
  INV_X1 U13593 ( .A(n11349), .ZN(n11064) );
  NAND2_X1 U13594 ( .A1(n13172), .A2(n13200), .ZN(n11062) );
  NAND2_X1 U13595 ( .A1(n13173), .A2(n13198), .ZN(n11061) );
  AND2_X1 U13596 ( .A1(n11062), .A2(n11061), .ZN(n11346) );
  OAI22_X1 U13597 ( .A1(n14822), .A2(n11346), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14905), .ZN(n11063) );
  AOI21_X1 U13598 ( .B1(n11064), .B2(n13174), .A(n11063), .ZN(n11065) );
  OAI211_X1 U13599 ( .C1(n11348), .C2(n13133), .A(n11066), .B(n11065), .ZN(
        P2_U3189) );
  INV_X1 U13600 ( .A(n11067), .ZN(n11070) );
  OAI222_X1 U13601 ( .A1(n14216), .A2(n11068), .B1(n14225), .B2(n11070), .C1(
        P1_U3086), .C2(n13895), .ZN(P1_U3337) );
  INV_X1 U13602 ( .A(n13265), .ZN(n13269) );
  OAI222_X1 U13603 ( .A1(n13269), .A2(P2_U3088), .B1(n13708), .B2(n11070), 
        .C1(n11069), .C2(n13705), .ZN(P2_U3309) );
  INV_X1 U13604 ( .A(n14107), .ZN(n14527) );
  XNOR2_X1 U13605 ( .A(n14749), .B(n14598), .ZN(n12276) );
  XNOR2_X1 U13606 ( .A(n11071), .B(n12276), .ZN(n14752) );
  OAI211_X1 U13607 ( .C1(n14728), .C2(n14749), .A(n14705), .B(n14726), .ZN(
        n14748) );
  INV_X1 U13608 ( .A(n14719), .ZN(n14702) );
  INV_X1 U13609 ( .A(n11072), .ZN(n11073) );
  AOI22_X1 U13610 ( .A1(n14723), .A2(n12110), .B1(n14702), .B2(n11073), .ZN(
        n11074) );
  OAI21_X1 U13611 ( .B1(n14088), .B2(n14748), .A(n11074), .ZN(n11081) );
  INV_X1 U13612 ( .A(n12276), .ZN(n11075) );
  XNOR2_X1 U13613 ( .A(n11076), .B(n11075), .ZN(n11077) );
  NAND2_X1 U13614 ( .A1(n11077), .A2(n14716), .ZN(n11079) );
  NAND2_X1 U13615 ( .A1(n11079), .A2(n11078), .ZN(n14750) );
  MUX2_X1 U13616 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n14750), .S(n14721), .Z(
        n11080) );
  AOI211_X1 U13617 ( .C1(n14527), .C2(n14752), .A(n11081), .B(n11080), .ZN(
        n11082) );
  INV_X1 U13618 ( .A(n11082), .ZN(P1_U3289) );
  INV_X1 U13619 ( .A(n11083), .ZN(n11090) );
  AOI22_X1 U13620 ( .A1(n13517), .A2(P2_REG2_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n13511), .ZN(n11084) );
  OAI21_X1 U13621 ( .B1(n6909), .B2(n13461), .A(n11084), .ZN(n11085) );
  AOI21_X1 U13622 ( .B1(n13529), .B2(n11086), .A(n11085), .ZN(n11089) );
  NAND2_X1 U13623 ( .A1(n11087), .A2(n13519), .ZN(n11088) );
  OAI211_X1 U13624 ( .C1(n13467), .C2(n11090), .A(n11089), .B(n11088), .ZN(
        P2_U3263) );
  INV_X1 U13625 ( .A(n11091), .ZN(n11099) );
  INV_X1 U13626 ( .A(n11092), .ZN(n11093) );
  MUX2_X1 U13627 ( .A(n11094), .B(n11093), .S(n13519), .Z(n11098) );
  OAI22_X1 U13628 ( .A1(n13461), .A2(n11223), .B1(n11219), .B2(n13521), .ZN(
        n11095) );
  AOI21_X1 U13629 ( .B1(n11096), .B2(n13529), .A(n11095), .ZN(n11097) );
  OAI211_X1 U13630 ( .C1(n13467), .C2(n11099), .A(n11098), .B(n11097), .ZN(
        P2_U3261) );
  INV_X1 U13631 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11100) );
  MUX2_X1 U13632 ( .A(n11100), .B(P2_REG1_REG_13__SCAN_IN), .S(n11482), .Z(
        n11104) );
  OAI21_X1 U13633 ( .B1(n11102), .B2(P2_REG1_REG_12__SCAN_IN), .A(n11101), 
        .ZN(n11103) );
  AOI211_X1 U13634 ( .C1(n11104), .C2(n11103), .A(n14932), .B(n11481), .ZN(
        n11113) );
  AOI21_X1 U13635 ( .B1(n11584), .B2(n11106), .A(n11105), .ZN(n11108) );
  MUX2_X1 U13636 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n11669), .S(n11482), .Z(
        n11107) );
  NAND2_X1 U13637 ( .A1(n11108), .A2(n11107), .ZN(n11476) );
  OAI211_X1 U13638 ( .C1(n11108), .C2(n11107), .A(n11476), .B(n14941), .ZN(
        n11111) );
  NOR2_X1 U13639 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14820), .ZN(n11109) );
  AOI21_X1 U13640 ( .B1(n14924), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n11109), 
        .ZN(n11110) );
  OAI211_X1 U13641 ( .C1(n14930), .C2(n11477), .A(n11111), .B(n11110), .ZN(
        n11112) );
  OR2_X1 U13642 ( .A1(n11113), .A2(n11112), .ZN(P2_U3227) );
  XOR2_X1 U13643 ( .A(n11114), .B(n11120), .Z(n14970) );
  INV_X1 U13644 ( .A(n14970), .ZN(n11128) );
  XNOR2_X1 U13645 ( .A(n11115), .B(n12350), .ZN(n11117) );
  NAND2_X1 U13646 ( .A1(n11117), .A2(n11269), .ZN(n14966) );
  INV_X1 U13647 ( .A(n14966), .ZN(n11119) );
  OAI22_X1 U13648 ( .A1(n13461), .A2(n12350), .B1(n13521), .B2(n12347), .ZN(
        n11118) );
  AOI21_X1 U13649 ( .B1(n13529), .B2(n11119), .A(n11118), .ZN(n11127) );
  XNOR2_X1 U13650 ( .A(n11121), .B(n11120), .ZN(n11124) );
  NAND2_X1 U13651 ( .A1(n13173), .A2(n13203), .ZN(n11123) );
  NAND2_X1 U13652 ( .A1(n13172), .A2(n13205), .ZN(n11122) );
  NAND2_X1 U13653 ( .A1(n11123), .A2(n11122), .ZN(n12348) );
  AOI21_X1 U13654 ( .B1(n11124), .B2(n13484), .A(n12348), .ZN(n14967) );
  MUX2_X1 U13655 ( .A(n11125), .B(n14967), .S(n13519), .Z(n11126) );
  OAI211_X1 U13656 ( .C1(n11128), .C2(n13467), .A(n11127), .B(n11126), .ZN(
        P2_U3260) );
  INV_X1 U13657 ( .A(n11129), .ZN(n11139) );
  OAI22_X1 U13658 ( .A1(n13461), .A2(n11131), .B1(n11130), .B2(n13521), .ZN(
        n11132) );
  AOI21_X1 U13659 ( .B1(n13529), .B2(n11133), .A(n11132), .ZN(n11138) );
  INV_X1 U13660 ( .A(n11134), .ZN(n11136) );
  MUX2_X1 U13661 ( .A(n11136), .B(n11135), .S(n13517), .Z(n11137) );
  OAI211_X1 U13662 ( .C1(n13467), .C2(n11139), .A(n11138), .B(n11137), .ZN(
        P2_U3264) );
  INV_X1 U13663 ( .A(n13167), .ZN(n13140) );
  OAI22_X1 U13664 ( .A1(n13140), .A2(n11140), .B1(n11146), .B2(n14824), .ZN(
        n11142) );
  NAND2_X1 U13665 ( .A1(n11142), .A2(n11141), .ZN(n11145) );
  AOI22_X1 U13666 ( .A1(n13159), .A2(n11143), .B1(n11161), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n11144) );
  OAI211_X1 U13667 ( .C1(n13133), .C2(n11146), .A(n11145), .B(n11144), .ZN(
        P2_U3204) );
  NAND2_X1 U13668 ( .A1(n12563), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n11147) );
  OAI21_X1 U13669 ( .B1(n12405), .B2(n12563), .A(n11147), .ZN(P3_U3520) );
  NAND2_X1 U13670 ( .A1(n12563), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n11148) );
  OAI21_X1 U13671 ( .B1(n11149), .B2(n12563), .A(n11148), .ZN(P3_U3521) );
  NAND2_X1 U13672 ( .A1(n11151), .A2(n11150), .ZN(n11153) );
  OAI211_X1 U13673 ( .C1(n11154), .C2(n11761), .A(n11153), .B(n11152), .ZN(
        P3_U3272) );
  OAI22_X1 U13674 ( .A1(n13140), .A2(n11156), .B1(n11155), .B2(n14824), .ZN(
        n11160) );
  INV_X1 U13675 ( .A(n11157), .ZN(n11159) );
  NAND3_X1 U13676 ( .A1(n11160), .A2(n11159), .A3(n11158), .ZN(n11168) );
  INV_X1 U13677 ( .A(n11161), .ZN(n11163) );
  OAI22_X1 U13678 ( .A1(n14822), .A2(n11164), .B1(n11163), .B2(n11162), .ZN(
        n11165) );
  AOI21_X1 U13679 ( .B1(n11166), .B2(n14829), .A(n11165), .ZN(n11167) );
  OAI211_X1 U13680 ( .C1(n14824), .C2(n11169), .A(n11168), .B(n11167), .ZN(
        P2_U3209) );
  INV_X1 U13681 ( .A(n11188), .ZN(n11173) );
  NOR3_X1 U13682 ( .A1(n13140), .A2(n11171), .A3(n11170), .ZN(n11172) );
  AOI21_X1 U13683 ( .B1(n11173), .B2(n13148), .A(n11172), .ZN(n11183) );
  NAND2_X1 U13684 ( .A1(n13172), .A2(n13202), .ZN(n11175) );
  NAND2_X1 U13685 ( .A1(n13173), .A2(n13200), .ZN(n11174) );
  AND2_X1 U13686 ( .A1(n11175), .A2(n11174), .ZN(n11426) );
  INV_X1 U13687 ( .A(n11426), .ZN(n11176) );
  NAND2_X1 U13688 ( .A1(n13159), .A2(n11176), .ZN(n11177) );
  NAND2_X1 U13689 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n14893) );
  OAI211_X1 U13690 ( .C1(n14832), .C2(n11430), .A(n11177), .B(n14893), .ZN(
        n11179) );
  NOR2_X1 U13691 ( .A1(n11260), .A2(n14824), .ZN(n11178) );
  AOI211_X1 U13692 ( .C1(n11180), .C2(n14829), .A(n11179), .B(n11178), .ZN(
        n11181) );
  OAI21_X1 U13693 ( .B1(n11183), .B2(n11182), .A(n11181), .ZN(P2_U3193) );
  INV_X1 U13694 ( .A(n11184), .ZN(n11185) );
  AOI21_X1 U13695 ( .B1(n11186), .B2(n11185), .A(n14824), .ZN(n11190) );
  NOR3_X1 U13696 ( .A1(n13140), .A2(n11191), .A3(n11187), .ZN(n11189) );
  OAI21_X1 U13697 ( .B1(n11190), .B2(n11189), .A(n11188), .ZN(n11196) );
  INV_X1 U13698 ( .A(n11306), .ZN(n11194) );
  OAI22_X1 U13699 ( .A1(n11256), .A2(n13136), .B1(n11191), .B2(n13135), .ZN(
        n11299) );
  INV_X1 U13700 ( .A(n11299), .ZN(n11192) );
  INV_X1 U13701 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n11914) );
  OAI22_X1 U13702 ( .A1(n14822), .A2(n11192), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11914), .ZN(n11193) );
  AOI21_X1 U13703 ( .B1(n11194), .B2(n13174), .A(n11193), .ZN(n11195) );
  OAI211_X1 U13704 ( .C1(n14980), .C2(n13133), .A(n11196), .B(n11195), .ZN(
        P2_U3185) );
  XNOR2_X1 U13705 ( .A(n11197), .B(n11201), .ZN(n14779) );
  INV_X1 U13706 ( .A(n14779), .ZN(n11211) );
  INV_X1 U13707 ( .A(n11198), .ZN(n11199) );
  AOI211_X1 U13708 ( .C1(n11201), .C2(n11200), .A(n14691), .B(n11199), .ZN(
        n14777) );
  NAND2_X1 U13709 ( .A1(n13856), .A2(n14596), .ZN(n11203) );
  NAND2_X1 U13710 ( .A1(n13854), .A2(n14498), .ZN(n11202) );
  AND2_X1 U13711 ( .A1(n11203), .A2(n11202), .ZN(n14774) );
  INV_X1 U13712 ( .A(n14774), .ZN(n11204) );
  OAI21_X1 U13713 ( .B1(n14777), .B2(n11204), .A(n14721), .ZN(n11210) );
  OAI22_X1 U13714 ( .A1(n14721), .A2(n11206), .B1(n11205), .B2(n14719), .ZN(
        n11208) );
  OAI211_X1 U13715 ( .C1(n14682), .C2(n14776), .A(n14726), .B(n14667), .ZN(
        n14775) );
  NOR2_X1 U13716 ( .A1(n14775), .A2(n14088), .ZN(n11207) );
  AOI211_X1 U13717 ( .C1(n14723), .C2(n12127), .A(n11208), .B(n11207), .ZN(
        n11209) );
  OAI211_X1 U13718 ( .C1(n11211), .C2(n14107), .A(n11210), .B(n11209), .ZN(
        P1_U3285) );
  INV_X1 U13719 ( .A(n11212), .ZN(n14813) );
  NOR3_X1 U13720 ( .A1(n13140), .A2(n11214), .A3(n11213), .ZN(n11215) );
  AOI21_X1 U13721 ( .B1(n13148), .B2(n14813), .A(n11215), .ZN(n11227) );
  INV_X1 U13722 ( .A(n11216), .ZN(n12354) );
  INV_X1 U13723 ( .A(n11217), .ZN(n11218) );
  AOI22_X1 U13724 ( .A1(n13159), .A2(n11218), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11222) );
  INV_X1 U13725 ( .A(n11219), .ZN(n11220) );
  NAND2_X1 U13726 ( .A1(n13174), .A2(n11220), .ZN(n11221) );
  OAI211_X1 U13727 ( .C1(n11223), .C2(n13133), .A(n11222), .B(n11221), .ZN(
        n11224) );
  AOI21_X1 U13728 ( .B1(n12354), .B2(n13148), .A(n11224), .ZN(n11225) );
  OAI21_X1 U13729 ( .B1(n11227), .B2(n11226), .A(n11225), .ZN(P2_U3202) );
  NAND2_X1 U13730 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n11771)
         );
  INV_X1 U13731 ( .A(n11771), .ZN(n11228) );
  AOI21_X1 U13732 ( .B1(n14615), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n11228), 
        .ZN(n11229) );
  INV_X1 U13733 ( .A(n11229), .ZN(n11235) );
  OAI21_X1 U13734 ( .B1(n11236), .B2(P1_REG1_REG_12__SCAN_IN), .A(n11230), 
        .ZN(n11233) );
  INV_X1 U13735 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11231) );
  MUX2_X1 U13736 ( .A(n11231), .B(P1_REG1_REG_13__SCAN_IN), .S(n11375), .Z(
        n11232) );
  NOR2_X1 U13737 ( .A1(n11233), .A2(n11232), .ZN(n11374) );
  AOI211_X1 U13738 ( .C1(n11233), .C2(n11232), .A(n11374), .B(n13911), .ZN(
        n11234) );
  AOI211_X1 U13739 ( .C1(n14645), .C2(n11375), .A(n11235), .B(n11234), .ZN(
        n11243) );
  NOR2_X1 U13740 ( .A1(n11236), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11238) );
  NOR2_X1 U13741 ( .A1(n11238), .A2(n11237), .ZN(n11241) );
  MUX2_X1 U13742 ( .A(n11655), .B(P1_REG2_REG_13__SCAN_IN), .S(n11375), .Z(
        n11239) );
  INV_X1 U13743 ( .A(n11239), .ZN(n11240) );
  NAND2_X1 U13744 ( .A1(n11240), .A2(n11241), .ZN(n11369) );
  OAI211_X1 U13745 ( .C1(n11241), .C2(n11240), .A(n14649), .B(n11369), .ZN(
        n11242) );
  NAND2_X1 U13746 ( .A1(n11243), .A2(n11242), .ZN(P1_U3256) );
  INV_X1 U13747 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n11245) );
  NAND2_X1 U13748 ( .A1(n12739), .A2(P3_U3897), .ZN(n11244) );
  OAI21_X1 U13749 ( .B1(P3_U3897), .B2(n11245), .A(n11244), .ZN(P3_U3517) );
  INV_X1 U13750 ( .A(n11246), .ZN(n11248) );
  OAI222_X1 U13751 ( .A1(n13276), .A2(P2_U3088), .B1(n13708), .B2(n11248), 
        .C1(n11247), .C2(n13705), .ZN(P2_U3308) );
  OAI222_X1 U13752 ( .A1(n14216), .A2(n11249), .B1(n14225), .B2(n11248), .C1(
        n13915), .C2(P1_U3086), .ZN(P1_U3336) );
  NOR2_X1 U13753 ( .A1(n14832), .A2(n11507), .ZN(n11254) );
  NAND2_X1 U13754 ( .A1(n13172), .A2(n13201), .ZN(n11251) );
  NAND2_X1 U13755 ( .A1(n13173), .A2(n13199), .ZN(n11250) );
  AND2_X1 U13756 ( .A1(n11251), .A2(n11250), .ZN(n11361) );
  OAI21_X1 U13757 ( .B1(n14822), .B2(n11361), .A(n11252), .ZN(n11253) );
  AOI211_X1 U13758 ( .C1(n11363), .C2(n14829), .A(n11254), .B(n11253), .ZN(
        n11262) );
  INV_X1 U13759 ( .A(n11255), .ZN(n11259) );
  OAI22_X1 U13760 ( .A1(n11257), .A2(n14824), .B1(n11256), .B2(n13140), .ZN(
        n11258) );
  NAND3_X1 U13761 ( .A1(n11260), .A2(n11259), .A3(n11258), .ZN(n11261) );
  OAI211_X1 U13762 ( .C1(n11263), .C2(n14824), .A(n11262), .B(n11261), .ZN(
        P2_U3203) );
  XNOR2_X1 U13763 ( .A(n13526), .B(n6469), .ZN(n11266) );
  NAND2_X1 U13764 ( .A1(n13198), .A2(n13490), .ZN(n11267) );
  XNOR2_X1 U13765 ( .A(n11266), .B(n11267), .ZN(n12423) );
  AND2_X1 U13766 ( .A1(n12423), .A2(n11264), .ZN(n11265) );
  INV_X1 U13767 ( .A(n11266), .ZN(n11277) );
  NAND2_X1 U13768 ( .A1(n11277), .A2(n11267), .ZN(n11268) );
  XNOR2_X1 U13769 ( .A(n11741), .B(n6469), .ZN(n11553) );
  NAND2_X1 U13770 ( .A1(n13197), .A2(n13490), .ZN(n11554) );
  XNOR2_X1 U13771 ( .A(n11553), .B(n11554), .ZN(n11275) );
  NOR2_X1 U13772 ( .A1(n14832), .A2(n11583), .ZN(n11274) );
  NAND2_X1 U13773 ( .A1(n13173), .A2(n11566), .ZN(n11271) );
  NAND2_X1 U13774 ( .A1(n13172), .A2(n13198), .ZN(n11270) );
  AND2_X1 U13775 ( .A1(n11271), .A2(n11270), .ZN(n11579) );
  OAI21_X1 U13776 ( .B1(n14822), .B2(n11579), .A(n11272), .ZN(n11273) );
  AOI211_X1 U13777 ( .C1(n11741), .C2(n14829), .A(n11274), .B(n11273), .ZN(
        n11281) );
  INV_X1 U13778 ( .A(n11275), .ZN(n11279) );
  OAI22_X1 U13779 ( .A1(n11277), .A2(n14824), .B1(n11276), .B2(n13140), .ZN(
        n11278) );
  NAND3_X1 U13780 ( .A1(n12432), .A2(n11279), .A3(n11278), .ZN(n11280) );
  OAI211_X1 U13781 ( .C1(n11557), .C2(n14824), .A(n11281), .B(n11280), .ZN(
        P2_U3196) );
  OAI21_X1 U13782 ( .B1(n6665), .B2(n11283), .A(n11282), .ZN(n11285) );
  AOI21_X1 U13783 ( .B1(n11285), .B2(n13484), .A(n11284), .ZN(n14974) );
  MUX2_X1 U13784 ( .A(n11286), .B(n14974), .S(n13519), .Z(n11296) );
  XNOR2_X1 U13785 ( .A(n11287), .B(n11288), .ZN(n14977) );
  INV_X1 U13786 ( .A(n11289), .ZN(n11291) );
  INV_X1 U13787 ( .A(n11305), .ZN(n11290) );
  OAI211_X1 U13788 ( .C1(n14975), .C2(n11291), .A(n11290), .B(n11269), .ZN(
        n14973) );
  NOR2_X1 U13789 ( .A1(n14973), .A2(n13498), .ZN(n11294) );
  OAI22_X1 U13790 ( .A1(n13461), .A2(n14975), .B1(n13521), .B2(n11292), .ZN(
        n11293) );
  AOI211_X1 U13791 ( .C1(n14977), .C2(n13527), .A(n11294), .B(n11293), .ZN(
        n11295) );
  NAND2_X1 U13792 ( .A1(n11296), .A2(n11295), .ZN(P2_U3259) );
  XNOR2_X1 U13793 ( .A(n11298), .B(n11297), .ZN(n11300) );
  AOI21_X1 U13794 ( .B1(n11300), .B2(n13484), .A(n11299), .ZN(n14979) );
  MUX2_X1 U13795 ( .A(n11301), .B(n14979), .S(n13519), .Z(n11310) );
  XNOR2_X1 U13796 ( .A(n11302), .B(n11303), .ZN(n14983) );
  INV_X1 U13797 ( .A(n11429), .ZN(n11304) );
  OAI211_X1 U13798 ( .C1(n14980), .C2(n11305), .A(n11304), .B(n11269), .ZN(
        n14978) );
  NOR2_X1 U13799 ( .A1(n14978), .A2(n13498), .ZN(n11308) );
  OAI22_X1 U13800 ( .A1(n13461), .A2(n14980), .B1(n13521), .B2(n11306), .ZN(
        n11307) );
  AOI211_X1 U13801 ( .C1(n14983), .C2(n13527), .A(n11308), .B(n11307), .ZN(
        n11309) );
  NAND2_X1 U13802 ( .A1(n11310), .A2(n11309), .ZN(P2_U3258) );
  XNOR2_X1 U13803 ( .A(n12386), .B(n11459), .ZN(n11409) );
  XNOR2_X1 U13804 ( .A(n11409), .B(n12560), .ZN(n11326) );
  AOI21_X1 U13805 ( .B1(n15207), .B2(n11314), .A(n11465), .ZN(n11312) );
  NAND2_X1 U13806 ( .A1(n11313), .A2(n7488), .ZN(n11324) );
  INV_X1 U13807 ( .A(n11314), .ZN(n11315) );
  NAND2_X1 U13808 ( .A1(n11315), .A2(n12562), .ZN(n11334) );
  NOR2_X1 U13809 ( .A1(n11317), .A2(n11334), .ZN(n11319) );
  OAI21_X1 U13810 ( .B1(n11317), .B2(n11316), .A(n11465), .ZN(n11318) );
  OAI21_X1 U13811 ( .B1(n11319), .B2(n11465), .A(n11318), .ZN(n11322) );
  INV_X1 U13812 ( .A(n11320), .ZN(n11321) );
  AOI21_X1 U13813 ( .B1(n11326), .B2(n11325), .A(n11411), .ZN(n11333) );
  AOI22_X1 U13814 ( .A1(n12548), .A2(n11327), .B1(n12545), .B2(n12559), .ZN(
        n11330) );
  NOR2_X1 U13815 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11328), .ZN(n15085) );
  AOI21_X1 U13816 ( .B1(n12522), .B2(n12561), .A(n15085), .ZN(n11329) );
  OAI211_X1 U13817 ( .C1(n14379), .C2(n11460), .A(n11330), .B(n11329), .ZN(
        n11331) );
  INV_X1 U13818 ( .A(n11331), .ZN(n11332) );
  OAI21_X1 U13819 ( .B1(n11333), .B2(n12550), .A(n11332), .ZN(P3_U3171) );
  NAND2_X1 U13820 ( .A1(n11335), .A2(n11334), .ZN(n11466) );
  XNOR2_X1 U13821 ( .A(n11466), .B(n11465), .ZN(n11340) );
  AOI22_X1 U13822 ( .A1(n12548), .A2(n11336), .B1(n12545), .B2(n12561), .ZN(
        n11338) );
  AOI22_X1 U13823 ( .A1(n12522), .A2(n12562), .B1(P3_REG3_REG_7__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11337) );
  OAI211_X1 U13824 ( .C1(n14379), .C2(n11392), .A(n11338), .B(n11337), .ZN(
        n11339) );
  AOI21_X1 U13825 ( .B1(n11340), .B2(n14376), .A(n11339), .ZN(n11341) );
  INV_X1 U13826 ( .A(n11341), .ZN(P3_U3153) );
  XNOR2_X1 U13827 ( .A(n11342), .B(n11344), .ZN(n11491) );
  INV_X1 U13828 ( .A(n11491), .ZN(n11354) );
  OAI211_X1 U13829 ( .C1(n11345), .C2(n11344), .A(n11343), .B(n13484), .ZN(
        n11347) );
  NAND2_X1 U13830 ( .A1(n11347), .A2(n11346), .ZN(n11489) );
  NAND2_X1 U13831 ( .A1(n11489), .A2(n13519), .ZN(n11353) );
  AOI211_X1 U13832 ( .C1(n11493), .C2(n11357), .A(n13490), .B(n11598), .ZN(
        n11490) );
  NOR2_X1 U13833 ( .A1(n11348), .A2(n13461), .ZN(n11351) );
  OAI22_X1 U13834 ( .A1(n13519), .A2(n10738), .B1(n11349), .B2(n13521), .ZN(
        n11350) );
  AOI211_X1 U13835 ( .C1(n11490), .C2(n13529), .A(n11351), .B(n11350), .ZN(
        n11352) );
  OAI211_X1 U13836 ( .C1(n11354), .C2(n13467), .A(n11353), .B(n11352), .ZN(
        P2_U3255) );
  XNOR2_X1 U13837 ( .A(n11355), .B(n7204), .ZN(n11504) );
  INV_X1 U13838 ( .A(n11357), .ZN(n11358) );
  AOI211_X1 U13839 ( .C1(n11363), .C2(n11356), .A(n13490), .B(n11358), .ZN(
        n11510) );
  OAI211_X1 U13840 ( .C1(n11360), .C2(n7204), .A(n11359), .B(n13484), .ZN(
        n11362) );
  NAND2_X1 U13841 ( .A1(n11362), .A2(n11361), .ZN(n11505) );
  AOI211_X1 U13842 ( .C1(n14982), .C2(n11504), .A(n11510), .B(n11505), .ZN(
        n11368) );
  INV_X1 U13843 ( .A(n11363), .ZN(n11506) );
  OAI22_X1 U13844 ( .A1(n13630), .A2(n11506), .B1(n15002), .B2(n10087), .ZN(
        n11364) );
  INV_X1 U13845 ( .A(n11364), .ZN(n11365) );
  OAI21_X1 U13846 ( .B1(n11368), .B2(n6478), .A(n11365), .ZN(P2_U3508) );
  OAI22_X1 U13847 ( .A1(n13677), .A2(n11506), .B1(n14995), .B2(n9225), .ZN(
        n11366) );
  INV_X1 U13848 ( .A(n11366), .ZN(n11367) );
  OAI21_X1 U13849 ( .B1(n11368), .B2(n14994), .A(n11367), .ZN(P2_U3457) );
  NAND2_X1 U13850 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n11375), .ZN(n11370) );
  NAND2_X1 U13851 ( .A1(n11370), .A2(n11369), .ZN(n11372) );
  MUX2_X1 U13852 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n14119), .S(n11781), .Z(
        n11371) );
  NAND2_X1 U13853 ( .A1(n11371), .A2(n11372), .ZN(n11790) );
  OAI211_X1 U13854 ( .C1(n11372), .C2(n11371), .A(n14649), .B(n11790), .ZN(
        n11383) );
  MUX2_X1 U13855 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n11373), .S(n11781), .Z(
        n11377) );
  OAI21_X1 U13856 ( .B1(n11377), .B2(n11376), .A(n11780), .ZN(n11381) );
  NAND2_X1 U13857 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n13716)
         );
  INV_X1 U13858 ( .A(n13716), .ZN(n11378) );
  AOI21_X1 U13859 ( .B1(n14615), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n11378), 
        .ZN(n11379) );
  OAI21_X1 U13860 ( .B1(n14634), .B2(n11791), .A(n11379), .ZN(n11380) );
  AOI21_X1 U13861 ( .B1(n14648), .B2(n11381), .A(n11380), .ZN(n11382) );
  NAND2_X1 U13862 ( .A1(n11383), .A2(n11382), .ZN(P1_U3257) );
  XNOR2_X1 U13863 ( .A(n11384), .B(n11386), .ZN(n15298) );
  AOI22_X1 U13864 ( .A1(n12561), .A2(n15259), .B1(n15256), .B2(n12562), .ZN(
        n11389) );
  OAI211_X1 U13865 ( .C1(n11387), .C2(n11386), .A(n11385), .B(n15262), .ZN(
        n11388) );
  OAI211_X1 U13866 ( .C1(n15298), .C2(n15266), .A(n11389), .B(n11388), .ZN(
        n15299) );
  INV_X1 U13867 ( .A(n15299), .ZN(n11390) );
  MUX2_X1 U13868 ( .A(n11390), .B(n12624), .S(n12719), .Z(n11395) );
  NOR2_X1 U13869 ( .A1(n11391), .A2(n15253), .ZN(n15300) );
  INV_X1 U13870 ( .A(n11392), .ZN(n11393) );
  AOI22_X1 U13871 ( .A1(n15227), .A2(n15300), .B1(n15226), .B2(n11393), .ZN(
        n11394) );
  OAI211_X1 U13872 ( .C1(n15298), .C2(n15270), .A(n11395), .B(n11394), .ZN(
        P3_U3226) );
  XOR2_X1 U13873 ( .A(n11397), .B(n11396), .Z(n11401) );
  AOI22_X1 U13874 ( .A1(n15256), .A2(n15190), .B1(n12560), .B2(n15259), .ZN(
        n11400) );
  XNOR2_X1 U13875 ( .A(n11398), .B(n11397), .ZN(n15305) );
  INV_X1 U13876 ( .A(n15266), .ZN(n15246) );
  NAND2_X1 U13877 ( .A1(n15305), .A2(n15246), .ZN(n11399) );
  OAI211_X1 U13878 ( .C1(n11401), .C2(n15249), .A(n11400), .B(n11399), .ZN(
        n15303) );
  INV_X1 U13879 ( .A(n15303), .ZN(n11407) );
  INV_X1 U13880 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n12622) );
  NOR2_X1 U13881 ( .A1(n11402), .A2(n15253), .ZN(n15304) );
  AOI22_X1 U13882 ( .A1(n15227), .A2(n15304), .B1(n15226), .B2(n11403), .ZN(
        n11404) );
  OAI21_X1 U13883 ( .B1(n12622), .B2(n15273), .A(n11404), .ZN(n11405) );
  AOI21_X1 U13884 ( .B1(n15305), .B2(n11530), .A(n11405), .ZN(n11406) );
  OAI21_X1 U13885 ( .B1(n11407), .B2(n12719), .A(n11406), .ZN(P3_U3225) );
  XNOR2_X1 U13886 ( .A(n12386), .B(n11408), .ZN(n11639) );
  XNOR2_X1 U13887 ( .A(n11639), .B(n14453), .ZN(n11412) );
  NOR2_X1 U13888 ( .A1(n11409), .A2(n12560), .ZN(n11413) );
  OAI21_X1 U13889 ( .B1(n11411), .B2(n11413), .A(n11412), .ZN(n11414) );
  NAND3_X1 U13890 ( .A1(n6667), .A2(n14376), .A3(n11414), .ZN(n11418) );
  NAND2_X1 U13891 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n15099)
         );
  INV_X1 U13892 ( .A(n15099), .ZN(n11416) );
  OAI22_X1 U13893 ( .A1(n14373), .A2(n11524), .B1(n12507), .B2(n11727), .ZN(
        n11415) );
  AOI211_X1 U13894 ( .C1(n12522), .C2(n12560), .A(n11416), .B(n11415), .ZN(
        n11417) );
  OAI211_X1 U13895 ( .C1(n11525), .C2(n14379), .A(n11418), .B(n11417), .ZN(
        P3_U3157) );
  INV_X1 U13896 ( .A(n11419), .ZN(n11421) );
  OAI21_X1 U13897 ( .B1(n11421), .B2(n11422), .A(n11420), .ZN(n14985) );
  NAND2_X1 U13898 ( .A1(n11423), .A2(n11422), .ZN(n11424) );
  NAND3_X1 U13899 ( .A1(n11425), .A2(n13484), .A3(n11424), .ZN(n11427) );
  NAND2_X1 U13900 ( .A1(n11427), .A2(n11426), .ZN(n14992) );
  INV_X1 U13901 ( .A(n14992), .ZN(n11428) );
  MUX2_X1 U13902 ( .A(n11428), .B(n10104), .S(n13517), .Z(n11434) );
  OAI211_X1 U13903 ( .C1(n11429), .C2(n14990), .A(n11269), .B(n11356), .ZN(
        n14988) );
  INV_X1 U13904 ( .A(n14988), .ZN(n11432) );
  OAI22_X1 U13905 ( .A1(n14990), .A2(n13461), .B1(n11430), .B2(n13521), .ZN(
        n11431) );
  AOI21_X1 U13906 ( .B1(n11432), .B2(n13529), .A(n11431), .ZN(n11433) );
  OAI211_X1 U13907 ( .C1(n13467), .C2(n14985), .A(n11434), .B(n11433), .ZN(
        P2_U3257) );
  NAND2_X1 U13908 ( .A1(n12438), .A2(P3_U3897), .ZN(n11435) );
  OAI21_X1 U13909 ( .B1(P3_U3897), .B2(n11436), .A(n11435), .ZN(P3_U3519) );
  INV_X1 U13910 ( .A(n14665), .ZN(n14782) );
  NAND2_X1 U13911 ( .A1(n11438), .A2(n11437), .ZN(n11439) );
  AOI22_X1 U13912 ( .A1(n14665), .A2(n12028), .B1(n12039), .B2(n13854), .ZN(
        n11677) );
  INV_X1 U13913 ( .A(n11677), .ZN(n11441) );
  AOI22_X1 U13914 ( .A1(n14665), .A2(n12035), .B1(n6542), .B2(n13854), .ZN(
        n11442) );
  XOR2_X1 U13915 ( .A(n12332), .B(n11442), .Z(n11443) );
  OAI211_X1 U13916 ( .C1(n11444), .C2(n11443), .A(n11680), .B(n14488), .ZN(
        n11449) );
  INV_X1 U13917 ( .A(n14606), .ZN(n13834) );
  INV_X1 U13918 ( .A(n11445), .ZN(n14664) );
  AOI22_X1 U13919 ( .A1(n14596), .A2(n13855), .B1(n13853), .B2(n14597), .ZN(
        n14657) );
  OAI21_X1 U13920 ( .B1(n14657), .B2(n13836), .A(n11446), .ZN(n11447) );
  AOI21_X1 U13921 ( .B1(n13834), .B2(n14664), .A(n11447), .ZN(n11448) );
  OAI211_X1 U13922 ( .C1(n14782), .C2(n13817), .A(n11449), .B(n11448), .ZN(
        P1_U3231) );
  XNOR2_X1 U13923 ( .A(n11450), .B(n11455), .ZN(n15307) );
  NAND2_X1 U13924 ( .A1(n12559), .A2(n15259), .ZN(n11451) );
  OAI21_X1 U13925 ( .B1(n11452), .B2(n15243), .A(n11451), .ZN(n11453) );
  AOI21_X1 U13926 ( .B1(n15307), .B2(n15246), .A(n11453), .ZN(n11458) );
  XNOR2_X1 U13927 ( .A(n11454), .B(n11455), .ZN(n11456) );
  NAND2_X1 U13928 ( .A1(n11456), .A2(n15262), .ZN(n11457) );
  AND2_X1 U13929 ( .A1(n11458), .A2(n11457), .ZN(n15309) );
  NOR2_X1 U13930 ( .A1(n11459), .A2(n15253), .ZN(n15306) );
  INV_X1 U13931 ( .A(n11460), .ZN(n11461) );
  AOI22_X1 U13932 ( .A1(n15227), .A2(n15306), .B1(n15226), .B2(n11461), .ZN(
        n11462) );
  OAI21_X1 U13933 ( .B1(n12620), .B2(n15273), .A(n11462), .ZN(n11463) );
  AOI21_X1 U13934 ( .B1(n15307), .B2(n11530), .A(n11463), .ZN(n11464) );
  OAI21_X1 U13935 ( .B1(n15309), .B2(n12719), .A(n11464), .ZN(P3_U3224) );
  MUX2_X1 U13936 ( .A(n11466), .B(n15190), .S(n11465), .Z(n11468) );
  XNOR2_X1 U13937 ( .A(n11468), .B(n11467), .ZN(n11475) );
  AOI22_X1 U13938 ( .A1(n12548), .A2(n7322), .B1(n12545), .B2(n12560), .ZN(
        n11471) );
  NAND2_X1 U13939 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n15074) );
  INV_X1 U13940 ( .A(n15074), .ZN(n11469) );
  AOI21_X1 U13941 ( .B1(n12522), .B2(n15190), .A(n11469), .ZN(n11470) );
  OAI211_X1 U13942 ( .C1(n14379), .C2(n11472), .A(n11471), .B(n11470), .ZN(
        n11473) );
  INV_X1 U13943 ( .A(n11473), .ZN(n11474) );
  OAI21_X1 U13944 ( .B1(n11475), .B2(n12550), .A(n11474), .ZN(P3_U3161) );
  OAI21_X1 U13945 ( .B1(n11669), .B2(n11477), .A(n11476), .ZN(n13223) );
  XNOR2_X1 U13946 ( .A(n13223), .B(n13238), .ZN(n13225) );
  XNOR2_X1 U13947 ( .A(n13225), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n11487) );
  NOR2_X1 U13948 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11567), .ZN(n11478) );
  AOI21_X1 U13949 ( .B1(n14924), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n11478), 
        .ZN(n11479) );
  OAI21_X1 U13950 ( .B1(n11480), .B2(n14930), .A(n11479), .ZN(n11486) );
  XNOR2_X1 U13951 ( .A(n13238), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n11483) );
  AOI211_X1 U13952 ( .C1(n11484), .C2(n11483), .A(n14932), .B(n13237), .ZN(
        n11485) );
  AOI211_X1 U13953 ( .C1(n14941), .C2(n11487), .A(n11486), .B(n11485), .ZN(
        n11488) );
  INV_X1 U13954 ( .A(n11488), .ZN(P2_U3228) );
  AOI211_X1 U13955 ( .C1(n14982), .C2(n11491), .A(n11490), .B(n11489), .ZN(
        n11495) );
  AOI22_X1 U13956 ( .A1(n13634), .A2(n11493), .B1(n6478), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n11492) );
  OAI21_X1 U13957 ( .B1(n11495), .B2(n6478), .A(n11492), .ZN(P2_U3509) );
  AOI22_X1 U13958 ( .A1(n13680), .A2(n11493), .B1(n14994), .B2(
        P2_REG0_REG_10__SCAN_IN), .ZN(n11494) );
  OAI21_X1 U13959 ( .B1(n11495), .B2(n14994), .A(n11494), .ZN(P2_U3460) );
  INV_X1 U13960 ( .A(n11496), .ZN(n11498) );
  INV_X1 U13961 ( .A(n13461), .ZN(n13525) );
  AOI22_X1 U13962 ( .A1(n13525), .A2(n14818), .B1(n9148), .B2(n13511), .ZN(
        n11497) );
  OAI21_X1 U13963 ( .B1(n11498), .B2(n13498), .A(n11497), .ZN(n11501) );
  MUX2_X1 U13964 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11499), .S(n13519), .Z(
        n11500) );
  AOI211_X1 U13965 ( .C1(n13527), .C2(n11502), .A(n11501), .B(n11500), .ZN(
        n11503) );
  INV_X1 U13966 ( .A(n11503), .ZN(P2_U3262) );
  INV_X1 U13967 ( .A(n11504), .ZN(n11513) );
  NAND2_X1 U13968 ( .A1(n11505), .A2(n13519), .ZN(n11512) );
  NOR2_X1 U13969 ( .A1(n11506), .A2(n13461), .ZN(n11509) );
  OAI22_X1 U13970 ( .A1(n13519), .A2(n10106), .B1(n11507), .B2(n13521), .ZN(
        n11508) );
  AOI211_X1 U13971 ( .C1(n11510), .C2(n13529), .A(n11509), .B(n11508), .ZN(
        n11511) );
  OAI211_X1 U13972 ( .C1(n11513), .C2(n13467), .A(n11512), .B(n11511), .ZN(
        P2_U3256) );
  XNOR2_X1 U13973 ( .A(n11514), .B(n11519), .ZN(n15313) );
  NAND2_X1 U13974 ( .A1(n12558), .A2(n15259), .ZN(n11516) );
  NAND2_X1 U13975 ( .A1(n12560), .A2(n15256), .ZN(n11515) );
  NAND2_X1 U13976 ( .A1(n11516), .A2(n11515), .ZN(n11517) );
  AOI21_X1 U13977 ( .B1(n15313), .B2(n15246), .A(n11517), .ZN(n11523) );
  INV_X1 U13978 ( .A(n11519), .ZN(n11520) );
  XNOR2_X1 U13979 ( .A(n11518), .B(n11520), .ZN(n11521) );
  NAND2_X1 U13980 ( .A1(n11521), .A2(n15262), .ZN(n11522) );
  NOR2_X1 U13981 ( .A1(n11524), .A2(n15253), .ZN(n15311) );
  INV_X1 U13982 ( .A(n11525), .ZN(n11526) );
  AOI22_X1 U13983 ( .A1(n15227), .A2(n15311), .B1(n15226), .B2(n11526), .ZN(
        n11527) );
  OAI21_X1 U13984 ( .B1(n11528), .B2(n15273), .A(n11527), .ZN(n11529) );
  AOI21_X1 U13985 ( .B1(n15313), .B2(n11530), .A(n11529), .ZN(n11531) );
  OAI21_X1 U13986 ( .B1(n15315), .B2(n12719), .A(n11531), .ZN(P3_U3223) );
  XNOR2_X1 U13987 ( .A(n11532), .B(n12284), .ZN(n14796) );
  INV_X1 U13988 ( .A(n14796), .ZN(n11544) );
  INV_X1 U13989 ( .A(n11533), .ZN(n11534) );
  AOI211_X1 U13990 ( .C1(n12284), .C2(n11535), .A(n14691), .B(n11534), .ZN(
        n14794) );
  NAND2_X1 U13991 ( .A1(n13854), .A2(n14596), .ZN(n14487) );
  INV_X1 U13992 ( .A(n14487), .ZN(n11536) );
  OAI21_X1 U13993 ( .B1(n14794), .B2(n11536), .A(n14721), .ZN(n11543) );
  NAND2_X1 U13994 ( .A1(n13852), .A2(n14498), .ZN(n14486) );
  INV_X1 U13995 ( .A(n14492), .ZN(n11537) );
  AOI22_X1 U13996 ( .A1(n14701), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n11537), 
        .B2(n14702), .ZN(n11538) );
  OAI21_X1 U13997 ( .B1(n14088), .B2(n14486), .A(n11538), .ZN(n11541) );
  XNOR2_X1 U13998 ( .A(n14668), .B(n14478), .ZN(n14793) );
  AND2_X1 U13999 ( .A1(n14731), .A2(n14726), .ZN(n13974) );
  INV_X1 U14000 ( .A(n13974), .ZN(n11539) );
  NOR2_X1 U14001 ( .A1(n14793), .A2(n11539), .ZN(n11540) );
  AOI211_X1 U14002 ( .C1(n14723), .C2(n14478), .A(n11541), .B(n11540), .ZN(
        n11542) );
  OAI211_X1 U14003 ( .C1(n11544), .C2(n14107), .A(n11543), .B(n11542), .ZN(
        P1_U3283) );
  INV_X1 U14004 ( .A(n11545), .ZN(n11551) );
  OAI222_X1 U14005 ( .A1(n14225), .A2(n11551), .B1(P1_U3086), .B2(n12255), 
        .C1(n11546), .C2(n14216), .ZN(P1_U3335) );
  INV_X1 U14006 ( .A(n11547), .ZN(n11549) );
  OAI222_X1 U14007 ( .A1(P3_U3151), .A2(n8985), .B1(n13021), .B2(n11549), .C1(
        n11548), .C2(n11761), .ZN(P3_U3271) );
  OAI222_X1 U14008 ( .A1(P2_U3088), .A2(n11552), .B1(n13708), .B2(n11551), 
        .C1(n11550), .C2(n13705), .ZN(P2_U3307) );
  INV_X1 U14009 ( .A(n11553), .ZN(n11555) );
  NAND2_X1 U14010 ( .A1(n11555), .A2(n11554), .ZN(n11556) );
  NAND2_X1 U14011 ( .A1(n11557), .A2(n11556), .ZN(n14825) );
  XNOR2_X1 U14012 ( .A(n14830), .B(n6469), .ZN(n11563) );
  AND2_X1 U14013 ( .A1(n11566), .A2(n13490), .ZN(n11558) );
  NAND2_X1 U14014 ( .A1(n11563), .A2(n11558), .ZN(n11702) );
  INV_X1 U14015 ( .A(n11563), .ZN(n11560) );
  INV_X1 U14016 ( .A(n11558), .ZN(n11559) );
  NAND2_X1 U14017 ( .A1(n11560), .A2(n11559), .ZN(n11561) );
  NAND2_X1 U14018 ( .A1(n11702), .A2(n11561), .ZN(n14826) );
  NAND2_X1 U14019 ( .A1(n13196), .A2(n13490), .ZN(n11703) );
  INV_X1 U14020 ( .A(n11701), .ZN(n11562) );
  XOR2_X1 U14021 ( .A(n11703), .B(n11562), .Z(n11571) );
  INV_X1 U14022 ( .A(n11804), .ZN(n11574) );
  NAND3_X1 U14023 ( .A1(n11563), .A2(n13167), .A3(n11566), .ZN(n11564) );
  OAI21_X1 U14024 ( .B1(n11699), .B2(n14824), .A(n11564), .ZN(n11572) );
  INV_X1 U14025 ( .A(n11565), .ZN(n13512) );
  AOI22_X1 U14026 ( .A1(n13172), .A2(n11566), .B1(n13173), .B2(n13195), .ZN(
        n13503) );
  OAI22_X1 U14027 ( .A1(n14822), .A2(n13503), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11567), .ZN(n11568) );
  AOI21_X1 U14028 ( .B1(n13512), .B2(n13174), .A(n11568), .ZN(n11569) );
  OAI21_X1 U14029 ( .B1(n13678), .B2(n13133), .A(n11569), .ZN(n11570) );
  AOI21_X1 U14030 ( .B1(n11572), .B2(n11571), .A(n11570), .ZN(n11573) );
  OAI21_X1 U14031 ( .B1(n11574), .B2(n14824), .A(n11573), .ZN(P2_U3187) );
  OAI21_X1 U14032 ( .B1(n11576), .B2(n9272), .A(n11575), .ZN(n11736) );
  INV_X1 U14033 ( .A(n11736), .ZN(n11589) );
  OAI211_X1 U14034 ( .C1(n6658), .C2(n11578), .A(n13484), .B(n11577), .ZN(
        n11580) );
  NAND2_X1 U14035 ( .A1(n11580), .A2(n11579), .ZN(n11734) );
  NAND2_X1 U14036 ( .A1(n11734), .A2(n13519), .ZN(n11588) );
  INV_X1 U14037 ( .A(n11599), .ZN(n11582) );
  INV_X1 U14038 ( .A(n11667), .ZN(n11581) );
  AOI211_X1 U14039 ( .C1(n11741), .C2(n11582), .A(n13490), .B(n11581), .ZN(
        n11735) );
  NOR2_X1 U14040 ( .A1(n11738), .A2(n13461), .ZN(n11586) );
  OAI22_X1 U14041 ( .A1(n13519), .A2(n11584), .B1(n11583), .B2(n13521), .ZN(
        n11585) );
  AOI211_X1 U14042 ( .C1(n11735), .C2(n13529), .A(n11586), .B(n11585), .ZN(
        n11587) );
  OAI211_X1 U14043 ( .C1(n11589), .C2(n13467), .A(n11588), .B(n11587), .ZN(
        P2_U3253) );
  INV_X1 U14044 ( .A(n11590), .ZN(n11591) );
  OAI222_X1 U14045 ( .A1(n11593), .A2(P3_U3151), .B1(n11761), .B2(n11592), 
        .C1(n13021), .C2(n11591), .ZN(P3_U3270) );
  INV_X1 U14046 ( .A(n11594), .ZN(n12418) );
  OAI222_X1 U14047 ( .A1(n14216), .A2(n11595), .B1(n14225), .B2(n12418), .C1(
        n12248), .C2(P1_U3086), .ZN(P1_U3334) );
  XNOR2_X1 U14048 ( .A(n11597), .B(n11596), .ZN(n13528) );
  OAI21_X1 U14049 ( .B1(n11606), .B2(n11598), .A(n11269), .ZN(n11600) );
  NOR2_X1 U14050 ( .A1(n11600), .A2(n11599), .ZN(n13530) );
  INV_X1 U14051 ( .A(n11601), .ZN(n11602) );
  AOI21_X1 U14052 ( .B1(n11604), .B2(n11603), .A(n11602), .ZN(n11605) );
  AOI22_X1 U14053 ( .A1(n13172), .A2(n13199), .B1(n13173), .B2(n13197), .ZN(
        n12427) );
  OAI21_X1 U14054 ( .B1(n11605), .B2(n13504), .A(n12427), .ZN(n13520) );
  AOI211_X1 U14055 ( .C1(n13528), .C2(n14982), .A(n13530), .B(n13520), .ZN(
        n11610) );
  OAI22_X1 U14056 ( .A1(n11606), .A2(n13677), .B1(n14995), .B2(n9250), .ZN(
        n11607) );
  INV_X1 U14057 ( .A(n11607), .ZN(n11608) );
  OAI21_X1 U14058 ( .B1(n11610), .B2(n14994), .A(n11608), .ZN(P2_U3463) );
  AOI22_X1 U14059 ( .A1(n13526), .A2(n13634), .B1(n6478), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n11609) );
  OAI21_X1 U14060 ( .B1(n11610), .B2(n6478), .A(n11609), .ZN(P2_U3510) );
  AOI21_X1 U14061 ( .B1(n11611), .B2(n11615), .A(n15249), .ZN(n11614) );
  OAI22_X1 U14062 ( .A1(n11727), .A2(n15243), .B1(n12363), .B2(n15241), .ZN(
        n11612) );
  AOI21_X1 U14063 ( .B1(n11614), .B2(n11613), .A(n11612), .ZN(n14464) );
  XNOR2_X1 U14064 ( .A(n11616), .B(n11615), .ZN(n14467) );
  NAND2_X1 U14065 ( .A1(n15266), .A2(n11617), .ZN(n15209) );
  INV_X1 U14066 ( .A(n12863), .ZN(n12818) );
  NOR2_X1 U14067 ( .A1(n15273), .A2(n11618), .ZN(n11621) );
  NAND2_X1 U14068 ( .A1(n11731), .A2(n12888), .ZN(n14463) );
  OAI22_X1 U14069 ( .A1(n11619), .A2(n14463), .B1(n11728), .B2(n15268), .ZN(
        n11620) );
  AOI211_X1 U14070 ( .C1(n14467), .C2(n12818), .A(n11621), .B(n11620), .ZN(
        n11622) );
  OAI21_X1 U14071 ( .B1(n14464), .B2(n12719), .A(n11622), .ZN(P3_U3221) );
  XNOR2_X1 U14072 ( .A(n11623), .B(n11625), .ZN(n14361) );
  INV_X1 U14073 ( .A(n14361), .ZN(n11638) );
  INV_X1 U14074 ( .A(n11624), .ZN(n11626) );
  AOI21_X1 U14075 ( .B1(n11626), .B2(n11625), .A(n14691), .ZN(n11630) );
  NAND2_X1 U14076 ( .A1(n14114), .A2(n14498), .ZN(n11628) );
  NAND2_X1 U14077 ( .A1(n13852), .A2(n14596), .ZN(n11627) );
  NAND2_X1 U14078 ( .A1(n11628), .A2(n11627), .ZN(n11757) );
  AOI21_X1 U14079 ( .B1(n11630), .B2(n11629), .A(n11757), .ZN(n14358) );
  INV_X1 U14080 ( .A(n14358), .ZN(n11636) );
  NAND2_X1 U14081 ( .A1(n14524), .A2(n12147), .ZN(n11631) );
  NAND3_X1 U14082 ( .A1(n11653), .A2(n14726), .A3(n11631), .ZN(n14357) );
  OAI22_X1 U14083 ( .A1(n14721), .A2(n11632), .B1(n11754), .B2(n14719), .ZN(
        n11633) );
  AOI21_X1 U14084 ( .B1(n12147), .B2(n14723), .A(n11633), .ZN(n11634) );
  OAI21_X1 U14085 ( .B1(n14357), .B2(n14088), .A(n11634), .ZN(n11635) );
  AOI21_X1 U14086 ( .B1(n11636), .B2(n14721), .A(n11635), .ZN(n11637) );
  OAI21_X1 U14087 ( .B1(n14107), .B2(n11638), .A(n11637), .ZN(P1_U3281) );
  INV_X1 U14088 ( .A(n11639), .ZN(n11640) );
  XNOR2_X1 U14089 ( .A(n12386), .B(n11641), .ZN(n11722) );
  XNOR2_X1 U14090 ( .A(n11723), .B(n12558), .ZN(n11645) );
  AOI22_X1 U14091 ( .A1(n12548), .A2(n11641), .B1(n12545), .B2(n12557), .ZN(
        n11643) );
  AND2_X1 U14092 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n15115) );
  AOI21_X1 U14093 ( .B1(n12522), .B2(n12559), .A(n15115), .ZN(n11642) );
  OAI211_X1 U14094 ( .C1(n14379), .C2(n14456), .A(n11643), .B(n11642), .ZN(
        n11644) );
  AOI21_X1 U14095 ( .B1(n11645), .B2(n14376), .A(n11644), .ZN(n11646) );
  INV_X1 U14096 ( .A(n11646), .ZN(P3_U3176) );
  XNOR2_X1 U14097 ( .A(n11647), .B(n11648), .ZN(n14550) );
  INV_X1 U14098 ( .A(n14550), .ZN(n11660) );
  OAI211_X1 U14099 ( .C1(n11650), .C2(n12286), .A(n11649), .B(n14716), .ZN(
        n11652) );
  AOI22_X1 U14100 ( .A1(n11945), .A2(n14498), .B1(n14596), .B2(n13851), .ZN(
        n11651) );
  NAND2_X1 U14101 ( .A1(n11652), .A2(n11651), .ZN(n14555) );
  AOI21_X1 U14102 ( .B1(n12151), .B2(n11653), .A(n14792), .ZN(n11654) );
  NAND2_X1 U14103 ( .A1(n11654), .A2(n14125), .ZN(n14551) );
  OAI22_X1 U14104 ( .A1(n14721), .A2(n11655), .B1(n11775), .B2(n14719), .ZN(
        n11656) );
  AOI21_X1 U14105 ( .B1(n12151), .B2(n14723), .A(n11656), .ZN(n11657) );
  OAI21_X1 U14106 ( .B1(n14551), .B2(n14088), .A(n11657), .ZN(n11658) );
  AOI21_X1 U14107 ( .B1(n14555), .B2(n14721), .A(n11658), .ZN(n11659) );
  OAI21_X1 U14108 ( .B1(n14107), .B2(n11660), .A(n11659), .ZN(P1_U3280) );
  INV_X1 U14109 ( .A(n11663), .ZN(n11662) );
  XNOR2_X1 U14110 ( .A(n11661), .B(n11662), .ZN(n13633) );
  INV_X1 U14111 ( .A(n13633), .ZN(n11674) );
  XNOR2_X1 U14112 ( .A(n11664), .B(n11663), .ZN(n11665) );
  AOI22_X1 U14113 ( .A1(n13172), .A2(n13197), .B1(n13173), .B2(n13196), .ZN(
        n14821) );
  OAI21_X1 U14114 ( .B1(n11665), .B2(n13504), .A(n14821), .ZN(n13631) );
  NAND2_X1 U14115 ( .A1(n13631), .A2(n13519), .ZN(n11673) );
  INV_X1 U14116 ( .A(n13509), .ZN(n11666) );
  AOI211_X1 U14117 ( .C1(n14830), .C2(n11667), .A(n13490), .B(n11666), .ZN(
        n13632) );
  INV_X1 U14118 ( .A(n14830), .ZN(n11668) );
  NOR2_X1 U14119 ( .A1(n11668), .A2(n13461), .ZN(n11671) );
  OAI22_X1 U14120 ( .A1(n13519), .A2(n11669), .B1(n14833), .B2(n13521), .ZN(
        n11670) );
  AOI211_X1 U14121 ( .C1(n13632), .C2(n13529), .A(n11671), .B(n11670), .ZN(
        n11672) );
  OAI211_X1 U14122 ( .C1(n11674), .C2(n13467), .A(n11673), .B(n11672), .ZN(
        P2_U3252) );
  OAI22_X1 U14123 ( .A1(n14558), .A2(n10660), .B1(n11676), .B2(n12331), .ZN(
        n11675) );
  XNOR2_X1 U14124 ( .A(n11675), .B(n12332), .ZN(n11749) );
  INV_X1 U14125 ( .A(n11944), .ZN(n12330) );
  OAI22_X1 U14126 ( .A1(n14558), .A2(n12334), .B1(n11676), .B2(n12330), .ZN(
        n11748) );
  XNOR2_X1 U14127 ( .A(n11749), .B(n11748), .ZN(n11686) );
  OR2_X1 U14128 ( .A1(n11678), .A2(n11677), .ZN(n11679) );
  INV_X1 U14129 ( .A(n14478), .ZN(n11682) );
  OAI22_X1 U14130 ( .A1(n11682), .A2(n12334), .B1(n11681), .B2(n12330), .ZN(
        n14483) );
  AOI22_X1 U14131 ( .A1(n14478), .A2(n12035), .B1(n10693), .B2(n13853), .ZN(
        n11683) );
  XOR2_X1 U14132 ( .A(n12332), .B(n11683), .Z(n14484) );
  INV_X1 U14133 ( .A(n14483), .ZN(n11684) );
  AOI21_X1 U14134 ( .B1(n11686), .B2(n11685), .A(n6564), .ZN(n11693) );
  NAND2_X1 U14135 ( .A1(n13851), .A2(n14498), .ZN(n11688) );
  NAND2_X1 U14136 ( .A1(n13853), .A2(n14596), .ZN(n11687) );
  NAND2_X1 U14137 ( .A1(n11688), .A2(n11687), .ZN(n14516) );
  NAND2_X1 U14138 ( .A1(n14601), .A2(n14516), .ZN(n11689) );
  OAI211_X1 U14139 ( .C1(n14606), .C2(n14519), .A(n11690), .B(n11689), .ZN(
        n11691) );
  AOI21_X1 U14140 ( .B1(n14521), .B2(n13794), .A(n11691), .ZN(n11692) );
  OAI21_X1 U14141 ( .B1(n11693), .B2(n14593), .A(n11692), .ZN(P1_U3236) );
  INV_X1 U14142 ( .A(n11694), .ZN(n11695) );
  OAI222_X1 U14143 ( .A1(n11697), .A2(P3_U3151), .B1(n11761), .B2(n11696), 
        .C1(n13021), .C2(n11695), .ZN(P3_U3269) );
  XNOR2_X1 U14144 ( .A(n13672), .B(n6469), .ZN(n11708) );
  INV_X1 U14145 ( .A(n11708), .ZN(n11700) );
  NAND2_X1 U14146 ( .A1(n11701), .A2(n11703), .ZN(n11707) );
  NAND3_X1 U14147 ( .A1(n14823), .A2(n11700), .A3(n11707), .ZN(n11711) );
  INV_X1 U14148 ( .A(n11703), .ZN(n11706) );
  INV_X1 U14149 ( .A(n11702), .ZN(n11705) );
  AOI21_X1 U14150 ( .B1(n11703), .B2(n11702), .A(n11701), .ZN(n11704) );
  AOI211_X1 U14151 ( .C1(n11706), .C2(n11705), .A(n11708), .B(n11704), .ZN(
        n11709) );
  AND2_X1 U14152 ( .A1(n11708), .A2(n11707), .ZN(n11802) );
  INV_X1 U14153 ( .A(n11807), .ZN(n11721) );
  AOI22_X1 U14154 ( .A1(n6716), .A2(n13148), .B1(n13167), .B2(n13195), .ZN(
        n11720) );
  NAND2_X1 U14155 ( .A1(n13173), .A2(n13194), .ZN(n11716) );
  NAND2_X1 U14156 ( .A1(n13172), .A2(n13196), .ZN(n11715) );
  NAND2_X1 U14157 ( .A1(n11716), .A2(n11715), .ZN(n13491) );
  AOI22_X1 U14158 ( .A1(n13159), .A2(n13491), .B1(P2_U3088), .B2(
        P2_REG3_REG_15__SCAN_IN), .ZN(n11717) );
  OAI21_X1 U14159 ( .B1(n13494), .B2(n14832), .A(n11717), .ZN(n11718) );
  AOI21_X1 U14160 ( .B1(n13672), .B2(n14829), .A(n11718), .ZN(n11719) );
  OAI21_X1 U14161 ( .B1(n11721), .B2(n11720), .A(n11719), .ZN(P2_U3213) );
  OAI22_X1 U14162 ( .A1(n11723), .A2(n11727), .B1(n7489), .B2(n11722), .ZN(
        n11816) );
  XNOR2_X1 U14163 ( .A(n11724), .B(n12386), .ZN(n11817) );
  XNOR2_X1 U14164 ( .A(n11817), .B(n14454), .ZN(n11725) );
  XNOR2_X1 U14165 ( .A(n11816), .B(n11725), .ZN(n11733) );
  AOI22_X1 U14166 ( .A1(n12545), .A2(n12556), .B1(P3_REG3_REG_12__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11726) );
  OAI21_X1 U14167 ( .B1(n11727), .B2(n12543), .A(n11726), .ZN(n11730) );
  NOR2_X1 U14168 ( .A1(n14379), .A2(n11728), .ZN(n11729) );
  AOI211_X1 U14169 ( .C1(n11731), .C2(n12548), .A(n11730), .B(n11729), .ZN(
        n11732) );
  OAI21_X1 U14170 ( .B1(n11733), .B2(n12550), .A(n11732), .ZN(P3_U3164) );
  AOI211_X1 U14171 ( .C1(n14982), .C2(n11736), .A(n11735), .B(n11734), .ZN(
        n11743) );
  INV_X1 U14172 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n11737) );
  OAI22_X1 U14173 ( .A1(n11738), .A2(n13677), .B1(n14995), .B2(n11737), .ZN(
        n11739) );
  INV_X1 U14174 ( .A(n11739), .ZN(n11740) );
  OAI21_X1 U14175 ( .B1(n11743), .B2(n14994), .A(n11740), .ZN(P2_U3466) );
  AOI22_X1 U14176 ( .A1(n11741), .A2(n13634), .B1(n6478), .B2(
        P2_REG1_REG_12__SCAN_IN), .ZN(n11742) );
  OAI21_X1 U14177 ( .B1(n11743), .B2(n6478), .A(n11742), .ZN(P2_U3511) );
  INV_X1 U14178 ( .A(n12147), .ZN(n14359) );
  NAND2_X1 U14179 ( .A1(n12147), .A2(n12035), .ZN(n11745) );
  NAND2_X1 U14180 ( .A1(n13851), .A2(n10693), .ZN(n11744) );
  NAND2_X1 U14181 ( .A1(n11745), .A2(n11744), .ZN(n11746) );
  XNOR2_X1 U14182 ( .A(n11746), .B(n12025), .ZN(n11764) );
  AND2_X1 U14183 ( .A1(n12039), .A2(n13851), .ZN(n11747) );
  AOI21_X1 U14184 ( .B1(n12147), .B2(n10693), .A(n11747), .ZN(n11765) );
  XNOR2_X1 U14185 ( .A(n11764), .B(n11765), .ZN(n11750) );
  NOR2_X1 U14186 ( .A1(n11749), .A2(n11748), .ZN(n11751) );
  INV_X1 U14187 ( .A(n11768), .ZN(n11753) );
  OAI21_X1 U14188 ( .B1(n6564), .B2(n11751), .A(n11750), .ZN(n11752) );
  NAND3_X1 U14189 ( .A1(n11753), .A2(n14488), .A3(n11752), .ZN(n11759) );
  NOR2_X1 U14190 ( .A1(n14606), .A2(n11754), .ZN(n11755) );
  AOI211_X1 U14191 ( .C1(n14601), .C2(n11757), .A(n11756), .B(n11755), .ZN(
        n11758) );
  OAI211_X1 U14192 ( .C1(n14359), .C2(n13817), .A(n11759), .B(n11758), .ZN(
        P1_U3224) );
  INV_X1 U14193 ( .A(n11760), .ZN(n11763) );
  OAI222_X1 U14194 ( .A1(n12670), .A2(P3_U3151), .B1(n13021), .B2(n11763), 
        .C1(n11762), .C2(n11761), .ZN(P3_U3268) );
  INV_X1 U14195 ( .A(n11764), .ZN(n11767) );
  INV_X1 U14196 ( .A(n11765), .ZN(n11766) );
  AND2_X1 U14197 ( .A1(n12039), .A2(n14114), .ZN(n11769) );
  AOI21_X1 U14198 ( .B1(n12151), .B2(n10693), .A(n11769), .ZN(n11940) );
  INV_X1 U14199 ( .A(n12151), .ZN(n14552) );
  INV_X1 U14200 ( .A(n10664), .ZN(n12334) );
  OAI22_X1 U14201 ( .A1(n14552), .A2(n10660), .B1(n12152), .B2(n12334), .ZN(
        n11770) );
  XNOR2_X1 U14202 ( .A(n11770), .B(n12332), .ZN(n11938) );
  XOR2_X1 U14203 ( .A(n11940), .B(n11938), .Z(n11941) );
  XNOR2_X1 U14204 ( .A(n11942), .B(n11941), .ZN(n11778) );
  OAI21_X1 U14205 ( .B1(n13811), .B2(n11772), .A(n11771), .ZN(n11773) );
  AOI21_X1 U14206 ( .B1(n13814), .B2(n13851), .A(n11773), .ZN(n11774) );
  OAI21_X1 U14207 ( .B1(n14606), .B2(n11775), .A(n11774), .ZN(n11776) );
  AOI21_X1 U14208 ( .B1(n12151), .B2(n13794), .A(n11776), .ZN(n11777) );
  OAI21_X1 U14209 ( .B1(n11778), .B2(n14593), .A(n11777), .ZN(P1_U3234) );
  INV_X1 U14210 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n11779) );
  NAND2_X1 U14211 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13761)
         );
  OAI21_X1 U14212 ( .B1(n14653), .B2(n11779), .A(n13761), .ZN(n11789) );
  NAND2_X1 U14213 ( .A1(n11793), .A2(n11782), .ZN(n11783) );
  NAND2_X1 U14214 ( .A1(n14644), .A2(n7875), .ZN(n14643) );
  NAND2_X1 U14215 ( .A1(n11783), .A2(n14643), .ZN(n11787) );
  NOR2_X1 U14216 ( .A1(n11885), .A2(n11784), .ZN(n11785) );
  AOI21_X1 U14217 ( .B1(n11885), .B2(n11784), .A(n11785), .ZN(n11786) );
  NOR2_X1 U14218 ( .A1(n11787), .A2(n11786), .ZN(n11884) );
  AOI211_X1 U14219 ( .C1(n11787), .C2(n11786), .A(n13911), .B(n11884), .ZN(
        n11788) );
  AOI211_X1 U14220 ( .C1(n14645), .C2(n11885), .A(n11789), .B(n11788), .ZN(
        n11801) );
  OAI21_X1 U14221 ( .B1(n14119), .B2(n11791), .A(n11790), .ZN(n11792) );
  NOR2_X1 U14222 ( .A1(n14646), .A2(n11792), .ZN(n11794) );
  XOR2_X1 U14223 ( .A(n11793), .B(n11792), .Z(n14641) );
  NOR2_X1 U14224 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14641), .ZN(n14640) );
  NOR2_X1 U14225 ( .A1(n11794), .A2(n14640), .ZN(n11799) );
  MUX2_X1 U14226 ( .A(P1_REG2_REG_16__SCAN_IN), .B(n11795), .S(n11885), .Z(
        n11798) );
  NAND2_X1 U14227 ( .A1(n11796), .A2(n11795), .ZN(n11797) );
  NAND2_X1 U14228 ( .A1(n11885), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11891) );
  NAND3_X1 U14229 ( .A1(n11799), .A2(n11797), .A3(n11891), .ZN(n11892) );
  OAI211_X1 U14230 ( .C1(n11799), .C2(n11798), .A(n11892), .B(n14649), .ZN(
        n11800) );
  NAND2_X1 U14231 ( .A1(n11801), .A2(n11800), .ZN(P1_U3259) );
  NAND2_X1 U14232 ( .A1(n13194), .A2(n13490), .ZN(n12068) );
  XNOR2_X1 U14233 ( .A(n13477), .B(n6469), .ZN(n12074) );
  XOR2_X1 U14234 ( .A(n12068), .B(n12074), .Z(n11809) );
  INV_X1 U14235 ( .A(n11802), .ZN(n11803) );
  NOR2_X1 U14236 ( .A1(n11804), .A2(n11803), .ZN(n11805) );
  INV_X1 U14237 ( .A(n11805), .ZN(n11806) );
  AOI21_X1 U14238 ( .B1(n11809), .B2(n11808), .A(n12077), .ZN(n11815) );
  NOR2_X1 U14239 ( .A1(n14832), .A2(n13471), .ZN(n11813) );
  NAND2_X1 U14240 ( .A1(n13172), .A2(n13195), .ZN(n11811) );
  NAND2_X1 U14241 ( .A1(n13173), .A2(n13193), .ZN(n11810) );
  AND2_X1 U14242 ( .A1(n11811), .A2(n11810), .ZN(n13611) );
  OAI22_X1 U14243 ( .A1(n14822), .A2(n13611), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14931), .ZN(n11812) );
  AOI211_X1 U14244 ( .C1(n13477), .C2(n14829), .A(n11813), .B(n11812), .ZN(
        n11814) );
  OAI21_X1 U14245 ( .B1(n11815), .B2(n14824), .A(n11814), .ZN(P2_U3198) );
  INV_X1 U14246 ( .A(n11816), .ZN(n11820) );
  NAND2_X1 U14247 ( .A1(n11817), .A2(n12557), .ZN(n11819) );
  INV_X1 U14248 ( .A(n11817), .ZN(n11818) );
  XNOR2_X1 U14249 ( .A(n11833), .B(n12386), .ZN(n12362) );
  XNOR2_X1 U14250 ( .A(n12362), .B(n12363), .ZN(n11821) );
  XNOR2_X1 U14251 ( .A(n12361), .B(n11821), .ZN(n11827) );
  NOR2_X1 U14252 ( .A1(n14373), .A2(n11833), .ZN(n11824) );
  AOI22_X1 U14253 ( .A1(n12545), .A2(n12856), .B1(P3_REG3_REG_13__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11822) );
  OAI21_X1 U14254 ( .B1(n14454), .B2(n12543), .A(n11822), .ZN(n11823) );
  AOI211_X1 U14255 ( .C1(n11825), .C2(n12535), .A(n11824), .B(n11823), .ZN(
        n11826) );
  OAI21_X1 U14256 ( .B1(n11827), .B2(n12550), .A(n11826), .ZN(P3_U3174) );
  XNOR2_X1 U14257 ( .A(n11829), .B(n11828), .ZN(n14462) );
  INV_X1 U14258 ( .A(n14462), .ZN(n11839) );
  XNOR2_X1 U14259 ( .A(n11831), .B(n11830), .ZN(n11832) );
  OAI222_X1 U14260 ( .A1(n15243), .A2(n14454), .B1(n15241), .B2(n12542), .C1(
        n11832), .C2(n15249), .ZN(n14460) );
  NAND2_X1 U14261 ( .A1(n14460), .A2(n15273), .ZN(n11838) );
  NOR2_X1 U14262 ( .A1(n11833), .A2(n15253), .ZN(n14461) );
  OAI22_X1 U14263 ( .A1(n15273), .A2(n11835), .B1(n11834), .B2(n15268), .ZN(
        n11836) );
  AOI21_X1 U14264 ( .B1(n15227), .B2(n14461), .A(n11836), .ZN(n11837) );
  OAI211_X1 U14265 ( .C1(n12863), .C2(n11839), .A(n11838), .B(n11837), .ZN(
        P3_U3220) );
  INV_X1 U14266 ( .A(n11840), .ZN(n11841) );
  AOI21_X1 U14267 ( .B1(n11848), .B2(n11842), .A(n11841), .ZN(n14538) );
  INV_X1 U14268 ( .A(n14505), .ZN(n11844) );
  AOI211_X1 U14269 ( .C1(n11950), .C2(n14124), .A(n14792), .B(n11844), .ZN(
        n14540) );
  INV_X1 U14270 ( .A(n11950), .ZN(n13832) );
  AOI22_X1 U14271 ( .A1(n14701), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n13833), 
        .B2(n14702), .ZN(n11845) );
  OAI21_X1 U14272 ( .B1(n13832), .B2(n14103), .A(n11845), .ZN(n11846) );
  AOI21_X1 U14273 ( .B1(n14540), .B2(n14731), .A(n11846), .ZN(n11852) );
  OAI211_X1 U14274 ( .C1(n11849), .C2(n11848), .A(n11847), .B(n14716), .ZN(
        n11850) );
  AOI22_X1 U14275 ( .A1(n11945), .A2(n14596), .B1(n14498), .B2(n13850), .ZN(
        n13837) );
  NAND2_X1 U14276 ( .A1(n11850), .A2(n13837), .ZN(n14539) );
  NAND2_X1 U14277 ( .A1(n14539), .A2(n14721), .ZN(n11851) );
  OAI211_X1 U14278 ( .C1(n14538), .C2(n14107), .A(n11852), .B(n11851), .ZN(
        P1_U3278) );
  NAND2_X1 U14279 ( .A1(n11855), .A2(n14210), .ZN(n11853) );
  OAI211_X1 U14280 ( .C1(n11854), .C2(n14216), .A(n11853), .B(n12324), .ZN(
        P1_U3332) );
  NAND2_X1 U14281 ( .A1(n11855), .A2(n13694), .ZN(n11857) );
  OAI211_X1 U14282 ( .C1(n11858), .C2(n13705), .A(n11857), .B(n11856), .ZN(
        P2_U3304) );
  INV_X1 U14283 ( .A(n11859), .ZN(n11863) );
  OAI222_X1 U14284 ( .A1(n14216), .A2(n11861), .B1(n14225), .B2(n11863), .C1(
        n11860), .C2(P1_U3086), .ZN(P1_U3331) );
  OAI222_X1 U14285 ( .A1(n11864), .A2(P2_U3088), .B1(n13708), .B2(n11863), 
        .C1(n11862), .C2(n13705), .ZN(P2_U3303) );
  INV_X1 U14286 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12608) );
  XNOR2_X1 U14287 ( .A(n11865), .B(n11868), .ZN(n11866) );
  OAI22_X1 U14288 ( .A1(n12476), .A2(n15241), .B1(n12363), .B2(n15243), .ZN(
        n14371) );
  AOI21_X1 U14289 ( .B1(n11866), .B2(n15262), .A(n14371), .ZN(n11875) );
  MUX2_X1 U14290 ( .A(n12608), .B(n11875), .S(n15331), .Z(n11870) );
  OAI21_X1 U14291 ( .B1(n6656), .B2(n11868), .A(n11867), .ZN(n11874) );
  INV_X1 U14292 ( .A(n12903), .ZN(n12919) );
  NAND2_X1 U14293 ( .A1(n11874), .A2(n12919), .ZN(n11869) );
  OAI211_X1 U14294 ( .C1(n12907), .C2(n14374), .A(n11870), .B(n11869), .ZN(
        P3_U3473) );
  MUX2_X1 U14295 ( .A(n11871), .B(n11875), .S(n15318), .Z(n11873) );
  INV_X1 U14296 ( .A(n12975), .ZN(n13006) );
  NAND2_X1 U14297 ( .A1(n11874), .A2(n13006), .ZN(n11872) );
  OAI211_X1 U14298 ( .C1(n12983), .C2(n14374), .A(n11873), .B(n11872), .ZN(
        P3_U3432) );
  INV_X1 U14299 ( .A(n11874), .ZN(n11880) );
  MUX2_X1 U14300 ( .A(n8438), .B(n11875), .S(n15273), .Z(n11879) );
  INV_X1 U14301 ( .A(n14374), .ZN(n11877) );
  AOI22_X1 U14302 ( .A1(n11877), .A2(n12860), .B1(n15226), .B2(n11876), .ZN(
        n11878) );
  OAI211_X1 U14303 ( .C1(n11880), .C2(n12863), .A(n11879), .B(n11878), .ZN(
        P3_U3219) );
  INV_X1 U14304 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n11883) );
  NOR2_X1 U14305 ( .A1(n11881), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13776) );
  INV_X1 U14306 ( .A(n13776), .ZN(n11882) );
  OAI21_X1 U14307 ( .B1(n14653), .B2(n11883), .A(n11882), .ZN(n11889) );
  AOI21_X1 U14308 ( .B1(n11885), .B2(P1_REG1_REG_16__SCAN_IN), .A(n11884), 
        .ZN(n11887) );
  XNOR2_X1 U14309 ( .A(n13890), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n11886) );
  AOI211_X1 U14310 ( .C1(n11887), .C2(n11886), .A(n13911), .B(n13889), .ZN(
        n11888) );
  AOI211_X1 U14311 ( .C1(n14645), .C2(n13890), .A(n11889), .B(n11888), .ZN(
        n11898) );
  INV_X1 U14312 ( .A(n11892), .ZN(n11896) );
  NAND2_X1 U14313 ( .A1(n13887), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n11890) );
  OAI211_X1 U14314 ( .C1(n13887), .C2(P1_REG2_REG_17__SCAN_IN), .A(n11890), 
        .B(n11891), .ZN(n11895) );
  NAND2_X1 U14315 ( .A1(n11892), .A2(n11891), .ZN(n11894) );
  NAND2_X1 U14316 ( .A1(n13890), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n11893) );
  OAI211_X1 U14317 ( .C1(n13890), .C2(P1_REG2_REG_17__SCAN_IN), .A(n11894), 
        .B(n11893), .ZN(n13886) );
  OAI211_X1 U14318 ( .C1(n11896), .C2(n11895), .A(n13886), .B(n14649), .ZN(
        n11897) );
  NAND2_X1 U14319 ( .A1(n11898), .A2(n11897), .ZN(P1_U3260) );
  MUX2_X1 U14320 ( .A(n11899), .B(P1_REG2_REG_1__SCAN_IN), .S(n14736), .Z(
        n11908) );
  NAND2_X1 U14321 ( .A1(n13974), .A2(n11900), .ZN(n11905) );
  INV_X1 U14322 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n11901) );
  OAI22_X1 U14323 ( .A1(n14103), .A2(n11902), .B1(n11901), .B2(n14719), .ZN(
        n11903) );
  INV_X1 U14324 ( .A(n11903), .ZN(n11904) );
  OAI211_X1 U14325 ( .C1(n11906), .C2(n14094), .A(n11905), .B(n11904), .ZN(
        n11907) );
  OR2_X1 U14326 ( .A1(n11908), .A2(n11907), .ZN(P1_U3292) );
  INV_X1 U14327 ( .A(n11909), .ZN(n13707) );
  OAI222_X1 U14328 ( .A1(n14216), .A2(n11910), .B1(n14225), .B2(n13707), .C1(
        n11911), .C2(P1_U3086), .ZN(P1_U3330) );
  INV_X1 U14329 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n11913) );
  AOI22_X1 U14330 ( .A1(n6674), .A2(n11913), .B1(n11912), .B2(n11911), .ZN(
        P1_U3446) );
  NOR2_X1 U14331 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11914), .ZN(n11919) );
  AOI211_X1 U14332 ( .C1(n11917), .C2(n11916), .A(n14932), .B(n11915), .ZN(
        n11918) );
  AOI211_X1 U14333 ( .C1(n14924), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n11919), .B(
        n11918), .ZN(n11926) );
  INV_X1 U14334 ( .A(n11920), .ZN(n11924) );
  NAND3_X1 U14335 ( .A1(n14884), .A2(n11922), .A3(n11921), .ZN(n11923) );
  NAND3_X1 U14336 ( .A1(n14941), .A2(n11924), .A3(n11923), .ZN(n11925) );
  OAI211_X1 U14337 ( .C1(n14930), .C2(n11927), .A(n11926), .B(n11925), .ZN(
        P2_U3221) );
  INV_X1 U14338 ( .A(n11928), .ZN(n13692) );
  OAI222_X1 U14339 ( .A1(n14225), .A2(n13692), .B1(n11930), .B2(P1_U3086), 
        .C1(n11929), .C2(n14216), .ZN(P1_U3326) );
  INV_X1 U14340 ( .A(n14137), .ZN(n13938) );
  NAND2_X1 U14341 ( .A1(n14137), .A2(n12035), .ZN(n11932) );
  NAND2_X1 U14342 ( .A1(n13844), .A2(n12028), .ZN(n11931) );
  NAND2_X1 U14343 ( .A1(n11932), .A2(n11931), .ZN(n11933) );
  XNOR2_X1 U14344 ( .A(n11933), .B(n12332), .ZN(n11937) );
  NAND2_X1 U14345 ( .A1(n14137), .A2(n12028), .ZN(n11935) );
  NAND2_X1 U14346 ( .A1(n13844), .A2(n11944), .ZN(n11934) );
  NAND2_X1 U14347 ( .A1(n11935), .A2(n11934), .ZN(n11936) );
  NOR2_X1 U14348 ( .A1(n11937), .A2(n11936), .ZN(n12329) );
  AOI21_X1 U14349 ( .B1(n11937), .B2(n11936), .A(n12329), .ZN(n12046) );
  INV_X1 U14350 ( .A(n11938), .ZN(n11939) );
  AOI22_X1 U14351 ( .A1(n14545), .A2(n12035), .B1(n12028), .B2(n11945), .ZN(
        n11943) );
  XNOR2_X1 U14352 ( .A(n11943), .B(n12332), .ZN(n11947) );
  AOI22_X1 U14353 ( .A1(n14545), .A2(n10693), .B1(n12039), .B2(n11945), .ZN(
        n11946) );
  NAND2_X1 U14354 ( .A1(n11947), .A2(n11946), .ZN(n11948) );
  OAI21_X1 U14355 ( .B1(n11947), .B2(n11946), .A(n11948), .ZN(n13715) );
  INV_X1 U14356 ( .A(n11948), .ZN(n11949) );
  AOI22_X1 U14357 ( .A1(n11950), .A2(n12035), .B1(n10693), .B2(n14499), .ZN(
        n11951) );
  XOR2_X1 U14358 ( .A(n12332), .B(n11951), .Z(n11952) );
  OAI22_X1 U14359 ( .A1(n13832), .A2(n12334), .B1(n14113), .B2(n12330), .ZN(
        n13831) );
  NAND2_X1 U14360 ( .A1(n14531), .A2(n12035), .ZN(n11956) );
  NAND2_X1 U14361 ( .A1(n13850), .A2(n10693), .ZN(n11955) );
  NAND2_X1 U14362 ( .A1(n11956), .A2(n11955), .ZN(n11957) );
  XNOR2_X1 U14363 ( .A(n11957), .B(n12025), .ZN(n11960) );
  AND2_X1 U14364 ( .A1(n12039), .A2(n13850), .ZN(n11958) );
  AOI21_X1 U14365 ( .B1(n14531), .B2(n10693), .A(n11958), .ZN(n11959) );
  NAND2_X1 U14366 ( .A1(n11960), .A2(n11959), .ZN(n11961) );
  OAI21_X1 U14367 ( .B1(n11960), .B2(n11959), .A(n11961), .ZN(n13759) );
  INV_X1 U14368 ( .A(n11961), .ZN(n13770) );
  INV_X1 U14369 ( .A(n14497), .ZN(n12167) );
  OAI22_X1 U14370 ( .A1(n14104), .A2(n10660), .B1(n12167), .B2(n12334), .ZN(
        n11962) );
  XNOR2_X1 U14371 ( .A(n11962), .B(n12025), .ZN(n11965) );
  OR2_X1 U14372 ( .A1(n14104), .A2(n12334), .ZN(n11964) );
  NAND2_X1 U14373 ( .A1(n14497), .A2(n12039), .ZN(n11963) );
  AND2_X1 U14374 ( .A1(n11964), .A2(n11963), .ZN(n11966) );
  NAND2_X1 U14375 ( .A1(n11965), .A2(n11966), .ZN(n11970) );
  INV_X1 U14376 ( .A(n11965), .ZN(n11968) );
  INV_X1 U14377 ( .A(n11966), .ZN(n11967) );
  NAND2_X1 U14378 ( .A1(n11968), .A2(n11967), .ZN(n11969) );
  AND2_X1 U14379 ( .A1(n11970), .A2(n11969), .ZN(n13769) );
  OR2_X1 U14380 ( .A1(n14188), .A2(n12334), .ZN(n11972) );
  NAND2_X1 U14381 ( .A1(n14066), .A2(n12039), .ZN(n11971) );
  NAND2_X1 U14382 ( .A1(n11972), .A2(n11971), .ZN(n11977) );
  INV_X1 U14383 ( .A(n14066), .ZN(n12187) );
  OAI22_X1 U14384 ( .A1(n14188), .A2(n10660), .B1(n12187), .B2(n12334), .ZN(
        n11973) );
  XNOR2_X1 U14385 ( .A(n11973), .B(n12332), .ZN(n11976) );
  XOR2_X1 U14386 ( .A(n11977), .B(n11976), .Z(n13807) );
  AND2_X1 U14387 ( .A1(n14081), .A2(n12039), .ZN(n11974) );
  AOI21_X1 U14388 ( .B1(n14181), .B2(n10693), .A(n11974), .ZN(n11981) );
  AOI22_X1 U14389 ( .A1(n14181), .A2(n12035), .B1(n6542), .B2(n14081), .ZN(
        n11975) );
  XNOR2_X1 U14390 ( .A(n11975), .B(n12332), .ZN(n11980) );
  XOR2_X1 U14391 ( .A(n11981), .B(n11980), .Z(n13733) );
  INV_X1 U14392 ( .A(n11976), .ZN(n11979) );
  INV_X1 U14393 ( .A(n11977), .ZN(n11978) );
  NAND2_X1 U14394 ( .A1(n11979), .A2(n11978), .ZN(n13731) );
  INV_X1 U14395 ( .A(n11981), .ZN(n11982) );
  OAI22_X1 U14396 ( .A1(n14177), .A2(n12334), .B1(n14034), .B2(n12330), .ZN(
        n11985) );
  OAI22_X1 U14397 ( .A1(n14177), .A2(n10660), .B1(n14034), .B2(n12334), .ZN(
        n11984) );
  XNOR2_X1 U14398 ( .A(n11984), .B(n12332), .ZN(n11986) );
  XOR2_X1 U14399 ( .A(n11985), .B(n11986), .Z(n13787) );
  NAND2_X1 U14400 ( .A1(n14044), .A2(n12035), .ZN(n11988) );
  NAND2_X1 U14401 ( .A1(n14050), .A2(n10693), .ZN(n11987) );
  NAND2_X1 U14402 ( .A1(n11988), .A2(n11987), .ZN(n11989) );
  XNOR2_X1 U14403 ( .A(n11989), .B(n12332), .ZN(n11993) );
  NAND2_X1 U14404 ( .A1(n14044), .A2(n12028), .ZN(n11991) );
  NAND2_X1 U14405 ( .A1(n14050), .A2(n12039), .ZN(n11990) );
  NAND2_X1 U14406 ( .A1(n11991), .A2(n11990), .ZN(n11992) );
  NOR2_X1 U14407 ( .A1(n11993), .A2(n11992), .ZN(n11994) );
  AOI21_X1 U14408 ( .B1(n11993), .B2(n11992), .A(n11994), .ZN(n13740) );
  INV_X1 U14409 ( .A(n11994), .ZN(n11995) );
  NAND2_X1 U14410 ( .A1(n13739), .A2(n11995), .ZN(n13798) );
  NAND2_X1 U14411 ( .A1(n14165), .A2(n12035), .ZN(n11997) );
  NAND2_X1 U14412 ( .A1(n14032), .A2(n6542), .ZN(n11996) );
  NAND2_X1 U14413 ( .A1(n11997), .A2(n11996), .ZN(n11998) );
  XNOR2_X1 U14414 ( .A(n11998), .B(n12332), .ZN(n12002) );
  NAND2_X1 U14415 ( .A1(n14165), .A2(n10693), .ZN(n12000) );
  NAND2_X1 U14416 ( .A1(n14032), .A2(n12039), .ZN(n11999) );
  NAND2_X1 U14417 ( .A1(n12000), .A2(n11999), .ZN(n12001) );
  NOR2_X1 U14418 ( .A1(n12002), .A2(n12001), .ZN(n12003) );
  AOI21_X1 U14419 ( .B1(n12002), .B2(n12001), .A(n12003), .ZN(n13799) );
  NAND2_X1 U14420 ( .A1(n13798), .A2(n13799), .ZN(n13797) );
  INV_X1 U14421 ( .A(n12003), .ZN(n12004) );
  NAND2_X1 U14422 ( .A1(n14160), .A2(n12035), .ZN(n12006) );
  NAND2_X1 U14423 ( .A1(n13848), .A2(n10693), .ZN(n12005) );
  NAND2_X1 U14424 ( .A1(n12006), .A2(n12005), .ZN(n12007) );
  XNOR2_X1 U14425 ( .A(n12007), .B(n12332), .ZN(n12011) );
  NAND2_X1 U14426 ( .A1(n14160), .A2(n10693), .ZN(n12009) );
  NAND2_X1 U14427 ( .A1(n13848), .A2(n12039), .ZN(n12008) );
  NAND2_X1 U14428 ( .A1(n12009), .A2(n12008), .ZN(n12010) );
  NOR2_X1 U14429 ( .A1(n12011), .A2(n12010), .ZN(n12012) );
  AOI21_X1 U14430 ( .B1(n12011), .B2(n12010), .A(n12012), .ZN(n13724) );
  INV_X1 U14431 ( .A(n12012), .ZN(n13780) );
  NAND2_X1 U14432 ( .A1(n14155), .A2(n12035), .ZN(n12014) );
  NAND2_X1 U14433 ( .A1(n13847), .A2(n10693), .ZN(n12013) );
  NAND2_X1 U14434 ( .A1(n12014), .A2(n12013), .ZN(n12015) );
  XNOR2_X1 U14435 ( .A(n12015), .B(n12025), .ZN(n12017) );
  AND2_X1 U14436 ( .A1(n11944), .A2(n13847), .ZN(n12016) );
  AOI21_X1 U14437 ( .B1(n14155), .B2(n6542), .A(n12016), .ZN(n12018) );
  NAND2_X1 U14438 ( .A1(n12017), .A2(n12018), .ZN(n12022) );
  INV_X1 U14439 ( .A(n12017), .ZN(n12020) );
  INV_X1 U14440 ( .A(n12018), .ZN(n12019) );
  NAND2_X1 U14441 ( .A1(n12020), .A2(n12019), .ZN(n12021) );
  NAND2_X1 U14442 ( .A1(n12022), .A2(n12021), .ZN(n13779) );
  INV_X1 U14443 ( .A(n12022), .ZN(n13750) );
  NAND2_X1 U14444 ( .A1(n14147), .A2(n12035), .ZN(n12024) );
  NAND2_X1 U14445 ( .A1(n13846), .A2(n10693), .ZN(n12023) );
  NAND2_X1 U14446 ( .A1(n12024), .A2(n12023), .ZN(n12026) );
  XNOR2_X1 U14447 ( .A(n12026), .B(n12025), .ZN(n12029) );
  AND2_X1 U14448 ( .A1(n11944), .A2(n13846), .ZN(n12027) );
  AOI21_X1 U14449 ( .B1(n14147), .B2(n6542), .A(n12027), .ZN(n12030) );
  NAND2_X1 U14450 ( .A1(n12029), .A2(n12030), .ZN(n12034) );
  INV_X1 U14451 ( .A(n12029), .ZN(n12032) );
  INV_X1 U14452 ( .A(n12030), .ZN(n12031) );
  NAND2_X1 U14453 ( .A1(n12032), .A2(n12031), .ZN(n12033) );
  NAND2_X1 U14454 ( .A1(n13960), .A2(n12035), .ZN(n12037) );
  NAND2_X1 U14455 ( .A1(n13845), .A2(n6542), .ZN(n12036) );
  NAND2_X1 U14456 ( .A1(n12037), .A2(n12036), .ZN(n12038) );
  XNOR2_X1 U14457 ( .A(n12038), .B(n12332), .ZN(n12043) );
  NAND2_X1 U14458 ( .A1(n13960), .A2(n12028), .ZN(n12041) );
  NAND2_X1 U14459 ( .A1(n13845), .A2(n11944), .ZN(n12040) );
  NAND2_X1 U14460 ( .A1(n12041), .A2(n12040), .ZN(n12042) );
  NOR2_X1 U14461 ( .A1(n12043), .A2(n12042), .ZN(n12044) );
  AOI21_X1 U14462 ( .B1(n12043), .B2(n12042), .A(n12044), .ZN(n13820) );
  INV_X1 U14463 ( .A(n12044), .ZN(n12045) );
  INV_X1 U14464 ( .A(n12048), .ZN(n13936) );
  AOI22_X1 U14465 ( .A1(n14596), .A2(n13845), .B1(n13843), .B2(n14597), .ZN(
        n13932) );
  OAI22_X1 U14466 ( .A1(n13932), .A2(n13836), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12049), .ZN(n12050) );
  AOI21_X1 U14467 ( .B1(n13834), .B2(n13936), .A(n12050), .ZN(n12051) );
  INV_X1 U14468 ( .A(n14721), .ZN(n14701) );
  OAI22_X1 U14469 ( .A1(n14721), .A2(n12052), .B1(n12342), .B2(n14719), .ZN(
        n12055) );
  NOR2_X1 U14470 ( .A1(n12053), .A2(n14088), .ZN(n12054) );
  AOI211_X1 U14471 ( .C1(n14723), .C2(n12344), .A(n12055), .B(n12054), .ZN(
        n12059) );
  NAND3_X1 U14472 ( .A1(n12057), .A2(n14527), .A3(n12056), .ZN(n12058) );
  OAI211_X1 U14473 ( .C1(n12060), .C2(n14701), .A(n12059), .B(n12058), .ZN(
        P1_U3265) );
  INV_X1 U14474 ( .A(n13695), .ZN(n12063) );
  OAI222_X1 U14475 ( .A1(n14225), .A2(n12063), .B1(n12062), .B2(P1_U3086), 
        .C1(n12061), .C2(n14216), .ZN(P1_U3327) );
  INV_X1 U14476 ( .A(n12064), .ZN(n12066) );
  OAI222_X1 U14477 ( .A1(n13705), .A2(n12067), .B1(n13708), .B2(n12066), .C1(
        P2_U3088), .C2(n12065), .ZN(P2_U3305) );
  INV_X1 U14478 ( .A(n12068), .ZN(n12069) );
  XNOR2_X1 U14479 ( .A(n12073), .B(n6469), .ZN(n13027) );
  NAND2_X1 U14480 ( .A1(n13193), .A2(n13490), .ZN(n13025) );
  XNOR2_X1 U14481 ( .A(n13027), .B(n13025), .ZN(n12075) );
  NOR2_X1 U14482 ( .A1(n14832), .A2(n13462), .ZN(n12072) );
  AOI22_X1 U14483 ( .A1(n13192), .A2(n13173), .B1(n13172), .B2(n13194), .ZN(
        n13456) );
  OAI22_X1 U14484 ( .A1(n14822), .A2(n13456), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12070), .ZN(n12071) );
  AOI211_X1 U14485 ( .C1(n12073), .C2(n14829), .A(n12072), .B(n12071), .ZN(
        n12079) );
  AOI22_X1 U14486 ( .A1(n12074), .A2(n13148), .B1(n13167), .B2(n13194), .ZN(
        n12076) );
  OR3_X1 U14487 ( .A1(n12077), .A2(n12076), .A3(n12075), .ZN(n12078) );
  OAI211_X1 U14488 ( .C1(n13026), .C2(n14824), .A(n12079), .B(n12078), .ZN(
        P2_U3200) );
  OAI21_X1 U14489 ( .B1(n12248), .B2(n13915), .A(n12264), .ZN(n12080) );
  NAND2_X1 U14490 ( .A1(n12080), .A2(n12249), .ZN(n12083) );
  NAND2_X1 U14491 ( .A1(n12249), .A2(n12247), .ZN(n12081) );
  NAND2_X1 U14492 ( .A1(n12081), .A2(n12255), .ZN(n12082) );
  NAND2_X1 U14493 ( .A1(n12274), .A2(n12086), .ZN(n12087) );
  NAND3_X1 U14494 ( .A1(n12087), .A2(n12273), .A3(n12094), .ZN(n12102) );
  MUX2_X1 U14495 ( .A(n12090), .B(n12089), .S(n12239), .Z(n12098) );
  INV_X1 U14496 ( .A(n12091), .ZN(n12093) );
  NAND3_X1 U14497 ( .A1(n12096), .A2(n12239), .A3(n12095), .ZN(n12097) );
  INV_X1 U14498 ( .A(n12100), .ZN(n12101) );
  OAI211_X1 U14499 ( .C1(n12103), .C2(n12102), .A(n12101), .B(n14714), .ZN(
        n12109) );
  NAND2_X1 U14500 ( .A1(n14724), .A2(n12239), .ZN(n12107) );
  NAND2_X1 U14501 ( .A1(n12105), .A2(n12227), .ZN(n12106) );
  MUX2_X1 U14502 ( .A(n12107), .B(n12106), .S(n13859), .Z(n12108) );
  NAND2_X1 U14503 ( .A1(n12109), .A2(n12108), .ZN(n12112) );
  MUX2_X1 U14504 ( .A(n14598), .B(n12110), .S(n12239), .Z(n12113) );
  MUX2_X1 U14505 ( .A(n12110), .B(n14598), .S(n12239), .Z(n12111) );
  MUX2_X1 U14506 ( .A(n14704), .B(n13858), .S(n12239), .Z(n12116) );
  MUX2_X1 U14507 ( .A(n13858), .B(n14704), .S(n12239), .Z(n12114) );
  MUX2_X1 U14508 ( .A(n14762), .B(n13857), .S(n12227), .Z(n12118) );
  MUX2_X1 U14509 ( .A(n14762), .B(n13857), .S(n12239), .Z(n12117) );
  MUX2_X1 U14510 ( .A(n14681), .B(n13856), .S(n12239), .Z(n12122) );
  NAND2_X1 U14511 ( .A1(n12121), .A2(n12122), .ZN(n12120) );
  MUX2_X1 U14512 ( .A(n13856), .B(n14681), .S(n12239), .Z(n12119) );
  NAND2_X1 U14513 ( .A1(n12120), .A2(n12119), .ZN(n12126) );
  INV_X1 U14514 ( .A(n12121), .ZN(n12124) );
  INV_X1 U14515 ( .A(n12122), .ZN(n12123) );
  NAND2_X1 U14516 ( .A1(n12124), .A2(n12123), .ZN(n12125) );
  NAND2_X1 U14517 ( .A1(n12126), .A2(n12125), .ZN(n12129) );
  MUX2_X1 U14518 ( .A(n13855), .B(n12127), .S(n12239), .Z(n12130) );
  MUX2_X1 U14519 ( .A(n13855), .B(n12127), .S(n12227), .Z(n12128) );
  MUX2_X1 U14520 ( .A(n13854), .B(n14665), .S(n12227), .Z(n12134) );
  MUX2_X1 U14521 ( .A(n13854), .B(n14665), .S(n12239), .Z(n12131) );
  NAND2_X1 U14522 ( .A1(n12132), .A2(n12131), .ZN(n12137) );
  INV_X1 U14523 ( .A(n12133), .ZN(n12135) );
  NAND2_X1 U14524 ( .A1(n12135), .A2(n7145), .ZN(n12136) );
  MUX2_X1 U14525 ( .A(n13853), .B(n14478), .S(n12239), .Z(n12139) );
  MUX2_X1 U14526 ( .A(n13853), .B(n14478), .S(n12227), .Z(n12138) );
  MUX2_X1 U14527 ( .A(n13852), .B(n14521), .S(n12227), .Z(n12142) );
  MUX2_X1 U14528 ( .A(n13852), .B(n14521), .S(n12239), .Z(n12140) );
  INV_X1 U14529 ( .A(n12141), .ZN(n12144) );
  INV_X1 U14530 ( .A(n12142), .ZN(n12143) );
  NAND2_X1 U14531 ( .A1(n12144), .A2(n12143), .ZN(n12145) );
  NAND2_X1 U14532 ( .A1(n12146), .A2(n12145), .ZN(n12149) );
  MUX2_X1 U14533 ( .A(n13851), .B(n12147), .S(n12239), .Z(n12150) );
  MUX2_X1 U14534 ( .A(n13851), .B(n12147), .S(n12227), .Z(n12148) );
  MUX2_X1 U14535 ( .A(n14114), .B(n12151), .S(n12227), .Z(n12154) );
  MUX2_X1 U14536 ( .A(n12152), .B(n14552), .S(n12239), .Z(n12153) );
  NAND2_X1 U14537 ( .A1(n12160), .A2(n12155), .ZN(n12158) );
  NAND2_X1 U14538 ( .A1(n12159), .A2(n12156), .ZN(n12157) );
  MUX2_X1 U14539 ( .A(n12158), .B(n12157), .S(n12239), .Z(n12162) );
  MUX2_X1 U14540 ( .A(n12160), .B(n12159), .S(n12227), .Z(n12161) );
  MUX2_X1 U14541 ( .A(n13850), .B(n14531), .S(n12239), .Z(n12180) );
  NAND2_X1 U14542 ( .A1(n12180), .A2(n14497), .ZN(n12164) );
  NAND2_X1 U14543 ( .A1(n12163), .A2(n12239), .ZN(n12166) );
  AOI21_X1 U14544 ( .B1(n12164), .B2(n12166), .A(n14104), .ZN(n12171) );
  NAND2_X1 U14545 ( .A1(n12180), .A2(n12167), .ZN(n12165) );
  OR2_X1 U14546 ( .A1(n14531), .A2(n12239), .ZN(n12172) );
  AOI21_X1 U14547 ( .B1(n12165), .B2(n12172), .A(n14192), .ZN(n12170) );
  NAND2_X1 U14548 ( .A1(n14497), .A2(n12227), .ZN(n12173) );
  OR2_X1 U14549 ( .A1(n14531), .A2(n12173), .ZN(n12169) );
  INV_X1 U14550 ( .A(n12166), .ZN(n12176) );
  NAND2_X1 U14551 ( .A1(n12176), .A2(n12167), .ZN(n12168) );
  NAND2_X1 U14552 ( .A1(n12169), .A2(n12168), .ZN(n12179) );
  INV_X1 U14553 ( .A(n12172), .ZN(n12175) );
  INV_X1 U14554 ( .A(n12173), .ZN(n12174) );
  AOI21_X1 U14555 ( .B1(n12180), .B2(n12175), .A(n12174), .ZN(n12183) );
  NAND2_X1 U14556 ( .A1(n12180), .A2(n12176), .ZN(n12177) );
  OAI21_X1 U14557 ( .B1(n12227), .B2(n14497), .A(n12177), .ZN(n12178) );
  NAND2_X1 U14558 ( .A1(n12178), .A2(n14192), .ZN(n12182) );
  NAND2_X1 U14559 ( .A1(n12180), .A2(n12179), .ZN(n12181) );
  OAI211_X1 U14560 ( .C1(n12183), .C2(n14192), .A(n12182), .B(n12181), .ZN(
        n12184) );
  INV_X1 U14561 ( .A(n12184), .ZN(n12185) );
  MUX2_X1 U14562 ( .A(n12187), .B(n14188), .S(n12227), .Z(n12188) );
  NAND2_X1 U14563 ( .A1(n12191), .A2(n12190), .ZN(n12192) );
  MUX2_X1 U14564 ( .A(n12194), .B(n12193), .S(n12239), .Z(n12195) );
  MUX2_X1 U14565 ( .A(n14034), .B(n14177), .S(n12239), .Z(n12197) );
  MUX2_X1 U14566 ( .A(n14067), .B(n14058), .S(n12227), .Z(n12196) );
  MUX2_X1 U14567 ( .A(n14044), .B(n14050), .S(n12239), .Z(n12200) );
  MUX2_X1 U14568 ( .A(n14050), .B(n14044), .S(n12239), .Z(n12198) );
  NAND2_X1 U14569 ( .A1(n12199), .A2(n12198), .ZN(n12202) );
  NAND2_X1 U14570 ( .A1(n6622), .A2(n7150), .ZN(n12201) );
  MUX2_X1 U14571 ( .A(n14032), .B(n14165), .S(n12239), .Z(n12204) );
  MUX2_X1 U14572 ( .A(n14032), .B(n14165), .S(n12227), .Z(n12203) );
  MUX2_X1 U14573 ( .A(n13848), .B(n14160), .S(n12104), .Z(n12207) );
  MUX2_X1 U14574 ( .A(n13848), .B(n14160), .S(n12239), .Z(n12205) );
  MUX2_X1 U14575 ( .A(n13847), .B(n14155), .S(n12239), .Z(n12209) );
  MUX2_X1 U14576 ( .A(n13847), .B(n14155), .S(n12104), .Z(n12208) );
  MUX2_X1 U14577 ( .A(n13846), .B(n14147), .S(n12104), .Z(n12213) );
  NAND2_X1 U14578 ( .A1(n12212), .A2(n12213), .ZN(n12211) );
  MUX2_X1 U14579 ( .A(n13846), .B(n14147), .S(n12239), .Z(n12210) );
  NAND2_X1 U14580 ( .A1(n12211), .A2(n12210), .ZN(n12217) );
  INV_X1 U14581 ( .A(n12212), .ZN(n12215) );
  INV_X1 U14582 ( .A(n12213), .ZN(n12214) );
  NAND2_X1 U14583 ( .A1(n12215), .A2(n12214), .ZN(n12216) );
  MUX2_X1 U14584 ( .A(n13845), .B(n13960), .S(n12239), .Z(n12219) );
  MUX2_X1 U14585 ( .A(n13845), .B(n13960), .S(n12227), .Z(n12218) );
  MUX2_X1 U14586 ( .A(n13844), .B(n14137), .S(n12104), .Z(n12222) );
  MUX2_X1 U14587 ( .A(n13844), .B(n14137), .S(n12239), .Z(n12220) );
  INV_X1 U14588 ( .A(n12221), .ZN(n12224) );
  INV_X1 U14589 ( .A(n12222), .ZN(n12223) );
  NAND2_X1 U14590 ( .A1(n12224), .A2(n12223), .ZN(n12225) );
  NAND2_X1 U14591 ( .A1(n12226), .A2(n12225), .ZN(n12229) );
  MUX2_X1 U14592 ( .A(n13843), .B(n12344), .S(n12239), .Z(n12230) );
  MUX2_X1 U14593 ( .A(n13843), .B(n12344), .S(n12227), .Z(n12228) );
  MUX2_X1 U14594 ( .A(n13842), .B(n12231), .S(n12104), .Z(n12235) );
  INV_X1 U14595 ( .A(n13842), .ZN(n12233) );
  MUX2_X1 U14596 ( .A(n12233), .B(n12232), .S(n12239), .Z(n12234) );
  OR2_X1 U14597 ( .A1(n7673), .A2(n14217), .ZN(n12237) );
  NAND2_X1 U14598 ( .A1(n12299), .A2(n12239), .ZN(n12254) );
  INV_X1 U14599 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n12240) );
  NOR2_X1 U14600 ( .A1(n12241), .A2(n12240), .ZN(n12246) );
  INV_X1 U14601 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n13919) );
  NOR2_X1 U14602 ( .A1(n12242), .A2(n13919), .ZN(n12245) );
  INV_X1 U14603 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n12243) );
  NOR2_X1 U14604 ( .A1(n6541), .A2(n12243), .ZN(n12244) );
  NAND2_X1 U14605 ( .A1(n13920), .A2(n12104), .ZN(n12251) );
  NAND3_X1 U14606 ( .A1(n12249), .A2(n12248), .A3(n12247), .ZN(n12250) );
  NAND2_X1 U14607 ( .A1(n12251), .A2(n12250), .ZN(n12252) );
  NAND2_X1 U14608 ( .A1(n12252), .A2(n13841), .ZN(n12253) );
  NAND2_X1 U14609 ( .A1(n12254), .A2(n12253), .ZN(n12258) );
  OAI21_X1 U14610 ( .B1(n13920), .B2(n12255), .A(n13841), .ZN(n12256) );
  MUX2_X1 U14611 ( .A(n12256), .B(n14134), .S(n12104), .Z(n12257) );
  NAND2_X1 U14612 ( .A1(n13683), .A2(n12260), .ZN(n12262) );
  INV_X1 U14613 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14215) );
  OR2_X1 U14614 ( .A1(n7673), .A2(n14215), .ZN(n12261) );
  OR2_X1 U14615 ( .A1(n13923), .A2(n12104), .ZN(n12309) );
  INV_X1 U14616 ( .A(n13920), .ZN(n12268) );
  NAND2_X1 U14617 ( .A1(n12264), .A2(n12263), .ZN(n12266) );
  NAND2_X1 U14618 ( .A1(n12266), .A2(n12265), .ZN(n12316) );
  AND2_X1 U14619 ( .A1(n12316), .A2(n12314), .ZN(n12304) );
  OAI21_X1 U14620 ( .B1(n12309), .B2(n12268), .A(n12304), .ZN(n12267) );
  INV_X1 U14621 ( .A(n12267), .ZN(n12270) );
  NOR2_X1 U14622 ( .A1(n14131), .A2(n12239), .ZN(n12307) );
  XOR2_X1 U14623 ( .A(n13920), .B(n14131), .Z(n12315) );
  NAND2_X1 U14624 ( .A1(n12272), .A2(n12271), .ZN(n14106) );
  NAND4_X1 U14625 ( .A1(n12273), .A2(n12274), .A3(n12275), .A4(n14714), .ZN(
        n12277) );
  NOR3_X1 U14626 ( .A1(n12277), .A2(n12276), .A3(n14689), .ZN(n12280) );
  NAND4_X1 U14627 ( .A1(n12281), .A2(n12280), .A3(n12279), .A4(n12278), .ZN(
        n12282) );
  NOR4_X1 U14628 ( .A1(n12284), .A2(n12283), .A3(n14523), .A4(n12282), .ZN(
        n12287) );
  NAND4_X1 U14629 ( .A1(n14106), .A2(n12287), .A3(n12286), .A4(n12285), .ZN(
        n12289) );
  NOR4_X1 U14630 ( .A1(n14503), .A2(n12290), .A3(n12289), .A4(n12288), .ZN(
        n12291) );
  NAND4_X1 U14631 ( .A1(n14056), .A2(n14074), .A3(n12291), .A4(n14079), .ZN(
        n12292) );
  NOR4_X1 U14632 ( .A1(n12294), .A2(n12293), .A3(n14027), .A4(n12292), .ZN(
        n12295) );
  NAND3_X1 U14633 ( .A1(n12295), .A2(n13994), .A3(n14002), .ZN(n12296) );
  NOR4_X1 U14634 ( .A1(n12298), .A2(n12297), .A3(n13946), .A4(n12296), .ZN(
        n12302) );
  XNOR2_X1 U14635 ( .A(n12299), .B(n13841), .ZN(n12300) );
  NAND4_X1 U14636 ( .A1(n12315), .A2(n12302), .A3(n12301), .A4(n12300), .ZN(
        n12303) );
  NOR2_X1 U14637 ( .A1(n13920), .A2(n12316), .ZN(n12308) );
  INV_X1 U14638 ( .A(n12304), .ZN(n12305) );
  NOR4_X1 U14639 ( .A1(n12307), .A2(n14131), .A3(n13920), .A4(n12305), .ZN(
        n12306) );
  AOI21_X1 U14640 ( .B1(n12308), .B2(n12307), .A(n12306), .ZN(n12313) );
  INV_X1 U14641 ( .A(n12309), .ZN(n12310) );
  XOR2_X1 U14642 ( .A(n12316), .B(n12310), .Z(n12311) );
  NAND4_X1 U14643 ( .A1(n12311), .A2(n14131), .A3(n13920), .A4(n12314), .ZN(
        n12312) );
  INV_X1 U14644 ( .A(n12315), .ZN(n12317) );
  NOR2_X1 U14645 ( .A1(n12317), .A2(n12316), .ZN(n12318) );
  NOR3_X1 U14646 ( .A1(n12321), .A2(n6538), .A3(n14696), .ZN(n12323) );
  OAI21_X1 U14647 ( .B1(n12324), .B2(n14227), .A(P1_B_REG_SCAN_IN), .ZN(n12322) );
  OAI22_X1 U14648 ( .A1(n6587), .A2(n12324), .B1(n12323), .B2(n12322), .ZN(
        P1_U3242) );
  INV_X1 U14649 ( .A(n12325), .ZN(n12326) );
  OAI222_X1 U14650 ( .A1(P3_U3151), .A2(n12328), .B1(n13023), .B2(n12327), 
        .C1(n13021), .C2(n12326), .ZN(P3_U3267) );
  OAI22_X1 U14651 ( .A1(n12336), .A2(n12331), .B1(n12335), .B2(n12330), .ZN(
        n12333) );
  XNOR2_X1 U14652 ( .A(n12333), .B(n12332), .ZN(n12338) );
  OAI22_X1 U14653 ( .A1(n12336), .A2(n10660), .B1(n12335), .B2(n12334), .ZN(
        n12337) );
  XNOR2_X1 U14654 ( .A(n12338), .B(n12337), .ZN(n12339) );
  AOI22_X1 U14655 ( .A1(n13814), .A2(n13844), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12341) );
  NAND2_X1 U14656 ( .A1(n13789), .A2(n13842), .ZN(n12340) );
  OAI211_X1 U14657 ( .C1(n14606), .C2(n12342), .A(n12341), .B(n12340), .ZN(
        n12343) );
  AOI21_X1 U14658 ( .B1(n12344), .B2(n13794), .A(n12343), .ZN(n12345) );
  OAI21_X1 U14659 ( .B1(n12346), .B2(n14593), .A(n12345), .ZN(P1_U3220) );
  INV_X1 U14660 ( .A(n12347), .ZN(n12357) );
  AOI22_X1 U14661 ( .A1(n13159), .A2(n12348), .B1(P2_REG3_REG_5__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12349) );
  OAI21_X1 U14662 ( .B1(n12350), .B2(n13133), .A(n12349), .ZN(n12356) );
  AOI22_X1 U14663 ( .A1(n13167), .A2(n13205), .B1(n13148), .B2(n12351), .ZN(
        n12353) );
  NOR3_X1 U14664 ( .A1(n12354), .A2(n12353), .A3(n12352), .ZN(n12355) );
  AOI211_X1 U14665 ( .C1(n13174), .C2(n12357), .A(n12356), .B(n12355), .ZN(
        n12358) );
  OAI21_X1 U14666 ( .B1(n12359), .B2(n14824), .A(n12358), .ZN(P2_U3199) );
  INV_X1 U14667 ( .A(n12362), .ZN(n12364) );
  XNOR2_X1 U14668 ( .A(n14374), .B(n12386), .ZN(n12366) );
  XNOR2_X1 U14669 ( .A(n12366), .B(n12542), .ZN(n14368) );
  XNOR2_X1 U14670 ( .A(n13004), .B(n12386), .ZN(n12367) );
  XNOR2_X1 U14671 ( .A(n12367), .B(n12476), .ZN(n12540) );
  XNOR2_X1 U14672 ( .A(n12998), .B(n12386), .ZN(n12368) );
  XNOR2_X1 U14673 ( .A(n12368), .B(n12855), .ZN(n12474) );
  INV_X1 U14674 ( .A(n12368), .ZN(n12369) );
  XNOR2_X1 U14675 ( .A(n12992), .B(n12386), .ZN(n12370) );
  XNOR2_X1 U14676 ( .A(n12370), .B(n12371), .ZN(n12482) );
  XNOR2_X1 U14677 ( .A(n12986), .B(n12386), .ZN(n12372) );
  XNOR2_X1 U14678 ( .A(n12372), .B(n12833), .ZN(n12520) );
  INV_X1 U14679 ( .A(n12372), .ZN(n12373) );
  XNOR2_X1 U14680 ( .A(n12982), .B(n12386), .ZN(n12374) );
  XNOR2_X1 U14681 ( .A(n12374), .B(n12824), .ZN(n12449) );
  INV_X1 U14682 ( .A(n12374), .ZN(n12375) );
  XNOR2_X1 U14683 ( .A(n12972), .B(n12386), .ZN(n12377) );
  XNOR2_X1 U14684 ( .A(n12377), .B(n12555), .ZN(n12504) );
  XNOR2_X1 U14685 ( .A(n12966), .B(n10969), .ZN(n12378) );
  NOR2_X1 U14686 ( .A1(n12378), .A2(n12796), .ZN(n12379) );
  AOI21_X1 U14687 ( .B1(n12378), .B2(n12796), .A(n12379), .ZN(n12457) );
  XNOR2_X1 U14688 ( .A(n12960), .B(n12386), .ZN(n12381) );
  NAND2_X1 U14689 ( .A1(n12380), .A2(n12381), .ZN(n12385) );
  INV_X1 U14690 ( .A(n12380), .ZN(n12383) );
  INV_X1 U14691 ( .A(n12381), .ZN(n12382) );
  NAND2_X1 U14692 ( .A1(n12383), .A2(n12382), .ZN(n12384) );
  XNOR2_X1 U14693 ( .A(n12954), .B(n12386), .ZN(n12387) );
  XNOR2_X1 U14694 ( .A(n12887), .B(n12386), .ZN(n12389) );
  NAND2_X1 U14695 ( .A1(n12389), .A2(n12763), .ZN(n12467) );
  INV_X1 U14696 ( .A(n12389), .ZN(n12390) );
  NAND2_X1 U14697 ( .A1(n12390), .A2(n12738), .ZN(n12391) );
  NAND2_X1 U14698 ( .A1(n12494), .A2(n12467), .ZN(n12397) );
  XNOR2_X1 U14699 ( .A(n12944), .B(n12386), .ZN(n12394) );
  NAND2_X1 U14700 ( .A1(n12394), .A2(n12393), .ZN(n12398) );
  INV_X1 U14701 ( .A(n12394), .ZN(n12395) );
  NAND2_X1 U14702 ( .A1(n12395), .A2(n12553), .ZN(n12396) );
  NAND2_X1 U14703 ( .A1(n12397), .A2(n12465), .ZN(n12469) );
  XNOR2_X1 U14704 ( .A(n12880), .B(n10969), .ZN(n12399) );
  NOR2_X1 U14705 ( .A1(n12399), .A2(n12739), .ZN(n12400) );
  AOI21_X1 U14706 ( .B1(n12399), .B2(n12739), .A(n12400), .ZN(n12530) );
  NAND2_X1 U14707 ( .A1(n12529), .A2(n12530), .ZN(n12528) );
  INV_X1 U14708 ( .A(n12400), .ZN(n12401) );
  XNOR2_X1 U14709 ( .A(n12433), .B(n10969), .ZN(n12402) );
  NOR2_X1 U14710 ( .A1(n12402), .A2(n12552), .ZN(n12403) );
  AOI21_X1 U14711 ( .B1(n12402), .B2(n12552), .A(n12403), .ZN(n12435) );
  XNOR2_X1 U14712 ( .A(n12702), .B(n12386), .ZN(n12404) );
  OR2_X1 U14713 ( .A1(n12405), .A2(n15241), .ZN(n12408) );
  OR2_X1 U14714 ( .A1(n12406), .A2(n15243), .ZN(n12407) );
  NAND2_X1 U14715 ( .A1(n12408), .A2(n12407), .ZN(n12706) );
  INV_X1 U14716 ( .A(n12533), .ZN(n14370) );
  AOI22_X1 U14717 ( .A1(n12706), .A2(n14370), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12409) );
  OAI21_X1 U14718 ( .B1(n14379), .B2(n12701), .A(n12409), .ZN(n12410) );
  AOI21_X1 U14719 ( .B1(n12872), .B2(n12548), .A(n12410), .ZN(n12411) );
  OAI21_X1 U14720 ( .B1(n12412), .B2(n12550), .A(n12411), .ZN(P3_U3160) );
  INV_X1 U14721 ( .A(SI_30_), .ZN(n12415) );
  INV_X1 U14722 ( .A(n12413), .ZN(n12414) );
  OAI222_X1 U14723 ( .A1(P3_U3151), .A2(n12416), .B1(n13023), .B2(n12415), 
        .C1(n13021), .C2(n12414), .ZN(P3_U3265) );
  OAI222_X1 U14724 ( .A1(n12419), .A2(P2_U3088), .B1(n13708), .B2(n12418), 
        .C1(n12417), .C2(n13705), .ZN(P2_U3306) );
  NAND3_X1 U14725 ( .A1(n12420), .A2(n13167), .A3(n13199), .ZN(n12421) );
  OAI21_X1 U14726 ( .B1(n12422), .B2(n14824), .A(n12421), .ZN(n12425) );
  INV_X1 U14727 ( .A(n12423), .ZN(n12424) );
  NAND2_X1 U14728 ( .A1(n12425), .A2(n12424), .ZN(n12431) );
  NOR2_X1 U14729 ( .A1(n14832), .A2(n13522), .ZN(n12429) );
  OAI22_X1 U14730 ( .A1(n14822), .A2(n12427), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12426), .ZN(n12428) );
  AOI211_X1 U14731 ( .C1(n13526), .C2(n14829), .A(n12429), .B(n12428), .ZN(
        n12430) );
  OAI211_X1 U14732 ( .C1(n12432), .C2(n14824), .A(n12431), .B(n12430), .ZN(
        P2_U3208) );
  NAND2_X1 U14733 ( .A1(n12436), .A2(n14376), .ZN(n12442) );
  INV_X1 U14734 ( .A(n12437), .ZN(n12718) );
  AOI22_X1 U14735 ( .A1(n15259), .A2(n12438), .B1(n12739), .B2(n15256), .ZN(
        n12713) );
  OAI22_X1 U14736 ( .A1(n12713), .A2(n12533), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12439), .ZN(n12440) );
  AOI21_X1 U14737 ( .B1(n12718), .B2(n12535), .A(n12440), .ZN(n12441) );
  OAI211_X1 U14738 ( .C1(n12937), .C2(n14373), .A(n12442), .B(n12441), .ZN(
        P3_U3154) );
  AOI21_X1 U14739 ( .B1(n12776), .B2(n12443), .A(n6571), .ZN(n12448) );
  AOI22_X1 U14740 ( .A1(n12522), .A2(n12554), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12445) );
  NAND2_X1 U14741 ( .A1(n12545), .A2(n12738), .ZN(n12444) );
  OAI211_X1 U14742 ( .C1(n14379), .C2(n12769), .A(n12445), .B(n12444), .ZN(
        n12446) );
  AOI21_X1 U14743 ( .B1(n12954), .B2(n12548), .A(n12446), .ZN(n12447) );
  OAI21_X1 U14744 ( .B1(n12448), .B2(n12550), .A(n12447), .ZN(P3_U3156) );
  XNOR2_X1 U14745 ( .A(n12450), .B(n12449), .ZN(n12455) );
  AOI22_X1 U14746 ( .A1(n12522), .A2(n12833), .B1(P3_REG3_REG_19__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12451) );
  OAI21_X1 U14747 ( .B1(n12808), .B2(n12507), .A(n12451), .ZN(n12453) );
  NOR2_X1 U14748 ( .A1(n12982), .A2(n14373), .ZN(n12452) );
  AOI211_X1 U14749 ( .C1(n12814), .C2(n12535), .A(n12453), .B(n12452), .ZN(
        n12454) );
  OAI21_X1 U14750 ( .B1(n12455), .B2(n12550), .A(n12454), .ZN(P3_U3159) );
  OAI21_X1 U14751 ( .B1(n12457), .B2(n6661), .A(n12456), .ZN(n12458) );
  NAND2_X1 U14752 ( .A1(n12458), .A2(n14376), .ZN(n12462) );
  OAI22_X1 U14753 ( .A1(n12808), .A2(n15243), .B1(n12764), .B2(n15241), .ZN(
        n12786) );
  AOI22_X1 U14754 ( .A1(n12786), .A2(n14370), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12461) );
  NAND2_X1 U14755 ( .A1(n12966), .A2(n12548), .ZN(n12460) );
  NAND2_X1 U14756 ( .A1(n12535), .A2(n12789), .ZN(n12459) );
  NAND4_X1 U14757 ( .A1(n12462), .A2(n12461), .A3(n12460), .A4(n12459), .ZN(
        P3_U3163) );
  AOI22_X1 U14758 ( .A1(n12522), .A2(n12738), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12464) );
  NAND2_X1 U14759 ( .A1(n12545), .A2(n12739), .ZN(n12463) );
  OAI211_X1 U14760 ( .C1(n14379), .C2(n12742), .A(n12464), .B(n12463), .ZN(
        n12471) );
  INV_X1 U14761 ( .A(n12465), .ZN(n12466) );
  NAND3_X1 U14762 ( .A1(n12494), .A2(n12467), .A3(n12466), .ZN(n12468) );
  AOI21_X1 U14763 ( .B1(n12469), .B2(n12468), .A(n12550), .ZN(n12470) );
  AOI211_X1 U14764 ( .C1(n12944), .C2(n12548), .A(n12471), .B(n12470), .ZN(
        n12472) );
  INV_X1 U14765 ( .A(n12472), .ZN(P3_U3165) );
  XNOR2_X1 U14766 ( .A(n12473), .B(n12474), .ZN(n12481) );
  OAI22_X1 U14767 ( .A1(n12543), .A2(n12476), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12475), .ZN(n12477) );
  AOI21_X1 U14768 ( .B1(n12545), .B2(n12844), .A(n12477), .ZN(n12478) );
  OAI21_X1 U14769 ( .B1(n12847), .B2(n14379), .A(n12478), .ZN(n12479) );
  AOI21_X1 U14770 ( .B1(n12998), .B2(n12548), .A(n12479), .ZN(n12480) );
  OAI21_X1 U14771 ( .B1(n12481), .B2(n12550), .A(n12480), .ZN(P3_U3166) );
  XNOR2_X1 U14772 ( .A(n12483), .B(n12482), .ZN(n12490) );
  INV_X1 U14773 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n12484) );
  OAI22_X1 U14774 ( .A1(n12543), .A2(n12485), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12484), .ZN(n12486) );
  AOI21_X1 U14775 ( .B1(n12545), .B2(n12833), .A(n12486), .ZN(n12487) );
  OAI21_X1 U14776 ( .B1(n12835), .B2(n14379), .A(n12487), .ZN(n12488) );
  AOI21_X1 U14777 ( .B1(n12992), .B2(n12548), .A(n12488), .ZN(n12489) );
  OAI21_X1 U14778 ( .B1(n12490), .B2(n12550), .A(n12489), .ZN(P3_U3168) );
  INV_X1 U14779 ( .A(n12887), .ZN(n12502) );
  INV_X1 U14780 ( .A(n12491), .ZN(n12493) );
  NOR3_X1 U14781 ( .A1(n6571), .A2(n12493), .A3(n12492), .ZN(n12496) );
  INV_X1 U14782 ( .A(n12494), .ZN(n12495) );
  OAI21_X1 U14783 ( .B1(n12496), .B2(n12495), .A(n14376), .ZN(n12501) );
  INV_X1 U14784 ( .A(n12751), .ZN(n12499) );
  AOI22_X1 U14785 ( .A1(n15256), .A2(n12776), .B1(n12553), .B2(n15259), .ZN(
        n12756) );
  INV_X1 U14786 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n12497) );
  OAI22_X1 U14787 ( .A1(n12756), .A2(n12533), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12497), .ZN(n12498) );
  AOI21_X1 U14788 ( .B1(n12499), .B2(n12535), .A(n12498), .ZN(n12500) );
  OAI211_X1 U14789 ( .C1(n12502), .C2(n14373), .A(n12501), .B(n12500), .ZN(
        P3_U3169) );
  XNOR2_X1 U14790 ( .A(n12503), .B(n12504), .ZN(n12511) );
  NAND2_X1 U14791 ( .A1(n12535), .A2(n12799), .ZN(n12506) );
  AOI22_X1 U14792 ( .A1(n12522), .A2(n12824), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12505) );
  OAI211_X1 U14793 ( .C1(n12508), .C2(n12507), .A(n12506), .B(n12505), .ZN(
        n12509) );
  AOI21_X1 U14794 ( .B1(n12972), .B2(n12548), .A(n12509), .ZN(n12510) );
  OAI21_X1 U14795 ( .B1(n12511), .B2(n12550), .A(n12510), .ZN(P3_U3173) );
  INV_X1 U14796 ( .A(n12512), .ZN(n12513) );
  AOI21_X1 U14797 ( .B1(n12554), .B2(n12514), .A(n12513), .ZN(n12519) );
  AOI22_X1 U14798 ( .A1(n12522), .A2(n12796), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12516) );
  NAND2_X1 U14799 ( .A1(n12545), .A2(n12776), .ZN(n12515) );
  OAI211_X1 U14800 ( .C1(n14379), .C2(n12779), .A(n12516), .B(n12515), .ZN(
        n12517) );
  AOI21_X1 U14801 ( .B1(n12960), .B2(n12548), .A(n12517), .ZN(n12518) );
  OAI21_X1 U14802 ( .B1(n12519), .B2(n12550), .A(n12518), .ZN(P3_U3175) );
  XNOR2_X1 U14803 ( .A(n12521), .B(n12520), .ZN(n12527) );
  AOI22_X1 U14804 ( .A1(n12522), .A2(n12844), .B1(P3_REG3_REG_18__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12524) );
  NAND2_X1 U14805 ( .A1(n12545), .A2(n12824), .ZN(n12523) );
  OAI211_X1 U14806 ( .C1(n14379), .C2(n12826), .A(n12524), .B(n12523), .ZN(
        n12525) );
  AOI21_X1 U14807 ( .B1(n12986), .B2(n12548), .A(n12525), .ZN(n12526) );
  OAI21_X1 U14808 ( .B1(n12527), .B2(n12550), .A(n12526), .ZN(P3_U3178) );
  INV_X1 U14809 ( .A(n12880), .ZN(n12539) );
  OAI21_X1 U14810 ( .B1(n12530), .B2(n12529), .A(n12528), .ZN(n12531) );
  NAND2_X1 U14811 ( .A1(n12531), .A2(n14376), .ZN(n12538) );
  INV_X1 U14812 ( .A(n12729), .ZN(n12536) );
  AOI22_X1 U14813 ( .A1(n15256), .A2(n12553), .B1(n12552), .B2(n15259), .ZN(
        n12727) );
  INV_X1 U14814 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n12532) );
  OAI22_X1 U14815 ( .A1(n12727), .A2(n12533), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12532), .ZN(n12534) );
  AOI21_X1 U14816 ( .B1(n12536), .B2(n12535), .A(n12534), .ZN(n12537) );
  OAI211_X1 U14817 ( .C1(n12539), .C2(n14373), .A(n12538), .B(n12537), .ZN(
        P3_U3180) );
  XNOR2_X1 U14818 ( .A(n12541), .B(n12540), .ZN(n12551) );
  OAI22_X1 U14819 ( .A1(n12543), .A2(n12542), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14386), .ZN(n12544) );
  AOI21_X1 U14820 ( .B1(n12545), .B2(n12855), .A(n12544), .ZN(n12546) );
  OAI21_X1 U14821 ( .B1(n14379), .B2(n12858), .A(n12546), .ZN(n12547) );
  AOI21_X1 U14822 ( .B1(n13004), .B2(n12548), .A(n12547), .ZN(n12549) );
  OAI21_X1 U14823 ( .B1(n12551), .B2(n12550), .A(n12549), .ZN(P3_U3181) );
  MUX2_X1 U14824 ( .A(n12683), .B(P3_DATAO_REG_31__SCAN_IN), .S(n12563), .Z(
        P3_U3522) );
  MUX2_X1 U14825 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12552), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14826 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12553), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14827 ( .A(n12738), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12563), .Z(
        P3_U3515) );
  MUX2_X1 U14828 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n12776), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U14829 ( .A(n12554), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12563), .Z(
        P3_U3513) );
  MUX2_X1 U14830 ( .A(n12796), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12563), .Z(
        P3_U3512) );
  MUX2_X1 U14831 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12555), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14832 ( .A(n12824), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12563), .Z(
        P3_U3510) );
  MUX2_X1 U14833 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12833), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14834 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12844), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14835 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12855), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14836 ( .A(n12856), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12563), .Z(
        P3_U3505) );
  MUX2_X1 U14837 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12556), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14838 ( .A(n12557), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12563), .Z(
        P3_U3503) );
  MUX2_X1 U14839 ( .A(n12558), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12563), .Z(
        P3_U3502) );
  MUX2_X1 U14840 ( .A(n12559), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12563), .Z(
        P3_U3501) );
  MUX2_X1 U14841 ( .A(n12560), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12563), .Z(
        P3_U3500) );
  MUX2_X1 U14842 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12561), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14843 ( .A(n15190), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12563), .Z(
        P3_U3498) );
  MUX2_X1 U14844 ( .A(n12562), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12563), .Z(
        P3_U3497) );
  MUX2_X1 U14845 ( .A(n15189), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12563), .Z(
        P3_U3496) );
  MUX2_X1 U14846 ( .A(n15217), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12563), .Z(
        P3_U3495) );
  MUX2_X1 U14847 ( .A(n15258), .B(P3_DATAO_REG_2__SCAN_IN), .S(n12563), .Z(
        P3_U3493) );
  MUX2_X1 U14848 ( .A(n12564), .B(P3_DATAO_REG_1__SCAN_IN), .S(n12563), .Z(
        P3_U3492) );
  NAND2_X1 U14849 ( .A1(n15169), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12662) );
  INV_X1 U14850 ( .A(n15151), .ZN(n12657) );
  INV_X1 U14851 ( .A(n15117), .ZN(n12650) );
  NAND2_X1 U14852 ( .A1(n12626), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n12565) );
  NAND2_X1 U14853 ( .A1(n12566), .A2(n12565), .ZN(n12567) );
  INV_X1 U14854 ( .A(n15014), .ZN(n12596) );
  XNOR2_X1 U14855 ( .A(n12567), .B(n12596), .ZN(n15003) );
  NAND2_X1 U14856 ( .A1(n15003), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n15006) );
  INV_X1 U14857 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n15200) );
  AOI22_X1 U14858 ( .A1(n12632), .A2(P3_REG2_REG_6__SCAN_IN), .B1(n15200), 
        .B2(n15028), .ZN(n15026) );
  NAND2_X1 U14859 ( .A1(n12569), .A2(n15052), .ZN(n12568) );
  INV_X1 U14860 ( .A(n12568), .ZN(n12570) );
  OAI21_X1 U14861 ( .B1(n12569), .B2(n15052), .A(n12568), .ZN(n15041) );
  NOR2_X1 U14862 ( .A1(n12624), .A2(n15041), .ZN(n15040) );
  NOR2_X1 U14863 ( .A1(n12570), .A2(n15040), .ZN(n15069) );
  AOI22_X1 U14864 ( .A1(n12640), .A2(P3_REG2_REG_8__SCAN_IN), .B1(n12622), 
        .B2(n15066), .ZN(n15068) );
  NAND2_X1 U14865 ( .A1(n12572), .A2(n15083), .ZN(n12571) );
  INV_X1 U14866 ( .A(n12571), .ZN(n12573) );
  OAI21_X1 U14867 ( .B1(n12572), .B2(n15083), .A(n12571), .ZN(n15078) );
  NOR2_X1 U14868 ( .A1(n12620), .A2(n15078), .ZN(n15077) );
  INV_X1 U14869 ( .A(n15100), .ZN(n12646) );
  AOI22_X1 U14870 ( .A1(n12646), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n11528), 
        .B2(n15100), .ZN(n15093) );
  NOR2_X1 U14871 ( .A1(n12650), .A2(n12574), .ZN(n12575) );
  NAND2_X1 U14872 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n15135), .ZN(n12576) );
  OAI21_X1 U14873 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n15135), .A(n12576), 
        .ZN(n15128) );
  NOR2_X1 U14874 ( .A1(n12657), .A2(n12577), .ZN(n12578) );
  OAI21_X1 U14875 ( .B1(n15169), .B2(P3_REG2_REG_14__SCAN_IN), .A(n12662), 
        .ZN(n15164) );
  AND2_X1 U14876 ( .A1(n14389), .A2(n12579), .ZN(n12580) );
  OR2_X1 U14877 ( .A1(n14399), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12582) );
  NAND2_X1 U14878 ( .A1(n14399), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12581) );
  AND2_X1 U14879 ( .A1(n12582), .A2(n12581), .ZN(n14409) );
  NAND2_X1 U14880 ( .A1(n14431), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12586) );
  INV_X1 U14881 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12584) );
  NAND2_X1 U14882 ( .A1(n12617), .A2(n12584), .ZN(n12585) );
  AND2_X1 U14883 ( .A1(n12586), .A2(n12585), .ZN(n14441) );
  AOI21_X1 U14884 ( .B1(P3_REG2_REG_18__SCAN_IN), .B2(n12617), .A(n14443), 
        .ZN(n12587) );
  MUX2_X1 U14885 ( .A(P3_REG2_REG_19__SCAN_IN), .B(n12811), .S(n12676), .Z(
        n12672) );
  XNOR2_X1 U14886 ( .A(n12587), .B(n12672), .ZN(n12680) );
  NAND2_X1 U14887 ( .A1(n15169), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12661) );
  NAND2_X1 U14888 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n15135), .ZN(n12605) );
  MUX2_X1 U14889 ( .A(P3_REG1_REG_12__SCAN_IN), .B(n12588), .S(n15135), .Z(
        n15131) );
  MUX2_X1 U14890 ( .A(P3_REG1_REG_10__SCAN_IN), .B(n12589), .S(n15100), .Z(
        n15096) );
  AOI22_X1 U14891 ( .A1(n12640), .A2(n12621), .B1(P3_REG1_REG_8__SCAN_IN), 
        .B2(n15066), .ZN(n15061) );
  OR2_X1 U14892 ( .A1(n12632), .A2(n12625), .ZN(n12598) );
  AOI22_X1 U14893 ( .A1(n12632), .A2(n12625), .B1(P3_REG1_REG_6__SCAN_IN), 
        .B2(n15028), .ZN(n15023) );
  INV_X1 U14894 ( .A(n12626), .ZN(n12591) );
  OAI22_X1 U14895 ( .A1(n12593), .A2(n12592), .B1(n12591), .B2(n12590), .ZN(
        n12594) );
  XNOR2_X1 U14896 ( .A(n12594), .B(n15014), .ZN(n15017) );
  INV_X1 U14897 ( .A(n12594), .ZN(n12595) );
  OAI22_X1 U14898 ( .A1(n15017), .A2(n12597), .B1(n12596), .B2(n12595), .ZN(
        n15024) );
  NAND2_X1 U14899 ( .A1(n15023), .A2(n15024), .ZN(n15022) );
  NAND2_X1 U14900 ( .A1(n12598), .A2(n15022), .ZN(n12599) );
  NAND2_X1 U14901 ( .A1(n12599), .A2(n15052), .ZN(n12600) );
  INV_X1 U14902 ( .A(n15052), .ZN(n12636) );
  XNOR2_X1 U14903 ( .A(n12636), .B(n12599), .ZN(n15044) );
  NAND2_X1 U14904 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n15044), .ZN(n15043) );
  NAND2_X1 U14905 ( .A1(n12600), .A2(n15043), .ZN(n15060) );
  NAND2_X1 U14906 ( .A1(n15061), .A2(n15060), .ZN(n15059) );
  OAI21_X1 U14907 ( .B1(n12640), .B2(n12621), .A(n15059), .ZN(n12601) );
  INV_X1 U14908 ( .A(n12601), .ZN(n12602) );
  INV_X1 U14909 ( .A(n15083), .ZN(n12643) );
  XNOR2_X1 U14910 ( .A(n12601), .B(n12643), .ZN(n15087) );
  NAND2_X1 U14911 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n15087), .ZN(n15086) );
  OAI21_X1 U14912 ( .B1(n12602), .B2(n12643), .A(n15086), .ZN(n15097) );
  NAND2_X1 U14913 ( .A1(n15096), .A2(n15097), .ZN(n15095) );
  OAI21_X1 U14914 ( .B1(n12646), .B2(n12589), .A(n15095), .ZN(n12603) );
  NAND2_X1 U14915 ( .A1(n15117), .A2(n12603), .ZN(n12604) );
  XNOR2_X1 U14916 ( .A(n12650), .B(n12603), .ZN(n15113) );
  NAND2_X1 U14917 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n15113), .ZN(n15112) );
  NAND2_X1 U14918 ( .A1(n12604), .A2(n15112), .ZN(n15132) );
  NAND2_X1 U14919 ( .A1(n15131), .A2(n15132), .ZN(n15130) );
  NAND2_X1 U14920 ( .A1(n12605), .A2(n15130), .ZN(n12606) );
  NAND2_X1 U14921 ( .A1(n15151), .A2(n12606), .ZN(n12607) );
  XNOR2_X1 U14922 ( .A(n12606), .B(n12657), .ZN(n15147) );
  NAND2_X1 U14923 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n15147), .ZN(n15146) );
  NAND2_X1 U14924 ( .A1(n12607), .A2(n15146), .ZN(n15167) );
  INV_X1 U14925 ( .A(n15169), .ZN(n12609) );
  NAND2_X1 U14926 ( .A1(n12609), .A2(n12608), .ZN(n12610) );
  AND2_X1 U14927 ( .A1(n12610), .A2(n12661), .ZN(n15168) );
  NAND2_X1 U14928 ( .A1(n15167), .A2(n15168), .ZN(n15166) );
  NAND2_X1 U14929 ( .A1(n12661), .A2(n15166), .ZN(n12611) );
  NAND2_X1 U14930 ( .A1(n14389), .A2(n12611), .ZN(n12612) );
  XOR2_X1 U14931 ( .A(n14389), .B(n12611), .Z(n14385) );
  NAND2_X1 U14932 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n14385), .ZN(n14384) );
  NAND2_X1 U14933 ( .A1(n12612), .A2(n14384), .ZN(n14406) );
  XNOR2_X1 U14934 ( .A(n14399), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n14405) );
  AOI22_X1 U14935 ( .A1(n14406), .A2(n14405), .B1(P3_REG1_REG_16__SCAN_IN), 
        .B2(n12613), .ZN(n12614) );
  INV_X1 U14936 ( .A(n12614), .ZN(n12615) );
  NAND2_X1 U14937 ( .A1(n12666), .A2(n12615), .ZN(n12616) );
  XOR2_X1 U14938 ( .A(n12666), .B(n12615), .Z(n14418) );
  NAND2_X1 U14939 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n14418), .ZN(n14417) );
  NAND2_X1 U14940 ( .A1(n12616), .A2(n14417), .ZN(n14434) );
  XNOR2_X1 U14941 ( .A(n14431), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n14433) );
  AOI22_X1 U14942 ( .A1(n14434), .A2(n14433), .B1(P3_REG1_REG_18__SCAN_IN), 
        .B2(n12617), .ZN(n12618) );
  XNOR2_X1 U14943 ( .A(n12676), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12669) );
  XNOR2_X1 U14944 ( .A(n12618), .B(n12669), .ZN(n12678) );
  MUX2_X1 U14945 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12670), .Z(n12667) );
  MUX2_X1 U14946 ( .A(n12846), .B(n12914), .S(n12670), .Z(n12665) );
  NOR2_X1 U14947 ( .A1(n12665), .A2(n14399), .ZN(n14400) );
  MUX2_X1 U14948 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n12670), .Z(n12645) );
  XNOR2_X1 U14949 ( .A(n12645), .B(n12646), .ZN(n15104) );
  MUX2_X1 U14950 ( .A(n12620), .B(n12619), .S(n12670), .Z(n12644) );
  MUX2_X1 U14951 ( .A(n12622), .B(n12621), .S(n12670), .Z(n12641) );
  NAND2_X1 U14952 ( .A1(n12641), .A2(n12640), .ZN(n12639) );
  INV_X1 U14953 ( .A(n12639), .ZN(n12642) );
  MUX2_X1 U14954 ( .A(n12624), .B(n12623), .S(n12670), .Z(n12637) );
  NAND2_X1 U14955 ( .A1(n12637), .A2(n12636), .ZN(n12635) );
  INV_X1 U14956 ( .A(n12635), .ZN(n12638) );
  MUX2_X1 U14957 ( .A(n15200), .B(n12625), .S(n12670), .Z(n12633) );
  NAND2_X1 U14958 ( .A1(n12633), .A2(n12632), .ZN(n12631) );
  INV_X1 U14959 ( .A(n12631), .ZN(n12634) );
  MUX2_X1 U14960 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12670), .Z(n12630) );
  NAND2_X1 U14961 ( .A1(n12630), .A2(n15014), .ZN(n15007) );
  NOR2_X1 U14962 ( .A1(n12630), .A2(n15014), .ZN(n15009) );
  AOI21_X1 U14963 ( .B1(n15011), .B2(n15007), .A(n15009), .ZN(n15032) );
  OAI21_X1 U14964 ( .B1(n12633), .B2(n12632), .A(n12631), .ZN(n15031) );
  NOR2_X1 U14965 ( .A1(n15032), .A2(n15031), .ZN(n15030) );
  NOR2_X1 U14966 ( .A1(n12634), .A2(n15030), .ZN(n15046) );
  OAI21_X1 U14967 ( .B1(n12637), .B2(n12636), .A(n12635), .ZN(n15047) );
  NOR2_X1 U14968 ( .A1(n15046), .A2(n15047), .ZN(n15045) );
  NOR2_X1 U14969 ( .A1(n12638), .A2(n15045), .ZN(n15063) );
  OAI21_X1 U14970 ( .B1(n12641), .B2(n12640), .A(n12639), .ZN(n15064) );
  NOR2_X1 U14971 ( .A1(n15063), .A2(n15064), .ZN(n15062) );
  XNOR2_X1 U14972 ( .A(n12644), .B(n12643), .ZN(n15081) );
  NAND2_X1 U14973 ( .A1(n15104), .A2(n15105), .ZN(n15103) );
  INV_X1 U14974 ( .A(n12645), .ZN(n12647) );
  NAND2_X1 U14975 ( .A1(n12647), .A2(n12646), .ZN(n12648) );
  NAND2_X1 U14976 ( .A1(n15103), .A2(n12648), .ZN(n15122) );
  MUX2_X1 U14977 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12670), .Z(n12649) );
  XNOR2_X1 U14978 ( .A(n12649), .B(n12650), .ZN(n15121) );
  NAND2_X1 U14979 ( .A1(n15122), .A2(n15121), .ZN(n15120) );
  INV_X1 U14980 ( .A(n12649), .ZN(n12651) );
  NAND2_X1 U14981 ( .A1(n12651), .A2(n12650), .ZN(n12652) );
  MUX2_X1 U14982 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12670), .Z(n12654) );
  XNOR2_X1 U14983 ( .A(n12654), .B(n12653), .ZN(n15139) );
  NAND2_X1 U14984 ( .A1(n12654), .A2(n15135), .ZN(n12655) );
  MUX2_X1 U14985 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12670), .Z(n12656) );
  XNOR2_X1 U14986 ( .A(n12656), .B(n15151), .ZN(n15157) );
  INV_X1 U14987 ( .A(n12656), .ZN(n12658) );
  NAND2_X1 U14988 ( .A1(n12658), .A2(n12657), .ZN(n12659) );
  INV_X1 U14989 ( .A(n15164), .ZN(n12660) );
  MUX2_X1 U14990 ( .A(n12660), .B(n15168), .S(n12670), .Z(n15180) );
  NAND2_X1 U14991 ( .A1(n15181), .A2(n15180), .ZN(n15179) );
  MUX2_X1 U14992 ( .A(n12662), .B(n12661), .S(n12670), .Z(n12663) );
  MUX2_X1 U14993 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12670), .Z(n14394) );
  NOR2_X1 U14994 ( .A1(n12664), .A2(n14392), .ZN(n14404) );
  NAND2_X1 U14995 ( .A1(n12665), .A2(n14399), .ZN(n14402) );
  OAI21_X1 U14996 ( .B1(n14400), .B2(n14404), .A(n14402), .ZN(n14421) );
  XNOR2_X1 U14997 ( .A(n12667), .B(n12666), .ZN(n14420) );
  NOR2_X1 U14998 ( .A1(n14421), .A2(n14420), .ZN(n14419) );
  AOI21_X1 U14999 ( .B1(n12667), .B2(n12666), .A(n14419), .ZN(n12668) );
  XNOR2_X1 U15000 ( .A(n12668), .B(n14431), .ZN(n14436) );
  MUX2_X1 U15001 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12670), .Z(n14437) );
  NOR2_X1 U15002 ( .A1(n14436), .A2(n14437), .ZN(n14435) );
  INV_X1 U15003 ( .A(n12669), .ZN(n12671) );
  MUX2_X1 U15004 ( .A(n12672), .B(n12671), .S(n12670), .Z(n12673) );
  NAND2_X1 U15005 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(P3_U3151), .ZN(n12675)
         );
  NAND2_X1 U15006 ( .A1(n15149), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12674) );
  OAI211_X1 U15007 ( .C1(n15170), .C2(n12676), .A(n12675), .B(n12674), .ZN(
        n12677) );
  OAI21_X1 U15008 ( .B1(n12680), .B2(n15184), .A(n12679), .ZN(P3_U3201) );
  INV_X1 U15009 ( .A(n12860), .ZN(n12816) );
  INV_X1 U15010 ( .A(n15273), .ZN(n12719) );
  INV_X1 U15011 ( .A(n12682), .ZN(n12684) );
  NAND2_X1 U15012 ( .A1(n12684), .A2(n12683), .ZN(n12922) );
  OR2_X1 U15013 ( .A1(n15268), .A2(n12685), .ZN(n12691) );
  OAI21_X1 U15014 ( .B1(n12719), .B2(n12922), .A(n12691), .ZN(n12687) );
  AOI21_X1 U15015 ( .B1(P3_REG2_REG_31__SCAN_IN), .B2(n12719), .A(n12687), 
        .ZN(n12686) );
  OAI21_X1 U15016 ( .B1(n12924), .B2(n12816), .A(n12686), .ZN(P3_U3202) );
  AOI21_X1 U15017 ( .B1(P3_REG2_REG_30__SCAN_IN), .B2(n12719), .A(n12687), 
        .ZN(n12688) );
  OAI21_X1 U15018 ( .B1(n12689), .B2(n12816), .A(n12688), .ZN(P3_U3203) );
  NAND2_X1 U15019 ( .A1(n12690), .A2(n15273), .ZN(n12696) );
  OAI21_X1 U15020 ( .B1(n15273), .B2(n12692), .A(n12691), .ZN(n12693) );
  AOI21_X1 U15021 ( .B1(n12694), .B2(n12860), .A(n12693), .ZN(n12695) );
  OAI211_X1 U15022 ( .C1(n12697), .C2(n12863), .A(n12696), .B(n12695), .ZN(
        P3_U3204) );
  OAI21_X1 U15023 ( .B1(n12700), .B2(n12699), .A(n12698), .ZN(n12869) );
  INV_X1 U15024 ( .A(n12872), .ZN(n12930) );
  OAI22_X1 U15025 ( .A1(n12930), .A2(n12816), .B1(n12701), .B2(n15268), .ZN(
        n12710) );
  NOR2_X1 U15026 ( .A1(n12703), .A2(n12702), .ZN(n12705) );
  INV_X1 U15027 ( .A(n12706), .ZN(n12707) );
  INV_X1 U15028 ( .A(n12711), .ZN(P3_U3205) );
  XNOR2_X1 U15029 ( .A(n12712), .B(n12716), .ZN(n12714) );
  OAI21_X1 U15030 ( .B1(n12714), .B2(n15249), .A(n12713), .ZN(n12875) );
  INV_X1 U15031 ( .A(n12875), .ZN(n12723) );
  OAI21_X1 U15032 ( .B1(n12717), .B2(n12716), .A(n12715), .ZN(n12876) );
  AOI22_X1 U15033 ( .A1(n12719), .A2(P3_REG2_REG_27__SCAN_IN), .B1(n15226), 
        .B2(n12718), .ZN(n12720) );
  OAI21_X1 U15034 ( .B1(n12937), .B2(n12816), .A(n12720), .ZN(n12721) );
  AOI21_X1 U15035 ( .B1(n12876), .B2(n12818), .A(n12721), .ZN(n12722) );
  OAI21_X1 U15036 ( .B1(n12723), .B2(n12719), .A(n12722), .ZN(P3_U3206) );
  XOR2_X1 U15037 ( .A(n12724), .B(n12726), .Z(n12941) );
  XOR2_X1 U15038 ( .A(n12726), .B(n12725), .Z(n12728) );
  OAI21_X1 U15039 ( .B1(n12728), .B2(n15249), .A(n12727), .ZN(n12879) );
  NAND2_X1 U15040 ( .A1(n12879), .A2(n15273), .ZN(n12733) );
  INV_X1 U15041 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12730) );
  OAI22_X1 U15042 ( .A1(n15273), .A2(n12730), .B1(n12729), .B2(n15268), .ZN(
        n12731) );
  AOI21_X1 U15043 ( .B1(n12880), .B2(n12860), .A(n12731), .ZN(n12732) );
  OAI211_X1 U15044 ( .C1(n12941), .C2(n12863), .A(n12733), .B(n12732), .ZN(
        P3_U3207) );
  XNOR2_X1 U15045 ( .A(n12735), .B(n12734), .ZN(n12947) );
  INV_X1 U15046 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n12741) );
  XNOR2_X1 U15047 ( .A(n12736), .B(n12737), .ZN(n12740) );
  AOI222_X1 U15048 ( .A1(n15262), .A2(n12740), .B1(n12739), .B2(n15259), .C1(
        n12738), .C2(n15256), .ZN(n12942) );
  MUX2_X1 U15049 ( .A(n12741), .B(n12942), .S(n15273), .Z(n12745) );
  INV_X1 U15050 ( .A(n12742), .ZN(n12743) );
  AOI22_X1 U15051 ( .A1(n12944), .A2(n12860), .B1(n15226), .B2(n12743), .ZN(
        n12744) );
  OAI211_X1 U15052 ( .C1(n12947), .C2(n12863), .A(n12745), .B(n12744), .ZN(
        P3_U3208) );
  NAND2_X1 U15053 ( .A1(n12746), .A2(n12747), .ZN(n12750) );
  INV_X1 U15054 ( .A(n12748), .ZN(n12749) );
  AOI21_X1 U15055 ( .B1(n12754), .B2(n12750), .A(n12749), .ZN(n12951) );
  INV_X1 U15056 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12752) );
  OAI22_X1 U15057 ( .A1(n15273), .A2(n12752), .B1(n12751), .B2(n15268), .ZN(
        n12753) );
  AOI21_X1 U15058 ( .B1(n12887), .B2(n12860), .A(n12753), .ZN(n12759) );
  XNOR2_X1 U15059 ( .A(n12755), .B(n12754), .ZN(n12757) );
  OAI21_X1 U15060 ( .B1(n12757), .B2(n15249), .A(n12756), .ZN(n12886) );
  NAND2_X1 U15061 ( .A1(n12886), .A2(n15273), .ZN(n12758) );
  OAI211_X1 U15062 ( .C1(n12951), .C2(n12863), .A(n12759), .B(n12758), .ZN(
        P3_U3209) );
  OAI21_X1 U15063 ( .B1(n12760), .B2(n12761), .A(n12746), .ZN(n12957) );
  AOI21_X1 U15064 ( .B1(n12762), .B2(n12761), .A(n15249), .ZN(n12767) );
  OAI22_X1 U15065 ( .A1(n12764), .A2(n15243), .B1(n12763), .B2(n15241), .ZN(
        n12765) );
  AOI21_X1 U15066 ( .B1(n12767), .B2(n12766), .A(n12765), .ZN(n12952) );
  MUX2_X1 U15067 ( .A(n12768), .B(n12952), .S(n15273), .Z(n12772) );
  INV_X1 U15068 ( .A(n12769), .ZN(n12770) );
  AOI22_X1 U15069 ( .A1(n12954), .A2(n12860), .B1(n15226), .B2(n12770), .ZN(
        n12771) );
  OAI211_X1 U15070 ( .C1(n12957), .C2(n12863), .A(n12772), .B(n12771), .ZN(
        P3_U3210) );
  XNOR2_X1 U15071 ( .A(n12773), .B(n12774), .ZN(n12963) );
  INV_X1 U15072 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n12778) );
  XNOR2_X1 U15073 ( .A(n12775), .B(n12774), .ZN(n12777) );
  AOI222_X1 U15074 ( .A1(n15262), .A2(n12777), .B1(n12796), .B2(n15256), .C1(
        n12776), .C2(n15259), .ZN(n12958) );
  MUX2_X1 U15075 ( .A(n12778), .B(n12958), .S(n15273), .Z(n12782) );
  INV_X1 U15076 ( .A(n12779), .ZN(n12780) );
  AOI22_X1 U15077 ( .A1(n12960), .A2(n12860), .B1(n15226), .B2(n12780), .ZN(
        n12781) );
  OAI211_X1 U15078 ( .C1(n12963), .C2(n12863), .A(n12782), .B(n12781), .ZN(
        P3_U3211) );
  XNOR2_X1 U15079 ( .A(n12783), .B(n12785), .ZN(n12969) );
  XNOR2_X1 U15080 ( .A(n12784), .B(n12785), .ZN(n12787) );
  AOI21_X1 U15081 ( .B1(n12787), .B2(n15262), .A(n12786), .ZN(n12964) );
  MUX2_X1 U15082 ( .A(n12788), .B(n12964), .S(n15273), .Z(n12791) );
  AOI22_X1 U15083 ( .A1(n12966), .A2(n12860), .B1(n15226), .B2(n12789), .ZN(
        n12790) );
  OAI211_X1 U15084 ( .C1(n12969), .C2(n12863), .A(n12791), .B(n12790), .ZN(
        P3_U3212) );
  OAI21_X1 U15085 ( .B1(n12793), .B2(n12794), .A(n12792), .ZN(n12976) );
  INV_X1 U15086 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12798) );
  XNOR2_X1 U15087 ( .A(n12795), .B(n12794), .ZN(n12797) );
  AOI222_X1 U15088 ( .A1(n15262), .A2(n12797), .B1(n12796), .B2(n15259), .C1(
        n12824), .C2(n15256), .ZN(n12970) );
  MUX2_X1 U15089 ( .A(n12798), .B(n12970), .S(n15273), .Z(n12801) );
  AOI22_X1 U15090 ( .A1(n12972), .A2(n12860), .B1(n15226), .B2(n12799), .ZN(
        n12800) );
  OAI211_X1 U15091 ( .C1(n12976), .C2(n12863), .A(n12801), .B(n12800), .ZN(
        P3_U3213) );
  INV_X1 U15092 ( .A(n12802), .ZN(n12806) );
  AOI21_X1 U15093 ( .B1(n12803), .B2(n12804), .A(n12812), .ZN(n12805) );
  NOR3_X1 U15094 ( .A1(n12806), .A2(n12805), .A3(n15249), .ZN(n12810) );
  OAI22_X1 U15095 ( .A1(n12808), .A2(n15241), .B1(n12807), .B2(n15243), .ZN(
        n12809) );
  NOR2_X1 U15096 ( .A1(n12810), .A2(n12809), .ZN(n12977) );
  MUX2_X1 U15097 ( .A(n12811), .B(n12977), .S(n15273), .Z(n12820) );
  XNOR2_X1 U15098 ( .A(n12813), .B(n12812), .ZN(n12979) );
  INV_X1 U15099 ( .A(n12814), .ZN(n12815) );
  OAI22_X1 U15100 ( .A1(n12982), .A2(n12816), .B1(n12815), .B2(n15268), .ZN(
        n12817) );
  AOI21_X1 U15101 ( .B1(n12979), .B2(n12818), .A(n12817), .ZN(n12819) );
  NAND2_X1 U15102 ( .A1(n12820), .A2(n12819), .ZN(P3_U3214) );
  XNOR2_X1 U15103 ( .A(n12822), .B(n12821), .ZN(n12987) );
  INV_X1 U15104 ( .A(n12987), .ZN(n12830) );
  OAI21_X1 U15105 ( .B1(n6657), .B2(n12823), .A(n12803), .ZN(n12825) );
  AOI222_X1 U15106 ( .A1(n15262), .A2(n12825), .B1(n12844), .B2(n15256), .C1(
        n12824), .C2(n15259), .ZN(n12984) );
  MUX2_X1 U15107 ( .A(n12584), .B(n12984), .S(n15273), .Z(n12829) );
  INV_X1 U15108 ( .A(n12826), .ZN(n12827) );
  AOI22_X1 U15109 ( .A1(n12986), .A2(n12860), .B1(n15226), .B2(n12827), .ZN(
        n12828) );
  OAI211_X1 U15110 ( .C1(n12830), .C2(n12863), .A(n12829), .B(n12828), .ZN(
        P3_U3215) );
  XNOR2_X1 U15111 ( .A(n12831), .B(n7345), .ZN(n12993) );
  INV_X1 U15112 ( .A(n12993), .ZN(n12839) );
  XNOR2_X1 U15113 ( .A(n12832), .B(n7345), .ZN(n12834) );
  AOI222_X1 U15114 ( .A1(n15262), .A2(n12834), .B1(n12855), .B2(n15256), .C1(
        n12833), .C2(n15259), .ZN(n12990) );
  MUX2_X1 U15115 ( .A(n14425), .B(n12990), .S(n15273), .Z(n12838) );
  INV_X1 U15116 ( .A(n12835), .ZN(n12836) );
  AOI22_X1 U15117 ( .A1(n12992), .A2(n12860), .B1(n15226), .B2(n12836), .ZN(
        n12837) );
  OAI211_X1 U15118 ( .C1(n12839), .C2(n12863), .A(n12838), .B(n12837), .ZN(
        P3_U3216) );
  OAI21_X1 U15119 ( .B1(n12841), .B2(n12843), .A(n12840), .ZN(n12999) );
  INV_X1 U15120 ( .A(n12999), .ZN(n12851) );
  XNOR2_X1 U15121 ( .A(n12842), .B(n12843), .ZN(n12845) );
  AOI222_X1 U15122 ( .A1(n15262), .A2(n12845), .B1(n7302), .B2(n15256), .C1(
        n12844), .C2(n15259), .ZN(n12996) );
  MUX2_X1 U15123 ( .A(n12846), .B(n12996), .S(n15273), .Z(n12850) );
  INV_X1 U15124 ( .A(n12847), .ZN(n12848) );
  AOI22_X1 U15125 ( .A1(n12998), .A2(n12860), .B1(n15226), .B2(n12848), .ZN(
        n12849) );
  OAI211_X1 U15126 ( .C1(n12851), .C2(n12863), .A(n12850), .B(n12849), .ZN(
        P3_U3217) );
  XNOR2_X1 U15127 ( .A(n12852), .B(n12854), .ZN(n13007) );
  INV_X1 U15128 ( .A(n13007), .ZN(n12864) );
  XNOR2_X1 U15129 ( .A(n12853), .B(n12854), .ZN(n12857) );
  AOI222_X1 U15130 ( .A1(n15262), .A2(n12857), .B1(n12856), .B2(n15256), .C1(
        n12855), .C2(n15259), .ZN(n13002) );
  MUX2_X1 U15131 ( .A(n14383), .B(n13002), .S(n15273), .Z(n12862) );
  INV_X1 U15132 ( .A(n12858), .ZN(n12859) );
  AOI22_X1 U15133 ( .A1(n13004), .A2(n12860), .B1(n12859), .B2(n15226), .ZN(
        n12861) );
  OAI211_X1 U15134 ( .C1(n12864), .C2(n12863), .A(n12862), .B(n12861), .ZN(
        P3_U3218) );
  NOR2_X1 U15135 ( .A1(n15329), .A2(n12922), .ZN(n12866) );
  AOI21_X1 U15136 ( .B1(P3_REG1_REG_31__SCAN_IN), .B2(n15329), .A(n12866), 
        .ZN(n12865) );
  OAI21_X1 U15137 ( .B1(n12924), .B2(n12907), .A(n12865), .ZN(P3_U3490) );
  NAND2_X1 U15138 ( .A1(n12925), .A2(n12918), .ZN(n12868) );
  INV_X1 U15139 ( .A(n12866), .ZN(n12867) );
  OAI211_X1 U15140 ( .C1(n15331), .C2(n8677), .A(n12868), .B(n12867), .ZN(
        P3_U3489) );
  INV_X1 U15141 ( .A(n12869), .ZN(n12931) );
  INV_X1 U15142 ( .A(n12929), .ZN(n12870) );
  NAND2_X1 U15143 ( .A1(n12872), .A2(n12918), .ZN(n12873) );
  OAI211_X1 U15144 ( .C1(n12931), .C2(n12903), .A(n12874), .B(n12873), .ZN(
        P3_U3487) );
  AOI21_X1 U15145 ( .B1(n15293), .B2(n12876), .A(n12875), .ZN(n12934) );
  MUX2_X1 U15146 ( .A(n12877), .B(n12934), .S(n15331), .Z(n12878) );
  OAI21_X1 U15147 ( .B1(n12937), .B2(n12907), .A(n12878), .ZN(P3_U3486) );
  AOI21_X1 U15148 ( .B1(n12888), .B2(n12880), .A(n12879), .ZN(n12938) );
  MUX2_X1 U15149 ( .A(n12881), .B(n12938), .S(n15331), .Z(n12882) );
  OAI21_X1 U15150 ( .B1(n12903), .B2(n12941), .A(n12882), .ZN(P3_U3485) );
  MUX2_X1 U15151 ( .A(n12883), .B(n12942), .S(n15331), .Z(n12885) );
  NAND2_X1 U15152 ( .A1(n12944), .A2(n12918), .ZN(n12884) );
  OAI211_X1 U15153 ( .C1(n12903), .C2(n12947), .A(n12885), .B(n12884), .ZN(
        P3_U3484) );
  AOI21_X1 U15154 ( .B1(n12888), .B2(n12887), .A(n12886), .ZN(n12948) );
  MUX2_X1 U15155 ( .A(n12889), .B(n12948), .S(n15331), .Z(n12890) );
  OAI21_X1 U15156 ( .B1(n12951), .B2(n12903), .A(n12890), .ZN(P3_U3483) );
  INV_X1 U15157 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12891) );
  MUX2_X1 U15158 ( .A(n12891), .B(n12952), .S(n15331), .Z(n12893) );
  NAND2_X1 U15159 ( .A1(n12954), .A2(n12918), .ZN(n12892) );
  OAI211_X1 U15160 ( .C1(n12903), .C2(n12957), .A(n12893), .B(n12892), .ZN(
        P3_U3482) );
  MUX2_X1 U15161 ( .A(n12894), .B(n12958), .S(n15331), .Z(n12896) );
  NAND2_X1 U15162 ( .A1(n12960), .A2(n12918), .ZN(n12895) );
  OAI211_X1 U15163 ( .C1(n12963), .C2(n12903), .A(n12896), .B(n12895), .ZN(
        P3_U3481) );
  MUX2_X1 U15164 ( .A(n12897), .B(n12964), .S(n15331), .Z(n12899) );
  NAND2_X1 U15165 ( .A1(n12966), .A2(n12918), .ZN(n12898) );
  OAI211_X1 U15166 ( .C1(n12903), .C2(n12969), .A(n12899), .B(n12898), .ZN(
        P3_U3480) );
  INV_X1 U15167 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12900) );
  MUX2_X1 U15168 ( .A(n12900), .B(n12970), .S(n15331), .Z(n12902) );
  NAND2_X1 U15169 ( .A1(n12972), .A2(n12918), .ZN(n12901) );
  OAI211_X1 U15170 ( .C1(n12903), .C2(n12976), .A(n12902), .B(n12901), .ZN(
        P3_U3479) );
  MUX2_X1 U15171 ( .A(n12904), .B(n12977), .S(n15331), .Z(n12906) );
  NAND2_X1 U15172 ( .A1(n12979), .A2(n12919), .ZN(n12905) );
  OAI211_X1 U15173 ( .C1(n12907), .C2(n12982), .A(n12906), .B(n12905), .ZN(
        P3_U3478) );
  MUX2_X1 U15174 ( .A(n12908), .B(n12984), .S(n15331), .Z(n12910) );
  AOI22_X1 U15175 ( .A1(n12987), .A2(n12919), .B1(n12918), .B2(n12986), .ZN(
        n12909) );
  NAND2_X1 U15176 ( .A1(n12910), .A2(n12909), .ZN(P3_U3477) );
  MUX2_X1 U15177 ( .A(n12911), .B(n12990), .S(n15331), .Z(n12913) );
  AOI22_X1 U15178 ( .A1(n12993), .A2(n12919), .B1(n12918), .B2(n12992), .ZN(
        n12912) );
  NAND2_X1 U15179 ( .A1(n12913), .A2(n12912), .ZN(P3_U3476) );
  MUX2_X1 U15180 ( .A(n12914), .B(n12996), .S(n15331), .Z(n12916) );
  AOI22_X1 U15181 ( .A1(n12999), .A2(n12919), .B1(n12918), .B2(n12998), .ZN(
        n12915) );
  NAND2_X1 U15182 ( .A1(n12916), .A2(n12915), .ZN(P3_U3475) );
  MUX2_X1 U15183 ( .A(n12917), .B(n13002), .S(n15331), .Z(n12921) );
  AOI22_X1 U15184 ( .A1(n13007), .A2(n12919), .B1(n12918), .B2(n13004), .ZN(
        n12920) );
  NAND2_X1 U15185 ( .A1(n12921), .A2(n12920), .ZN(P3_U3474) );
  NOR2_X1 U15186 ( .A1(n15316), .A2(n12922), .ZN(n12926) );
  AOI21_X1 U15187 ( .B1(P3_REG0_REG_31__SCAN_IN), .B2(n15316), .A(n12926), 
        .ZN(n12923) );
  OAI21_X1 U15188 ( .B1(n12924), .B2(n12983), .A(n12923), .ZN(P3_U3458) );
  NAND2_X1 U15189 ( .A1(n12925), .A2(n13005), .ZN(n12928) );
  INV_X1 U15190 ( .A(n12926), .ZN(n12927) );
  OAI211_X1 U15191 ( .C1(n8678), .C2(n15318), .A(n12928), .B(n12927), .ZN(
        P3_U3457) );
  MUX2_X1 U15192 ( .A(n12929), .B(P3_REG0_REG_28__SCAN_IN), .S(n15316), .Z(
        n12933) );
  OAI22_X1 U15193 ( .A1(n12931), .A2(n12975), .B1(n12930), .B2(n12983), .ZN(
        n12932) );
  OR2_X1 U15194 ( .A1(n12933), .A2(n12932), .ZN(P3_U3455) );
  MUX2_X1 U15195 ( .A(n12935), .B(n12934), .S(n15318), .Z(n12936) );
  OAI21_X1 U15196 ( .B1(n12937), .B2(n12983), .A(n12936), .ZN(P3_U3454) );
  MUX2_X1 U15197 ( .A(n12939), .B(n12938), .S(n15318), .Z(n12940) );
  OAI21_X1 U15198 ( .B1(n12941), .B2(n12975), .A(n12940), .ZN(P3_U3453) );
  MUX2_X1 U15199 ( .A(n12943), .B(n12942), .S(n15318), .Z(n12946) );
  NAND2_X1 U15200 ( .A1(n12944), .A2(n13005), .ZN(n12945) );
  OAI211_X1 U15201 ( .C1(n12947), .C2(n12975), .A(n12946), .B(n12945), .ZN(
        P3_U3452) );
  MUX2_X1 U15202 ( .A(n12949), .B(n12948), .S(n15318), .Z(n12950) );
  OAI21_X1 U15203 ( .B1(n12951), .B2(n12975), .A(n12950), .ZN(P3_U3451) );
  MUX2_X1 U15204 ( .A(n12953), .B(n12952), .S(n15318), .Z(n12956) );
  NAND2_X1 U15205 ( .A1(n12954), .A2(n13005), .ZN(n12955) );
  OAI211_X1 U15206 ( .C1(n12957), .C2(n12975), .A(n12956), .B(n12955), .ZN(
        P3_U3450) );
  MUX2_X1 U15207 ( .A(n12959), .B(n12958), .S(n15318), .Z(n12962) );
  NAND2_X1 U15208 ( .A1(n12960), .A2(n13005), .ZN(n12961) );
  OAI211_X1 U15209 ( .C1(n12963), .C2(n12975), .A(n12962), .B(n12961), .ZN(
        P3_U3449) );
  MUX2_X1 U15210 ( .A(n12965), .B(n12964), .S(n15318), .Z(n12968) );
  NAND2_X1 U15211 ( .A1(n12966), .A2(n13005), .ZN(n12967) );
  OAI211_X1 U15212 ( .C1(n12969), .C2(n12975), .A(n12968), .B(n12967), .ZN(
        P3_U3448) );
  INV_X1 U15213 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12971) );
  MUX2_X1 U15214 ( .A(n12971), .B(n12970), .S(n15318), .Z(n12974) );
  NAND2_X1 U15215 ( .A1(n12972), .A2(n13005), .ZN(n12973) );
  OAI211_X1 U15216 ( .C1(n12976), .C2(n12975), .A(n12974), .B(n12973), .ZN(
        P3_U3447) );
  MUX2_X1 U15217 ( .A(n12978), .B(n12977), .S(n15318), .Z(n12981) );
  NAND2_X1 U15218 ( .A1(n12979), .A2(n13006), .ZN(n12980) );
  OAI211_X1 U15219 ( .C1(n12983), .C2(n12982), .A(n12981), .B(n12980), .ZN(
        P3_U3446) );
  MUX2_X1 U15220 ( .A(n12985), .B(n12984), .S(n15318), .Z(n12989) );
  AOI22_X1 U15221 ( .A1(n12987), .A2(n13006), .B1(n13005), .B2(n12986), .ZN(
        n12988) );
  NAND2_X1 U15222 ( .A1(n12989), .A2(n12988), .ZN(P3_U3444) );
  INV_X1 U15223 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12991) );
  MUX2_X1 U15224 ( .A(n12991), .B(n12990), .S(n15318), .Z(n12995) );
  AOI22_X1 U15225 ( .A1(n12993), .A2(n13006), .B1(n13005), .B2(n12992), .ZN(
        n12994) );
  NAND2_X1 U15226 ( .A1(n12995), .A2(n12994), .ZN(P3_U3441) );
  INV_X1 U15227 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12997) );
  MUX2_X1 U15228 ( .A(n12997), .B(n12996), .S(n15318), .Z(n13001) );
  AOI22_X1 U15229 ( .A1(n12999), .A2(n13006), .B1(n13005), .B2(n12998), .ZN(
        n13000) );
  NAND2_X1 U15230 ( .A1(n13001), .A2(n13000), .ZN(P3_U3438) );
  MUX2_X1 U15231 ( .A(n13003), .B(n13002), .S(n15318), .Z(n13009) );
  AOI22_X1 U15232 ( .A1(n13007), .A2(n13006), .B1(n13005), .B2(n13004), .ZN(
        n13008) );
  NAND2_X1 U15233 ( .A1(n13009), .A2(n13008), .ZN(P3_U3435) );
  INV_X1 U15234 ( .A(n13010), .ZN(n13016) );
  NOR4_X1 U15235 ( .A1(n13012), .A2(P3_IR_REG_30__SCAN_IN), .A3(P3_U3151), 
        .A4(n13011), .ZN(n13013) );
  AOI21_X1 U15236 ( .B1(SI_31_), .B2(n13014), .A(n13013), .ZN(n13015) );
  OAI21_X1 U15237 ( .B1(n13016), .B2(n13021), .A(n13015), .ZN(P3_U3264) );
  INV_X1 U15238 ( .A(n13017), .ZN(n13020) );
  OAI222_X1 U15239 ( .A1(n13023), .A2(n13022), .B1(n13021), .B2(n13020), .C1(
        P3_U3151), .C2(n13018), .ZN(P3_U3266) );
  MUX2_X1 U15240 ( .A(n13024), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  XNOR2_X1 U15241 ( .A(n13404), .B(n6469), .ZN(n13035) );
  NAND2_X1 U15242 ( .A1(n13189), .A2(n13490), .ZN(n13036) );
  XNOR2_X1 U15243 ( .A(n13590), .B(n13044), .ZN(n13034) );
  NAND2_X1 U15244 ( .A1(n13190), .A2(n13490), .ZN(n13033) );
  XNOR2_X1 U15245 ( .A(n13596), .B(n13044), .ZN(n13142) );
  NAND2_X1 U15246 ( .A1(n13191), .A2(n13490), .ZN(n13032) );
  INV_X1 U15247 ( .A(n13025), .ZN(n13028) );
  XNOR2_X1 U15248 ( .A(n13601), .B(n6469), .ZN(n13083) );
  AND2_X1 U15249 ( .A1(n13192), .A2(n13490), .ZN(n13029) );
  NAND2_X1 U15250 ( .A1(n13083), .A2(n13029), .ZN(n13030) );
  OAI21_X1 U15251 ( .B1(n13083), .B2(n13029), .A(n13030), .ZN(n13162) );
  INV_X1 U15252 ( .A(n13030), .ZN(n13031) );
  XNOR2_X1 U15253 ( .A(n13142), .B(n13032), .ZN(n13086) );
  XNOR2_X1 U15254 ( .A(n13034), .B(n13033), .ZN(n13144) );
  XNOR2_X1 U15255 ( .A(n13035), .B(n13036), .ZN(n13105) );
  NAND2_X1 U15256 ( .A1(n13106), .A2(n13105), .ZN(n13104) );
  AND2_X1 U15257 ( .A1(n13188), .A2(n13490), .ZN(n13037) );
  INV_X1 U15258 ( .A(n13038), .ZN(n13039) );
  NAND2_X2 U15259 ( .A1(n13150), .A2(n13040), .ZN(n13042) );
  XNOR2_X2 U15260 ( .A(n13042), .B(n7487), .ZN(n13071) );
  INV_X1 U15261 ( .A(n13042), .ZN(n13043) );
  XNOR2_X1 U15262 ( .A(n13567), .B(n13044), .ZN(n13113) );
  NAND2_X1 U15263 ( .A1(n13186), .A2(n13490), .ZN(n13045) );
  NOR2_X1 U15264 ( .A1(n13113), .A2(n13045), .ZN(n13046) );
  AOI21_X1 U15265 ( .B1(n13113), .B2(n13045), .A(n13046), .ZN(n13125) );
  INV_X1 U15266 ( .A(n13046), .ZN(n13047) );
  XNOR2_X1 U15267 ( .A(n13562), .B(n6469), .ZN(n13168) );
  AND2_X1 U15268 ( .A1(n13185), .A2(n13490), .ZN(n13048) );
  NAND2_X1 U15269 ( .A1(n13168), .A2(n13048), .ZN(n13053) );
  INV_X1 U15270 ( .A(n13168), .ZN(n13050) );
  INV_X1 U15271 ( .A(n13048), .ZN(n13049) );
  NAND2_X1 U15272 ( .A1(n13050), .A2(n13049), .ZN(n13051) );
  NAND2_X1 U15273 ( .A1(n13184), .A2(n13490), .ZN(n13056) );
  XNOR2_X1 U15274 ( .A(n13557), .B(n6469), .ZN(n13058) );
  XOR2_X1 U15275 ( .A(n13056), .B(n13058), .Z(n13170) );
  INV_X1 U15276 ( .A(n13053), .ZN(n13054) );
  NOR2_X1 U15277 ( .A1(n13170), .A2(n13054), .ZN(n13055) );
  INV_X1 U15278 ( .A(n13056), .ZN(n13057) );
  XNOR2_X1 U15279 ( .A(n13317), .B(n6469), .ZN(n13061) );
  AND2_X1 U15280 ( .A1(n13183), .A2(n13490), .ZN(n13060) );
  NAND2_X1 U15281 ( .A1(n13061), .A2(n13060), .ZN(n13090) );
  OAI21_X1 U15282 ( .B1(n13061), .B2(n13060), .A(n13090), .ZN(n13063) );
  AOI21_X1 U15283 ( .B1(n13062), .B2(n13063), .A(n14824), .ZN(n13064) );
  NAND2_X1 U15284 ( .A1(n13064), .A2(n13091), .ZN(n13070) );
  AND2_X1 U15285 ( .A1(n13184), .A2(n13172), .ZN(n13065) );
  AOI21_X1 U15286 ( .B1(n13182), .B2(n13173), .A(n13065), .ZN(n13314) );
  INV_X1 U15287 ( .A(n13314), .ZN(n13068) );
  OAI22_X1 U15288 ( .A1(n13318), .A2(n14832), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13066), .ZN(n13067) );
  AOI21_X1 U15289 ( .B1(n13068), .B2(n13159), .A(n13067), .ZN(n13069) );
  OAI211_X1 U15290 ( .C1(n13647), .C2(n13133), .A(n13070), .B(n13069), .ZN(
        P2_U3186) );
  AOI22_X1 U15291 ( .A1(n13071), .A2(n13148), .B1(n13167), .B2(n13187), .ZN(
        n13079) );
  INV_X1 U15292 ( .A(n13072), .ZN(n13078) );
  AND2_X1 U15293 ( .A1(n13188), .A2(n13172), .ZN(n13073) );
  AOI21_X1 U15294 ( .B1(n13186), .B2(n13173), .A(n13073), .ZN(n13573) );
  INV_X1 U15295 ( .A(n13074), .ZN(n13370) );
  AOI22_X1 U15296 ( .A1(n13370), .A2(n13174), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13075) );
  OAI21_X1 U15297 ( .B1(n13573), .B2(n14822), .A(n13075), .ZN(n13076) );
  AOI21_X1 U15298 ( .B1(n13375), .B2(n14829), .A(n13076), .ZN(n13077) );
  OAI21_X1 U15299 ( .B1(n13079), .B2(n13078), .A(n13077), .ZN(P2_U3188) );
  NOR2_X1 U15300 ( .A1(n14832), .A2(n13431), .ZN(n13082) );
  AOI22_X1 U15301 ( .A1(n13190), .A2(n13173), .B1(n13172), .B2(n13192), .ZN(
        n13427) );
  OAI22_X1 U15302 ( .A1(n14822), .A2(n13427), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13080), .ZN(n13081) );
  AOI211_X1 U15303 ( .C1(n13596), .C2(n14829), .A(n13082), .B(n13081), .ZN(
        n13089) );
  INV_X1 U15304 ( .A(n13161), .ZN(n13085) );
  NAND3_X1 U15305 ( .A1(n13083), .A2(n13167), .A3(n13192), .ZN(n13084) );
  OAI21_X1 U15306 ( .B1(n13085), .B2(n14824), .A(n13084), .ZN(n13087) );
  NAND2_X1 U15307 ( .A1(n13087), .A2(n13086), .ZN(n13088) );
  OAI211_X1 U15308 ( .C1(n7237), .C2(n14824), .A(n13089), .B(n13088), .ZN(
        P2_U3191) );
  NAND2_X1 U15309 ( .A1(n13091), .A2(n13090), .ZN(n13096) );
  NAND2_X1 U15310 ( .A1(n13182), .A2(n13490), .ZN(n13093) );
  XNOR2_X1 U15311 ( .A(n13093), .B(n6469), .ZN(n13094) );
  XNOR2_X1 U15312 ( .A(n13548), .B(n13094), .ZN(n13095) );
  XNOR2_X1 U15313 ( .A(n13096), .B(n13095), .ZN(n13103) );
  NAND2_X1 U15314 ( .A1(n13181), .A2(n13173), .ZN(n13098) );
  NAND2_X1 U15315 ( .A1(n13183), .A2(n13172), .ZN(n13097) );
  NAND2_X1 U15316 ( .A1(n13098), .A2(n13097), .ZN(n13303) );
  OAI22_X1 U15317 ( .A1(n13297), .A2(n14832), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13099), .ZN(n13101) );
  NOR2_X1 U15318 ( .A1(n6912), .A2(n13133), .ZN(n13100) );
  AOI211_X1 U15319 ( .C1(n13159), .C2(n13303), .A(n13101), .B(n13100), .ZN(
        n13102) );
  OAI21_X1 U15320 ( .B1(n13103), .B2(n14824), .A(n13102), .ZN(P2_U3192) );
  OAI211_X1 U15321 ( .C1(n13106), .C2(n13105), .A(n13104), .B(n13148), .ZN(
        n13110) );
  AOI22_X1 U15322 ( .A1(n13188), .A2(n13173), .B1(n13172), .B2(n13190), .ZN(
        n13397) );
  OAI22_X1 U15323 ( .A1(n13397), .A2(n14822), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13107), .ZN(n13108) );
  AOI21_X1 U15324 ( .B1(n13405), .B2(n13174), .A(n13108), .ZN(n13109) );
  OAI211_X1 U15325 ( .C1(n9542), .C2(n13133), .A(n13110), .B(n13109), .ZN(
        P2_U3195) );
  INV_X1 U15326 ( .A(n13111), .ZN(n13112) );
  AOI21_X1 U15327 ( .B1(n13124), .B2(n13112), .A(n14824), .ZN(n13116) );
  NOR3_X1 U15328 ( .A1(n13113), .A2(n13117), .A3(n13140), .ZN(n13115) );
  OAI21_X1 U15329 ( .B1(n13116), .B2(n13115), .A(n13114), .ZN(n13123) );
  OAI22_X1 U15330 ( .A1(n13118), .A2(n13136), .B1(n13117), .B2(n13135), .ZN(
        n13341) );
  INV_X1 U15331 ( .A(n13347), .ZN(n13120) );
  OAI22_X1 U15332 ( .A1(n13120), .A2(n14832), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13119), .ZN(n13121) );
  AOI21_X1 U15333 ( .B1(n13341), .B2(n13159), .A(n13121), .ZN(n13122) );
  OAI211_X1 U15334 ( .C1(n7215), .C2(n13133), .A(n13123), .B(n13122), .ZN(
        P2_U3197) );
  OAI211_X1 U15335 ( .C1(n13126), .C2(n13125), .A(n13124), .B(n13148), .ZN(
        n13132) );
  OAI22_X1 U15336 ( .A1(n13128), .A2(n13136), .B1(n13127), .B2(n13135), .ZN(
        n13353) );
  OAI22_X1 U15337 ( .A1(n13361), .A2(n14832), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13129), .ZN(n13130) );
  AOI21_X1 U15338 ( .B1(n13353), .B2(n13159), .A(n13130), .ZN(n13131) );
  OAI211_X1 U15339 ( .C1(n13359), .C2(n13133), .A(n13132), .B(n13131), .ZN(
        P2_U3201) );
  INV_X1 U15340 ( .A(n13134), .ZN(n13147) );
  OAI22_X1 U15341 ( .A1(n13137), .A2(n13136), .B1(n13141), .B2(n13135), .ZN(
        n13412) );
  AOI22_X1 U15342 ( .A1(n13412), .A2(n13159), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13138) );
  OAI21_X1 U15343 ( .B1(n13415), .B2(n14832), .A(n13138), .ZN(n13139) );
  AOI21_X1 U15344 ( .B1(n13590), .B2(n14829), .A(n13139), .ZN(n13146) );
  OAI22_X1 U15345 ( .A1(n13142), .A2(n14824), .B1(n13141), .B2(n13140), .ZN(
        n13143) );
  NAND3_X1 U15346 ( .A1(n7237), .A2(n13144), .A3(n13143), .ZN(n13145) );
  OAI211_X1 U15347 ( .C1(n13147), .C2(n14824), .A(n13146), .B(n13145), .ZN(
        P2_U3205) );
  AOI22_X1 U15348 ( .A1(n13149), .A2(n13148), .B1(n13167), .B2(n13188), .ZN(
        n13156) );
  INV_X1 U15349 ( .A(n13150), .ZN(n13155) );
  AOI22_X1 U15350 ( .A1(n13187), .A2(n13173), .B1(n13172), .B2(n13189), .ZN(
        n13381) );
  INV_X1 U15351 ( .A(n13151), .ZN(n13389) );
  AOI22_X1 U15352 ( .A1(n13174), .A2(n13389), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13152) );
  OAI21_X1 U15353 ( .B1(n13381), .B2(n14822), .A(n13152), .ZN(n13153) );
  AOI21_X1 U15354 ( .B1(n13580), .B2(n14829), .A(n13153), .ZN(n13154) );
  OAI21_X1 U15355 ( .B1(n13156), .B2(n13155), .A(n13154), .ZN(P2_U3207) );
  NAND2_X1 U15356 ( .A1(n13191), .A2(n13173), .ZN(n13158) );
  NAND2_X1 U15357 ( .A1(n13172), .A2(n13193), .ZN(n13157) );
  NAND2_X1 U15358 ( .A1(n13158), .A2(n13157), .ZN(n13439) );
  NAND2_X1 U15359 ( .A1(n13159), .A2(n13439), .ZN(n13160) );
  NAND2_X1 U15360 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13253)
         );
  OAI211_X1 U15361 ( .C1(n14832), .C2(n13442), .A(n13160), .B(n13253), .ZN(
        n13165) );
  AOI211_X1 U15362 ( .C1(n13163), .C2(n13162), .A(n14824), .B(n13161), .ZN(
        n13164) );
  AOI211_X1 U15363 ( .C1(n13601), .C2(n14829), .A(n13165), .B(n13164), .ZN(
        n13166) );
  INV_X1 U15364 ( .A(n13166), .ZN(P2_U3210) );
  NAND3_X1 U15365 ( .A1(n13168), .A2(n13167), .A3(n13185), .ZN(n13169) );
  OAI21_X1 U15366 ( .B1(n13114), .B2(n14824), .A(n13169), .ZN(n13171) );
  NAND2_X1 U15367 ( .A1(n13171), .A2(n13170), .ZN(n13178) );
  AOI22_X1 U15368 ( .A1(n13183), .A2(n13173), .B1(n13172), .B2(n13185), .ZN(
        n13326) );
  AOI22_X1 U15369 ( .A1(n13331), .A2(n13174), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13175) );
  OAI21_X1 U15370 ( .B1(n13326), .B2(n14822), .A(n13175), .ZN(n13176) );
  AOI21_X1 U15371 ( .B1(n13557), .B2(n14829), .A(n13176), .ZN(n13177) );
  OAI211_X1 U15372 ( .C1(n14824), .C2(n13179), .A(n13178), .B(n13177), .ZN(
        P2_U3212) );
  MUX2_X1 U15373 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13283), .S(n13208), .Z(
        P2_U3562) );
  MUX2_X1 U15374 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13180), .S(n13208), .Z(
        P2_U3561) );
  MUX2_X1 U15375 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13181), .S(n13208), .Z(
        P2_U3560) );
  MUX2_X1 U15376 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13182), .S(P2_U3947), .Z(
        P2_U3559) );
  MUX2_X1 U15377 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13183), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U15378 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13184), .S(P2_U3947), .Z(
        P2_U3557) );
  MUX2_X1 U15379 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13185), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U15380 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13186), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U15381 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13187), .S(n13208), .Z(
        P2_U3554) );
  MUX2_X1 U15382 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13188), .S(n13208), .Z(
        P2_U3553) );
  MUX2_X1 U15383 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13189), .S(n13208), .Z(
        P2_U3552) );
  MUX2_X1 U15384 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13190), .S(n13208), .Z(
        P2_U3551) );
  MUX2_X1 U15385 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13191), .S(n13208), .Z(
        P2_U3550) );
  MUX2_X1 U15386 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13192), .S(n13208), .Z(
        P2_U3549) );
  MUX2_X1 U15387 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13193), .S(n13208), .Z(
        P2_U3548) );
  MUX2_X1 U15388 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13194), .S(n13208), .Z(
        P2_U3547) );
  MUX2_X1 U15389 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13195), .S(n13208), .Z(
        P2_U3546) );
  MUX2_X1 U15390 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13196), .S(n13208), .Z(
        P2_U3545) );
  MUX2_X1 U15391 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13197), .S(n13208), .Z(
        P2_U3543) );
  MUX2_X1 U15392 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13198), .S(n13208), .Z(
        P2_U3542) );
  MUX2_X1 U15393 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13199), .S(n13208), .Z(
        P2_U3541) );
  MUX2_X1 U15394 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13200), .S(n13208), .Z(
        P2_U3540) );
  MUX2_X1 U15395 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13201), .S(n13208), .Z(
        P2_U3539) );
  MUX2_X1 U15396 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13202), .S(n13208), .Z(
        P2_U3538) );
  MUX2_X1 U15397 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13203), .S(n13208), .Z(
        P2_U3537) );
  MUX2_X1 U15398 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13204), .S(n13208), .Z(
        P2_U3536) );
  MUX2_X1 U15399 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13205), .S(n13208), .Z(
        P2_U3535) );
  MUX2_X1 U15400 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13206), .S(n13208), .Z(
        P2_U3534) );
  MUX2_X1 U15401 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13207), .S(n13208), .Z(
        P2_U3533) );
  MUX2_X1 U15402 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n9552), .S(n13208), .Z(
        P2_U3532) );
  MUX2_X1 U15403 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n9559), .S(n13208), .Z(
        P2_U3531) );
  INV_X1 U15404 ( .A(n14930), .ZN(n14939) );
  AND3_X1 U15405 ( .A1(n14855), .A2(n13210), .A3(n13209), .ZN(n13211) );
  NOR3_X1 U15406 ( .A1(n14913), .A2(n13212), .A3(n13211), .ZN(n13213) );
  AOI21_X1 U15407 ( .B1(n14939), .B2(n13214), .A(n13213), .ZN(n13221) );
  NOR2_X1 U15408 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9148), .ZN(n13215) );
  AOI21_X1 U15409 ( .B1(n14924), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n13215), .ZN(
        n13220) );
  OAI211_X1 U15410 ( .C1(n13218), .C2(n13217), .A(n14863), .B(n13216), .ZN(
        n13219) );
  NAND3_X1 U15411 ( .A1(n13221), .A2(n13220), .A3(n13219), .ZN(P2_U3217) );
  NAND2_X1 U15412 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n14938), .ZN(n13231) );
  MUX2_X1 U15413 ( .A(n9317), .B(P2_REG2_REG_16__SCAN_IN), .S(n14938), .Z(
        n13222) );
  INV_X1 U15414 ( .A(n13222), .ZN(n14942) );
  NAND2_X1 U15415 ( .A1(n13238), .A2(n13223), .ZN(n13227) );
  NAND2_X1 U15416 ( .A1(n13227), .A2(n13226), .ZN(n13229) );
  NAND2_X1 U15417 ( .A1(n13228), .A2(n13229), .ZN(n13230) );
  XNOR2_X1 U15418 ( .A(n14929), .B(n13229), .ZN(n14926) );
  NAND2_X1 U15419 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n14926), .ZN(n14925) );
  NAND2_X1 U15420 ( .A1(n13230), .A2(n14925), .ZN(n14943) );
  NAND2_X1 U15421 ( .A1(n14942), .A2(n14943), .ZN(n14940) );
  NAND2_X1 U15422 ( .A1(n13231), .A2(n14940), .ZN(n13235) );
  INV_X1 U15423 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13251) );
  NAND2_X1 U15424 ( .A1(n13255), .A2(n13251), .ZN(n13232) );
  OAI21_X1 U15425 ( .B1(n13255), .B2(n13251), .A(n13232), .ZN(n13234) );
  NAND2_X1 U15426 ( .A1(n13250), .A2(n13251), .ZN(n13233) );
  OAI211_X1 U15427 ( .C1(n13251), .C2(n13250), .A(n13235), .B(n13233), .ZN(
        n13249) );
  OAI211_X1 U15428 ( .C1(n13235), .C2(n13234), .A(n13249), .B(n14941), .ZN(
        n13248) );
  AND2_X1 U15429 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13236) );
  AOI21_X1 U15430 ( .B1(n14924), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n13236), 
        .ZN(n13247) );
  NAND2_X1 U15431 ( .A1(n14939), .A2(n13255), .ZN(n13246) );
  XNOR2_X1 U15432 ( .A(n13255), .B(n13609), .ZN(n13244) );
  NAND2_X1 U15433 ( .A1(n14938), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n13242) );
  NOR2_X1 U15434 ( .A1(n13239), .A2(n14929), .ZN(n13240) );
  XNOR2_X1 U15435 ( .A(n13239), .B(n14929), .ZN(n14921) );
  NOR2_X1 U15436 ( .A1(n14920), .A2(n14921), .ZN(n14919) );
  NOR2_X1 U15437 ( .A1(n13240), .A2(n14919), .ZN(n14935) );
  XNOR2_X1 U15438 ( .A(n14938), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n14934) );
  NOR2_X1 U15439 ( .A1(n14935), .A2(n14934), .ZN(n14933) );
  INV_X1 U15440 ( .A(n14933), .ZN(n13241) );
  NAND2_X1 U15441 ( .A1(n13242), .A2(n13241), .ZN(n13243) );
  NAND2_X1 U15442 ( .A1(n13243), .A2(n13244), .ZN(n13257) );
  OAI211_X1 U15443 ( .C1(n13244), .C2(n13243), .A(n14863), .B(n13257), .ZN(
        n13245) );
  NAND4_X1 U15444 ( .A1(n13248), .A2(n13247), .A3(n13246), .A4(n13245), .ZN(
        P2_U3231) );
  OAI21_X1 U15445 ( .B1(n13251), .B2(n13250), .A(n13249), .ZN(n13264) );
  XNOR2_X1 U15446 ( .A(n13264), .B(n13265), .ZN(n13252) );
  NOR2_X1 U15447 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n13252), .ZN(n13267) );
  AOI21_X1 U15448 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n13252), .A(n13267), 
        .ZN(n13263) );
  INV_X1 U15449 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n13254) );
  OAI21_X1 U15450 ( .B1(n14946), .B2(n13254), .A(n13253), .ZN(n13261) );
  NAND2_X1 U15451 ( .A1(n13255), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n13256) );
  XNOR2_X1 U15452 ( .A(n13270), .B(n13269), .ZN(n13259) );
  INV_X1 U15453 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n13258) );
  NOR2_X1 U15454 ( .A1(n13258), .A2(n13259), .ZN(n13272) );
  AOI211_X1 U15455 ( .C1(n13259), .C2(n13258), .A(n13272), .B(n14932), .ZN(
        n13260) );
  AOI211_X1 U15456 ( .C1(n14939), .C2(n13265), .A(n13261), .B(n13260), .ZN(
        n13262) );
  OAI21_X1 U15457 ( .B1(n13263), .B2(n14913), .A(n13262), .ZN(P2_U3232) );
  NOR2_X1 U15458 ( .A1(n13265), .A2(n13264), .ZN(n13266) );
  NOR2_X1 U15459 ( .A1(n13267), .A2(n13266), .ZN(n13268) );
  XOR2_X1 U15460 ( .A(n13268), .B(P2_REG2_REG_19__SCAN_IN), .Z(n13275) );
  NOR2_X1 U15461 ( .A1(n13270), .A2(n13269), .ZN(n13271) );
  NOR2_X1 U15462 ( .A1(n13272), .A2(n13271), .ZN(n13273) );
  XNOR2_X1 U15463 ( .A(n13273), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n13274) );
  AOI22_X1 U15464 ( .A1(n13275), .A2(n14941), .B1(n14863), .B2(n13274), .ZN(
        n13277) );
  MUX2_X1 U15465 ( .A(n13278), .B(n13277), .S(n13276), .Z(n13280) );
  NAND2_X1 U15466 ( .A1(n14924), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n13279) );
  OAI211_X1 U15467 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n13080), .A(n13280), .B(
        n13279), .ZN(P2_U3233) );
  NAND2_X1 U15468 ( .A1(n13284), .A2(n13283), .ZN(n13537) );
  NOR2_X1 U15469 ( .A1(n13517), .A2(n13537), .ZN(n13290) );
  AOI21_X1 U15470 ( .B1(n13517), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13290), 
        .ZN(n13286) );
  NAND2_X1 U15471 ( .A1(n9821), .A2(n13525), .ZN(n13285) );
  OAI211_X1 U15472 ( .C1(n13535), .C2(n13498), .A(n13286), .B(n13285), .ZN(
        P2_U3234) );
  OAI211_X1 U15473 ( .C1(n13641), .C2(n13288), .A(n11269), .B(n13287), .ZN(
        n13538) );
  NOR2_X1 U15474 ( .A1(n13641), .A2(n13461), .ZN(n13289) );
  AOI211_X1 U15475 ( .C1(n13517), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13290), 
        .B(n13289), .ZN(n13291) );
  OAI21_X1 U15476 ( .B1(n13498), .B2(n13538), .A(n13291), .ZN(P2_U3235) );
  XNOR2_X1 U15477 ( .A(n13293), .B(n13292), .ZN(n13549) );
  INV_X1 U15478 ( .A(n13294), .ZN(n13295) );
  AOI211_X1 U15479 ( .C1(n13548), .C2(n13316), .A(n13490), .B(n13295), .ZN(
        n13547) );
  NOR2_X1 U15480 ( .A1(n6912), .A2(n13461), .ZN(n13299) );
  OAI22_X1 U15481 ( .A1(n13297), .A2(n13521), .B1(n13296), .B2(n13519), .ZN(
        n13298) );
  AOI211_X1 U15482 ( .C1(n13547), .C2(n13529), .A(n13299), .B(n13298), .ZN(
        n13307) );
  AOI21_X1 U15483 ( .B1(n13310), .B2(n13301), .A(n13300), .ZN(n13305) );
  INV_X1 U15484 ( .A(n13303), .ZN(n13304) );
  NAND2_X1 U15485 ( .A1(n13546), .A2(n13519), .ZN(n13306) );
  OAI211_X1 U15486 ( .C1(n13549), .C2(n13467), .A(n13307), .B(n13306), .ZN(
        P2_U3237) );
  XNOR2_X1 U15487 ( .A(n13309), .B(n13308), .ZN(n13552) );
  INV_X1 U15488 ( .A(n13552), .ZN(n13324) );
  OAI21_X1 U15489 ( .B1(n13312), .B2(n13311), .A(n13310), .ZN(n13313) );
  NAND2_X1 U15490 ( .A1(n13313), .A2(n13484), .ZN(n13315) );
  NAND2_X1 U15491 ( .A1(n13315), .A2(n13314), .ZN(n13550) );
  AOI211_X1 U15492 ( .C1(n13317), .C2(n13329), .A(n13490), .B(n6913), .ZN(
        n13551) );
  NAND2_X1 U15493 ( .A1(n13551), .A2(n13529), .ZN(n13321) );
  INV_X1 U15494 ( .A(n13318), .ZN(n13319) );
  AOI22_X1 U15495 ( .A1(n13319), .A2(n13511), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n13517), .ZN(n13320) );
  OAI211_X1 U15496 ( .C1(n13647), .C2(n13461), .A(n13321), .B(n13320), .ZN(
        n13322) );
  AOI21_X1 U15497 ( .B1(n13550), .B2(n13519), .A(n13322), .ZN(n13323) );
  OAI21_X1 U15498 ( .B1(n13324), .B2(n13467), .A(n13323), .ZN(P2_U3238) );
  XOR2_X1 U15499 ( .A(n13335), .B(n13325), .Z(n13327) );
  OAI21_X1 U15500 ( .B1(n13327), .B2(n13504), .A(n13326), .ZN(n13555) );
  INV_X1 U15501 ( .A(n13328), .ZN(n13345) );
  AOI21_X1 U15502 ( .B1(n13345), .B2(n13557), .A(n13490), .ZN(n13330) );
  NAND2_X1 U15503 ( .A1(n13556), .A2(n13529), .ZN(n13333) );
  AOI22_X1 U15504 ( .A1(n13331), .A2(n13511), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n13517), .ZN(n13332) );
  OAI211_X1 U15505 ( .C1(n13334), .C2(n13461), .A(n13333), .B(n13332), .ZN(
        n13338) );
  XNOR2_X1 U15506 ( .A(n13336), .B(n13335), .ZN(n13559) );
  NOR2_X1 U15507 ( .A1(n13559), .A2(n13467), .ZN(n13337) );
  AOI211_X1 U15508 ( .C1(n13519), .C2(n13555), .A(n13338), .B(n13337), .ZN(
        n13339) );
  INV_X1 U15509 ( .A(n13339), .ZN(P2_U3239) );
  XNOR2_X1 U15510 ( .A(n13340), .B(n7216), .ZN(n13342) );
  AOI21_X1 U15511 ( .B1(n13342), .B2(n13484), .A(n13341), .ZN(n13564) );
  OAI21_X1 U15512 ( .B1(n6593), .B2(n13344), .A(n13343), .ZN(n13560) );
  AOI21_X1 U15513 ( .B1(n13358), .B2(n13562), .A(n13490), .ZN(n13346) );
  AND2_X1 U15514 ( .A1(n13346), .A2(n13345), .ZN(n13561) );
  NAND2_X1 U15515 ( .A1(n13561), .A2(n13529), .ZN(n13349) );
  AOI22_X1 U15516 ( .A1(n13347), .A2(n13511), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n13517), .ZN(n13348) );
  OAI211_X1 U15517 ( .C1(n7215), .C2(n13461), .A(n13349), .B(n13348), .ZN(
        n13350) );
  AOI21_X1 U15518 ( .B1(n13560), .B2(n13527), .A(n13350), .ZN(n13351) );
  OAI21_X1 U15519 ( .B1(n13517), .B2(n13564), .A(n13351), .ZN(P2_U3240) );
  XNOR2_X1 U15520 ( .A(n13352), .B(n13357), .ZN(n13354) );
  AOI21_X1 U15521 ( .B1(n13354), .B2(n13484), .A(n13353), .ZN(n13570) );
  AOI21_X1 U15522 ( .B1(n13357), .B2(n13356), .A(n13355), .ZN(n13566) );
  OAI211_X1 U15523 ( .C1(n6579), .C2(n13359), .A(n11269), .B(n13358), .ZN(
        n13569) );
  INV_X1 U15524 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13360) );
  OAI22_X1 U15525 ( .A1(n13361), .A2(n13521), .B1(n13360), .B2(n13519), .ZN(
        n13362) );
  AOI21_X1 U15526 ( .B1(n13567), .B2(n13525), .A(n13362), .ZN(n13363) );
  OAI21_X1 U15527 ( .B1(n13569), .B2(n13498), .A(n13363), .ZN(n13364) );
  AOI21_X1 U15528 ( .B1(n13566), .B2(n13527), .A(n13364), .ZN(n13365) );
  OAI21_X1 U15529 ( .B1(n13517), .B2(n13570), .A(n13365), .ZN(P2_U3241) );
  INV_X1 U15530 ( .A(n13573), .ZN(n13369) );
  XOR2_X1 U15531 ( .A(n13371), .B(n13366), .Z(n13367) );
  NAND2_X1 U15532 ( .A1(n13367), .A2(n13484), .ZN(n13574) );
  INV_X1 U15533 ( .A(n13574), .ZN(n13368) );
  AOI211_X1 U15534 ( .C1(n13511), .C2(n13370), .A(n13369), .B(n13368), .ZN(
        n13379) );
  XNOR2_X1 U15535 ( .A(n13372), .B(n13371), .ZN(n13576) );
  NAND2_X1 U15536 ( .A1(n13375), .A2(n13387), .ZN(n13373) );
  NAND2_X1 U15537 ( .A1(n13373), .A2(n11269), .ZN(n13374) );
  OR2_X1 U15538 ( .A1(n6579), .A2(n13374), .ZN(n13572) );
  AOI22_X1 U15539 ( .A1(n13375), .A2(n13525), .B1(n13517), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n13376) );
  OAI21_X1 U15540 ( .B1(n13572), .B2(n13498), .A(n13376), .ZN(n13377) );
  AOI21_X1 U15541 ( .B1(n13576), .B2(n13527), .A(n13377), .ZN(n13378) );
  OAI21_X1 U15542 ( .B1(n13379), .B2(n13517), .A(n13378), .ZN(P2_U3242) );
  XNOR2_X1 U15543 ( .A(n13380), .B(n13385), .ZN(n13383) );
  INV_X1 U15544 ( .A(n13381), .ZN(n13382) );
  AOI21_X1 U15545 ( .B1(n13383), .B2(n13484), .A(n13382), .ZN(n13582) );
  OAI21_X1 U15546 ( .B1(n13386), .B2(n13385), .A(n13384), .ZN(n13583) );
  INV_X1 U15547 ( .A(n13583), .ZN(n13394) );
  AOI21_X1 U15548 ( .B1(n13580), .B2(n13402), .A(n13490), .ZN(n13388) );
  AND2_X1 U15549 ( .A1(n13388), .A2(n13387), .ZN(n13579) );
  NAND2_X1 U15550 ( .A1(n13579), .A2(n13529), .ZN(n13391) );
  AOI22_X1 U15551 ( .A1(P2_REG2_REG_22__SCAN_IN), .A2(n13517), .B1(n13389), 
        .B2(n13511), .ZN(n13390) );
  OAI211_X1 U15552 ( .C1(n13392), .C2(n13461), .A(n13391), .B(n13390), .ZN(
        n13393) );
  AOI21_X1 U15553 ( .B1(n13394), .B2(n13527), .A(n13393), .ZN(n13395) );
  OAI21_X1 U15554 ( .B1(n13517), .B2(n13582), .A(n13395), .ZN(P2_U3243) );
  XNOR2_X1 U15555 ( .A(n13396), .B(n13399), .ZN(n13398) );
  OAI21_X1 U15556 ( .B1(n13398), .B2(n13504), .A(n13397), .ZN(n13584) );
  INV_X1 U15557 ( .A(n13584), .ZN(n13410) );
  XNOR2_X1 U15558 ( .A(n13400), .B(n13399), .ZN(n13586) );
  INV_X1 U15559 ( .A(n13402), .ZN(n13403) );
  AOI211_X1 U15560 ( .C1(n13404), .C2(n13414), .A(n13490), .B(n13403), .ZN(
        n13585) );
  NAND2_X1 U15561 ( .A1(n13585), .A2(n13529), .ZN(n13407) );
  AOI22_X1 U15562 ( .A1(n13517), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13405), 
        .B2(n13511), .ZN(n13406) );
  OAI211_X1 U15563 ( .C1(n9542), .C2(n13461), .A(n13407), .B(n13406), .ZN(
        n13408) );
  AOI21_X1 U15564 ( .B1(n13586), .B2(n13527), .A(n13408), .ZN(n13409) );
  OAI21_X1 U15565 ( .B1(n13517), .B2(n13410), .A(n13409), .ZN(P2_U3244) );
  XNOR2_X1 U15566 ( .A(n13411), .B(n13420), .ZN(n13413) );
  AOI21_X1 U15567 ( .B1(n13413), .B2(n13484), .A(n13412), .ZN(n13592) );
  AOI211_X1 U15568 ( .C1(n13590), .C2(n13429), .A(n13490), .B(n13401), .ZN(
        n13589) );
  INV_X1 U15569 ( .A(n13415), .ZN(n13416) );
  AOI22_X1 U15570 ( .A1(n13517), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13416), 
        .B2(n13511), .ZN(n13417) );
  OAI21_X1 U15571 ( .B1(n13418), .B2(n13461), .A(n13417), .ZN(n13422) );
  XNOR2_X1 U15572 ( .A(n13419), .B(n13420), .ZN(n13593) );
  NOR2_X1 U15573 ( .A1(n13593), .A2(n13467), .ZN(n13421) );
  AOI211_X1 U15574 ( .C1(n13589), .C2(n13529), .A(n13422), .B(n13421), .ZN(
        n13423) );
  OAI21_X1 U15575 ( .B1(n13517), .B2(n13592), .A(n13423), .ZN(P2_U3245) );
  XNOR2_X1 U15576 ( .A(n13424), .B(n13426), .ZN(n13598) );
  XOR2_X1 U15577 ( .A(n13426), .B(n13425), .Z(n13428) );
  OAI21_X1 U15578 ( .B1(n13428), .B2(n13504), .A(n13427), .ZN(n13594) );
  NAND2_X1 U15579 ( .A1(n13594), .A2(n13519), .ZN(n13437) );
  INV_X1 U15580 ( .A(n13429), .ZN(n13430) );
  AOI211_X1 U15581 ( .C1(n13596), .C2(n7495), .A(n13490), .B(n13430), .ZN(
        n13595) );
  INV_X1 U15582 ( .A(n13431), .ZN(n13432) );
  AOI22_X1 U15583 ( .A1(n13517), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13432), 
        .B2(n13511), .ZN(n13433) );
  OAI21_X1 U15584 ( .B1(n13434), .B2(n13461), .A(n13433), .ZN(n13435) );
  AOI21_X1 U15585 ( .B1(n13595), .B2(n13529), .A(n13435), .ZN(n13436) );
  OAI211_X1 U15586 ( .C1(n13467), .C2(n13598), .A(n13437), .B(n13436), .ZN(
        P2_U3246) );
  XNOR2_X1 U15587 ( .A(n13438), .B(n13447), .ZN(n13440) );
  AOI21_X1 U15588 ( .B1(n13440), .B2(n13484), .A(n13439), .ZN(n13603) );
  AOI211_X1 U15589 ( .C1(n13601), .C2(n13460), .A(n13490), .B(n6911), .ZN(
        n13600) );
  INV_X1 U15590 ( .A(n13601), .ZN(n13441) );
  NOR2_X1 U15591 ( .A1(n13441), .A2(n13461), .ZN(n13445) );
  INV_X1 U15592 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n13443) );
  OAI22_X1 U15593 ( .A1(n13519), .A2(n13443), .B1(n13442), .B2(n13521), .ZN(
        n13444) );
  AOI211_X1 U15594 ( .C1(n13600), .C2(n13529), .A(n13445), .B(n13444), .ZN(
        n13450) );
  OAI21_X1 U15595 ( .B1(n13448), .B2(n13447), .A(n13446), .ZN(n13599) );
  NAND2_X1 U15596 ( .A1(n13599), .A2(n13527), .ZN(n13449) );
  OAI211_X1 U15597 ( .C1(n13603), .C2(n13517), .A(n13450), .B(n13449), .ZN(
        P2_U3247) );
  INV_X1 U15598 ( .A(n13451), .ZN(n13453) );
  XNOR2_X1 U15599 ( .A(n13452), .B(n13453), .ZN(n13605) );
  INV_X1 U15600 ( .A(n13605), .ZN(n13468) );
  XNOR2_X1 U15601 ( .A(n13454), .B(n13453), .ZN(n13455) );
  NAND2_X1 U15602 ( .A1(n13455), .A2(n13484), .ZN(n13457) );
  NAND2_X1 U15603 ( .A1(n13457), .A2(n13456), .ZN(n13607) );
  NAND2_X1 U15604 ( .A1(n13607), .A2(n13519), .ZN(n13466) );
  OR2_X1 U15605 ( .A1(n13458), .A2(n13665), .ZN(n13459) );
  AND3_X1 U15606 ( .A1(n13460), .A2(n11269), .A3(n13459), .ZN(n13606) );
  NOR2_X1 U15607 ( .A1(n13665), .A2(n13461), .ZN(n13464) );
  OAI22_X1 U15608 ( .A1(n13519), .A2(n13251), .B1(n13462), .B2(n13521), .ZN(
        n13463) );
  AOI211_X1 U15609 ( .C1(n13606), .C2(n13529), .A(n13464), .B(n13463), .ZN(
        n13465) );
  OAI211_X1 U15610 ( .C1(n13468), .C2(n13467), .A(n13466), .B(n13465), .ZN(
        P2_U3248) );
  XNOR2_X1 U15611 ( .A(n13469), .B(n13474), .ZN(n13470) );
  NAND2_X1 U15612 ( .A1(n13470), .A2(n13484), .ZN(n13616) );
  OAI211_X1 U15613 ( .C1(n13521), .C2(n13471), .A(n13616), .B(n13611), .ZN(
        n13481) );
  INV_X1 U15614 ( .A(n13477), .ZN(n13669) );
  XNOR2_X1 U15615 ( .A(n13492), .B(n13669), .ZN(n13472) );
  NAND2_X1 U15616 ( .A1(n13472), .A2(n11269), .ZN(n13612) );
  NAND2_X1 U15617 ( .A1(n13473), .A2(n13474), .ZN(n13475) );
  AND2_X1 U15618 ( .A1(n13476), .A2(n13475), .ZN(n13614) );
  NAND2_X1 U15619 ( .A1(n13614), .A2(n13527), .ZN(n13479) );
  AOI22_X1 U15620 ( .A1(n13477), .A2(n13525), .B1(P2_REG2_REG_16__SCAN_IN), 
        .B2(n13517), .ZN(n13478) );
  OAI211_X1 U15621 ( .C1(n13612), .C2(n13498), .A(n13479), .B(n13478), .ZN(
        n13480) );
  AOI21_X1 U15622 ( .B1(n13481), .B2(n13519), .A(n13480), .ZN(n13482) );
  INV_X1 U15623 ( .A(n13482), .ZN(P2_U3249) );
  XNOR2_X1 U15624 ( .A(n13483), .B(n13486), .ZN(n13485) );
  NAND2_X1 U15625 ( .A1(n13485), .A2(n13484), .ZN(n13620) );
  XNOR2_X1 U15626 ( .A(n13488), .B(n13487), .ZN(n13621) );
  INV_X1 U15627 ( .A(n13621), .ZN(n13500) );
  AOI21_X1 U15628 ( .B1(n13672), .B2(n13508), .A(n13490), .ZN(n13493) );
  AOI21_X1 U15629 ( .B1(n13493), .B2(n13492), .A(n13491), .ZN(n13619) );
  OAI22_X1 U15630 ( .A1(n13519), .A2(n13495), .B1(n13494), .B2(n13521), .ZN(
        n13496) );
  AOI21_X1 U15631 ( .B1(n13672), .B2(n13525), .A(n13496), .ZN(n13497) );
  OAI21_X1 U15632 ( .B1(n13619), .B2(n13498), .A(n13497), .ZN(n13499) );
  AOI21_X1 U15633 ( .B1(n13500), .B2(n13527), .A(n13499), .ZN(n13501) );
  OAI21_X1 U15634 ( .B1(n13620), .B2(n13517), .A(n13501), .ZN(P2_U3250) );
  XOR2_X1 U15635 ( .A(n13506), .B(n13502), .Z(n13505) );
  OAI21_X1 U15636 ( .B1(n13505), .B2(n13504), .A(n13503), .ZN(n13625) );
  INV_X1 U15637 ( .A(n13625), .ZN(n13518) );
  XNOR2_X1 U15638 ( .A(n13507), .B(n13506), .ZN(n13627) );
  AOI211_X1 U15639 ( .C1(n13510), .C2(n13509), .A(n13490), .B(n13489), .ZN(
        n13626) );
  NAND2_X1 U15640 ( .A1(n13626), .A2(n13529), .ZN(n13514) );
  AOI22_X1 U15641 ( .A1(n13517), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n13512), 
        .B2(n13511), .ZN(n13513) );
  OAI211_X1 U15642 ( .C1(n13678), .C2(n13461), .A(n13514), .B(n13513), .ZN(
        n13515) );
  AOI21_X1 U15643 ( .B1(n13527), .B2(n13627), .A(n13515), .ZN(n13516) );
  OAI21_X1 U15644 ( .B1(n13518), .B2(n13517), .A(n13516), .ZN(P2_U3251) );
  NAND2_X1 U15645 ( .A1(n13520), .A2(n13519), .ZN(n13534) );
  OAI22_X1 U15646 ( .A1(n13519), .A2(n13523), .B1(n13522), .B2(n13521), .ZN(
        n13524) );
  AOI21_X1 U15647 ( .B1(n13526), .B2(n13525), .A(n13524), .ZN(n13533) );
  NAND2_X1 U15648 ( .A1(n13528), .A2(n13527), .ZN(n13532) );
  NAND2_X1 U15649 ( .A1(n13530), .A2(n13529), .ZN(n13531) );
  NAND4_X1 U15650 ( .A1(n13534), .A2(n13533), .A3(n13532), .A4(n13531), .ZN(
        P2_U3254) );
  NAND2_X1 U15651 ( .A1(n13535), .A2(n13537), .ZN(n13636) );
  MUX2_X1 U15652 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13636), .S(n15002), .Z(
        n13536) );
  MUX2_X1 U15653 ( .A(n13639), .B(n13539), .S(n6478), .Z(n13540) );
  OAI21_X1 U15654 ( .B1(n13641), .B2(n13630), .A(n13540), .ZN(P2_U3529) );
  AOI21_X1 U15655 ( .B1(n14972), .B2(n13542), .A(n13541), .ZN(n13543) );
  MUX2_X1 U15656 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13643), .S(n15002), .Z(
        P2_U3527) );
  AOI211_X1 U15657 ( .C1(n13552), .C2(n14982), .A(n13551), .B(n13550), .ZN(
        n13644) );
  MUX2_X1 U15658 ( .A(n13553), .B(n13644), .S(n15002), .Z(n13554) );
  OAI21_X1 U15659 ( .B1(n13647), .B2(n13630), .A(n13554), .ZN(P2_U3526) );
  AOI211_X1 U15660 ( .C1(n14972), .C2(n13557), .A(n13556), .B(n13555), .ZN(
        n13558) );
  OAI21_X1 U15661 ( .B1(n13559), .B2(n13622), .A(n13558), .ZN(n13648) );
  MUX2_X1 U15662 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13648), .S(n15002), .Z(
        P2_U3525) );
  INV_X1 U15663 ( .A(n13560), .ZN(n13565) );
  AOI21_X1 U15664 ( .B1(n14972), .B2(n13562), .A(n13561), .ZN(n13563) );
  OAI211_X1 U15665 ( .C1(n13565), .C2(n13622), .A(n13564), .B(n13563), .ZN(
        n13649) );
  MUX2_X1 U15666 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13649), .S(n15002), .Z(
        P2_U3524) );
  NAND2_X1 U15667 ( .A1(n13566), .A2(n14982), .ZN(n13571) );
  NAND2_X1 U15668 ( .A1(n13567), .A2(n14972), .ZN(n13568) );
  NAND4_X1 U15669 ( .A1(n13571), .A2(n13570), .A3(n13569), .A4(n13568), .ZN(
        n13650) );
  MUX2_X1 U15670 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13650), .S(n15002), .Z(
        P2_U3523) );
  INV_X1 U15671 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n13577) );
  NAND3_X1 U15672 ( .A1(n13574), .A2(n13573), .A3(n13572), .ZN(n13575) );
  AOI21_X1 U15673 ( .B1(n13576), .B2(n14982), .A(n13575), .ZN(n13651) );
  MUX2_X1 U15674 ( .A(n13577), .B(n13651), .S(n15002), .Z(n13578) );
  OAI21_X1 U15675 ( .B1(n13654), .B2(n13630), .A(n13578), .ZN(P2_U3522) );
  AOI21_X1 U15676 ( .B1(n14972), .B2(n13580), .A(n13579), .ZN(n13581) );
  OAI211_X1 U15677 ( .C1(n13583), .C2(n13622), .A(n13582), .B(n13581), .ZN(
        n13655) );
  MUX2_X1 U15678 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13655), .S(n15002), .Z(
        P2_U3521) );
  AOI211_X1 U15679 ( .C1(n13586), .C2(n14982), .A(n13585), .B(n13584), .ZN(
        n13656) );
  MUX2_X1 U15680 ( .A(n13587), .B(n13656), .S(n15002), .Z(n13588) );
  OAI21_X1 U15681 ( .B1(n9542), .B2(n13630), .A(n13588), .ZN(P2_U3520) );
  AOI21_X1 U15682 ( .B1(n14972), .B2(n13590), .A(n13589), .ZN(n13591) );
  OAI211_X1 U15683 ( .C1(n13593), .C2(n13622), .A(n13592), .B(n13591), .ZN(
        n13659) );
  MUX2_X1 U15684 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13659), .S(n15002), .Z(
        P2_U3519) );
  AOI211_X1 U15685 ( .C1(n14972), .C2(n13596), .A(n13595), .B(n13594), .ZN(
        n13597) );
  OAI21_X1 U15686 ( .B1(n13622), .B2(n13598), .A(n13597), .ZN(n13660) );
  MUX2_X1 U15687 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13660), .S(n15002), .Z(
        P2_U3518) );
  INV_X1 U15688 ( .A(n13599), .ZN(n13604) );
  AOI21_X1 U15689 ( .B1(n14972), .B2(n13601), .A(n13600), .ZN(n13602) );
  OAI211_X1 U15690 ( .C1(n13604), .C2(n13622), .A(n13603), .B(n13602), .ZN(
        n13661) );
  MUX2_X1 U15691 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13661), .S(n15002), .Z(
        P2_U3517) );
  AND2_X1 U15692 ( .A1(n13605), .A2(n14982), .ZN(n13608) );
  NOR3_X1 U15693 ( .A1(n13608), .A2(n13607), .A3(n13606), .ZN(n13663) );
  MUX2_X1 U15694 ( .A(n13663), .B(n13609), .S(n6478), .Z(n13610) );
  OAI21_X1 U15695 ( .B1(n13665), .B2(n13630), .A(n13610), .ZN(P2_U3516) );
  INV_X1 U15696 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n13617) );
  NAND2_X1 U15697 ( .A1(n13612), .A2(n13611), .ZN(n13613) );
  AOI21_X1 U15698 ( .B1(n13614), .B2(n14982), .A(n13613), .ZN(n13615) );
  AND2_X1 U15699 ( .A1(n13616), .A2(n13615), .ZN(n13666) );
  MUX2_X1 U15700 ( .A(n13617), .B(n13666), .S(n15002), .Z(n13618) );
  OAI21_X1 U15701 ( .B1(n13669), .B2(n13630), .A(n13618), .ZN(P2_U3515) );
  OAI211_X1 U15702 ( .C1(n13622), .C2(n13621), .A(n13620), .B(n13619), .ZN(
        n13670) );
  MUX2_X1 U15703 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13670), .S(n15002), .Z(
        n13623) );
  AOI21_X1 U15704 ( .B1(n13634), .B2(n13672), .A(n13623), .ZN(n13624) );
  INV_X1 U15705 ( .A(n13624), .ZN(P2_U3514) );
  INV_X1 U15706 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n13628) );
  AOI211_X1 U15707 ( .C1(n13627), .C2(n14982), .A(n13626), .B(n13625), .ZN(
        n13674) );
  MUX2_X1 U15708 ( .A(n13628), .B(n13674), .S(n15002), .Z(n13629) );
  OAI21_X1 U15709 ( .B1(n13678), .B2(n13630), .A(n13629), .ZN(P2_U3513) );
  AOI211_X1 U15710 ( .C1(n13633), .C2(n14982), .A(n13632), .B(n13631), .ZN(
        n13682) );
  AOI22_X1 U15711 ( .A1(n14830), .A2(n13634), .B1(n6478), .B2(
        P2_REG1_REG_13__SCAN_IN), .ZN(n13635) );
  OAI21_X1 U15712 ( .B1(n13682), .B2(n6478), .A(n13635), .ZN(P2_U3512) );
  MUX2_X1 U15713 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13636), .S(n14995), .Z(
        n13637) );
  INV_X1 U15714 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n13638) );
  MUX2_X1 U15715 ( .A(n13639), .B(n13638), .S(n14994), .Z(n13640) );
  OAI21_X1 U15716 ( .B1(n13641), .B2(n13677), .A(n13640), .ZN(P2_U3497) );
  MUX2_X1 U15717 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13642), .S(n14995), .Z(
        P2_U3496) );
  MUX2_X1 U15718 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13643), .S(n14995), .Z(
        P2_U3495) );
  INV_X1 U15719 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n13645) );
  MUX2_X1 U15720 ( .A(n13645), .B(n13644), .S(n14995), .Z(n13646) );
  OAI21_X1 U15721 ( .B1(n13647), .B2(n13677), .A(n13646), .ZN(P2_U3494) );
  MUX2_X1 U15722 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13648), .S(n14995), .Z(
        P2_U3493) );
  MUX2_X1 U15723 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13649), .S(n14995), .Z(
        P2_U3492) );
  MUX2_X1 U15724 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13650), .S(n14995), .Z(
        P2_U3491) );
  MUX2_X1 U15725 ( .A(n13652), .B(n13651), .S(n14995), .Z(n13653) );
  OAI21_X1 U15726 ( .B1(n13654), .B2(n13677), .A(n13653), .ZN(P2_U3490) );
  MUX2_X1 U15727 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13655), .S(n14995), .Z(
        P2_U3489) );
  INV_X1 U15728 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n13657) );
  MUX2_X1 U15729 ( .A(n13657), .B(n13656), .S(n14995), .Z(n13658) );
  OAI21_X1 U15730 ( .B1(n9542), .B2(n13677), .A(n13658), .ZN(P2_U3488) );
  MUX2_X1 U15731 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13659), .S(n14995), .Z(
        P2_U3487) );
  MUX2_X1 U15732 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13660), .S(n14995), .Z(
        P2_U3486) );
  MUX2_X1 U15733 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13661), .S(n14995), .Z(
        P2_U3484) );
  INV_X1 U15734 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n13662) );
  MUX2_X1 U15735 ( .A(n13663), .B(n13662), .S(n14994), .Z(n13664) );
  OAI21_X1 U15736 ( .B1(n13665), .B2(n13677), .A(n13664), .ZN(P2_U3481) );
  MUX2_X1 U15737 ( .A(n13667), .B(n13666), .S(n14995), .Z(n13668) );
  OAI21_X1 U15738 ( .B1(n13669), .B2(n13677), .A(n13668), .ZN(P2_U3478) );
  MUX2_X1 U15739 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13670), .S(n14995), .Z(
        n13671) );
  AOI21_X1 U15740 ( .B1(n13680), .B2(n13672), .A(n13671), .ZN(n13673) );
  INV_X1 U15741 ( .A(n13673), .ZN(P2_U3475) );
  MUX2_X1 U15742 ( .A(n13675), .B(n13674), .S(n14995), .Z(n13676) );
  OAI21_X1 U15743 ( .B1(n13678), .B2(n13677), .A(n13676), .ZN(P2_U3472) );
  NOR2_X1 U15744 ( .A1(n14995), .A2(n9280), .ZN(n13679) );
  AOI21_X1 U15745 ( .B1(n14830), .B2(n13680), .A(n13679), .ZN(n13681) );
  OAI21_X1 U15746 ( .B1(n13682), .B2(n14994), .A(n13681), .ZN(P2_U3469) );
  NAND3_X1 U15747 ( .A1(n13685), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n13687) );
  OAI22_X1 U15748 ( .A1(n13684), .A2(n13687), .B1(n13686), .B2(n13705), .ZN(
        n13688) );
  AOI21_X1 U15749 ( .B1(n13683), .B2(n13694), .A(n13688), .ZN(n13689) );
  INV_X1 U15750 ( .A(n13689), .ZN(P2_U3296) );
  OAI222_X1 U15751 ( .A1(P2_U3088), .A2(n9062), .B1(n13708), .B2(n14219), .C1(
        n13690), .C2(n13705), .ZN(P2_U3297) );
  OAI222_X1 U15752 ( .A1(P2_U3088), .A2(n13693), .B1(n13708), .B2(n13692), 
        .C1(n13691), .C2(n13705), .ZN(P2_U3298) );
  NAND2_X1 U15753 ( .A1(n13695), .A2(n13694), .ZN(n13697) );
  OAI211_X1 U15754 ( .C1(n13705), .C2(n13698), .A(n13697), .B(n13696), .ZN(
        P2_U3299) );
  INV_X1 U15755 ( .A(n13699), .ZN(n14221) );
  INV_X1 U15756 ( .A(n13702), .ZN(n14224) );
  OAI222_X1 U15757 ( .A1(P2_U3088), .A2(n13704), .B1(n13708), .B2(n14224), 
        .C1(n13703), .C2(n13705), .ZN(P2_U3301) );
  OAI222_X1 U15758 ( .A1(n13710), .A2(P2_U3088), .B1(n13708), .B2(n13707), 
        .C1(n13706), .C2(n13705), .ZN(P2_U3302) );
  INV_X1 U15759 ( .A(n13711), .ZN(n13712) );
  MUX2_X1 U15760 ( .A(n13712), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  AOI21_X1 U15761 ( .B1(n13715), .B2(n13714), .A(n13713), .ZN(n13721) );
  OAI21_X1 U15762 ( .B1(n13811), .B2(n14113), .A(n13716), .ZN(n13717) );
  AOI21_X1 U15763 ( .B1(n13814), .B2(n14114), .A(n13717), .ZN(n13718) );
  OAI21_X1 U15764 ( .B1(n14606), .B2(n14118), .A(n13718), .ZN(n13719) );
  AOI21_X1 U15765 ( .B1(n14545), .B2(n13794), .A(n13719), .ZN(n13720) );
  OAI21_X1 U15766 ( .B1(n13721), .B2(n14593), .A(n13720), .ZN(P1_U3215) );
  OAI21_X1 U15767 ( .B1(n13724), .B2(n13723), .A(n13722), .ZN(n13725) );
  NAND2_X1 U15768 ( .A1(n13725), .A2(n14488), .ZN(n13730) );
  INV_X1 U15769 ( .A(n14007), .ZN(n13728) );
  AOI22_X1 U15770 ( .A1(n14596), .A2(n14032), .B1(n13847), .B2(n14597), .ZN(
        n14004) );
  INV_X1 U15771 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n13726) );
  OAI22_X1 U15772 ( .A1(n14004), .A2(n13836), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13726), .ZN(n13727) );
  AOI21_X1 U15773 ( .B1(n13834), .B2(n13728), .A(n13727), .ZN(n13729) );
  OAI211_X1 U15774 ( .C1(n14012), .C2(n13817), .A(n13730), .B(n13729), .ZN(
        P1_U3216) );
  INV_X1 U15775 ( .A(n14181), .ZN(n14072) );
  AND2_X1 U15776 ( .A1(n13806), .A2(n13731), .ZN(n13734) );
  OAI211_X1 U15777 ( .C1(n13734), .C2(n13733), .A(n14488), .B(n13732), .ZN(
        n13738) );
  NOR2_X1 U15778 ( .A1(n14606), .A2(n14069), .ZN(n13736) );
  NAND2_X1 U15779 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13917)
         );
  OAI21_X1 U15780 ( .B1(n14034), .B2(n13811), .A(n13917), .ZN(n13735) );
  AOI211_X1 U15781 ( .C1(n13814), .C2(n14066), .A(n13736), .B(n13735), .ZN(
        n13737) );
  OAI211_X1 U15782 ( .C1(n14072), .C2(n13817), .A(n13738), .B(n13737), .ZN(
        P1_U3219) );
  OAI21_X1 U15783 ( .B1(n13741), .B2(n13740), .A(n13739), .ZN(n13742) );
  NAND2_X1 U15784 ( .A1(n13742), .A2(n14488), .ZN(n13746) );
  AOI22_X1 U15785 ( .A1(n13789), .A2(n14032), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13743) );
  OAI21_X1 U15786 ( .B1(n14034), .B2(n13763), .A(n13743), .ZN(n13744) );
  AOI21_X1 U15787 ( .B1(n14043), .B2(n13834), .A(n13744), .ZN(n13745) );
  OAI211_X1 U15788 ( .C1(n6939), .C2(n13817), .A(n13746), .B(n13745), .ZN(
        P1_U3223) );
  INV_X1 U15789 ( .A(n14147), .ZN(n13972) );
  INV_X1 U15790 ( .A(n13747), .ZN(n13752) );
  NOR3_X1 U15791 ( .A1(n13748), .A2(n13750), .A3(n13749), .ZN(n13751) );
  OAI21_X1 U15792 ( .B1(n13752), .B2(n13751), .A(n14488), .ZN(n13757) );
  INV_X1 U15793 ( .A(n13753), .ZN(n13969) );
  AOI22_X1 U15794 ( .A1(n14596), .A2(n13847), .B1(n13845), .B2(n14597), .ZN(
        n13965) );
  OAI22_X1 U15795 ( .A1(n13965), .A2(n13836), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13754), .ZN(n13755) );
  AOI21_X1 U15796 ( .B1(n13834), .B2(n13969), .A(n13755), .ZN(n13756) );
  OAI211_X1 U15797 ( .C1(n13972), .C2(n13817), .A(n13757), .B(n13756), .ZN(
        P1_U3225) );
  AOI21_X1 U15798 ( .B1(n6676), .B2(n13759), .A(n13758), .ZN(n13767) );
  NAND2_X1 U15799 ( .A1(n13789), .A2(n14497), .ZN(n13762) );
  OAI211_X1 U15800 ( .C1(n13763), .C2(n14113), .A(n13762), .B(n13761), .ZN(
        n13764) );
  AOI21_X1 U15801 ( .B1(n14508), .B2(n13834), .A(n13764), .ZN(n13766) );
  NAND2_X1 U15802 ( .A1(n14531), .A2(n13794), .ZN(n13765) );
  OAI211_X1 U15803 ( .C1(n13767), .C2(n14593), .A(n13766), .B(n13765), .ZN(
        P1_U3226) );
  INV_X1 U15804 ( .A(n13768), .ZN(n13772) );
  NOR3_X1 U15805 ( .A1(n13758), .A2(n13770), .A3(n13769), .ZN(n13771) );
  OAI21_X1 U15806 ( .B1(n13772), .B2(n13771), .A(n14488), .ZN(n13778) );
  NAND2_X1 U15807 ( .A1(n14066), .A2(n14597), .ZN(n13774) );
  NAND2_X1 U15808 ( .A1(n13850), .A2(n14596), .ZN(n13773) );
  NAND2_X1 U15809 ( .A1(n13774), .A2(n13773), .ZN(n14097) );
  NOR2_X1 U15810 ( .A1(n14606), .A2(n14100), .ZN(n13775) );
  AOI211_X1 U15811 ( .C1(n14601), .C2(n14097), .A(n13776), .B(n13775), .ZN(
        n13777) );
  OAI211_X1 U15812 ( .C1(n14104), .C2(n13817), .A(n13778), .B(n13777), .ZN(
        P1_U3228) );
  AND3_X1 U15813 ( .A1(n13722), .A2(n13780), .A3(n13779), .ZN(n13781) );
  OAI21_X1 U15814 ( .B1(n13748), .B2(n13781), .A(n14488), .ZN(n13786) );
  INV_X1 U15815 ( .A(n13782), .ZN(n13988) );
  AOI22_X1 U15816 ( .A1(n14596), .A2(n13848), .B1(n13846), .B2(n14597), .ZN(
        n13983) );
  INV_X1 U15817 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n13783) );
  OAI22_X1 U15818 ( .A1(n13983), .A2(n13836), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13783), .ZN(n13784) );
  AOI21_X1 U15819 ( .B1(n13834), .B2(n13988), .A(n13784), .ZN(n13785) );
  OAI211_X1 U15820 ( .C1(n13990), .C2(n13817), .A(n13786), .B(n13785), .ZN(
        P1_U3229) );
  XNOR2_X1 U15821 ( .A(n13788), .B(n13787), .ZN(n13796) );
  AOI22_X1 U15822 ( .A1(n14050), .A2(n13789), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13791) );
  NAND2_X1 U15823 ( .A1(n13814), .A2(n14081), .ZN(n13790) );
  OAI211_X1 U15824 ( .C1(n14606), .C2(n13792), .A(n13791), .B(n13790), .ZN(
        n13793) );
  AOI21_X1 U15825 ( .B1(n14058), .B2(n13794), .A(n13793), .ZN(n13795) );
  OAI21_X1 U15826 ( .B1(n13796), .B2(n14593), .A(n13795), .ZN(P1_U3233) );
  OAI21_X1 U15827 ( .B1(n13799), .B2(n13798), .A(n13797), .ZN(n13800) );
  NAND2_X1 U15828 ( .A1(n13800), .A2(n14488), .ZN(n13805) );
  INV_X1 U15829 ( .A(n13801), .ZN(n14023) );
  AOI22_X1 U15830 ( .A1(n14050), .A2(n14596), .B1(n14597), .B2(n13848), .ZN(
        n14017) );
  INV_X1 U15831 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13802) );
  OAI22_X1 U15832 ( .A1(n14017), .A2(n13836), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13802), .ZN(n13803) );
  AOI21_X1 U15833 ( .B1(n14023), .B2(n13834), .A(n13803), .ZN(n13804) );
  OAI211_X1 U15834 ( .C1(n13817), .C2(n14025), .A(n13805), .B(n13804), .ZN(
        P1_U3235) );
  OAI21_X1 U15835 ( .B1(n13808), .B2(n13807), .A(n13806), .ZN(n13809) );
  NAND2_X1 U15836 ( .A1(n13809), .A2(n14488), .ZN(n13816) );
  NOR2_X1 U15837 ( .A1(n14606), .A2(n14085), .ZN(n13813) );
  NAND2_X1 U15838 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13894)
         );
  OAI21_X1 U15839 ( .B1(n13811), .B2(n13810), .A(n13894), .ZN(n13812) );
  AOI211_X1 U15840 ( .C1(n13814), .C2(n14497), .A(n13813), .B(n13812), .ZN(
        n13815) );
  OAI211_X1 U15841 ( .C1(n14188), .C2(n13817), .A(n13816), .B(n13815), .ZN(
        P1_U3238) );
  NAND2_X1 U15842 ( .A1(n13960), .A2(n14761), .ZN(n14141) );
  INV_X1 U15843 ( .A(n14592), .ZN(n14480) );
  OAI21_X1 U15844 ( .B1(n13820), .B2(n13819), .A(n13818), .ZN(n13821) );
  NAND2_X1 U15845 ( .A1(n13821), .A2(n14488), .ZN(n13828) );
  INV_X1 U15846 ( .A(n13954), .ZN(n13826) );
  NAND2_X1 U15847 ( .A1(n13844), .A2(n14498), .ZN(n13823) );
  NAND2_X1 U15848 ( .A1(n13846), .A2(n14596), .ZN(n13822) );
  AND2_X1 U15849 ( .A1(n13823), .A2(n13822), .ZN(n14143) );
  OAI22_X1 U15850 ( .A1(n13836), .A2(n14143), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13824), .ZN(n13825) );
  AOI21_X1 U15851 ( .B1(n13834), .B2(n13826), .A(n13825), .ZN(n13827) );
  OAI211_X1 U15852 ( .C1(n14141), .C2(n14480), .A(n13828), .B(n13827), .ZN(
        P1_U3240) );
  AOI21_X1 U15853 ( .B1(n13831), .B2(n13830), .A(n13829), .ZN(n13840) );
  NOR2_X1 U15854 ( .A1(n13832), .A2(n14781), .ZN(n14541) );
  NAND2_X1 U15855 ( .A1(n13834), .A2(n13833), .ZN(n13835) );
  NAND2_X1 U15856 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14651)
         );
  OAI211_X1 U15857 ( .C1(n13837), .C2(n13836), .A(n13835), .B(n14651), .ZN(
        n13838) );
  AOI21_X1 U15858 ( .B1(n14541), .B2(n14592), .A(n13838), .ZN(n13839) );
  OAI21_X1 U15859 ( .B1(n13840), .B2(n14593), .A(n13839), .ZN(P1_U3241) );
  MUX2_X1 U15860 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13920), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15861 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13841), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15862 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13842), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15863 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13843), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15864 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13844), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15865 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13845), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15866 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13846), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15867 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13847), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15868 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13848), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15869 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14032), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15870 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14050), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15871 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14067), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15872 ( .A(n14081), .B(P1_DATAO_REG_19__SCAN_IN), .S(n13849), .Z(
        P1_U3579) );
  MUX2_X1 U15873 ( .A(n14066), .B(P1_DATAO_REG_18__SCAN_IN), .S(n13849), .Z(
        P1_U3578) );
  MUX2_X1 U15874 ( .A(n14497), .B(P1_DATAO_REG_17__SCAN_IN), .S(n13849), .Z(
        P1_U3577) );
  MUX2_X1 U15875 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13850), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U15876 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14499), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15877 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14114), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U15878 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13851), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U15879 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13852), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U15880 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13853), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U15881 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13854), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U15882 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13855), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U15883 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13856), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U15884 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13857), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U15885 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13858), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U15886 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14598), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U15887 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13859), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U15888 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n12090), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U15889 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n13860), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U15890 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n13861), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI211_X1 U15891 ( .C1(n13864), .C2(n13863), .A(n14648), .B(n13862), .ZN(
        n13873) );
  OAI211_X1 U15892 ( .C1(n9982), .C2(n13867), .A(n14649), .B(n13866), .ZN(
        n13872) );
  AOI22_X1 U15893 ( .A1(n14615), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n13871) );
  INV_X1 U15894 ( .A(n13868), .ZN(n13869) );
  NAND2_X1 U15895 ( .A1(n14645), .A2(n13869), .ZN(n13870) );
  NAND4_X1 U15896 ( .A1(n13873), .A2(n13872), .A3(n13871), .A4(n13870), .ZN(
        P1_U3244) );
  AND2_X1 U15897 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n13875) );
  NOR2_X1 U15898 ( .A1(n14634), .A2(n13878), .ZN(n13874) );
  AOI211_X1 U15899 ( .C1(n14615), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n13875), .B(
        n13874), .ZN(n13885) );
  OAI211_X1 U15900 ( .C1(n13877), .C2(n13876), .A(n14648), .B(n14628), .ZN(
        n13884) );
  MUX2_X1 U15901 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n14720), .S(n13878), .Z(
        n13879) );
  NAND3_X1 U15902 ( .A1(n13881), .A2(n13880), .A3(n13879), .ZN(n13882) );
  NAND3_X1 U15903 ( .A1(n14649), .A2(n14622), .A3(n13882), .ZN(n13883) );
  NAND3_X1 U15904 ( .A1(n13885), .A2(n13884), .A3(n13883), .ZN(P1_U3246) );
  INV_X1 U15905 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n13888) );
  OAI21_X1 U15906 ( .B1(n13888), .B2(n13887), .A(n13886), .ZN(n13904) );
  XNOR2_X1 U15907 ( .A(n13904), .B(n13903), .ZN(n13901) );
  INV_X1 U15908 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14086) );
  XNOR2_X1 U15909 ( .A(n13901), .B(n14086), .ZN(n13900) );
  AND2_X1 U15910 ( .A1(n13892), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n13909) );
  INV_X1 U15911 ( .A(n13909), .ZN(n13891) );
  OAI211_X1 U15912 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n13892), .A(n13891), 
        .B(n14648), .ZN(n13898) );
  NAND2_X1 U15913 ( .A1(n14615), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n13893) );
  OAI211_X1 U15914 ( .C1(n14634), .C2(n13895), .A(n13894), .B(n13893), .ZN(
        n13896) );
  INV_X1 U15915 ( .A(n13896), .ZN(n13897) );
  OAI211_X1 U15916 ( .C1(n13900), .C2(n13899), .A(n13898), .B(n13897), .ZN(
        P1_U3261) );
  INV_X1 U15917 ( .A(n13901), .ZN(n13902) );
  NAND2_X1 U15918 ( .A1(n13902), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n13906) );
  NAND2_X1 U15919 ( .A1(n13904), .A2(n13903), .ZN(n13905) );
  NAND2_X1 U15920 ( .A1(n13906), .A2(n13905), .ZN(n13907) );
  XOR2_X1 U15921 ( .A(n13907), .B(P1_REG2_REG_19__SCAN_IN), .Z(n13914) );
  INV_X1 U15922 ( .A(n13914), .ZN(n13912) );
  NOR2_X1 U15923 ( .A1(n13909), .A2(n13908), .ZN(n13910) );
  XNOR2_X1 U15924 ( .A(n13910), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n13913) );
  AOI22_X1 U15925 ( .A1(n13914), .A2(n14649), .B1(n14648), .B2(n13913), .ZN(
        n13916) );
  NAND2_X1 U15926 ( .A1(n13926), .A2(n14134), .ZN(n13925) );
  XNOR2_X1 U15927 ( .A(n14131), .B(n13925), .ZN(n13918) );
  NOR2_X1 U15929 ( .A1(n14721), .A2(n13919), .ZN(n13922) );
  NAND2_X1 U15930 ( .A1(n13921), .A2(n13920), .ZN(n14132) );
  NOR2_X1 U15931 ( .A1(n14701), .A2(n14132), .ZN(n13928) );
  AOI211_X1 U15932 ( .C1(n13923), .C2(n14723), .A(n13922), .B(n13928), .ZN(
        n13924) );
  OAI21_X1 U15933 ( .B1(n14130), .B2(n14088), .A(n13924), .ZN(P1_U3263) );
  OAI211_X1 U15934 ( .C1(n13926), .C2(n14134), .A(n14726), .B(n13925), .ZN(
        n14133) );
  NOR2_X1 U15935 ( .A1(n14134), .A2(n14103), .ZN(n13927) );
  AOI211_X1 U15936 ( .C1(n14736), .C2(P1_REG2_REG_30__SCAN_IN), .A(n13928), 
        .B(n13927), .ZN(n13929) );
  OAI21_X1 U15937 ( .B1(n14088), .B2(n14133), .A(n13929), .ZN(P1_U3264) );
  OAI21_X1 U15938 ( .B1(n13941), .B2(n13931), .A(n13930), .ZN(n13934) );
  INV_X1 U15939 ( .A(n13932), .ZN(n13933) );
  AOI211_X1 U15940 ( .C1(n14137), .C2(n13956), .A(n14792), .B(n6944), .ZN(
        n14136) );
  AOI22_X1 U15941 ( .A1(n14701), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n13936), 
        .B2(n14702), .ZN(n13937) );
  OAI21_X1 U15942 ( .B1(n13938), .B2(n14103), .A(n13937), .ZN(n13943) );
  AOI21_X1 U15943 ( .B1(n13941), .B2(n13940), .A(n13939), .ZN(n14140) );
  NOR2_X1 U15944 ( .A1(n14140), .A2(n14107), .ZN(n13942) );
  AOI211_X1 U15945 ( .C1(n14136), .C2(n14731), .A(n13943), .B(n13942), .ZN(
        n13944) );
  OAI21_X1 U15946 ( .B1(n14736), .B2(n14139), .A(n13944), .ZN(P1_U3266) );
  OAI21_X1 U15947 ( .B1(n13947), .B2(n13946), .A(n13945), .ZN(n14146) );
  OAI21_X1 U15948 ( .B1(n13950), .B2(n13949), .A(n13948), .ZN(n13951) );
  NAND2_X1 U15949 ( .A1(n13951), .A2(n14716), .ZN(n14144) );
  INV_X1 U15950 ( .A(n14144), .ZN(n13953) );
  INV_X1 U15951 ( .A(n14143), .ZN(n13952) );
  OAI21_X1 U15952 ( .B1(n13953), .B2(n13952), .A(n14721), .ZN(n13962) );
  INV_X1 U15953 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n13955) );
  OAI22_X1 U15954 ( .A1(n14721), .A2(n13955), .B1(n13954), .B2(n14719), .ZN(
        n13959) );
  AOI21_X1 U15955 ( .B1(n13960), .B2(n13970), .A(n14792), .ZN(n13957) );
  NAND2_X1 U15956 ( .A1(n13957), .A2(n13956), .ZN(n14142) );
  NOR2_X1 U15957 ( .A1(n14142), .A2(n14088), .ZN(n13958) );
  AOI211_X1 U15958 ( .C1(n14723), .C2(n13960), .A(n13959), .B(n13958), .ZN(
        n13961) );
  OAI211_X1 U15959 ( .C1(n14146), .C2(n14107), .A(n13962), .B(n13961), .ZN(
        P1_U3267) );
  OAI21_X1 U15960 ( .B1(n13975), .B2(n13964), .A(n13963), .ZN(n13967) );
  INV_X1 U15961 ( .A(n13965), .ZN(n13966) );
  AOI21_X1 U15962 ( .B1(n13967), .B2(n14716), .A(n13966), .ZN(n14153) );
  INV_X1 U15963 ( .A(n14153), .ZN(n13968) );
  AOI21_X1 U15964 ( .B1(n13969), .B2(n14702), .A(n13968), .ZN(n13979) );
  AOI21_X1 U15965 ( .B1(n14147), .B2(n13986), .A(n6946), .ZN(n14148) );
  OAI22_X1 U15966 ( .A1(n13972), .A2(n14103), .B1(n13971), .B2(n14721), .ZN(
        n13973) );
  AOI21_X1 U15967 ( .B1(n14148), .B2(n13974), .A(n13973), .ZN(n13978) );
  NAND2_X1 U15968 ( .A1(n13976), .A2(n13975), .ZN(n14149) );
  NAND3_X1 U15969 ( .A1(n14150), .A2(n14149), .A3(n14527), .ZN(n13977) );
  OAI211_X1 U15970 ( .C1(n13979), .C2(n14701), .A(n13978), .B(n13977), .ZN(
        P1_U3268) );
  AOI211_X1 U15971 ( .C1(n13982), .C2(n13981), .A(n14691), .B(n13980), .ZN(
        n13985) );
  INV_X1 U15972 ( .A(n13983), .ZN(n13984) );
  NOR2_X1 U15973 ( .A1(n13985), .A2(n13984), .ZN(n14157) );
  INV_X1 U15974 ( .A(n13986), .ZN(n13987) );
  AOI211_X1 U15975 ( .C1(n14155), .C2(n14009), .A(n14792), .B(n13987), .ZN(
        n14154) );
  AOI22_X1 U15976 ( .A1(n14701), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n13988), 
        .B2(n14702), .ZN(n13989) );
  OAI21_X1 U15977 ( .B1(n13990), .B2(n14103), .A(n13989), .ZN(n13996) );
  INV_X1 U15978 ( .A(n13991), .ZN(n13992) );
  AOI21_X1 U15979 ( .B1(n13994), .B2(n13993), .A(n13992), .ZN(n14158) );
  NOR2_X1 U15980 ( .A1(n14158), .A2(n14107), .ZN(n13995) );
  AOI211_X1 U15981 ( .C1(n14154), .C2(n14731), .A(n13996), .B(n13995), .ZN(
        n13997) );
  OAI21_X1 U15982 ( .B1(n14157), .B2(n14701), .A(n13997), .ZN(P1_U3269) );
  NAND2_X1 U15983 ( .A1(n13998), .A2(n14002), .ZN(n13999) );
  NAND2_X1 U15984 ( .A1(n14000), .A2(n13999), .ZN(n14163) );
  OAI21_X1 U15985 ( .B1(n14003), .B2(n14002), .A(n14001), .ZN(n14006) );
  INV_X1 U15986 ( .A(n14004), .ZN(n14005) );
  AOI21_X1 U15987 ( .B1(n14006), .B2(n14716), .A(n14005), .ZN(n14162) );
  OAI21_X1 U15988 ( .B1(n14007), .B2(n14719), .A(n14162), .ZN(n14008) );
  NAND2_X1 U15989 ( .A1(n14008), .A2(n14721), .ZN(n14015) );
  INV_X1 U15990 ( .A(n14009), .ZN(n14010) );
  AOI211_X1 U15991 ( .C1(n14160), .C2(n14021), .A(n14792), .B(n14010), .ZN(
        n14159) );
  OAI22_X1 U15992 ( .A1(n14012), .A2(n14103), .B1(n14011), .B2(n14721), .ZN(
        n14013) );
  AOI21_X1 U15993 ( .B1(n14159), .B2(n14731), .A(n14013), .ZN(n14014) );
  OAI211_X1 U15994 ( .C1(n14163), .C2(n14107), .A(n14015), .B(n14014), .ZN(
        P1_U3270) );
  XNOR2_X1 U15995 ( .A(n14016), .B(n14027), .ZN(n14019) );
  INV_X1 U15996 ( .A(n14017), .ZN(n14018) );
  AOI21_X1 U15997 ( .B1(n14019), .B2(n14716), .A(n14018), .ZN(n14167) );
  INV_X1 U15998 ( .A(n14020), .ZN(n14042) );
  INV_X1 U15999 ( .A(n14021), .ZN(n14022) );
  AOI211_X1 U16000 ( .C1(n14165), .C2(n14042), .A(n14792), .B(n14022), .ZN(
        n14164) );
  AOI22_X1 U16001 ( .A1(n14701), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n14023), 
        .B2(n14702), .ZN(n14024) );
  OAI21_X1 U16002 ( .B1(n14025), .B2(n14103), .A(n14024), .ZN(n14029) );
  XOR2_X1 U16003 ( .A(n14026), .B(n14027), .Z(n14168) );
  NOR2_X1 U16004 ( .A1(n14168), .A2(n14107), .ZN(n14028) );
  AOI211_X1 U16005 ( .C1(n14164), .C2(n14731), .A(n14029), .B(n14028), .ZN(
        n14030) );
  OAI21_X1 U16006 ( .B1(n14736), .B2(n14167), .A(n14030), .ZN(P1_U3271) );
  XNOR2_X1 U16007 ( .A(n14031), .B(n14037), .ZN(n14036) );
  INV_X1 U16008 ( .A(n14032), .ZN(n14033) );
  OAI22_X1 U16009 ( .A1(n14034), .A2(n14696), .B1(n14033), .B2(n14694), .ZN(
        n14035) );
  AOI21_X1 U16010 ( .B1(n14036), .B2(n14716), .A(n14035), .ZN(n14173) );
  NAND2_X1 U16011 ( .A1(n14038), .A2(n14037), .ZN(n14039) );
  NAND2_X1 U16012 ( .A1(n14040), .A2(n14039), .ZN(n14171) );
  NAND2_X1 U16013 ( .A1(n14044), .A2(n14054), .ZN(n14041) );
  NAND3_X1 U16014 ( .A1(n14042), .A2(n14726), .A3(n14041), .ZN(n14169) );
  AOI22_X1 U16015 ( .A1(n14701), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n14043), 
        .B2(n14702), .ZN(n14046) );
  NAND2_X1 U16016 ( .A1(n14044), .A2(n14723), .ZN(n14045) );
  OAI211_X1 U16017 ( .C1(n14169), .C2(n14088), .A(n14046), .B(n14045), .ZN(
        n14047) );
  AOI21_X1 U16018 ( .B1(n14171), .B2(n14527), .A(n14047), .ZN(n14048) );
  OAI21_X1 U16019 ( .B1(n14173), .B2(n14701), .A(n14048), .ZN(P1_U3272) );
  OAI211_X1 U16020 ( .C1(n6566), .C2(n14056), .A(n14049), .B(n14716), .ZN(
        n14052) );
  AOI22_X1 U16021 ( .A1(n14050), .A2(n14498), .B1(n14596), .B2(n14081), .ZN(
        n14051) );
  NAND2_X1 U16022 ( .A1(n14052), .A2(n14051), .ZN(n14179) );
  AOI21_X1 U16023 ( .B1(n14053), .B2(n14702), .A(n14179), .ZN(n14063) );
  OAI211_X1 U16024 ( .C1(n14177), .C2(n6650), .A(n14726), .B(n14054), .ZN(
        n14175) );
  NAND2_X1 U16025 ( .A1(n14057), .A2(n14056), .ZN(n14174) );
  NAND3_X1 U16026 ( .A1(n14055), .A2(n14174), .A3(n14527), .ZN(n14060) );
  AOI22_X1 U16027 ( .A1(n14058), .A2(n14723), .B1(n14736), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n14059) );
  OAI211_X1 U16028 ( .C1(n14175), .C2(n14088), .A(n14060), .B(n14059), .ZN(
        n14061) );
  INV_X1 U16029 ( .A(n14061), .ZN(n14062) );
  OAI21_X1 U16030 ( .B1(n14063), .B2(n14701), .A(n14062), .ZN(P1_U3273) );
  XNOR2_X1 U16031 ( .A(n14065), .B(n14064), .ZN(n14068) );
  AOI222_X1 U16032 ( .A1(n14068), .A2(n14716), .B1(n14067), .B2(n14498), .C1(
        n14066), .C2(n14596), .ZN(n14183) );
  AOI211_X1 U16033 ( .C1(n14181), .C2(n14087), .A(n14792), .B(n6650), .ZN(
        n14180) );
  INV_X1 U16034 ( .A(n14069), .ZN(n14070) );
  AOI22_X1 U16035 ( .A1(n14701), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14070), 
        .B2(n14702), .ZN(n14071) );
  OAI21_X1 U16036 ( .B1(n14072), .B2(n14103), .A(n14071), .ZN(n14076) );
  XNOR2_X1 U16037 ( .A(n14073), .B(n14074), .ZN(n14184) );
  NOR2_X1 U16038 ( .A1(n14184), .A2(n14107), .ZN(n14075) );
  AOI211_X1 U16039 ( .C1(n14180), .C2(n14731), .A(n14076), .B(n14075), .ZN(
        n14077) );
  OAI21_X1 U16040 ( .B1(n14736), .B2(n14183), .A(n14077), .ZN(P1_U3274) );
  XNOR2_X1 U16041 ( .A(n14078), .B(n14079), .ZN(n14185) );
  INV_X1 U16042 ( .A(n14185), .ZN(n14095) );
  XNOR2_X1 U16043 ( .A(n14080), .B(n14079), .ZN(n14084) );
  AOI22_X1 U16044 ( .A1(n14081), .A2(n14498), .B1(n14596), .B2(n14497), .ZN(
        n14083) );
  NAND2_X1 U16045 ( .A1(n14185), .A2(n14718), .ZN(n14082) );
  OAI211_X1 U16046 ( .C1(n14084), .C2(n14691), .A(n14083), .B(n14082), .ZN(
        n14190) );
  NAND2_X1 U16047 ( .A1(n14190), .A2(n14721), .ZN(n14093) );
  OAI22_X1 U16048 ( .A1(n14721), .A2(n14086), .B1(n14085), .B2(n14719), .ZN(
        n14090) );
  OAI211_X1 U16049 ( .C1(n14099), .C2(n14188), .A(n14726), .B(n14087), .ZN(
        n14186) );
  NOR2_X1 U16050 ( .A1(n14186), .A2(n14088), .ZN(n14089) );
  AOI211_X1 U16051 ( .C1(n14723), .C2(n14091), .A(n14090), .B(n14089), .ZN(
        n14092) );
  OAI211_X1 U16052 ( .C1(n14095), .C2(n14094), .A(n14093), .B(n14092), .ZN(
        P1_U3275) );
  XNOR2_X1 U16053 ( .A(n14096), .B(n14106), .ZN(n14098) );
  AOI21_X1 U16054 ( .B1(n14098), .B2(n14716), .A(n14097), .ZN(n14194) );
  AOI211_X1 U16055 ( .C1(n14192), .C2(n14506), .A(n14792), .B(n14099), .ZN(
        n14191) );
  INV_X1 U16056 ( .A(n14100), .ZN(n14101) );
  AOI22_X1 U16057 ( .A1(n14701), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n14101), 
        .B2(n14702), .ZN(n14102) );
  OAI21_X1 U16058 ( .B1(n14104), .B2(n14103), .A(n14102), .ZN(n14109) );
  XNOR2_X1 U16059 ( .A(n14105), .B(n14106), .ZN(n14195) );
  NOR2_X1 U16060 ( .A1(n14195), .A2(n14107), .ZN(n14108) );
  AOI211_X1 U16061 ( .C1(n14191), .C2(n14731), .A(n14109), .B(n14108), .ZN(
        n14110) );
  OAI21_X1 U16062 ( .B1(n14736), .B2(n14194), .A(n14110), .ZN(P1_U3276) );
  OAI211_X1 U16063 ( .C1(n14112), .C2(n14122), .A(n14716), .B(n14111), .ZN(
        n14548) );
  INV_X1 U16064 ( .A(n14548), .ZN(n14117) );
  OR2_X1 U16065 ( .A1(n14113), .A2(n14694), .ZN(n14116) );
  NAND2_X1 U16066 ( .A1(n14114), .A2(n14596), .ZN(n14115) );
  NAND2_X1 U16067 ( .A1(n14116), .A2(n14115), .ZN(n14544) );
  OAI21_X1 U16068 ( .B1(n14117), .B2(n14544), .A(n14721), .ZN(n14129) );
  OAI22_X1 U16069 ( .A1(n14721), .A2(n14119), .B1(n14118), .B2(n14719), .ZN(
        n14120) );
  AOI21_X1 U16070 ( .B1(n14545), .B2(n14723), .A(n14120), .ZN(n14128) );
  NAND2_X1 U16071 ( .A1(n14123), .A2(n14122), .ZN(n14546) );
  NAND3_X1 U16072 ( .A1(n14121), .A2(n14546), .A3(n14527), .ZN(n14127) );
  AOI211_X1 U16073 ( .C1(n14545), .C2(n14125), .A(n14792), .B(n11843), .ZN(
        n14543) );
  NAND2_X1 U16074 ( .A1(n14543), .A2(n14731), .ZN(n14126) );
  NAND4_X1 U16075 ( .A1(n14129), .A2(n14128), .A3(n14127), .A4(n14126), .ZN(
        P1_U3279) );
  OAI211_X1 U16076 ( .C1(n14131), .C2(n14781), .A(n14130), .B(n14132), .ZN(
        n14197) );
  MUX2_X1 U16077 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14197), .S(n14811), .Z(
        P1_U3559) );
  OAI211_X1 U16078 ( .C1(n14134), .C2(n14781), .A(n14133), .B(n14132), .ZN(
        n14198) );
  MUX2_X1 U16079 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14198), .S(n14811), .Z(
        P1_U3558) );
  MUX2_X1 U16080 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14135), .S(n14811), .Z(
        P1_U3556) );
  AOI21_X1 U16081 ( .B1(n14137), .B2(n14761), .A(n14136), .ZN(n14138) );
  OAI211_X1 U16082 ( .C1(n14537), .C2(n14140), .A(n14139), .B(n14138), .ZN(
        n14199) );
  MUX2_X1 U16083 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14199), .S(n14811), .Z(
        P1_U3555) );
  OAI21_X1 U16084 ( .B1(n14537), .B2(n14146), .A(n14145), .ZN(n14200) );
  MUX2_X1 U16085 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14200), .S(n14811), .Z(
        P1_U3554) );
  AOI22_X1 U16086 ( .A1(n14148), .A2(n14726), .B1(n14147), .B2(n14761), .ZN(
        n14152) );
  NAND3_X1 U16087 ( .A1(n14150), .A2(n14797), .A3(n14149), .ZN(n14151) );
  NAND3_X1 U16088 ( .A1(n14153), .A2(n14152), .A3(n14151), .ZN(n14201) );
  MUX2_X1 U16089 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14201), .S(n14811), .Z(
        P1_U3553) );
  AOI21_X1 U16090 ( .B1(n14155), .B2(n14761), .A(n14154), .ZN(n14156) );
  OAI211_X1 U16091 ( .C1(n14537), .C2(n14158), .A(n14157), .B(n14156), .ZN(
        n14202) );
  MUX2_X1 U16092 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14202), .S(n14811), .Z(
        P1_U3552) );
  AOI21_X1 U16093 ( .B1(n14160), .B2(n14761), .A(n14159), .ZN(n14161) );
  OAI211_X1 U16094 ( .C1(n14537), .C2(n14163), .A(n14162), .B(n14161), .ZN(
        n14203) );
  MUX2_X1 U16095 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14203), .S(n14811), .Z(
        P1_U3551) );
  AOI21_X1 U16096 ( .B1(n14165), .B2(n14761), .A(n14164), .ZN(n14166) );
  OAI211_X1 U16097 ( .C1(n14537), .C2(n14168), .A(n14167), .B(n14166), .ZN(
        n14204) );
  MUX2_X1 U16098 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14204), .S(n14811), .Z(
        P1_U3550) );
  OAI21_X1 U16099 ( .B1(n6939), .B2(n14781), .A(n14169), .ZN(n14170) );
  AOI21_X1 U16100 ( .B1(n14171), .B2(n14797), .A(n14170), .ZN(n14172) );
  NAND2_X1 U16101 ( .A1(n14173), .A2(n14172), .ZN(n14205) );
  MUX2_X1 U16102 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14205), .S(n14811), .Z(
        P1_U3549) );
  NAND3_X1 U16103 ( .A1(n14055), .A2(n14174), .A3(n14797), .ZN(n14176) );
  OAI211_X1 U16104 ( .C1(n14177), .C2(n14781), .A(n14176), .B(n14175), .ZN(
        n14178) );
  INV_X1 U16105 ( .A(n14811), .ZN(n14809) );
  MUX2_X1 U16106 ( .A(n14206), .B(P1_REG1_REG_20__SCAN_IN), .S(n14809), .Z(
        P1_U3548) );
  AOI21_X1 U16107 ( .B1(n14181), .B2(n14761), .A(n14180), .ZN(n14182) );
  OAI211_X1 U16108 ( .C1(n14537), .C2(n14184), .A(n14183), .B(n14182), .ZN(
        n14207) );
  MUX2_X1 U16109 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14207), .S(n14811), .Z(
        P1_U3547) );
  NAND2_X1 U16110 ( .A1(n14185), .A2(n14787), .ZN(n14187) );
  OAI211_X1 U16111 ( .C1(n14188), .C2(n14781), .A(n14187), .B(n14186), .ZN(
        n14189) );
  OR2_X1 U16112 ( .A1(n14190), .A2(n14189), .ZN(n14208) );
  MUX2_X1 U16113 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14208), .S(n14811), .Z(
        P1_U3546) );
  AOI21_X1 U16114 ( .B1(n14192), .B2(n14761), .A(n14191), .ZN(n14193) );
  OAI211_X1 U16115 ( .C1(n14537), .C2(n14195), .A(n14194), .B(n14193), .ZN(
        n14209) );
  MUX2_X1 U16116 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14209), .S(n14811), .Z(
        P1_U3545) );
  MUX2_X1 U16117 ( .A(n14196), .B(P1_REG1_REG_0__SCAN_IN), .S(n14809), .Z(
        P1_U3528) );
  MUX2_X1 U16118 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14197), .S(n14799), .Z(
        P1_U3527) );
  MUX2_X1 U16119 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14198), .S(n14799), .Z(
        P1_U3526) );
  MUX2_X1 U16120 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14199), .S(n14799), .Z(
        P1_U3523) );
  MUX2_X1 U16121 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14200), .S(n14799), .Z(
        P1_U3522) );
  MUX2_X1 U16122 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14201), .S(n14799), .Z(
        P1_U3521) );
  MUX2_X1 U16123 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14202), .S(n14799), .Z(
        P1_U3520) );
  MUX2_X1 U16124 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14203), .S(n14799), .Z(
        P1_U3519) );
  MUX2_X1 U16125 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14204), .S(n14799), .Z(
        P1_U3518) );
  MUX2_X1 U16126 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14205), .S(n14799), .Z(
        P1_U3517) );
  MUX2_X1 U16127 ( .A(n14206), .B(P1_REG0_REG_20__SCAN_IN), .S(n14798), .Z(
        P1_U3516) );
  MUX2_X1 U16128 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14207), .S(n14799), .Z(
        P1_U3515) );
  MUX2_X1 U16129 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14208), .S(n14799), .Z(
        P1_U3513) );
  MUX2_X1 U16130 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14209), .S(n14799), .Z(
        P1_U3510) );
  NAND2_X1 U16131 ( .A1(n13683), .A2(n14210), .ZN(n14214) );
  NAND2_X1 U16132 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_STATE_REG_SCAN_IN), 
        .ZN(n14211) );
  OR3_X1 U16133 ( .A1(n14212), .A2(P1_IR_REG_30__SCAN_IN), .A3(n14211), .ZN(
        n14213) );
  OAI211_X1 U16134 ( .C1(n14215), .C2(n14216), .A(n14214), .B(n14213), .ZN(
        P1_U3324) );
  OAI222_X1 U16135 ( .A1(n14225), .A2(n14219), .B1(n14218), .B2(P1_U3086), 
        .C1(n14217), .C2(n14216), .ZN(P1_U3325) );
  OAI222_X1 U16136 ( .A1(n14225), .A2(n14221), .B1(n6538), .B2(P1_U3086), .C1(
        n14220), .C2(n14216), .ZN(P1_U3328) );
  OAI222_X1 U16137 ( .A1(n14225), .A2(n14224), .B1(P1_U3086), .B2(n14223), 
        .C1(n14222), .C2(n14216), .ZN(P1_U3329) );
  MUX2_X1 U16138 ( .A(n14227), .B(n14226), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16139 ( .A(n14228), .ZN(n14229) );
  MUX2_X1 U16140 ( .A(n14229), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AND2_X1 U16141 ( .A1(n11779), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n14264) );
  INV_X1 U16142 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14230) );
  NAND2_X1 U16143 ( .A1(n14230), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n14262) );
  INV_X1 U16144 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15172) );
  OR2_X1 U16145 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(n15172), .ZN(n14261) );
  INV_X1 U16146 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14259) );
  INV_X1 U16147 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14257) );
  INV_X1 U16148 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14255) );
  INV_X1 U16149 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n14249) );
  INV_X1 U16150 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15076) );
  AOI22_X1 U16151 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n15076), .B1(
        P3_ADDR_REG_8__SCAN_IN), .B2(n14249), .ZN(n14302) );
  INV_X1 U16152 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14244) );
  XNOR2_X1 U16153 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n14278) );
  NAND2_X1 U16154 ( .A1(n14283), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14282) );
  NAND2_X1 U16155 ( .A1(n14281), .A2(n14280), .ZN(n14231) );
  NAND2_X1 U16156 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14233), .ZN(n14236) );
  INV_X1 U16157 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14234) );
  NAND2_X1 U16158 ( .A1(n14277), .A2(n14234), .ZN(n14235) );
  NAND2_X1 U16159 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14237), .ZN(n14238) );
  INV_X1 U16160 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14639) );
  NAND2_X1 U16161 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14239), .ZN(n14242) );
  INV_X1 U16162 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14240) );
  NAND2_X1 U16163 ( .A1(n14275), .A2(n14240), .ZN(n14241) );
  INV_X1 U16164 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n15039) );
  NAND2_X1 U16165 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n15039), .ZN(n14243) );
  INV_X1 U16166 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n15058) );
  NAND2_X1 U16167 ( .A1(n14245), .A2(n15058), .ZN(n14247) );
  XNOR2_X1 U16168 ( .A(n14245), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n14298) );
  NAND2_X1 U16169 ( .A1(n14298), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n14246) );
  NAND2_X1 U16170 ( .A1(n14247), .A2(n14246), .ZN(n14303) );
  NAND2_X1 U16171 ( .A1(n14302), .A2(n14303), .ZN(n14248) );
  XOR2_X1 U16172 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(P3_ADDR_REG_9__SCAN_IN), .Z(
        n14273) );
  NAND2_X1 U16173 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14252), .ZN(n14312) );
  XNOR2_X1 U16174 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n14271) );
  NAND2_X1 U16175 ( .A1(n14272), .A2(n14271), .ZN(n14254) );
  XOR2_X1 U16176 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .Z(n14269) );
  AND2_X1 U16177 ( .A1(n14259), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n14258) );
  OAI22_X1 U16178 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14259), .B1(n14315), 
        .B2(n14258), .ZN(n14260) );
  INV_X1 U16179 ( .A(n14260), .ZN(n14317) );
  AOI22_X1 U16180 ( .A1(n14261), .A2(n14317), .B1(n15172), .B2(
        P1_ADDR_REG_14__SCAN_IN), .ZN(n14268) );
  INV_X1 U16181 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14654) );
  AOI22_X1 U16182 ( .A1(n14262), .A2(n14268), .B1(n14654), .B2(
        P3_ADDR_REG_15__SCAN_IN), .ZN(n14265) );
  INV_X1 U16183 ( .A(n14265), .ZN(n14263) );
  OAI22_X1 U16184 ( .A1(n14264), .A2(n14263), .B1(P3_ADDR_REG_16__SCAN_IN), 
        .B2(n11779), .ZN(n14322) );
  XNOR2_X1 U16185 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14322), .ZN(n14323) );
  XNOR2_X1 U16186 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14323), .ZN(n14366) );
  XNOR2_X1 U16187 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n14266) );
  XNOR2_X1 U16188 ( .A(n14266), .B(n14265), .ZN(n14590) );
  XOR2_X1 U16189 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .Z(n14267) );
  XOR2_X1 U16190 ( .A(n14268), .B(n14267), .Z(n14319) );
  XOR2_X1 U16191 ( .A(n14270), .B(n14269), .Z(n14572) );
  XNOR2_X1 U16192 ( .A(n14272), .B(n14271), .ZN(n14569) );
  XOR2_X1 U16193 ( .A(n14274), .B(n14273), .Z(n14307) );
  XNOR2_X1 U16194 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n14275), .ZN(n14291) );
  XNOR2_X1 U16195 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n14276), .ZN(n14289) );
  NAND2_X1 U16196 ( .A1(n14289), .A2(n14876), .ZN(n14290) );
  XNOR2_X1 U16197 ( .A(n14277), .B(P1_ADDR_REG_3__SCAN_IN), .ZN(n15344) );
  XOR2_X1 U16198 ( .A(n14279), .B(n14278), .Z(n14343) );
  INV_X1 U16199 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n14285) );
  NOR2_X1 U16200 ( .A1(n14284), .A2(n14285), .ZN(n14286) );
  OAI21_X1 U16201 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n14283), .A(n14282), .ZN(
        n15338) );
  NAND2_X1 U16202 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15338), .ZN(n15348) );
  NOR2_X1 U16203 ( .A1(n15348), .A2(n15347), .ZN(n15346) );
  NOR2_X1 U16204 ( .A1(n14343), .A2(n14342), .ZN(n14287) );
  NAND2_X1 U16205 ( .A1(n14343), .A2(n14342), .ZN(n14341) );
  NAND2_X1 U16206 ( .A1(n15344), .A2(n15343), .ZN(n14288) );
  NOR2_X1 U16207 ( .A1(n15344), .A2(n15343), .ZN(n15342) );
  XNOR2_X1 U16208 ( .A(P2_ADDR_REG_4__SCAN_IN), .B(n14289), .ZN(n15333) );
  NAND2_X1 U16209 ( .A1(n15334), .A2(n15333), .ZN(n15332) );
  NAND2_X1 U16210 ( .A1(n14291), .A2(n14292), .ZN(n14293) );
  INV_X1 U16211 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15336) );
  INV_X1 U16212 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n14889) );
  NOR2_X1 U16213 ( .A1(n14294), .A2(n14889), .ZN(n14297) );
  XOR2_X1 U16214 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), .Z(
        n14295) );
  XNOR2_X1 U16215 ( .A(n14296), .B(n14295), .ZN(n14346) );
  INV_X1 U16216 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n14300) );
  NOR2_X1 U16217 ( .A1(n14299), .A2(n14300), .ZN(n14301) );
  XNOR2_X1 U16218 ( .A(n14298), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15341) );
  XNOR2_X1 U16219 ( .A(n14303), .B(n14302), .ZN(n14305) );
  NAND2_X1 U16220 ( .A1(n14304), .A2(n14305), .ZN(n14306) );
  INV_X1 U16221 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14904) );
  NOR2_X1 U16222 ( .A1(n14307), .A2(n14308), .ZN(n14309) );
  INV_X1 U16223 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14352) );
  INV_X1 U16224 ( .A(n14310), .ZN(n14311) );
  NAND2_X1 U16225 ( .A1(n14312), .A2(n14311), .ZN(n14313) );
  XNOR2_X1 U16226 ( .A(n14313), .B(P3_ADDR_REG_10__SCAN_IN), .ZN(n14354) );
  NAND2_X1 U16227 ( .A1(n14355), .A2(n14354), .ZN(n14353) );
  XOR2_X1 U16228 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .Z(n14314) );
  XOR2_X1 U16229 ( .A(n14315), .B(n14314), .Z(n14576) );
  NAND2_X1 U16230 ( .A1(n14577), .A2(n14576), .ZN(n14316) );
  XNOR2_X1 U16231 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n14318) );
  XNOR2_X1 U16232 ( .A(n14318), .B(n14317), .ZN(n14581) );
  INV_X1 U16233 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n14587) );
  NAND2_X1 U16234 ( .A1(n14320), .A2(n14319), .ZN(n14586) );
  NAND2_X1 U16235 ( .A1(n14366), .A2(n14365), .ZN(n14321) );
  XNOR2_X1 U16236 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n14327) );
  NOR2_X1 U16237 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14322), .ZN(n14326) );
  NOR2_X1 U16238 ( .A1(n14324), .A2(n14323), .ZN(n14325) );
  NOR2_X1 U16239 ( .A1(n14326), .A2(n14325), .ZN(n14330) );
  XNOR2_X1 U16240 ( .A(n14327), .B(n14330), .ZN(n14337) );
  INV_X1 U16241 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n14328) );
  OR2_X1 U16242 ( .A1(n14328), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n14329) );
  AOI22_X1 U16243 ( .A1(n14330), .A2(n14329), .B1(P1_ADDR_REG_18__SCAN_IN), 
        .B2(n14328), .ZN(n14331) );
  XNOR2_X1 U16244 ( .A(n14332), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n14333) );
  XNOR2_X1 U16245 ( .A(n14333), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n14334) );
  OAI21_X1 U16246 ( .B1(n14337), .B2(n14336), .A(n14335), .ZN(n14338) );
  XNOR2_X1 U16247 ( .A(n14338), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16248 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14339) );
  OAI21_X1 U16249 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14339), 
        .ZN(U28) );
  AOI21_X1 U16250 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14340) );
  OAI21_X1 U16251 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14340), 
        .ZN(U29) );
  OAI21_X1 U16252 ( .B1(n14343), .B2(n14342), .A(n14341), .ZN(n14344) );
  XNOR2_X1 U16253 ( .A(n14344), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  AOI21_X1 U16254 ( .B1(n14347), .B2(n14346), .A(n14345), .ZN(SUB_1596_U57) );
  OAI21_X1 U16255 ( .B1(n14349), .B2(n14904), .A(n14348), .ZN(SUB_1596_U55) );
  AOI21_X1 U16256 ( .B1(n14352), .B2(n14351), .A(n14350), .ZN(SUB_1596_U54) );
  OAI21_X1 U16257 ( .B1(n14355), .B2(n14354), .A(n14353), .ZN(n14356) );
  XNOR2_X1 U16258 ( .A(n14356), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  OAI211_X1 U16259 ( .C1(n14359), .C2(n14781), .A(n14358), .B(n14357), .ZN(
        n14360) );
  AOI21_X1 U16260 ( .B1(n14361), .B2(n14797), .A(n14360), .ZN(n14363) );
  AOI22_X1 U16261 ( .A1(n14799), .A2(n14363), .B1(n14362), .B2(n14798), .ZN(
        P1_U3495) );
  AOI22_X1 U16262 ( .A1(n14811), .A2(n14363), .B1(n10831), .B2(n14809), .ZN(
        P1_U3540) );
  AOI21_X1 U16263 ( .B1(n14366), .B2(n14365), .A(n14364), .ZN(n14367) );
  XOR2_X1 U16264 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n14367), .Z(SUB_1596_U63)
         );
  XOR2_X1 U16265 ( .A(n6717), .B(n14368), .Z(n14377) );
  NAND2_X1 U16266 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(P3_U3151), .ZN(n15171)
         );
  NAND2_X1 U16267 ( .A1(n14371), .A2(n14370), .ZN(n14372) );
  OAI211_X1 U16268 ( .C1(n14374), .C2(n14373), .A(n15171), .B(n14372), .ZN(
        n14375) );
  AOI21_X1 U16269 ( .B1(n14377), .B2(n14376), .A(n14375), .ZN(n14378) );
  OAI21_X1 U16270 ( .B1(n14380), .B2(n14379), .A(n14378), .ZN(P3_U3155) );
  AOI21_X1 U16271 ( .B1(n14383), .B2(n14382), .A(n14381), .ZN(n14398) );
  OAI21_X1 U16272 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n14385), .A(n14384), 
        .ZN(n14391) );
  NOR2_X1 U16273 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14386), .ZN(n14387) );
  AOI21_X1 U16274 ( .B1(n15149), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n14387), 
        .ZN(n14388) );
  OAI21_X1 U16275 ( .B1(n15170), .B2(n14389), .A(n14388), .ZN(n14390) );
  AOI21_X1 U16276 ( .B1(n14391), .B2(n15176), .A(n14390), .ZN(n14397) );
  AOI21_X1 U16277 ( .B1(n14394), .B2(n14393), .A(n14392), .ZN(n14395) );
  OR2_X1 U16278 ( .A1(n14395), .A2(n15158), .ZN(n14396) );
  OAI211_X1 U16279 ( .C1(n14398), .C2(n15184), .A(n14397), .B(n14396), .ZN(
        P3_U3197) );
  INV_X1 U16280 ( .A(n15170), .ZN(n14432) );
  AOI22_X1 U16281 ( .A1(n14432), .A2(n14399), .B1(n15149), .B2(
        P3_ADDR_REG_16__SCAN_IN), .ZN(n14415) );
  INV_X1 U16282 ( .A(n14400), .ZN(n14401) );
  NAND2_X1 U16283 ( .A1(n14402), .A2(n14401), .ZN(n14403) );
  XNOR2_X1 U16284 ( .A(n14404), .B(n14403), .ZN(n14408) );
  XNOR2_X1 U16285 ( .A(n14406), .B(n14405), .ZN(n14407) );
  AOI22_X1 U16286 ( .A1(n14408), .A2(n15178), .B1(n15176), .B2(n14407), .ZN(
        n14414) );
  NAND2_X1 U16287 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P3_U3151), .ZN(n14413)
         );
  OAI221_X1 U16288 ( .B1(n14411), .B2(n14410), .C1(n14411), .C2(n14409), .A(
        n15054), .ZN(n14412) );
  NAND4_X1 U16289 ( .A1(n14415), .A2(n14414), .A3(n14413), .A4(n14412), .ZN(
        P3_U3198) );
  AOI22_X1 U16290 ( .A1(n14432), .A2(n14416), .B1(n15149), .B2(
        P3_ADDR_REG_17__SCAN_IN), .ZN(n14430) );
  OAI21_X1 U16291 ( .B1(P3_REG1_REG_17__SCAN_IN), .B2(n14418), .A(n14417), 
        .ZN(n14423) );
  AOI211_X1 U16292 ( .C1(n14421), .C2(n14420), .A(n14419), .B(n15158), .ZN(
        n14422) );
  AOI21_X1 U16293 ( .B1(n15176), .B2(n14423), .A(n14422), .ZN(n14429) );
  NAND2_X1 U16294 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(P3_U3151), .ZN(n14428)
         );
  OAI221_X1 U16295 ( .B1(n14426), .B2(n14425), .C1(n14426), .C2(n14424), .A(
        n15054), .ZN(n14427) );
  NAND4_X1 U16296 ( .A1(n14430), .A2(n14429), .A3(n14428), .A4(n14427), .ZN(
        P3_U3199) );
  AOI22_X1 U16297 ( .A1(n14432), .A2(n14431), .B1(n15149), .B2(
        P3_ADDR_REG_18__SCAN_IN), .ZN(n14447) );
  XNOR2_X1 U16298 ( .A(n14434), .B(n14433), .ZN(n14440) );
  AOI21_X1 U16299 ( .B1(n14437), .B2(n14436), .A(n14435), .ZN(n14438) );
  NOR2_X1 U16300 ( .A1(n14438), .A2(n15158), .ZN(n14439) );
  AOI21_X1 U16301 ( .B1(n14440), .B2(n15176), .A(n14439), .ZN(n14446) );
  NAND2_X1 U16302 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(P3_U3151), .ZN(n14445)
         );
  OAI221_X1 U16303 ( .B1(n14443), .B2(n14442), .C1(n14443), .C2(n14441), .A(
        n15054), .ZN(n14444) );
  NAND4_X1 U16304 ( .A1(n14447), .A2(n14446), .A3(n14445), .A4(n14444), .ZN(
        P3_U3200) );
  XNOR2_X1 U16305 ( .A(n14449), .B(n14448), .ZN(n14470) );
  XNOR2_X1 U16306 ( .A(n14450), .B(n14451), .ZN(n14452) );
  OAI222_X1 U16307 ( .A1(n15241), .A2(n14454), .B1(n15243), .B2(n14453), .C1(
        n14452), .C2(n15249), .ZN(n14468) );
  AOI21_X1 U16308 ( .B1(n14470), .B2(n15209), .A(n14468), .ZN(n14459) );
  NOR2_X1 U16309 ( .A1(n14455), .A2(n15253), .ZN(n14469) );
  INV_X1 U16310 ( .A(n14456), .ZN(n14457) );
  AOI22_X1 U16311 ( .A1(n15227), .A2(n14469), .B1(n15226), .B2(n14457), .ZN(
        n14458) );
  OAI221_X1 U16312 ( .B1(n12719), .B2(n14459), .C1(n15273), .C2(n8366), .A(
        n14458), .ZN(P3_U3222) );
  AOI211_X1 U16313 ( .C1(n14462), .C2(n15293), .A(n14461), .B(n14460), .ZN(
        n14473) );
  AOI22_X1 U16314 ( .A1(n15331), .A2(n14473), .B1(n8418), .B2(n15329), .ZN(
        P3_U3472) );
  INV_X1 U16315 ( .A(n14463), .ZN(n14466) );
  INV_X1 U16316 ( .A(n14464), .ZN(n14465) );
  AOI211_X1 U16317 ( .C1(n14467), .C2(n15293), .A(n14466), .B(n14465), .ZN(
        n14475) );
  AOI22_X1 U16318 ( .A1(n15331), .A2(n14475), .B1(n12588), .B2(n15329), .ZN(
        P3_U3471) );
  AOI211_X1 U16319 ( .C1(n14470), .C2(n15293), .A(n14469), .B(n14468), .ZN(
        n14477) );
  INV_X1 U16320 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14471) );
  AOI22_X1 U16321 ( .A1(n15331), .A2(n14477), .B1(n14471), .B2(n15329), .ZN(
        P3_U3470) );
  INV_X1 U16322 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14472) );
  AOI22_X1 U16323 ( .A1(n15318), .A2(n14473), .B1(n14472), .B2(n15316), .ZN(
        P3_U3429) );
  INV_X1 U16324 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14474) );
  AOI22_X1 U16325 ( .A1(n15318), .A2(n14475), .B1(n14474), .B2(n15316), .ZN(
        P3_U3426) );
  INV_X1 U16326 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14476) );
  AOI22_X1 U16327 ( .A1(n15318), .A2(n14477), .B1(n14476), .B2(n15316), .ZN(
        P3_U3423) );
  NAND2_X1 U16328 ( .A1(n14478), .A2(n14761), .ZN(n14790) );
  INV_X1 U16329 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n14479) );
  OAI22_X1 U16330 ( .A1(n14790), .A2(n14480), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14479), .ZN(n14481) );
  INV_X1 U16331 ( .A(n14481), .ZN(n14491) );
  XNOR2_X1 U16332 ( .A(n14484), .B(n14483), .ZN(n14485) );
  XNOR2_X1 U16333 ( .A(n14482), .B(n14485), .ZN(n14489) );
  NAND2_X1 U16334 ( .A1(n14487), .A2(n14486), .ZN(n14789) );
  AOI22_X1 U16335 ( .A1(n14489), .A2(n14488), .B1(n14601), .B2(n14789), .ZN(
        n14490) );
  OAI211_X1 U16336 ( .C1(n14492), .C2(n14606), .A(n14491), .B(n14490), .ZN(
        P1_U3217) );
  NAND2_X1 U16337 ( .A1(n14493), .A2(n14503), .ZN(n14494) );
  NAND2_X1 U16338 ( .A1(n14495), .A2(n14494), .ZN(n14496) );
  NAND2_X1 U16339 ( .A1(n14496), .A2(n14716), .ZN(n14501) );
  AOI22_X1 U16340 ( .A1(n14499), .A2(n14596), .B1(n14498), .B2(n14497), .ZN(
        n14500) );
  NAND2_X1 U16341 ( .A1(n14501), .A2(n14500), .ZN(n14536) );
  XNOR2_X1 U16342 ( .A(n14502), .B(n14503), .ZN(n14530) );
  AND2_X1 U16343 ( .A1(n14530), .A2(n14504), .ZN(n14513) );
  AOI21_X1 U16344 ( .B1(n14505), .B2(n14531), .A(n14792), .ZN(n14507) );
  NAND2_X1 U16345 ( .A1(n14507), .A2(n14506), .ZN(n14532) );
  AOI22_X1 U16346 ( .A1(n14531), .A2(n14509), .B1(n14508), .B2(n14702), .ZN(
        n14510) );
  OAI21_X1 U16347 ( .B1(n14532), .B2(n14511), .A(n14510), .ZN(n14512) );
  AOI22_X1 U16348 ( .A1(n14736), .A2(n11795), .B1(n7497), .B2(n14721), .ZN(
        P1_U3277) );
  INV_X1 U16349 ( .A(n14514), .ZN(n14515) );
  AOI21_X1 U16350 ( .B1(n14515), .B2(n14523), .A(n14691), .ZN(n14518) );
  AOI21_X1 U16351 ( .B1(n14518), .B2(n14517), .A(n14516), .ZN(n14557) );
  INV_X1 U16352 ( .A(n14519), .ZN(n14520) );
  AOI222_X1 U16353 ( .A1(n14521), .A2(n14723), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n14701), .C1(n14520), .C2(n14702), .ZN(n14529) );
  XNOR2_X1 U16354 ( .A(n14522), .B(n14523), .ZN(n14560) );
  OAI211_X1 U16355 ( .C1(n14558), .C2(n14525), .A(n14726), .B(n14524), .ZN(
        n14556) );
  INV_X1 U16356 ( .A(n14556), .ZN(n14526) );
  AOI22_X1 U16357 ( .A1(n14560), .A2(n14527), .B1(n14731), .B2(n14526), .ZN(
        n14528) );
  OAI211_X1 U16358 ( .C1(n14701), .C2(n14557), .A(n14529), .B(n14528), .ZN(
        P1_U3282) );
  AND2_X1 U16359 ( .A1(n14530), .A2(n14797), .ZN(n14535) );
  INV_X1 U16360 ( .A(n14531), .ZN(n14533) );
  OAI21_X1 U16361 ( .B1(n14533), .B2(n14781), .A(n14532), .ZN(n14534) );
  AOI22_X1 U16362 ( .A1(n14811), .A2(n7496), .B1(n11784), .B2(n14809), .ZN(
        P1_U3544) );
  NOR2_X1 U16363 ( .A1(n14538), .A2(n14537), .ZN(n14542) );
  NOR4_X1 U16364 ( .A1(n14542), .A2(n14541), .A3(n14540), .A4(n14539), .ZN(
        n14561) );
  AOI22_X1 U16365 ( .A1(n14811), .A2(n14561), .B1(n7875), .B2(n14809), .ZN(
        P1_U3543) );
  AOI211_X1 U16366 ( .C1(n14545), .C2(n14761), .A(n14544), .B(n14543), .ZN(
        n14549) );
  NAND3_X1 U16367 ( .A1(n14121), .A2(n14546), .A3(n14797), .ZN(n14547) );
  AOI22_X1 U16368 ( .A1(n14811), .A2(n14563), .B1(n11373), .B2(n14809), .ZN(
        P1_U3542) );
  AND2_X1 U16369 ( .A1(n14550), .A2(n14797), .ZN(n14554) );
  OAI21_X1 U16370 ( .B1(n14552), .B2(n14781), .A(n14551), .ZN(n14553) );
  NOR3_X1 U16371 ( .A1(n14555), .A2(n14554), .A3(n14553), .ZN(n14564) );
  AOI22_X1 U16372 ( .A1(n14811), .A2(n14564), .B1(n11231), .B2(n14809), .ZN(
        P1_U3541) );
  OAI211_X1 U16373 ( .C1(n14558), .C2(n14781), .A(n14557), .B(n14556), .ZN(
        n14559) );
  AOI21_X1 U16374 ( .B1(n14797), .B2(n14560), .A(n14559), .ZN(n14566) );
  AOI22_X1 U16375 ( .A1(n14811), .A2(n14566), .B1(n10587), .B2(n14809), .ZN(
        P1_U3539) );
  AOI22_X1 U16376 ( .A1(n14799), .A2(n7496), .B1(n7892), .B2(n14798), .ZN(
        P1_U3507) );
  AOI22_X1 U16377 ( .A1(n14799), .A2(n14561), .B1(n7877), .B2(n14798), .ZN(
        P1_U3504) );
  INV_X1 U16378 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14562) );
  AOI22_X1 U16379 ( .A1(n14799), .A2(n14563), .B1(n14562), .B2(n14798), .ZN(
        P1_U3501) );
  AOI22_X1 U16380 ( .A1(n14799), .A2(n14564), .B1(n7844), .B2(n14798), .ZN(
        P1_U3498) );
  INV_X1 U16381 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14565) );
  AOI22_X1 U16382 ( .A1(n14799), .A2(n14566), .B1(n14565), .B2(n14798), .ZN(
        P1_U3492) );
  OAI21_X1 U16383 ( .B1(n14569), .B2(n14568), .A(n14567), .ZN(n14570) );
  XNOR2_X1 U16384 ( .A(n14570), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  OAI21_X1 U16385 ( .B1(n14573), .B2(n14572), .A(n14571), .ZN(n14574) );
  XNOR2_X1 U16386 ( .A(n14574), .B(P2_ADDR_REG_12__SCAN_IN), .ZN(SUB_1596_U68)
         );
  AOI21_X1 U16387 ( .B1(n14577), .B2(n14576), .A(n14575), .ZN(n14578) );
  XOR2_X1 U16388 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n14578), .Z(SUB_1596_U67)
         );
  OAI21_X1 U16389 ( .B1(n14581), .B2(n14580), .A(n14579), .ZN(n14582) );
  XNOR2_X1 U16390 ( .A(n14582), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  OAI222_X1 U16391 ( .A1(n14587), .A2(n14586), .B1(n14587), .B2(n14585), .C1(
        n14584), .C2(n14583), .ZN(SUB_1596_U65) );
  OAI21_X1 U16392 ( .B1(n14590), .B2(n14589), .A(n14588), .ZN(n14591) );
  XNOR2_X1 U16393 ( .A(n14591), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  AND2_X1 U16394 ( .A1(n14724), .A2(n14761), .ZN(n14740) );
  AOI22_X1 U16395 ( .A1(n14592), .A2(n14740), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14605) );
  AOI21_X1 U16396 ( .B1(n14595), .B2(n14594), .A(n14593), .ZN(n14603) );
  NAND2_X1 U16397 ( .A1(n12090), .A2(n14596), .ZN(n14600) );
  NAND2_X1 U16398 ( .A1(n14598), .A2(n14597), .ZN(n14599) );
  NAND2_X1 U16399 ( .A1(n14600), .A2(n14599), .ZN(n14741) );
  AOI22_X1 U16400 ( .A1(n14603), .A2(n14602), .B1(n14601), .B2(n14741), .ZN(
        n14604) );
  OAI211_X1 U16401 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n14606), .A(n14605), .B(
        n14604), .ZN(P1_U3218) );
  INV_X1 U16402 ( .A(n14607), .ZN(n14614) );
  NAND2_X1 U16403 ( .A1(n6538), .A2(n14608), .ZN(n14612) );
  NAND2_X1 U16404 ( .A1(n14610), .A2(n14612), .ZN(n14611) );
  MUX2_X1 U16405 ( .A(n14612), .B(n14611), .S(P1_IR_REG_0__SCAN_IN), .Z(n14613) );
  NAND2_X1 U16406 ( .A1(n14614), .A2(n14613), .ZN(n14617) );
  AOI22_X1 U16407 ( .A1(n14615), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14616) );
  OAI21_X1 U16408 ( .B1(n14618), .B2(n14617), .A(n14616), .ZN(P1_U3243) );
  INV_X1 U16409 ( .A(n14619), .ZN(n14625) );
  MUX2_X1 U16410 ( .A(n9981), .B(P1_REG2_REG_4__SCAN_IN), .S(n14620), .Z(
        n14623) );
  NAND3_X1 U16411 ( .A1(n14623), .A2(n14622), .A3(n14621), .ZN(n14624) );
  NAND3_X1 U16412 ( .A1(n14649), .A2(n14625), .A3(n14624), .ZN(n14633) );
  INV_X1 U16413 ( .A(n14626), .ZN(n14631) );
  NAND3_X1 U16414 ( .A1(n6885), .A2(n14629), .A3(n14628), .ZN(n14630) );
  NAND3_X1 U16415 ( .A1(n14648), .A2(n14631), .A3(n14630), .ZN(n14632) );
  OAI211_X1 U16416 ( .C1(n14634), .C2(n6884), .A(n14633), .B(n14632), .ZN(
        n14635) );
  NOR2_X1 U16417 ( .A1(n14636), .A2(n14635), .ZN(n14638) );
  OAI211_X1 U16418 ( .C1(n14653), .C2(n14639), .A(n14638), .B(n14637), .ZN(
        P1_U3247) );
  AOI21_X1 U16419 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14641), .A(n14640), 
        .ZN(n14642) );
  INV_X1 U16420 ( .A(n14642), .ZN(n14650) );
  OAI21_X1 U16421 ( .B1(n14644), .B2(n7875), .A(n14643), .ZN(n14647) );
  AOI222_X1 U16422 ( .A1(n14650), .A2(n14649), .B1(n14648), .B2(n14647), .C1(
        n14646), .C2(n14645), .ZN(n14652) );
  OAI211_X1 U16423 ( .C1(n14654), .C2(n14653), .A(n14652), .B(n14651), .ZN(
        P1_U3258) );
  OAI21_X1 U16424 ( .B1(n14656), .B2(n14659), .A(n14655), .ZN(n14663) );
  INV_X1 U16425 ( .A(n14657), .ZN(n14662) );
  XNOR2_X1 U16426 ( .A(n14658), .B(n14659), .ZN(n14666) );
  NOR2_X1 U16427 ( .A1(n14666), .A2(n14660), .ZN(n14661) );
  AOI211_X1 U16428 ( .C1(n14716), .C2(n14663), .A(n14662), .B(n14661), .ZN(
        n14783) );
  AOI222_X1 U16429 ( .A1(n14665), .A2(n14723), .B1(n14664), .B2(n14702), .C1(
        P1_REG2_REG_9__SCAN_IN), .C2(n14701), .ZN(n14672) );
  INV_X1 U16430 ( .A(n14666), .ZN(n14786) );
  INV_X1 U16431 ( .A(n14667), .ZN(n14669) );
  OAI211_X1 U16432 ( .C1(n14669), .C2(n14782), .A(n14726), .B(n14668), .ZN(
        n14780) );
  INV_X1 U16433 ( .A(n14780), .ZN(n14670) );
  AOI22_X1 U16434 ( .A1(n14786), .A2(n14732), .B1(n14731), .B2(n14670), .ZN(
        n14671) );
  OAI211_X1 U16435 ( .C1(n14701), .C2(n14783), .A(n14672), .B(n14671), .ZN(
        P1_U3284) );
  XNOR2_X1 U16436 ( .A(n14673), .B(n14674), .ZN(n14773) );
  XNOR2_X1 U16437 ( .A(n14675), .B(n14674), .ZN(n14676) );
  NOR2_X1 U16438 ( .A1(n14676), .A2(n14691), .ZN(n14677) );
  AOI211_X1 U16439 ( .C1(n14773), .C2(n14718), .A(n14678), .B(n14677), .ZN(
        n14770) );
  INV_X1 U16440 ( .A(n14679), .ZN(n14680) );
  AOI222_X1 U16441 ( .A1(n14681), .A2(n14723), .B1(n14680), .B2(n14702), .C1(
        P1_REG2_REG_7__SCAN_IN), .C2(n14701), .ZN(n14687) );
  INV_X1 U16442 ( .A(n14682), .ZN(n14683) );
  OAI211_X1 U16443 ( .C1(n14769), .C2(n14684), .A(n14683), .B(n14726), .ZN(
        n14768) );
  INV_X1 U16444 ( .A(n14768), .ZN(n14685) );
  AOI22_X1 U16445 ( .A1(n14773), .A2(n14732), .B1(n14731), .B2(n14685), .ZN(
        n14686) );
  OAI211_X1 U16446 ( .C1(n14701), .C2(n14770), .A(n14687), .B(n14686), .ZN(
        P1_U3286) );
  XNOR2_X1 U16447 ( .A(n14688), .B(n14689), .ZN(n14758) );
  NAND2_X1 U16448 ( .A1(n14690), .A2(n14689), .ZN(n14692) );
  AOI21_X1 U16449 ( .B1(n14693), .B2(n14692), .A(n14691), .ZN(n14699) );
  OAI22_X1 U16450 ( .A1(n14697), .A2(n14696), .B1(n14695), .B2(n14694), .ZN(
        n14698) );
  AOI211_X1 U16451 ( .C1(n14758), .C2(n14718), .A(n14699), .B(n14698), .ZN(
        n14755) );
  INV_X1 U16452 ( .A(n14700), .ZN(n14703) );
  AOI222_X1 U16453 ( .A1(n14704), .A2(n14723), .B1(n14703), .B2(n14702), .C1(
        P1_REG2_REG_5__SCAN_IN), .C2(n14701), .ZN(n14710) );
  INV_X1 U16454 ( .A(n14705), .ZN(n14707) );
  OAI211_X1 U16455 ( .C1(n14707), .C2(n14754), .A(n14726), .B(n14706), .ZN(
        n14753) );
  INV_X1 U16456 ( .A(n14753), .ZN(n14708) );
  AOI22_X1 U16457 ( .A1(n14758), .A2(n14732), .B1(n14731), .B2(n14708), .ZN(
        n14709) );
  OAI211_X1 U16458 ( .C1(n14701), .C2(n14755), .A(n14710), .B(n14709), .ZN(
        P1_U3288) );
  OAI21_X1 U16459 ( .B1(n14713), .B2(n14712), .A(n14711), .ZN(n14746) );
  XNOR2_X1 U16460 ( .A(n14715), .B(n14714), .ZN(n14717) );
  AND2_X1 U16461 ( .A1(n14717), .A2(n14716), .ZN(n14744) );
  AOI211_X1 U16462 ( .C1(n14718), .C2(n14746), .A(n14741), .B(n14744), .ZN(
        n14735) );
  OAI22_X1 U16463 ( .A1(n14721), .A2(n14720), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14719), .ZN(n14722) );
  AOI21_X1 U16464 ( .B1(n14723), .B2(n14724), .A(n14722), .ZN(n14734) );
  NAND2_X1 U16465 ( .A1(n14725), .A2(n14724), .ZN(n14727) );
  NAND2_X1 U16466 ( .A1(n14727), .A2(n14726), .ZN(n14729) );
  OR2_X1 U16467 ( .A1(n14729), .A2(n14728), .ZN(n14743) );
  INV_X1 U16468 ( .A(n14743), .ZN(n14730) );
  AOI22_X1 U16469 ( .A1(n14746), .A2(n14732), .B1(n14731), .B2(n14730), .ZN(
        n14733) );
  OAI211_X1 U16470 ( .C1(n14736), .C2(n14735), .A(n14734), .B(n14733), .ZN(
        P1_U3290) );
  AND2_X1 U16471 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14739), .ZN(P1_U3294) );
  AND2_X1 U16472 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14739), .ZN(P1_U3295) );
  AND2_X1 U16473 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14739), .ZN(P1_U3296) );
  AND2_X1 U16474 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14739), .ZN(P1_U3297) );
  AND2_X1 U16475 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14739), .ZN(P1_U3298) );
  AND2_X1 U16476 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14739), .ZN(P1_U3299) );
  AND2_X1 U16477 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14739), .ZN(P1_U3300) );
  AND2_X1 U16478 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14739), .ZN(P1_U3301) );
  AND2_X1 U16479 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14739), .ZN(P1_U3302) );
  AND2_X1 U16480 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14739), .ZN(P1_U3303) );
  AND2_X1 U16481 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14739), .ZN(P1_U3304) );
  AND2_X1 U16482 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14739), .ZN(P1_U3305) );
  AND2_X1 U16483 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14739), .ZN(P1_U3306) );
  AND2_X1 U16484 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14739), .ZN(P1_U3307) );
  AND2_X1 U16485 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14739), .ZN(P1_U3308) );
  AND2_X1 U16486 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14739), .ZN(P1_U3309) );
  AND2_X1 U16487 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14739), .ZN(P1_U3310) );
  AND2_X1 U16488 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n6674), .ZN(P1_U3311) );
  AND2_X1 U16489 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n6674), .ZN(P1_U3312) );
  AND2_X1 U16490 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n6674), .ZN(P1_U3313) );
  AND2_X1 U16491 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n6674), .ZN(P1_U3314) );
  INV_X1 U16492 ( .A(n6674), .ZN(n14738) );
  NOR2_X1 U16493 ( .A1(n14738), .A2(n14737), .ZN(P1_U3315) );
  AND2_X1 U16494 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n6674), .ZN(P1_U3316) );
  AND2_X1 U16495 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n6674), .ZN(P1_U3317) );
  AND2_X1 U16496 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n6674), .ZN(P1_U3318) );
  AND2_X1 U16497 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n6674), .ZN(P1_U3319) );
  AND2_X1 U16498 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n6674), .ZN(P1_U3320) );
  AND2_X1 U16499 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n6674), .ZN(P1_U3321) );
  AND2_X1 U16500 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n6674), .ZN(P1_U3322) );
  AND2_X1 U16501 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n6674), .ZN(P1_U3323) );
  NOR2_X1 U16502 ( .A1(n14741), .A2(n14740), .ZN(n14742) );
  NAND2_X1 U16503 ( .A1(n14743), .A2(n14742), .ZN(n14745) );
  AOI211_X1 U16504 ( .C1(n14797), .C2(n14746), .A(n14745), .B(n14744), .ZN(
        n14800) );
  INV_X1 U16505 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14747) );
  AOI22_X1 U16506 ( .A1(n14799), .A2(n14800), .B1(n14747), .B2(n14798), .ZN(
        P1_U3468) );
  OAI21_X1 U16507 ( .B1(n14749), .B2(n14781), .A(n14748), .ZN(n14751) );
  AOI211_X1 U16508 ( .C1(n14752), .C2(n14797), .A(n14751), .B(n14750), .ZN(
        n14802) );
  AOI22_X1 U16509 ( .A1(n14799), .A2(n14802), .B1(n7692), .B2(n14798), .ZN(
        P1_U3471) );
  OAI21_X1 U16510 ( .B1(n14754), .B2(n14781), .A(n14753), .ZN(n14757) );
  INV_X1 U16511 ( .A(n14755), .ZN(n14756) );
  AOI211_X1 U16512 ( .C1(n14787), .C2(n14758), .A(n14757), .B(n14756), .ZN(
        n14803) );
  INV_X1 U16513 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14759) );
  AOI22_X1 U16514 ( .A1(n14799), .A2(n14803), .B1(n14759), .B2(n14798), .ZN(
        P1_U3474) );
  AOI21_X1 U16515 ( .B1(n14762), .B2(n14761), .A(n14760), .ZN(n14763) );
  OAI211_X1 U16516 ( .C1(n14766), .C2(n14765), .A(n14764), .B(n14763), .ZN(
        n14767) );
  INV_X1 U16517 ( .A(n14767), .ZN(n14805) );
  AOI22_X1 U16518 ( .A1(n14799), .A2(n14805), .B1(n7726), .B2(n14798), .ZN(
        P1_U3477) );
  OAI21_X1 U16519 ( .B1(n14769), .B2(n14781), .A(n14768), .ZN(n14772) );
  INV_X1 U16520 ( .A(n14770), .ZN(n14771) );
  AOI211_X1 U16521 ( .C1(n14787), .C2(n14773), .A(n14772), .B(n14771), .ZN(
        n14806) );
  AOI22_X1 U16522 ( .A1(n14799), .A2(n14806), .B1(n7743), .B2(n14798), .ZN(
        P1_U3480) );
  OAI211_X1 U16523 ( .C1(n14776), .C2(n14781), .A(n14775), .B(n14774), .ZN(
        n14778) );
  AOI211_X1 U16524 ( .C1(n14779), .C2(n14797), .A(n14778), .B(n14777), .ZN(
        n14807) );
  AOI22_X1 U16525 ( .A1(n14799), .A2(n14807), .B1(n7761), .B2(n14798), .ZN(
        P1_U3483) );
  OAI21_X1 U16526 ( .B1(n14782), .B2(n14781), .A(n14780), .ZN(n14785) );
  INV_X1 U16527 ( .A(n14783), .ZN(n14784) );
  AOI211_X1 U16528 ( .C1(n14787), .C2(n14786), .A(n14785), .B(n14784), .ZN(
        n14808) );
  INV_X1 U16529 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14788) );
  AOI22_X1 U16530 ( .A1(n14799), .A2(n14808), .B1(n14788), .B2(n14798), .ZN(
        P1_U3486) );
  INV_X1 U16531 ( .A(n14789), .ZN(n14791) );
  OAI211_X1 U16532 ( .C1(n14793), .C2(n14792), .A(n14791), .B(n14790), .ZN(
        n14795) );
  AOI211_X1 U16533 ( .C1(n14797), .C2(n14796), .A(n14795), .B(n14794), .ZN(
        n14810) );
  AOI22_X1 U16534 ( .A1(n14799), .A2(n14810), .B1(n7796), .B2(n14798), .ZN(
        P1_U3489) );
  AOI22_X1 U16535 ( .A1(n14811), .A2(n14800), .B1(n9972), .B2(n14809), .ZN(
        P1_U3531) );
  AOI22_X1 U16536 ( .A1(n14811), .A2(n14802), .B1(n14801), .B2(n14809), .ZN(
        P1_U3532) );
  AOI22_X1 U16537 ( .A1(n14811), .A2(n14803), .B1(n9973), .B2(n14809), .ZN(
        P1_U3533) );
  INV_X1 U16538 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n14804) );
  AOI22_X1 U16539 ( .A1(n14811), .A2(n14805), .B1(n14804), .B2(n14809), .ZN(
        P1_U3534) );
  AOI22_X1 U16540 ( .A1(n14811), .A2(n14806), .B1(n9974), .B2(n14809), .ZN(
        P1_U3535) );
  AOI22_X1 U16541 ( .A1(n14811), .A2(n14807), .B1(n10037), .B2(n14809), .ZN(
        P1_U3536) );
  AOI22_X1 U16542 ( .A1(n14811), .A2(n14808), .B1(n10196), .B2(n14809), .ZN(
        P1_U3537) );
  AOI22_X1 U16543 ( .A1(n14811), .A2(n14810), .B1(n10514), .B2(n14809), .ZN(
        P1_U3538) );
  NOR2_X1 U16544 ( .A1(n14924), .A2(P2_U3947), .ZN(P2_U3087) );
  OAI22_X1 U16545 ( .A1(n14822), .A2(n14812), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9148), .ZN(n14817) );
  AOI211_X1 U16546 ( .C1(n14815), .C2(n14814), .A(n14824), .B(n14813), .ZN(
        n14816) );
  AOI211_X1 U16547 ( .C1(n14818), .C2(n14829), .A(n14817), .B(n14816), .ZN(
        n14819) );
  OAI21_X1 U16548 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n14832), .A(n14819), .ZN(
        P2_U3190) );
  OAI22_X1 U16549 ( .A1(n14822), .A2(n14821), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14820), .ZN(n14828) );
  AOI211_X1 U16550 ( .C1(n14826), .C2(n14825), .A(n14824), .B(n14823), .ZN(
        n14827) );
  AOI211_X1 U16551 ( .C1(n14830), .C2(n14829), .A(n14828), .B(n14827), .ZN(
        n14831) );
  OAI21_X1 U16552 ( .B1(n14833), .B2(n14832), .A(n14831), .ZN(P2_U3206) );
  AOI22_X1 U16553 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n14941), .B1(n14863), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n14837) );
  AOI22_X1 U16554 ( .A1(n14924), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n14836) );
  OAI22_X1 U16555 ( .A1(n14932), .A2(P2_REG1_REG_0__SCAN_IN), .B1(
        P2_REG2_REG_0__SCAN_IN), .B2(n14913), .ZN(n14834) );
  OAI21_X1 U16556 ( .B1(n14939), .B2(n14834), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n14835) );
  OAI211_X1 U16557 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n14837), .A(n14836), .B(
        n14835), .ZN(P2_U3214) );
  AOI22_X1 U16558 ( .A1(n14924), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n14848) );
  XOR2_X1 U16559 ( .A(n14839), .B(n14838), .Z(n14842) );
  INV_X1 U16560 ( .A(n14895), .ZN(n14841) );
  AOI22_X1 U16561 ( .A1(n14863), .A2(n14842), .B1(n14841), .B2(n14840), .ZN(
        n14847) );
  AND2_X1 U16562 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n14845) );
  OAI211_X1 U16563 ( .C1(n14845), .C2(n14844), .A(n14941), .B(n14843), .ZN(
        n14846) );
  NAND3_X1 U16564 ( .A1(n14848), .A2(n14847), .A3(n14846), .ZN(P2_U3215) );
  AOI22_X1 U16565 ( .A1(n14924), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n14860) );
  OAI211_X1 U16566 ( .C1(n14851), .C2(n14850), .A(n14863), .B(n14849), .ZN(
        n14852) );
  OAI21_X1 U16567 ( .B1(n14930), .B2(n14853), .A(n14852), .ZN(n14854) );
  INV_X1 U16568 ( .A(n14854), .ZN(n14859) );
  OAI211_X1 U16569 ( .C1(n14857), .C2(n14856), .A(n14941), .B(n14855), .ZN(
        n14858) );
  NAND3_X1 U16570 ( .A1(n14860), .A2(n14859), .A3(n14858), .ZN(P2_U3216) );
  INV_X1 U16571 ( .A(n14861), .ZN(n14862) );
  OAI211_X1 U16572 ( .C1(n14865), .C2(n14864), .A(n14863), .B(n14862), .ZN(
        n14867) );
  NAND2_X1 U16573 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n14866) );
  OAI211_X1 U16574 ( .C1(n14930), .C2(n14868), .A(n14867), .B(n14866), .ZN(
        n14869) );
  INV_X1 U16575 ( .A(n14869), .ZN(n14875) );
  AOI211_X1 U16576 ( .C1(n14872), .C2(n14871), .A(n14870), .B(n14913), .ZN(
        n14873) );
  INV_X1 U16577 ( .A(n14873), .ZN(n14874) );
  OAI211_X1 U16578 ( .C1(n14946), .C2(n14876), .A(n14875), .B(n14874), .ZN(
        P2_U3218) );
  INV_X1 U16579 ( .A(n14877), .ZN(n14882) );
  AOI211_X1 U16580 ( .C1(n14880), .C2(n14879), .A(n14878), .B(n14932), .ZN(
        n14881) );
  AOI211_X1 U16581 ( .C1(n14939), .C2(n14883), .A(n14882), .B(n14881), .ZN(
        n14888) );
  OAI211_X1 U16582 ( .C1(n14886), .C2(n14885), .A(n14941), .B(n14884), .ZN(
        n14887) );
  OAI211_X1 U16583 ( .C1(n14946), .C2(n14889), .A(n14888), .B(n14887), .ZN(
        P2_U3220) );
  AOI211_X1 U16584 ( .C1(n14892), .C2(n14891), .A(n14932), .B(n14890), .ZN(
        n14897) );
  OAI21_X1 U16585 ( .B1(n14895), .B2(n14894), .A(n14893), .ZN(n14896) );
  NOR2_X1 U16586 ( .A1(n14897), .A2(n14896), .ZN(n14903) );
  AOI211_X1 U16587 ( .C1(n14900), .C2(n14899), .A(n14913), .B(n14898), .ZN(
        n14901) );
  INV_X1 U16588 ( .A(n14901), .ZN(n14902) );
  OAI211_X1 U16589 ( .C1(n14946), .C2(n14904), .A(n14903), .B(n14902), .ZN(
        P2_U3222) );
  NOR2_X1 U16590 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14905), .ZN(n14910) );
  AOI211_X1 U16591 ( .C1(n14908), .C2(n14907), .A(n14932), .B(n14906), .ZN(
        n14909) );
  AOI211_X1 U16592 ( .C1(n14939), .C2(n14911), .A(n14910), .B(n14909), .ZN(
        n14918) );
  AOI211_X1 U16593 ( .C1(n14915), .C2(n14914), .A(n14913), .B(n14912), .ZN(
        n14916) );
  INV_X1 U16594 ( .A(n14916), .ZN(n14917) );
  OAI211_X1 U16595 ( .C1(n14946), .C2(n6704), .A(n14918), .B(n14917), .ZN(
        P2_U3224) );
  NOR2_X1 U16596 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9304), .ZN(n14923) );
  AOI211_X1 U16597 ( .C1(n14921), .C2(n14920), .A(n14919), .B(n14932), .ZN(
        n14922) );
  AOI211_X1 U16598 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n14924), .A(n14923), 
        .B(n14922), .ZN(n14928) );
  OAI211_X1 U16599 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n14926), .A(n14941), 
        .B(n14925), .ZN(n14927) );
  OAI211_X1 U16600 ( .C1(n14930), .C2(n14929), .A(n14928), .B(n14927), .ZN(
        P2_U3229) );
  NOR2_X1 U16601 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14931), .ZN(n14937) );
  AOI211_X1 U16602 ( .C1(n14935), .C2(n14934), .A(n14933), .B(n14932), .ZN(
        n14936) );
  AOI211_X1 U16603 ( .C1(n14939), .C2(n14938), .A(n14937), .B(n14936), .ZN(
        n14945) );
  OAI211_X1 U16604 ( .C1(n14943), .C2(n14942), .A(n14941), .B(n14940), .ZN(
        n14944) );
  OAI211_X1 U16605 ( .C1(n14946), .C2(n6917), .A(n14945), .B(n14944), .ZN(
        P2_U3230) );
  NOR2_X1 U16606 ( .A1(n14957), .A2(n14947), .ZN(n14950) );
  AND2_X1 U16607 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14951), .ZN(P2_U3266) );
  AND2_X1 U16608 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14951), .ZN(P2_U3267) );
  AND2_X1 U16609 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14951), .ZN(P2_U3268) );
  AND2_X1 U16610 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14951), .ZN(P2_U3269) );
  AND2_X1 U16611 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14951), .ZN(P2_U3270) );
  AND2_X1 U16612 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14951), .ZN(P2_U3271) );
  AND2_X1 U16613 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14951), .ZN(P2_U3272) );
  AND2_X1 U16614 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14951), .ZN(P2_U3273) );
  AND2_X1 U16615 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14951), .ZN(P2_U3274) );
  AND2_X1 U16616 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14951), .ZN(P2_U3275) );
  AND2_X1 U16617 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14951), .ZN(P2_U3276) );
  AND2_X1 U16618 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14951), .ZN(P2_U3277) );
  AND2_X1 U16619 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14951), .ZN(P2_U3278) );
  AND2_X1 U16620 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14951), .ZN(P2_U3279) );
  AND2_X1 U16621 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14951), .ZN(P2_U3280) );
  AND2_X1 U16622 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14951), .ZN(P2_U3281) );
  NOR2_X1 U16623 ( .A1(n14950), .A2(n14948), .ZN(P2_U3282) );
  AND2_X1 U16624 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14951), .ZN(P2_U3283) );
  AND2_X1 U16625 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14951), .ZN(P2_U3284) );
  AND2_X1 U16626 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14951), .ZN(P2_U3285) );
  AND2_X1 U16627 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14951), .ZN(P2_U3286) );
  AND2_X1 U16628 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14951), .ZN(P2_U3287) );
  AND2_X1 U16629 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14951), .ZN(P2_U3288) );
  AND2_X1 U16630 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14951), .ZN(P2_U3289) );
  AND2_X1 U16631 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14951), .ZN(P2_U3290) );
  AND2_X1 U16632 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14951), .ZN(P2_U3291) );
  NOR2_X1 U16633 ( .A1(n14950), .A2(n14949), .ZN(P2_U3292) );
  AND2_X1 U16634 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14951), .ZN(P2_U3293) );
  AND2_X1 U16635 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14951), .ZN(P2_U3294) );
  AND2_X1 U16636 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14951), .ZN(P2_U3295) );
  AOI22_X1 U16637 ( .A1(n14954), .A2(n14953), .B1(n14952), .B2(n14957), .ZN(
        P2_U3416) );
  INV_X1 U16638 ( .A(n14955), .ZN(n14956) );
  AOI21_X1 U16639 ( .B1(n14958), .B2(n14957), .A(n14956), .ZN(P2_U3417) );
  OAI211_X1 U16640 ( .C1(n14987), .C2(n14961), .A(n14960), .B(n14959), .ZN(
        n14996) );
  OAI22_X1 U16641 ( .A1(n14994), .A2(n14996), .B1(P2_REG0_REG_0__SCAN_IN), 
        .B2(n14995), .ZN(n14962) );
  INV_X1 U16642 ( .A(n14962), .ZN(P2_U3430) );
  INV_X1 U16643 ( .A(n14986), .ZN(n14971) );
  NAND2_X1 U16644 ( .A1(n14970), .A2(n14963), .ZN(n14968) );
  NAND2_X1 U16645 ( .A1(n14964), .A2(n14972), .ZN(n14965) );
  NAND4_X1 U16646 ( .A1(n14968), .A2(n14967), .A3(n14966), .A4(n14965), .ZN(
        n14969) );
  AOI21_X1 U16647 ( .B1(n14971), .B2(n14970), .A(n14969), .ZN(n14998) );
  AOI22_X1 U16648 ( .A1(n14995), .A2(n14998), .B1(n9172), .B2(n14994), .ZN(
        P2_U3445) );
  INV_X1 U16649 ( .A(n14972), .ZN(n14989) );
  OAI211_X1 U16650 ( .C1(n14975), .C2(n14989), .A(n14974), .B(n14973), .ZN(
        n14976) );
  AOI21_X1 U16651 ( .B1(n14982), .B2(n14977), .A(n14976), .ZN(n14999) );
  AOI22_X1 U16652 ( .A1(n14995), .A2(n14999), .B1(n9184), .B2(n14994), .ZN(
        P2_U3448) );
  OAI211_X1 U16653 ( .C1(n14980), .C2(n14989), .A(n14979), .B(n14978), .ZN(
        n14981) );
  AOI21_X1 U16654 ( .B1(n14983), .B2(n14982), .A(n14981), .ZN(n15000) );
  INV_X1 U16655 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n14984) );
  AOI22_X1 U16656 ( .A1(n14995), .A2(n15000), .B1(n14984), .B2(n14994), .ZN(
        P2_U3451) );
  AOI21_X1 U16657 ( .B1(n14987), .B2(n14986), .A(n14985), .ZN(n14993) );
  OAI21_X1 U16658 ( .B1(n14990), .B2(n14989), .A(n14988), .ZN(n14991) );
  NOR3_X1 U16659 ( .A1(n14993), .A2(n14992), .A3(n14991), .ZN(n15001) );
  AOI22_X1 U16660 ( .A1(n14995), .A2(n15001), .B1(n9209), .B2(n14994), .ZN(
        P2_U3454) );
  OAI22_X1 U16661 ( .A1(n6478), .A2(n14996), .B1(P2_REG1_REG_0__SCAN_IN), .B2(
        n15002), .ZN(n14997) );
  INV_X1 U16662 ( .A(n14997), .ZN(P2_U3499) );
  AOI22_X1 U16663 ( .A1(n15002), .A2(n14998), .B1(n10084), .B2(n6478), .ZN(
        P2_U3504) );
  AOI22_X1 U16664 ( .A1(n15002), .A2(n14999), .B1(n9182), .B2(n6478), .ZN(
        P2_U3505) );
  AOI22_X1 U16665 ( .A1(n15002), .A2(n15000), .B1(n10085), .B2(n6478), .ZN(
        P2_U3506) );
  AOI22_X1 U16666 ( .A1(n15002), .A2(n15001), .B1(n10086), .B2(n6478), .ZN(
        P2_U3507) );
  NOR2_X1 U16667 ( .A1(P3_U3897), .A2(n15149), .ZN(P3_U3150) );
  INV_X1 U16668 ( .A(n6464), .ZN(n15004) );
  INV_X1 U16669 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n15214) );
  NAND2_X1 U16670 ( .A1(n15004), .A2(n15214), .ZN(n15005) );
  AND2_X1 U16671 ( .A1(n15006), .A2(n15005), .ZN(n15021) );
  INV_X1 U16672 ( .A(n15007), .ZN(n15008) );
  NOR2_X1 U16673 ( .A1(n15009), .A2(n15008), .ZN(n15010) );
  XNOR2_X1 U16674 ( .A(n15011), .B(n15010), .ZN(n15016) );
  AOI21_X1 U16675 ( .B1(n15149), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n15012), .ZN(
        n15013) );
  OAI21_X1 U16676 ( .B1(n15170), .B2(n15014), .A(n15013), .ZN(n15015) );
  AOI21_X1 U16677 ( .B1(n15016), .B2(n15178), .A(n15015), .ZN(n15020) );
  XOR2_X1 U16678 ( .A(P3_REG1_REG_5__SCAN_IN), .B(n15017), .Z(n15018) );
  NAND2_X1 U16679 ( .A1(n15176), .A2(n15018), .ZN(n15019) );
  OAI211_X1 U16680 ( .C1(n15021), .C2(n15184), .A(n15020), .B(n15019), .ZN(
        P3_U3187) );
  OAI21_X1 U16681 ( .B1(n15024), .B2(n15023), .A(n15022), .ZN(n15036) );
  AOI21_X1 U16682 ( .B1(n15027), .B2(n15026), .A(n15025), .ZN(n15029) );
  OAI22_X1 U16683 ( .A1(n15184), .A2(n15029), .B1(n15028), .B2(n15170), .ZN(
        n15035) );
  AOI21_X1 U16684 ( .B1(n15032), .B2(n15031), .A(n15030), .ZN(n15033) );
  NOR2_X1 U16685 ( .A1(n15033), .A2(n15158), .ZN(n15034) );
  AOI211_X1 U16686 ( .C1(n15176), .C2(n15036), .A(n15035), .B(n15034), .ZN(
        n15038) );
  OAI211_X1 U16687 ( .C1(n15039), .C2(n15173), .A(n15038), .B(n15037), .ZN(
        P3_U3188) );
  AOI21_X1 U16688 ( .B1(n15041), .B2(n12624), .A(n15040), .ZN(n15042) );
  INV_X1 U16689 ( .A(n15042), .ZN(n15055) );
  OAI21_X1 U16690 ( .B1(n15044), .B2(P3_REG1_REG_7__SCAN_IN), .A(n15043), .ZN(
        n15050) );
  AOI21_X1 U16691 ( .B1(n15047), .B2(n15046), .A(n15045), .ZN(n15048) );
  NOR2_X1 U16692 ( .A1(n15048), .A2(n15158), .ZN(n15049) );
  AOI21_X1 U16693 ( .B1(n15176), .B2(n15050), .A(n15049), .ZN(n15051) );
  OAI21_X1 U16694 ( .B1(n15052), .B2(n15170), .A(n15051), .ZN(n15053) );
  AOI21_X1 U16695 ( .B1(n15055), .B2(n15054), .A(n15053), .ZN(n15057) );
  NAND2_X1 U16696 ( .A1(P3_REG3_REG_7__SCAN_IN), .A2(P3_U3151), .ZN(n15056) );
  OAI211_X1 U16697 ( .C1(n15058), .C2(n15173), .A(n15057), .B(n15056), .ZN(
        P3_U3189) );
  OAI21_X1 U16698 ( .B1(n15061), .B2(n15060), .A(n15059), .ZN(n15073) );
  AOI21_X1 U16699 ( .B1(n15064), .B2(n15063), .A(n15062), .ZN(n15065) );
  OAI22_X1 U16700 ( .A1(n15170), .A2(n15066), .B1(n15065), .B2(n15158), .ZN(
        n15072) );
  AOI21_X1 U16701 ( .B1(n15069), .B2(n15068), .A(n15067), .ZN(n15070) );
  NOR2_X1 U16702 ( .A1(n15070), .A2(n15184), .ZN(n15071) );
  AOI211_X1 U16703 ( .C1(n15176), .C2(n15073), .A(n15072), .B(n15071), .ZN(
        n15075) );
  OAI211_X1 U16704 ( .C1(n15076), .C2(n15173), .A(n15075), .B(n15074), .ZN(
        P3_U3190) );
  AOI21_X1 U16705 ( .B1(n12620), .B2(n15078), .A(n15077), .ZN(n15091) );
  AOI21_X1 U16706 ( .B1(n15081), .B2(n15080), .A(n15079), .ZN(n15082) );
  OAI22_X1 U16707 ( .A1(n15170), .A2(n15083), .B1(n15082), .B2(n15158), .ZN(
        n15084) );
  AOI211_X1 U16708 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n15149), .A(n15085), .B(
        n15084), .ZN(n15090) );
  OAI21_X1 U16709 ( .B1(n15087), .B2(P3_REG1_REG_9__SCAN_IN), .A(n15086), .ZN(
        n15088) );
  NAND2_X1 U16710 ( .A1(n15088), .A2(n15176), .ZN(n15089) );
  OAI211_X1 U16711 ( .C1(n15091), .C2(n15184), .A(n15090), .B(n15089), .ZN(
        P3_U3191) );
  AOI21_X1 U16712 ( .B1(n15094), .B2(n15093), .A(n15092), .ZN(n15109) );
  OAI21_X1 U16713 ( .B1(n15097), .B2(n15096), .A(n15095), .ZN(n15098) );
  AND2_X1 U16714 ( .A1(n15098), .A2(n15176), .ZN(n15102) );
  OAI21_X1 U16715 ( .B1(n15170), .B2(n15100), .A(n15099), .ZN(n15101) );
  AOI211_X1 U16716 ( .C1(P3_ADDR_REG_10__SCAN_IN), .C2(n15149), .A(n15102), 
        .B(n15101), .ZN(n15108) );
  OAI21_X1 U16717 ( .B1(n15105), .B2(n15104), .A(n15103), .ZN(n15106) );
  NAND2_X1 U16718 ( .A1(n15106), .A2(n15178), .ZN(n15107) );
  OAI211_X1 U16719 ( .C1(n15109), .C2(n15184), .A(n15108), .B(n15107), .ZN(
        P3_U3192) );
  AOI21_X1 U16720 ( .B1(n8366), .B2(n15111), .A(n15110), .ZN(n15126) );
  OAI21_X1 U16721 ( .B1(n15113), .B2(P3_REG1_REG_11__SCAN_IN), .A(n15112), 
        .ZN(n15114) );
  AND2_X1 U16722 ( .A1(n15176), .A2(n15114), .ZN(n15119) );
  INV_X1 U16723 ( .A(n15115), .ZN(n15116) );
  OAI21_X1 U16724 ( .B1(n15170), .B2(n15117), .A(n15116), .ZN(n15118) );
  AOI211_X1 U16725 ( .C1(P3_ADDR_REG_11__SCAN_IN), .C2(n15149), .A(n15119), 
        .B(n15118), .ZN(n15125) );
  OAI21_X1 U16726 ( .B1(n15122), .B2(n15121), .A(n15120), .ZN(n15123) );
  NAND2_X1 U16727 ( .A1(n15123), .A2(n15178), .ZN(n15124) );
  OAI211_X1 U16728 ( .C1(n15126), .C2(n15184), .A(n15125), .B(n15124), .ZN(
        P3_U3193) );
  AOI21_X1 U16729 ( .B1(n15129), .B2(n15128), .A(n15127), .ZN(n15143) );
  OAI21_X1 U16730 ( .B1(n15132), .B2(n15131), .A(n15130), .ZN(n15133) );
  AND2_X1 U16731 ( .A1(n15133), .A2(n15176), .ZN(n15137) );
  NAND2_X1 U16732 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(P3_U3151), .ZN(n15134)
         );
  OAI21_X1 U16733 ( .B1(n15170), .B2(n15135), .A(n15134), .ZN(n15136) );
  AOI211_X1 U16734 ( .C1(P3_ADDR_REG_12__SCAN_IN), .C2(n15149), .A(n15137), 
        .B(n15136), .ZN(n15142) );
  OAI211_X1 U16735 ( .C1(n15140), .C2(n15139), .A(n15138), .B(n15178), .ZN(
        n15141) );
  OAI211_X1 U16736 ( .C1(n15143), .C2(n15184), .A(n15142), .B(n15141), .ZN(
        P3_U3194) );
  AOI21_X1 U16737 ( .B1(n11835), .B2(n15145), .A(n15144), .ZN(n15162) );
  OAI21_X1 U16738 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n15147), .A(n15146), 
        .ZN(n15153) );
  AND2_X1 U16739 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n15148) );
  AOI21_X1 U16740 ( .B1(n15149), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n15148), 
        .ZN(n15150) );
  OAI21_X1 U16741 ( .B1(n15170), .B2(n15151), .A(n15150), .ZN(n15152) );
  AOI21_X1 U16742 ( .B1(n15153), .B2(n15176), .A(n15152), .ZN(n15161) );
  INV_X1 U16743 ( .A(n15154), .ZN(n15155) );
  AOI21_X1 U16744 ( .B1(n15157), .B2(n15156), .A(n15155), .ZN(n15159) );
  OR2_X1 U16745 ( .A1(n15159), .A2(n15158), .ZN(n15160) );
  OAI211_X1 U16746 ( .C1(n15162), .C2(n15184), .A(n15161), .B(n15160), .ZN(
        P3_U3195) );
  AOI21_X1 U16747 ( .B1(n15165), .B2(n15164), .A(n15163), .ZN(n15185) );
  OAI21_X1 U16748 ( .B1(n15168), .B2(n15167), .A(n15166), .ZN(n15177) );
  NOR2_X1 U16749 ( .A1(n15170), .A2(n15169), .ZN(n15175) );
  OAI21_X1 U16750 ( .B1(n15173), .B2(n15172), .A(n15171), .ZN(n15174) );
  AOI211_X1 U16751 ( .C1(n15177), .C2(n15176), .A(n15175), .B(n15174), .ZN(
        n15183) );
  OAI211_X1 U16752 ( .C1(n15181), .C2(n15180), .A(n15179), .B(n15178), .ZN(
        n15182) );
  OAI211_X1 U16753 ( .C1(n15185), .C2(n15184), .A(n15183), .B(n15182), .ZN(
        P3_U3196) );
  OAI21_X1 U16754 ( .B1(n15188), .B2(n15187), .A(n15186), .ZN(n15297) );
  INV_X1 U16755 ( .A(n15297), .ZN(n15195) );
  AOI22_X1 U16756 ( .A1(n15259), .A2(n15190), .B1(n15189), .B2(n15256), .ZN(
        n15194) );
  OAI211_X1 U16757 ( .C1(n6666), .C2(n15192), .A(n15262), .B(n15191), .ZN(
        n15193) );
  OAI211_X1 U16758 ( .C1(n15195), .C2(n15266), .A(n15194), .B(n15193), .ZN(
        n15295) );
  AOI21_X1 U16759 ( .B1(n15251), .B2(n15297), .A(n15295), .ZN(n15201) );
  NOR2_X1 U16760 ( .A1(n15196), .A2(n15253), .ZN(n15296) );
  INV_X1 U16761 ( .A(n15197), .ZN(n15198) );
  AOI22_X1 U16762 ( .A1(n15227), .A2(n15296), .B1(n15226), .B2(n15198), .ZN(
        n15199) );
  OAI221_X1 U16763 ( .B1(n12719), .B2(n15201), .C1(n15273), .C2(n15200), .A(
        n15199), .ZN(P3_U3227) );
  XNOR2_X1 U16764 ( .A(n15203), .B(n15202), .ZN(n15294) );
  XNOR2_X1 U16765 ( .A(n15204), .B(n15205), .ZN(n15206) );
  OAI222_X1 U16766 ( .A1(n15243), .A2(n15208), .B1(n15241), .B2(n15207), .C1(
        n15206), .C2(n15249), .ZN(n15291) );
  AOI21_X1 U16767 ( .B1(n15294), .B2(n15209), .A(n15291), .ZN(n15215) );
  NOR2_X1 U16768 ( .A1(n15210), .A2(n15253), .ZN(n15292) );
  INV_X1 U16769 ( .A(n15211), .ZN(n15212) );
  AOI22_X1 U16770 ( .A1(n15227), .A2(n15292), .B1(n15226), .B2(n15212), .ZN(
        n15213) );
  OAI221_X1 U16771 ( .B1(n12719), .B2(n15215), .C1(n15273), .C2(n15214), .A(
        n15213), .ZN(P3_U3228) );
  XNOR2_X1 U16772 ( .A(n15216), .B(n15219), .ZN(n15223) );
  INV_X1 U16773 ( .A(n15223), .ZN(n15286) );
  AOI22_X1 U16774 ( .A1(n15256), .A2(n15258), .B1(n15217), .B2(n15259), .ZN(
        n15222) );
  OAI211_X1 U16775 ( .C1(n15220), .C2(n15219), .A(n15218), .B(n15262), .ZN(
        n15221) );
  OAI211_X1 U16776 ( .C1(n15223), .C2(n15266), .A(n15222), .B(n15221), .ZN(
        n15284) );
  AOI21_X1 U16777 ( .B1(n15251), .B2(n15286), .A(n15284), .ZN(n15229) );
  NOR2_X1 U16778 ( .A1(n15224), .A2(n15253), .ZN(n15285) );
  AOI22_X1 U16779 ( .A1(n15227), .A2(n15285), .B1(n15226), .B2(n15225), .ZN(
        n15228) );
  OAI221_X1 U16780 ( .B1(n12719), .B2(n15229), .C1(n15273), .C2(n8216), .A(
        n15228), .ZN(P3_U3230) );
  NAND3_X1 U16781 ( .A1(n15232), .A2(n15231), .A3(n15230), .ZN(n15233) );
  NAND2_X1 U16782 ( .A1(n15234), .A2(n15233), .ZN(n15282) );
  NOR2_X1 U16783 ( .A1(n15235), .A2(n15253), .ZN(n15281) );
  INV_X1 U16784 ( .A(n15281), .ZN(n15238) );
  OAI22_X1 U16785 ( .A1(n15238), .A2(n15237), .B1(n15236), .B2(n15268), .ZN(
        n15250) );
  XNOR2_X1 U16786 ( .A(n15240), .B(n15239), .ZN(n15248) );
  OAI22_X1 U16787 ( .A1(n15244), .A2(n15243), .B1(n15242), .B2(n15241), .ZN(
        n15245) );
  AOI21_X1 U16788 ( .B1(n15282), .B2(n15246), .A(n15245), .ZN(n15247) );
  OAI21_X1 U16789 ( .B1(n15249), .B2(n15248), .A(n15247), .ZN(n15280) );
  AOI211_X1 U16790 ( .C1(n15251), .C2(n15282), .A(n15250), .B(n15280), .ZN(
        n15252) );
  AOI22_X1 U16791 ( .A1(n12719), .A2(n8174), .B1(n15252), .B2(n15273), .ZN(
        P3_U3231) );
  NOR2_X1 U16792 ( .A1(n15254), .A2(n15253), .ZN(n15278) );
  XNOR2_X1 U16793 ( .A(n15255), .B(n15261), .ZN(n15276) );
  AOI22_X1 U16794 ( .A1(n15259), .A2(n15258), .B1(n15257), .B2(n15256), .ZN(
        n15265) );
  XNOR2_X1 U16795 ( .A(n15261), .B(n15260), .ZN(n15263) );
  NAND2_X1 U16796 ( .A1(n15263), .A2(n15262), .ZN(n15264) );
  OAI211_X1 U16797 ( .C1(n15276), .C2(n15266), .A(n15265), .B(n15264), .ZN(
        n15277) );
  AOI21_X1 U16798 ( .B1(n15278), .B2(n15267), .A(n15277), .ZN(n15274) );
  OAI22_X1 U16799 ( .A1(n15270), .A2(n15276), .B1(n15269), .B2(n15268), .ZN(
        n15271) );
  INV_X1 U16800 ( .A(n15271), .ZN(n15272) );
  OAI221_X1 U16801 ( .B1(n12719), .B2(n15274), .C1(n15273), .C2(n8203), .A(
        n15272), .ZN(P3_U3232) );
  INV_X1 U16802 ( .A(n15276), .ZN(n15279) );
  AOI211_X1 U16803 ( .C1(n15312), .C2(n15279), .A(n15278), .B(n15277), .ZN(
        n15319) );
  AOI22_X1 U16804 ( .A1(n15318), .A2(n15319), .B1(n8202), .B2(n15316), .ZN(
        P3_U3393) );
  AOI211_X1 U16805 ( .C1(n15312), .C2(n15282), .A(n15281), .B(n15280), .ZN(
        n15320) );
  INV_X1 U16806 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15283) );
  AOI22_X1 U16807 ( .A1(n15318), .A2(n15320), .B1(n15283), .B2(n15316), .ZN(
        P3_U3396) );
  AOI211_X1 U16808 ( .C1(n15286), .C2(n15312), .A(n15285), .B(n15284), .ZN(
        n15322) );
  AOI22_X1 U16809 ( .A1(n15318), .A2(n15322), .B1(n8215), .B2(n15316), .ZN(
        P3_U3399) );
  INV_X1 U16810 ( .A(n15287), .ZN(n15289) );
  AOI211_X1 U16811 ( .C1(n15290), .C2(n15312), .A(n15289), .B(n15288), .ZN(
        n15323) );
  AOI22_X1 U16812 ( .A1(n15318), .A2(n15323), .B1(n8233), .B2(n15316), .ZN(
        P3_U3402) );
  AOI211_X1 U16813 ( .C1(n15294), .C2(n15293), .A(n15292), .B(n15291), .ZN(
        n15324) );
  AOI22_X1 U16814 ( .A1(n15318), .A2(n15324), .B1(n8252), .B2(n15316), .ZN(
        P3_U3405) );
  AOI211_X1 U16815 ( .C1(n15312), .C2(n15297), .A(n15296), .B(n15295), .ZN(
        n15325) );
  AOI22_X1 U16816 ( .A1(n15318), .A2(n15325), .B1(n8269), .B2(n15316), .ZN(
        P3_U3408) );
  INV_X1 U16817 ( .A(n15298), .ZN(n15301) );
  AOI211_X1 U16818 ( .C1(n15301), .C2(n15312), .A(n15300), .B(n15299), .ZN(
        n15326) );
  INV_X1 U16819 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15302) );
  AOI22_X1 U16820 ( .A1(n15318), .A2(n15326), .B1(n15302), .B2(n15316), .ZN(
        P3_U3411) );
  AOI211_X1 U16821 ( .C1(n15312), .C2(n15305), .A(n15304), .B(n15303), .ZN(
        n15327) );
  AOI22_X1 U16822 ( .A1(n15318), .A2(n15327), .B1(n8311), .B2(n15316), .ZN(
        P3_U3414) );
  AOI21_X1 U16823 ( .B1(n15307), .B2(n15312), .A(n15306), .ZN(n15308) );
  AND2_X1 U16824 ( .A1(n15309), .A2(n15308), .ZN(n15328) );
  INV_X1 U16825 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15310) );
  AOI22_X1 U16826 ( .A1(n15318), .A2(n15328), .B1(n15310), .B2(n15316), .ZN(
        P3_U3417) );
  AOI21_X1 U16827 ( .B1(n15313), .B2(n15312), .A(n15311), .ZN(n15314) );
  INV_X1 U16828 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15317) );
  AOI22_X1 U16829 ( .A1(n15318), .A2(n15330), .B1(n15317), .B2(n15316), .ZN(
        P3_U3420) );
  AOI22_X1 U16830 ( .A1(n15331), .A2(n15319), .B1(n10782), .B2(n15329), .ZN(
        P3_U3460) );
  AOI22_X1 U16831 ( .A1(n15331), .A2(n15320), .B1(n10447), .B2(n15329), .ZN(
        P3_U3461) );
  INV_X1 U16832 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15321) );
  AOI22_X1 U16833 ( .A1(n15331), .A2(n15322), .B1(n15321), .B2(n15329), .ZN(
        P3_U3462) );
  AOI22_X1 U16834 ( .A1(n15331), .A2(n15323), .B1(n12590), .B2(n15329), .ZN(
        P3_U3463) );
  AOI22_X1 U16835 ( .A1(n15331), .A2(n15324), .B1(n12597), .B2(n15329), .ZN(
        P3_U3464) );
  AOI22_X1 U16836 ( .A1(n15331), .A2(n15325), .B1(n12625), .B2(n15329), .ZN(
        P3_U3465) );
  AOI22_X1 U16837 ( .A1(n15331), .A2(n15326), .B1(n12623), .B2(n15329), .ZN(
        P3_U3466) );
  AOI22_X1 U16838 ( .A1(n15331), .A2(n15327), .B1(n12621), .B2(n15329), .ZN(
        P3_U3467) );
  AOI22_X1 U16839 ( .A1(n15331), .A2(n15328), .B1(n12619), .B2(n15329), .ZN(
        P3_U3468) );
  AOI22_X1 U16840 ( .A1(n15331), .A2(n15330), .B1(n12589), .B2(n15329), .ZN(
        P3_U3469) );
  OAI21_X1 U16841 ( .B1(n15334), .B2(n15333), .A(n15332), .ZN(SUB_1596_U59) );
  OAI21_X1 U16842 ( .B1(n15337), .B2(n15336), .A(n15335), .ZN(SUB_1596_U58) );
  XOR2_X1 U16843 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15338), .Z(SUB_1596_U53) );
  AOI21_X1 U16844 ( .B1(n15341), .B2(n15340), .A(n15339), .ZN(SUB_1596_U56) );
  AOI21_X1 U16845 ( .B1(n15344), .B2(n15343), .A(n15342), .ZN(n15345) );
  XOR2_X1 U16846 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15345), .Z(SUB_1596_U60) );
  AOI21_X1 U16847 ( .B1(n15348), .B2(n15347), .A(n15346), .ZN(SUB_1596_U5) );
  OAI21_X2 U7255 ( .B1(n7578), .B2(P1_IR_REG_27__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7577) );
  NOR2_X2 U8319 ( .A1(n14524), .A2(n12147), .ZN(n6943) );
  OR2_X2 U8566 ( .A1(n14505), .A2(n14531), .ZN(n14506) );
  OR2_X1 U9926 ( .A1(n7673), .A2(n9876), .ZN(n7659) );
  OR2_X1 U10487 ( .A1(n14705), .A2(n14704), .ZN(n14706) );
  AND2_X2 U10490 ( .A1(n14684), .A2(n14769), .ZN(n14682) );
  OR2_X1 U10484 ( .A1(n10191), .A2(n12089), .ZN(n14725) );
  INV_X1 U7228 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9454) );
  NAND2_X2 U9855 ( .A1(n7676), .A2(n9854), .ZN(n12236) );
  INV_X1 U9935 ( .A(n12092), .ZN(n12089) );
  AND2_X1 U9366 ( .A1(n14099), .A2(n6563), .ZN(n14020) );
  NAND2_X1 U7322 ( .A1(n12698), .A2(n8848), .ZN(n9015) );
  CLKBUF_X3 U7320 ( .A(n8569), .Z(n6477) );
  INV_X1 U7514 ( .A(n7676), .ZN(n7936) );
  CLKBUF_X1 U7588 ( .A(n13760), .Z(n6676) );
  OAI211_X1 U8797 ( .C1(n7676), .C2(n13878), .A(n7675), .B(n7674), .ZN(n14724)
         );
  NAND2_X1 U9154 ( .A1(n13918), .A2(n14726), .ZN(n14130) );
endmodule

