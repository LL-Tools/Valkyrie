

module b21_C_gen_AntiSAT_k_256_10 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2, 
        keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7, 
        keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12, 
        keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17, 
        keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22, 
        keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27, 
        keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32, 
        keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37, 
        keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42, 
        keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47, 
        keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52, 
        keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57, 
        keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62, 
        keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67, 
        keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72, 
        keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77, 
        keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82, 
        keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87, 
        keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92, 
        keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97, 
        keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4475, n4476, n4478, n4479, n4480, n4481, n4482, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10484;

  INV_X1 U4980 ( .A(P1_STATE_REG_SCAN_IN), .ZN(n10484) );
  NOR2_X1 U4981 ( .A1(n5960), .A2(n5961), .ZN(n8688) );
  OR2_X1 U4982 ( .A1(n8861), .A2(n8654), .ZN(n5964) );
  INV_X1 U4983 ( .A(n5312), .ZN(n5604) );
  CLKBUF_X2 U4984 ( .A(n6128), .Z(n6666) );
  CLKBUF_X1 U4985 ( .A(n6127), .Z(n6458) );
  CLKBUF_X1 U4986 ( .A(n6118), .Z(n4481) );
  CLKBUF_X1 U4987 ( .A(n6118), .Z(n4485) );
  BUF_X1 U4988 ( .A(n7377), .Z(n4479) );
  BUF_X1 U4989 ( .A(n6675), .Z(n4487) );
  INV_X1 U4990 ( .A(n10484), .ZN(n4475) );
  INV_X1 U4991 ( .A(n4475), .ZN(n4476) );
  INV_X1 U4992 ( .A(n4475), .ZN(P1_U3084) );
  INV_X1 U4993 ( .A(n5981), .ZN(n4635) );
  OR2_X1 U4995 ( .A1(n9928), .A2(n9927), .ZN(n9929) );
  NOR2_X1 U4996 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5314) );
  BUF_X1 U5000 ( .A(n6180), .Z(n8134) );
  OR2_X1 U5001 ( .A1(n6059), .A2(n9536), .ZN(n6061) );
  INV_X1 U5002 ( .A(n7337), .ZN(n5743) );
  CLKBUF_X3 U5003 ( .A(n5305), .Z(n5834) );
  INV_X1 U5004 ( .A(n8835), .ZN(n8797) );
  AND2_X1 U5005 ( .A1(n9194), .A2(n9198), .ZN(n9195) );
  NAND2_X1 U5006 ( .A1(n6673), .A2(n6672), .ZN(n7492) );
  INV_X1 U5007 ( .A(n6702), .ZN(n9811) );
  NAND2_X1 U5008 ( .A1(n6048), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6074) );
  INV_X4 U5009 ( .A(n6835), .ZN(n8129) );
  XNOR2_X1 U5010 ( .A(n5248), .B(P2_IR_REG_21__SCAN_IN), .ZN(n5868) );
  NAND2_X2 U5011 ( .A1(n6675), .A2(n8430), .ZN(n8130) );
  OR3_X1 U5012 ( .A1(n9552), .A2(n8005), .A3(n8069), .ZN(n6800) );
  XNOR2_X1 U5013 ( .A(n6074), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6656) );
  NAND2_X1 U5014 ( .A1(n6592), .A2(n6591), .ZN(n9252) );
  XNOR2_X1 U5015 ( .A(n6053), .B(n6052), .ZN(n9552) );
  INV_X1 U5016 ( .A(n9317), .ZN(n9331) );
  NOR2_X2 U5017 ( .A1(n5517), .A2(n10318), .ZN(n5539) );
  AND2_X1 U5018 ( .A1(n9947), .A2(n7741), .ZN(n4478) );
  AND2_X1 U5019 ( .A1(n9947), .A2(n7741), .ZN(n6882) );
  OAI21_X2 U5020 ( .B1(n9228), .B2(n5086), .A(n5084), .ZN(n5093) );
  NAND2_X2 U5021 ( .A1(n6734), .A2(n6733), .ZN(n9228) );
  OAI22_X2 U5023 ( .A1(n7890), .A2(n6277), .B1(n7888), .B2(n7887), .ZN(n7932)
         );
  NOR2_X2 U5024 ( .A1(n9196), .A2(n9195), .ZN(n9410) );
  OAI211_X2 U5025 ( .C1(n8130), .C2(n7075), .A(n6201), .B(n6200), .ZN(n7784)
         );
  NAND4_X1 U5026 ( .A1(n6042), .A2(n6041), .A3(n6040), .A4(n6039), .ZN(n6695)
         );
  OAI211_X1 U5027 ( .C1(n8130), .C2(n6962), .A(n6109), .B(n6108), .ZN(n7377)
         );
  NAND2_X2 U5028 ( .A1(n4800), .A2(n4798), .ZN(n6694) );
  XNOR2_X2 U5029 ( .A(n4755), .B(n4754), .ZN(n9542) );
  NOR2_X2 U5030 ( .A1(n6794), .A2(n6795), .ZN(n5634) );
  OAI21_X2 U5031 ( .B1(n5601), .B2(n5024), .A(n5022), .ZN(n6794) );
  AND2_X1 U5032 ( .A1(n8085), .A2(n8970), .ZN(n4480) );
  AND2_X1 U5033 ( .A1(n8085), .A2(n8970), .ZN(n5290) );
  INV_X2 U5034 ( .A(n5868), .ZN(n7782) );
  XNOR2_X2 U5035 ( .A(n5236), .B(n5265), .ZN(n5793) );
  AND2_X1 U5036 ( .A1(n6070), .A2(n6800), .ZN(n6118) );
  OAI222_X1 U5037 ( .A1(n9552), .A2(n4476), .B1(n8089), .B2(n9551), .C1(n9550), 
        .C2(n9549), .ZN(P1_U3327) );
  NAND2_X1 U5038 ( .A1(n6717), .A2(n6716), .ZN(n9617) );
  OAI21_X1 U5039 ( .B1(n7976), .B2(n4804), .A(n4801), .ZN(n9621) );
  OR2_X1 U5040 ( .A1(n5710), .A2(n8537), .ZN(n5735) );
  AND2_X1 U5041 ( .A1(n8459), .A2(n5336), .ZN(n8510) );
  INV_X2 U5042 ( .A(n7784), .ZN(n7682) );
  INV_X1 U5043 ( .A(n7661), .ZN(n7363) );
  CLKBUF_X2 U5044 ( .A(n6486), .Z(n6628) );
  CLKBUF_X2 U5045 ( .A(n6160), .Z(n6556) );
  NAND4_X1 U5046 ( .A1(n6114), .A2(n6113), .A3(n6112), .A4(n6111), .ZN(n9138)
         );
  INV_X2 U5047 ( .A(n6694), .ZN(n6742) );
  CLKBUF_X2 U5048 ( .A(n6125), .Z(n6587) );
  CLKBUF_X2 U5049 ( .A(n6126), .Z(n6501) );
  NAND2_X2 U5050 ( .A1(n5782), .A2(n7782), .ZN(n5020) );
  INV_X1 U5051 ( .A(n5778), .ZN(n5782) );
  XNOR2_X1 U5052 ( .A(n6061), .B(n6060), .ZN(n6675) );
  OAI21_X1 U5053 ( .B1(n4824), .B2(n9833), .A(n4767), .ZN(n6785) );
  NOR2_X1 U5054 ( .A1(n9191), .A2(n4531), .ZN(n4768) );
  OR2_X1 U5055 ( .A1(n4831), .A2(n4830), .ZN(n4659) );
  OAI21_X1 U5056 ( .B1(n5827), .B2(n5826), .A(n5974), .ZN(n5844) );
  OAI211_X1 U5057 ( .C1(n5672), .C2(n4698), .A(n4695), .B(n4694), .ZN(n8487)
         );
  NAND2_X1 U5058 ( .A1(n5672), .A2(n5671), .ZN(n4703) );
  OAI21_X1 U5059 ( .B1(n8240), .B2(n8239), .A(n8238), .ZN(n8251) );
  NAND2_X1 U5060 ( .A1(n8684), .A2(n5104), .ZN(n8687) );
  NAND2_X1 U5061 ( .A1(n8696), .A2(n8697), .ZN(n8684) );
  NAND2_X1 U5062 ( .A1(n5241), .A2(n5240), .ZN(n5817) );
  NAND2_X1 U5063 ( .A1(n6714), .A2(n5102), .ZN(n5045) );
  NAND2_X1 U5064 ( .A1(n6543), .A2(n6542), .ZN(n9428) );
  NAND2_X1 U5065 ( .A1(n5077), .A2(n5076), .ZN(n7967) );
  OR2_X1 U5066 ( .A1(n7545), .A2(n7546), .ZN(n7596) );
  NOR2_X1 U5067 ( .A1(n4530), .A2(n5044), .ZN(n5043) );
  NAND2_X1 U5068 ( .A1(n6412), .A2(n6411), .ZN(n9465) );
  INV_X2 U5069 ( .A(n8839), .ZN(n9936) );
  NAND2_X1 U5070 ( .A1(n9660), .A2(n7505), .ZN(n9654) );
  NAND2_X1 U5071 ( .A1(n6132), .A2(n4520), .ZN(n6701) );
  NAND4_X1 U5072 ( .A1(n6151), .A2(n6150), .A3(n6149), .A4(n6148), .ZN(n9137)
         );
  NAND4_X1 U5073 ( .A1(n6089), .A2(n6088), .A3(n6087), .A4(n6086), .ZN(n6696)
         );
  AND4_X1 U5074 ( .A1(n5343), .A2(n5342), .A3(n5341), .A4(n5340), .ZN(n5809)
         );
  AND4_X1 U5075 ( .A1(n5375), .A2(n5374), .A3(n5373), .A4(n5372), .ZN(n7410)
         );
  AND2_X2 U5076 ( .A1(n6808), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  AND2_X1 U5077 ( .A1(n6656), .A2(n8339), .ZN(n6070) );
  AND3_X2 U5078 ( .A1(n5301), .A2(n5300), .A3(n5299), .ZN(n7141) );
  NAND4_X1 U5079 ( .A1(n5294), .A2(n5293), .A3(n5292), .A4(n5291), .ZN(n5805)
         );
  NAND2_X1 U5080 ( .A1(n6049), .A2(n6048), .ZN(n8339) );
  INV_X2 U5081 ( .A(n5289), .ZN(n5843) );
  NAND2_X1 U5082 ( .A1(n6051), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6053) );
  XNOR2_X1 U5083 ( .A(n5749), .B(P2_IR_REG_22__SCAN_IN), .ZN(n5778) );
  NAND2_X1 U5084 ( .A1(n6409), .A2(n4994), .ZN(n6048) );
  XNOR2_X1 U5085 ( .A(n6056), .B(n6055), .ZN(n8005) );
  XNOR2_X1 U5086 ( .A(n6058), .B(n6057), .ZN(n8069) );
  NOR2_X1 U5087 ( .A1(n6387), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n6409) );
  NAND2_X1 U5088 ( .A1(n4655), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5267) );
  NAND2_X1 U5089 ( .A1(n6050), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6058) );
  OR2_X1 U5090 ( .A1(n5266), .A2(n5386), .ZN(n5236) );
  AND2_X1 U5091 ( .A1(n5063), .A2(n4746), .ZN(n6034) );
  AND2_X1 U5092 ( .A1(n6054), .A2(n5063), .ZN(n6059) );
  NOR2_X1 U5093 ( .A1(n5441), .A2(n10102), .ZN(n5460) );
  NOR3_X1 U5094 ( .A1(n5529), .A2(n4850), .A3(P2_IR_REG_29__SCAN_IN), .ZN(
        n4653) );
  NAND2_X2 U5095 ( .A1(n4779), .A2(n4778), .ZN(n5216) );
  AND4_X1 U5096 ( .A1(n5229), .A2(n5356), .A3(n5228), .A4(n4569), .ZN(n5587)
         );
  NOR2_X1 U5097 ( .A1(n4501), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5064) );
  NOR2_X1 U5098 ( .A1(n5015), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5014) );
  AND4_X1 U5099 ( .A1(n6027), .A2(n6302), .A3(n6028), .A4(n6263), .ZN(n6029)
         );
  NAND3_X1 U5100 ( .A1(n5108), .A2(n4622), .A3(n4621), .ZN(n4779) );
  NAND3_X1 U5101 ( .A1(n4620), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4778) );
  AND2_X1 U5102 ( .A1(n5227), .A2(n5226), .ZN(n5228) );
  INV_X1 U5103 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6198) );
  INV_X1 U5104 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6052) );
  NOR2_X1 U5105 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5221) );
  NOR2_X1 U5106 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5222) );
  NOR2_X1 U5107 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5223) );
  INV_X1 U5108 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4621) );
  INV_X1 U5109 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5108) );
  INV_X1 U5110 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6057) );
  INV_X1 U5111 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6428) );
  NOR2_X1 U5112 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n6302) );
  NOR2_X1 U5113 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n6028) );
  INV_X1 U5114 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6073) );
  AND2_X1 U5115 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5359) );
  NOR2_X1 U5116 ( .A1(n8817), .A2(n8816), .ZN(n8815) );
  NOR2_X2 U5117 ( .A1(n8861), .A2(n8678), .ZN(n8661) );
  AOI21_X2 U5118 ( .B1(n6718), .B2(n4497), .A(n4533), .ZN(n8091) );
  XNOR2_X2 U5119 ( .A(n6695), .B(n6742), .ZN(n6741) );
  INV_X2 U5120 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  OAI21_X1 U5121 ( .B1(n8026), .B2(n4646), .A(n5927), .ZN(n4645) );
  INV_X1 U5122 ( .A(n5925), .ZN(n4646) );
  AND4_X1 U5123 ( .A1(n6025), .A2(n6024), .A3(n6198), .A4(n6023), .ZN(n6026)
         );
  INV_X1 U5124 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6025) );
  INV_X1 U5125 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6024) );
  INV_X1 U5126 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U5127 ( .A1(n5471), .A2(n5154), .ZN(n4957) );
  INV_X1 U5128 ( .A(n5834), .ZN(n5546) );
  INV_X1 U5129 ( .A(n8688), .ZN(n4897) );
  AND2_X1 U5130 ( .A1(n5007), .A2(n4678), .ZN(n4677) );
  NAND2_X1 U5131 ( .A1(n5104), .A2(n8621), .ZN(n4678) );
  NOR2_X1 U5132 ( .A1(n8651), .A2(n5008), .ZN(n5007) );
  INV_X1 U5133 ( .A(n5816), .ZN(n5008) );
  OR2_X1 U5134 ( .A1(n9609), .A2(n8061), .ZN(n5922) );
  NAND2_X1 U5135 ( .A1(n7993), .A2(n4983), .ZN(n4982) );
  NOR2_X1 U5136 ( .A1(n8036), .A2(n4984), .ZN(n4983) );
  INV_X1 U5137 ( .A(n6326), .ZN(n4984) );
  AND2_X1 U5138 ( .A1(n8138), .A2(n8137), .ZN(n8378) );
  INV_X1 U5139 ( .A(n6735), .ZN(n5092) );
  NAND2_X1 U5140 ( .A1(n6711), .A2(n5083), .ZN(n5082) );
  NAND2_X1 U5141 ( .A1(n4934), .A2(n4933), .ZN(n5831) );
  AOI21_X1 U5142 ( .B1(n4511), .B2(n4938), .A(n4590), .ZN(n4933) );
  NAND2_X1 U5143 ( .A1(n5721), .A2(n4511), .ZN(n4934) );
  INV_X1 U5144 ( .A(n5220), .ZN(n4938) );
  AND2_X1 U5145 ( .A1(n5187), .A2(n5186), .ZN(n5618) );
  NAND2_X1 U5146 ( .A1(n5793), .A2(n8977), .ZN(n5313) );
  AND2_X1 U5147 ( .A1(n6658), .A2(n6659), .ZN(n8987) );
  NAND2_X1 U5148 ( .A1(n8130), .A2(n8129), .ZN(n6155) );
  NAND2_X1 U5149 ( .A1(n8130), .A2(n6835), .ZN(n6180) );
  NAND2_X1 U5150 ( .A1(n5811), .A2(n5892), .ZN(n4640) );
  NOR2_X1 U5151 ( .A1(n4846), .A2(n5941), .ZN(n4845) );
  OAI21_X1 U5152 ( .B1(n5926), .B2(n4642), .A(n4641), .ZN(n5939) );
  NAND2_X1 U5153 ( .A1(n4647), .A2(n4644), .ZN(n4641) );
  NAND2_X1 U5154 ( .A1(n4647), .A2(n4643), .ZN(n4642) );
  INV_X1 U5155 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n6263) );
  NAND2_X1 U5156 ( .A1(n5133), .A2(n10430), .ZN(n5136) );
  NAND2_X1 U5157 ( .A1(n4898), .A2(n8651), .ZN(n4894) );
  NAND2_X1 U5158 ( .A1(n8664), .A2(n8654), .ZN(n4899) );
  AND2_X1 U5159 ( .A1(n8867), .A2(n8670), .ZN(n5961) );
  NOR2_X1 U5160 ( .A1(n8727), .A2(n5019), .ZN(n5018) );
  NAND2_X1 U5161 ( .A1(n8883), .A2(n8752), .ZN(n4882) );
  NOR2_X1 U5162 ( .A1(n8747), .A2(n4881), .ZN(n4880) );
  INV_X1 U5163 ( .A(n8615), .ZN(n4881) );
  NAND2_X1 U5164 ( .A1(n8909), .A2(n8611), .ZN(n4913) );
  INV_X1 U5165 ( .A(n5917), .ZN(n4669) );
  AND2_X1 U5166 ( .A1(n5917), .A2(n5918), .ZN(n7917) );
  OR2_X1 U5167 ( .A1(n9927), .A2(n7548), .ZN(n5894) );
  NOR2_X1 U5168 ( .A1(n7408), .A2(n4871), .ZN(n4870) );
  INV_X1 U5169 ( .A(n7402), .ZN(n4871) );
  INV_X1 U5170 ( .A(n9542), .ZN(n6037) );
  AOI21_X1 U5171 ( .B1(n5080), .B2(n5079), .A(n4538), .ZN(n5078) );
  INV_X1 U5172 ( .A(n5083), .ZN(n5079) );
  AND2_X1 U5173 ( .A1(n6026), .A2(n4560), .ZN(n4748) );
  AND2_X1 U5174 ( .A1(n5098), .A2(n10403), .ZN(n4995) );
  AOI21_X1 U5175 ( .B1(n4493), .B2(n4712), .A(n4550), .ZN(n4705) );
  NAND2_X1 U5176 ( .A1(n4929), .A2(n4930), .ZN(n5381) );
  AOI21_X1 U5177 ( .B1(n4931), .B2(n5364), .A(n4544), .ZN(n4930) );
  OAI211_X1 U5178 ( .C1(n4629), .C2(n4628), .A(n4521), .B(n4627), .ZN(n4929)
         );
  INV_X1 U5179 ( .A(n6106), .ZN(n6022) );
  NAND2_X1 U5180 ( .A1(n8523), .A2(n8522), .ZN(n5672) );
  NAND2_X1 U5181 ( .A1(n5670), .A2(n5669), .ZN(n5671) );
  NAND2_X1 U5182 ( .A1(n8053), .A2(n5559), .ZN(n5028) );
  AOI21_X1 U5183 ( .B1(n5614), .B2(n5023), .A(n4500), .ZN(n5022) );
  AND2_X1 U5184 ( .A1(n5451), .A2(n5435), .ZN(n5036) );
  NAND2_X1 U5185 ( .A1(n4612), .A2(n4611), .ZN(n4610) );
  INV_X1 U5186 ( .A(n7195), .ZN(n4611) );
  INV_X1 U5187 ( .A(n7196), .ZN(n4612) );
  AND4_X1 U5188 ( .A1(n5550), .A2(n5549), .A3(n5548), .A4(n5547), .ZN(n8061)
         );
  AND4_X1 U5189 ( .A1(n5399), .A2(n5398), .A3(n5397), .A4(n5396), .ZN(n7485)
         );
  INV_X1 U5190 ( .A(n8085), .ZN(n4680) );
  NAND2_X1 U5192 ( .A1(n5003), .A2(n5104), .ZN(n4676) );
  NAND2_X1 U5193 ( .A1(n4675), .A2(n5003), .ZN(n4674) );
  AND2_X1 U5194 ( .A1(n5005), .A2(n5818), .ZN(n5003) );
  OR2_X1 U5195 ( .A1(n8867), .A2(n8622), .ZN(n4900) );
  NAND2_X1 U5196 ( .A1(n4885), .A2(n4895), .ZN(n4901) );
  OR2_X1 U5197 ( .A1(n8889), .A2(n8763), .ZN(n5935) );
  OAI21_X1 U5198 ( .B1(n8025), .B2(n4552), .A(n5009), .ZN(n8817) );
  NAND2_X1 U5199 ( .A1(n5010), .A2(n4525), .ZN(n5009) );
  NAND2_X1 U5200 ( .A1(n8828), .A2(n5012), .ZN(n5010) );
  INV_X1 U5201 ( .A(n8795), .ZN(n9917) );
  NAND2_X1 U5202 ( .A1(n5621), .A2(n5620), .ZN(n8900) );
  NAND2_X1 U5203 ( .A1(n4982), .A2(n4985), .ZN(n6363) );
  XNOR2_X1 U5204 ( .A(n6080), .B(n7492), .ZN(n6100) );
  NAND2_X1 U5205 ( .A1(n6072), .A2(n6071), .ZN(n6080) );
  OAI211_X1 U5206 ( .C1(n8378), .C2(n8268), .A(n4918), .B(n4916), .ZN(n8427)
         );
  NAND2_X1 U5207 ( .A1(n4919), .A2(n4528), .ZN(n4918) );
  OAI21_X1 U5208 ( .B1(n8378), .B2(n4917), .A(n8262), .ZN(n4916) );
  AND2_X1 U5209 ( .A1(n9172), .A2(n9175), .ZN(n8426) );
  INV_X1 U5210 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6060) );
  INV_X1 U5211 ( .A(n9198), .ZN(n5087) );
  AND2_X1 U5212 ( .A1(n9203), .A2(n9217), .ZN(n5094) );
  NAND2_X1 U5213 ( .A1(n6726), .A2(n6729), .ZN(n5073) );
  NAND2_X1 U5214 ( .A1(n7976), .A2(n8361), .ZN(n4807) );
  NAND2_X1 U5215 ( .A1(n6739), .A2(n6738), .ZN(n6774) );
  INV_X1 U5216 ( .A(n6600), .ZN(n4990) );
  NAND2_X1 U5217 ( .A1(n4548), .A2(n4635), .ZN(n4634) );
  INV_X1 U5218 ( .A(n4640), .ZN(n4639) );
  NOR2_X1 U5219 ( .A1(n4640), .A2(n5889), .ZN(n4637) );
  INV_X1 U5220 ( .A(n4840), .ZN(n4839) );
  OAI21_X1 U5221 ( .B1(n4848), .B2(n4841), .A(n4535), .ZN(n4840) );
  NAND2_X1 U5222 ( .A1(n4649), .A2(n4635), .ZN(n4648) );
  INV_X1 U5223 ( .A(n5946), .ZN(n4649) );
  NAND2_X1 U5224 ( .A1(n4651), .A2(n4519), .ZN(n4650) );
  NAND2_X1 U5225 ( .A1(n5945), .A2(n4652), .ZN(n4651) );
  AND2_X1 U5226 ( .A1(n5943), .A2(n5944), .ZN(n4652) );
  OAI21_X1 U5227 ( .B1(n5955), .B2(n4546), .A(n4856), .ZN(n4855) );
  NOR2_X1 U5228 ( .A1(n5959), .A2(n5960), .ZN(n4856) );
  NOR2_X1 U5229 ( .A1(n5962), .A2(n5963), .ZN(n4854) );
  OR2_X1 U5230 ( .A1(n9428), .A2(n9038), .ZN(n8318) );
  OAI21_X1 U5231 ( .B1(n4626), .B2(n4543), .A(n4623), .ZN(n4826) );
  AOI21_X1 U5232 ( .B1(n5972), .B2(n4624), .A(n5976), .ZN(n4623) );
  AOI21_X1 U5233 ( .B1(n5972), .B2(n8671), .A(n8626), .ZN(n4626) );
  OR2_X1 U5234 ( .A1(n8852), .A2(n8653), .ZN(n5973) );
  AND2_X1 U5235 ( .A1(n9180), .A2(n8260), .ZN(n8265) );
  OR2_X1 U5236 ( .A1(n9180), .A2(n8335), .ZN(n8372) );
  AND2_X1 U5237 ( .A1(n4944), .A2(n4948), .ZN(n4943) );
  NOR2_X1 U5238 ( .A1(n5690), .A2(n4949), .ZN(n4948) );
  NAND2_X1 U5239 ( .A1(n4946), .A2(n5674), .ZN(n4944) );
  INV_X1 U5240 ( .A(n5204), .ZN(n4949) );
  INV_X1 U5241 ( .A(n4946), .ZN(n4945) );
  INV_X1 U5242 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5165) );
  INV_X1 U5243 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5149) );
  NOR2_X1 U5244 ( .A1(n7388), .A2(n5034), .ZN(n5033) );
  INV_X1 U5245 ( .A(n5379), .ZN(n5034) );
  NAND2_X1 U5246 ( .A1(n8687), .A2(n5816), .ZN(n8665) );
  NOR2_X1 U5247 ( .A1(n8883), .A2(n4791), .ZN(n4790) );
  INV_X1 U5248 ( .A(n4792), .ZN(n4791) );
  INV_X1 U5249 ( .A(n4515), .ZN(n5001) );
  NOR2_X1 U5250 ( .A1(n8889), .A2(n8895), .ZN(n4792) );
  XNOR2_X1 U5251 ( .A(n7467), .B(n5807), .ZN(n7160) );
  OR2_X1 U5252 ( .A1(n5546), .A2(n6902), .ZN(n5340) );
  OR2_X1 U5253 ( .A1(n5806), .A2(n9952), .ZN(n5874) );
  NAND2_X1 U5254 ( .A1(n5994), .A2(n6883), .ZN(n5867) );
  INV_X1 U5255 ( .A(n7328), .ZN(n7332) );
  INV_X1 U5256 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5235) );
  NAND2_X1 U5257 ( .A1(n5750), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5774) );
  INV_X1 U5258 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5748) );
  INV_X1 U5259 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5246) );
  AOI21_X1 U5260 ( .B1(n6447), .B2(n4725), .A(n4723), .ZN(n4722) );
  NAND2_X1 U5261 ( .A1(n6473), .A2(n4724), .ZN(n4723) );
  NAND2_X1 U5262 ( .A1(n4726), .A2(n4725), .ZN(n4724) );
  NAND2_X1 U5263 ( .A1(n8377), .A2(n8336), .ZN(n8375) );
  OR2_X1 U5264 ( .A1(n9742), .A2(n4717), .ZN(n7716) );
  AND2_X1 U5265 ( .A1(n9747), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4717) );
  OR2_X1 U5266 ( .A1(n9203), .A2(n8993), .ZN(n8330) );
  OR2_X1 U5267 ( .A1(n9423), .A2(n9106), .ZN(n8269) );
  INV_X1 U5268 ( .A(n6731), .ZN(n5075) );
  NOR2_X1 U5269 ( .A1(n4771), .A2(n9443), .ZN(n4770) );
  INV_X1 U5270 ( .A(n4772), .ZN(n4771) );
  NOR2_X1 U5271 ( .A1(n9455), .A2(n9449), .ZN(n4772) );
  INV_X1 U5272 ( .A(n9349), .ZN(n4816) );
  OR2_X1 U5273 ( .A1(n7895), .A2(n9645), .ZN(n8292) );
  NAND2_X1 U5274 ( .A1(n8287), .A2(n8379), .ZN(n8145) );
  NOR2_X1 U5275 ( .A1(n8142), .A2(n8387), .ZN(n8383) );
  OR2_X1 U5276 ( .A1(n9134), .A2(n7622), .ZN(n8275) );
  AND2_X1 U5277 ( .A1(n8199), .A2(n8198), .ZN(n9364) );
  AND2_X1 U5278 ( .A1(n8339), .A2(n9331), .ZN(n6678) );
  INV_X1 U5279 ( .A(n8339), .ZN(n8417) );
  AOI21_X1 U5280 ( .B1(n4924), .B2(n4926), .A(n4922), .ZN(n4921) );
  INV_X1 U5281 ( .A(n5187), .ZN(n4922) );
  OAI21_X1 U5282 ( .B1(n5552), .B2(n5551), .A(n5164), .ZN(n5528) );
  OAI21_X1 U5283 ( .B1(n4955), .B2(n4710), .A(n4952), .ZN(n4709) );
  OR2_X1 U5284 ( .A1(n4495), .A2(n4711), .ZN(n4710) );
  NAND2_X1 U5285 ( .A1(n4956), .A2(n5148), .ZN(n4712) );
  NAND2_X1 U5286 ( .A1(n5151), .A2(n5150), .ZN(n5154) );
  INV_X1 U5287 ( .A(SI_12_), .ZN(n5150) );
  NAND2_X1 U5288 ( .A1(n4707), .A2(n5148), .ZN(n5472) );
  OAI21_X1 U5289 ( .B1(n4686), .B2(n4685), .A(n4683), .ZN(n5436) );
  INV_X1 U5290 ( .A(n5132), .ZN(n4686) );
  AOI21_X1 U5291 ( .B1(n4689), .B2(n4691), .A(n4684), .ZN(n4683) );
  INV_X1 U5292 ( .A(n5136), .ZN(n4691) );
  NAND2_X1 U5293 ( .A1(n4693), .A2(n5131), .ZN(n4692) );
  INV_X1 U5294 ( .A(n5405), .ZN(n4693) );
  INV_X1 U5295 ( .A(n5344), .ZN(n4632) );
  AOI21_X1 U5296 ( .B1(n4631), .B2(n5344), .A(n4549), .ZN(n4630) );
  INV_X1 U5297 ( .A(n5121), .ZN(n4631) );
  AND2_X1 U5298 ( .A1(n4602), .A2(n8486), .ZN(n4601) );
  INV_X1 U5299 ( .A(n8533), .ZN(n4602) );
  AND3_X1 U5300 ( .A1(n4617), .A2(n4614), .A3(n4613), .ZN(n8455) );
  NAND2_X1 U5301 ( .A1(n5603), .A2(n9849), .ZN(n4613) );
  NAND2_X1 U5302 ( .A1(n5604), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n4617) );
  NAND2_X1 U5303 ( .A1(n4616), .A2(n4615), .ZN(n4614) );
  NAND2_X1 U5304 ( .A1(n8121), .A2(n5613), .ZN(n5024) );
  XNOR2_X1 U5305 ( .A(n5617), .B(n5615), .ZN(n8121) );
  OAI21_X1 U5306 ( .B1(n8487), .B2(n4598), .A(n4595), .ZN(n4603) );
  AOI21_X1 U5307 ( .B1(n4599), .B2(n4597), .A(n4596), .ZN(n4595) );
  INV_X1 U5308 ( .A(n4599), .ZN(n4598) );
  INV_X1 U5309 ( .A(n4601), .ZN(n4597) );
  INV_X1 U5310 ( .A(n8495), .ZN(n4700) );
  INV_X1 U5311 ( .A(n8498), .ZN(n4699) );
  INV_X1 U5312 ( .A(n4701), .ZN(n4604) );
  AOI22_X1 U5313 ( .A1(n5687), .A2(n4702), .B1(n5689), .B2(n5688), .ZN(n4701)
         );
  INV_X1 U5314 ( .A(n5671), .ZN(n4696) );
  NAND3_X1 U5315 ( .A1(n5020), .A2(n7782), .A3(n6885), .ZN(n5257) );
  XNOR2_X1 U5316 ( .A(n8455), .B(n5744), .ZN(n5333) );
  INV_X1 U5317 ( .A(n5033), .ZN(n5032) );
  INV_X1 U5318 ( .A(n4609), .ZN(n4607) );
  AOI21_X1 U5319 ( .B1(n5033), .B2(n5031), .A(n5030), .ZN(n5029) );
  INV_X1 U5320 ( .A(n5404), .ZN(n5030) );
  INV_X1 U5321 ( .A(n7301), .ZN(n5031) );
  OR2_X1 U5322 ( .A1(n5608), .A2(n5607), .ZN(n5622) );
  NOR2_X1 U5323 ( .A1(n6789), .A2(n5040), .ZN(n5039) );
  NAND2_X1 U5324 ( .A1(n8468), .A2(n5651), .ZN(n5668) );
  NAND2_X1 U5325 ( .A1(n5260), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5608) );
  INV_X1 U5326 ( .A(n5592), .ZN(n5260) );
  NAND2_X1 U5327 ( .A1(n8074), .A2(n5584), .ZN(n5601) );
  NAND2_X1 U5328 ( .A1(n7196), .A2(n7195), .ZN(n4609) );
  INV_X1 U5329 ( .A(n6014), .ZN(n4829) );
  AND4_X1 U5330 ( .A1(n5538), .A2(n5537), .A3(n5536), .A4(n5535), .ZN(n8607)
         );
  NAND2_X1 U5331 ( .A1(n8649), .A2(n4785), .ZN(n4784) );
  NOR2_X1 U5332 ( .A1(n4894), .A2(n4896), .ZN(n4890) );
  OAI21_X1 U5333 ( .B1(n4894), .B2(n4888), .A(n4892), .ZN(n4887) );
  AOI21_X1 U5334 ( .B1(n4898), .B2(n4893), .A(n4545), .ZN(n4892) );
  NAND2_X1 U5335 ( .A1(n4895), .A2(n4513), .ZN(n4888) );
  NAND2_X1 U5336 ( .A1(n4673), .A2(n4677), .ZN(n5004) );
  OR2_X1 U5337 ( .A1(n8696), .A2(n4679), .ZN(n4673) );
  NAND2_X1 U5338 ( .A1(n8623), .A2(n5006), .ZN(n5005) );
  INV_X1 U5339 ( .A(n5964), .ZN(n5006) );
  AND2_X1 U5340 ( .A1(n8665), .A2(n5964), .ZN(n8652) );
  NAND2_X1 U5341 ( .A1(n8666), .A2(n4899), .ZN(n4898) );
  NAND2_X1 U5342 ( .A1(n8876), .A2(n8619), .ZN(n8620) );
  AND2_X1 U5343 ( .A1(n5702), .A2(n5701), .ZN(n8715) );
  AND2_X1 U5344 ( .A1(n8712), .A2(n5950), .ZN(n5016) );
  NAND2_X1 U5345 ( .A1(n4875), .A2(n4882), .ZN(n4873) );
  INV_X1 U5346 ( .A(n4878), .ZN(n4877) );
  OAI22_X1 U5347 ( .A1(n8747), .A2(n4879), .B1(n8889), .B2(n8616), .ZN(n4878)
         );
  INV_X1 U5348 ( .A(n4884), .ZN(n4879) );
  NAND2_X1 U5349 ( .A1(n8758), .A2(n4880), .ZN(n4876) );
  NOR2_X1 U5350 ( .A1(n8895), .A2(n8749), .ZN(n4884) );
  AND2_X1 U5351 ( .A1(n5667), .A2(n5666), .ZN(n8763) );
  AND2_X1 U5352 ( .A1(n5629), .A2(n5628), .ZN(n8762) );
  NOR2_X1 U5353 ( .A1(n8760), .A2(n4846), .ZN(n5002) );
  NAND2_X1 U5354 ( .A1(n8781), .A2(n8613), .ZN(n8786) );
  AOI21_X1 U5355 ( .B1(n4489), .B2(n4908), .A(n4556), .ZN(n4903) );
  NAND2_X1 U5356 ( .A1(n4910), .A2(n4541), .ZN(n4909) );
  INV_X1 U5357 ( .A(n4914), .ZN(n4910) );
  NAND2_X1 U5358 ( .A1(n8064), .A2(n8607), .ZN(n5012) );
  NAND2_X1 U5359 ( .A1(n4863), .A2(n4581), .ZN(n4862) );
  AOI21_X1 U5360 ( .B1(n4671), .B2(n4670), .A(n4669), .ZN(n4664) );
  INV_X1 U5361 ( .A(n4671), .ZN(n4665) );
  INV_X1 U5362 ( .A(n4667), .ZN(n4666) );
  OAI21_X1 U5363 ( .B1(n4671), .B2(n4669), .A(n7941), .ZN(n4667) );
  AND2_X1 U5364 ( .A1(n5922), .A2(n5921), .ZN(n7941) );
  AND2_X1 U5365 ( .A1(n5912), .A2(n7917), .ZN(n4671) );
  NAND2_X1 U5366 ( .A1(n7872), .A2(n7871), .ZN(n4672) );
  INV_X1 U5367 ( .A(n7917), .ZN(n7924) );
  OAI21_X1 U5368 ( .B1(n7649), .B2(n4860), .A(n4858), .ZN(n7869) );
  AOI21_X1 U5369 ( .B1(n4861), .B2(n4859), .A(n4537), .ZN(n4858) );
  INV_X1 U5370 ( .A(n4861), .ZN(n4860) );
  AND4_X1 U5371 ( .A1(n5503), .A2(n5502), .A3(n5501), .A4(n5500), .ZN(n7918)
         );
  INV_X1 U5372 ( .A(n4868), .ZN(n4867) );
  AOI21_X1 U5373 ( .B1(n4868), .B2(n4866), .A(n4540), .ZN(n4865) );
  NOR2_X1 U5374 ( .A1(n5811), .A2(n4869), .ZN(n4868) );
  OAI211_X1 U5375 ( .C1(n5103), .C2(n4997), .A(n4996), .B(n5997), .ZN(n7417)
         );
  NAND2_X1 U5376 ( .A1(n5882), .A2(n7440), .ZN(n4996) );
  INV_X1 U5377 ( .A(n8750), .ZN(n8818) );
  OR2_X1 U5378 ( .A1(n6915), .A2(n5798), .ZN(n8820) );
  NAND2_X1 U5379 ( .A1(n5874), .A2(n5877), .ZN(n7328) );
  NAND2_X1 U5380 ( .A1(n6885), .A2(n6884), .ZN(n8795) );
  OR2_X1 U5381 ( .A1(n8561), .A2(n7203), .ZN(n6883) );
  NAND2_X1 U5382 ( .A1(n5606), .A2(n5605), .ZN(n8906) );
  NAND2_X1 U5383 ( .A1(n7669), .A2(n4616), .ZN(n5606) );
  AND2_X1 U5384 ( .A1(n5761), .A2(n5759), .ZN(n9937) );
  NAND2_X1 U5385 ( .A1(n5014), .A2(n5265), .ZN(n4850) );
  NOR2_X1 U5386 ( .A1(n5529), .A2(n4850), .ZN(n4654) );
  NAND2_X1 U5387 ( .A1(n5774), .A2(n5773), .ZN(n5776) );
  INV_X1 U5388 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5255) );
  INV_X1 U5389 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5251) );
  INV_X1 U5390 ( .A(n7521), .ZN(n4753) );
  INV_X1 U5391 ( .A(n6189), .ZN(n4750) );
  INV_X1 U5392 ( .A(n4732), .ZN(n4731) );
  INV_X1 U5393 ( .A(n7585), .ZN(n4963) );
  NOR2_X1 U5394 ( .A1(n7795), .A2(n4966), .ZN(n4965) );
  OR2_X1 U5395 ( .A1(n6448), .A2(n4727), .ZN(n4725) );
  NAND2_X1 U5396 ( .A1(n4993), .A2(n4992), .ZN(n9042) );
  AND2_X1 U5397 ( .A1(n6407), .A2(n6386), .ZN(n4992) );
  AOI21_X1 U5398 ( .B1(n4742), .B2(n4743), .A(n4576), .ZN(n4740) );
  NOR2_X1 U5399 ( .A1(n4741), .A2(n4737), .ZN(n4736) );
  INV_X1 U5400 ( .A(n4742), .ZN(n4739) );
  NOR2_X1 U5401 ( .A1(n7832), .A2(n4733), .ZN(n4732) );
  INV_X1 U5402 ( .A(n4964), .ZN(n4733) );
  AND2_X1 U5403 ( .A1(n6094), .A2(n6093), .ZN(n6805) );
  NAND2_X1 U5404 ( .A1(n4976), .A2(n6472), .ZN(n9019) );
  INV_X1 U5405 ( .A(n9021), .ZN(n4976) );
  NAND2_X1 U5406 ( .A1(n6325), .A2(n6324), .ZN(n7993) );
  NAND2_X1 U5407 ( .A1(n9028), .A2(n9027), .ZN(n6510) );
  AND2_X1 U5408 ( .A1(n4960), .A2(n6169), .ZN(n4959) );
  NAND2_X1 U5409 ( .A1(n7308), .A2(n6187), .ZN(n4960) );
  INV_X1 U5410 ( .A(n6070), .ZN(n6672) );
  NAND2_X1 U5411 ( .A1(n8433), .A2(n9331), .ZN(n6673) );
  OR2_X1 U5412 ( .A1(n6127), .A2(n6035), .ZN(n6042) );
  OR2_X1 U5413 ( .A1(n6125), .A2(n7513), .ZN(n6041) );
  NOR2_X1 U5414 ( .A1(n7085), .A2(n4574), .ZN(n7131) );
  OR2_X1 U5415 ( .A1(n7131), .A2(n7130), .ZN(n4716) );
  OR2_X1 U5416 ( .A1(n6327), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6346) );
  NOR2_X1 U5417 ( .A1(n9744), .A2(n9743), .ZN(n9742) );
  AOI21_X1 U5418 ( .B1(n5091), .B2(n6736), .A(n4539), .ZN(n5089) );
  AND2_X1 U5419 ( .A1(n8330), .A2(n8329), .ZN(n9198) );
  NAND2_X1 U5420 ( .A1(n6583), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6621) );
  AND2_X1 U5421 ( .A1(n8232), .A2(n8228), .ZN(n9275) );
  AOI21_X1 U5422 ( .B1(n4492), .B2(n5051), .A(n4578), .ZN(n5047) );
  AOI21_X1 U5423 ( .B1(n9308), .B2(n8219), .A(n8221), .ZN(n4797) );
  OR2_X1 U5424 ( .A1(n6753), .A2(n9309), .ZN(n4796) );
  AND2_X1 U5425 ( .A1(n8213), .A2(n8218), .ZN(n9333) );
  NAND2_X1 U5426 ( .A1(n8096), .A2(n8315), .ZN(n9350) );
  AOI21_X1 U5427 ( .B1(n5057), .B2(n5060), .A(n4584), .ZN(n5054) );
  OR2_X1 U5428 ( .A1(n6770), .A2(n9381), .ZN(n5062) );
  NAND2_X1 U5429 ( .A1(n6770), .A2(n9381), .ZN(n5061) );
  NAND2_X1 U5430 ( .A1(n4510), .A2(n4773), .ZN(n9388) );
  NOR2_X1 U5431 ( .A1(n4776), .A2(n9390), .ZN(n4775) );
  NOR2_X1 U5432 ( .A1(n8360), .A2(n4806), .ZN(n4805) );
  INV_X1 U5433 ( .A(n8172), .ZN(n4806) );
  NAND2_X1 U5434 ( .A1(n4807), .A2(n8172), .ZN(n8006) );
  AOI21_X1 U5435 ( .B1(n4551), .B2(n5078), .A(n4498), .ZN(n5076) );
  INV_X1 U5436 ( .A(n8134), .ZN(n6450) );
  INV_X1 U5437 ( .A(n8130), .ZN(n6449) );
  NAND2_X1 U5438 ( .A1(n6758), .A2(n8132), .ZN(n9649) );
  OR2_X1 U5439 ( .A1(n8425), .A2(n9687), .ZN(n9646) );
  OR2_X1 U5440 ( .A1(n8425), .A2(n4487), .ZN(n9644) );
  INV_X1 U5441 ( .A(n9649), .ZN(n9326) );
  INV_X1 U5442 ( .A(n9646), .ZN(n9379) );
  NAND2_X1 U5443 ( .A1(n6775), .A2(n9808), .ZN(n7151) );
  AND2_X1 U5444 ( .A1(n9175), .A2(n9174), .ZN(n9403) );
  OR2_X1 U5445 ( .A1(n6155), .A2(n6853), .ZN(n6201) );
  AND4_X1 U5446 ( .A1(n4592), .A2(n4748), .A3(n6029), .A4(n4747), .ZN(n4746)
         );
  AND2_X1 U5447 ( .A1(n6022), .A2(n6060), .ZN(n4747) );
  XNOR2_X1 U5448 ( .A(n6032), .B(P1_IR_REG_29__SCAN_IN), .ZN(n6036) );
  OR2_X1 U5449 ( .A1(n6034), .A2(n9536), .ZN(n6032) );
  NAND2_X1 U5450 ( .A1(n5215), .A2(n5214), .ZN(n5721) );
  AND2_X1 U5451 ( .A1(n5220), .A2(n5219), .ZN(n5720) );
  XNOR2_X1 U5452 ( .A(n5691), .B(n5690), .ZN(n8067) );
  NAND2_X1 U5453 ( .A1(n4950), .A2(n5204), .ZN(n5691) );
  NAND2_X1 U5454 ( .A1(n5676), .A2(n4946), .ZN(n4950) );
  AND2_X1 U5455 ( .A1(n6409), .A2(n4995), .ZN(n6045) );
  AND2_X1 U5456 ( .A1(n4995), .A2(n6044), .ZN(n4994) );
  NAND2_X1 U5457 ( .A1(n4923), .A2(n5183), .ZN(n5619) );
  NAND2_X1 U5458 ( .A1(n5178), .A2(n4927), .ZN(n4923) );
  XNOR2_X1 U5459 ( .A(n5406), .B(n5405), .ZN(n6865) );
  XNOR2_X1 U5460 ( .A(n5128), .B(n5127), .ZN(n5364) );
  XNOR2_X1 U5461 ( .A(n5125), .B(n10413), .ZN(n5353) );
  OR3_X1 U5462 ( .A1(n7991), .A2(n8982), .A3(n8070), .ZN(n6916) );
  NAND2_X1 U5463 ( .A1(n4594), .A2(n4599), .ZN(n8438) );
  NAND2_X1 U5464 ( .A1(n8487), .A2(n4601), .ZN(n4594) );
  INV_X1 U5465 ( .A(n5024), .ZN(n5614) );
  AND2_X1 U5466 ( .A1(n5817), .A2(n5026), .ZN(n5025) );
  NAND2_X1 U5467 ( .A1(n5785), .A2(n8542), .ZN(n5026) );
  NAND2_X1 U5468 ( .A1(n7482), .A2(n5431), .ZN(n7572) );
  AND4_X1 U5469 ( .A1(n5522), .A2(n5521), .A3(n5520), .A4(n5519), .ZN(n7950)
         );
  NAND2_X1 U5470 ( .A1(n5601), .A2(n8073), .ZN(n8120) );
  NAND2_X1 U5471 ( .A1(n5709), .A2(n5708), .ZN(n8867) );
  AND2_X1 U5472 ( .A1(n7741), .A2(n8835), .ZN(n6017) );
  NAND2_X1 U5473 ( .A1(n7407), .A2(n5891), .ZN(n9916) );
  NOR2_X1 U5474 ( .A1(n4583), .A2(n4508), .ZN(n4989) );
  NAND2_X1 U5475 ( .A1(n6512), .A2(n6511), .ZN(n9438) );
  NAND2_X1 U5476 ( .A1(n6664), .A2(n9655), .ZN(n9095) );
  INV_X1 U5477 ( .A(n9267), .ZN(n9106) );
  AOI21_X1 U5478 ( .B1(n4980), .B2(n4527), .A(n4977), .ZN(n9101) );
  NAND2_X1 U5479 ( .A1(n4978), .A2(n4582), .ZN(n4977) );
  OAI211_X1 U5480 ( .C1(n4523), .C2(n8428), .A(n4488), .B(n4491), .ZN(n8429)
         );
  NAND2_X1 U5481 ( .A1(n6054), .A2(n5064), .ZN(n6062) );
  NAND2_X1 U5482 ( .A1(n6627), .A2(n6626), .ZN(n9217) );
  NAND2_X1 U5483 ( .A1(n6535), .A2(n6534), .ZN(n9303) );
  NAND4_X1 U5484 ( .A1(n6197), .A2(n6196), .A3(n6195), .A4(n6194), .ZN(n9135)
         );
  OR2_X1 U5485 ( .A1(n6663), .A2(n7845), .ZN(n9655) );
  NAND2_X1 U5486 ( .A1(n4825), .A2(n4768), .ZN(n4824) );
  INV_X1 U5487 ( .A(n9185), .ZN(n4825) );
  INV_X1 U5488 ( .A(n4832), .ZN(n5873) );
  OAI21_X1 U5489 ( .B1(n5883), .B2(n4542), .A(n4833), .ZN(n4832) );
  NOR2_X1 U5490 ( .A1(n5865), .A2(n5866), .ZN(n4833) );
  OAI21_X1 U5491 ( .B1(n5882), .B2(n4635), .A(n4834), .ZN(n5883) );
  NAND2_X1 U5492 ( .A1(n4835), .A2(n4635), .ZN(n4834) );
  NAND2_X1 U5493 ( .A1(n5997), .A2(n5864), .ZN(n4835) );
  NAND2_X1 U5494 ( .A1(n4638), .A2(n4636), .ZN(n5901) );
  NOR2_X1 U5495 ( .A1(n4837), .A2(n4637), .ZN(n4636) );
  NAND2_X1 U5496 ( .A1(n5896), .A2(n7603), .ZN(n4837) );
  OAI21_X1 U5497 ( .B1(n5916), .B2(n4670), .A(n5915), .ZN(n5920) );
  INV_X1 U5498 ( .A(n4645), .ZN(n4643) );
  INV_X1 U5499 ( .A(n5932), .ZN(n4647) );
  MUX2_X1 U5500 ( .A(n8177), .B(n8300), .S(n8262), .Z(n8196) );
  NAND2_X1 U5501 ( .A1(n4515), .A2(n5940), .ZN(n4848) );
  OR2_X1 U5502 ( .A1(n4845), .A2(n4847), .ZN(n4841) );
  AND2_X1 U5503 ( .A1(n4849), .A2(n5944), .ZN(n4847) );
  NOR2_X1 U5504 ( .A1(n5933), .A2(n8791), .ZN(n4849) );
  NOR2_X1 U5505 ( .A1(n4848), .A2(n4843), .ZN(n4842) );
  OR2_X1 U5506 ( .A1(n4845), .A2(n4844), .ZN(n4843) );
  OAI21_X1 U5507 ( .B1(n5939), .B2(n4844), .A(n5938), .ZN(n5942) );
  MUX2_X1 U5508 ( .A(n8212), .B(n8211), .S(n8267), .Z(n8216) );
  MUX2_X1 U5509 ( .A(n4635), .B(n5936), .S(n5935), .Z(n5947) );
  AND2_X1 U5510 ( .A1(n8175), .A2(n8172), .ZN(n8299) );
  NAND2_X1 U5511 ( .A1(n4855), .A2(n4854), .ZN(n5970) );
  INV_X1 U5512 ( .A(n4625), .ZN(n4624) );
  OAI21_X1 U5513 ( .B1(n5817), .B2(n4635), .A(n5971), .ZN(n4625) );
  OAI21_X1 U5514 ( .B1(n8251), .B2(n8250), .A(n8249), .ZN(n8252) );
  NAND2_X1 U5515 ( .A1(n5979), .A2(n4828), .ZN(n4827) );
  INV_X1 U5516 ( .A(n5975), .ZN(n4828) );
  AND2_X1 U5517 ( .A1(n8666), .A2(n8667), .ZN(n5816) );
  OR2_X1 U5518 ( .A1(n9600), .A2(n7950), .ZN(n5917) );
  NOR3_X1 U5519 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n5233) );
  NAND2_X1 U5520 ( .A1(n8231), .A2(n8243), .ZN(n8400) );
  NOR2_X1 U5521 ( .A1(n9415), .A2(n4764), .ZN(n4762) );
  OAI21_X1 U5522 ( .B1(n5831), .B2(n5830), .A(n5829), .ZN(n5847) );
  NAND2_X1 U5523 ( .A1(n4937), .A2(n5220), .ZN(n4936) );
  INV_X1 U5524 ( .A(n5720), .ZN(n4937) );
  INV_X1 U5525 ( .A(n4925), .ZN(n4924) );
  OAI21_X1 U5526 ( .B1(n4927), .B2(n4926), .A(n5618), .ZN(n4925) );
  INV_X1 U5527 ( .A(n5183), .ZN(n4926) );
  INV_X1 U5528 ( .A(n5148), .ZN(n4711) );
  AOI21_X1 U5529 ( .B1(n4956), .B2(n4954), .A(n4953), .ZN(n4952) );
  INV_X1 U5530 ( .A(n5158), .ZN(n4953) );
  INV_X1 U5531 ( .A(n5154), .ZN(n4954) );
  AOI21_X1 U5532 ( .B1(n4692), .B2(n5136), .A(n4690), .ZN(n4689) );
  INV_X1 U5533 ( .A(n5101), .ZN(n4690) );
  INV_X1 U5534 ( .A(n5140), .ZN(n4684) );
  INV_X1 U5535 ( .A(n4630), .ZN(n4628) );
  NAND2_X1 U5536 ( .A1(n4630), .A2(n4632), .ZN(n4627) );
  INV_X1 U5537 ( .A(n5126), .ZN(n4931) );
  INV_X1 U5538 ( .A(n6845), .ZN(n4615) );
  INV_X1 U5539 ( .A(n8439), .ZN(n4596) );
  XNOR2_X1 U5540 ( .A(n8906), .B(n5724), .ZN(n5617) );
  NOR4_X1 U5541 ( .A1(n6010), .A2(n6009), .A3(n8626), .A4(n6008), .ZN(n6011)
         );
  OR2_X1 U5542 ( .A1(n5420), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5477) );
  INV_X1 U5543 ( .A(n4677), .ZN(n4675) );
  NOR2_X1 U5544 ( .A1(n8623), .A2(n4517), .ZN(n4893) );
  NAND2_X1 U5545 ( .A1(n4907), .A2(n4909), .ZN(n4906) );
  NAND2_X1 U5546 ( .A1(n8020), .A2(n4864), .ZN(n4863) );
  INV_X1 U5547 ( .A(n7939), .ZN(n4864) );
  NOR2_X1 U5548 ( .A1(n4670), .A2(n4669), .ZN(n4668) );
  INV_X1 U5549 ( .A(n7652), .ZN(n4859) );
  NOR2_X1 U5550 ( .A1(n7909), .A2(n7776), .ZN(n4787) );
  INV_X1 U5551 ( .A(n7542), .ZN(n4869) );
  INV_X1 U5552 ( .A(n4870), .ZN(n4866) );
  INV_X1 U5553 ( .A(n5893), .ZN(n7603) );
  AND2_X1 U5554 ( .A1(n5998), .A2(n7280), .ZN(n5882) );
  NAND2_X1 U5555 ( .A1(n8775), .A2(n4788), .ZN(n8716) );
  NOR2_X1 U5556 ( .A1(n8617), .A2(n4789), .ZN(n4788) );
  INV_X1 U5557 ( .A(n4790), .ZN(n4789) );
  INV_X1 U5558 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5265) );
  NAND2_X1 U5559 ( .A1(n5235), .A2(n4857), .ZN(n5015) );
  INV_X1 U5560 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5773) );
  INV_X1 U5561 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5042) );
  INV_X1 U5562 ( .A(n9090), .ZN(n4727) );
  NAND2_X1 U5563 ( .A1(n4969), .A2(n4744), .ZN(n4743) );
  INV_X1 U5564 ( .A(n4518), .ZN(n4744) );
  INV_X1 U5565 ( .A(n9071), .ZN(n4737) );
  INV_X1 U5566 ( .A(n4743), .ZN(n4741) );
  NAND2_X1 U5567 ( .A1(n4505), .A2(n9027), .ZN(n4742) );
  MUX2_X1 U5568 ( .A(n8267), .B(n8259), .S(n9189), .Z(n8261) );
  AND2_X1 U5569 ( .A1(n8407), .A2(n8263), .ZN(n4917) );
  OR2_X1 U5570 ( .A1(n8266), .A2(n8265), .ZN(n4919) );
  NAND2_X1 U5571 ( .A1(n6128), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6040) );
  OR2_X1 U5572 ( .A1(n9415), .A2(n6737), .ZN(n8326) );
  NAND2_X1 U5573 ( .A1(n4796), .A2(n4496), .ZN(n9274) );
  NAND2_X1 U5574 ( .A1(n5050), .A2(n6725), .ZN(n5049) );
  INV_X1 U5575 ( .A(n6724), .ZN(n5050) );
  INV_X1 U5576 ( .A(n6725), .ZN(n5051) );
  AND2_X1 U5577 ( .A1(n9376), .A2(n5058), .ZN(n5057) );
  NAND2_X1 U5578 ( .A1(n5059), .A2(n5061), .ZN(n5058) );
  INV_X1 U5579 ( .A(n5062), .ZN(n5059) );
  INV_X1 U5580 ( .A(n5061), .ZN(n5060) );
  INV_X1 U5581 ( .A(n6715), .ZN(n5044) );
  NAND2_X1 U5582 ( .A1(n9528), .A2(n4777), .ZN(n4776) );
  INV_X1 U5583 ( .A(n8178), .ZN(n4813) );
  INV_X1 U5584 ( .A(n8181), .ZN(n4810) );
  INV_X1 U5585 ( .A(n8292), .ZN(n4809) );
  OR2_X1 U5586 ( .A1(n6267), .A2(n7126), .ZN(n6287) );
  NAND2_X1 U5587 ( .A1(n4794), .A2(n4534), .ZN(n7752) );
  AND2_X1 U5588 ( .A1(n7682), .A2(n7501), .ZN(n4758) );
  NOR2_X1 U5589 ( .A1(n7840), .A2(n7625), .ZN(n4757) );
  OR2_X1 U5590 ( .A1(n9135), .A2(n7682), .ZN(n8158) );
  OR2_X1 U5591 ( .A1(n9136), .A2(n9818), .ZN(n8146) );
  AND2_X1 U5592 ( .A1(n9259), .A2(n4760), .ZN(n9206) );
  AND2_X1 U5593 ( .A1(n4762), .A2(n4761), .ZN(n4760) );
  NAND2_X1 U5594 ( .A1(n9259), .A2(n4762), .ZN(n9221) );
  NAND2_X1 U5595 ( .A1(n4942), .A2(n4940), .ZN(n5707) );
  AOI21_X1 U5596 ( .B1(n4943), .B2(n4945), .A(n4941), .ZN(n4940) );
  INV_X1 U5597 ( .A(n5210), .ZN(n4941) );
  AND2_X1 U5598 ( .A1(n5214), .A2(n5213), .ZN(n5706) );
  NOR2_X1 U5599 ( .A1(n5205), .A2(n4947), .ZN(n4946) );
  INV_X1 U5600 ( .A(n5201), .ZN(n4947) );
  NOR2_X1 U5601 ( .A1(n5106), .A2(n5190), .ZN(n5652) );
  NOR2_X1 U5602 ( .A1(n5602), .A2(n4928), .ZN(n4927) );
  INV_X1 U5603 ( .A(n5177), .ZN(n4928) );
  NAND2_X1 U5604 ( .A1(n5586), .A2(n5175), .ZN(n5178) );
  INV_X1 U5605 ( .A(SI_17_), .ZN(n5171) );
  INV_X1 U5606 ( .A(SI_16_), .ZN(n5166) );
  INV_X1 U5607 ( .A(n6152), .ZN(n5053) );
  AND2_X1 U5608 ( .A1(n6026), .A2(n6153), .ZN(n5052) );
  INV_X1 U5609 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6020) );
  INV_X1 U5610 ( .A(SI_9_), .ZN(n10418) );
  INV_X1 U5611 ( .A(SI_8_), .ZN(n10430) );
  INV_X1 U5612 ( .A(SI_22_), .ZN(n10343) );
  NAND2_X1 U5613 ( .A1(n7302), .A2(n7301), .ZN(n5035) );
  AOI21_X1 U5614 ( .B1(n8482), .B2(n4601), .A(n4600), .ZN(n4599) );
  NOR2_X1 U5615 ( .A1(n5719), .A2(n5718), .ZN(n4600) );
  NAND2_X1 U5616 ( .A1(n5035), .A2(n5033), .ZN(n7480) );
  NAND2_X1 U5617 ( .A1(n5020), .A2(n6885), .ZN(n4830) );
  OR2_X1 U5618 ( .A1(n5987), .A2(n7275), .ZN(n4831) );
  AND2_X1 U5619 ( .A1(n5983), .A2(n4635), .ZN(n5984) );
  AND3_X1 U5620 ( .A1(n5837), .A2(n5836), .A3(n5835), .ZN(n6854) );
  AND3_X1 U5621 ( .A1(n5596), .A2(n5595), .A3(n5594), .ZN(n8610) );
  INV_X1 U5622 ( .A(n4784), .ZN(n4782) );
  INV_X1 U5623 ( .A(n5961), .ZN(n8667) );
  AND2_X1 U5624 ( .A1(n5735), .A2(n5711), .ZN(n8681) );
  NOR2_X1 U5625 ( .A1(n8782), .A2(n5001), .ZN(n5000) );
  NAND2_X1 U5626 ( .A1(n8775), .A2(n8770), .ZN(n8764) );
  NAND2_X1 U5627 ( .A1(n8775), .A2(n4792), .ZN(n8740) );
  NAND2_X1 U5628 ( .A1(n5261), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5640) );
  OR2_X1 U5629 ( .A1(n5640), .A2(n8471), .ZN(n5660) );
  NOR2_X1 U5630 ( .A1(n8906), .A2(n8807), .ZN(n8774) );
  AND2_X1 U5631 ( .A1(n8780), .A2(n8774), .ZN(n8775) );
  AND2_X1 U5632 ( .A1(n8609), .A2(n8831), .ZN(n8806) );
  NOR2_X1 U5633 ( .A1(n8914), .A2(n8546), .ZN(n4914) );
  NAND2_X1 U5634 ( .A1(n5259), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5573) );
  OR2_X1 U5635 ( .A1(n8025), .A2(n8026), .ZN(n5013) );
  INV_X1 U5636 ( .A(n8827), .ZN(n4912) );
  AND2_X1 U5637 ( .A1(n7613), .A2(n9997), .ZN(n7732) );
  NAND2_X1 U5638 ( .A1(n7732), .A2(n4787), .ZN(n7880) );
  AND2_X1 U5639 ( .A1(n7730), .A2(n7727), .ZN(n4861) );
  NAND2_X1 U5640 ( .A1(n7649), .A2(n7652), .ZN(n7728) );
  INV_X1 U5641 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10102) );
  AND4_X1 U5642 ( .A1(n5429), .A2(n5428), .A3(n5427), .A4(n5426), .ZN(n7601)
         );
  OR2_X1 U5643 ( .A1(n5424), .A2(n5423), .ZN(n5441) );
  AND2_X1 U5644 ( .A1(n5992), .A2(n7603), .ZN(n7546) );
  AND4_X1 U5645 ( .A1(n5446), .A2(n5445), .A3(n5444), .A4(n5443), .ZN(n7772)
         );
  NAND2_X1 U5646 ( .A1(n7407), .A2(n4529), .ZN(n9919) );
  AND4_X1 U5647 ( .A1(n5414), .A2(n5413), .A3(n5412), .A4(n5411), .ZN(n7548)
         );
  NAND2_X1 U5648 ( .A1(n4780), .A2(n9966), .ZN(n7425) );
  INV_X1 U5649 ( .A(n7442), .ZN(n4780) );
  NOR2_X1 U5650 ( .A1(n7425), .A2(n7431), .ZN(n7426) );
  AND2_X1 U5651 ( .A1(n5884), .A2(n5887), .ZN(n7424) );
  NAND2_X1 U5652 ( .A1(n8559), .A2(n9958), .ZN(n7280) );
  NAND2_X1 U5653 ( .A1(n4512), .A2(n9958), .ZN(n7442) );
  INV_X1 U5654 ( .A(n7440), .ZN(n5810) );
  NAND2_X1 U5655 ( .A1(n7163), .A2(n7160), .ZN(n5808) );
  NAND2_X1 U5656 ( .A1(n7280), .A2(n5864), .ZN(n7440) );
  OR2_X1 U5657 ( .A1(n4662), .A2(n8513), .ZN(n5342) );
  OR2_X1 U5658 ( .A1(n5843), .A2(n6934), .ZN(n5341) );
  AND2_X1 U5659 ( .A1(n9937), .A2(n9941), .ZN(n5760) );
  AND2_X1 U5660 ( .A1(n7877), .A2(n8939), .ZN(n8934) );
  AND2_X1 U5661 ( .A1(n5480), .A2(n5479), .ZN(n10012) );
  INV_X1 U5662 ( .A(n8455), .ZN(n7467) );
  AND2_X1 U5663 ( .A1(n9947), .A2(n5791), .ZN(n8930) );
  AND2_X1 U5664 ( .A1(n5867), .A2(n5993), .ZN(n7331) );
  OR2_X1 U5665 ( .A1(n5297), .A2(n6837), .ZN(n5301) );
  INV_X1 U5666 ( .A(n8930), .ZN(n10011) );
  NOR2_X1 U5667 ( .A1(n6878), .A2(n6877), .ZN(n7063) );
  XNOR2_X1 U5668 ( .A(n5754), .B(P2_IR_REG_26__SCAN_IN), .ZN(n5761) );
  INV_X1 U5669 ( .A(n5755), .ZN(n5756) );
  NAND2_X1 U5670 ( .A1(n5249), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5248) );
  NOR2_X1 U5671 ( .A1(n4514), .A2(n4575), .ZN(n4981) );
  INV_X1 U5672 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7126) );
  AND2_X1 U5673 ( .A1(n6448), .A2(n4727), .ZN(n4726) );
  NAND2_X1 U5674 ( .A1(n9111), .A2(n6383), .ZN(n4993) );
  XNOR2_X1 U5675 ( .A(n4756), .B(n7492), .ZN(n7308) );
  NAND2_X1 U5676 ( .A1(n6184), .A2(n6183), .ZN(n4756) );
  NAND2_X1 U5677 ( .A1(n6391), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6414) );
  INV_X1 U5678 ( .A(n6392), .ZN(n6391) );
  NAND2_X1 U5679 ( .A1(n9042), .A2(n6408), .ZN(n9052) );
  NAND2_X1 U5680 ( .A1(n6528), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6546) );
  INV_X1 U5681 ( .A(n6529), .ZN(n6528) );
  NAND2_X1 U5682 ( .A1(n4980), .A2(n6559), .ZN(n9059) );
  XNOR2_X1 U5683 ( .A(n6138), .B(n7492), .ZN(n6140) );
  NAND2_X1 U5684 ( .A1(n7795), .A2(n4966), .ZN(n4964) );
  NAND2_X1 U5685 ( .A1(n6226), .A2(n4490), .ZN(n4734) );
  OR2_X1 U5686 ( .A1(n6455), .A2(n6454), .ZN(n6479) );
  INV_X1 U5687 ( .A(n4974), .ZN(n4973) );
  OAI21_X1 U5688 ( .B1(n6472), .B2(n4975), .A(n9069), .ZN(n4974) );
  OR2_X1 U5689 ( .A1(n6332), .A2(n6331), .ZN(n6352) );
  OR2_X1 U5690 ( .A1(n6804), .A2(n6160), .ZN(n6098) );
  INV_X1 U5691 ( .A(n9058), .ZN(n4980) );
  NAND2_X1 U5692 ( .A1(n9035), .A2(n4979), .ZN(n4978) );
  INV_X1 U5693 ( .A(n6562), .ZN(n4979) );
  NAND2_X1 U5694 ( .A1(n6350), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6373) );
  INV_X1 U5695 ( .A(n6352), .ZN(n6350) );
  INV_X1 U5696 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6372) );
  OR2_X1 U5697 ( .A1(n8426), .A2(n4593), .ZN(n4915) );
  AND2_X1 U5698 ( .A1(n5064), .A2(n6063), .ZN(n5063) );
  AND2_X1 U5699 ( .A1(n6029), .A2(n6022), .ZN(n4745) );
  OR2_X1 U5700 ( .A1(n6501), .A2(n7018), .ZN(n6131) );
  OR2_X1 U5701 ( .A1(n6216), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n6227) );
  NOR2_X1 U5702 ( .A1(n7066), .A2(n4714), .ZN(n7024) );
  AND2_X1 U5703 ( .A1(n7023), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4714) );
  NAND2_X1 U5704 ( .A1(n7024), .A2(n7025), .ZN(n7049) );
  NAND2_X1 U5705 ( .A1(n7049), .A2(n4713), .ZN(n9719) );
  OR2_X1 U5706 ( .A1(n7050), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4713) );
  NAND2_X1 U5707 ( .A1(n9719), .A2(n9718), .ZN(n9717) );
  AND2_X1 U5708 ( .A1(n4716), .A2(n4715), .ZN(n7056) );
  NAND2_X1 U5709 ( .A1(n7055), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4715) );
  NAND2_X1 U5710 ( .A1(n7056), .A2(n7057), .ZN(n7713) );
  NOR2_X1 U5711 ( .A1(n9729), .A2(n4718), .ZN(n9744) );
  AND2_X1 U5712 ( .A1(n9734), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4718) );
  INV_X1 U5713 ( .A(n7716), .ZN(n9140) );
  NOR2_X1 U5714 ( .A1(n9776), .A2(n4721), .ZN(n9793) );
  AND2_X1 U5715 ( .A1(n9781), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4721) );
  NOR2_X1 U5716 ( .A1(n9793), .A2(n9792), .ZN(n9791) );
  XNOR2_X1 U5717 ( .A(n4719), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9166) );
  OR2_X1 U5718 ( .A1(n9791), .A2(n4720), .ZN(n4719) );
  AND2_X1 U5719 ( .A1(n9797), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4720) );
  AND2_X1 U5720 ( .A1(n9189), .A2(n9206), .ZN(n9179) );
  AND2_X1 U5721 ( .A1(n8326), .A2(n8325), .ZN(n9215) );
  AND2_X1 U5722 ( .A1(n8270), .A2(n8324), .ZN(n9229) );
  OAI21_X1 U5723 ( .B1(n9250), .B2(n6755), .A(n8269), .ZN(n9231) );
  NAND2_X1 U5724 ( .A1(n9264), .A2(n8234), .ZN(n9250) );
  NAND2_X1 U5725 ( .A1(n9259), .A2(n9249), .ZN(n9244) );
  NAND2_X1 U5726 ( .A1(n5065), .A2(n5066), .ZN(n9243) );
  AOI21_X1 U5727 ( .B1(n5067), .B2(n5074), .A(n4547), .ZN(n5066) );
  NAND2_X1 U5728 ( .A1(n9266), .A2(n9265), .ZN(n9264) );
  NOR2_X1 U5729 ( .A1(n9283), .A2(n9428), .ZN(n9259) );
  OR2_X1 U5730 ( .A1(n6495), .A2(n9029), .ZN(n6513) );
  AND2_X1 U5731 ( .A1(n9339), .A2(n4561), .ZN(n9295) );
  INV_X1 U5732 ( .A(n9438), .ZN(n4769) );
  NAND2_X1 U5733 ( .A1(n9339), .A2(n4770), .ZN(n9314) );
  NAND2_X1 U5734 ( .A1(n6752), .A2(n9347), .ZN(n9352) );
  AOI21_X1 U5735 ( .B1(n4819), .B2(n8315), .A(n4816), .ZN(n4815) );
  INV_X1 U5736 ( .A(n8315), .ZN(n4817) );
  NAND2_X1 U5737 ( .A1(n9339), .A2(n9346), .ZN(n9340) );
  NAND2_X1 U5738 ( .A1(n6434), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6455) );
  INV_X1 U5739 ( .A(n6436), .ZN(n6434) );
  NAND2_X1 U5740 ( .A1(n6751), .A2(n4818), .ZN(n8096) );
  AND2_X1 U5741 ( .A1(n9360), .A2(n8093), .ZN(n9339) );
  NOR2_X1 U5742 ( .A1(n9388), .A2(n9465), .ZN(n9360) );
  INV_X1 U5743 ( .A(n9364), .ZN(n9359) );
  NAND2_X1 U5744 ( .A1(n4773), .A2(n4774), .ZN(n9618) );
  NOR2_X1 U5745 ( .A1(n6770), .A2(n4776), .ZN(n4774) );
  INV_X1 U5746 ( .A(n4805), .ZN(n4804) );
  AOI21_X1 U5747 ( .B1(n4805), .B2(n4803), .A(n4802), .ZN(n4801) );
  INV_X1 U5748 ( .A(n8173), .ZN(n4802) );
  NOR2_X1 U5749 ( .A1(n7981), .A2(n4776), .ZN(n9619) );
  NOR2_X1 U5750 ( .A1(n7981), .A2(n8167), .ZN(n8012) );
  OAI21_X1 U5751 ( .B1(n7852), .B2(n4811), .A(n4808), .ZN(n9643) );
  INV_X1 U5752 ( .A(n4812), .ZN(n4811) );
  AOI21_X1 U5753 ( .B1(n4812), .B2(n4810), .A(n4809), .ZN(n4808) );
  NOR2_X1 U5754 ( .A1(n7806), .A2(n4813), .ZN(n4812) );
  OAI21_X1 U5755 ( .B1(n7851), .B2(n5081), .A(n5078), .ZN(n9635) );
  OR2_X1 U5756 ( .A1(n9825), .A2(n9132), .ZN(n5083) );
  NAND2_X1 U5757 ( .A1(n4814), .A2(n8178), .ZN(n7807) );
  NAND2_X1 U5758 ( .A1(n7852), .A2(n8181), .ZN(n4814) );
  INV_X1 U5759 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6248) );
  OR2_X1 U5760 ( .A1(n6249), .A2(n6248), .ZN(n6267) );
  AND2_X1 U5761 ( .A1(n8169), .A2(n8178), .ZN(n8352) );
  INV_X1 U5762 ( .A(n9131), .ZN(n9645) );
  AND2_X1 U5763 ( .A1(n8164), .A2(n8276), .ZN(n8351) );
  AND2_X1 U5764 ( .A1(n7501), .A2(n7682), .ZN(n7680) );
  XNOR2_X1 U5765 ( .A(n6701), .B(n9811), .ZN(n8343) );
  NOR2_X1 U5766 ( .A1(n7376), .A2(n4479), .ZN(n7695) );
  NAND2_X1 U5767 ( .A1(n6741), .A2(n7188), .ZN(n7187) );
  MUX2_X1 U5768 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8962), .S(n8129), .Z(n8131) );
  NAND2_X1 U5769 ( .A1(n8136), .A2(n8135), .ZN(n9180) );
  NAND2_X1 U5770 ( .A1(n6751), .A2(n8306), .ZN(n9365) );
  OR2_X1 U5771 ( .A1(n9488), .A2(n6678), .ZN(n9826) );
  OR2_X1 U5772 ( .A1(n9488), .A2(n8417), .ZN(n9827) );
  INV_X1 U5773 ( .A(n9827), .ZN(n9467) );
  OR2_X1 U5774 ( .A1(n8267), .A2(n8417), .ZN(n7845) );
  NOR2_X1 U5775 ( .A1(n6782), .A2(n7151), .ZN(n7491) );
  NAND2_X1 U5776 ( .A1(n9652), .A2(n7845), .ZN(n9822) );
  NAND2_X1 U5777 ( .A1(n6651), .A2(n6650), .ZN(n7490) );
  XNOR2_X1 U5778 ( .A(n5845), .B(SI_30_), .ZN(n8133) );
  XNOR2_X1 U5779 ( .A(n5831), .B(n5823), .ZN(n8082) );
  XNOR2_X1 U5780 ( .A(n5243), .B(n5242), .ZN(n7989) );
  NAND2_X1 U5781 ( .A1(n5676), .A2(n5201), .ZN(n5243) );
  NAND2_X1 U5782 ( .A1(n5656), .A2(n5195), .ZN(n5673) );
  XNOR2_X1 U5783 ( .A(n6079), .B(P1_IR_REG_19__SCAN_IN), .ZN(n9317) );
  NAND2_X1 U5784 ( .A1(n6409), .A2(n5098), .ZN(n6078) );
  XNOR2_X1 U5785 ( .A(n4681), .B(n5602), .ZN(n7669) );
  NAND2_X1 U5786 ( .A1(n5178), .A2(n5177), .ZN(n4681) );
  NAND2_X1 U5787 ( .A1(n4706), .A2(n4708), .ZN(n5511) );
  OR2_X1 U5788 ( .A1(n5145), .A2(n4712), .ZN(n4706) );
  OAI21_X1 U5789 ( .B1(n5472), .B2(n5471), .A(n5154), .ZN(n5493) );
  OR2_X1 U5790 ( .A1(n6304), .A2(n6303), .ZN(n6327) );
  INV_X1 U5791 ( .A(n4687), .ZN(n5419) );
  INV_X1 U5792 ( .A(n4692), .ZN(n4688) );
  NAND2_X1 U5793 ( .A1(n6022), .A2(n6021), .ZN(n6152) );
  NAND2_X1 U5794 ( .A1(n5035), .A2(n5379), .ZN(n7389) );
  AND2_X1 U5795 ( .A1(n5742), .A2(n5741), .ZN(n8671) );
  NAND2_X1 U5796 ( .A1(n5723), .A2(n5722), .ZN(n8861) );
  AND2_X1 U5797 ( .A1(n9598), .A2(n5509), .ZN(n5037) );
  AND2_X1 U5798 ( .A1(n5038), .A2(n5509), .ZN(n9599) );
  NAND2_X1 U5799 ( .A1(n5679), .A2(n5678), .ZN(n8883) );
  NAND2_X1 U5800 ( .A1(n7572), .A2(n5435), .ZN(n7825) );
  INV_X1 U5801 ( .A(n8457), .ZN(n4619) );
  NAND2_X1 U5802 ( .A1(n7232), .A2(n5323), .ZN(n8458) );
  INV_X1 U5803 ( .A(n5635), .ZN(n4682) );
  INV_X1 U5804 ( .A(n5634), .ZN(n8466) );
  AND4_X1 U5805 ( .A1(n5465), .A2(n5464), .A3(n5463), .A4(n5462), .ZN(n7899)
         );
  INV_X1 U5806 ( .A(n10012), .ZN(n7909) );
  NAND2_X1 U5807 ( .A1(n5693), .A2(n5692), .ZN(n8873) );
  AOI21_X1 U5808 ( .B1(n4696), .B2(n4697), .A(n4555), .ZN(n4695) );
  AND2_X1 U5809 ( .A1(n5583), .A2(n5565), .ZN(n5027) );
  NAND2_X1 U5810 ( .A1(n5028), .A2(n5565), .ZN(n8045) );
  NOR2_X1 U5811 ( .A1(n4703), .A2(n4702), .ZN(n8493) );
  NAND2_X1 U5812 ( .A1(n4558), .A2(n5029), .ZN(n4605) );
  INV_X1 U5813 ( .A(n5029), .ZN(n4606) );
  MUX2_X1 U5814 ( .A(n5286), .B(n8984), .S(n5313), .Z(n7203) );
  NAND2_X1 U5815 ( .A1(n5287), .A2(n7337), .ZN(n7205) );
  NAND2_X1 U5816 ( .A1(n9606), .A2(n8750), .ZN(n8526) );
  NAND2_X1 U5817 ( .A1(n5659), .A2(n5658), .ZN(n8889) );
  AND3_X1 U5818 ( .A1(n5318), .A2(n5317), .A3(n5316), .ZN(n9952) );
  NAND2_X1 U5819 ( .A1(n5591), .A2(n5590), .ZN(n8909) );
  NAND2_X1 U5820 ( .A1(n4608), .A2(n4609), .ZN(n7302) );
  OAI21_X1 U5821 ( .B1(n8487), .B2(n8482), .A(n8486), .ZN(n8534) );
  NAND2_X1 U5822 ( .A1(n5795), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9616) );
  INV_X1 U5823 ( .A(n8481), .ZN(n9606) );
  NAND2_X1 U5824 ( .A1(n5558), .A2(n5557), .ZN(n9609) );
  AND2_X1 U5825 ( .A1(n5799), .A2(n5798), .ZN(n8750) );
  INV_X1 U5826 ( .A(n8763), .ZN(n8616) );
  AND3_X1 U5827 ( .A1(n5612), .A2(n5611), .A3(n5610), .ZN(n8821) );
  NAND4_X1 U5828 ( .A1(n5363), .A2(n5362), .A3(n5361), .A4(n5360), .ZN(n8558)
         );
  INV_X1 U5829 ( .A(n5809), .ZN(n8559) );
  NAND2_X1 U5830 ( .A1(n5328), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5308) );
  NAND4_X1 U5831 ( .A1(n5281), .A2(n5280), .A3(n5279), .A4(n5278), .ZN(n8561)
         );
  INV_X2 U5832 ( .A(P2_U3966), .ZN(n8560) );
  NAND2_X1 U5833 ( .A1(n5853), .A2(n5852), .ZN(n8844) );
  XNOR2_X1 U5834 ( .A(n8848), .B(n8844), .ZN(n8846) );
  NAND2_X1 U5835 ( .A1(n8661), .A2(n4783), .ZN(n8848) );
  NOR2_X1 U5836 ( .A1(n5839), .A2(n4784), .ZN(n4783) );
  AOI21_X1 U5837 ( .B1(n8634), .B2(n8795), .A(n8633), .ZN(n8855) );
  NAND2_X1 U5838 ( .A1(n4889), .A2(n4886), .ZN(n8625) );
  INV_X1 U5839 ( .A(n4887), .ZN(n4886) );
  NAND2_X1 U5840 ( .A1(n5004), .A2(n5005), .ZN(n8650) );
  NAND2_X1 U5841 ( .A1(n4891), .A2(n4898), .ZN(n8642) );
  NAND2_X1 U5842 ( .A1(n4901), .A2(n4517), .ZN(n4891) );
  NAND2_X1 U5843 ( .A1(n4901), .A2(n4900), .ZN(n8660) );
  AOI21_X1 U5844 ( .B1(n8695), .B2(n8621), .A(n4513), .ZN(n8677) );
  NAND2_X1 U5845 ( .A1(n4876), .A2(n4877), .ZN(n8735) );
  AOI21_X1 U5846 ( .B1(n8758), .B2(n8615), .A(n4884), .ZN(n8739) );
  NAND2_X1 U5847 ( .A1(n8786), .A2(n5944), .ZN(n8759) );
  NAND2_X1 U5848 ( .A1(n8827), .A2(n4905), .ZN(n4904) );
  INV_X1 U5849 ( .A(n4909), .ZN(n4905) );
  NAND2_X1 U5850 ( .A1(n5533), .A2(n5532), .ZN(n8064) );
  OAI21_X1 U5851 ( .B1(n7872), .B2(n4665), .A(n4664), .ZN(n7948) );
  NAND2_X1 U5852 ( .A1(n8839), .A2(n7276), .ZN(n8813) );
  NAND2_X1 U5853 ( .A1(n7940), .A2(n7939), .ZN(n8021) );
  AND2_X1 U5854 ( .A1(n7923), .A2(n7922), .ZN(n7925) );
  NAND2_X1 U5855 ( .A1(n4672), .A2(n4671), .ZN(n7919) );
  NAND2_X1 U5856 ( .A1(n9938), .A2(n7269), .ZN(n8836) );
  NAND2_X1 U5857 ( .A1(n4633), .A2(n5408), .ZN(n9927) );
  NAND2_X1 U5858 ( .A1(n6865), .A2(n4616), .ZN(n4633) );
  NAND2_X1 U5859 ( .A1(n7543), .A2(n7542), .ZN(n9914) );
  AND2_X1 U5860 ( .A1(n7421), .A2(n7402), .ZN(n7404) );
  INV_X1 U5861 ( .A(n7141), .ZN(n7352) );
  NAND2_X1 U5862 ( .A1(n8839), .A2(n7271), .ZN(n8843) );
  INV_X1 U5863 ( .A(n8813), .ZN(n9926) );
  INV_X1 U5864 ( .A(n8717), .ZN(n9932) );
  AND2_X2 U5865 ( .A1(n7063), .A2(n7267), .ZN(n10021) );
  AND2_X1 U5866 ( .A1(n6015), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9945) );
  NAND2_X1 U5867 ( .A1(n9939), .A2(n9938), .ZN(n9942) );
  INV_X1 U5868 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8964) );
  INV_X1 U5869 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5269) );
  NAND2_X1 U5870 ( .A1(n5268), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5270) );
  NAND2_X1 U5871 ( .A1(n4853), .A2(n4654), .ZN(n5268) );
  NAND2_X1 U5872 ( .A1(n5239), .A2(n5238), .ZN(n8977) );
  MUX2_X1 U5873 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5237), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5239) );
  NAND2_X1 U5874 ( .A1(n4618), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5237) );
  INV_X1 U5875 ( .A(n5761), .ZN(n8982) );
  INV_X1 U5876 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7990) );
  NAND2_X1 U5877 ( .A1(n5776), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5752) );
  INV_X1 U5878 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7781) );
  INV_X1 U5879 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7740) );
  XNOR2_X1 U5880 ( .A(n5256), .B(n5255), .ZN(n7741) );
  INV_X1 U5881 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7671) );
  OR2_X1 U5882 ( .A1(n5252), .A2(n5251), .ZN(n5253) );
  INV_X1 U5883 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7260) );
  INV_X1 U5884 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7184) );
  INV_X1 U5885 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7175) );
  INV_X1 U5886 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7137) );
  INV_X1 U5887 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6874) );
  INV_X1 U5888 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6870) );
  NOR2_X1 U5889 ( .A1(n6800), .A2(n7956), .ZN(n6808) );
  INV_X1 U5890 ( .A(n4752), .ZN(n4751) );
  AOI21_X1 U5891 ( .B1(n4750), .B2(n4752), .A(n4557), .ZN(n4749) );
  OR2_X1 U5892 ( .A1(n7522), .A2(n4753), .ZN(n4752) );
  INV_X1 U5893 ( .A(n9217), .ZN(n8993) );
  NAND2_X1 U5894 ( .A1(n6527), .A2(n6526), .ZN(n9286) );
  INV_X1 U5895 ( .A(n4729), .ZN(n4728) );
  OAI21_X1 U5896 ( .B1(n4731), .B2(n4490), .A(n6262), .ZN(n4729) );
  NAND2_X1 U5897 ( .A1(n6265), .A2(n6264), .ZN(n7895) );
  OAI21_X1 U5898 ( .B1(n6447), .B2(n4726), .A(n4725), .ZN(n9021) );
  NAND2_X1 U5899 ( .A1(n4967), .A2(n6243), .ZN(n7794) );
  INV_X1 U5900 ( .A(n6100), .ZN(n7241) );
  NAND2_X1 U5901 ( .A1(n6307), .A2(n6306), .ZN(n7999) );
  NAND2_X1 U5902 ( .A1(n9059), .A2(n6562), .ZN(n9034) );
  NAND2_X1 U5903 ( .A1(n6564), .A2(n6563), .ZN(n9423) );
  NAND2_X1 U5904 ( .A1(n4993), .A2(n6386), .ZN(n9045) );
  NAND2_X1 U5905 ( .A1(n6390), .A2(n6389), .ZN(n9390) );
  NAND2_X1 U5906 ( .A1(n7319), .A2(n6169), .ZN(n4961) );
  NAND2_X1 U5907 ( .A1(n9019), .A2(n6473), .ZN(n9068) );
  NAND2_X1 U5908 ( .A1(n7993), .A2(n6326), .ZN(n8038) );
  NAND2_X1 U5909 ( .A1(n6510), .A2(n4518), .ZN(n9079) );
  NAND2_X1 U5910 ( .A1(n6510), .A2(n6509), .ZN(n4971) );
  XNOR2_X1 U5911 ( .A(n6524), .B(n7492), .ZN(n9081) );
  NAND2_X1 U5912 ( .A1(n6283), .A2(n6282), .ZN(n7935) );
  NAND2_X1 U5913 ( .A1(n6447), .A2(n6448), .ZN(n9088) );
  NAND2_X1 U5914 ( .A1(n6433), .A2(n6432), .ZN(n9462) );
  NAND2_X1 U5915 ( .A1(n4958), .A2(n6189), .ZN(n7524) );
  INV_X1 U5916 ( .A(n9120), .ZN(n9105) );
  AND2_X1 U5917 ( .A1(n6686), .A2(n9687), .ZN(n9120) );
  AND2_X1 U5918 ( .A1(n6671), .A2(n6680), .ZN(n9115) );
  OR2_X1 U5919 ( .A1(n6673), .A2(n6672), .ZN(n8431) );
  XNOR2_X1 U5920 ( .A(n6077), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8433) );
  OR3_X1 U5921 ( .A1(n7179), .A2(n7178), .A3(n7177), .ZN(n9175) );
  NAND2_X1 U5922 ( .A1(n6609), .A2(n6608), .ZN(n9233) );
  NAND2_X1 U5923 ( .A1(n6573), .A2(n6572), .ZN(n9267) );
  OR2_X1 U5924 ( .A1(n6127), .A2(n6961), .ZN(n6113) );
  CLKBUF_X1 U5925 ( .A(n6695), .Z(n9139) );
  INV_X1 U5926 ( .A(n4716), .ZN(n7129) );
  AOI21_X1 U5927 ( .B1(n5085), .B2(n5090), .A(n5094), .ZN(n5084) );
  AND2_X1 U5928 ( .A1(n5088), .A2(n5085), .ZN(n9196) );
  NAND2_X1 U5929 ( .A1(n5088), .A2(n5089), .ZN(n9194) );
  NAND2_X1 U5930 ( .A1(n5068), .A2(n5071), .ZN(n9257) );
  NAND2_X1 U5931 ( .A1(n9294), .A2(n5069), .ZN(n5068) );
  NAND2_X1 U5932 ( .A1(n5070), .A2(n6729), .ZN(n9272) );
  NAND2_X1 U5933 ( .A1(n6728), .A2(n6727), .ZN(n5070) );
  NAND2_X1 U5934 ( .A1(n4796), .A2(n4797), .ZN(n9300) );
  NAND2_X1 U5935 ( .A1(n5048), .A2(n6725), .ZN(n9307) );
  NAND2_X1 U5936 ( .A1(n9332), .A2(n6724), .ZN(n5048) );
  NAND2_X1 U5937 ( .A1(n6753), .A2(n8218), .ZN(n9310) );
  NAND2_X1 U5938 ( .A1(n6475), .A2(n6474), .ZN(n9449) );
  NAND2_X1 U5939 ( .A1(n5056), .A2(n5061), .ZN(n9386) );
  NAND2_X1 U5940 ( .A1(n9617), .A2(n5062), .ZN(n5056) );
  NAND2_X1 U5941 ( .A1(n5045), .A2(n6715), .ZN(n8011) );
  NAND2_X1 U5942 ( .A1(n4807), .A2(n4805), .ZN(n8008) );
  NOR2_X1 U5943 ( .A1(n7537), .A2(n9317), .ZN(n9395) );
  NAND2_X1 U5944 ( .A1(n4794), .A2(n8381), .ZN(n7565) );
  AND2_X1 U5945 ( .A1(n9395), .A2(n9467), .ZN(n9640) );
  NAND2_X1 U5946 ( .A1(n4799), .A2(n8130), .ZN(n4798) );
  OAI21_X1 U5947 ( .B1(n6837), .B2(n6835), .A(n4554), .ZN(n4799) );
  AND2_X2 U5948 ( .A1(n6778), .A2(n6783), .ZN(n9840) );
  AOI21_X1 U5949 ( .B1(n9410), .B2(n9822), .A(n9409), .ZN(n9497) );
  OR2_X1 U5950 ( .A1(n9408), .A2(n9407), .ZN(n9409) );
  INV_X1 U5951 ( .A(n9286), .ZN(n9509) );
  AND2_X1 U5952 ( .A1(n6800), .A2(n6655), .ZN(n9808) );
  XNOR2_X1 U5953 ( .A(n5820), .B(n5819), .ZN(n6615) );
  NAND2_X1 U5954 ( .A1(n4935), .A2(n5220), .ZN(n5820) );
  INV_X1 U5955 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8003) );
  INV_X1 U5956 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7914) );
  INV_X1 U5957 ( .A(n8433), .ZN(n7915) );
  INV_X1 U5958 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8087) );
  INV_X1 U5959 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10419) );
  NAND2_X1 U5960 ( .A1(n6044), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6046) );
  INV_X1 U5961 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10375) );
  INV_X1 U5962 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7185) );
  INV_X1 U5963 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10316) );
  INV_X1 U5964 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6871) );
  INV_X1 U5965 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6866) );
  XNOR2_X1 U5966 ( .A(n5365), .B(n5364), .ZN(n6853) );
  NAND2_X1 U5967 ( .A1(n4932), .A2(n5126), .ZN(n5365) );
  NAND2_X1 U5968 ( .A1(n8120), .A2(n5614), .ZN(n8128) );
  OAI21_X1 U5969 ( .B1(n5781), .B2(n9610), .A(n5025), .ZN(n5802) );
  AND2_X1 U5970 ( .A1(n6692), .A2(n4987), .ZN(n4986) );
  NAND2_X1 U5971 ( .A1(n4991), .A2(n4508), .ZN(n4987) );
  NOR2_X1 U5972 ( .A1(n4580), .A2(n4822), .ZN(n4821) );
  NAND2_X1 U5973 ( .A1(n9833), .A2(n6784), .ZN(n4767) );
  INV_X2 U5974 ( .A(n5297), .ZN(n4616) );
  AND4_X1 U5975 ( .A1(n8423), .A2(n8422), .A3(n8421), .A4(n8420), .ZN(n4488)
         );
  INV_X1 U5976 ( .A(n5234), .ZN(n4853) );
  AND2_X1 U5977 ( .A1(n4906), .A2(n8612), .ZN(n4489) );
  INV_X1 U5978 ( .A(n8026), .ZN(n5011) );
  OR2_X1 U5979 ( .A1(n5817), .A2(n8671), .ZN(n5818) );
  NAND2_X1 U5980 ( .A1(n5313), .A2(n6835), .ZN(n5297) );
  AND3_X1 U5981 ( .A1(n4592), .A2(n4748), .A3(n4745), .ZN(n6054) );
  NOR2_X1 U5982 ( .A1(n4965), .A2(n4963), .ZN(n4490) );
  OR2_X1 U5983 ( .A1(n8427), .A2(n4915), .ZN(n4491) );
  AND2_X1 U5984 ( .A1(n9309), .A2(n5049), .ZN(n4492) );
  AND2_X1 U5985 ( .A1(n4708), .A2(n5510), .ZN(n4493) );
  NOR2_X1 U5986 ( .A1(n4579), .A2(n4914), .ZN(n4494) );
  AND2_X1 U5987 ( .A1(n5144), .A2(n5453), .ZN(n4495) );
  OR2_X1 U5988 ( .A1(n8900), .A2(n8762), .ZN(n5944) );
  INV_X1 U5989 ( .A(n5944), .ZN(n4846) );
  AND2_X1 U5990 ( .A1(n4797), .A2(n4795), .ZN(n4496) );
  AND2_X1 U5991 ( .A1(n5913), .A2(n5912), .ZN(n7871) );
  INV_X1 U5992 ( .A(n7871), .ZN(n4670) );
  NAND2_X1 U5993 ( .A1(n5571), .A2(n5570), .ZN(n8914) );
  INV_X1 U5994 ( .A(n4908), .ZN(n4907) );
  OAI21_X1 U5995 ( .B1(n4909), .B2(n4911), .A(n4913), .ZN(n4908) );
  NAND2_X1 U5996 ( .A1(n9465), .A2(n9380), .ZN(n4497) );
  NOR2_X1 U5997 ( .A1(n9215), .A2(n5092), .ZN(n5091) );
  NAND2_X1 U5998 ( .A1(n6603), .A2(n6602), .ZN(n9415) );
  NAND2_X1 U5999 ( .A1(n9259), .A2(n4763), .ZN(n4766) );
  AND2_X1 U6000 ( .A1(n7935), .A2(n9130), .ZN(n4498) );
  AND3_X1 U6001 ( .A1(n5330), .A2(n5329), .A3(n5331), .ZN(n4499) );
  INV_X1 U6002 ( .A(n5074), .ZN(n5069) );
  NAND2_X1 U6003 ( .A1(n5075), .A2(n6729), .ZN(n5074) );
  AND2_X1 U6004 ( .A1(n5617), .A2(n5616), .ZN(n4500) );
  NAND2_X1 U6005 ( .A1(n6052), .A2(n6057), .ZN(n4501) );
  OR2_X1 U6006 ( .A1(n7935), .A2(n9130), .ZN(n4502) );
  AND2_X1 U6007 ( .A1(n4787), .A2(n4786), .ZN(n4503) );
  OR2_X1 U6008 ( .A1(n6447), .A2(n6448), .ZN(n4504) );
  NAND2_X1 U6009 ( .A1(n4968), .A2(n4970), .ZN(n4505) );
  INV_X1 U6010 ( .A(n8895), .ZN(n8770) );
  NAND2_X1 U6011 ( .A1(n5639), .A2(n5638), .ZN(n8895) );
  AND3_X1 U6012 ( .A1(n6030), .A2(n6043), .A3(n10403), .ZN(n4506) );
  AND3_X1 U6013 ( .A1(n5356), .A2(n5228), .A3(n4567), .ZN(n4507) );
  INV_X1 U6014 ( .A(n5688), .ZN(n4702) );
  NAND2_X1 U6015 ( .A1(n6226), .A2(n7585), .ZN(n4967) );
  OR2_X1 U6016 ( .A1(n8987), .A2(n4990), .ZN(n4508) );
  NAND2_X1 U6017 ( .A1(n7728), .A2(n4861), .ZN(n7867) );
  OR2_X1 U6018 ( .A1(n4967), .A2(n6243), .ZN(n7793) );
  NAND2_X1 U6019 ( .A1(n4672), .A2(n5912), .ZN(n4509) );
  AND2_X1 U6020 ( .A1(n9663), .A2(n4775), .ZN(n4510) );
  NAND2_X1 U6021 ( .A1(n6348), .A2(n6347), .ZN(n9007) );
  AND2_X1 U6022 ( .A1(n5819), .A2(n4936), .ZN(n4511) );
  NAND2_X1 U6023 ( .A1(n4734), .A2(n4964), .ZN(n7831) );
  AND2_X1 U6024 ( .A1(n7340), .A2(n8455), .ZN(n4512) );
  NAND2_X2 U6025 ( .A1(n5313), .A2(n8129), .ZN(n5312) );
  AND2_X1 U6026 ( .A1(n8705), .A2(n8715), .ZN(n4513) );
  AND2_X1 U6027 ( .A1(n4680), .A2(n5271), .ZN(n5328) );
  AND2_X1 U6028 ( .A1(n6345), .A2(n6344), .ZN(n4514) );
  OR2_X1 U6029 ( .A1(n8770), .A2(n8749), .ZN(n4515) );
  NAND4_X1 U6030 ( .A1(n5309), .A2(n5308), .A3(n5307), .A4(n5306), .ZN(n5806)
         );
  XNOR2_X1 U6031 ( .A(n8914), .B(n8546), .ZN(n8828) );
  INV_X1 U6032 ( .A(n8828), .ZN(n4911) );
  NOR2_X2 U6033 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6067) );
  INV_X1 U6034 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9536) );
  AND2_X1 U6035 ( .A1(n7924), .A2(n7922), .ZN(n4516) );
  AND2_X1 U6036 ( .A1(n4899), .A2(n4900), .ZN(n4517) );
  AND2_X1 U6037 ( .A1(n6509), .A2(n4970), .ZN(n4518) );
  AND3_X1 U6038 ( .A1(n4515), .A2(n5981), .A3(n5946), .ZN(n4519) );
  AND2_X1 U6039 ( .A1(n4851), .A2(n4853), .ZN(n5266) );
  AND3_X1 U6040 ( .A1(n6131), .A2(n6130), .A3(n6129), .ZN(n4520) );
  AND2_X1 U6041 ( .A1(n5364), .A2(n5353), .ZN(n4521) );
  INV_X1 U6042 ( .A(n5081), .ZN(n5080) );
  NAND2_X1 U6043 ( .A1(n7806), .A2(n5082), .ZN(n5081) );
  NOR2_X1 U6044 ( .A1(n6152), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6178) );
  AND2_X1 U6045 ( .A1(n5053), .A2(n5052), .ZN(n4522) );
  AND2_X1 U6046 ( .A1(n8085), .A2(n5271), .ZN(n5289) );
  OR3_X1 U6047 ( .A1(n8426), .A2(n8433), .A3(n8132), .ZN(n4523) );
  INV_X1 U6048 ( .A(n8138), .ZN(n9172) );
  OR2_X1 U6049 ( .A1(n5948), .A2(n5981), .ZN(n4524) );
  OR2_X1 U6050 ( .A1(n8914), .A2(n8819), .ZN(n4525) );
  XNOR2_X1 U6051 ( .A(n5721), .B(n5720), .ZN(n6601) );
  AND4_X1 U6052 ( .A1(n6428), .A2(n6076), .A3(n6073), .A4(n6044), .ZN(n4526)
         );
  NAND2_X1 U6053 ( .A1(n6036), .A2(n9542), .ZN(n6127) );
  AND2_X1 U6054 ( .A1(n6559), .A2(n9035), .ZN(n4527) );
  AND2_X1 U6055 ( .A1(n8374), .A2(n8267), .ZN(n4528) );
  NAND2_X1 U6056 ( .A1(n6452), .A2(n6451), .ZN(n9455) );
  AND2_X1 U6057 ( .A1(n5811), .A2(n5891), .ZN(n4529) );
  NAND2_X1 U6058 ( .A1(n4735), .A2(n4740), .ZN(n9010) );
  NOR2_X1 U6059 ( .A1(n9007), .A2(n9127), .ZN(n4530) );
  AND2_X1 U6060 ( .A1(n9184), .A2(n9822), .ZN(n4531) );
  AND2_X1 U6061 ( .A1(n5358), .A2(n5357), .ZN(n9966) );
  AND2_X1 U6062 ( .A1(n5245), .A2(n5244), .ZN(n8876) );
  INV_X1 U6063 ( .A(n8727), .ZN(n8734) );
  AND2_X1 U6064 ( .A1(n7232), .A2(n5323), .ZN(n4532) );
  AND2_X1 U6065 ( .A1(n5815), .A2(n5957), .ZN(n8697) );
  NOR2_X1 U6066 ( .A1(n9465), .A2(n9380), .ZN(n4533) );
  INV_X1 U6067 ( .A(n5104), .ZN(n4679) );
  AND2_X1 U6068 ( .A1(n5818), .A2(n5971), .ZN(n8623) );
  AND2_X1 U6069 ( .A1(n4793), .A2(n8381), .ZN(n4534) );
  AND2_X1 U6070 ( .A1(n5944), .A2(n5940), .ZN(n8613) );
  INV_X1 U6071 ( .A(n8613), .ZN(n8782) );
  AND2_X1 U6072 ( .A1(n5943), .A2(n4635), .ZN(n4535) );
  INV_X1 U6073 ( .A(n8341), .ZN(n4795) );
  INV_X1 U6074 ( .A(n5072), .ZN(n5071) );
  OAI21_X1 U6075 ( .B1(n6731), .B2(n5073), .A(n6730), .ZN(n5072) );
  OAI21_X1 U6076 ( .B1(n4645), .B2(n5011), .A(n8828), .ZN(n4644) );
  AND2_X1 U6077 ( .A1(n5891), .A2(n5890), .ZN(n7408) );
  INV_X1 U6078 ( .A(n5091), .ZN(n5090) );
  INV_X1 U6079 ( .A(n5839), .ZN(n8851) );
  NAND2_X1 U6080 ( .A1(n5833), .A2(n5832), .ZN(n5839) );
  AND2_X1 U6081 ( .A1(n8786), .A2(n5002), .ZN(n4536) );
  INV_X1 U6082 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4857) );
  INV_X1 U6083 ( .A(n4896), .ZN(n4895) );
  OAI21_X1 U6084 ( .B1(n8621), .B2(n4513), .A(n4897), .ZN(n4896) );
  NOR2_X1 U6085 ( .A1(n7909), .A2(n8551), .ZN(n4537) );
  NOR2_X1 U6086 ( .A1(n7895), .A2(n9131), .ZN(n4538) );
  NOR2_X1 U6087 ( .A1(n9415), .A2(n9233), .ZN(n4539) );
  AND2_X1 U6088 ( .A1(n9927), .A2(n8555), .ZN(n4540) );
  NAND2_X1 U6089 ( .A1(n8814), .A2(n8610), .ZN(n4541) );
  AND2_X1 U6090 ( .A1(n5863), .A2(n5864), .ZN(n4542) );
  INV_X1 U6091 ( .A(n4514), .ZN(n4985) );
  AND2_X1 U6092 ( .A1(n5973), .A2(n4635), .ZN(n4543) );
  AND2_X1 U6093 ( .A1(n5128), .A2(SI_6_), .ZN(n4544) );
  AOI21_X1 U6094 ( .B1(n9028), .B2(n4739), .A(n4741), .ZN(n4738) );
  NOR2_X1 U6095 ( .A1(n5817), .A2(n8628), .ZN(n4545) );
  NAND2_X1 U6096 ( .A1(n8697), .A2(n4524), .ZN(n4546) );
  INV_X1 U6097 ( .A(n4764), .ZN(n4763) );
  NAND2_X1 U6098 ( .A1(n9249), .A2(n4765), .ZN(n4764) );
  NOR2_X1 U6099 ( .A1(n9428), .A2(n9280), .ZN(n4547) );
  INV_X1 U6100 ( .A(n4969), .ZN(n4968) );
  OR2_X1 U6101 ( .A1(n5886), .A2(n5885), .ZN(n4548) );
  INV_X1 U6102 ( .A(n6473), .ZN(n4975) );
  AND2_X1 U6103 ( .A1(n5124), .A2(SI_4_), .ZN(n4549) );
  AND2_X1 U6104 ( .A1(n5160), .A2(SI_14_), .ZN(n4550) );
  AND2_X1 U6105 ( .A1(n5081), .A2(n4502), .ZN(n4551) );
  NAND2_X1 U6106 ( .A1(n4525), .A2(n5011), .ZN(n4552) );
  AND2_X1 U6107 ( .A1(n5356), .A2(n5228), .ZN(n4553) );
  NAND2_X1 U6108 ( .A1(n6835), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4554) );
  AND2_X1 U6109 ( .A1(n4700), .A2(n4699), .ZN(n4555) );
  NOR2_X1 U6110 ( .A1(n8802), .A2(n8821), .ZN(n4556) );
  AND2_X1 U6111 ( .A1(n7522), .A2(n4753), .ZN(n4557) );
  INV_X1 U6112 ( .A(n4819), .ZN(n4818) );
  OR2_X1 U6113 ( .A1(n8139), .A2(n4820), .ZN(n4819) );
  AND2_X1 U6114 ( .A1(n4957), .A2(n5099), .ZN(n4956) );
  INV_X1 U6115 ( .A(n4698), .ZN(n4697) );
  NAND2_X1 U6116 ( .A1(n5687), .A2(n5688), .ZN(n4698) );
  INV_X1 U6117 ( .A(n4875), .ZN(n4874) );
  NAND2_X1 U6118 ( .A1(n4877), .A2(n8727), .ZN(n4875) );
  OR2_X1 U6119 ( .A1(n5032), .A2(n4607), .ZN(n4558) );
  NAND2_X1 U6120 ( .A1(n4939), .A2(n5170), .ZN(n5566) );
  OR2_X1 U6121 ( .A1(n8873), .A2(n8715), .ZN(n5815) );
  AND2_X1 U6122 ( .A1(n5078), .A2(n4502), .ZN(n4559) );
  AND3_X1 U6123 ( .A1(n6153), .A2(n6021), .A3(n6031), .ZN(n4560) );
  XNOR2_X1 U6124 ( .A(n5270), .B(n5269), .ZN(n8970) );
  AND2_X1 U6125 ( .A1(n4770), .A2(n4769), .ZN(n4561) );
  AND2_X1 U6126 ( .A1(n8020), .A2(n4516), .ZN(n4562) );
  AND2_X1 U6127 ( .A1(n4880), .A2(n4882), .ZN(n4563) );
  OR2_X1 U6128 ( .A1(n5002), .A2(n5001), .ZN(n4564) );
  NOR2_X1 U6129 ( .A1(n5072), .A2(n6732), .ZN(n5067) );
  AND2_X1 U6130 ( .A1(n5856), .A2(n4827), .ZN(n4565) );
  AND2_X1 U6131 ( .A1(n8734), .A2(n4648), .ZN(n4566) );
  AND2_X1 U6132 ( .A1(n5235), .A2(n4857), .ZN(n4567) );
  AND2_X1 U6133 ( .A1(n5017), .A2(n5950), .ZN(n4568) );
  AND2_X1 U6134 ( .A1(n5042), .A2(n5041), .ZN(n4569) );
  INV_X1 U6135 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n10403) );
  INV_X1 U6136 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U6137 ( .A1(n5516), .A2(n5515), .ZN(n9600) );
  INV_X1 U6138 ( .A(n5086), .ZN(n5085) );
  NAND2_X1 U6139 ( .A1(n5089), .A2(n5087), .ZN(n5086) );
  OR2_X1 U6140 ( .A1(n9171), .A2(n9170), .ZN(P1_U3260) );
  NAND2_X1 U6141 ( .A1(n6582), .A2(n6581), .ZN(n9236) );
  INV_X1 U6142 ( .A(n9236), .ZN(n4765) );
  NAND2_X1 U6143 ( .A1(n6617), .A2(n6616), .ZN(n9203) );
  INV_X1 U6144 ( .A(n9203), .ZN(n4761) );
  INV_X1 U6145 ( .A(n6125), .ZN(n6453) );
  AND2_X1 U6146 ( .A1(n7732), .A2(n4503), .ZN(n4571) );
  AND2_X1 U6147 ( .A1(n8775), .A2(n4790), .ZN(n4572) );
  NAND2_X1 U6148 ( .A1(n6370), .A2(n6369), .ZN(n6770) );
  NAND2_X1 U6149 ( .A1(n6247), .A2(n6246), .ZN(n9825) );
  NAND2_X1 U6150 ( .A1(n9339), .A2(n4772), .ZN(n4573) );
  AND2_X1 U6151 ( .A1(n7053), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4574) );
  INV_X1 U6152 ( .A(n8306), .ZN(n4820) );
  NAND2_X1 U6153 ( .A1(n5055), .A2(n5054), .ZN(n9358) );
  XOR2_X1 U6154 ( .A(n6360), .B(n6556), .Z(n4575) );
  NAND2_X1 U6155 ( .A1(n8998), .A2(n6364), .ZN(n9111) );
  XOR2_X1 U6156 ( .A(n6538), .B(n6556), .Z(n4576) );
  AND2_X1 U6157 ( .A1(n4904), .A2(n4907), .ZN(n4577) );
  INV_X1 U6158 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U6159 ( .A1(n7923), .A2(n4516), .ZN(n7940) );
  NAND2_X1 U6160 ( .A1(n4553), .A2(n5229), .ZN(n5529) );
  AND2_X1 U6161 ( .A1(n9443), .A2(n9302), .ZN(n4578) );
  AND2_X1 U6162 ( .A1(n4912), .A2(n4911), .ZN(n4579) );
  NAND2_X1 U6163 ( .A1(n4982), .A2(n4981), .ZN(n8997) );
  NOR2_X1 U6164 ( .A1(n9189), .A2(n9486), .ZN(n4580) );
  NAND2_X1 U6165 ( .A1(n5825), .A2(n5824), .ZN(n8852) );
  INV_X1 U6166 ( .A(n8852), .ZN(n4785) );
  OR2_X1 U6167 ( .A1(n9609), .A2(n8548), .ZN(n4581) );
  AND2_X1 U6168 ( .A1(n5647), .A2(n5646), .ZN(n8784) );
  NAND2_X1 U6169 ( .A1(n6580), .A2(n6579), .ZN(n4582) );
  INV_X1 U6170 ( .A(n9443), .ZN(n6771) );
  NAND2_X1 U6171 ( .A1(n6494), .A2(n6493), .ZN(n9443) );
  NAND2_X1 U6172 ( .A1(n6662), .A2(n9115), .ZN(n4583) );
  AND2_X1 U6173 ( .A1(n9390), .A2(n9366), .ZN(n4584) );
  NAND2_X1 U6174 ( .A1(n4876), .A2(n4874), .ZN(n4883) );
  INV_X1 U6175 ( .A(n5937), .ZN(n4844) );
  INV_X1 U6176 ( .A(n6770), .ZN(n9663) );
  AND2_X1 U6177 ( .A1(n5567), .A2(n5170), .ZN(n4585) );
  AND2_X1 U6178 ( .A1(n5013), .A2(n5012), .ZN(n4586) );
  AND2_X1 U6179 ( .A1(n7728), .A2(n7727), .ZN(n4587) );
  INV_X1 U6180 ( .A(n6693), .ZN(n4991) );
  INV_X1 U6181 ( .A(n8361), .ZN(n4803) );
  INV_X2 U6182 ( .A(n9833), .ZN(n9835) );
  NAND2_X1 U6183 ( .A1(n5496), .A2(n5495), .ZN(n7921) );
  INV_X1 U6184 ( .A(n7921), .ZN(n4786) );
  NAND2_X1 U6185 ( .A1(n6330), .A2(n6329), .ZN(n8167) );
  INV_X1 U6186 ( .A(n8167), .ZN(n4777) );
  OAI211_X1 U6187 ( .C1(n4608), .C2(n4606), .A(n4605), .B(n7478), .ZN(n7482)
         );
  NOR2_X1 U6188 ( .A1(n5529), .A2(n5234), .ZN(n5755) );
  INV_X1 U6189 ( .A(n8542), .ZN(n9611) );
  NAND2_X1 U6190 ( .A1(n7330), .A2(n5874), .ZN(n7163) );
  INV_X1 U6191 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5041) );
  NAND2_X1 U6192 ( .A1(n7421), .A2(n4870), .ZN(n7543) );
  OR2_X1 U6193 ( .A1(n9638), .A2(n7999), .ZN(n7981) );
  INV_X1 U6194 ( .A(n7981), .ZN(n4773) );
  INV_X1 U6195 ( .A(n8073), .ZN(n5023) );
  NAND2_X1 U6196 ( .A1(n5755), .A2(n5235), .ZN(n5753) );
  AND2_X1 U6197 ( .A1(n7732), .A2(n10005), .ZN(n4588) );
  AND2_X1 U6198 ( .A1(n4734), .A2(n4732), .ZN(n4589) );
  AND2_X1 U6199 ( .A1(n5821), .A2(n10390), .ZN(n4590) );
  NAND2_X1 U6200 ( .A1(n4758), .A2(n4757), .ZN(n4759) );
  NAND4_X1 U6201 ( .A1(n4592), .A2(n5052), .A3(n5053), .A4(n6029), .ZN(n4591)
         );
  AND2_X1 U6202 ( .A1(n4526), .A2(n4506), .ZN(n4592) );
  NAND2_X1 U6203 ( .A1(n7915), .A2(n9317), .ZN(n8267) );
  INV_X1 U6204 ( .A(n4781), .ZN(n7340) );
  OR2_X1 U6205 ( .A1(n7344), .A2(n7339), .ZN(n4781) );
  OR2_X1 U6206 ( .A1(n8425), .A2(n8424), .ZN(n4593) );
  INV_X1 U6207 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5497) );
  INV_X1 U6208 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6055) );
  INV_X1 U6209 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6043) );
  INV_X1 U6210 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4754) );
  INV_X1 U6211 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4620) );
  NAND2_X1 U6212 ( .A1(n5254), .A2(n5253), .ZN(n8835) );
  INV_X1 U6213 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4622) );
  MUX2_X1 U6214 ( .A(n5911), .B(n5910), .S(n5981), .Z(n5916) );
  MUX2_X1 U6215 ( .A(n5905), .B(n5904), .S(n5981), .Z(n5907) );
  INV_X1 U6216 ( .A(n4689), .ZN(n4685) );
  INV_X1 U6217 ( .A(n4956), .ZN(n4955) );
  NAND2_X1 U6218 ( .A1(n5174), .A2(n5173), .ZN(n5586) );
  NAND2_X1 U6219 ( .A1(n5528), .A2(n5527), .ZN(n4939) );
  INV_X1 U6220 ( .A(n4709), .ZN(n4708) );
  NAND2_X1 U6221 ( .A1(n4603), .A2(n5732), .ZN(n5747) );
  NAND3_X1 U6222 ( .A1(n5672), .A2(n5671), .A3(n4604), .ZN(n4694) );
  XNOR2_X2 U6223 ( .A(n5668), .B(n5669), .ZN(n8523) );
  NAND2_X1 U6224 ( .A1(n7198), .A2(n4610), .ZN(n4608) );
  NAND2_X2 U6225 ( .A1(n5028), .A2(n5027), .ZN(n8074) );
  NAND2_X2 U6226 ( .A1(n9597), .A2(n5526), .ZN(n8053) );
  NAND3_X1 U6227 ( .A1(n4853), .A2(n5229), .A3(n4507), .ZN(n4618) );
  NAND2_X1 U6228 ( .A1(n4619), .A2(n4532), .ZN(n8459) );
  AND2_X1 U6229 ( .A1(n5216), .A2(SI_0_), .ZN(n6090) );
  INV_X1 U6230 ( .A(n5122), .ZN(n4629) );
  OAI21_X1 U6231 ( .B1(n5122), .B2(n4632), .A(n4630), .ZN(n5354) );
  NAND2_X1 U6232 ( .A1(n5122), .A2(n5121), .ZN(n5345) );
  NAND3_X1 U6233 ( .A1(n4836), .A2(n4639), .A3(n4634), .ZN(n4638) );
  NAND3_X1 U6234 ( .A1(n5947), .A2(n4650), .A3(n4566), .ZN(n5949) );
  NAND2_X1 U6235 ( .A1(n4853), .A2(n4653), .ZN(n4655) );
  INV_X1 U6236 ( .A(n4655), .ZN(n8963) );
  NAND2_X1 U6237 ( .A1(n4656), .A2(n6019), .ZN(P2_U3244) );
  NAND2_X1 U6238 ( .A1(n4657), .A2(n6016), .ZN(n4656) );
  NAND3_X1 U6239 ( .A1(n4660), .A2(n4659), .A3(n4658), .ZN(n4657) );
  NAND2_X1 U6240 ( .A1(n4831), .A2(n4829), .ZN(n4658) );
  NAND2_X1 U6241 ( .A1(n4998), .A2(n5861), .ZN(n4660) );
  NAND3_X1 U6242 ( .A1(n5874), .A2(n5867), .A3(n4661), .ZN(n7330) );
  OAI21_X2 U6243 ( .B1(n4662), .B2(P2_REG3_REG_3__SCAN_IN), .A(n4499), .ZN(
        n5807) );
  INV_X2 U6244 ( .A(n5328), .ZN(n4662) );
  AND2_X1 U6245 ( .A1(n5993), .A2(n5877), .ZN(n4661) );
  NAND2_X1 U6246 ( .A1(n7872), .A2(n4668), .ZN(n4663) );
  NAND2_X1 U6247 ( .A1(n4663), .A2(n4666), .ZN(n7951) );
  OAI21_X1 U6248 ( .B1(n8696), .B2(n4676), .A(n4674), .ZN(n8627) );
  OAI21_X2 U6249 ( .B1(n5634), .B2(n4682), .A(n8464), .ZN(n8468) );
  AOI21_X1 U6250 ( .B1(n5132), .B2(n4688), .A(n4691), .ZN(n4687) );
  NAND2_X1 U6251 ( .A1(n5132), .A2(n5131), .ZN(n5406) );
  XNOR2_X2 U6252 ( .A(n4703), .B(n5688), .ZN(n8446) );
  NAND2_X1 U6253 ( .A1(n5145), .A2(n4493), .ZN(n4704) );
  NAND2_X1 U6254 ( .A1(n4704), .A2(n4705), .ZN(n5552) );
  NAND2_X1 U6255 ( .A1(n5145), .A2(n4495), .ZN(n4707) );
  NAND2_X1 U6256 ( .A1(n5145), .A2(n5144), .ZN(n5454) );
  MUX2_X1 U6257 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n6835), .Z(n5125) );
  MUX2_X1 U6258 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n6835), .Z(n5128) );
  INV_X1 U6259 ( .A(n4722), .ZN(n4972) );
  NAND2_X1 U6260 ( .A1(n4962), .A2(n4732), .ZN(n4730) );
  NAND2_X1 U6261 ( .A1(n4730), .A2(n4728), .ZN(n7890) );
  NAND2_X1 U6262 ( .A1(n9067), .A2(n9071), .ZN(n9028) );
  NAND2_X1 U6263 ( .A1(n9067), .A2(n4736), .ZN(n4735) );
  OAI21_X1 U6264 ( .B1(n4958), .B2(n4751), .A(n4749), .ZN(n7584) );
  NAND3_X1 U6265 ( .A1(n4758), .A2(n4757), .A3(n6769), .ZN(n7861) );
  NAND3_X1 U6266 ( .A1(n7622), .A2(n7501), .A3(n7682), .ZN(n7759) );
  INV_X1 U6267 ( .A(n4759), .ZN(n7758) );
  INV_X1 U6268 ( .A(n4766), .ZN(n9220) );
  INV_X2 U6269 ( .A(n5216), .ZN(n6835) );
  NAND3_X1 U6270 ( .A1(n4779), .A2(n4778), .A3(n5110), .ZN(n5284) );
  AND2_X1 U6271 ( .A1(n8661), .A2(n4782), .ZN(n8635) );
  NAND2_X1 U6272 ( .A1(n8661), .A2(n8649), .ZN(n8643) );
  NAND3_X1 U6273 ( .A1(n7732), .A2(n4503), .A3(n7942), .ZN(n7944) );
  INV_X1 U6274 ( .A(n8155), .ZN(n4793) );
  NAND2_X1 U6275 ( .A1(n8383), .A2(n8145), .ZN(n4794) );
  NAND3_X1 U6276 ( .A1(n4487), .A2(n8430), .A3(n7032), .ZN(n4800) );
  OAI21_X1 U6277 ( .B1(n6751), .B2(n4817), .A(n4815), .ZN(n6752) );
  INV_X1 U6278 ( .A(n6741), .ZN(n8345) );
  OAI21_X1 U6279 ( .B1(n6741), .B2(n7188), .A(n7187), .ZN(n7510) );
  XNOR2_X1 U6280 ( .A(n7530), .B(n6741), .ZN(n7190) );
  NAND2_X1 U6281 ( .A1(n4823), .A2(n4821), .ZN(P1_U3552) );
  NOR2_X1 U6282 ( .A1(n9840), .A2(n6779), .ZN(n4822) );
  NAND2_X1 U6283 ( .A1(n4824), .A2(n9840), .ZN(n4823) );
  XNOR2_X2 U6284 ( .A(n5267), .B(n8964), .ZN(n8085) );
  NAND2_X1 U6285 ( .A1(n4826), .A2(n4565), .ZN(n5978) );
  NAND3_X1 U6286 ( .A1(n5880), .A2(n5879), .A3(n5884), .ZN(n4836) );
  NAND2_X1 U6287 ( .A1(n4838), .A2(n4839), .ZN(n5936) );
  NAND2_X1 U6288 ( .A1(n5939), .A2(n4842), .ZN(n4838) );
  NOR2_X1 U6289 ( .A1(n5529), .A2(n4852), .ZN(n4851) );
  INV_X1 U6290 ( .A(n5014), .ZN(n4852) );
  NAND2_X1 U6291 ( .A1(n5970), .A2(n5969), .ZN(n5972) );
  AOI21_X1 U6292 ( .B1(n5906), .B2(n5988), .A(n5908), .ZN(n5911) );
  AOI21_X1 U6293 ( .B1(n5986), .B2(n5985), .A(n5984), .ZN(n5987) );
  NAND2_X1 U6294 ( .A1(n7398), .A2(n7272), .ZN(n5997) );
  NOR2_X2 U6295 ( .A1(n8064), .A2(n8030), .ZN(n8831) );
  NOR2_X2 U6296 ( .A1(n8873), .A2(n8716), .ZN(n8700) );
  AOI21_X1 U6297 ( .B1(n7923), .B2(n4562), .A(n4862), .ZN(n8022) );
  OAI21_X1 U6298 ( .B1(n7421), .B2(n4867), .A(n4865), .ZN(n7545) );
  NAND2_X1 U6299 ( .A1(n4872), .A2(n4873), .ZN(n8710) );
  NAND2_X1 U6300 ( .A1(n8758), .A2(n4563), .ZN(n4872) );
  INV_X1 U6301 ( .A(n4883), .ZN(n8888) );
  OR2_X1 U6302 ( .A1(n8695), .A2(n4513), .ZN(n4885) );
  NAND2_X1 U6303 ( .A1(n8695), .A2(n4890), .ZN(n4889) );
  NAND2_X1 U6304 ( .A1(n8827), .A2(n4489), .ZN(n4902) );
  NAND2_X1 U6305 ( .A1(n4902), .A2(n4903), .ZN(n8773) );
  NAND2_X1 U6306 ( .A1(n5178), .A2(n4924), .ZN(n4920) );
  NAND2_X1 U6307 ( .A1(n4920), .A2(n4921), .ZN(n5637) );
  NAND2_X1 U6308 ( .A1(n5354), .A2(n5353), .ZN(n4932) );
  NAND2_X1 U6309 ( .A1(n5721), .A2(n5720), .ZN(n4935) );
  NAND2_X1 U6310 ( .A1(n4939), .A2(n4585), .ZN(n5174) );
  NAND2_X1 U6311 ( .A1(n5673), .A2(n4943), .ZN(n4942) );
  NAND2_X1 U6312 ( .A1(n5673), .A2(n5200), .ZN(n5676) );
  XNOR2_X1 U6313 ( .A(n4951), .B(n5850), .ZN(n8962) );
  OAI21_X1 U6314 ( .B1(n5845), .B2(n10098), .A(n5848), .ZN(n4951) );
  NAND2_X1 U6315 ( .A1(n7319), .A2(n4959), .ZN(n4958) );
  XNOR2_X1 U6316 ( .A(n4961), .B(n7309), .ZN(n7315) );
  INV_X1 U6317 ( .A(n6226), .ZN(n4962) );
  INV_X1 U6318 ( .A(n6243), .ZN(n4966) );
  OAI21_X1 U6319 ( .B1(n6509), .B2(n4970), .A(n9081), .ZN(n4969) );
  INV_X1 U6320 ( .A(n6525), .ZN(n4970) );
  NAND2_X1 U6321 ( .A1(n4971), .A2(n6525), .ZN(n9078) );
  NAND2_X1 U6322 ( .A1(n4972), .A2(n4973), .ZN(n9067) );
  OAI211_X1 U6323 ( .C1(n9099), .C2(n6693), .A(n4988), .B(n4986), .ZN(P1_U3218) );
  NAND2_X1 U6324 ( .A1(n9099), .A2(n4989), .ZN(n4988) );
  NAND2_X1 U6325 ( .A1(n9099), .A2(n6600), .ZN(n8990) );
  NAND3_X1 U6326 ( .A1(n5053), .A2(n6029), .A3(n5052), .ZN(n6387) );
  NAND2_X1 U6327 ( .A1(n5103), .A2(n5810), .ZN(n7436) );
  INV_X1 U6328 ( .A(n5882), .ZN(n4997) );
  AND2_X1 U6329 ( .A1(n5808), .A2(n5863), .ZN(n5103) );
  XNOR2_X1 U6330 ( .A(n5860), .B(n8797), .ZN(n4998) );
  NAND2_X1 U6331 ( .A1(n4999), .A2(n4564), .ZN(n8748) );
  NAND2_X1 U6332 ( .A1(n8781), .A2(n5000), .ZN(n4999) );
  NAND2_X1 U6333 ( .A1(n7409), .A2(n7408), .ZN(n7407) );
  INV_X1 U6334 ( .A(n5013), .ZN(n8024) );
  NAND2_X1 U6335 ( .A1(n8746), .A2(n5018), .ZN(n5017) );
  NAND2_X1 U6336 ( .A1(n5017), .A2(n5016), .ZN(n8711) );
  NAND2_X1 U6337 ( .A1(n8746), .A2(n5935), .ZN(n8726) );
  INV_X1 U6338 ( .A(n5017), .ZN(n8725) );
  INV_X1 U6339 ( .A(n5935), .ZN(n5019) );
  INV_X1 U6340 ( .A(n5020), .ZN(n9947) );
  NAND2_X1 U6341 ( .A1(n5303), .A2(n5021), .ZN(n5304) );
  XNOR2_X1 U6342 ( .A(n5302), .B(n5021), .ZN(n7143) );
  OAI22_X1 U6343 ( .A1(n8505), .A2(n5804), .B1(n8542), .B2(n5021), .ZN(n7229)
         );
  XNOR2_X2 U6344 ( .A(n5744), .B(n7141), .ZN(n5021) );
  XNOR2_X1 U6345 ( .A(n5747), .B(n5746), .ZN(n5781) );
  NAND2_X1 U6346 ( .A1(n7572), .A2(n5036), .ZN(n7823) );
  NAND2_X1 U6347 ( .A1(n7906), .A2(n5039), .ZN(n5038) );
  NAND2_X1 U6348 ( .A1(n5038), .A2(n5037), .ZN(n9597) );
  NAND2_X1 U6349 ( .A1(n7906), .A2(n5492), .ZN(n6788) );
  INV_X1 U6350 ( .A(n5038), .ZN(n6787) );
  INV_X1 U6351 ( .A(n5492), .ZN(n5040) );
  NAND4_X1 U6352 ( .A1(n5229), .A2(n5356), .A3(n5228), .A4(n5042), .ZN(n5568)
         );
  NAND2_X1 U6353 ( .A1(n5045), .A2(n5043), .ZN(n6717) );
  NAND2_X1 U6354 ( .A1(n9332), .A2(n4492), .ZN(n5046) );
  NAND2_X1 U6355 ( .A1(n5046), .A2(n5047), .ZN(n9294) );
  NAND2_X1 U6356 ( .A1(n9617), .A2(n5057), .ZN(n5055) );
  NAND2_X1 U6357 ( .A1(n6054), .A2(n6055), .ZN(n6050) );
  NAND2_X1 U6358 ( .A1(n6728), .A2(n5067), .ZN(n5065) );
  NAND2_X1 U6359 ( .A1(n7851), .A2(n4559), .ZN(n5077) );
  OAI21_X1 U6360 ( .B1(n7851), .B2(n6711), .A(n5083), .ZN(n7805) );
  OAI21_X1 U6361 ( .B1(n9228), .B2(n6736), .A(n6735), .ZN(n9213) );
  NAND2_X1 U6362 ( .A1(n9228), .A2(n5091), .ZN(n5088) );
  INV_X1 U6363 ( .A(n5093), .ZN(n6740) );
  INV_X1 U6364 ( .A(n5673), .ZN(n5675) );
  INV_X1 U6365 ( .A(n9180), .ZN(n9496) );
  XNOR2_X1 U6366 ( .A(n5113), .B(n5112), .ZN(n5296) );
  NAND2_X1 U6367 ( .A1(n5305), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5306) );
  NAND2_X1 U6368 ( .A1(n5305), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5294) );
  NAND2_X1 U6369 ( .A1(n5805), .A2(n7141), .ZN(n5993) );
  OR2_X1 U6370 ( .A1(n5805), .A2(n7352), .ZN(n7157) );
  XNOR2_X1 U6371 ( .A(n8627), .B(n8624), .ZN(n8634) );
  NAND2_X1 U6372 ( .A1(n5328), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6373 ( .A1(n5352), .A2(n8509), .ZN(n7198) );
  OR2_X1 U6374 ( .A1(n6126), .A2(n6038), .ZN(n6039) );
  AND2_X1 U6375 ( .A1(n8131), .A2(n8130), .ZN(n8138) );
  XNOR2_X1 U6376 ( .A(n6117), .B(n7492), .ZN(n6120) );
  NAND2_X1 U6377 ( .A1(n7144), .A2(n7143), .ZN(n7227) );
  INV_X1 U6378 ( .A(n6036), .ZN(n8084) );
  NAND2_X1 U6379 ( .A1(n6037), .A2(n8084), .ZN(n6126) );
  NAND2_X1 U6380 ( .A1(n6037), .A2(n6036), .ZN(n6125) );
  AND2_X1 U6381 ( .A1(n7138), .A2(n5784), .ZN(n9610) );
  INV_X1 U6382 ( .A(n9610), .ZN(n5785) );
  NAND2_X2 U6383 ( .A1(n7338), .A2(n8836), .ZN(n8839) );
  INV_X1 U6384 ( .A(n8351), .ZN(n6708) );
  INV_X1 U6385 ( .A(n9915), .ZN(n5811) );
  NAND2_X2 U6386 ( .A1(n7537), .A2(n9655), .ZN(n9660) );
  INV_X1 U6387 ( .A(n6656), .ZN(n6657) );
  INV_X1 U6388 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5386) );
  OR2_X1 U6389 ( .A1(n8919), .A2(n8607), .ZN(n5095) );
  OR2_X1 U6390 ( .A1(n9189), .A2(n9532), .ZN(n5096) );
  AND2_X1 U6391 ( .A1(n5251), .A2(n5255), .ZN(n5097) );
  AND2_X1 U6392 ( .A1(n6043), .A2(n6428), .ZN(n5098) );
  AND2_X1 U6393 ( .A1(n5158), .A2(n5157), .ZN(n5099) );
  AND2_X1 U6394 ( .A1(n5144), .A2(n5143), .ZN(n5100) );
  INV_X1 U6395 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n5657) );
  INV_X1 U6396 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5423) );
  INV_X1 U6397 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5572) );
  AND2_X1 U6398 ( .A1(n5140), .A2(n5139), .ZN(n5101) );
  NAND2_X1 U6399 ( .A1(n8167), .A2(n9128), .ZN(n5102) );
  AND2_X1 U6400 ( .A1(n8688), .A2(n5815), .ZN(n5104) );
  INV_X1 U6401 ( .A(n8618), .ZN(n8619) );
  OR2_X1 U6402 ( .A1(n8654), .A2(n8526), .ZN(n5105) );
  INV_X1 U6403 ( .A(n8876), .ZN(n8617) );
  AND2_X1 U6404 ( .A1(n5109), .A2(SI_21_), .ZN(n5106) );
  INV_X1 U6405 ( .A(n8626), .ZN(n8624) );
  AND2_X1 U6406 ( .A1(n9136), .A2(n6768), .ZN(n5107) );
  NAND2_X1 U6407 ( .A1(n5865), .A2(n4635), .ZN(n5888) );
  AND2_X1 U6408 ( .A1(n7408), .A2(n5888), .ZN(n5889) );
  AND2_X1 U6409 ( .A1(n7917), .A2(n5914), .ZN(n5915) );
  INV_X1 U6410 ( .A(n5968), .ZN(n5969) );
  INV_X1 U6411 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U6412 ( .A1(n6010), .A2(n5981), .ZN(n5977) );
  OAI21_X1 U6413 ( .B1(n5976), .B2(n5857), .A(n5856), .ZN(n5858) );
  OR4_X1 U6414 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6645) );
  NOR2_X1 U6415 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n6027) );
  INV_X1 U6416 ( .A(n9415), .ZN(n6772) );
  INV_X1 U6417 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6031) );
  INV_X1 U6418 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n6021) );
  INV_X1 U6419 ( .A(SI_27_), .ZN(n10387) );
  INV_X1 U6420 ( .A(SI_13_), .ZN(n10345) );
  INV_X1 U6421 ( .A(n5660), .ZN(n5262) );
  INV_X1 U6422 ( .A(n7408), .ZN(n7403) );
  INV_X1 U6423 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6331) );
  INV_X1 U6424 ( .A(n6479), .ZN(n6478) );
  INV_X1 U6425 ( .A(n6287), .ZN(n6285) );
  INV_X1 U6426 ( .A(n9825), .ZN(n6769) );
  INV_X1 U6427 ( .A(SI_26_), .ZN(n10358) );
  INV_X1 U6428 ( .A(SI_19_), .ZN(n5179) );
  INV_X1 U6429 ( .A(SI_15_), .ZN(n10348) );
  INV_X1 U6430 ( .A(SI_10_), .ZN(n10202) );
  INV_X1 U6431 ( .A(n5622), .ZN(n5261) );
  NAND2_X1 U6432 ( .A1(n5262), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5680) );
  OR2_X1 U6433 ( .A1(n5695), .A2(n5694), .ZN(n5710) );
  OR2_X1 U6434 ( .A1(n5680), .A2(n8449), .ZN(n5682) );
  NAND2_X1 U6435 ( .A1(n5481), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5498) );
  AND2_X1 U6436 ( .A1(n7117), .A2(n7116), .ZN(n7213) );
  AND2_X1 U6437 ( .A1(n5460), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5481) );
  INV_X1 U6438 ( .A(n7941), .ZN(n8020) );
  AOI21_X1 U6439 ( .B1(n7417), .B2(n7424), .A(n5865), .ZN(n7409) );
  OR2_X1 U6440 ( .A1(n5772), .A2(n5758), .ZN(n5759) );
  INV_X1 U6441 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5388) );
  INV_X1 U6442 ( .A(n7321), .ZN(n6163) );
  INV_X1 U6443 ( .A(n9061), .ZN(n6559) );
  OR2_X1 U6444 ( .A1(n6621), .A2(n6620), .ZN(n6665) );
  OR2_X1 U6445 ( .A1(n6566), .A2(n6565), .ZN(n6585) );
  INV_X1 U6446 ( .A(n6501), .ZN(n6667) );
  OR2_X1 U6447 ( .A1(n6513), .A2(n9082), .ZN(n6529) );
  NAND2_X1 U6448 ( .A1(n6478), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6495) );
  OR2_X1 U6449 ( .A1(n6414), .A2(n6413), .ZN(n6436) );
  OR2_X1 U6450 ( .A1(n6373), .A2(n6372), .ZN(n6392) );
  NAND2_X1 U6451 ( .A1(n6285), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6309) );
  AND2_X1 U6452 ( .A1(n9374), .A2(n8302), .ZN(n9622) );
  NAND2_X1 U6453 ( .A1(n8433), .A2(n6656), .ZN(n8425) );
  INV_X1 U6454 ( .A(SI_11_), .ZN(n5146) );
  INV_X1 U6455 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10318) );
  INV_X1 U6456 ( .A(n5744), .ZN(n5724) );
  INV_X1 U6457 ( .A(n8044), .ZN(n5583) );
  INV_X1 U6458 ( .A(n6881), .ZN(n5287) );
  OR2_X1 U6459 ( .A1(n5498), .A2(n5497), .ZN(n5517) );
  OR2_X1 U6460 ( .A1(n5792), .A2(n5791), .ZN(n8481) );
  OR2_X1 U6461 ( .A1(n8646), .A2(n4662), .ZN(n5742) );
  OR2_X1 U6462 ( .A1(n5573), .A2(n5572), .ZN(n5592) );
  AND2_X1 U6463 ( .A1(n9938), .A2(n6875), .ZN(n7266) );
  NAND2_X1 U6464 ( .A1(n8632), .A2(n8631), .ZN(n8633) );
  INV_X1 U6465 ( .A(n9103), .ZN(n9118) );
  AND2_X1 U6466 ( .A1(n6622), .A2(n6665), .ZN(n9207) );
  AND2_X1 U6467 ( .A1(n6585), .A2(n6567), .ZN(n9247) );
  INV_X1 U6468 ( .A(n9126), .ZN(n9328) );
  OR2_X1 U6469 ( .A1(n6857), .A2(n6780), .ZN(n6776) );
  INV_X1 U6470 ( .A(n6774), .ZN(n9189) );
  INV_X1 U6471 ( .A(n9644), .ZN(n9382) );
  INV_X1 U6472 ( .A(n7935), .ZN(n9673) );
  INV_X1 U6473 ( .A(n7625), .ZN(n7622) );
  OR2_X1 U6474 ( .A1(n9807), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6651) );
  INV_X1 U6475 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6044) );
  AND2_X1 U6476 ( .A1(n5170), .A2(n5169), .ZN(n5527) );
  NAND2_X1 U6477 ( .A1(n5284), .A2(n5111), .ZN(n5113) );
  NOR2_X1 U6478 ( .A1(n8481), .A2(n8820), .ZN(n8516) );
  OR2_X1 U6479 ( .A1(n5783), .A2(n5777), .ZN(n5792) );
  AOI21_X1 U6480 ( .B1(n8681), .B2(n5328), .A(n5715), .ZN(n8670) );
  INV_X1 U6481 ( .A(n9842), .ZN(n9905) );
  AND2_X1 U6482 ( .A1(n6922), .A2(n6921), .ZN(n9901) );
  INV_X1 U6483 ( .A(n8623), .ZN(n8651) );
  AND2_X1 U6484 ( .A1(n5935), .A2(n5946), .ZN(n8747) );
  INV_X1 U6485 ( .A(n8612), .ZN(n8792) );
  AND2_X1 U6486 ( .A1(n8608), .A2(n8023), .ZN(n8918) );
  NAND2_X1 U6487 ( .A1(n7597), .A2(n7605), .ZN(n7648) );
  AND2_X1 U6488 ( .A1(n8839), .A2(n7464), .ZN(n9933) );
  INV_X1 U6489 ( .A(n8843), .ZN(n8736) );
  NOR2_X1 U6490 ( .A1(n9940), .A2(n5760), .ZN(n7062) );
  INV_X1 U6491 ( .A(n6882), .ZN(n10013) );
  AND3_X1 U6492 ( .A1(n5782), .A2(n8797), .A3(n7741), .ZN(n10002) );
  INV_X1 U6493 ( .A(n8934), .ZN(n10018) );
  AND2_X1 U6494 ( .A1(n6916), .A2(n9945), .ZN(n9938) );
  INV_X1 U6495 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5751) );
  INV_X1 U6496 ( .A(n8968), .ZN(n8972) );
  INV_X1 U6497 ( .A(n9117), .ZN(n9108) );
  OR2_X1 U6498 ( .A1(n9102), .A2(n6587), .ZN(n6592) );
  OR2_X1 U6499 ( .A1(n9287), .A2(n6587), .ZN(n6535) );
  INV_X1 U6500 ( .A(n9790), .ZN(n9720) );
  AND2_X1 U6501 ( .A1(n9149), .A2(n6821), .ZN(n9783) );
  AND2_X1 U6502 ( .A1(n9149), .A2(n6810), .ZN(n9796) );
  AND2_X1 U6503 ( .A1(n8208), .A2(n8272), .ZN(n9347) );
  AND2_X1 U6504 ( .A1(n7749), .A2(n7751), .ZN(n7839) );
  NOR2_X1 U6505 ( .A1(n9399), .A2(n7659), .ZN(n9641) );
  INV_X1 U6506 ( .A(n9654), .ZN(n9334) );
  INV_X1 U6507 ( .A(n9822), .ZN(n9471) );
  INV_X1 U6508 ( .A(n9826), .ZN(n9466) );
  AND2_X1 U6509 ( .A1(n6777), .A2(n7490), .ZN(n6783) );
  OR2_X1 U6510 ( .A1(n6637), .A2(n9552), .ZN(n9807) );
  INV_X1 U6511 ( .A(n9544), .ZN(n9539) );
  INV_X1 U6512 ( .A(n9945), .ZN(n6786) );
  INV_X1 U6513 ( .A(n8516), .ZN(n8527) );
  INV_X1 U6514 ( .A(n8671), .ZN(n8628) );
  INV_X1 U6515 ( .A(n8784), .ZN(n8749) );
  INV_X1 U6516 ( .A(n9901), .ZN(n9841) );
  OR2_X1 U6517 ( .A1(n7338), .A2(n7337), .ZN(n8717) );
  INV_X1 U6518 ( .A(n10036), .ZN(n10033) );
  AND2_X2 U6519 ( .A1(n7063), .A2(n7062), .ZN(n10036) );
  INV_X1 U6520 ( .A(n10021), .ZN(n10019) );
  AND2_X1 U6521 ( .A1(n7991), .A2(n8982), .ZN(n9940) );
  XNOR2_X1 U6522 ( .A(n5752), .B(n5751), .ZN(n7991) );
  INV_X1 U6523 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7358) );
  INV_X1 U6524 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6868) );
  OR2_X1 U6525 ( .A1(n6676), .A2(n9687), .ZN(n9117) );
  INV_X1 U6526 ( .A(n9115), .ZN(n9097) );
  OR3_X1 U6527 ( .A1(n6765), .A2(n6764), .A3(n6763), .ZN(n9124) );
  NAND2_X1 U6528 ( .A1(n6553), .A2(n6552), .ZN(n9280) );
  INV_X1 U6529 ( .A(n9783), .ZN(n9802) );
  OR2_X1 U6530 ( .A1(P1_U3083), .A2(n6808), .ZN(n9806) );
  NAND2_X1 U6531 ( .A1(n9660), .A2(n7493), .ZN(n9373) );
  NAND2_X1 U6532 ( .A1(n9840), .A2(n9466), .ZN(n9486) );
  INV_X1 U6533 ( .A(n9840), .ZN(n9838) );
  INV_X1 U6534 ( .A(n9007), .ZN(n9528) );
  NAND2_X1 U6535 ( .A1(n7491), .A2(n6783), .ZN(n9833) );
  INV_X1 U6536 ( .A(n9810), .ZN(n9809) );
  INV_X1 U6537 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8117) );
  INV_X1 U6538 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n10402) );
  INV_X1 U6539 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10213) );
  INV_X1 U6540 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10230) );
  NOR2_X2 U6541 ( .A1(n6916), .A2(n6786), .ZN(P2_U3966) );
  MUX2_X1 U6542 ( .A(n7781), .B(n8087), .S(n8129), .Z(n5188) );
  INV_X1 U6543 ( .A(n5188), .ZN(n5109) );
  AND2_X1 U6544 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5110) );
  NAND2_X1 U6545 ( .A1(n6090), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5111) );
  INV_X1 U6546 ( .A(SI_1_), .ZN(n5112) );
  MUX2_X1 U6547 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5216), .Z(n5295) );
  NAND2_X1 U6548 ( .A1(n5296), .A2(n5295), .ZN(n5115) );
  NAND2_X1 U6549 ( .A1(n5113), .A2(SI_1_), .ZN(n5114) );
  NAND2_X1 U6550 ( .A1(n5115), .A2(n5114), .ZN(n5311) );
  MUX2_X1 U6551 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5216), .Z(n5117) );
  INV_X1 U6552 ( .A(SI_2_), .ZN(n5116) );
  XNOR2_X1 U6553 ( .A(n5117), .B(n5116), .ZN(n5310) );
  NAND2_X1 U6554 ( .A1(n5311), .A2(n5310), .ZN(n5119) );
  NAND2_X1 U6555 ( .A1(n5117), .A2(SI_2_), .ZN(n5118) );
  NAND2_X1 U6556 ( .A1(n5119), .A2(n5118), .ZN(n5327) );
  MUX2_X1 U6557 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n5216), .Z(n5120) );
  INV_X1 U6558 ( .A(SI_3_), .ZN(n10371) );
  XNOR2_X1 U6559 ( .A(n5120), .B(n10371), .ZN(n5326) );
  NAND2_X1 U6560 ( .A1(n5327), .A2(n5326), .ZN(n5122) );
  NAND2_X1 U6561 ( .A1(n5120), .A2(SI_3_), .ZN(n5121) );
  INV_X1 U6562 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6843) );
  INV_X1 U6563 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6840) );
  MUX2_X1 U6564 ( .A(n6843), .B(n6840), .S(n5216), .Z(n5123) );
  XNOR2_X1 U6565 ( .A(n5123), .B(SI_4_), .ZN(n5344) );
  INV_X1 U6566 ( .A(n5123), .ZN(n5124) );
  INV_X1 U6567 ( .A(SI_5_), .ZN(n10413) );
  NAND2_X1 U6568 ( .A1(n5125), .A2(SI_5_), .ZN(n5126) );
  INV_X1 U6569 ( .A(SI_6_), .ZN(n5127) );
  MUX2_X1 U6570 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n8129), .Z(n5130) );
  XNOR2_X1 U6571 ( .A(n5130), .B(SI_7_), .ZN(n5380) );
  INV_X1 U6572 ( .A(n5380), .ZN(n5129) );
  NAND2_X1 U6573 ( .A1(n5381), .A2(n5129), .ZN(n5132) );
  NAND2_X1 U6574 ( .A1(n5130), .A2(SI_7_), .ZN(n5131) );
  MUX2_X1 U6575 ( .A(n6868), .B(n6866), .S(n8129), .Z(n5133) );
  INV_X1 U6576 ( .A(n5133), .ZN(n5134) );
  NAND2_X1 U6577 ( .A1(n5134), .A2(SI_8_), .ZN(n5135) );
  NAND2_X1 U6578 ( .A1(n5136), .A2(n5135), .ZN(n5405) );
  MUX2_X1 U6579 ( .A(n6870), .B(n6871), .S(n8129), .Z(n5137) );
  NAND2_X1 U6580 ( .A1(n5137), .A2(n10418), .ZN(n5140) );
  INV_X1 U6581 ( .A(n5137), .ZN(n5138) );
  NAND2_X1 U6582 ( .A1(n5138), .A2(SI_9_), .ZN(n5139) );
  MUX2_X1 U6583 ( .A(n6874), .B(n10230), .S(n8129), .Z(n5141) );
  NAND2_X1 U6584 ( .A1(n5141), .A2(n10202), .ZN(n5144) );
  INV_X1 U6585 ( .A(n5141), .ZN(n5142) );
  NAND2_X1 U6586 ( .A1(n5142), .A2(SI_10_), .ZN(n5143) );
  NAND2_X1 U6587 ( .A1(n5436), .A2(n5100), .ZN(n5145) );
  MUX2_X1 U6588 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n5216), .Z(n5147) );
  XNOR2_X1 U6589 ( .A(n5147), .B(n5146), .ZN(n5453) );
  NAND2_X1 U6590 ( .A1(n5147), .A2(SI_11_), .ZN(n5148) );
  MUX2_X1 U6591 ( .A(n7137), .B(n5149), .S(n8129), .Z(n5151) );
  INV_X1 U6592 ( .A(n5151), .ZN(n5152) );
  NAND2_X1 U6593 ( .A1(n5152), .A2(SI_12_), .ZN(n5153) );
  NAND2_X1 U6594 ( .A1(n5154), .A2(n5153), .ZN(n5471) );
  MUX2_X1 U6595 ( .A(n7175), .B(n10316), .S(n8129), .Z(n5155) );
  NAND2_X1 U6596 ( .A1(n5155), .A2(n10345), .ZN(n5158) );
  INV_X1 U6597 ( .A(n5155), .ZN(n5156) );
  NAND2_X1 U6598 ( .A1(n5156), .A2(SI_13_), .ZN(n5157) );
  MUX2_X1 U6599 ( .A(n7184), .B(n7185), .S(n8129), .Z(n5159) );
  XNOR2_X1 U6600 ( .A(n5159), .B(SI_14_), .ZN(n5510) );
  INV_X1 U6601 ( .A(n5159), .ZN(n5160) );
  MUX2_X1 U6602 ( .A(n7260), .B(n10213), .S(n5216), .Z(n5161) );
  NAND2_X1 U6603 ( .A1(n5161), .A2(n10348), .ZN(n5164) );
  INV_X1 U6604 ( .A(n5161), .ZN(n5162) );
  NAND2_X1 U6605 ( .A1(n5162), .A2(SI_15_), .ZN(n5163) );
  NAND2_X1 U6606 ( .A1(n5164), .A2(n5163), .ZN(n5551) );
  MUX2_X1 U6607 ( .A(n7358), .B(n5165), .S(n8129), .Z(n5167) );
  NAND2_X1 U6608 ( .A1(n5167), .A2(n5166), .ZN(n5170) );
  INV_X1 U6609 ( .A(n5167), .ZN(n5168) );
  NAND2_X1 U6610 ( .A1(n5168), .A2(SI_16_), .ZN(n5169) );
  MUX2_X1 U6611 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n8129), .Z(n5172) );
  XNOR2_X1 U6612 ( .A(n5172), .B(n5171), .ZN(n5567) );
  NAND2_X1 U6613 ( .A1(n5172), .A2(SI_17_), .ZN(n5173) );
  MUX2_X1 U6614 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n8129), .Z(n5176) );
  XNOR2_X1 U6615 ( .A(n5176), .B(SI_18_), .ZN(n5585) );
  INV_X1 U6616 ( .A(n5585), .ZN(n5175) );
  NAND2_X1 U6617 ( .A1(n5176), .A2(SI_18_), .ZN(n5177) );
  MUX2_X1 U6618 ( .A(n7671), .B(n10375), .S(n8129), .Z(n5180) );
  NAND2_X1 U6619 ( .A1(n5180), .A2(n5179), .ZN(n5183) );
  INV_X1 U6620 ( .A(n5180), .ZN(n5181) );
  NAND2_X1 U6621 ( .A1(n5181), .A2(SI_19_), .ZN(n5182) );
  NAND2_X1 U6622 ( .A1(n5183), .A2(n5182), .ZN(n5602) );
  MUX2_X1 U6623 ( .A(n7740), .B(n10419), .S(n8129), .Z(n5184) );
  INV_X1 U6624 ( .A(SI_20_), .ZN(n10389) );
  NAND2_X1 U6625 ( .A1(n5184), .A2(n10389), .ZN(n5187) );
  INV_X1 U6626 ( .A(n5184), .ZN(n5185) );
  NAND2_X1 U6627 ( .A1(n5185), .A2(SI_20_), .ZN(n5186) );
  XNOR2_X1 U6628 ( .A(n5188), .B(SI_21_), .ZN(n5636) );
  INV_X1 U6629 ( .A(n5636), .ZN(n5189) );
  NOR2_X1 U6630 ( .A1(n5637), .A2(n5189), .ZN(n5190) );
  MUX2_X1 U6631 ( .A(n5657), .B(n7914), .S(n8129), .Z(n5191) );
  NAND2_X1 U6632 ( .A1(n5191), .A2(n10343), .ZN(n5195) );
  INV_X1 U6633 ( .A(n5191), .ZN(n5192) );
  NAND2_X1 U6634 ( .A1(n5192), .A2(SI_22_), .ZN(n5193) );
  NAND2_X1 U6635 ( .A1(n5195), .A2(n5193), .ZN(n5653) );
  INV_X1 U6636 ( .A(n5653), .ZN(n5194) );
  NAND2_X1 U6637 ( .A1(n5652), .A2(n5194), .ZN(n5656) );
  INV_X1 U6638 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7961) );
  MUX2_X1 U6639 ( .A(n7961), .B(n10402), .S(n5216), .Z(n5197) );
  INV_X1 U6640 ( .A(SI_23_), .ZN(n5196) );
  NAND2_X1 U6641 ( .A1(n5197), .A2(n5196), .ZN(n5201) );
  INV_X1 U6642 ( .A(n5197), .ZN(n5198) );
  NAND2_X1 U6643 ( .A1(n5198), .A2(SI_23_), .ZN(n5199) );
  NAND2_X1 U6644 ( .A1(n5201), .A2(n5199), .ZN(n5674) );
  INV_X1 U6645 ( .A(n5674), .ZN(n5200) );
  MUX2_X1 U6646 ( .A(n7990), .B(n8003), .S(n8129), .Z(n5202) );
  XNOR2_X1 U6647 ( .A(n5202), .B(SI_24_), .ZN(n5242) );
  INV_X1 U6648 ( .A(n5242), .ZN(n5205) );
  INV_X1 U6649 ( .A(n5202), .ZN(n5203) );
  NAND2_X1 U6650 ( .A1(n5203), .A2(SI_24_), .ZN(n5204) );
  INV_X1 U6651 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8072) );
  INV_X1 U6652 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8068) );
  MUX2_X1 U6653 ( .A(n8072), .B(n8068), .S(n8129), .Z(n5207) );
  INV_X1 U6654 ( .A(SI_25_), .ZN(n5206) );
  NAND2_X1 U6655 ( .A1(n5207), .A2(n5206), .ZN(n5210) );
  INV_X1 U6656 ( .A(n5207), .ZN(n5208) );
  NAND2_X1 U6657 ( .A1(n5208), .A2(SI_25_), .ZN(n5209) );
  NAND2_X1 U6658 ( .A1(n5210), .A2(n5209), .ZN(n5690) );
  INV_X1 U6659 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8981) );
  INV_X1 U6660 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9550) );
  MUX2_X1 U6661 ( .A(n8981), .B(n9550), .S(n8129), .Z(n5211) );
  NAND2_X1 U6662 ( .A1(n5211), .A2(n10358), .ZN(n5214) );
  INV_X1 U6663 ( .A(n5211), .ZN(n5212) );
  NAND2_X1 U6664 ( .A1(n5212), .A2(SI_26_), .ZN(n5213) );
  NAND2_X1 U6665 ( .A1(n5707), .A2(n5706), .ZN(n5215) );
  INV_X1 U6666 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8976) );
  INV_X1 U6667 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9548) );
  MUX2_X1 U6668 ( .A(n8976), .B(n9548), .S(n5216), .Z(n5217) );
  NAND2_X1 U6669 ( .A1(n5217), .A2(n10387), .ZN(n5220) );
  INV_X1 U6670 ( .A(n5217), .ZN(n5218) );
  NAND2_X1 U6671 ( .A1(n5218), .A2(SI_27_), .ZN(n5219) );
  INV_X1 U6672 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8975) );
  MUX2_X1 U6673 ( .A(n8975), .B(n8117), .S(n8129), .Z(n5821) );
  XNOR2_X1 U6674 ( .A(n5821), .B(SI_28_), .ZN(n5819) );
  NOR2_X1 U6675 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5224) );
  AND4_X2 U6676 ( .A1(n5224), .A2(n5223), .A3(n5222), .A4(n5221), .ZN(n5229)
         );
  NOR2_X1 U6677 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5225) );
  AND2_X2 U6678 ( .A1(n5314), .A2(n5225), .ZN(n5356) );
  NOR2_X1 U6679 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5227) );
  NOR2_X1 U6680 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5226) );
  NOR2_X1 U6681 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5232) );
  NOR2_X1 U6682 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5231) );
  NOR2_X1 U6683 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5230) );
  NAND4_X1 U6684 ( .A1(n5233), .A2(n5232), .A3(n5231), .A4(n5230), .ZN(n5234)
         );
  INV_X1 U6685 ( .A(n5266), .ZN(n5238) );
  NAND2_X1 U6686 ( .A1(n6615), .A2(n4616), .ZN(n5241) );
  OR2_X1 U6687 ( .A1(n5312), .A2(n8975), .ZN(n5240) );
  NAND2_X1 U6688 ( .A1(n7989), .A2(n4616), .ZN(n5245) );
  OR2_X1 U6689 ( .A1(n5312), .A2(n7990), .ZN(n5244) );
  NAND2_X1 U6690 ( .A1(n5587), .A2(n5246), .ZN(n5250) );
  INV_X1 U6691 ( .A(n5250), .ZN(n5247) );
  NAND2_X1 U6692 ( .A1(n5247), .A2(n5097), .ZN(n5249) );
  OAI21_X2 U6693 ( .B1(n5249), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5749) );
  NAND2_X1 U6694 ( .A1(n5250), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U6695 ( .A1(n5252), .A2(n5251), .ZN(n5254) );
  NAND2_X1 U6696 ( .A1(n5778), .A2(n8797), .ZN(n6885) );
  NAND2_X1 U6697 ( .A1(n5254), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5256) );
  NAND2_X1 U6698 ( .A1(n7741), .A2(n5868), .ZN(n7270) );
  NAND2_X4 U6699 ( .A1(n5257), .A2(n7270), .ZN(n5744) );
  XNOR2_X1 U6700 ( .A(n8876), .B(n5744), .ZN(n8495) );
  NAND2_X1 U6701 ( .A1(n5359), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5393) );
  NAND2_X1 U6702 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n5258) );
  NOR2_X1 U6703 ( .A1(n5393), .A2(n5258), .ZN(n5409) );
  NAND2_X1 U6704 ( .A1(n5409), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5424) );
  NAND2_X1 U6705 ( .A1(n5539), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5543) );
  INV_X1 U6706 ( .A(n5543), .ZN(n5259) );
  INV_X1 U6707 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5607) );
  INV_X1 U6708 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8471) );
  INV_X1 U6709 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8449) );
  INV_X1 U6710 ( .A(n5682), .ZN(n5263) );
  NAND2_X1 U6711 ( .A1(n5263), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5695) );
  INV_X1 U6712 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10361) );
  NAND2_X1 U6713 ( .A1(n5682), .A2(n10361), .ZN(n5264) );
  NAND2_X1 U6714 ( .A1(n5695), .A2(n5264), .ZN(n8718) );
  OR2_X1 U6715 ( .A1(n8718), .A2(n4662), .ZN(n5277) );
  INV_X1 U6716 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n5274) );
  INV_X1 U6717 ( .A(n8970), .ZN(n5271) );
  NOR2_X2 U6718 ( .A1(n8085), .A2(n5271), .ZN(n5305) );
  NAND2_X1 U6719 ( .A1(n5305), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5273) );
  NAND2_X1 U6720 ( .A1(n4480), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5272) );
  OAI211_X1 U6721 ( .C1(n5274), .C2(n5843), .A(n5273), .B(n5272), .ZN(n5275)
         );
  INV_X1 U6722 ( .A(n5275), .ZN(n5276) );
  NAND2_X1 U6723 ( .A1(n5277), .A2(n5276), .ZN(n8618) );
  NAND2_X2 U6724 ( .A1(n4478), .A2(n8835), .ZN(n7337) );
  NAND2_X1 U6725 ( .A1(n8618), .A2(n7337), .ZN(n8498) );
  NAND2_X1 U6726 ( .A1(n5328), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5281) );
  NAND2_X1 U6727 ( .A1(n4480), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5280) );
  NAND2_X1 U6728 ( .A1(n5289), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5279) );
  NAND2_X1 U6729 ( .A1(n5305), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5278) );
  INV_X1 U6730 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U6731 ( .A1(n6835), .A2(SI_0_), .ZN(n5283) );
  INV_X1 U6732 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5282) );
  NAND2_X1 U6733 ( .A1(n5283), .A2(n5282), .ZN(n5285) );
  NAND2_X1 U6734 ( .A1(n5285), .A2(n5284), .ZN(n8984) );
  INV_X1 U6735 ( .A(n7203), .ZN(n9946) );
  NAND2_X1 U6736 ( .A1(n8561), .A2(n9946), .ZN(n6881) );
  NAND2_X1 U6737 ( .A1(n5724), .A2(n7203), .ZN(n5288) );
  AND2_X1 U6738 ( .A1(n7205), .A2(n5288), .ZN(n7144) );
  NAND2_X1 U6739 ( .A1(n5289), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5292) );
  NAND2_X1 U6740 ( .A1(n5290), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5291) );
  AND2_X1 U6741 ( .A1(n5805), .A2(n7337), .ZN(n5302) );
  XNOR2_X1 U6742 ( .A(n5296), .B(n5295), .ZN(n6837) );
  INV_X1 U6743 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6838) );
  OR2_X1 U6744 ( .A1(n5312), .A2(n6838), .ZN(n5300) );
  NAND2_X1 U6745 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5298) );
  XNOR2_X1 U6746 ( .A(n5298), .B(P2_IR_REG_1__SCAN_IN), .ZN(n9568) );
  INV_X1 U6747 ( .A(n9568), .ZN(n6836) );
  OR2_X1 U6748 ( .A1(n5313), .A2(n6836), .ZN(n5299) );
  INV_X1 U6749 ( .A(n5302), .ZN(n5303) );
  NAND2_X1 U6750 ( .A1(n7227), .A2(n5304), .ZN(n5319) );
  NAND2_X1 U6751 ( .A1(n4480), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5309) );
  NAND2_X1 U6752 ( .A1(n5289), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5307) );
  AND2_X1 U6753 ( .A1(n5806), .A2(n7337), .ZN(n5320) );
  XNOR2_X1 U6754 ( .A(n5311), .B(n5310), .ZN(n6848) );
  OR2_X1 U6755 ( .A1(n5297), .A2(n6848), .ZN(n5318) );
  INV_X1 U6756 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6849) );
  OR2_X1 U6757 ( .A1(n5312), .A2(n6849), .ZN(n5317) );
  OR2_X1 U6758 ( .A1(n5314), .A2(n5386), .ZN(n5315) );
  XNOR2_X1 U6759 ( .A(n5315), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9578) );
  INV_X1 U6760 ( .A(n9578), .ZN(n6847) );
  OR2_X1 U6761 ( .A1(n6945), .A2(n6847), .ZN(n5316) );
  XNOR2_X1 U6762 ( .A(n5744), .B(n9952), .ZN(n5322) );
  XNOR2_X1 U6763 ( .A(n5320), .B(n5322), .ZN(n7226) );
  NAND2_X1 U6764 ( .A1(n5319), .A2(n7226), .ZN(n7232) );
  INV_X1 U6765 ( .A(n5320), .ZN(n5321) );
  NAND2_X1 U6766 ( .A1(n5322), .A2(n5321), .ZN(n5323) );
  OR3_X1 U6767 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n5324) );
  NAND2_X1 U6768 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5324), .ZN(n5325) );
  XNOR2_X1 U6769 ( .A(n5325), .B(P2_IR_REG_3__SCAN_IN), .ZN(n9849) );
  INV_X1 U6770 ( .A(n9849), .ZN(n6844) );
  XNOR2_X1 U6771 ( .A(n5327), .B(n5326), .ZN(n6845) );
  INV_X1 U6772 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6846) );
  NAND2_X1 U6773 ( .A1(n4480), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5331) );
  INV_X1 U6774 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7465) );
  NAND2_X1 U6775 ( .A1(n5289), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5330) );
  NAND2_X1 U6776 ( .A1(n5834), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5329) );
  NAND2_X1 U6777 ( .A1(n5807), .A2(n7337), .ZN(n5332) );
  XNOR2_X1 U6778 ( .A(n5333), .B(n5332), .ZN(n8457) );
  INV_X1 U6779 ( .A(n5332), .ZN(n5335) );
  INV_X1 U6780 ( .A(n5333), .ZN(n5334) );
  NAND2_X1 U6781 ( .A1(n5335), .A2(n5334), .ZN(n5336) );
  NAND2_X1 U6782 ( .A1(n4480), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5343) );
  INV_X1 U6783 ( .A(n5359), .ZN(n5339) );
  INV_X1 U6784 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5337) );
  NAND2_X1 U6785 ( .A1(n7465), .A2(n5337), .ZN(n5338) );
  NAND2_X1 U6786 ( .A1(n5339), .A2(n5338), .ZN(n8513) );
  INV_X1 U6787 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6934) );
  INV_X1 U6788 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6902) );
  NOR2_X1 U6789 ( .A1(n5809), .A2(n5743), .ZN(n5349) );
  XNOR2_X1 U6790 ( .A(n5345), .B(n5344), .ZN(n6842) );
  OR2_X1 U6791 ( .A1(n6842), .A2(n5297), .ZN(n5348) );
  INV_X2 U6792 ( .A(n6945), .ZN(n5603) );
  OR2_X1 U6793 ( .A1(n5356), .A2(n5386), .ZN(n5346) );
  XNOR2_X1 U6794 ( .A(n5346), .B(P2_IR_REG_4__SCAN_IN), .ZN(n9861) );
  AOI22_X1 U6795 ( .A1(n5604), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n5603), .B2(
        n9861), .ZN(n5347) );
  NAND2_X1 U6796 ( .A1(n5348), .A2(n5347), .ZN(n8515) );
  XNOR2_X1 U6797 ( .A(n8515), .B(n5744), .ZN(n5350) );
  NAND2_X1 U6798 ( .A1(n5349), .A2(n5350), .ZN(n8508) );
  NAND2_X1 U6799 ( .A1(n8510), .A2(n8508), .ZN(n5352) );
  INV_X1 U6800 ( .A(n5349), .ZN(n5351) );
  INV_X1 U6801 ( .A(n5350), .ZN(n8504) );
  NAND2_X1 U6802 ( .A1(n5351), .A2(n8504), .ZN(n8509) );
  XNOR2_X1 U6803 ( .A(n5354), .B(n5353), .ZN(n6851) );
  OR2_X1 U6804 ( .A1(n6851), .A2(n5297), .ZN(n5358) );
  INV_X1 U6805 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5355) );
  NAND2_X1 U6806 ( .A1(n5356), .A2(n5355), .ZN(n5385) );
  NAND2_X1 U6807 ( .A1(n5385), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5366) );
  XNOR2_X1 U6808 ( .A(n5366), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9555) );
  AOI22_X1 U6809 ( .A1(n5604), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n5603), .B2(
        n9555), .ZN(n5357) );
  XNOR2_X1 U6810 ( .A(n9966), .B(n5744), .ZN(n7196) );
  OAI21_X1 U6811 ( .B1(n5359), .B2(P2_REG3_REG_5__SCAN_IN), .A(n5393), .ZN(
        n7277) );
  OR2_X1 U6812 ( .A1(n4662), .A2(n7277), .ZN(n5363) );
  NAND2_X1 U6813 ( .A1(n5834), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6814 ( .A1(n4480), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6815 ( .A1(n5289), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5360) );
  NAND2_X1 U6816 ( .A1(n8558), .A2(n7337), .ZN(n7195) );
  OR2_X1 U6817 ( .A1(n6853), .A2(n5297), .ZN(n5370) );
  INV_X1 U6818 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5383) );
  NAND2_X1 U6819 ( .A1(n5366), .A2(n5383), .ZN(n5367) );
  NAND2_X1 U6820 ( .A1(n5367), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5368) );
  XNOR2_X1 U6821 ( .A(n5368), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9874) );
  AOI22_X1 U6822 ( .A1(n5604), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n5603), .B2(
        n9874), .ZN(n5369) );
  NAND2_X1 U6823 ( .A1(n5370), .A2(n5369), .ZN(n7431) );
  XNOR2_X1 U6824 ( .A(n7431), .B(n5744), .ZN(n5376) );
  NAND2_X1 U6825 ( .A1(n4480), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5375) );
  INV_X1 U6826 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6894) );
  OR2_X1 U6827 ( .A1(n5546), .A2(n6894), .ZN(n5374) );
  INV_X1 U6828 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5371) );
  XNOR2_X1 U6829 ( .A(n5393), .B(n5371), .ZN(n7429) );
  OR2_X1 U6830 ( .A1(n4662), .A2(n7429), .ZN(n5373) );
  INV_X1 U6831 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6927) );
  OR2_X1 U6832 ( .A1(n5843), .A2(n6927), .ZN(n5372) );
  INV_X1 U6833 ( .A(n7410), .ZN(n8557) );
  NAND2_X1 U6834 ( .A1(n8557), .A2(n7337), .ZN(n5377) );
  XNOR2_X1 U6835 ( .A(n5376), .B(n5377), .ZN(n7301) );
  INV_X1 U6836 ( .A(n5376), .ZN(n5378) );
  NAND2_X1 U6837 ( .A1(n5378), .A2(n5377), .ZN(n5379) );
  XNOR2_X1 U6838 ( .A(n5381), .B(n5380), .ZN(n6861) );
  NAND2_X1 U6839 ( .A1(n6861), .A2(n4616), .ZN(n5392) );
  INV_X1 U6840 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5382) );
  NAND2_X1 U6841 ( .A1(n5383), .A2(n5382), .ZN(n5384) );
  NOR2_X1 U6842 ( .A1(n5385), .A2(n5384), .ZN(n5389) );
  OR2_X1 U6843 ( .A1(n5389), .A2(n5386), .ZN(n5387) );
  MUX2_X1 U6844 ( .A(n5387), .B(P2_IR_REG_31__SCAN_IN), .S(n5388), .Z(n5390)
         );
  NAND2_X1 U6845 ( .A1(n5389), .A2(n5388), .ZN(n5420) );
  AND2_X1 U6846 ( .A1(n5390), .A2(n5420), .ZN(n7098) );
  AOI22_X1 U6847 ( .A1(n5604), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5603), .B2(
        n7098), .ZN(n5391) );
  NAND2_X1 U6848 ( .A1(n5392), .A2(n5391), .ZN(n7541) );
  XNOR2_X1 U6849 ( .A(n7541), .B(n5744), .ZN(n5400) );
  NAND2_X1 U6850 ( .A1(n4480), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5399) );
  INV_X1 U6851 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6908) );
  OR2_X1 U6852 ( .A1(n5546), .A2(n6908), .ZN(n5398) );
  INV_X1 U6853 ( .A(n5393), .ZN(n5394) );
  AOI21_X1 U6854 ( .B1(n5394), .B2(P2_REG3_REG_6__SCAN_IN), .A(
        P2_REG3_REG_7__SCAN_IN), .ZN(n5395) );
  OR2_X1 U6855 ( .A1(n5395), .A2(n5409), .ZN(n7390) );
  OR2_X1 U6856 ( .A1(n4662), .A2(n7390), .ZN(n5397) );
  INV_X1 U6857 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6940) );
  OR2_X1 U6858 ( .A1(n5843), .A2(n6940), .ZN(n5396) );
  NOR2_X1 U6859 ( .A1(n7485), .A2(n5743), .ZN(n5401) );
  NAND2_X1 U6860 ( .A1(n5400), .A2(n5401), .ZN(n5404) );
  INV_X1 U6861 ( .A(n5400), .ZN(n7481) );
  INV_X1 U6862 ( .A(n5401), .ZN(n5402) );
  NAND2_X1 U6863 ( .A1(n7481), .A2(n5402), .ZN(n5403) );
  NAND2_X1 U6864 ( .A1(n5404), .A2(n5403), .ZN(n7388) );
  NAND2_X1 U6865 ( .A1(n5420), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5407) );
  XNOR2_X1 U6866 ( .A(n5407), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9886) );
  AOI22_X1 U6867 ( .A1(n5604), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5603), .B2(
        n9886), .ZN(n5408) );
  XNOR2_X1 U6868 ( .A(n9927), .B(n5744), .ZN(n5415) );
  NAND2_X1 U6869 ( .A1(n5834), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5414) );
  NAND2_X1 U6870 ( .A1(n4480), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5413) );
  OR2_X1 U6871 ( .A1(n5409), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5410) );
  NAND2_X1 U6872 ( .A1(n5424), .A2(n5410), .ZN(n9923) );
  OR2_X1 U6873 ( .A1(n4662), .A2(n9923), .ZN(n5412) );
  INV_X1 U6874 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6926) );
  OR2_X1 U6875 ( .A1(n5843), .A2(n6926), .ZN(n5411) );
  NOR2_X1 U6876 ( .A1(n7548), .A2(n5743), .ZN(n5416) );
  NAND2_X1 U6877 ( .A1(n5415), .A2(n5416), .ZN(n5430) );
  INV_X1 U6878 ( .A(n5415), .ZN(n7573) );
  INV_X1 U6879 ( .A(n5416), .ZN(n5417) );
  NAND2_X1 U6880 ( .A1(n7573), .A2(n5417), .ZN(n5418) );
  AND2_X1 U6881 ( .A1(n5430), .A2(n5418), .ZN(n7478) );
  XNOR2_X1 U6882 ( .A(n5419), .B(n5101), .ZN(n6869) );
  NAND2_X1 U6883 ( .A1(n6869), .A2(n4616), .ZN(n5422) );
  NAND2_X1 U6884 ( .A1(n5477), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5437) );
  XNOR2_X1 U6885 ( .A(n5437), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6985) );
  AOI22_X1 U6886 ( .A1(n5604), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5603), .B2(
        n6985), .ZN(n5421) );
  NAND2_X1 U6887 ( .A1(n5422), .A2(n5421), .ZN(n7594) );
  XNOR2_X1 U6888 ( .A(n7594), .B(n5744), .ZN(n5432) );
  NAND2_X1 U6889 ( .A1(n4480), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5429) );
  INV_X1 U6890 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7552) );
  OR2_X1 U6891 ( .A1(n5546), .A2(n7552), .ZN(n5428) );
  NAND2_X1 U6892 ( .A1(n5424), .A2(n5423), .ZN(n5425) );
  NAND2_X1 U6893 ( .A1(n5441), .A2(n5425), .ZN(n7577) );
  OR2_X1 U6894 ( .A1(n4662), .A2(n7577), .ZN(n5427) );
  INV_X1 U6895 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6925) );
  OR2_X1 U6896 ( .A1(n5843), .A2(n6925), .ZN(n5426) );
  INV_X1 U6897 ( .A(n7601), .ZN(n8554) );
  NAND2_X1 U6898 ( .A1(n8554), .A2(n7337), .ZN(n5433) );
  XNOR2_X1 U6899 ( .A(n5432), .B(n5433), .ZN(n7574) );
  AND2_X1 U6900 ( .A1(n7574), .A2(n5430), .ZN(n5431) );
  INV_X1 U6901 ( .A(n5432), .ZN(n5434) );
  NAND2_X1 U6902 ( .A1(n5434), .A2(n5433), .ZN(n5435) );
  XNOR2_X1 U6903 ( .A(n5436), .B(n5100), .ZN(n6873) );
  NAND2_X1 U6904 ( .A1(n6873), .A2(n4616), .ZN(n5440) );
  INV_X1 U6905 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U6906 ( .A1(n5437), .A2(n5474), .ZN(n5438) );
  NAND2_X1 U6907 ( .A1(n5438), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5455) );
  XNOR2_X1 U6908 ( .A(n5455), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7000) );
  AOI22_X1 U6909 ( .A1(n5604), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5603), .B2(
        n7000), .ZN(n5439) );
  NAND2_X1 U6910 ( .A1(n5440), .A2(n5439), .ZN(n7829) );
  XNOR2_X1 U6911 ( .A(n7829), .B(n5744), .ZN(n5447) );
  NAND2_X1 U6912 ( .A1(n4480), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5446) );
  INV_X1 U6913 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7611) );
  OR2_X1 U6914 ( .A1(n5546), .A2(n7611), .ZN(n5445) );
  AND2_X1 U6915 ( .A1(n5441), .A2(n10102), .ZN(n5442) );
  OR2_X1 U6916 ( .A1(n5442), .A2(n5460), .ZN(n7822) );
  OR2_X1 U6917 ( .A1(n4662), .A2(n7822), .ZN(n5444) );
  INV_X1 U6918 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6924) );
  OR2_X1 U6919 ( .A1(n5843), .A2(n6924), .ZN(n5443) );
  NOR2_X1 U6920 ( .A1(n7772), .A2(n5743), .ZN(n5448) );
  NAND2_X1 U6921 ( .A1(n5447), .A2(n5448), .ZN(n5452) );
  INV_X1 U6922 ( .A(n5447), .ZN(n7767) );
  INV_X1 U6923 ( .A(n5448), .ZN(n5449) );
  NAND2_X1 U6924 ( .A1(n7767), .A2(n5449), .ZN(n5450) );
  NAND2_X1 U6925 ( .A1(n5452), .A2(n5450), .ZN(n7826) );
  INV_X1 U6926 ( .A(n7826), .ZN(n5451) );
  NAND2_X1 U6927 ( .A1(n7823), .A2(n5452), .ZN(n5470) );
  XNOR2_X1 U6928 ( .A(n5454), .B(n5453), .ZN(n6975) );
  NAND2_X1 U6929 ( .A1(n6975), .A2(n4616), .ZN(n5459) );
  INV_X1 U6930 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U6931 ( .A1(n5455), .A2(n5475), .ZN(n5456) );
  NAND2_X1 U6932 ( .A1(n5456), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5457) );
  XNOR2_X1 U6933 ( .A(n5457), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7106) );
  AOI22_X1 U6934 ( .A1(n5604), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7106), .B2(
        n5603), .ZN(n5458) );
  NAND2_X1 U6935 ( .A1(n5459), .A2(n5458), .ZN(n7776) );
  XNOR2_X1 U6936 ( .A(n7776), .B(n5744), .ZN(n5466) );
  NAND2_X1 U6937 ( .A1(n4480), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5465) );
  INV_X1 U6938 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7654) );
  OR2_X1 U6939 ( .A1(n5546), .A2(n7654), .ZN(n5464) );
  NOR2_X1 U6940 ( .A1(n5460), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5461) );
  OR2_X1 U6941 ( .A1(n5481), .A2(n5461), .ZN(n7771) );
  OR2_X1 U6942 ( .A1(n4662), .A2(n7771), .ZN(n5463) );
  INV_X1 U6943 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6944) );
  OR2_X1 U6944 ( .A1(n5843), .A2(n6944), .ZN(n5462) );
  NOR2_X1 U6945 ( .A1(n7899), .A2(n5743), .ZN(n5467) );
  NAND2_X1 U6946 ( .A1(n5466), .A2(n5467), .ZN(n5487) );
  INV_X1 U6947 ( .A(n5466), .ZN(n7900) );
  INV_X1 U6948 ( .A(n5467), .ZN(n5468) );
  NAND2_X1 U6949 ( .A1(n7900), .A2(n5468), .ZN(n5469) );
  AND2_X1 U6950 ( .A1(n5487), .A2(n5469), .ZN(n7765) );
  NAND2_X1 U6951 ( .A1(n5470), .A2(n7765), .ZN(n7768) );
  XNOR2_X1 U6952 ( .A(n5472), .B(n5471), .ZN(n7104) );
  NAND2_X1 U6953 ( .A1(n7104), .A2(n4616), .ZN(n5480) );
  INV_X1 U6954 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5473) );
  NAND3_X1 U6955 ( .A1(n5475), .A2(n5474), .A3(n5473), .ZN(n5476) );
  OR2_X1 U6956 ( .A1(n5477), .A2(n5476), .ZN(n5494) );
  NAND2_X1 U6957 ( .A1(n5494), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5478) );
  XNOR2_X1 U6958 ( .A(n5478), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7111) );
  AOI22_X1 U6959 ( .A1(n5604), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5603), .B2(
        n7111), .ZN(n5479) );
  XNOR2_X1 U6960 ( .A(n10012), .B(n5724), .ZN(n5489) );
  OR2_X1 U6961 ( .A1(n5481), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5482) );
  NAND2_X1 U6962 ( .A1(n5498), .A2(n5482), .ZN(n7905) );
  OR2_X1 U6963 ( .A1(n4662), .A2(n7905), .ZN(n5486) );
  NAND2_X1 U6964 ( .A1(n5834), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5485) );
  NAND2_X1 U6965 ( .A1(n5290), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U6966 ( .A1(n5289), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5483) );
  NAND4_X1 U6967 ( .A1(n5486), .A2(n5485), .A3(n5484), .A4(n5483), .ZN(n8551)
         );
  NAND2_X1 U6968 ( .A1(n8551), .A2(n7337), .ZN(n5490) );
  XNOR2_X1 U6969 ( .A(n5489), .B(n5490), .ZN(n7911) );
  AND2_X1 U6970 ( .A1(n7911), .A2(n5487), .ZN(n5488) );
  NAND2_X1 U6971 ( .A1(n7768), .A2(n5488), .ZN(n7906) );
  INV_X1 U6972 ( .A(n5489), .ZN(n5491) );
  NAND2_X1 U6973 ( .A1(n5491), .A2(n5490), .ZN(n5492) );
  XNOR2_X1 U6974 ( .A(n5493), .B(n5099), .ZN(n7174) );
  NAND2_X1 U6975 ( .A1(n7174), .A2(n4616), .ZN(n5496) );
  OAI21_X1 U6976 ( .B1(n5494), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5513) );
  XNOR2_X1 U6977 ( .A(n5513), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7221) );
  AOI22_X1 U6978 ( .A1(n5604), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5603), .B2(
        n7221), .ZN(n5495) );
  XNOR2_X1 U6979 ( .A(n7921), .B(n5744), .ZN(n5504) );
  NAND2_X1 U6980 ( .A1(n5290), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5503) );
  INV_X1 U6981 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7879) );
  OR2_X1 U6982 ( .A1(n5546), .A2(n7879), .ZN(n5502) );
  NAND2_X1 U6983 ( .A1(n5498), .A2(n5497), .ZN(n5499) );
  NAND2_X1 U6984 ( .A1(n5517), .A2(n5499), .ZN(n7878) );
  OR2_X1 U6985 ( .A1(n4662), .A2(n7878), .ZN(n5501) );
  INV_X1 U6986 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7290) );
  OR2_X1 U6987 ( .A1(n5843), .A2(n7290), .ZN(n5500) );
  NOR2_X1 U6988 ( .A1(n7918), .A2(n5743), .ZN(n5505) );
  NAND2_X1 U6989 ( .A1(n5504), .A2(n5505), .ZN(n5509) );
  INV_X1 U6990 ( .A(n5504), .ZN(n5507) );
  INV_X1 U6991 ( .A(n5505), .ZN(n5506) );
  NAND2_X1 U6992 ( .A1(n5507), .A2(n5506), .ZN(n5508) );
  NAND2_X1 U6993 ( .A1(n5509), .A2(n5508), .ZN(n6789) );
  XNOR2_X1 U6994 ( .A(n5511), .B(n5510), .ZN(n7183) );
  NAND2_X1 U6995 ( .A1(n7183), .A2(n4616), .ZN(n5516) );
  INV_X1 U6996 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5512) );
  NAND2_X1 U6997 ( .A1(n5513), .A2(n5512), .ZN(n5514) );
  NAND2_X1 U6998 ( .A1(n5514), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5554) );
  XNOR2_X1 U6999 ( .A(n5554), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7448) );
  AOI22_X1 U7000 ( .A1(n7448), .A2(n5603), .B1(n5604), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5515) );
  XNOR2_X1 U7001 ( .A(n9600), .B(n5744), .ZN(n5523) );
  NAND2_X1 U7002 ( .A1(n5290), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5522) );
  AND2_X1 U7003 ( .A1(n5517), .A2(n10318), .ZN(n5518) );
  OR2_X1 U7004 ( .A1(n5539), .A2(n5518), .ZN(n9604) );
  OR2_X1 U7005 ( .A1(n4662), .A2(n9604), .ZN(n5521) );
  INV_X1 U7006 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7453) );
  OR2_X1 U7007 ( .A1(n5843), .A2(n7453), .ZN(n5520) );
  INV_X1 U7008 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7926) );
  OR2_X1 U7009 ( .A1(n5546), .A2(n7926), .ZN(n5519) );
  INV_X1 U7010 ( .A(n7950), .ZN(n8549) );
  NAND2_X1 U7011 ( .A1(n8549), .A2(n7337), .ZN(n5524) );
  XNOR2_X1 U7012 ( .A(n5523), .B(n5524), .ZN(n9598) );
  INV_X1 U7013 ( .A(n5523), .ZN(n5525) );
  NAND2_X1 U7014 ( .A1(n5525), .A2(n5524), .ZN(n5526) );
  XNOR2_X1 U7015 ( .A(n5528), .B(n5527), .ZN(n7316) );
  NAND2_X1 U7016 ( .A1(n7316), .A2(n4616), .ZN(n5533) );
  NAND2_X1 U7017 ( .A1(n5529), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5530) );
  MUX2_X1 U7018 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5530), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5531) );
  AND2_X1 U7019 ( .A1(n5531), .A2(n5568), .ZN(n7640) );
  AOI22_X1 U7020 ( .A1(n5604), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5603), .B2(
        n7640), .ZN(n5532) );
  XNOR2_X1 U7021 ( .A(n8064), .B(n5744), .ZN(n8056) );
  INV_X1 U7022 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10435) );
  NAND2_X1 U7023 ( .A1(n5543), .A2(n10435), .ZN(n5534) );
  NAND2_X1 U7024 ( .A1(n5573), .A2(n5534), .ZN(n8060) );
  OR2_X1 U7025 ( .A1(n8060), .A2(n4662), .ZN(n5538) );
  NAND2_X1 U7026 ( .A1(n5290), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5537) );
  INV_X1 U7027 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8576) );
  OR2_X1 U7028 ( .A1(n5546), .A2(n8576), .ZN(n5536) );
  INV_X1 U7029 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8564) );
  OR2_X1 U7030 ( .A1(n5843), .A2(n8564), .ZN(n5535) );
  NOR2_X1 U7031 ( .A1(n8607), .A2(n5743), .ZN(n5560) );
  NAND2_X1 U7032 ( .A1(n5290), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5550) );
  INV_X1 U7033 ( .A(n5539), .ZN(n5541) );
  INV_X1 U7034 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5540) );
  NAND2_X1 U7035 ( .A1(n5541), .A2(n5540), .ZN(n5542) );
  NAND2_X1 U7036 ( .A1(n5543), .A2(n5542), .ZN(n9615) );
  OR2_X1 U7037 ( .A1(n4662), .A2(n9615), .ZN(n5549) );
  INV_X1 U7038 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n5544) );
  OR2_X1 U7039 ( .A1(n5843), .A2(n5544), .ZN(n5548) );
  INV_X1 U7040 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n5545) );
  OR2_X1 U7041 ( .A1(n5546), .A2(n5545), .ZN(n5547) );
  NOR2_X1 U7042 ( .A1(n8061), .A2(n5743), .ZN(n5561) );
  XNOR2_X1 U7043 ( .A(n5552), .B(n5551), .ZN(n7259) );
  NAND2_X1 U7044 ( .A1(n7259), .A2(n4616), .ZN(n5558) );
  INV_X1 U7045 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5553) );
  NAND2_X1 U7046 ( .A1(n5554), .A2(n5553), .ZN(n5555) );
  NAND2_X1 U7047 ( .A1(n5555), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5556) );
  XNOR2_X1 U7048 ( .A(n5556), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7636) );
  AOI22_X1 U7049 ( .A1(n7636), .A2(n5603), .B1(n5604), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5557) );
  XNOR2_X1 U7050 ( .A(n9609), .B(n5744), .ZN(n8052) );
  AOI22_X1 U7051 ( .A1(n8056), .A2(n5560), .B1(n5561), .B2(n8052), .ZN(n5559)
         );
  INV_X1 U7052 ( .A(n8056), .ZN(n5564) );
  OAI21_X1 U7053 ( .B1(n8052), .B2(n5561), .A(n5560), .ZN(n5563) );
  INV_X1 U7054 ( .A(n8052), .ZN(n8054) );
  INV_X1 U7055 ( .A(n5560), .ZN(n8055) );
  INV_X1 U7056 ( .A(n5561), .ZN(n9607) );
  AND2_X1 U7057 ( .A1(n8055), .A2(n9607), .ZN(n5562) );
  AOI22_X1 U7058 ( .A1(n5564), .A2(n5563), .B1(n8054), .B2(n5562), .ZN(n5565)
         );
  XNOR2_X1 U7059 ( .A(n5566), .B(n5567), .ZN(n7386) );
  NAND2_X1 U7060 ( .A1(n7386), .A2(n4616), .ZN(n5571) );
  NAND2_X1 U7061 ( .A1(n5568), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5569) );
  XNOR2_X1 U7062 ( .A(n5569), .B(n5041), .ZN(n8573) );
  INV_X1 U7063 ( .A(n8573), .ZN(n9904) );
  AOI22_X1 U7064 ( .A1(n5604), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5603), .B2(
        n9904), .ZN(n5570) );
  XNOR2_X1 U7065 ( .A(n8914), .B(n5744), .ZN(n5579) );
  NAND2_X1 U7066 ( .A1(n5573), .A2(n5572), .ZN(n5574) );
  NAND2_X1 U7067 ( .A1(n5592), .A2(n5574), .ZN(n8837) );
  NAND2_X1 U7068 ( .A1(n5834), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U7069 ( .A1(n5290), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5575) );
  AND2_X1 U7070 ( .A1(n5576), .A2(n5575), .ZN(n5578) );
  NAND2_X1 U7071 ( .A1(n5289), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5577) );
  OAI211_X1 U7072 ( .C1(n8837), .C2(n4662), .A(n5578), .B(n5577), .ZN(n8546)
         );
  AND2_X1 U7073 ( .A1(n8546), .A2(n7337), .ZN(n5580) );
  NAND2_X1 U7074 ( .A1(n5579), .A2(n5580), .ZN(n5584) );
  INV_X1 U7075 ( .A(n5579), .ZN(n8075) );
  INV_X1 U7076 ( .A(n5580), .ZN(n5581) );
  NAND2_X1 U7077 ( .A1(n8075), .A2(n5581), .ZN(n5582) );
  NAND2_X1 U7078 ( .A1(n5584), .A2(n5582), .ZN(n8044) );
  XNOR2_X1 U7079 ( .A(n5586), .B(n5585), .ZN(n7519) );
  NAND2_X1 U7080 ( .A1(n7519), .A2(n4616), .ZN(n5591) );
  INV_X1 U7081 ( .A(n5587), .ZN(n5588) );
  NAND2_X1 U7082 ( .A1(n5588), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5589) );
  XNOR2_X1 U7083 ( .A(n5589), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8578) );
  AOI22_X1 U7084 ( .A1(n5604), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5603), .B2(
        n8578), .ZN(n5590) );
  XNOR2_X1 U7085 ( .A(n8909), .B(n5744), .ZN(n8118) );
  INV_X1 U7086 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10427) );
  NAND2_X1 U7087 ( .A1(n5592), .A2(n10427), .ZN(n5593) );
  NAND2_X1 U7088 ( .A1(n5608), .A2(n5593), .ZN(n8810) );
  OR2_X1 U7089 ( .A1(n8810), .A2(n4662), .ZN(n5596) );
  AOI22_X1 U7090 ( .A1(n5834), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n5290), .B2(
        P2_REG0_REG_18__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U7091 ( .A1(n5289), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5594) );
  NOR2_X1 U7092 ( .A1(n8610), .A2(n5743), .ZN(n5597) );
  NAND2_X1 U7093 ( .A1(n8118), .A2(n5597), .ZN(n5613) );
  INV_X1 U7094 ( .A(n8118), .ZN(n5599) );
  INV_X1 U7095 ( .A(n5597), .ZN(n5598) );
  NAND2_X1 U7096 ( .A1(n5599), .A2(n5598), .ZN(n5600) );
  AND2_X1 U7097 ( .A1(n5613), .A2(n5600), .ZN(n8073) );
  AOI22_X1 U7098 ( .A1(n5604), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8797), .B2(
        n5603), .ZN(n5605) );
  NAND2_X1 U7099 ( .A1(n5608), .A2(n5607), .ZN(n5609) );
  AND2_X1 U7100 ( .A1(n5622), .A2(n5609), .ZN(n8800) );
  NAND2_X1 U7101 ( .A1(n8800), .A2(n5328), .ZN(n5612) );
  AOI22_X1 U7102 ( .A1(n5305), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n5290), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U7103 ( .A1(n5289), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5610) );
  NOR2_X1 U7104 ( .A1(n8821), .A2(n5743), .ZN(n5615) );
  INV_X1 U7105 ( .A(n5615), .ZN(n5616) );
  XNOR2_X1 U7106 ( .A(n5619), .B(n5618), .ZN(n7739) );
  NAND2_X1 U7107 ( .A1(n7739), .A2(n4616), .ZN(n5621) );
  OR2_X1 U7108 ( .A1(n5312), .A2(n7740), .ZN(n5620) );
  XNOR2_X1 U7109 ( .A(n8900), .B(n5744), .ZN(n5630) );
  INV_X1 U7110 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10347) );
  NAND2_X1 U7111 ( .A1(n5622), .A2(n10347), .ZN(n5623) );
  NAND2_X1 U7112 ( .A1(n5640), .A2(n5623), .ZN(n8777) );
  OR2_X1 U7113 ( .A1(n8777), .A2(n4662), .ZN(n5629) );
  INV_X1 U7114 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U7115 ( .A1(n5834), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U7116 ( .A1(n4480), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5624) );
  OAI211_X1 U7117 ( .C1(n5626), .C2(n5843), .A(n5625), .B(n5624), .ZN(n5627)
         );
  INV_X1 U7118 ( .A(n5627), .ZN(n5628) );
  NOR2_X1 U7119 ( .A1(n8762), .A2(n5743), .ZN(n5631) );
  NAND2_X1 U7120 ( .A1(n5630), .A2(n5631), .ZN(n5635) );
  INV_X1 U7121 ( .A(n5630), .ZN(n8467) );
  INV_X1 U7122 ( .A(n5631), .ZN(n5632) );
  NAND2_X1 U7123 ( .A1(n8467), .A2(n5632), .ZN(n5633) );
  NAND2_X1 U7124 ( .A1(n5635), .A2(n5633), .ZN(n6795) );
  XNOR2_X1 U7125 ( .A(n5637), .B(n5636), .ZN(n7780) );
  NAND2_X1 U7126 ( .A1(n7780), .A2(n4616), .ZN(n5639) );
  OR2_X1 U7127 ( .A1(n5312), .A2(n7781), .ZN(n5638) );
  XNOR2_X1 U7128 ( .A(n8895), .B(n5724), .ZN(n5648) );
  NAND2_X1 U7129 ( .A1(n5640), .A2(n8471), .ZN(n5641) );
  AND2_X1 U7130 ( .A1(n5660), .A2(n5641), .ZN(n8767) );
  NAND2_X1 U7131 ( .A1(n8767), .A2(n5328), .ZN(n5647) );
  INV_X1 U7132 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U7133 ( .A1(n5305), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5643) );
  NAND2_X1 U7134 ( .A1(n5290), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5642) );
  OAI211_X1 U7135 ( .C1(n5644), .C2(n5843), .A(n5643), .B(n5642), .ZN(n5645)
         );
  INV_X1 U7136 ( .A(n5645), .ZN(n5646) );
  NOR2_X1 U7137 ( .A1(n8784), .A2(n5743), .ZN(n5649) );
  XNOR2_X1 U7138 ( .A(n5648), .B(n5649), .ZN(n8464) );
  INV_X1 U7139 ( .A(n5648), .ZN(n5650) );
  NAND2_X1 U7140 ( .A1(n5650), .A2(n5649), .ZN(n5651) );
  INV_X1 U7141 ( .A(n5652), .ZN(n5654) );
  NAND2_X1 U7142 ( .A1(n5654), .A2(n5653), .ZN(n5655) );
  NAND2_X1 U7143 ( .A1(n5656), .A2(n5655), .ZN(n7913) );
  NAND2_X1 U7144 ( .A1(n7913), .A2(n4616), .ZN(n5659) );
  OR2_X1 U7145 ( .A1(n5312), .A2(n5657), .ZN(n5658) );
  XNOR2_X1 U7146 ( .A(n8889), .B(n5724), .ZN(n5669) );
  INV_X1 U7147 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10085) );
  NAND2_X1 U7148 ( .A1(n5660), .A2(n10085), .ZN(n5661) );
  NAND2_X1 U7149 ( .A1(n5680), .A2(n5661), .ZN(n8742) );
  OR2_X1 U7150 ( .A1(n8742), .A2(n4662), .ZN(n5667) );
  INV_X1 U7151 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n5664) );
  NAND2_X1 U7152 ( .A1(n5834), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U7153 ( .A1(n5290), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5662) );
  OAI211_X1 U7154 ( .C1(n5664), .C2(n5843), .A(n5663), .B(n5662), .ZN(n5665)
         );
  INV_X1 U7155 ( .A(n5665), .ZN(n5666) );
  NAND2_X1 U7156 ( .A1(n8616), .A2(n7337), .ZN(n8522) );
  INV_X1 U7157 ( .A(n5668), .ZN(n5670) );
  NAND2_X1 U7158 ( .A1(n5675), .A2(n5674), .ZN(n5677) );
  NAND2_X1 U7159 ( .A1(n5677), .A2(n5676), .ZN(n7958) );
  NAND2_X1 U7160 ( .A1(n7958), .A2(n4616), .ZN(n5679) );
  OR2_X1 U7161 ( .A1(n5312), .A2(n7961), .ZN(n5678) );
  XNOR2_X1 U7162 ( .A(n8883), .B(n5744), .ZN(n5688) );
  NAND2_X1 U7163 ( .A1(n5680), .A2(n8449), .ZN(n5681) );
  AND2_X1 U7164 ( .A1(n5682), .A2(n5681), .ZN(n8730) );
  INV_X1 U7165 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U7166 ( .A1(n5834), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U7167 ( .A1(n4480), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5683) );
  OAI211_X1 U7168 ( .C1(n5685), .C2(n5843), .A(n5684), .B(n5683), .ZN(n5686)
         );
  AOI21_X1 U7169 ( .B1(n8730), .B2(n5328), .A(n5686), .ZN(n8528) );
  OR2_X1 U7170 ( .A1(n8528), .A2(n5743), .ZN(n8447) );
  AOI21_X1 U7171 ( .B1(n8495), .B2(n8619), .A(n8447), .ZN(n5687) );
  NAND2_X1 U7172 ( .A1(n8495), .A2(n8498), .ZN(n5689) );
  NAND2_X1 U7173 ( .A1(n8067), .A2(n4616), .ZN(n5693) );
  OR2_X1 U7174 ( .A1(n5312), .A2(n8072), .ZN(n5692) );
  XNOR2_X1 U7175 ( .A(n8873), .B(n5744), .ZN(n8484) );
  INV_X1 U7176 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5694) );
  NAND2_X1 U7177 ( .A1(n5695), .A2(n5694), .ZN(n5696) );
  NAND2_X1 U7178 ( .A1(n5710), .A2(n5696), .ZN(n8478) );
  OR2_X1 U7179 ( .A1(n8478), .A2(n4662), .ZN(n5702) );
  INV_X1 U7180 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n5699) );
  NAND2_X1 U7181 ( .A1(n5305), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5698) );
  NAND2_X1 U7182 ( .A1(n5290), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5697) );
  OAI211_X1 U7183 ( .C1(n5699), .C2(n5843), .A(n5698), .B(n5697), .ZN(n5700)
         );
  INV_X1 U7184 ( .A(n5700), .ZN(n5701) );
  NOR2_X1 U7185 ( .A1(n8715), .A2(n5743), .ZN(n5703) );
  AND2_X1 U7186 ( .A1(n8484), .A2(n5703), .ZN(n8482) );
  INV_X1 U7187 ( .A(n8484), .ZN(n5705) );
  INV_X1 U7188 ( .A(n5703), .ZN(n5704) );
  NAND2_X1 U7189 ( .A1(n5705), .A2(n5704), .ZN(n8486) );
  XNOR2_X1 U7190 ( .A(n5707), .B(n5706), .ZN(n8979) );
  NAND2_X1 U7191 ( .A1(n8979), .A2(n4616), .ZN(n5709) );
  OR2_X1 U7192 ( .A1(n5312), .A2(n8981), .ZN(n5708) );
  XNOR2_X1 U7193 ( .A(n8867), .B(n5744), .ZN(n5716) );
  INV_X1 U7194 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8537) );
  NAND2_X1 U7195 ( .A1(n5710), .A2(n8537), .ZN(n5711) );
  INV_X1 U7196 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n5714) );
  NAND2_X1 U7197 ( .A1(n5834), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5713) );
  NAND2_X1 U7198 ( .A1(n4480), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5712) );
  OAI211_X1 U7199 ( .C1(n5714), .C2(n5843), .A(n5713), .B(n5712), .ZN(n5715)
         );
  NOR2_X1 U7200 ( .A1(n8670), .A2(n5743), .ZN(n5717) );
  XNOR2_X1 U7201 ( .A(n5716), .B(n5717), .ZN(n8533) );
  INV_X1 U7202 ( .A(n5716), .ZN(n5719) );
  INV_X1 U7203 ( .A(n5717), .ZN(n5718) );
  NAND2_X1 U7204 ( .A1(n6601), .A2(n4616), .ZN(n5723) );
  OR2_X1 U7205 ( .A1(n5312), .A2(n8976), .ZN(n5722) );
  XNOR2_X1 U7206 ( .A(n8861), .B(n5724), .ZN(n5729) );
  XNOR2_X1 U7207 ( .A(n5735), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8662) );
  INV_X1 U7208 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n5727) );
  NAND2_X1 U7209 ( .A1(n5305), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5726) );
  NAND2_X1 U7210 ( .A1(n5290), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5725) );
  OAI211_X1 U7211 ( .C1(n5727), .C2(n5843), .A(n5726), .B(n5725), .ZN(n5728)
         );
  AOI21_X1 U7212 ( .B1(n8662), .B2(n5328), .A(n5728), .ZN(n8654) );
  NOR2_X1 U7213 ( .A1(n8654), .A2(n5743), .ZN(n5730) );
  XNOR2_X1 U7214 ( .A(n5729), .B(n5730), .ZN(n8439) );
  INV_X1 U7215 ( .A(n5729), .ZN(n5731) );
  NAND2_X1 U7216 ( .A1(n5731), .A2(n5730), .ZN(n5732) );
  INV_X1 U7217 ( .A(n5735), .ZN(n5734) );
  AND2_X1 U7218 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n5733) );
  NAND2_X1 U7219 ( .A1(n5734), .A2(n5733), .ZN(n5786) );
  INV_X1 U7220 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8440) );
  INV_X1 U7221 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5796) );
  OAI21_X1 U7222 ( .B1(n5735), .B2(n8440), .A(n5796), .ZN(n5736) );
  NAND2_X1 U7223 ( .A1(n5786), .A2(n5736), .ZN(n8646) );
  INV_X1 U7224 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n5739) );
  NAND2_X1 U7225 ( .A1(n5305), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5738) );
  NAND2_X1 U7226 ( .A1(n5290), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5737) );
  OAI211_X1 U7227 ( .C1(n5739), .C2(n5843), .A(n5738), .B(n5737), .ZN(n5740)
         );
  INV_X1 U7228 ( .A(n5740), .ZN(n5741) );
  NOR2_X1 U7229 ( .A1(n8671), .A2(n5743), .ZN(n5745) );
  XNOR2_X1 U7230 ( .A(n5745), .B(n5744), .ZN(n5746) );
  INV_X1 U7231 ( .A(n5781), .ZN(n5780) );
  NAND2_X1 U7232 ( .A1(n5749), .A2(n5748), .ZN(n5750) );
  NAND2_X1 U7233 ( .A1(n5753), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5754) );
  NAND2_X1 U7234 ( .A1(n5756), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5757) );
  XNOR2_X1 U7235 ( .A(n5757), .B(P2_IR_REG_25__SCAN_IN), .ZN(n5772) );
  XOR2_X1 U7236 ( .A(n7991), .B(P2_B_REG_SCAN_IN), .Z(n5758) );
  INV_X1 U7237 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9941) );
  INV_X1 U7238 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9943) );
  NOR2_X1 U7239 ( .A1(n5772), .A2(n5761), .ZN(n9944) );
  AOI21_X1 U7240 ( .B1(n9937), .B2(n9943), .A(n9944), .ZN(n6877) );
  NOR4_X1 U7241 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5765) );
  NOR4_X1 U7242 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5764) );
  NOR4_X1 U7243 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5763) );
  NOR4_X1 U7244 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5762) );
  NAND4_X1 U7245 ( .A1(n5765), .A2(n5764), .A3(n5763), .A4(n5762), .ZN(n5771)
         );
  NOR2_X1 U7246 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n5769) );
  NOR4_X1 U7247 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n5768) );
  NOR4_X1 U7248 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5767) );
  NOR4_X1 U7249 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5766) );
  NAND4_X1 U7250 ( .A1(n5769), .A2(n5768), .A3(n5767), .A4(n5766), .ZN(n5770)
         );
  OAI21_X1 U7251 ( .B1(n5771), .B2(n5770), .A(n9937), .ZN(n6876) );
  AND2_X1 U7252 ( .A1(n6877), .A2(n6876), .ZN(n7265) );
  NAND2_X1 U7253 ( .A1(n7062), .A2(n7265), .ZN(n5783) );
  INV_X1 U7254 ( .A(n5772), .ZN(n8070) );
  OR2_X1 U7255 ( .A1(n5774), .A2(n5773), .ZN(n5775) );
  NAND2_X1 U7256 ( .A1(n5776), .A2(n5775), .ZN(n6015) );
  INV_X1 U7257 ( .A(n9938), .ZN(n5777) );
  INV_X1 U7258 ( .A(n6017), .ZN(n5791) );
  NAND2_X1 U7259 ( .A1(n5778), .A2(n5868), .ZN(n6915) );
  INV_X1 U7260 ( .A(n6915), .ZN(n5799) );
  OR2_X1 U7261 ( .A1(n8930), .A2(n5799), .ZN(n5779) );
  OR2_X2 U7262 ( .A1(n5792), .A2(n5779), .ZN(n8542) );
  NAND2_X1 U7263 ( .A1(n5780), .A2(n9611), .ZN(n5803) );
  NAND2_X1 U7264 ( .A1(n10002), .A2(n7782), .ZN(n7268) );
  NAND2_X1 U7265 ( .A1(n5783), .A2(n7268), .ZN(n7138) );
  AND2_X1 U7266 ( .A1(n9938), .A2(n8930), .ZN(n5784) );
  INV_X1 U7267 ( .A(n5786), .ZN(n8636) );
  INV_X1 U7268 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U7269 ( .A1(n5834), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5788) );
  NAND2_X1 U7270 ( .A1(n4480), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5787) );
  OAI211_X1 U7271 ( .C1(n5789), .C2(n5843), .A(n5788), .B(n5787), .ZN(n5790)
         );
  AOI21_X1 U7272 ( .B1(n8636), .B2(n5328), .A(n5790), .ZN(n8653) );
  INV_X1 U7273 ( .A(n8653), .ZN(n8544) );
  INV_X1 U7274 ( .A(n5793), .ZN(n5798) );
  OR2_X1 U7275 ( .A1(n6915), .A2(n6017), .ZN(n6875) );
  AND3_X1 U7276 ( .A1(n6916), .A2(n6015), .A3(n6875), .ZN(n5794) );
  NAND2_X1 U7277 ( .A1(n7138), .A2(n5794), .ZN(n5795) );
  OAI22_X1 U7278 ( .A1(n8646), .A2(n9616), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5796), .ZN(n5797) );
  AOI21_X1 U7279 ( .B1(n8544), .B2(n8516), .A(n5797), .ZN(n5800) );
  AND2_X1 U7280 ( .A1(n5800), .A2(n5105), .ZN(n5801) );
  OAI211_X1 U7281 ( .C1(n5817), .C2(n5803), .A(n5802), .B(n5801), .ZN(P2_U3222) );
  INV_X1 U7282 ( .A(n5805), .ZN(n5804) );
  NAND2_X1 U7283 ( .A1(n5804), .A2(n7352), .ZN(n5994) );
  NAND2_X1 U7284 ( .A1(n5806), .A2(n9952), .ZN(n5877) );
  OR2_X1 U7285 ( .A1(n5807), .A2(n8455), .ZN(n5863) );
  INV_X1 U7286 ( .A(n8515), .ZN(n9958) );
  NAND2_X1 U7287 ( .A1(n5809), .A2(n8515), .ZN(n5864) );
  NAND2_X1 U7288 ( .A1(n9966), .A2(n8558), .ZN(n5998) );
  INV_X1 U7289 ( .A(n8558), .ZN(n7398) );
  INV_X1 U7290 ( .A(n9966), .ZN(n7272) );
  OR2_X1 U7291 ( .A1(n7431), .A2(n7410), .ZN(n5884) );
  NAND2_X1 U7292 ( .A1(n7431), .A2(n7410), .ZN(n5887) );
  INV_X1 U7293 ( .A(n5887), .ZN(n5865) );
  OR2_X1 U7294 ( .A1(n7541), .A2(n7485), .ZN(n5891) );
  NAND2_X1 U7295 ( .A1(n7541), .A2(n7485), .ZN(n5890) );
  NAND2_X1 U7296 ( .A1(n9927), .A2(n7548), .ZN(n5895) );
  NAND2_X1 U7297 ( .A1(n5894), .A2(n5895), .ZN(n9915) );
  NAND2_X1 U7298 ( .A1(n9919), .A2(n5895), .ZN(n7547) );
  OR2_X1 U7299 ( .A1(n7594), .A2(n7601), .ZN(n5992) );
  NAND2_X1 U7300 ( .A1(n7547), .A2(n5992), .ZN(n7604) );
  OR2_X1 U7301 ( .A1(n7829), .A2(n7772), .ZN(n7650) );
  NAND2_X1 U7302 ( .A1(n7829), .A2(n7772), .ZN(n5899) );
  NAND2_X1 U7303 ( .A1(n7650), .A2(n5899), .ZN(n7605) );
  AND2_X1 U7304 ( .A1(n7594), .A2(n7601), .ZN(n5893) );
  NOR2_X1 U7305 ( .A1(n7605), .A2(n5893), .ZN(n5812) );
  NAND2_X1 U7306 ( .A1(n7604), .A2(n5812), .ZN(n7607) );
  OR2_X1 U7307 ( .A1(n7776), .A2(n7899), .ZN(n5991) );
  AND2_X1 U7308 ( .A1(n5991), .A2(n7650), .ZN(n5902) );
  AND2_X1 U7309 ( .A1(n7776), .A2(n7899), .ZN(n5897) );
  AOI21_X2 U7310 ( .B1(n7607), .B2(n5902), .A(n5897), .ZN(n7729) );
  INV_X1 U7311 ( .A(n8551), .ZN(n7773) );
  NAND2_X1 U7312 ( .A1(n7909), .A2(n7773), .ZN(n5988) );
  AND2_X1 U7313 ( .A1(n10012), .A2(n8551), .ZN(n5908) );
  AOI21_X2 U7314 ( .B1(n7729), .B2(n5988), .A(n5908), .ZN(n7872) );
  OR2_X1 U7315 ( .A1(n7921), .A2(n7918), .ZN(n5913) );
  NAND2_X1 U7316 ( .A1(n7921), .A2(n7918), .ZN(n5912) );
  NAND2_X1 U7317 ( .A1(n9600), .A2(n7950), .ZN(n5918) );
  NAND2_X1 U7318 ( .A1(n9609), .A2(n8061), .ZN(n5921) );
  NAND2_X1 U7319 ( .A1(n7951), .A2(n5922), .ZN(n8025) );
  XNOR2_X1 U7320 ( .A(n8064), .B(n8607), .ZN(n8026) );
  INV_X1 U7321 ( .A(n8546), .ZN(n8819) );
  OR2_X1 U7322 ( .A1(n8909), .A2(n8610), .ZN(n5929) );
  NAND2_X1 U7323 ( .A1(n8909), .A2(n8610), .ZN(n5937) );
  NAND2_X1 U7324 ( .A1(n5929), .A2(n5937), .ZN(n8816) );
  INV_X1 U7325 ( .A(n5929), .ZN(n8791) );
  OR2_X1 U7326 ( .A1(n8906), .A2(n8821), .ZN(n5938) );
  NAND2_X1 U7327 ( .A1(n8906), .A2(n8821), .ZN(n5941) );
  NAND2_X1 U7328 ( .A1(n5938), .A2(n5941), .ZN(n8612) );
  NOR3_X1 U7329 ( .A1(n8815), .A2(n8791), .A3(n8612), .ZN(n5813) );
  INV_X1 U7330 ( .A(n5941), .ZN(n5934) );
  NOR2_X1 U7331 ( .A1(n5813), .A2(n5934), .ZN(n8781) );
  NAND2_X1 U7332 ( .A1(n8900), .A2(n8762), .ZN(n5940) );
  XNOR2_X1 U7333 ( .A(n8895), .B(n8784), .ZN(n8760) );
  NAND2_X1 U7334 ( .A1(n8889), .A2(n8763), .ZN(n5946) );
  NAND2_X1 U7335 ( .A1(n8748), .A2(n8747), .ZN(n8746) );
  OR2_X1 U7336 ( .A1(n8883), .A2(n8528), .ZN(n5951) );
  NAND2_X1 U7337 ( .A1(n8883), .A2(n8528), .ZN(n5950) );
  NAND2_X1 U7338 ( .A1(n5951), .A2(n5950), .ZN(n8727) );
  NOR2_X1 U7339 ( .A1(n8876), .A2(n8618), .ZN(n5956) );
  NOR2_X1 U7340 ( .A1(n8617), .A2(n8619), .ZN(n5814) );
  NOR2_X1 U7341 ( .A1(n5956), .A2(n5814), .ZN(n8712) );
  INV_X1 U7342 ( .A(n5814), .ZN(n5953) );
  NAND2_X1 U7343 ( .A1(n8711), .A2(n5953), .ZN(n8696) );
  NAND2_X1 U7344 ( .A1(n8873), .A2(n8715), .ZN(n5957) );
  NOR2_X1 U7345 ( .A1(n8867), .A2(n8670), .ZN(n5960) );
  NAND2_X1 U7346 ( .A1(n8861), .A2(n8654), .ZN(n5965) );
  AND2_X2 U7347 ( .A1(n5964), .A2(n5965), .ZN(n8666) );
  NAND2_X1 U7348 ( .A1(n5817), .A2(n8671), .ZN(n5971) );
  INV_X1 U7349 ( .A(n8627), .ZN(n5827) );
  INV_X1 U7350 ( .A(SI_28_), .ZN(n10390) );
  MUX2_X1 U7351 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n6835), .Z(n5828) );
  INV_X1 U7352 ( .A(SI_29_), .ZN(n5822) );
  XNOR2_X1 U7353 ( .A(n5828), .B(n5822), .ZN(n5823) );
  NAND2_X1 U7354 ( .A1(n8082), .A2(n4616), .ZN(n5825) );
  INV_X1 U7355 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8969) );
  OR2_X1 U7356 ( .A1(n5312), .A2(n8969), .ZN(n5824) );
  INV_X1 U7357 ( .A(n5973), .ZN(n5826) );
  NAND2_X1 U7358 ( .A1(n8852), .A2(n8653), .ZN(n5974) );
  NOR2_X1 U7359 ( .A1(n5828), .A2(SI_29_), .ZN(n5830) );
  NAND2_X1 U7360 ( .A1(n5828), .A2(SI_29_), .ZN(n5829) );
  MUX2_X1 U7361 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6835), .Z(n5846) );
  XNOR2_X1 U7362 ( .A(n5847), .B(n5846), .ZN(n5845) );
  NAND2_X1 U7363 ( .A1(n8133), .A2(n4616), .ZN(n5833) );
  INV_X1 U7364 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8086) );
  OR2_X1 U7365 ( .A1(n5312), .A2(n8086), .ZN(n5832) );
  NAND2_X1 U7366 ( .A1(n5289), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5837) );
  NAND2_X1 U7367 ( .A1(n5834), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n5836) );
  NAND2_X1 U7368 ( .A1(n4480), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5835) );
  OAI211_X1 U7369 ( .C1(n5844), .C2(n5839), .A(n6854), .B(n5868), .ZN(n5838)
         );
  INV_X1 U7370 ( .A(n5838), .ZN(n5859) );
  INV_X1 U7371 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n5842) );
  NAND2_X1 U7372 ( .A1(n5290), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5841) );
  NAND2_X1 U7373 ( .A1(n5305), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5840) );
  OAI211_X1 U7374 ( .C1(n5843), .C2(n5842), .A(n5841), .B(n5840), .ZN(n8629)
         );
  AND2_X1 U7375 ( .A1(n8851), .A2(n8629), .ZN(n5976) );
  INV_X1 U7376 ( .A(n5844), .ZN(n5857) );
  NAND2_X1 U7377 ( .A1(n5847), .A2(n5846), .ZN(n5848) );
  MUX2_X1 U7378 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6835), .Z(n5849) );
  XNOR2_X1 U7379 ( .A(n5849), .B(SI_31_), .ZN(n5850) );
  NAND2_X1 U7380 ( .A1(n8962), .A2(n4616), .ZN(n5853) );
  INV_X1 U7381 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5851) );
  OR2_X1 U7382 ( .A1(n5312), .A2(n5851), .ZN(n5852) );
  OR2_X1 U7383 ( .A1(n8844), .A2(n6854), .ZN(n5980) );
  INV_X1 U7384 ( .A(n8629), .ZN(n5854) );
  NAND2_X1 U7385 ( .A1(n5839), .A2(n5854), .ZN(n5855) );
  NAND2_X1 U7386 ( .A1(n5980), .A2(n5855), .ZN(n6010) );
  INV_X1 U7387 ( .A(n6010), .ZN(n5856) );
  NAND2_X1 U7388 ( .A1(n8844), .A2(n6854), .ZN(n5982) );
  OAI21_X1 U7389 ( .B1(n5859), .B2(n5858), .A(n5982), .ZN(n5860) );
  INV_X1 U7390 ( .A(n7741), .ZN(n7275) );
  NAND2_X1 U7391 ( .A1(n7275), .A2(n5868), .ZN(n6884) );
  NAND2_X1 U7392 ( .A1(n7337), .A2(n6884), .ZN(n5861) );
  NAND2_X1 U7393 ( .A1(n5868), .A2(n8797), .ZN(n5862) );
  OR2_X1 U7394 ( .A1(n5778), .A2(n5862), .ZN(n5981) );
  INV_X1 U7395 ( .A(n5997), .ZN(n5866) );
  NAND2_X1 U7396 ( .A1(n8561), .A2(n7203), .ZN(n5995) );
  AOI21_X1 U7397 ( .B1(n5868), .B2(n5995), .A(n5867), .ZN(n5870) );
  NAND2_X1 U7398 ( .A1(n5993), .A2(n5877), .ZN(n5869) );
  OAI211_X1 U7399 ( .C1(n5870), .C2(n5869), .A(n5981), .B(n5874), .ZN(n5871)
         );
  NAND2_X1 U7400 ( .A1(n5871), .A2(n7160), .ZN(n5872) );
  OAI22_X1 U7401 ( .A1(n5873), .A2(n4635), .B1(n5872), .B2(n5883), .ZN(n5880)
         );
  INV_X1 U7402 ( .A(n5993), .ZN(n5876) );
  INV_X1 U7403 ( .A(n5995), .ZN(n5875) );
  OAI211_X1 U7404 ( .C1(n5876), .C2(n5875), .A(n5994), .B(n5874), .ZN(n5878)
         );
  NAND3_X1 U7405 ( .A1(n5878), .A2(n4635), .A3(n5877), .ZN(n5879) );
  NAND2_X1 U7406 ( .A1(n5807), .A2(n8455), .ZN(n5881) );
  AOI22_X1 U7407 ( .A1(n5883), .A2(n5998), .B1(n5882), .B2(n5881), .ZN(n5886)
         );
  INV_X1 U7408 ( .A(n5884), .ZN(n5885) );
  MUX2_X1 U7409 ( .A(n5891), .B(n5890), .S(n5981), .Z(n5892) );
  MUX2_X1 U7410 ( .A(n5895), .B(n5894), .S(n5981), .Z(n5896) );
  NAND3_X1 U7411 ( .A1(n5901), .A2(n7650), .A3(n5992), .ZN(n5898) );
  INV_X1 U7412 ( .A(n5897), .ZN(n5990) );
  NAND3_X1 U7413 ( .A1(n5898), .A2(n5899), .A3(n5990), .ZN(n5905) );
  INV_X1 U7414 ( .A(n5992), .ZN(n5900) );
  OAI211_X1 U7415 ( .C1(n5901), .C2(n5900), .A(n5899), .B(n7603), .ZN(n5903)
         );
  NAND2_X1 U7416 ( .A1(n5903), .A2(n5902), .ZN(n5904) );
  NAND2_X1 U7417 ( .A1(n5907), .A2(n5991), .ZN(n5906) );
  NAND3_X1 U7418 ( .A1(n5907), .A2(n5990), .A3(n5988), .ZN(n5909) );
  INV_X1 U7419 ( .A(n5908), .ZN(n5989) );
  NAND2_X1 U7420 ( .A1(n5909), .A2(n5989), .ZN(n5910) );
  MUX2_X1 U7421 ( .A(n5913), .B(n5912), .S(n5981), .Z(n5914) );
  MUX2_X1 U7422 ( .A(n5918), .B(n5917), .S(n5981), .Z(n5919) );
  AOI21_X1 U7423 ( .B1(n5920), .B2(n5919), .A(n8020), .ZN(n5926) );
  INV_X1 U7424 ( .A(n5921), .ZN(n5924) );
  INV_X1 U7425 ( .A(n5922), .ZN(n5923) );
  MUX2_X1 U7426 ( .A(n5924), .B(n5923), .S(n5981), .Z(n5925) );
  NAND3_X1 U7427 ( .A1(n8064), .A2(n8607), .A3(n4635), .ZN(n5927) );
  AND2_X1 U7428 ( .A1(n8914), .A2(n8819), .ZN(n5931) );
  INV_X1 U7429 ( .A(n8064), .ZN(n8919) );
  INV_X1 U7430 ( .A(n8607), .ZN(n8547) );
  NAND3_X1 U7431 ( .A1(n8828), .A2(n8919), .A3(n8547), .ZN(n5928) );
  NAND3_X1 U7432 ( .A1(n5929), .A2(n5928), .A3(n4525), .ZN(n5930) );
  MUX2_X1 U7433 ( .A(n5931), .B(n5930), .S(n5981), .Z(n5932) );
  INV_X1 U7434 ( .A(n5938), .ZN(n5933) );
  NAND2_X1 U7435 ( .A1(n8770), .A2(n8749), .ZN(n5943) );
  NAND3_X1 U7436 ( .A1(n5942), .A2(n5941), .A3(n5940), .ZN(n5945) );
  INV_X1 U7437 ( .A(n5956), .ZN(n5948) );
  OAI211_X1 U7438 ( .C1(n4635), .C2(n5950), .A(n5949), .B(n5948), .ZN(n5954)
         );
  AOI21_X1 U7439 ( .B1(n5953), .B2(n5951), .A(n5981), .ZN(n5952) );
  AOI21_X1 U7440 ( .B1(n5954), .B2(n5953), .A(n5952), .ZN(n5955) );
  INV_X1 U7441 ( .A(n5815), .ZN(n8685) );
  NAND2_X1 U7442 ( .A1(n8667), .A2(n5957), .ZN(n5958) );
  MUX2_X1 U7443 ( .A(n8685), .B(n5958), .S(n5981), .Z(n5959) );
  MUX2_X1 U7444 ( .A(n5961), .B(n5960), .S(n5981), .Z(n5963) );
  INV_X1 U7445 ( .A(n8666), .ZN(n5962) );
  NAND2_X1 U7446 ( .A1(n5818), .A2(n5964), .ZN(n5967) );
  NAND2_X1 U7447 ( .A1(n8623), .A2(n5965), .ZN(n5966) );
  MUX2_X1 U7448 ( .A(n5967), .B(n5966), .S(n5981), .Z(n5968) );
  NAND2_X1 U7449 ( .A1(n5973), .A2(n5974), .ZN(n8626) );
  MUX2_X1 U7450 ( .A(n5974), .B(n5973), .S(n5981), .Z(n5975) );
  INV_X1 U7451 ( .A(n5976), .ZN(n5979) );
  NAND2_X1 U7452 ( .A1(n5978), .A2(n5977), .ZN(n5986) );
  NAND2_X1 U7453 ( .A1(n5982), .A2(n5979), .ZN(n6009) );
  NAND3_X1 U7454 ( .A1(n6009), .A2(n5981), .A3(n5980), .ZN(n5985) );
  INV_X1 U7455 ( .A(n5982), .ZN(n5983) );
  INV_X1 U7456 ( .A(n6885), .ZN(n6012) );
  INV_X1 U7457 ( .A(n8712), .ZN(n8709) );
  INV_X1 U7458 ( .A(n8697), .ZN(n8621) );
  NAND2_X1 U7459 ( .A1(n5989), .A2(n5988), .ZN(n7730) );
  NAND2_X1 U7460 ( .A1(n5991), .A2(n5990), .ZN(n7652) );
  INV_X1 U7461 ( .A(n7605), .ZN(n7598) );
  NAND2_X1 U7462 ( .A1(n5994), .A2(n5993), .ZN(n6880) );
  NAND2_X1 U7463 ( .A1(n6883), .A2(n5995), .ZN(n9948) );
  NOR4_X1 U7464 ( .A1(n7328), .A2(n6880), .A3(n9948), .A4(n7741), .ZN(n5996)
         );
  NAND3_X1 U7465 ( .A1(n5996), .A2(n5810), .A3(n7160), .ZN(n6000) );
  INV_X1 U7466 ( .A(n7424), .ZN(n5999) );
  NAND2_X1 U7467 ( .A1(n5998), .A2(n5997), .ZN(n7396) );
  NOR4_X1 U7468 ( .A1(n6000), .A2(n7403), .A3(n5999), .A4(n7396), .ZN(n6001)
         );
  NAND4_X1 U7469 ( .A1(n7598), .A2(n5811), .A3(n7546), .A4(n6001), .ZN(n6002)
         );
  NOR4_X1 U7470 ( .A1(n4670), .A2(n7730), .A3(n7652), .A4(n6002), .ZN(n6003)
         );
  NAND4_X1 U7471 ( .A1(n5011), .A2(n7941), .A3(n7917), .A4(n6003), .ZN(n6004)
         );
  NOR4_X1 U7472 ( .A1(n8612), .A2(n8816), .A3(n4911), .A4(n6004), .ZN(n6005)
         );
  NAND4_X1 U7473 ( .A1(n8734), .A2(n8613), .A3(n8747), .A4(n6005), .ZN(n6006)
         );
  NOR4_X1 U7474 ( .A1(n8709), .A2(n8621), .A3(n8760), .A4(n6006), .ZN(n6007)
         );
  NAND4_X1 U7475 ( .A1(n8666), .A2(n8623), .A3(n8688), .A4(n6007), .ZN(n6008)
         );
  XNOR2_X1 U7476 ( .A(n6011), .B(n8835), .ZN(n6013) );
  AOI22_X1 U7477 ( .A1(n6013), .A2(n7782), .B1(n6012), .B2(n7741), .ZN(n6014)
         );
  OR2_X1 U7478 ( .A1(n6015), .A2(P2_U3152), .ZN(n7959) );
  INV_X1 U7479 ( .A(n7959), .ZN(n6016) );
  INV_X1 U7480 ( .A(n8977), .ZN(n8599) );
  NAND4_X1 U7481 ( .A1(n9938), .A2(n6017), .A3(n8599), .A4(n8750), .ZN(n6018)
         );
  OAI211_X1 U7482 ( .C1(n5778), .C2(n7959), .A(n6018), .B(P2_B_REG_SCAN_IN), 
        .ZN(n6019) );
  NAND2_X1 U7483 ( .A1(n6067), .A2(n6020), .ZN(n6106) );
  INV_X1 U7484 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6033) );
  NAND2_X1 U7485 ( .A1(n6034), .A2(n6033), .ZN(n9537) );
  INV_X1 U7486 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6035) );
  INV_X1 U7487 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7513) );
  OR2_X2 U7488 ( .A1(n6037), .A2(n6036), .ZN(n6145) );
  INV_X1 U7489 ( .A(n6145), .ZN(n6128) );
  INV_X1 U7490 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6038) );
  OAI21_X1 U7491 ( .B1(n6045), .B2(n9536), .A(P1_IR_REG_20__SCAN_IN), .ZN(
        n6047) );
  NAND2_X1 U7492 ( .A1(n6047), .A2(n6046), .ZN(n6049) );
  NAND2_X1 U7493 ( .A1(n6058), .A2(n6057), .ZN(n6051) );
  INV_X1 U7494 ( .A(n6054), .ZN(n6653) );
  NAND2_X1 U7495 ( .A1(n6653), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6056) );
  NAND2_X1 U7496 ( .A1(n6695), .A2(n4481), .ZN(n6072) );
  NAND2_X1 U7497 ( .A1(n6062), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6064) );
  XNOR2_X2 U7498 ( .A(n6064), .B(n6063), .ZN(n8430) );
  INV_X1 U7499 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7500 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6066) );
  INV_X1 U7501 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n10369) );
  MUX2_X1 U7502 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6066), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n6069) );
  INV_X1 U7503 ( .A(n6067), .ZN(n6068) );
  NAND2_X1 U7504 ( .A1(n6069), .A2(n6068), .ZN(n6830) );
  AND2_X4 U7505 ( .A1(n6800), .A2(n6672), .ZN(n6521) );
  NAND2_X1 U7506 ( .A1(n6694), .A2(n6521), .ZN(n6071) );
  NAND2_X1 U7507 ( .A1(n6074), .A2(n6073), .ZN(n6075) );
  NAND2_X1 U7508 ( .A1(n6075), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U7509 ( .A1(n6078), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U7510 ( .A1(n7915), .A2(n6678), .ZN(n6081) );
  AND2_X2 U7511 ( .A1(n6521), .A2(n6081), .ZN(n6486) );
  NAND2_X1 U7512 ( .A1(n9139), .A2(n6486), .ZN(n6083) );
  NAND2_X1 U7513 ( .A1(n6694), .A2(n4486), .ZN(n6082) );
  NAND2_X1 U7514 ( .A1(n6083), .A2(n6082), .ZN(n6101) );
  NAND2_X1 U7515 ( .A1(n6100), .A2(n6101), .ZN(n6099) );
  INV_X1 U7516 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6084) );
  OR2_X1 U7517 ( .A1(n6126), .A2(n6084), .ZN(n6089) );
  INV_X1 U7518 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9688) );
  OR2_X1 U7519 ( .A1(n6127), .A2(n9688), .ZN(n6088) );
  NAND2_X1 U7520 ( .A1(n6453), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6087) );
  INV_X1 U7521 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6085) );
  OR2_X1 U7522 ( .A1(n6145), .A2(n6085), .ZN(n6086) );
  NAND2_X1 U7523 ( .A1(n6696), .A2(n6486), .ZN(n6094) );
  INV_X1 U7524 ( .A(n6090), .ZN(n6091) );
  XNOR2_X1 U7525 ( .A(n6091), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n6832) );
  MUX2_X1 U7526 ( .A(P1_IR_REG_0__SCAN_IN), .B(n6832), .S(n8130), .Z(n7538) );
  INV_X1 U7527 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10433) );
  NOR2_X1 U7528 ( .A1(n6800), .A2(n10433), .ZN(n6092) );
  AOI21_X1 U7529 ( .B1(n7538), .B2(n4484), .A(n6092), .ZN(n6093) );
  NAND2_X1 U7530 ( .A1(n6696), .A2(n4485), .ZN(n6097) );
  INV_X1 U7531 ( .A(n6800), .ZN(n6095) );
  AOI22_X1 U7532 ( .A1(n7538), .A2(n6521), .B1(n6095), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n6096) );
  NAND2_X1 U7533 ( .A1(n6097), .A2(n6096), .ZN(n6804) );
  NAND2_X1 U7534 ( .A1(n6805), .A2(n6804), .ZN(n6803) );
  INV_X1 U7535 ( .A(n7492), .ZN(n6160) );
  NAND2_X1 U7536 ( .A1(n6803), .A2(n6098), .ZN(n7239) );
  NAND2_X1 U7537 ( .A1(n6099), .A2(n7239), .ZN(n6103) );
  INV_X1 U7538 ( .A(n6101), .ZN(n7238) );
  NAND2_X1 U7539 ( .A1(n7241), .A2(n7238), .ZN(n6102) );
  NAND2_X1 U7540 ( .A1(n6103), .A2(n6102), .ZN(n7233) );
  NOR2_X1 U7541 ( .A1(n6067), .A2(n9536), .ZN(n6104) );
  MUX2_X1 U7542 ( .A(n9536), .B(n6104), .S(P1_IR_REG_2__SCAN_IN), .Z(n6105) );
  INV_X1 U7543 ( .A(n6105), .ZN(n6107) );
  NAND2_X1 U7544 ( .A1(n6107), .A2(n6106), .ZN(n6962) );
  INV_X1 U7545 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6834) );
  OR2_X1 U7546 ( .A1(n6180), .A2(n6834), .ZN(n6109) );
  OR2_X1 U7547 ( .A1(n6155), .A2(n6848), .ZN(n6108) );
  NAND2_X1 U7548 ( .A1(n4479), .A2(n6521), .ZN(n6116) );
  NAND2_X1 U7549 ( .A1(n6453), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6114) );
  INV_X1 U7550 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6961) );
  INV_X1 U7551 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6956) );
  OR2_X1 U7552 ( .A1(n6126), .A2(n6956), .ZN(n6112) );
  INV_X1 U7553 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6110) );
  OR2_X1 U7554 ( .A1(n6145), .A2(n6110), .ZN(n6111) );
  NAND2_X1 U7555 ( .A1(n9138), .A2(n4482), .ZN(n6115) );
  NAND2_X1 U7556 ( .A1(n6116), .A2(n6115), .ZN(n6117) );
  AND2_X1 U7557 ( .A1(n4479), .A2(n4486), .ZN(n6119) );
  AOI21_X1 U7558 ( .B1(n9138), .B2(n6486), .A(n6119), .ZN(n6121) );
  XNOR2_X1 U7559 ( .A(n6120), .B(n6121), .ZN(n7234) );
  NAND2_X1 U7560 ( .A1(n7233), .A2(n7234), .ZN(n6124) );
  INV_X1 U7561 ( .A(n6120), .ZN(n6122) );
  NAND2_X1 U7562 ( .A1(n6122), .A2(n6121), .ZN(n6123) );
  NAND2_X1 U7563 ( .A1(n6124), .A2(n6123), .ZN(n7246) );
  OR2_X1 U7564 ( .A1(n6587), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6132) );
  INV_X1 U7565 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7018) );
  INV_X1 U7566 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7003) );
  OR2_X1 U7567 ( .A1(n6127), .A2(n7003), .ZN(n6130) );
  NAND2_X1 U7568 ( .A1(n6128), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6129) );
  NAND2_X1 U7569 ( .A1(n6701), .A2(n4481), .ZN(n6137) );
  NAND2_X1 U7570 ( .A1(n6106), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6133) );
  XNOR2_X1 U7571 ( .A(n6133), .B(n6021), .ZN(n7017) );
  INV_X1 U7572 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6839) );
  OR2_X1 U7573 ( .A1(n6180), .A2(n6839), .ZN(n6135) );
  OR2_X1 U7574 ( .A1(n6155), .A2(n6845), .ZN(n6134) );
  OAI211_X1 U7575 ( .C1(n8130), .C2(n7017), .A(n6135), .B(n6134), .ZN(n6702)
         );
  NAND2_X1 U7576 ( .A1(n6702), .A2(n6521), .ZN(n6136) );
  NAND2_X1 U7577 ( .A1(n6137), .A2(n6136), .ZN(n6138) );
  AND2_X1 U7578 ( .A1(n6702), .A2(n4482), .ZN(n6139) );
  AOI21_X1 U7579 ( .B1(n6701), .B2(n6628), .A(n6139), .ZN(n6141) );
  XNOR2_X1 U7580 ( .A(n6140), .B(n6141), .ZN(n7247) );
  NAND2_X1 U7581 ( .A1(n7246), .A2(n7247), .ZN(n6144) );
  INV_X1 U7582 ( .A(n6140), .ZN(n6142) );
  NAND2_X1 U7583 ( .A1(n6142), .A2(n6141), .ZN(n6143) );
  NAND2_X1 U7584 ( .A1(n6144), .A2(n6143), .ZN(n7318) );
  INV_X1 U7585 ( .A(n7318), .ZN(n6164) );
  INV_X1 U7586 ( .A(n6127), .ZN(n6497) );
  NAND2_X1 U7587 ( .A1(n6497), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6151) );
  INV_X1 U7588 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6146) );
  OR2_X1 U7589 ( .A1(n6145), .A2(n6146), .ZN(n6150) );
  XNOR2_X1 U7590 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n7322) );
  OR2_X1 U7591 ( .A1(n6587), .A2(n7322), .ZN(n6149) );
  INV_X1 U7592 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6147) );
  OR2_X1 U7593 ( .A1(n6501), .A2(n6147), .ZN(n6148) );
  NAND2_X1 U7594 ( .A1(n9137), .A2(n4486), .ZN(n6159) );
  NAND2_X1 U7595 ( .A1(n6152), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6154) );
  INV_X1 U7596 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6153) );
  XNOR2_X1 U7597 ( .A(n6154), .B(n6153), .ZN(n7019) );
  OR2_X1 U7598 ( .A1(n6180), .A2(n6840), .ZN(n6157) );
  OR2_X1 U7599 ( .A1(n6155), .A2(n6842), .ZN(n6156) );
  OAI211_X1 U7600 ( .C1(n8130), .C2(n7019), .A(n6157), .B(n6156), .ZN(n7661)
         );
  NAND2_X1 U7601 ( .A1(n7661), .A2(n6521), .ZN(n6158) );
  NAND2_X1 U7602 ( .A1(n6159), .A2(n6158), .ZN(n6161) );
  XNOR2_X1 U7603 ( .A(n6161), .B(n6556), .ZN(n6165) );
  AND2_X1 U7604 ( .A1(n7661), .A2(n4484), .ZN(n6162) );
  AOI21_X1 U7605 ( .B1(n9137), .B2(n6628), .A(n6162), .ZN(n6166) );
  XNOR2_X1 U7606 ( .A(n6165), .B(n6166), .ZN(n7321) );
  NAND2_X1 U7607 ( .A1(n6164), .A2(n6163), .ZN(n7319) );
  INV_X1 U7608 ( .A(n6165), .ZN(n6168) );
  INV_X1 U7609 ( .A(n6166), .ZN(n6167) );
  NAND2_X1 U7610 ( .A1(n6168), .A2(n6167), .ZN(n6169) );
  NAND2_X1 U7611 ( .A1(n6128), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6177) );
  INV_X1 U7612 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6170) );
  OR2_X1 U7613 ( .A1(n6501), .A2(n6170), .ZN(n6176) );
  NAND3_X1 U7614 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6192) );
  INV_X1 U7615 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6172) );
  NAND2_X1 U7616 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6171) );
  NAND2_X1 U7617 ( .A1(n6172), .A2(n6171), .ZN(n6173) );
  NAND2_X1 U7618 ( .A1(n6192), .A2(n6173), .ZN(n7503) );
  OR2_X1 U7619 ( .A1(n6587), .A2(n7503), .ZN(n6175) );
  INV_X1 U7620 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7007) );
  OR2_X1 U7621 ( .A1(n6458), .A2(n7007), .ZN(n6174) );
  NAND4_X1 U7622 ( .A1(n6177), .A2(n6176), .A3(n6175), .A4(n6174), .ZN(n9136)
         );
  NAND2_X1 U7623 ( .A1(n9136), .A2(n4485), .ZN(n6184) );
  OR2_X1 U7624 ( .A1(n6178), .A2(n9536), .ZN(n6179) );
  XNOR2_X1 U7625 ( .A(n6179), .B(P1_IR_REG_5__SCAN_IN), .ZN(n7021) );
  INV_X1 U7626 ( .A(n7021), .ZN(n9696) );
  OR2_X1 U7627 ( .A1(n6155), .A2(n6851), .ZN(n6182) );
  INV_X1 U7628 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6850) );
  OR2_X1 U7629 ( .A1(n8134), .A2(n6850), .ZN(n6181) );
  OAI211_X1 U7630 ( .C1(n8130), .C2(n9696), .A(n6182), .B(n6181), .ZN(n6768)
         );
  NAND2_X1 U7631 ( .A1(n6768), .A2(n6521), .ZN(n6183) );
  NAND2_X1 U7632 ( .A1(n9136), .A2(n6486), .ZN(n6186) );
  NAND2_X1 U7633 ( .A1(n6768), .A2(n4482), .ZN(n6185) );
  NAND2_X1 U7634 ( .A1(n6186), .A2(n6185), .ZN(n6187) );
  INV_X1 U7635 ( .A(n7308), .ZN(n6188) );
  INV_X1 U7636 ( .A(n6187), .ZN(n7307) );
  NAND2_X1 U7637 ( .A1(n6188), .A2(n7307), .ZN(n6189) );
  NAND2_X1 U7638 ( .A1(n6666), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6197) );
  INV_X1 U7639 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6190) );
  OR2_X1 U7640 ( .A1(n6458), .A2(n6190), .ZN(n6196) );
  INV_X1 U7641 ( .A(n6192), .ZN(n6191) );
  NAND2_X1 U7642 ( .A1(n6191), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6210) );
  INV_X1 U7643 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7073) );
  NAND2_X1 U7644 ( .A1(n6192), .A2(n7073), .ZN(n6193) );
  NAND2_X1 U7645 ( .A1(n6210), .A2(n6193), .ZN(n7683) );
  OR2_X1 U7646 ( .A1(n6587), .A2(n7683), .ZN(n6195) );
  INV_X1 U7647 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7684) );
  OR2_X1 U7648 ( .A1(n6501), .A2(n7684), .ZN(n6194) );
  NAND2_X1 U7649 ( .A1(n9135), .A2(n4486), .ZN(n6203) );
  NAND2_X1 U7650 ( .A1(n6178), .A2(n6198), .ZN(n6216) );
  NAND2_X1 U7651 ( .A1(n6216), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6199) );
  XNOR2_X1 U7652 ( .A(n6199), .B(P1_IR_REG_6__SCAN_IN), .ZN(n7023) );
  INV_X1 U7653 ( .A(n7023), .ZN(n7075) );
  INV_X1 U7654 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10101) );
  OR2_X1 U7655 ( .A1(n8134), .A2(n10101), .ZN(n6200) );
  NAND2_X1 U7656 ( .A1(n7784), .A2(n6521), .ZN(n6202) );
  NAND2_X1 U7657 ( .A1(n6203), .A2(n6202), .ZN(n6204) );
  XNOR2_X1 U7658 ( .A(n6204), .B(n6556), .ZN(n7522) );
  NAND2_X1 U7659 ( .A1(n9135), .A2(n6486), .ZN(n6206) );
  NAND2_X1 U7660 ( .A1(n7784), .A2(n4481), .ZN(n6205) );
  NAND2_X1 U7661 ( .A1(n6206), .A2(n6205), .ZN(n7521) );
  NAND2_X1 U7662 ( .A1(n6666), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6215) );
  INV_X1 U7663 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6207) );
  OR2_X1 U7664 ( .A1(n6458), .A2(n6207), .ZN(n6214) );
  INV_X1 U7665 ( .A(n6210), .ZN(n6208) );
  NAND2_X1 U7666 ( .A1(n6208), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6232) );
  INV_X1 U7667 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U7668 ( .A1(n6210), .A2(n6209), .ZN(n6211) );
  NAND2_X1 U7669 ( .A1(n6232), .A2(n6211), .ZN(n7588) );
  OR2_X1 U7670 ( .A1(n6587), .A2(n7588), .ZN(n6213) );
  INV_X1 U7671 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7562) );
  OR2_X1 U7672 ( .A1(n6501), .A2(n7562), .ZN(n6212) );
  NAND4_X1 U7673 ( .A1(n6215), .A2(n6214), .A3(n6213), .A4(n6212), .ZN(n9134)
         );
  NAND2_X1 U7674 ( .A1(n9134), .A2(n4485), .ZN(n6222) );
  INV_X1 U7675 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10232) );
  NAND2_X1 U7676 ( .A1(n6227), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6217) );
  XNOR2_X1 U7677 ( .A(n6217), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7050) );
  INV_X1 U7678 ( .A(n7050), .ZN(n7010) );
  OAI22_X1 U7679 ( .A1(n8134), .A2(n10232), .B1(n8130), .B2(n7010), .ZN(n6218)
         );
  INV_X1 U7680 ( .A(n6218), .ZN(n6220) );
  INV_X2 U7681 ( .A(n6155), .ZN(n6244) );
  NAND2_X1 U7682 ( .A1(n6861), .A2(n6244), .ZN(n6219) );
  NAND2_X1 U7683 ( .A1(n6220), .A2(n6219), .ZN(n7625) );
  NAND2_X1 U7684 ( .A1(n7625), .A2(n6521), .ZN(n6221) );
  NAND2_X1 U7685 ( .A1(n6222), .A2(n6221), .ZN(n6223) );
  XNOR2_X1 U7686 ( .A(n6223), .B(n6556), .ZN(n6225) );
  AOI22_X1 U7687 ( .A1(n9134), .A2(n6486), .B1(n4482), .B2(n7625), .ZN(n6224)
         );
  OR2_X1 U7688 ( .A1(n6225), .A2(n6224), .ZN(n7586) );
  NAND2_X1 U7689 ( .A1(n7584), .A2(n7586), .ZN(n6226) );
  NAND2_X1 U7690 ( .A1(n6225), .A2(n6224), .ZN(n7585) );
  NAND2_X1 U7691 ( .A1(n6865), .A2(n6244), .ZN(n6230) );
  OAI21_X1 U7692 ( .B1(n6227), .B2(P1_IR_REG_7__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6228) );
  XNOR2_X1 U7693 ( .A(n6228), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7051) );
  AOI22_X1 U7694 ( .A1(n6450), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6449), .B2(
        n7051), .ZN(n6229) );
  NAND2_X1 U7695 ( .A1(n6230), .A2(n6229), .ZN(n7840) );
  NAND2_X1 U7696 ( .A1(n7840), .A2(n4481), .ZN(n6239) );
  NAND2_X1 U7697 ( .A1(n6666), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6237) );
  OR2_X1 U7698 ( .A1(n6458), .A2(n7847), .ZN(n6236) );
  INV_X1 U7699 ( .A(n6232), .ZN(n6231) );
  NAND2_X1 U7700 ( .A1(n6231), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6249) );
  INV_X1 U7701 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7798) );
  NAND2_X1 U7702 ( .A1(n6232), .A2(n7798), .ZN(n6233) );
  NAND2_X1 U7703 ( .A1(n6249), .A2(n6233), .ZN(n7800) );
  OR2_X1 U7704 ( .A1(n6587), .A2(n7800), .ZN(n6235) );
  INV_X1 U7705 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7760) );
  OR2_X1 U7706 ( .A1(n6501), .A2(n7760), .ZN(n6234) );
  NAND4_X1 U7707 ( .A1(n6237), .A2(n6236), .A3(n6235), .A4(n6234), .ZN(n9133)
         );
  NAND2_X1 U7708 ( .A1(n9133), .A2(n6486), .ZN(n6238) );
  AND2_X1 U7709 ( .A1(n6239), .A2(n6238), .ZN(n6243) );
  NAND2_X1 U7710 ( .A1(n7840), .A2(n6521), .ZN(n6241) );
  NAND2_X1 U7711 ( .A1(n9133), .A2(n4486), .ZN(n6240) );
  NAND2_X1 U7712 ( .A1(n6241), .A2(n6240), .ZN(n6242) );
  XNOR2_X1 U7713 ( .A(n6242), .B(n7492), .ZN(n7795) );
  NAND2_X1 U7714 ( .A1(n6869), .A2(n6244), .ZN(n6247) );
  OR2_X1 U7715 ( .A1(n4522), .A2(n9536), .ZN(n6245) );
  XNOR2_X1 U7716 ( .A(n6245), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7053) );
  AOI22_X1 U7717 ( .A1(n6450), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6449), .B2(
        n7053), .ZN(n6246) );
  NAND2_X1 U7718 ( .A1(n9825), .A2(n6521), .ZN(n6257) );
  NAND2_X1 U7719 ( .A1(n6666), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U7720 ( .A1(n6249), .A2(n6248), .ZN(n6250) );
  NAND2_X1 U7721 ( .A1(n6267), .A2(n6250), .ZN(n7858) );
  OR2_X1 U7722 ( .A1(n6587), .A2(n7858), .ZN(n6254) );
  INV_X1 U7723 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7859) );
  OR2_X1 U7724 ( .A1(n6501), .A2(n7859), .ZN(n6253) );
  INV_X1 U7725 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6251) );
  OR2_X1 U7726 ( .A1(n6458), .A2(n6251), .ZN(n6252) );
  NAND4_X1 U7727 ( .A1(n6255), .A2(n6254), .A3(n6253), .A4(n6252), .ZN(n9132)
         );
  NAND2_X1 U7728 ( .A1(n9132), .A2(n4484), .ZN(n6256) );
  NAND2_X1 U7729 ( .A1(n6257), .A2(n6256), .ZN(n6258) );
  XNOR2_X1 U7730 ( .A(n6258), .B(n6556), .ZN(n6261) );
  AND2_X1 U7731 ( .A1(n9132), .A2(n6628), .ZN(n6259) );
  AOI21_X1 U7732 ( .B1(n9825), .B2(n4486), .A(n6259), .ZN(n6260) );
  XNOR2_X1 U7733 ( .A(n6261), .B(n6260), .ZN(n7832) );
  NAND2_X1 U7734 ( .A1(n6261), .A2(n6260), .ZN(n6262) );
  NAND2_X1 U7735 ( .A1(n6873), .A2(n6244), .ZN(n6265) );
  NAND2_X1 U7736 ( .A1(n4522), .A2(n6263), .ZN(n6304) );
  NAND2_X1 U7737 ( .A1(n6304), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6279) );
  XNOR2_X1 U7738 ( .A(n6279), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7055) );
  AOI22_X1 U7739 ( .A1(n6450), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6449), .B2(
        n7055), .ZN(n6264) );
  NAND2_X1 U7740 ( .A1(n7895), .A2(n6521), .ZN(n6274) );
  NAND2_X1 U7741 ( .A1(n6666), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6272) );
  INV_X1 U7742 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6266) );
  OR2_X1 U7743 ( .A1(n6458), .A2(n6266), .ZN(n6271) );
  NAND2_X1 U7744 ( .A1(n6267), .A2(n7126), .ZN(n6268) );
  NAND2_X1 U7745 ( .A1(n6287), .A2(n6268), .ZN(n7892) );
  OR2_X1 U7746 ( .A1(n6587), .A2(n7892), .ZN(n6270) );
  INV_X1 U7747 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7813) );
  OR2_X1 U7748 ( .A1(n6501), .A2(n7813), .ZN(n6269) );
  NAND4_X1 U7749 ( .A1(n6272), .A2(n6271), .A3(n6270), .A4(n6269), .ZN(n9131)
         );
  NAND2_X1 U7750 ( .A1(n9131), .A2(n4486), .ZN(n6273) );
  NAND2_X1 U7751 ( .A1(n6274), .A2(n6273), .ZN(n6275) );
  XNOR2_X1 U7752 ( .A(n6275), .B(n6556), .ZN(n7888) );
  AND2_X1 U7753 ( .A1(n9131), .A2(n6628), .ZN(n6276) );
  AOI21_X1 U7754 ( .B1(n7895), .B2(n4485), .A(n6276), .ZN(n7887) );
  AND2_X1 U7755 ( .A1(n7888), .A2(n7887), .ZN(n6277) );
  NAND2_X1 U7756 ( .A1(n6975), .A2(n6244), .ZN(n6283) );
  INV_X1 U7757 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6278) );
  NAND2_X1 U7758 ( .A1(n6279), .A2(n6278), .ZN(n6280) );
  NAND2_X1 U7759 ( .A1(n6280), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6281) );
  XNOR2_X1 U7760 ( .A(n6281), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7714) );
  AOI22_X1 U7761 ( .A1(n6450), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6449), .B2(
        n7714), .ZN(n6282) );
  NAND2_X1 U7762 ( .A1(n7935), .A2(n6521), .ZN(n6294) );
  NAND2_X1 U7763 ( .A1(n6666), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6292) );
  INV_X1 U7764 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6284) );
  OR2_X1 U7765 ( .A1(n6458), .A2(n6284), .ZN(n6291) );
  INV_X1 U7766 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6286) );
  NAND2_X1 U7767 ( .A1(n6287), .A2(n6286), .ZN(n6288) );
  NAND2_X1 U7768 ( .A1(n6309), .A2(n6288), .ZN(n9656) );
  OR2_X1 U7769 ( .A1(n6587), .A2(n9656), .ZN(n6290) );
  INV_X1 U7770 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9657) );
  OR2_X1 U7771 ( .A1(n6501), .A2(n9657), .ZN(n6289) );
  NAND4_X1 U7772 ( .A1(n6292), .A2(n6291), .A3(n6290), .A4(n6289), .ZN(n9130)
         );
  NAND2_X1 U7773 ( .A1(n9130), .A2(n4484), .ZN(n6293) );
  NAND2_X1 U7774 ( .A1(n6294), .A2(n6293), .ZN(n6295) );
  XNOR2_X1 U7775 ( .A(n6295), .B(n7492), .ZN(n6299) );
  AND2_X1 U7776 ( .A1(n9130), .A2(n6628), .ZN(n6296) );
  AOI21_X1 U7777 ( .B1(n7935), .B2(n4486), .A(n6296), .ZN(n6297) );
  XNOR2_X1 U7778 ( .A(n6299), .B(n6297), .ZN(n7931) );
  NAND2_X1 U7779 ( .A1(n7932), .A2(n7931), .ZN(n6301) );
  INV_X1 U7780 ( .A(n6297), .ZN(n6298) );
  NAND2_X1 U7781 ( .A1(n6299), .A2(n6298), .ZN(n6300) );
  NAND2_X1 U7782 ( .A1(n6301), .A2(n6300), .ZN(n7992) );
  INV_X1 U7783 ( .A(n7992), .ZN(n6325) );
  NAND2_X1 U7784 ( .A1(n7104), .A2(n6244), .ZN(n6307) );
  INV_X1 U7785 ( .A(n6302), .ZN(n6303) );
  NAND2_X1 U7786 ( .A1(n6327), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6305) );
  XNOR2_X1 U7787 ( .A(n6305), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9734) );
  AOI22_X1 U7788 ( .A1(n6450), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6449), .B2(
        n9734), .ZN(n6306) );
  NAND2_X1 U7789 ( .A1(n7999), .A2(n6521), .ZN(n6316) );
  NAND2_X1 U7790 ( .A1(n6666), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6314) );
  INV_X1 U7791 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7969) );
  OR2_X1 U7792 ( .A1(n6501), .A2(n7969), .ZN(n6313) );
  INV_X1 U7793 ( .A(n6309), .ZN(n6308) );
  NAND2_X1 U7794 ( .A1(n6308), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6332) );
  INV_X1 U7795 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7996) );
  NAND2_X1 U7796 ( .A1(n6309), .A2(n7996), .ZN(n6310) );
  NAND2_X1 U7797 ( .A1(n6332), .A2(n6310), .ZN(n7997) );
  OR2_X1 U7798 ( .A1(n6587), .A2(n7997), .ZN(n6312) );
  INV_X1 U7799 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7706) );
  OR2_X1 U7800 ( .A1(n6458), .A2(n7706), .ZN(n6311) );
  NAND4_X1 U7801 ( .A1(n6314), .A2(n6313), .A3(n6312), .A4(n6311), .ZN(n9129)
         );
  NAND2_X1 U7802 ( .A1(n9129), .A2(n4481), .ZN(n6315) );
  NAND2_X1 U7803 ( .A1(n6316), .A2(n6315), .ZN(n6317) );
  XNOR2_X1 U7804 ( .A(n6317), .B(n6556), .ZN(n6319) );
  AND2_X1 U7805 ( .A1(n9129), .A2(n6628), .ZN(n6318) );
  AOI21_X1 U7806 ( .B1(n7999), .B2(n4482), .A(n6318), .ZN(n6320) );
  NAND2_X1 U7807 ( .A1(n6319), .A2(n6320), .ZN(n6326) );
  INV_X1 U7808 ( .A(n6319), .ZN(n6322) );
  INV_X1 U7809 ( .A(n6320), .ZN(n6321) );
  NAND2_X1 U7810 ( .A1(n6322), .A2(n6321), .ZN(n6323) );
  NAND2_X1 U7811 ( .A1(n6326), .A2(n6323), .ZN(n7995) );
  INV_X1 U7812 ( .A(n7995), .ZN(n6324) );
  NAND2_X1 U7813 ( .A1(n7174), .A2(n6244), .ZN(n6330) );
  NAND2_X1 U7814 ( .A1(n6346), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6328) );
  XNOR2_X1 U7815 ( .A(n6328), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9747) );
  AOI22_X1 U7816 ( .A1(n6450), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6449), .B2(
        n9747), .ZN(n6329) );
  NAND2_X1 U7817 ( .A1(n8167), .A2(n6521), .ZN(n6339) );
  NAND2_X1 U7818 ( .A1(n6666), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6337) );
  INV_X1 U7819 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7708) );
  OR2_X1 U7820 ( .A1(n6458), .A2(n7708), .ZN(n6336) );
  NAND2_X1 U7821 ( .A1(n6332), .A2(n6331), .ZN(n6333) );
  NAND2_X1 U7822 ( .A1(n6352), .A2(n6333), .ZN(n8040) );
  OR2_X1 U7823 ( .A1(n6587), .A2(n8040), .ZN(n6335) );
  INV_X1 U7824 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7983) );
  OR2_X1 U7825 ( .A1(n6501), .A2(n7983), .ZN(n6334) );
  NAND4_X1 U7826 ( .A1(n6337), .A2(n6336), .A3(n6335), .A4(n6334), .ZN(n9128)
         );
  NAND2_X1 U7827 ( .A1(n9128), .A2(n4486), .ZN(n6338) );
  NAND2_X1 U7828 ( .A1(n6339), .A2(n6338), .ZN(n6340) );
  XNOR2_X1 U7829 ( .A(n6340), .B(n6556), .ZN(n6342) );
  AND2_X1 U7830 ( .A1(n9128), .A2(n6628), .ZN(n6341) );
  AOI21_X1 U7831 ( .B1(n8167), .B2(n4485), .A(n6341), .ZN(n6343) );
  AND2_X1 U7832 ( .A1(n6342), .A2(n6343), .ZN(n8036) );
  INV_X1 U7833 ( .A(n6342), .ZN(n6345) );
  INV_X1 U7834 ( .A(n6343), .ZN(n6344) );
  NAND2_X1 U7835 ( .A1(n7183), .A2(n6244), .ZN(n6348) );
  OAI21_X1 U7836 ( .B1(n6346), .B2(P1_IR_REG_13__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6366) );
  XNOR2_X1 U7837 ( .A(n6366), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7720) );
  AOI22_X1 U7838 ( .A1(n6450), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6449), .B2(
        n7720), .ZN(n6347) );
  NAND2_X1 U7839 ( .A1(n9007), .A2(n6521), .ZN(n6359) );
  NAND2_X1 U7840 ( .A1(n6666), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6357) );
  INV_X1 U7841 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6349) );
  OR2_X1 U7842 ( .A1(n6458), .A2(n6349), .ZN(n6356) );
  INV_X1 U7843 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6351) );
  NAND2_X1 U7844 ( .A1(n6352), .A2(n6351), .ZN(n6353) );
  NAND2_X1 U7845 ( .A1(n6373), .A2(n6353), .ZN(n9004) );
  OR2_X1 U7846 ( .A1(n6587), .A2(n9004), .ZN(n6355) );
  INV_X1 U7847 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8014) );
  OR2_X1 U7848 ( .A1(n6501), .A2(n8014), .ZN(n6354) );
  NAND4_X1 U7849 ( .A1(n6357), .A2(n6356), .A3(n6355), .A4(n6354), .ZN(n9127)
         );
  NAND2_X1 U7850 ( .A1(n9127), .A2(n4484), .ZN(n6358) );
  NAND2_X1 U7851 ( .A1(n6359), .A2(n6358), .ZN(n6360) );
  NAND2_X1 U7852 ( .A1(n9007), .A2(n4485), .ZN(n6362) );
  NAND2_X1 U7853 ( .A1(n9127), .A2(n6486), .ZN(n6361) );
  NAND2_X1 U7854 ( .A1(n6362), .A2(n6361), .ZN(n9000) );
  NAND2_X1 U7855 ( .A1(n8997), .A2(n9000), .ZN(n6364) );
  NAND2_X1 U7856 ( .A1(n6363), .A2(n4575), .ZN(n8998) );
  NAND2_X1 U7857 ( .A1(n7259), .A2(n6244), .ZN(n6370) );
  INV_X1 U7858 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6365) );
  NAND2_X1 U7859 ( .A1(n6366), .A2(n6365), .ZN(n6367) );
  NAND2_X1 U7860 ( .A1(n6367), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6368) );
  XNOR2_X1 U7861 ( .A(n6368), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9759) );
  AOI22_X1 U7862 ( .A1(n6450), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6449), .B2(
        n9759), .ZN(n6369) );
  NAND2_X1 U7863 ( .A1(n6770), .A2(n6521), .ZN(n6380) );
  NAND2_X1 U7864 ( .A1(n6666), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6378) );
  INV_X1 U7865 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n6371) );
  OR2_X1 U7866 ( .A1(n6458), .A2(n6371), .ZN(n6377) );
  NAND2_X1 U7867 ( .A1(n6373), .A2(n6372), .ZN(n6374) );
  NAND2_X1 U7868 ( .A1(n6392), .A2(n6374), .ZN(n9629) );
  OR2_X1 U7869 ( .A1(n6587), .A2(n9629), .ZN(n6376) );
  INV_X1 U7870 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9630) );
  OR2_X1 U7871 ( .A1(n6501), .A2(n9630), .ZN(n6375) );
  NAND4_X1 U7872 ( .A1(n6378), .A2(n6377), .A3(n6376), .A4(n6375), .ZN(n9381)
         );
  NAND2_X1 U7873 ( .A1(n9381), .A2(n4481), .ZN(n6379) );
  NAND2_X1 U7874 ( .A1(n6380), .A2(n6379), .ZN(n6381) );
  XNOR2_X1 U7875 ( .A(n6381), .B(n6556), .ZN(n9113) );
  AND2_X1 U7876 ( .A1(n9381), .A2(n6628), .ZN(n6382) );
  AOI21_X1 U7877 ( .B1(n6770), .B2(n4485), .A(n6382), .ZN(n9112) );
  NAND2_X1 U7878 ( .A1(n9113), .A2(n9112), .ZN(n6383) );
  INV_X1 U7879 ( .A(n9113), .ZN(n6385) );
  INV_X1 U7880 ( .A(n9112), .ZN(n6384) );
  NAND2_X1 U7881 ( .A1(n6385), .A2(n6384), .ZN(n6386) );
  NAND2_X1 U7882 ( .A1(n7316), .A2(n6244), .ZN(n6390) );
  NAND2_X1 U7883 ( .A1(n6387), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6388) );
  XNOR2_X1 U7884 ( .A(n6388), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9770) );
  AOI22_X1 U7885 ( .A1(n6450), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6449), .B2(
        n9770), .ZN(n6389) );
  NAND2_X1 U7886 ( .A1(n9390), .A2(n6521), .ZN(n6399) );
  NAND2_X1 U7887 ( .A1(n6666), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6397) );
  INV_X1 U7888 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9476) );
  OR2_X1 U7889 ( .A1(n6458), .A2(n9476), .ZN(n6396) );
  INV_X1 U7890 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9046) );
  NAND2_X1 U7891 ( .A1(n6392), .A2(n9046), .ZN(n6393) );
  NAND2_X1 U7892 ( .A1(n6414), .A2(n6393), .ZN(n9391) );
  OR2_X1 U7893 ( .A1(n6587), .A2(n9391), .ZN(n6395) );
  INV_X1 U7894 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9392) );
  OR2_X1 U7895 ( .A1(n6501), .A2(n9392), .ZN(n6394) );
  NAND4_X1 U7896 ( .A1(n6397), .A2(n6396), .A3(n6395), .A4(n6394), .ZN(n9366)
         );
  NAND2_X1 U7897 ( .A1(n9366), .A2(n4486), .ZN(n6398) );
  NAND2_X1 U7898 ( .A1(n6399), .A2(n6398), .ZN(n6400) );
  XNOR2_X1 U7899 ( .A(n6400), .B(n6556), .ZN(n6402) );
  AND2_X1 U7900 ( .A1(n9366), .A2(n6628), .ZN(n6401) );
  AOI21_X1 U7901 ( .B1(n9390), .B2(n4482), .A(n6401), .ZN(n6403) );
  NAND2_X1 U7902 ( .A1(n6402), .A2(n6403), .ZN(n6408) );
  INV_X1 U7903 ( .A(n6402), .ZN(n6405) );
  INV_X1 U7904 ( .A(n6403), .ZN(n6404) );
  NAND2_X1 U7905 ( .A1(n6405), .A2(n6404), .ZN(n6406) );
  NAND2_X1 U7906 ( .A1(n6408), .A2(n6406), .ZN(n9044) );
  INV_X1 U7907 ( .A(n9044), .ZN(n6407) );
  NAND2_X1 U7908 ( .A1(n7386), .A2(n6244), .ZN(n6412) );
  INV_X1 U7909 ( .A(n6409), .ZN(n6410) );
  NAND2_X1 U7910 ( .A1(n6410), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6429) );
  XNOR2_X1 U7911 ( .A(n6429), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9781) );
  AOI22_X1 U7912 ( .A1(n6450), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6449), .B2(
        n9781), .ZN(n6411) );
  NAND2_X1 U7913 ( .A1(n9465), .A2(n6521), .ZN(n6421) );
  NAND2_X1 U7914 ( .A1(n6666), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6419) );
  INV_X1 U7915 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9157) );
  OR2_X1 U7916 ( .A1(n6458), .A2(n9157), .ZN(n6418) );
  INV_X1 U7917 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6413) );
  NAND2_X1 U7918 ( .A1(n6414), .A2(n6413), .ZN(n6415) );
  NAND2_X1 U7919 ( .A1(n6436), .A2(n6415), .ZN(n9369) );
  OR2_X1 U7920 ( .A1(n6587), .A2(n9369), .ZN(n6417) );
  INV_X1 U7921 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9361) );
  OR2_X1 U7922 ( .A1(n6501), .A2(n9361), .ZN(n6416) );
  NAND4_X1 U7923 ( .A1(n6419), .A2(n6418), .A3(n6417), .A4(n6416), .ZN(n9380)
         );
  NAND2_X1 U7924 ( .A1(n9380), .A2(n4486), .ZN(n6420) );
  NAND2_X1 U7925 ( .A1(n6421), .A2(n6420), .ZN(n6422) );
  XNOR2_X1 U7926 ( .A(n6422), .B(n7492), .ZN(n6424) );
  AND2_X1 U7927 ( .A1(n9380), .A2(n6628), .ZN(n6423) );
  AOI21_X1 U7928 ( .B1(n9465), .B2(n4484), .A(n6423), .ZN(n6425) );
  XNOR2_X1 U7929 ( .A(n6424), .B(n6425), .ZN(n9053) );
  NAND2_X1 U7930 ( .A1(n9052), .A2(n9053), .ZN(n9051) );
  INV_X1 U7931 ( .A(n6424), .ZN(n6426) );
  NAND2_X1 U7932 ( .A1(n6426), .A2(n6425), .ZN(n6427) );
  NAND2_X1 U7933 ( .A1(n9051), .A2(n6427), .ZN(n6447) );
  NAND2_X1 U7934 ( .A1(n7519), .A2(n6244), .ZN(n6433) );
  NAND2_X1 U7935 ( .A1(n6429), .A2(n6428), .ZN(n6430) );
  NAND2_X1 U7936 ( .A1(n6430), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6431) );
  XNOR2_X1 U7937 ( .A(n6431), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9797) );
  AOI22_X1 U7938 ( .A1(n6450), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6449), .B2(
        n9797), .ZN(n6432) );
  NAND2_X1 U7939 ( .A1(n9462), .A2(n6521), .ZN(n6443) );
  NAND2_X1 U7940 ( .A1(n6666), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6441) );
  INV_X1 U7941 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9159) );
  OR2_X1 U7942 ( .A1(n6458), .A2(n9159), .ZN(n6440) );
  INV_X1 U7943 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6435) );
  NAND2_X1 U7944 ( .A1(n6436), .A2(n6435), .ZN(n6437) );
  NAND2_X1 U7945 ( .A1(n6455), .A2(n6437), .ZN(n9091) );
  OR2_X1 U7946 ( .A1(n6587), .A2(n9091), .ZN(n6439) );
  INV_X1 U7947 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9147) );
  OR2_X1 U7948 ( .A1(n6501), .A2(n9147), .ZN(n6438) );
  NAND4_X1 U7949 ( .A1(n6441), .A2(n6440), .A3(n6439), .A4(n6438), .ZN(n9367)
         );
  NAND2_X1 U7950 ( .A1(n9367), .A2(n4484), .ZN(n6442) );
  NAND2_X1 U7951 ( .A1(n6443), .A2(n6442), .ZN(n6444) );
  XNOR2_X1 U7952 ( .A(n6444), .B(n6556), .ZN(n6448) );
  NAND2_X1 U7953 ( .A1(n9462), .A2(n4481), .ZN(n6446) );
  NAND2_X1 U7954 ( .A1(n9367), .A2(n6486), .ZN(n6445) );
  NAND2_X1 U7955 ( .A1(n6446), .A2(n6445), .ZN(n9090) );
  NAND2_X1 U7956 ( .A1(n7669), .A2(n6244), .ZN(n6452) );
  AOI22_X1 U7957 ( .A1(n6450), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9317), .B2(
        n6449), .ZN(n6451) );
  NAND2_X1 U7958 ( .A1(n9455), .A2(n6521), .ZN(n6464) );
  INV_X1 U7959 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6454) );
  NAND2_X1 U7960 ( .A1(n6455), .A2(n6454), .ZN(n6456) );
  AND2_X1 U7961 ( .A1(n6479), .A2(n6456), .ZN(n9344) );
  NAND2_X1 U7962 ( .A1(n6453), .A2(n9344), .ZN(n6462) );
  NAND2_X1 U7963 ( .A1(n6666), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6461) );
  INV_X1 U7964 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n6457) );
  OR2_X1 U7965 ( .A1(n6501), .A2(n6457), .ZN(n6460) );
  INV_X1 U7966 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9161) );
  OR2_X1 U7967 ( .A1(n6458), .A2(n9161), .ZN(n6459) );
  NAND4_X1 U7968 ( .A1(n6462), .A2(n6461), .A3(n6460), .A4(n6459), .ZN(n9126)
         );
  NAND2_X1 U7969 ( .A1(n9126), .A2(n4482), .ZN(n6463) );
  NAND2_X1 U7970 ( .A1(n6464), .A2(n6463), .ZN(n6465) );
  XNOR2_X1 U7971 ( .A(n6465), .B(n6556), .ZN(n6467) );
  AND2_X1 U7972 ( .A1(n9126), .A2(n6628), .ZN(n6466) );
  AOI21_X1 U7973 ( .B1(n9455), .B2(n4485), .A(n6466), .ZN(n6468) );
  NAND2_X1 U7974 ( .A1(n6467), .A2(n6468), .ZN(n6473) );
  INV_X1 U7975 ( .A(n6467), .ZN(n6470) );
  INV_X1 U7976 ( .A(n6468), .ZN(n6469) );
  NAND2_X1 U7977 ( .A1(n6470), .A2(n6469), .ZN(n6471) );
  NAND2_X1 U7978 ( .A1(n6473), .A2(n6471), .ZN(n9022) );
  INV_X1 U7979 ( .A(n9022), .ZN(n6472) );
  NAND2_X1 U7980 ( .A1(n7739), .A2(n6244), .ZN(n6475) );
  OR2_X1 U7981 ( .A1(n8134), .A2(n10419), .ZN(n6474) );
  NAND2_X1 U7982 ( .A1(n9449), .A2(n6521), .ZN(n6484) );
  INV_X1 U7983 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9453) );
  NAND2_X1 U7984 ( .A1(n6666), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6477) );
  NAND2_X1 U7985 ( .A1(n6667), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6476) );
  AND2_X1 U7986 ( .A1(n6477), .A2(n6476), .ZN(n6482) );
  INV_X1 U7987 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9073) );
  NAND2_X1 U7988 ( .A1(n6479), .A2(n9073), .ZN(n6480) );
  NAND2_X1 U7989 ( .A1(n6495), .A2(n6480), .ZN(n9324) );
  OR2_X1 U7990 ( .A1(n9324), .A2(n6587), .ZN(n6481) );
  OAI211_X1 U7991 ( .C1(n6458), .C2(n9453), .A(n6482), .B(n6481), .ZN(n9353)
         );
  NAND2_X1 U7992 ( .A1(n9353), .A2(n4486), .ZN(n6483) );
  NAND2_X1 U7993 ( .A1(n6484), .A2(n6483), .ZN(n6485) );
  XNOR2_X1 U7994 ( .A(n6485), .B(n7492), .ZN(n6489) );
  NAND2_X1 U7995 ( .A1(n9449), .A2(n4484), .ZN(n6488) );
  NAND2_X1 U7996 ( .A1(n9353), .A2(n6486), .ZN(n6487) );
  NAND2_X1 U7997 ( .A1(n6488), .A2(n6487), .ZN(n6490) );
  NAND2_X1 U7998 ( .A1(n6489), .A2(n6490), .ZN(n9069) );
  INV_X1 U7999 ( .A(n6489), .ZN(n6492) );
  INV_X1 U8000 ( .A(n6490), .ZN(n6491) );
  NAND2_X1 U8001 ( .A1(n6492), .A2(n6491), .ZN(n9071) );
  NAND2_X1 U8002 ( .A1(n7780), .A2(n6244), .ZN(n6494) );
  OR2_X1 U8003 ( .A1(n8134), .A2(n8087), .ZN(n6493) );
  NAND2_X1 U8004 ( .A1(n9443), .A2(n6521), .ZN(n6503) );
  INV_X1 U8005 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n6500) );
  INV_X1 U8006 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9029) );
  NAND2_X1 U8007 ( .A1(n6495), .A2(n9029), .ZN(n6496) );
  NAND2_X1 U8008 ( .A1(n6513), .A2(n6496), .ZN(n9316) );
  OR2_X1 U8009 ( .A1(n9316), .A2(n6587), .ZN(n6499) );
  AOI22_X1 U8010 ( .A1(n6497), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n6666), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n6498) );
  OAI211_X1 U8011 ( .C1(n6501), .C2(n6500), .A(n6499), .B(n6498), .ZN(n9302)
         );
  NAND2_X1 U8012 ( .A1(n9302), .A2(n4486), .ZN(n6502) );
  NAND2_X1 U8013 ( .A1(n6503), .A2(n6502), .ZN(n6504) );
  XNOR2_X1 U8014 ( .A(n6504), .B(n7492), .ZN(n6506) );
  AND2_X1 U8015 ( .A1(n9302), .A2(n6628), .ZN(n6505) );
  AOI21_X1 U8016 ( .B1(n9443), .B2(n4482), .A(n6505), .ZN(n6507) );
  XNOR2_X1 U8017 ( .A(n6506), .B(n6507), .ZN(n9027) );
  INV_X1 U8018 ( .A(n6506), .ZN(n6508) );
  NAND2_X1 U8019 ( .A1(n6508), .A2(n6507), .ZN(n6509) );
  NAND2_X1 U8020 ( .A1(n7913), .A2(n6244), .ZN(n6512) );
  OR2_X1 U8021 ( .A1(n8134), .A2(n7914), .ZN(n6511) );
  INV_X1 U8022 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9082) );
  NAND2_X1 U8023 ( .A1(n6513), .A2(n9082), .ZN(n6514) );
  NAND2_X1 U8024 ( .A1(n6529), .A2(n6514), .ZN(n9296) );
  INV_X1 U8025 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6517) );
  NAND2_X1 U8026 ( .A1(n6667), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6516) );
  NAND2_X1 U8027 ( .A1(n6666), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6515) );
  OAI211_X1 U8028 ( .C1(n6458), .C2(n6517), .A(n6516), .B(n6515), .ZN(n6518)
         );
  INV_X1 U8029 ( .A(n6518), .ZN(n6519) );
  OAI21_X1 U8030 ( .B1(n9296), .B2(n6587), .A(n6519), .ZN(n9279) );
  AND2_X1 U8031 ( .A1(n9279), .A2(n6628), .ZN(n6520) );
  AOI21_X1 U8032 ( .B1(n9438), .B2(n4484), .A(n6520), .ZN(n6525) );
  NAND2_X1 U8033 ( .A1(n9438), .A2(n6521), .ZN(n6523) );
  NAND2_X1 U8034 ( .A1(n9279), .A2(n4481), .ZN(n6522) );
  NAND2_X1 U8035 ( .A1(n6523), .A2(n6522), .ZN(n6524) );
  NAND2_X1 U8036 ( .A1(n7958), .A2(n6244), .ZN(n6527) );
  OR2_X1 U8037 ( .A1(n8134), .A2(n10402), .ZN(n6526) );
  NAND2_X1 U8038 ( .A1(n9286), .A2(n6521), .ZN(n6537) );
  INV_X1 U8039 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9014) );
  NAND2_X1 U8040 ( .A1(n6529), .A2(n9014), .ZN(n6530) );
  NAND2_X1 U8041 ( .A1(n6546), .A2(n6530), .ZN(n9287) );
  INV_X1 U8042 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9436) );
  NAND2_X1 U8043 ( .A1(n6666), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6532) );
  NAND2_X1 U8044 ( .A1(n6667), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6531) );
  OAI211_X1 U8045 ( .C1(n6458), .C2(n9436), .A(n6532), .B(n6531), .ZN(n6533)
         );
  INV_X1 U8046 ( .A(n6533), .ZN(n6534) );
  NAND2_X1 U8047 ( .A1(n9303), .A2(n4485), .ZN(n6536) );
  NAND2_X1 U8048 ( .A1(n6537), .A2(n6536), .ZN(n6538) );
  NAND2_X1 U8049 ( .A1(n9286), .A2(n4486), .ZN(n6540) );
  NAND2_X1 U8050 ( .A1(n9303), .A2(n6628), .ZN(n6539) );
  NAND2_X1 U8051 ( .A1(n6540), .A2(n6539), .ZN(n9013) );
  NAND2_X1 U8052 ( .A1(n9010), .A2(n9013), .ZN(n6541) );
  NAND2_X1 U8053 ( .A1(n4738), .A2(n4576), .ZN(n9011) );
  NAND2_X1 U8054 ( .A1(n6541), .A2(n9011), .ZN(n9058) );
  NAND2_X1 U8055 ( .A1(n7989), .A2(n6244), .ZN(n6543) );
  OR2_X1 U8056 ( .A1(n8134), .A2(n8003), .ZN(n6542) );
  NAND2_X1 U8057 ( .A1(n9428), .A2(n6521), .ZN(n6555) );
  INV_X1 U8058 ( .A(n6546), .ZN(n6544) );
  NAND2_X1 U8059 ( .A1(n6544), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6566) );
  INV_X1 U8060 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6545) );
  NAND2_X1 U8061 ( .A1(n6546), .A2(n6545), .ZN(n6547) );
  NAND2_X1 U8062 ( .A1(n6566), .A2(n6547), .ZN(n9260) );
  OR2_X1 U8063 ( .A1(n9260), .A2(n6587), .ZN(n6553) );
  INV_X1 U8064 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6550) );
  NAND2_X1 U8065 ( .A1(n6666), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6549) );
  NAND2_X1 U8066 ( .A1(n6667), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6548) );
  OAI211_X1 U8067 ( .C1(n6458), .C2(n6550), .A(n6549), .B(n6548), .ZN(n6551)
         );
  INV_X1 U8068 ( .A(n6551), .ZN(n6552) );
  NAND2_X1 U8069 ( .A1(n9280), .A2(n4486), .ZN(n6554) );
  NAND2_X1 U8070 ( .A1(n6555), .A2(n6554), .ZN(n6557) );
  XNOR2_X1 U8071 ( .A(n6557), .B(n6556), .ZN(n6561) );
  AND2_X1 U8072 ( .A1(n9280), .A2(n6628), .ZN(n6558) );
  AOI21_X1 U8073 ( .B1(n9428), .B2(n4482), .A(n6558), .ZN(n6560) );
  XNOR2_X1 U8074 ( .A(n6561), .B(n6560), .ZN(n9061) );
  NAND2_X1 U8075 ( .A1(n6561), .A2(n6560), .ZN(n6562) );
  NAND2_X1 U8076 ( .A1(n8067), .A2(n6244), .ZN(n6564) );
  OR2_X1 U8077 ( .A1(n8134), .A2(n8068), .ZN(n6563) );
  NAND2_X1 U8078 ( .A1(n9423), .A2(n6521), .ZN(n6575) );
  INV_X1 U8079 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6565) );
  NAND2_X1 U8080 ( .A1(n6566), .A2(n6565), .ZN(n6567) );
  NAND2_X1 U8081 ( .A1(n9247), .A2(n6453), .ZN(n6573) );
  INV_X1 U8082 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6570) );
  NAND2_X1 U8083 ( .A1(n6667), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6569) );
  NAND2_X1 U8084 ( .A1(n6666), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6568) );
  OAI211_X1 U8085 ( .C1(n6458), .C2(n6570), .A(n6569), .B(n6568), .ZN(n6571)
         );
  INV_X1 U8086 ( .A(n6571), .ZN(n6572) );
  NAND2_X1 U8087 ( .A1(n9267), .A2(n4481), .ZN(n6574) );
  NAND2_X1 U8088 ( .A1(n6575), .A2(n6574), .ZN(n6576) );
  XNOR2_X1 U8089 ( .A(n6576), .B(n7492), .ZN(n6578) );
  AND2_X1 U8090 ( .A1(n9267), .A2(n6628), .ZN(n6577) );
  AOI21_X1 U8091 ( .B1(n9423), .B2(n4482), .A(n6577), .ZN(n6579) );
  XNOR2_X1 U8092 ( .A(n6578), .B(n6579), .ZN(n9035) );
  INV_X1 U8093 ( .A(n6578), .ZN(n6580) );
  NAND2_X1 U8094 ( .A1(n8979), .A2(n6244), .ZN(n6582) );
  OR2_X1 U8095 ( .A1(n8134), .A2(n9550), .ZN(n6581) );
  NAND2_X1 U8096 ( .A1(n9236), .A2(n6521), .ZN(n6594) );
  INV_X1 U8097 ( .A(n6585), .ZN(n6583) );
  INV_X1 U8098 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6584) );
  NAND2_X1 U8099 ( .A1(n6585), .A2(n6584), .ZN(n6586) );
  NAND2_X1 U8100 ( .A1(n6621), .A2(n6586), .ZN(n9102) );
  INV_X1 U8101 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9421) );
  NAND2_X1 U8102 ( .A1(n6667), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6589) );
  NAND2_X1 U8103 ( .A1(n6666), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6588) );
  OAI211_X1 U8104 ( .C1(n6458), .C2(n9421), .A(n6589), .B(n6588), .ZN(n6590)
         );
  INV_X1 U8105 ( .A(n6590), .ZN(n6591) );
  NAND2_X1 U8106 ( .A1(n9252), .A2(n4482), .ZN(n6593) );
  NAND2_X1 U8107 ( .A1(n6594), .A2(n6593), .ZN(n6595) );
  XNOR2_X1 U8108 ( .A(n6595), .B(n7492), .ZN(n6599) );
  AND2_X1 U8109 ( .A1(n9252), .A2(n6628), .ZN(n6596) );
  AOI21_X1 U8110 ( .B1(n9236), .B2(n4485), .A(n6596), .ZN(n6597) );
  XNOR2_X1 U8111 ( .A(n6599), .B(n6597), .ZN(n9100) );
  NAND2_X1 U8112 ( .A1(n9101), .A2(n9100), .ZN(n9099) );
  INV_X1 U8113 ( .A(n6597), .ZN(n6598) );
  NAND2_X1 U8114 ( .A1(n6599), .A2(n6598), .ZN(n6600) );
  NAND2_X1 U8115 ( .A1(n6601), .A2(n6244), .ZN(n6603) );
  OR2_X1 U8116 ( .A1(n8134), .A2(n9548), .ZN(n6602) );
  NAND2_X1 U8117 ( .A1(n9415), .A2(n6521), .ZN(n6611) );
  XNOR2_X1 U8118 ( .A(n6621), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9223) );
  NAND2_X1 U8119 ( .A1(n9223), .A2(n6453), .ZN(n6609) );
  INV_X1 U8120 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n6606) );
  NAND2_X1 U8121 ( .A1(n6666), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6605) );
  NAND2_X1 U8122 ( .A1(n6667), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6604) );
  OAI211_X1 U8123 ( .C1(n6458), .C2(n6606), .A(n6605), .B(n6604), .ZN(n6607)
         );
  INV_X1 U8124 ( .A(n6607), .ZN(n6608) );
  NAND2_X1 U8125 ( .A1(n9233), .A2(n4485), .ZN(n6610) );
  NAND2_X1 U8126 ( .A1(n6611), .A2(n6610), .ZN(n6612) );
  XNOR2_X1 U8127 ( .A(n6612), .B(n7492), .ZN(n6658) );
  NAND2_X1 U8128 ( .A1(n9415), .A2(n4484), .ZN(n6614) );
  NAND2_X1 U8129 ( .A1(n9233), .A2(n6628), .ZN(n6613) );
  NAND2_X1 U8130 ( .A1(n6614), .A2(n6613), .ZN(n6659) );
  NAND2_X1 U8131 ( .A1(n6615), .A2(n6244), .ZN(n6617) );
  OR2_X1 U8132 ( .A1(n8134), .A2(n8117), .ZN(n6616) );
  NAND2_X1 U8133 ( .A1(n9203), .A2(n4484), .ZN(n6630) );
  INV_X1 U8134 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6619) );
  INV_X1 U8135 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6618) );
  OAI21_X1 U8136 ( .B1(n6621), .B2(n6619), .A(n6618), .ZN(n6622) );
  NAND2_X1 U8137 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .ZN(n6620) );
  NAND2_X1 U8138 ( .A1(n9207), .A2(n6453), .ZN(n6627) );
  INV_X1 U8139 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9411) );
  NAND2_X1 U8140 ( .A1(n6666), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6624) );
  NAND2_X1 U8141 ( .A1(n6667), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6623) );
  OAI211_X1 U8142 ( .C1(n6458), .C2(n9411), .A(n6624), .B(n6623), .ZN(n6625)
         );
  INV_X1 U8143 ( .A(n6625), .ZN(n6626) );
  NAND2_X1 U8144 ( .A1(n9217), .A2(n6628), .ZN(n6629) );
  NAND2_X1 U8145 ( .A1(n6630), .A2(n6629), .ZN(n6631) );
  XNOR2_X1 U8146 ( .A(n6631), .B(n7492), .ZN(n6633) );
  AOI22_X1 U8147 ( .A1(n9203), .A2(n6521), .B1(n4481), .B2(n9217), .ZN(n6632)
         );
  XNOR2_X1 U8148 ( .A(n6633), .B(n6632), .ZN(n6662) );
  INV_X1 U8149 ( .A(n6662), .ZN(n6689) );
  NAND3_X1 U8150 ( .A1(n8069), .A2(P1_B_REG_SCAN_IN), .A3(n8005), .ZN(n6636)
         );
  INV_X1 U8151 ( .A(n8005), .ZN(n6634) );
  INV_X1 U8152 ( .A(P1_B_REG_SCAN_IN), .ZN(n6760) );
  NAND2_X1 U8153 ( .A1(n6634), .A2(n6760), .ZN(n6635) );
  NAND2_X1 U8154 ( .A1(n6636), .A2(n6635), .ZN(n6637) );
  OR2_X1 U8155 ( .A1(n9807), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6639) );
  NAND2_X1 U8156 ( .A1(n9552), .A2(n8005), .ZN(n6638) );
  NAND2_X1 U8157 ( .A1(n6639), .A2(n6638), .ZN(n6857) );
  NOR4_X1 U8158 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6648) );
  NOR4_X1 U8159 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6647) );
  NOR4_X1 U8160 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6643) );
  NOR4_X1 U8161 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6642) );
  NOR4_X1 U8162 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6641) );
  NOR4_X1 U8163 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6640) );
  NAND4_X1 U8164 ( .A1(n6643), .A2(n6642), .A3(n6641), .A4(n6640), .ZN(n6644)
         );
  NOR4_X1 U8165 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n6645), .A4(n6644), .ZN(n6646) );
  AND3_X1 U8166 ( .A1(n6648), .A2(n6647), .A3(n6646), .ZN(n6649) );
  NOR2_X1 U8167 ( .A1(n9807), .A2(n6649), .ZN(n6780) );
  NAND2_X1 U8168 ( .A1(n9552), .A2(n8069), .ZN(n6650) );
  NOR2_X1 U8169 ( .A1(n6776), .A2(n7490), .ZN(n6677) );
  NAND2_X1 U8170 ( .A1(n4591), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6652) );
  MUX2_X1 U8171 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6652), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n6654) );
  NAND2_X1 U8172 ( .A1(n6654), .A2(n6653), .ZN(n6801) );
  AND2_X1 U8173 ( .A1(n6801), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6655) );
  AND2_X1 U8174 ( .A1(n6677), .A2(n9808), .ZN(n6671) );
  NAND2_X1 U8175 ( .A1(n7915), .A2(n6657), .ZN(n9488) );
  AND2_X1 U8176 ( .A1(n9826), .A2(n8425), .ZN(n6680) );
  INV_X1 U8177 ( .A(n6658), .ZN(n6661) );
  INV_X1 U8178 ( .A(n6659), .ZN(n6660) );
  NAND2_X1 U8179 ( .A1(n6661), .A2(n6660), .ZN(n8986) );
  NAND3_X1 U8180 ( .A1(n6689), .A2(n9115), .A3(n8986), .ZN(n6693) );
  OR2_X1 U8181 ( .A1(n9488), .A2(n8339), .ZN(n6682) );
  INV_X1 U8182 ( .A(n6682), .ZN(n7505) );
  NAND3_X1 U8183 ( .A1(n6677), .A2(n9808), .A3(n7505), .ZN(n6664) );
  NAND2_X1 U8184 ( .A1(n9808), .A2(n6657), .ZN(n6663) );
  INV_X1 U8185 ( .A(n6665), .ZN(n9186) );
  INV_X1 U8186 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6779) );
  NAND2_X1 U8187 ( .A1(n6666), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6669) );
  NAND2_X1 U8188 ( .A1(n6667), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6668) );
  OAI211_X1 U8189 ( .C1(n6458), .C2(n6779), .A(n6669), .B(n6668), .ZN(n6670)
         );
  AOI21_X1 U8190 ( .B1(n9186), .B2(n6453), .A(n6670), .ZN(n9125) );
  INV_X1 U8191 ( .A(n6671), .ZN(n6674) );
  NOR2_X1 U8192 ( .A1(n6674), .A2(n8431), .ZN(n6686) );
  INV_X1 U8193 ( .A(n6686), .ZN(n6676) );
  INV_X1 U8194 ( .A(n4487), .ZN(n9687) );
  INV_X1 U8195 ( .A(n6677), .ZN(n7149) );
  OR2_X1 U8196 ( .A1(n8425), .A2(n6678), .ZN(n6775) );
  NAND3_X1 U8197 ( .A1(n6775), .A2(n6800), .A3(n6801), .ZN(n6679) );
  AOI21_X1 U8198 ( .B1(n7149), .B2(n6680), .A(n6679), .ZN(n6681) );
  OR2_X1 U8199 ( .A1(n6681), .A2(n4476), .ZN(n6685) );
  NAND2_X1 U8200 ( .A1(n6682), .A2(n8431), .ZN(n6683) );
  AND2_X1 U8201 ( .A1(n6683), .A2(n9808), .ZN(n7150) );
  NAND2_X1 U8202 ( .A1(n7149), .A2(n7150), .ZN(n6684) );
  NAND2_X1 U8203 ( .A1(n6685), .A2(n6684), .ZN(n9103) );
  AOI22_X1 U8204 ( .A1(n9207), .A2(n9103), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        n4476), .ZN(n6688) );
  NAND2_X1 U8205 ( .A1(n9233), .A2(n9120), .ZN(n6687) );
  OAI211_X1 U8206 ( .C1(n9125), .C2(n9117), .A(n6688), .B(n6687), .ZN(n6691)
         );
  NOR3_X1 U8207 ( .A1(n6689), .A2(n9097), .A3(n8986), .ZN(n6690) );
  AOI211_X1 U8208 ( .C1(n9203), .C2(n9095), .A(n6691), .B(n6690), .ZN(n6692)
         );
  AND2_X1 U8209 ( .A1(n6696), .A2(n7538), .ZN(n7188) );
  NAND2_X1 U8210 ( .A1(n6695), .A2(n6694), .ZN(n6697) );
  NAND2_X1 U8211 ( .A1(n7187), .A2(n6697), .ZN(n7371) );
  INV_X1 U8212 ( .A(n7371), .ZN(n6699) );
  XNOR2_X2 U8213 ( .A(n9138), .B(n7377), .ZN(n8346) );
  INV_X1 U8214 ( .A(n8346), .ZN(n6698) );
  NAND2_X1 U8215 ( .A1(n6699), .A2(n6698), .ZN(n7369) );
  OR2_X1 U8216 ( .A1(n9138), .A2(n4479), .ZN(n6700) );
  NAND2_X1 U8217 ( .A1(n7369), .A2(n6700), .ZN(n7691) );
  NAND2_X1 U8218 ( .A1(n7691), .A2(n8343), .ZN(n7690) );
  OR2_X1 U8219 ( .A1(n6701), .A2(n6702), .ZN(n6703) );
  NAND2_X1 U8220 ( .A1(n7690), .A2(n6703), .ZN(n7359) );
  OR2_X1 U8221 ( .A1(n9137), .A2(n7363), .ZN(n7494) );
  NAND2_X1 U8222 ( .A1(n9137), .A2(n7363), .ZN(n8379) );
  NAND2_X1 U8223 ( .A1(n7494), .A2(n8379), .ZN(n8342) );
  NAND2_X1 U8224 ( .A1(n7359), .A2(n8342), .ZN(n7361) );
  OR2_X1 U8225 ( .A1(n9137), .A2(n7661), .ZN(n6704) );
  NAND2_X1 U8226 ( .A1(n7361), .A2(n6704), .ZN(n7489) );
  INV_X1 U8227 ( .A(n7489), .ZN(n6705) );
  INV_X1 U8228 ( .A(n6768), .ZN(n9818) );
  NAND2_X1 U8229 ( .A1(n9136), .A2(n9818), .ZN(n8148) );
  NAND2_X1 U8230 ( .A1(n8146), .A2(n8148), .ZN(n7497) );
  AOI21_X1 U8231 ( .B1(n6705), .B2(n7497), .A(n5107), .ZN(n7673) );
  NAND2_X1 U8232 ( .A1(n9135), .A2(n7682), .ZN(n8157) );
  NAND2_X1 U8233 ( .A1(n8158), .A2(n8157), .ZN(n8154) );
  NAND2_X1 U8234 ( .A1(n7673), .A2(n8154), .ZN(n7672) );
  OR2_X1 U8235 ( .A1(n9135), .A2(n7784), .ZN(n6706) );
  NAND2_X1 U8236 ( .A1(n7672), .A2(n6706), .ZN(n7559) );
  NAND2_X1 U8237 ( .A1(n9134), .A2(n7622), .ZN(n8380) );
  NAND2_X1 U8238 ( .A1(n8275), .A2(n8380), .ZN(n8155) );
  NAND2_X1 U8239 ( .A1(n7559), .A2(n8155), .ZN(n7558) );
  OR2_X1 U8240 ( .A1(n9134), .A2(n7625), .ZN(n6707) );
  NAND2_X1 U8241 ( .A1(n7558), .A2(n6707), .ZN(n7750) );
  INV_X1 U8242 ( .A(n7750), .ZN(n6709) );
  INV_X1 U8243 ( .A(n7840), .ZN(n7804) );
  NAND2_X1 U8244 ( .A1(n7804), .A2(n9133), .ZN(n8164) );
  INV_X1 U8245 ( .A(n9133), .ZN(n7854) );
  NAND2_X1 U8246 ( .A1(n7854), .A2(n7840), .ZN(n8276) );
  NAND2_X1 U8247 ( .A1(n6709), .A2(n6708), .ZN(n7749) );
  NAND2_X1 U8248 ( .A1(n7840), .A2(n9133), .ZN(n6710) );
  NAND2_X1 U8249 ( .A1(n7749), .A2(n6710), .ZN(n7851) );
  AND2_X1 U8250 ( .A1(n9825), .A2(n9132), .ZN(n6711) );
  NAND2_X1 U8251 ( .A1(n7895), .A2(n9645), .ZN(n8185) );
  NAND2_X1 U8252 ( .A1(n8292), .A2(n8185), .ZN(n7806) );
  INV_X1 U8253 ( .A(n9129), .ZN(n9647) );
  OR2_X1 U8254 ( .A1(n7999), .A2(n9647), .ZN(n8187) );
  NAND2_X1 U8255 ( .A1(n7999), .A2(n9647), .ZN(n8290) );
  NAND2_X1 U8256 ( .A1(n8187), .A2(n8290), .ZN(n8357) );
  NAND2_X1 U8257 ( .A1(n7967), .A2(n8357), .ZN(n6713) );
  NAND2_X1 U8258 ( .A1(n7999), .A2(n9129), .ZN(n6712) );
  NAND2_X1 U8259 ( .A1(n6713), .A2(n6712), .ZN(n7975) );
  INV_X1 U8260 ( .A(n7975), .ZN(n6714) );
  OR2_X1 U8261 ( .A1(n8167), .A2(n9128), .ZN(n6715) );
  NAND2_X1 U8262 ( .A1(n9007), .A2(n9127), .ZN(n6716) );
  INV_X1 U8263 ( .A(n9366), .ZN(n9623) );
  OR2_X1 U8264 ( .A1(n9390), .A2(n9623), .ZN(n8200) );
  NAND2_X1 U8265 ( .A1(n9390), .A2(n9623), .ZN(n8306) );
  NAND2_X1 U8266 ( .A1(n8200), .A2(n8306), .ZN(n9376) );
  INV_X1 U8267 ( .A(n9358), .ZN(n6718) );
  INV_X1 U8268 ( .A(n9367), .ZN(n6719) );
  OR2_X1 U8269 ( .A1(n9462), .A2(n6719), .ZN(n8206) );
  NAND2_X1 U8270 ( .A1(n9462), .A2(n6719), .ZN(n9349) );
  NAND2_X1 U8271 ( .A1(n8206), .A2(n9349), .ZN(n8097) );
  NAND2_X1 U8272 ( .A1(n8091), .A2(n8097), .ZN(n8090) );
  NAND2_X1 U8273 ( .A1(n9462), .A2(n9367), .ZN(n6720) );
  NAND2_X1 U8274 ( .A1(n8090), .A2(n6720), .ZN(n9338) );
  OR2_X1 U8275 ( .A1(n9455), .A2(n9126), .ZN(n6721) );
  NAND2_X1 U8276 ( .A1(n9338), .A2(n6721), .ZN(n6723) );
  NAND2_X1 U8277 ( .A1(n9455), .A2(n9126), .ZN(n6722) );
  NAND2_X1 U8278 ( .A1(n6723), .A2(n6722), .ZN(n9332) );
  OR2_X1 U8279 ( .A1(n9449), .A2(n9353), .ZN(n6724) );
  NAND2_X1 U8280 ( .A1(n9449), .A2(n9353), .ZN(n6725) );
  INV_X1 U8281 ( .A(n9302), .ZN(n9329) );
  OR2_X1 U8282 ( .A1(n9443), .A2(n9329), .ZN(n8313) );
  NAND2_X1 U8283 ( .A1(n9443), .A2(n9329), .ZN(n8220) );
  NAND2_X1 U8284 ( .A1(n8313), .A2(n8220), .ZN(n9309) );
  INV_X1 U8285 ( .A(n9294), .ZN(n6728) );
  AND2_X1 U8286 ( .A1(n9438), .A2(n9279), .ZN(n6726) );
  INV_X1 U8287 ( .A(n6726), .ZN(n6727) );
  OR2_X1 U8288 ( .A1(n9438), .A2(n9279), .ZN(n6729) );
  NOR2_X1 U8289 ( .A1(n9286), .A2(n9303), .ZN(n6731) );
  NAND2_X1 U8290 ( .A1(n9286), .A2(n9303), .ZN(n6730) );
  AND2_X1 U8291 ( .A1(n9428), .A2(n9280), .ZN(n6732) );
  NAND2_X1 U8292 ( .A1(n9423), .A2(n9106), .ZN(n8243) );
  NAND2_X1 U8293 ( .A1(n8269), .A2(n8243), .ZN(n9251) );
  NAND2_X1 U8294 ( .A1(n9243), .A2(n9251), .ZN(n6734) );
  OR2_X1 U8295 ( .A1(n9423), .A2(n9267), .ZN(n6733) );
  NOR2_X1 U8296 ( .A1(n9236), .A2(n9252), .ZN(n6736) );
  NAND2_X1 U8297 ( .A1(n9236), .A2(n9252), .ZN(n6735) );
  INV_X1 U8298 ( .A(n9233), .ZN(n6737) );
  NAND2_X1 U8299 ( .A1(n9415), .A2(n6737), .ZN(n8325) );
  NAND2_X1 U8300 ( .A1(n9203), .A2(n8993), .ZN(n8329) );
  NAND2_X1 U8301 ( .A1(n8082), .A2(n6244), .ZN(n6739) );
  INV_X1 U8302 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8083) );
  OR2_X1 U8303 ( .A1(n8134), .A2(n8083), .ZN(n6738) );
  OR2_X1 U8304 ( .A1(n6774), .A2(n9125), .ZN(n8331) );
  NAND2_X1 U8305 ( .A1(n6774), .A2(n9125), .ZN(n8406) );
  NAND2_X1 U8306 ( .A1(n8331), .A2(n8406), .ZN(n8371) );
  XNOR2_X1 U8307 ( .A(n6740), .B(n8371), .ZN(n9184) );
  NAND3_X1 U8308 ( .A1(n8431), .A2(n7492), .A3(n9331), .ZN(n9652) );
  INV_X1 U8309 ( .A(n7538), .ZN(n9489) );
  NOR2_X1 U8310 ( .A1(n6696), .A2(n9489), .ZN(n7530) );
  NAND2_X1 U8311 ( .A1(n8345), .A2(n7530), .ZN(n6744) );
  OR2_X1 U8312 ( .A1(n9139), .A2(n6742), .ZN(n6743) );
  NAND2_X1 U8313 ( .A1(n6744), .A2(n6743), .ZN(n7372) );
  NAND2_X1 U8314 ( .A1(n7372), .A2(n8346), .ZN(n6746) );
  INV_X1 U8315 ( .A(n4479), .ZN(n8281) );
  OR2_X1 U8316 ( .A1(n9138), .A2(n8281), .ZN(n6745) );
  NAND2_X1 U8317 ( .A1(n6746), .A2(n6745), .ZN(n7689) );
  NAND2_X1 U8318 ( .A1(n6701), .A2(n9811), .ZN(n8284) );
  NAND2_X1 U8319 ( .A1(n7689), .A2(n8284), .ZN(n8391) );
  OR2_X1 U8320 ( .A1(n6701), .A2(n9811), .ZN(n8382) );
  NAND2_X1 U8321 ( .A1(n8391), .A2(n8382), .ZN(n8287) );
  NAND2_X1 U8322 ( .A1(n8146), .A2(n7494), .ZN(n8142) );
  INV_X1 U8323 ( .A(n8158), .ZN(n8387) );
  INV_X1 U8324 ( .A(n8148), .ZN(n8143) );
  NAND2_X1 U8325 ( .A1(n8143), .A2(n8158), .ZN(n6747) );
  AND2_X1 U8326 ( .A1(n6747), .A2(n8157), .ZN(n8381) );
  INV_X1 U8327 ( .A(n8275), .ZN(n6748) );
  NOR2_X1 U8328 ( .A1(n6708), .A2(n6748), .ZN(n6749) );
  NAND2_X1 U8329 ( .A1(n7752), .A2(n6749), .ZN(n7852) );
  INV_X1 U8330 ( .A(n9132), .ZN(n7799) );
  OR2_X1 U8331 ( .A1(n9825), .A2(n7799), .ZN(n8169) );
  AND2_X1 U8332 ( .A1(n8169), .A2(n8164), .ZN(n8181) );
  NAND2_X1 U8333 ( .A1(n9825), .A2(n7799), .ZN(n8178) );
  INV_X1 U8334 ( .A(n9130), .ZN(n7891) );
  NAND2_X1 U8335 ( .A1(n7935), .A2(n7891), .ZN(n8355) );
  NAND2_X1 U8336 ( .A1(n9643), .A2(n8355), .ZN(n7962) );
  OR2_X1 U8337 ( .A1(n7935), .A2(n7891), .ZN(n8356) );
  AND2_X1 U8338 ( .A1(n8187), .A2(n8356), .ZN(n8297) );
  NAND2_X1 U8339 ( .A1(n7962), .A2(n8297), .ZN(n6750) );
  NAND2_X1 U8340 ( .A1(n6750), .A2(n8290), .ZN(n7976) );
  XNOR2_X1 U8341 ( .A(n8167), .B(n9128), .ZN(n8361) );
  INV_X1 U8342 ( .A(n9128), .ZN(n9002) );
  NAND2_X1 U8343 ( .A1(n8167), .A2(n9002), .ZN(n8172) );
  INV_X1 U8344 ( .A(n9127), .ZN(n9624) );
  OR2_X1 U8345 ( .A1(n9007), .A2(n9624), .ZN(n8173) );
  NAND2_X1 U8346 ( .A1(n9007), .A2(n9624), .ZN(n8175) );
  NAND2_X1 U8347 ( .A1(n8173), .A2(n8175), .ZN(n8360) );
  INV_X1 U8348 ( .A(n9381), .ZN(n9003) );
  NAND2_X1 U8349 ( .A1(n6770), .A2(n9003), .ZN(n8302) );
  NAND2_X1 U8350 ( .A1(n9621), .A2(n8302), .ZN(n9375) );
  OR2_X1 U8351 ( .A1(n6770), .A2(n9003), .ZN(n9374) );
  AND2_X1 U8352 ( .A1(n8200), .A2(n9374), .ZN(n8305) );
  NAND2_X1 U8353 ( .A1(n9375), .A2(n8305), .ZN(n6751) );
  INV_X1 U8354 ( .A(n9380), .ZN(n9092) );
  AND2_X1 U8355 ( .A1(n9465), .A2(n9092), .ZN(n8139) );
  OR2_X1 U8356 ( .A1(n9465), .A2(n9092), .ZN(n8198) );
  AND2_X1 U8357 ( .A1(n8206), .A2(n8198), .ZN(n8315) );
  OR2_X1 U8358 ( .A1(n9455), .A2(n9328), .ZN(n8208) );
  NAND2_X1 U8359 ( .A1(n9455), .A2(n9328), .ZN(n8272) );
  NAND2_X1 U8360 ( .A1(n9352), .A2(n8272), .ZN(n9325) );
  INV_X1 U8361 ( .A(n9353), .ZN(n9312) );
  OR2_X1 U8362 ( .A1(n9449), .A2(n9312), .ZN(n8213) );
  NAND2_X1 U8363 ( .A1(n9449), .A2(n9312), .ZN(n8218) );
  NAND2_X1 U8364 ( .A1(n9325), .A2(n9333), .ZN(n6753) );
  INV_X1 U8365 ( .A(n9309), .ZN(n9308) );
  INV_X1 U8366 ( .A(n9279), .ZN(n9313) );
  AND2_X1 U8367 ( .A1(n9438), .A2(n9313), .ZN(n8341) );
  INV_X1 U8368 ( .A(n9303), .ZN(n9083) );
  OR2_X1 U8369 ( .A1(n9286), .A2(n9083), .ZN(n8232) );
  OR2_X1 U8370 ( .A1(n9438), .A2(n9313), .ZN(n9273) );
  AND2_X1 U8371 ( .A1(n8232), .A2(n9273), .ZN(n8317) );
  NAND2_X1 U8372 ( .A1(n9274), .A2(n8317), .ZN(n6754) );
  NAND2_X1 U8373 ( .A1(n9286), .A2(n9083), .ZN(n8228) );
  NAND2_X1 U8374 ( .A1(n6754), .A2(n8228), .ZN(n9266) );
  XNOR2_X1 U8375 ( .A(n9428), .B(n9280), .ZN(n9265) );
  INV_X1 U8376 ( .A(n9280), .ZN(n9038) );
  NAND2_X1 U8377 ( .A1(n9428), .A2(n9038), .ZN(n8234) );
  INV_X1 U8378 ( .A(n8243), .ZN(n6755) );
  INV_X1 U8379 ( .A(n9252), .ZN(n8245) );
  OR2_X1 U8380 ( .A1(n9236), .A2(n8245), .ZN(n8270) );
  NAND2_X1 U8381 ( .A1(n9236), .A2(n8245), .ZN(n8324) );
  NAND2_X1 U8382 ( .A1(n9231), .A2(n9229), .ZN(n6756) );
  NAND2_X1 U8383 ( .A1(n6756), .A2(n8270), .ZN(n9216) );
  NAND2_X1 U8384 ( .A1(n9216), .A2(n9215), .ZN(n9214) );
  NAND2_X1 U8385 ( .A1(n9214), .A2(n8326), .ZN(n9199) );
  NAND2_X1 U8386 ( .A1(n9199), .A2(n9198), .ZN(n9197) );
  NAND2_X1 U8387 ( .A1(n9197), .A2(n8330), .ZN(n6757) );
  XNOR2_X1 U8388 ( .A(n6757), .B(n8371), .ZN(n6759) );
  OR2_X1 U8389 ( .A1(n7915), .A2(n9331), .ZN(n6758) );
  OR2_X1 U8390 ( .A1(n8339), .A2(n6657), .ZN(n8132) );
  NAND2_X1 U8391 ( .A1(n6759), .A2(n9649), .ZN(n6767) );
  NOR2_X1 U8392 ( .A1(n8430), .A2(n6760), .ZN(n6761) );
  NOR2_X1 U8393 ( .A1(n9646), .A2(n6761), .ZN(n9174) );
  INV_X1 U8394 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9405) );
  NOR2_X1 U8395 ( .A1(n6458), .A2(n9405), .ZN(n6765) );
  INV_X1 U8396 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n6762) );
  NOR2_X1 U8397 ( .A1(n6501), .A2(n6762), .ZN(n6764) );
  INV_X1 U8398 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9494) );
  NOR2_X1 U8399 ( .A1(n6145), .A2(n9494), .ZN(n6763) );
  AOI22_X1 U8400 ( .A1(n9217), .A2(n9382), .B1(n9174), .B2(n9124), .ZN(n6766)
         );
  NAND2_X1 U8401 ( .A1(n6767), .A2(n6766), .ZN(n9191) );
  INV_X1 U8402 ( .A(n9423), .ZN(n9249) );
  OR2_X1 U8403 ( .A1(n6694), .A2(n7538), .ZN(n7376) );
  NAND2_X1 U8404 ( .A1(n7695), .A2(n9811), .ZN(n7697) );
  OR2_X1 U8405 ( .A1(n7697), .A2(n7661), .ZN(n7500) );
  NOR2_X1 U8406 ( .A1(n7500), .A2(n6768), .ZN(n7501) );
  NOR2_X1 U8407 ( .A1(n7861), .A2(n7895), .ZN(n9636) );
  NAND2_X1 U8408 ( .A1(n9636), .A2(n9673), .ZN(n9638) );
  INV_X1 U8409 ( .A(n9462), .ZN(n8093) );
  INV_X1 U8410 ( .A(n9455), .ZN(n9346) );
  NAND2_X1 U8411 ( .A1(n9295), .A2(n9509), .ZN(n9283) );
  INV_X1 U8412 ( .A(n9206), .ZN(n6773) );
  AOI211_X1 U8413 ( .C1(n6774), .C2(n6773), .A(n9827), .B(n9179), .ZN(n9185)
         );
  NOR2_X1 U8414 ( .A1(n7151), .A2(n6776), .ZN(n6778) );
  OR2_X1 U8415 ( .A1(n7845), .A2(n6656), .ZN(n6777) );
  INV_X1 U8416 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6784) );
  INV_X1 U8417 ( .A(n6780), .ZN(n6781) );
  NAND2_X1 U8418 ( .A1(n6781), .A2(n6857), .ZN(n6782) );
  NAND2_X1 U8419 ( .A1(n9835), .A2(n9466), .ZN(n9532) );
  NAND2_X1 U8420 ( .A1(n6785), .A2(n5096), .ZN(P1_U3520) );
  INV_X1 U8421 ( .A(n6801), .ZN(n7956) );
  AOI211_X1 U8422 ( .C1(n6789), .C2(n6788), .A(n8542), .B(n6787), .ZN(n6793)
         );
  NOR2_X1 U8423 ( .A1(n4786), .A2(n5785), .ZN(n6792) );
  OAI22_X1 U8424 ( .A1(n9616), .A2(n7878), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5497), .ZN(n6791) );
  OAI22_X1 U8425 ( .A1(n8527), .A2(n7950), .B1(n7773), .B2(n8526), .ZN(n6790)
         );
  OR4_X1 U8426 ( .A1(n6793), .A2(n6792), .A3(n6791), .A4(n6790), .ZN(P2_U3236)
         );
  AOI211_X1 U8427 ( .C1(n6795), .C2(n6794), .A(n8542), .B(n5634), .ZN(n6799)
         );
  INV_X1 U8428 ( .A(n8900), .ZN(n8780) );
  NOR2_X1 U8429 ( .A1(n8780), .A2(n5785), .ZN(n6798) );
  OAI22_X1 U8430 ( .A1(n9616), .A2(n8777), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10347), .ZN(n6797) );
  OAI22_X1 U8431 ( .A1(n8527), .A2(n8784), .B1(n8821), .B2(n8526), .ZN(n6796)
         );
  OR4_X1 U8432 ( .A1(n6799), .A2(n6798), .A3(n6797), .A4(n6796), .ZN(P2_U3235)
         );
  NAND2_X1 U8433 ( .A1(n8425), .A2(n6800), .ZN(n6802) );
  NAND2_X1 U8434 ( .A1(n6802), .A2(n6801), .ZN(n9149) );
  NAND2_X1 U8435 ( .A1(n9149), .A2(n8130), .ZN(n9684) );
  NAND2_X1 U8436 ( .A1(n9684), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NAND2_X1 U8437 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6815) );
  OAI21_X1 U8438 ( .B1(n6805), .B2(n6804), .A(n6803), .ZN(n7148) );
  MUX2_X1 U8439 ( .A(n6815), .B(n7148), .S(n8430), .Z(n6807) );
  INV_X1 U8440 ( .A(n8430), .ZN(n9685) );
  OR2_X1 U8441 ( .A1(n4487), .A2(P1_U3084), .ZN(n8115) );
  AOI21_X1 U8442 ( .B1(n9685), .B2(n6084), .A(n8115), .ZN(n6806) );
  NOR2_X1 U8443 ( .A1(P1_U3084), .A2(n10433), .ZN(n6831) );
  OR2_X1 U8444 ( .A1(n6806), .A2(n6831), .ZN(n9690) );
  OAI211_X1 U8445 ( .C1(n6807), .C2(n4487), .A(n6808), .B(n9690), .ZN(n8113)
         );
  INV_X1 U8446 ( .A(n8113), .ZN(n6829) );
  INV_X1 U8447 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6809) );
  NOR2_X1 U8448 ( .A1(n9806), .A2(n6809), .ZN(n6828) );
  INV_X1 U8449 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6813) );
  OR2_X1 U8450 ( .A1(n8430), .A2(n4476), .ZN(n9546) );
  INV_X1 U8451 ( .A(n9546), .ZN(n9150) );
  AND2_X1 U8452 ( .A1(n9150), .A2(n4487), .ZN(n6810) );
  INV_X1 U8453 ( .A(n6962), .ZN(n6811) );
  NAND2_X1 U8454 ( .A1(n9796), .A2(n6811), .ZN(n6812) );
  OAI21_X1 U8455 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6813), .A(n6812), .ZN(n6827) );
  NOR2_X1 U8456 ( .A1(n8115), .A2(n8430), .ZN(n6814) );
  NAND2_X1 U8457 ( .A1(n9149), .A2(n6814), .ZN(n9790) );
  XNOR2_X1 U8458 ( .A(n6962), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n6818) );
  XNOR2_X1 U8459 ( .A(n6830), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n7035) );
  INV_X1 U8460 ( .A(n6815), .ZN(n7034) );
  NAND2_X1 U8461 ( .A1(n7035), .A2(n7034), .ZN(n7033) );
  INV_X1 U8462 ( .A(n6830), .ZN(n7032) );
  NAND2_X1 U8463 ( .A1(n7032), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6816) );
  NAND2_X1 U8464 ( .A1(n7033), .A2(n6816), .ZN(n6817) );
  NAND2_X1 U8465 ( .A1(n6818), .A2(n6817), .ZN(n6958) );
  OAI21_X1 U8466 ( .B1(n6818), .B2(n6817), .A(n6958), .ZN(n6825) );
  MUX2_X1 U8467 ( .A(n6961), .B(P1_REG1_REG_2__SCAN_IN), .S(n6962), .Z(n6823)
         );
  XNOR2_X1 U8468 ( .A(n6830), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n7031) );
  AND2_X1 U8469 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n7030) );
  NAND2_X1 U8470 ( .A1(n7031), .A2(n7030), .ZN(n6820) );
  NAND2_X1 U8471 ( .A1(n7032), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6819) );
  NAND2_X1 U8472 ( .A1(n6820), .A2(n6819), .ZN(n6822) );
  NOR2_X1 U8473 ( .A1(n8115), .A2(n9685), .ZN(n6821) );
  NAND2_X1 U8474 ( .A1(n6823), .A2(n6822), .ZN(n6967) );
  OAI211_X1 U8475 ( .C1(n6823), .C2(n6822), .A(n9783), .B(n6967), .ZN(n6824)
         );
  OAI21_X1 U8476 ( .B1(n9790), .B2(n6825), .A(n6824), .ZN(n6826) );
  OR4_X1 U8477 ( .A1(n6829), .A2(n6828), .A3(n6827), .A4(n6826), .ZN(P1_U3243)
         );
  NAND2_X1 U8478 ( .A1(n6835), .A2(P1_U3084), .ZN(n9544) );
  AND2_X1 U8479 ( .A1(n8129), .A2(n4476), .ZN(n9545) );
  INV_X2 U8480 ( .A(n9545), .ZN(n8089) );
  OAI222_X1 U8481 ( .A1(n9544), .A2(n6065), .B1(n8089), .B2(n6837), .C1(n6830), 
        .C2(n4476), .ZN(P1_U3352) );
  AOI21_X1 U8482 ( .B1(n6832), .B2(n4476), .A(n6831), .ZN(n6833) );
  INV_X1 U8483 ( .A(n6833), .ZN(P1_U3353) );
  OAI222_X1 U8484 ( .A1(n9544), .A2(n6834), .B1(n8089), .B2(n6848), .C1(n6962), 
        .C2(P1_U3084), .ZN(P1_U3351) );
  NOR2_X1 U8485 ( .A1(n6835), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8965) );
  INV_X2 U8486 ( .A(n8965), .ZN(n8980) );
  NAND2_X1 U8487 ( .A1(n6835), .A2(P2_U3152), .ZN(n8968) );
  OAI222_X1 U8488 ( .A1(n8980), .A2(n6838), .B1(n8968), .B2(n6837), .C1(
        P2_U3152), .C2(n6836), .ZN(P2_U3357) );
  OAI222_X1 U8489 ( .A1(n9544), .A2(n6839), .B1(n8089), .B2(n6845), .C1(n7017), 
        .C2(n4476), .ZN(P1_U3350) );
  OAI222_X1 U8490 ( .A1(n9544), .A2(n6840), .B1(n8089), .B2(n6842), .C1(n7019), 
        .C2(P1_U3084), .ZN(P1_U3349) );
  INV_X1 U8491 ( .A(n8972), .ZN(n8983) );
  AOI22_X1 U8492 ( .A1(n9555), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n8965), .ZN(n6841) );
  OAI21_X1 U8493 ( .B1(n6851), .B2(n8983), .A(n6841), .ZN(P2_U3353) );
  INV_X1 U8494 ( .A(n9861), .ZN(n6935) );
  OAI222_X1 U8495 ( .A1(n8980), .A2(n6843), .B1(n8983), .B2(n6842), .C1(
        P2_U3152), .C2(n6935), .ZN(P2_U3354) );
  OAI222_X1 U8496 ( .A1(n8980), .A2(n6846), .B1(n8983), .B2(n6845), .C1(
        P2_U3152), .C2(n6844), .ZN(P2_U3355) );
  OAI222_X1 U8497 ( .A1(n8980), .A2(n6849), .B1(n8983), .B2(n6848), .C1(
        P2_U3152), .C2(n6847), .ZN(P2_U3356) );
  OAI222_X1 U8498 ( .A1(n9696), .A2(P1_U3084), .B1(n8089), .B2(n6851), .C1(
        n6850), .C2(n9544), .ZN(P1_U3348) );
  AOI22_X1 U8499 ( .A1(n9874), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n8965), .ZN(n6852) );
  OAI21_X1 U8500 ( .B1(n6853), .B2(n8968), .A(n6852), .ZN(P2_U3352) );
  OAI222_X1 U8501 ( .A1(n7075), .A2(n4476), .B1(n8089), .B2(n6853), .C1(n10101), .C2(n9544), .ZN(P1_U3347) );
  INV_X1 U8502 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10416) );
  INV_X1 U8503 ( .A(n6854), .ZN(n8600) );
  NAND2_X1 U8504 ( .A1(n8600), .A2(P2_U3966), .ZN(n6855) );
  OAI21_X1 U8505 ( .B1(P2_U3966), .B2(n10416), .A(n6855), .ZN(P2_U3583) );
  INV_X1 U8506 ( .A(n9808), .ZN(n8432) );
  NAND2_X1 U8507 ( .A1(n8432), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6856) );
  OAI21_X1 U8508 ( .B1(n8432), .B2(n6857), .A(n6856), .ZN(P1_U3440) );
  NOR2_X1 U8509 ( .A1(n7959), .A2(n6945), .ZN(n6858) );
  OR2_X1 U8510 ( .A1(n9938), .A2(n6858), .ZN(n6860) );
  NAND2_X1 U8511 ( .A1(n6915), .A2(n6945), .ZN(n6859) );
  NAND2_X1 U8512 ( .A1(n6860), .A2(n6859), .ZN(n9566) );
  INV_X1 U8513 ( .A(n9566), .ZN(n9899) );
  NOR2_X1 U8514 ( .A1(n9899), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8515 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6862) );
  INV_X1 U8516 ( .A(n6861), .ZN(n6863) );
  INV_X1 U8517 ( .A(n7098), .ZN(n6939) );
  OAI222_X1 U8518 ( .A1(n8980), .A2(n6862), .B1(n8983), .B2(n6863), .C1(
        P2_U3152), .C2(n6939), .ZN(P2_U3351) );
  OAI222_X1 U8519 ( .A1(n7010), .A2(P1_U3084), .B1(n8089), .B2(n6863), .C1(
        n10232), .C2(n9544), .ZN(P1_U3346) );
  NAND2_X1 U8520 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n8560), .ZN(n6864) );
  OAI21_X1 U8521 ( .B1(n8821), .B2(n8560), .A(n6864), .ZN(P2_U3571) );
  INV_X1 U8522 ( .A(n7051), .ZN(n9712) );
  INV_X1 U8523 ( .A(n6865), .ZN(n6867) );
  OAI222_X1 U8524 ( .A1(n9712), .A2(n4476), .B1(n8089), .B2(n6867), .C1(n6866), 
        .C2(n9544), .ZN(P1_U3345) );
  INV_X1 U8525 ( .A(n9886), .ZN(n6910) );
  OAI222_X1 U8526 ( .A1(n8980), .A2(n6868), .B1(n8983), .B2(n6867), .C1(
        P2_U3152), .C2(n6910), .ZN(P2_U3350) );
  INV_X1 U8527 ( .A(n6869), .ZN(n6872) );
  INV_X1 U8528 ( .A(n6985), .ZN(n6942) );
  OAI222_X1 U8529 ( .A1(n8983), .A2(n6872), .B1(n6942), .B2(P2_U3152), .C1(
        n6870), .C2(n8980), .ZN(P2_U3349) );
  INV_X1 U8530 ( .A(n7053), .ZN(n7084) );
  INV_X1 U8531 ( .A(n9539), .ZN(n9549) );
  OAI222_X1 U8532 ( .A1(P1_U3084), .A2(n7084), .B1(n8089), .B2(n6872), .C1(
        n6871), .C2(n9549), .ZN(P1_U3344) );
  INV_X1 U8533 ( .A(n6873), .ZN(n6955) );
  INV_X1 U8534 ( .A(n7000), .ZN(n6943) );
  OAI222_X1 U8535 ( .A1(n8983), .A2(n6955), .B1(n6943), .B2(P2_U3152), .C1(
        n6874), .C2(n8980), .ZN(P2_U3348) );
  NAND3_X1 U8536 ( .A1(n6876), .A2(n7266), .A3(n7268), .ZN(n6878) );
  INV_X1 U8537 ( .A(n7062), .ZN(n7267) );
  XNOR2_X1 U8538 ( .A(n5778), .B(n7270), .ZN(n6879) );
  NAND2_X1 U8539 ( .A1(n6879), .A2(n8835), .ZN(n7877) );
  INV_X1 U8540 ( .A(n10002), .ZN(n8939) );
  NAND2_X1 U8541 ( .A1(n6880), .A2(n6881), .ZN(n7158) );
  OAI21_X1 U8542 ( .B1(n6880), .B2(n6881), .A(n7158), .ZN(n7353) );
  NAND2_X1 U8543 ( .A1(n7141), .A2(n7203), .ZN(n7339) );
  OAI21_X1 U8544 ( .B1(n7141), .B2(n7203), .A(n7339), .ZN(n7349) );
  OAI22_X1 U8545 ( .A1(n7349), .A2(n10013), .B1(n7141), .B2(n10011), .ZN(n6889) );
  XNOR2_X1 U8546 ( .A(n6880), .B(n6883), .ZN(n6886) );
  NAND2_X1 U8547 ( .A1(n6886), .A2(n8795), .ZN(n6888) );
  INV_X1 U8548 ( .A(n8820), .ZN(n8751) );
  AOI22_X1 U8549 ( .A1(n8750), .A2(n8561), .B1(n5806), .B2(n8751), .ZN(n6887)
         );
  NAND2_X1 U8550 ( .A1(n6888), .A2(n6887), .ZN(n7348) );
  AOI211_X1 U8551 ( .C1(n10018), .C2(n7353), .A(n6889), .B(n7348), .ZN(n7065)
         );
  INV_X1 U8552 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6890) );
  OR2_X1 U8553 ( .A1(n10021), .A2(n6890), .ZN(n6891) );
  OAI21_X1 U8554 ( .B1(n10019), .B2(n7065), .A(n6891), .ZN(P2_U3454) );
  INV_X1 U8555 ( .A(n7106), .ZN(n7113) );
  AOI22_X1 U8556 ( .A1(n7106), .A2(n7654), .B1(P2_REG2_REG_11__SCAN_IN), .B2(
        n7113), .ZN(n6914) );
  NAND2_X1 U8557 ( .A1(n7000), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6912) );
  MUX2_X1 U8558 ( .A(n7611), .B(P2_REG2_REG_10__SCAN_IN), .S(n7000), .Z(n6892)
         );
  INV_X1 U8559 ( .A(n6892), .ZN(n6992) );
  NAND2_X1 U8560 ( .A1(n6985), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6911) );
  MUX2_X1 U8561 ( .A(n7552), .B(P2_REG2_REG_9__SCAN_IN), .S(n6985), .Z(n6893)
         );
  INV_X1 U8562 ( .A(n6893), .ZN(n6987) );
  INV_X1 U8563 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6909) );
  MUX2_X1 U8564 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n6909), .S(n9886), .Z(n9891)
         );
  NAND2_X1 U8565 ( .A1(n9874), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6906) );
  MUX2_X1 U8566 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6894), .S(n9874), .Z(n9876)
         );
  NAND2_X1 U8567 ( .A1(n9555), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6905) );
  NAND2_X1 U8568 ( .A1(n9849), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6901) );
  INV_X1 U8569 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6895) );
  MUX2_X1 U8570 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6895), .S(n9849), .Z(n9854)
         );
  NAND2_X1 U8571 ( .A1(n9578), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6900) );
  INV_X1 U8572 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6896) );
  MUX2_X1 U8573 ( .A(n6896), .B(P2_REG2_REG_2__SCAN_IN), .S(n9578), .Z(n6897)
         );
  INV_X1 U8574 ( .A(n6897), .ZN(n9580) );
  NAND2_X1 U8575 ( .A1(n9568), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6899) );
  INV_X1 U8576 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6898) );
  MUX2_X1 U8577 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6898), .S(n9568), .Z(n9570)
         );
  NAND3_X1 U8578 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .A3(n9570), .ZN(n9569) );
  NAND2_X1 U8579 ( .A1(n6899), .A2(n9569), .ZN(n9581) );
  NAND2_X1 U8580 ( .A1(n9580), .A2(n9581), .ZN(n9579) );
  NAND2_X1 U8581 ( .A1(n6900), .A2(n9579), .ZN(n9855) );
  NAND2_X1 U8582 ( .A1(n9854), .A2(n9855), .ZN(n9853) );
  NAND2_X1 U8583 ( .A1(n6901), .A2(n9853), .ZN(n9864) );
  MUX2_X1 U8584 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6902), .S(n9861), .Z(n9863)
         );
  NAND2_X1 U8585 ( .A1(n9864), .A2(n9863), .ZN(n9862) );
  OAI21_X1 U8586 ( .B1(n6902), .B2(n6935), .A(n9862), .ZN(n9561) );
  INV_X1 U8587 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6903) );
  MUX2_X1 U8588 ( .A(n6903), .B(P2_REG2_REG_5__SCAN_IN), .S(n9555), .Z(n6904)
         );
  INV_X1 U8589 ( .A(n6904), .ZN(n9560) );
  NAND2_X1 U8590 ( .A1(n9561), .A2(n9560), .ZN(n9559) );
  NAND2_X1 U8591 ( .A1(n6905), .A2(n9559), .ZN(n9877) );
  NAND2_X1 U8592 ( .A1(n9876), .A2(n9877), .ZN(n9875) );
  AND2_X1 U8593 ( .A1(n6906), .A2(n9875), .ZN(n7094) );
  MUX2_X1 U8594 ( .A(n6908), .B(P2_REG2_REG_7__SCAN_IN), .S(n7098), .Z(n7093)
         );
  NOR2_X1 U8595 ( .A1(n7094), .A2(n7093), .ZN(n7092) );
  INV_X1 U8596 ( .A(n7092), .ZN(n6907) );
  OAI21_X1 U8597 ( .B1(n6908), .B2(n6939), .A(n6907), .ZN(n9892) );
  NAND2_X1 U8598 ( .A1(n9891), .A2(n9892), .ZN(n9890) );
  OAI21_X1 U8599 ( .B1(n6910), .B2(n6909), .A(n9890), .ZN(n6988) );
  NAND2_X1 U8600 ( .A1(n6987), .A2(n6988), .ZN(n6986) );
  NAND2_X1 U8601 ( .A1(n6911), .A2(n6986), .ZN(n6993) );
  NAND2_X1 U8602 ( .A1(n6992), .A2(n6993), .ZN(n6991) );
  NAND2_X1 U8603 ( .A1(n6912), .A2(n6991), .ZN(n6913) );
  NOR2_X1 U8604 ( .A1(n6913), .A2(n6914), .ZN(n7107) );
  AOI21_X1 U8605 ( .B1(n6914), .B2(n6913), .A(n7107), .ZN(n6954) );
  NAND2_X1 U8606 ( .A1(n9938), .A2(n6915), .ZN(n6919) );
  OR2_X1 U8607 ( .A1(n5793), .A2(P2_U3152), .ZN(n8973) );
  OAI21_X1 U8608 ( .B1(n6916), .B2(n8973), .A(n7959), .ZN(n6917) );
  INV_X1 U8609 ( .A(n6917), .ZN(n6918) );
  NAND2_X1 U8610 ( .A1(n6919), .A2(n6918), .ZN(n6947) );
  NAND2_X1 U8611 ( .A1(n6947), .A2(n6945), .ZN(n6920) );
  NAND2_X1 U8612 ( .A1(n6920), .A2(n8560), .ZN(n6922) );
  NOR2_X1 U8613 ( .A1(n5793), .A2(n8977), .ZN(n6921) );
  NAND2_X1 U8614 ( .A1(n6922), .A2(n5793), .ZN(n9842) );
  INV_X1 U8615 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10356) );
  NOR2_X1 U8616 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10356), .ZN(n6923) );
  AOI21_X1 U8617 ( .B1(n9899), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n6923), .ZN(
        n6951) );
  MUX2_X1 U8618 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n6924), .S(n7000), .Z(n6995)
         );
  MUX2_X1 U8619 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n6925), .S(n6985), .Z(n6981)
         );
  NAND2_X1 U8620 ( .A1(n9886), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6941) );
  MUX2_X1 U8621 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6926), .S(n9886), .Z(n9888)
         );
  NAND2_X1 U8622 ( .A1(n9874), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6938) );
  MUX2_X1 U8623 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6927), .S(n9874), .Z(n9879)
         );
  NAND2_X1 U8624 ( .A1(n9555), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6937) );
  NAND2_X1 U8625 ( .A1(n9849), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6933) );
  INV_X1 U8626 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6928) );
  MUX2_X1 U8627 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6928), .S(n9849), .Z(n9851)
         );
  NAND2_X1 U8628 ( .A1(n9578), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6932) );
  INV_X1 U8629 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6929) );
  MUX2_X1 U8630 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6929), .S(n9578), .Z(n9583)
         );
  NAND2_X1 U8631 ( .A1(n9568), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6931) );
  INV_X1 U8632 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6930) );
  MUX2_X1 U8633 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6930), .S(n9568), .Z(n9573)
         );
  NAND3_X1 U8634 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n9573), .ZN(n9572) );
  NAND2_X1 U8635 ( .A1(n6931), .A2(n9572), .ZN(n9584) );
  NAND2_X1 U8636 ( .A1(n9583), .A2(n9584), .ZN(n9582) );
  NAND2_X1 U8637 ( .A1(n6932), .A2(n9582), .ZN(n9852) );
  NAND2_X1 U8638 ( .A1(n9851), .A2(n9852), .ZN(n9850) );
  NAND2_X1 U8639 ( .A1(n6933), .A2(n9850), .ZN(n9867) );
  MUX2_X1 U8640 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6934), .S(n9861), .Z(n9866)
         );
  NAND2_X1 U8641 ( .A1(n9867), .A2(n9866), .ZN(n9865) );
  OAI21_X1 U8642 ( .B1(n6934), .B2(n6935), .A(n9865), .ZN(n9558) );
  INV_X1 U8643 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6936) );
  MUX2_X1 U8644 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6936), .S(n9555), .Z(n9557)
         );
  NAND2_X1 U8645 ( .A1(n9558), .A2(n9557), .ZN(n9556) );
  NAND2_X1 U8646 ( .A1(n6937), .A2(n9556), .ZN(n9880) );
  NAND2_X1 U8647 ( .A1(n9879), .A2(n9880), .ZN(n9878) );
  NAND2_X1 U8648 ( .A1(n6938), .A2(n9878), .ZN(n7097) );
  MUX2_X1 U8649 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6940), .S(n7098), .Z(n7096)
         );
  NAND2_X1 U8650 ( .A1(n7097), .A2(n7096), .ZN(n7095) );
  OAI21_X1 U8651 ( .B1(n6940), .B2(n6939), .A(n7095), .ZN(n9889) );
  NAND2_X1 U8652 ( .A1(n9888), .A2(n9889), .ZN(n9887) );
  NAND2_X1 U8653 ( .A1(n6941), .A2(n9887), .ZN(n6980) );
  NAND2_X1 U8654 ( .A1(n6981), .A2(n6980), .ZN(n6979) );
  OAI21_X1 U8655 ( .B1(n6942), .B2(n6925), .A(n6979), .ZN(n6996) );
  NAND2_X1 U8656 ( .A1(n6995), .A2(n6996), .ZN(n6994) );
  OAI21_X1 U8657 ( .B1(n6943), .B2(n6924), .A(n6994), .ZN(n6949) );
  MUX2_X1 U8658 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n6944), .S(n7106), .Z(n6948)
         );
  AND2_X1 U8659 ( .A1(n6945), .A2(n8977), .ZN(n6946) );
  NAND2_X1 U8660 ( .A1(n6947), .A2(n6946), .ZN(n9843) );
  INV_X1 U8661 ( .A(n9843), .ZN(n9906) );
  NAND2_X1 U8662 ( .A1(n6948), .A2(n6949), .ZN(n7112) );
  OAI211_X1 U8663 ( .C1(n6949), .C2(n6948), .A(n9906), .B(n7112), .ZN(n6950)
         );
  OAI211_X1 U8664 ( .C1(n9842), .C2(n7113), .A(n6951), .B(n6950), .ZN(n6952)
         );
  INV_X1 U8665 ( .A(n6952), .ZN(n6953) );
  OAI21_X1 U8666 ( .B1(n6954), .B2(n9841), .A(n6953), .ZN(P2_U3256) );
  INV_X1 U8667 ( .A(n7055), .ZN(n7128) );
  OAI222_X1 U8668 ( .A1(n4476), .A2(n7128), .B1(n8089), .B2(n6955), .C1(n10230), .C2(n9549), .ZN(P1_U3343) );
  INV_X1 U8669 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6974) );
  INV_X1 U8670 ( .A(n7017), .ZN(n6972) );
  AND2_X1 U8671 ( .A1(n4476), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7249) );
  XNOR2_X1 U8672 ( .A(n7017), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n6960) );
  OR2_X1 U8673 ( .A1(n6962), .A2(n6956), .ZN(n6957) );
  NAND2_X1 U8674 ( .A1(n6958), .A2(n6957), .ZN(n6959) );
  NAND2_X1 U8675 ( .A1(n6959), .A2(n6960), .ZN(n7016) );
  OAI21_X1 U8676 ( .B1(n6960), .B2(n6959), .A(n7016), .ZN(n6970) );
  OR2_X1 U8677 ( .A1(n6962), .A2(n6961), .ZN(n6966) );
  NAND2_X1 U8678 ( .A1(n6967), .A2(n6966), .ZN(n6964) );
  MUX2_X1 U8679 ( .A(n7003), .B(P1_REG1_REG_3__SCAN_IN), .S(n7017), .Z(n6963)
         );
  NAND2_X1 U8680 ( .A1(n6964), .A2(n6963), .ZN(n7005) );
  MUX2_X1 U8681 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n7003), .S(n7017), .Z(n6965)
         );
  NAND3_X1 U8682 ( .A1(n6967), .A2(n6966), .A3(n6965), .ZN(n6968) );
  NAND3_X1 U8683 ( .A1(n9783), .A2(n7005), .A3(n6968), .ZN(n6969) );
  OAI21_X1 U8684 ( .B1(n9790), .B2(n6970), .A(n6969), .ZN(n6971) );
  AOI211_X1 U8685 ( .C1(n6972), .C2(n9796), .A(n7249), .B(n6971), .ZN(n6973)
         );
  OAI21_X1 U8686 ( .B1(n9806), .B2(n6974), .A(n6973), .ZN(P1_U3244) );
  INV_X1 U8687 ( .A(n6975), .ZN(n6978) );
  INV_X1 U8688 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6976) );
  OAI222_X1 U8689 ( .A1(n8983), .A2(n6978), .B1(n7113), .B2(P2_U3152), .C1(
        n6976), .C2(n8980), .ZN(P2_U3347) );
  INV_X1 U8690 ( .A(n7714), .ZN(n7046) );
  INV_X1 U8691 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6977) );
  OAI222_X1 U8692 ( .A1(n4476), .A2(n7046), .B1(n8089), .B2(n6978), .C1(n6977), 
        .C2(n9549), .ZN(P1_U3342) );
  OAI21_X1 U8693 ( .B1(n6981), .B2(n6980), .A(n6979), .ZN(n6983) );
  NAND2_X1 U8694 ( .A1(n9899), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n6982) );
  NAND2_X1 U8695 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7576) );
  OAI211_X1 U8696 ( .C1(n9843), .C2(n6983), .A(n6982), .B(n7576), .ZN(n6984)
         );
  AOI21_X1 U8697 ( .B1(n9905), .B2(n6985), .A(n6984), .ZN(n6990) );
  OAI211_X1 U8698 ( .C1(n6988), .C2(n6987), .A(n9901), .B(n6986), .ZN(n6989)
         );
  NAND2_X1 U8699 ( .A1(n6990), .A2(n6989), .ZN(P2_U3254) );
  OAI211_X1 U8700 ( .C1(n6993), .C2(n6992), .A(n9901), .B(n6991), .ZN(n7002)
         );
  INV_X1 U8701 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n6998) );
  OAI211_X1 U8702 ( .C1(n6996), .C2(n6995), .A(n9906), .B(n6994), .ZN(n6997)
         );
  NAND2_X1 U8703 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n7820) );
  OAI211_X1 U8704 ( .C1(n9566), .C2(n6998), .A(n6997), .B(n7820), .ZN(n6999)
         );
  AOI21_X1 U8705 ( .B1(n7000), .B2(n9905), .A(n6999), .ZN(n7001) );
  NAND2_X1 U8706 ( .A1(n7002), .A2(n7001), .ZN(P2_U3255) );
  NOR2_X1 U8707 ( .A1(n7023), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7009) );
  NAND2_X1 U8708 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n7021), .ZN(n7008) );
  INV_X1 U8709 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7006) );
  OR2_X1 U8710 ( .A1(n7017), .A2(n7003), .ZN(n7004) );
  NAND2_X1 U8711 ( .A1(n7005), .A2(n7004), .ZN(n8104) );
  MUX2_X1 U8712 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n7006), .S(n7019), .Z(n8103)
         );
  NOR2_X1 U8713 ( .A1(n8104), .A2(n8103), .ZN(n8102) );
  AOI21_X1 U8714 ( .B1(n7006), .B2(n7019), .A(n8102), .ZN(n9707) );
  MUX2_X1 U8715 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n7007), .S(n7021), .Z(n9706)
         );
  NAND2_X1 U8716 ( .A1(n9707), .A2(n9706), .ZN(n9705) );
  NAND2_X1 U8717 ( .A1(n7008), .A2(n9705), .ZN(n7071) );
  AOI22_X1 U8718 ( .A1(n7023), .A2(n6190), .B1(P1_REG1_REG_6__SCAN_IN), .B2(
        n7075), .ZN(n7070) );
  NOR2_X1 U8719 ( .A1(n7071), .A2(n7070), .ZN(n7069) );
  NOR2_X1 U8720 ( .A1(n7009), .A2(n7069), .ZN(n7012) );
  AOI22_X1 U8721 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n7010), .B1(n7050), .B2(
        n6207), .ZN(n7011) );
  NOR2_X1 U8722 ( .A1(n7012), .A2(n7011), .ZN(n7041) );
  AOI21_X1 U8723 ( .B1(n7012), .B2(n7011), .A(n7041), .ZN(n7029) );
  AND2_X1 U8724 ( .A1(n4476), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7590) );
  INV_X1 U8725 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7013) );
  NOR2_X1 U8726 ( .A1(n9806), .A2(n7013), .ZN(n7014) );
  AOI211_X1 U8727 ( .C1(n9796), .C2(n7050), .A(n7590), .B(n7014), .ZN(n7028)
         );
  NOR2_X1 U8728 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n7050), .ZN(n7015) );
  AOI21_X1 U8729 ( .B1(n7050), .B2(P1_REG2_REG_7__SCAN_IN), .A(n7015), .ZN(
        n7025) );
  OAI21_X1 U8730 ( .B1(n7018), .B2(n7017), .A(n7016), .ZN(n8105) );
  MUX2_X1 U8731 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6147), .S(n7019), .Z(n8106)
         );
  NOR2_X1 U8732 ( .A1(n8105), .A2(n8106), .ZN(n9702) );
  INV_X1 U8733 ( .A(n7019), .ZN(n8111) );
  NOR2_X1 U8734 ( .A1(n8111), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9701) );
  NOR2_X1 U8735 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n7021), .ZN(n7020) );
  AOI21_X1 U8736 ( .B1(n7021), .B2(P1_REG2_REG_5__SCAN_IN), .A(n7020), .ZN(
        n9700) );
  OAI21_X1 U8737 ( .B1(n9702), .B2(n9701), .A(n9700), .ZN(n9699) );
  OAI21_X1 U8738 ( .B1(n7021), .B2(P1_REG2_REG_5__SCAN_IN), .A(n9699), .ZN(
        n7068) );
  NAND2_X1 U8739 ( .A1(n7023), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7022) );
  OAI21_X1 U8740 ( .B1(n7023), .B2(P1_REG2_REG_6__SCAN_IN), .A(n7022), .ZN(
        n7067) );
  NOR2_X1 U8741 ( .A1(n7068), .A2(n7067), .ZN(n7066) );
  OAI21_X1 U8742 ( .B1(n7025), .B2(n7024), .A(n7049), .ZN(n7026) );
  NAND2_X1 U8743 ( .A1(n7026), .A2(n9720), .ZN(n7027) );
  OAI211_X1 U8744 ( .C1(n7029), .C2(n9802), .A(n7028), .B(n7027), .ZN(P1_U3248) );
  INV_X1 U8745 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10038) );
  XNOR2_X1 U8746 ( .A(n7031), .B(n7030), .ZN(n7038) );
  AOI22_X1 U8747 ( .A1(n9796), .A2(n7032), .B1(n4476), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n7037) );
  OAI211_X1 U8748 ( .C1(n7035), .C2(n7034), .A(n9720), .B(n7033), .ZN(n7036)
         );
  OAI211_X1 U8749 ( .C1(n9802), .C2(n7038), .A(n7037), .B(n7036), .ZN(n7039)
         );
  INV_X1 U8750 ( .A(n7039), .ZN(n7040) );
  OAI21_X1 U8751 ( .B1(n10038), .B2(n9806), .A(n7040), .ZN(P1_U3242) );
  NOR2_X1 U8752 ( .A1(n7053), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7043) );
  INV_X1 U8753 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7847) );
  MUX2_X1 U8754 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n7847), .S(n7051), .Z(n9723)
         );
  NOR2_X1 U8755 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n7050), .ZN(n7042) );
  NOR2_X1 U8756 ( .A1(n7042), .A2(n7041), .ZN(n9724) );
  NAND2_X1 U8757 ( .A1(n9723), .A2(n9724), .ZN(n9722) );
  OAI21_X1 U8758 ( .B1(n7847), .B2(n9712), .A(n9722), .ZN(n7083) );
  AOI22_X1 U8759 ( .A1(n7053), .A2(n6251), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n7084), .ZN(n7082) );
  NOR2_X1 U8760 ( .A1(n7083), .A2(n7082), .ZN(n7081) );
  NOR2_X1 U8761 ( .A1(n7043), .A2(n7081), .ZN(n7125) );
  AOI22_X1 U8762 ( .A1(n7055), .A2(n6266), .B1(P1_REG1_REG_10__SCAN_IN), .B2(
        n7128), .ZN(n7124) );
  NOR2_X1 U8763 ( .A1(n7125), .A2(n7124), .ZN(n7123) );
  AOI21_X1 U8764 ( .B1(n7128), .B2(n6266), .A(n7123), .ZN(n7045) );
  AOI22_X1 U8765 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n7046), .B1(n7714), .B2(
        n6284), .ZN(n7044) );
  NOR2_X1 U8766 ( .A1(n7045), .A2(n7044), .ZN(n7705) );
  AOI21_X1 U8767 ( .B1(n7045), .B2(n7044), .A(n7705), .ZN(n7061) );
  INV_X1 U8768 ( .A(n9806), .ZN(n9694) );
  AND2_X1 U8769 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7934) );
  INV_X1 U8770 ( .A(n9796), .ZN(n9713) );
  NOR2_X1 U8771 ( .A1(n9713), .A2(n7046), .ZN(n7047) );
  AOI211_X1 U8772 ( .C1(n9694), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n7934), .B(
        n7047), .ZN(n7060) );
  NOR2_X1 U8773 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n7714), .ZN(n7048) );
  AOI21_X1 U8774 ( .B1(n7714), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7048), .ZN(
        n7057) );
  AOI22_X1 U8775 ( .A1(n7051), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7760), .B2(
        n9712), .ZN(n9718) );
  OAI21_X1 U8776 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n7051), .A(n9717), .ZN(
        n7087) );
  NAND2_X1 U8777 ( .A1(n7053), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7052) );
  OAI21_X1 U8778 ( .B1(n7053), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7052), .ZN(
        n7086) );
  NOR2_X1 U8779 ( .A1(n7087), .A2(n7086), .ZN(n7085) );
  NAND2_X1 U8780 ( .A1(n7055), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7054) );
  OAI21_X1 U8781 ( .B1(n7055), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7054), .ZN(
        n7130) );
  OAI21_X1 U8782 ( .B1(n7057), .B2(n7056), .A(n7713), .ZN(n7058) );
  NAND2_X1 U8783 ( .A1(n7058), .A2(n9720), .ZN(n7059) );
  OAI211_X1 U8784 ( .C1(n7061), .C2(n9802), .A(n7060), .B(n7059), .ZN(P1_U3252) );
  OR2_X1 U8785 ( .A1(n10036), .A2(n6930), .ZN(n7064) );
  OAI21_X1 U8786 ( .B1(n10033), .B2(n7065), .A(n7064), .ZN(P2_U3521) );
  INV_X1 U8787 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n7080) );
  AOI211_X1 U8788 ( .C1(n7068), .C2(n7067), .A(n7066), .B(n9790), .ZN(n7078)
         );
  AOI21_X1 U8789 ( .B1(n7071), .B2(n7070), .A(n7069), .ZN(n7072) );
  NOR2_X1 U8790 ( .A1(n9802), .A2(n7072), .ZN(n7077) );
  NOR2_X1 U8791 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7073), .ZN(n7527) );
  INV_X1 U8792 ( .A(n7527), .ZN(n7074) );
  OAI21_X1 U8793 ( .B1(n9713), .B2(n7075), .A(n7074), .ZN(n7076) );
  NOR3_X1 U8794 ( .A1(n7078), .A2(n7077), .A3(n7076), .ZN(n7079) );
  OAI21_X1 U8795 ( .B1(n9806), .B2(n7080), .A(n7079), .ZN(P1_U3247) );
  AOI21_X1 U8796 ( .B1(n7083), .B2(n7082), .A(n7081), .ZN(n7091) );
  NAND2_X1 U8797 ( .A1(n4476), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7833) );
  OAI21_X1 U8798 ( .B1(n9713), .B2(n7084), .A(n7833), .ZN(n7089) );
  AOI211_X1 U8799 ( .C1(n7087), .C2(n7086), .A(n7085), .B(n9790), .ZN(n7088)
         );
  AOI211_X1 U8800 ( .C1(n9694), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n7089), .B(
        n7088), .ZN(n7090) );
  OAI21_X1 U8801 ( .B1(n7091), .B2(n9802), .A(n7090), .ZN(P1_U3250) );
  AOI211_X1 U8802 ( .C1(n7094), .C2(n7093), .A(n7092), .B(n9841), .ZN(n7103)
         );
  OAI21_X1 U8803 ( .B1(n7097), .B2(n7096), .A(n7095), .ZN(n7101) );
  NAND2_X1 U8804 ( .A1(n9905), .A2(n7098), .ZN(n7100) );
  AND2_X1 U8805 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7391) );
  AOI21_X1 U8806 ( .B1(n9899), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7391), .ZN(
        n7099) );
  OAI211_X1 U8807 ( .C1(n9843), .C2(n7101), .A(n7100), .B(n7099), .ZN(n7102)
         );
  OR2_X1 U8808 ( .A1(n7103), .A2(n7102), .ZN(P2_U3252) );
  INV_X1 U8809 ( .A(n7104), .ZN(n7136) );
  AOI22_X1 U8810 ( .A1(n9734), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9539), .ZN(n7105) );
  OAI21_X1 U8811 ( .B1(n7136), .B2(n8089), .A(n7105), .ZN(P1_U3341) );
  INV_X1 U8812 ( .A(n7111), .ZN(n7214) );
  NOR2_X1 U8813 ( .A1(n7106), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7108) );
  NOR2_X1 U8814 ( .A1(n7108), .A2(n7107), .ZN(n7110) );
  INV_X1 U8815 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7733) );
  MUX2_X1 U8816 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n7733), .S(n7111), .Z(n7109)
         );
  NAND2_X1 U8817 ( .A1(n7111), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7210) );
  OAI211_X1 U8818 ( .C1(n7111), .C2(P2_REG2_REG_12__SCAN_IN), .A(n7110), .B(
        n7210), .ZN(n7209) );
  OAI211_X1 U8819 ( .C1(n7110), .C2(n7109), .A(n7209), .B(n9901), .ZN(n7122)
         );
  INV_X1 U8820 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10034) );
  MUX2_X1 U8821 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n10034), .S(n7111), .Z(n7117) );
  OAI21_X1 U8822 ( .B1(n6944), .B2(n7113), .A(n7112), .ZN(n7114) );
  INV_X1 U8823 ( .A(n7114), .ZN(n7116) );
  INV_X1 U8824 ( .A(n7213), .ZN(n7115) );
  OAI21_X1 U8825 ( .B1(n7117), .B2(n7116), .A(n7115), .ZN(n7120) );
  INV_X1 U8826 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7118) );
  NAND2_X1 U8827 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7903) );
  OAI21_X1 U8828 ( .B1(n9566), .B2(n7118), .A(n7903), .ZN(n7119) );
  AOI21_X1 U8829 ( .B1(n9906), .B2(n7120), .A(n7119), .ZN(n7121) );
  OAI211_X1 U8830 ( .C1(n9842), .C2(n7214), .A(n7122), .B(n7121), .ZN(P2_U3257) );
  AOI21_X1 U8831 ( .B1(n7125), .B2(n7124), .A(n7123), .ZN(n7135) );
  NOR2_X1 U8832 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7126), .ZN(n7894) );
  INV_X1 U8833 ( .A(n7894), .ZN(n7127) );
  OAI21_X1 U8834 ( .B1(n9713), .B2(n7128), .A(n7127), .ZN(n7133) );
  AOI211_X1 U8835 ( .C1(n7131), .C2(n7130), .A(n7129), .B(n9790), .ZN(n7132)
         );
  AOI211_X1 U8836 ( .C1(P1_ADDR_REG_10__SCAN_IN), .C2(n9694), .A(n7133), .B(
        n7132), .ZN(n7134) );
  OAI21_X1 U8837 ( .B1(n7135), .B2(n9802), .A(n7134), .ZN(P1_U3251) );
  OAI222_X1 U8838 ( .A1(n8980), .A2(n7137), .B1(n8968), .B2(n7136), .C1(
        P2_U3152), .C2(n7214), .ZN(P2_U3346) );
  INV_X1 U8839 ( .A(n8561), .ZN(n7204) );
  NAND2_X1 U8840 ( .A1(n7138), .A2(n7266), .ZN(n7225) );
  INV_X1 U8841 ( .A(n7225), .ZN(n7140) );
  INV_X1 U8842 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7139) );
  OAI22_X1 U8843 ( .A1(n5785), .A2(n7141), .B1(n7140), .B2(n7139), .ZN(n7142)
         );
  AOI21_X1 U8844 ( .B1(n8516), .B2(n5806), .A(n7142), .ZN(n7147) );
  OAI21_X1 U8845 ( .B1(n7144), .B2(n7143), .A(n7227), .ZN(n7145) );
  NAND2_X1 U8846 ( .A1(n9611), .A2(n7145), .ZN(n7146) );
  OAI211_X1 U8847 ( .C1(n7204), .C2(n8526), .A(n7147), .B(n7146), .ZN(P2_U3224) );
  INV_X1 U8848 ( .A(n9139), .ZN(n7156) );
  NAND2_X1 U8849 ( .A1(n7148), .A2(n9115), .ZN(n7155) );
  OAI21_X1 U8850 ( .B1(n7150), .B2(n9826), .A(n7149), .ZN(n7153) );
  INV_X1 U8851 ( .A(n7151), .ZN(n7152) );
  NAND2_X1 U8852 ( .A1(n7153), .A2(n7152), .ZN(n7242) );
  AOI22_X1 U8853 ( .A1(n7242), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n7538), .B2(
        n9095), .ZN(n7154) );
  OAI211_X1 U8854 ( .C1(n7156), .C2(n9117), .A(n7155), .B(n7154), .ZN(P1_U3230) );
  INV_X1 U8855 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7171) );
  NAND2_X1 U8856 ( .A1(n7158), .A2(n7157), .ZN(n7329) );
  NAND2_X1 U8857 ( .A1(n7329), .A2(n7328), .ZN(n7327) );
  INV_X1 U8858 ( .A(n9952), .ZN(n7344) );
  OR2_X1 U8859 ( .A1(n5806), .A2(n7344), .ZN(n7159) );
  NAND2_X1 U8860 ( .A1(n7327), .A2(n7159), .ZN(n7161) );
  INV_X1 U8861 ( .A(n7160), .ZN(n7164) );
  NAND2_X1 U8862 ( .A1(n7161), .A2(n7164), .ZN(n7263) );
  OAI21_X1 U8863 ( .B1(n7161), .B2(n7164), .A(n7263), .ZN(n7471) );
  INV_X1 U8864 ( .A(n7471), .ZN(n7169) );
  INV_X1 U8865 ( .A(n7877), .ZN(n9922) );
  INV_X1 U8866 ( .A(n5806), .ZN(n7162) );
  OAI22_X1 U8867 ( .A1(n7162), .A2(n8818), .B1(n5809), .B2(n8820), .ZN(n7167)
         );
  XNOR2_X1 U8868 ( .A(n7164), .B(n7163), .ZN(n7165) );
  NOR2_X1 U8869 ( .A1(n7165), .A2(n9917), .ZN(n7166) );
  AOI211_X1 U8870 ( .C1(n9922), .C2(n7471), .A(n7167), .B(n7166), .ZN(n7473)
         );
  AOI21_X1 U8871 ( .B1(n7467), .B2(n4781), .A(n4512), .ZN(n7466) );
  AOI22_X1 U8872 ( .A1(n7466), .A2(n6882), .B1(n8930), .B2(n7467), .ZN(n7168)
         );
  OAI211_X1 U8873 ( .C1(n7169), .C2(n8939), .A(n7473), .B(n7168), .ZN(n7172)
         );
  NAND2_X1 U8874 ( .A1(n7172), .A2(n10021), .ZN(n7170) );
  OAI21_X1 U8875 ( .B1(n10021), .B2(n7171), .A(n7170), .ZN(P2_U3460) );
  NAND2_X1 U8876 ( .A1(n7172), .A2(n10036), .ZN(n7173) );
  OAI21_X1 U8877 ( .B1(n10036), .B2(n6928), .A(n7173), .ZN(P2_U3523) );
  INV_X1 U8878 ( .A(n7174), .ZN(n7182) );
  INV_X1 U8879 ( .A(n7221), .ZN(n7291) );
  OAI222_X1 U8880 ( .A1(n8968), .A2(n7182), .B1(n7291), .B2(P2_U3152), .C1(
        n7175), .C2(n8980), .ZN(P2_U3345) );
  INV_X1 U8881 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9401) );
  NOR2_X1 U8882 ( .A1(n6458), .A2(n9401), .ZN(n7179) );
  INV_X1 U8883 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n7176) );
  NOR2_X1 U8884 ( .A1(n6501), .A2(n7176), .ZN(n7178) );
  INV_X1 U8885 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9491) );
  NOR2_X1 U8886 ( .A1(n6145), .A2(n9491), .ZN(n7177) );
  NAND2_X1 U8887 ( .A1(n9175), .A2(P1_U4006), .ZN(n7180) );
  OAI21_X1 U8888 ( .B1(P1_U4006), .B2(n5851), .A(n7180), .ZN(P1_U3586) );
  NAND2_X1 U8889 ( .A1(n9279), .A2(P1_U4006), .ZN(n7181) );
  OAI21_X1 U8890 ( .B1(n5657), .B2(P1_U4006), .A(n7181), .ZN(P1_U3577) );
  INV_X1 U8891 ( .A(n9747), .ZN(n7709) );
  OAI222_X1 U8892 ( .A1(P1_U3084), .A2(n7709), .B1(n8089), .B2(n7182), .C1(
        n10316), .C2(n9549), .ZN(P1_U3340) );
  INV_X1 U8893 ( .A(n7183), .ZN(n7186) );
  INV_X1 U8894 ( .A(n7448), .ZN(n7454) );
  OAI222_X1 U8895 ( .A1(n8968), .A2(n7186), .B1(n7454), .B2(P2_U3152), .C1(
        n7184), .C2(n8980), .ZN(P2_U3344) );
  INV_X1 U8896 ( .A(n7720), .ZN(n9152) );
  OAI222_X1 U8897 ( .A1(n4476), .A2(n9152), .B1(n8089), .B2(n7186), .C1(n7185), 
        .C2(n9549), .ZN(P1_U3339) );
  INV_X1 U8898 ( .A(n7510), .ZN(n7193) );
  NAND2_X1 U8899 ( .A1(n6694), .A2(n7538), .ZN(n7189) );
  AND3_X1 U8900 ( .A1(n7376), .A2(n9467), .A3(n7189), .ZN(n7511) );
  INV_X1 U8901 ( .A(n9138), .ZN(n7192) );
  INV_X1 U8902 ( .A(n6696), .ZN(n7191) );
  OAI222_X1 U8903 ( .A1(n9646), .A2(n7192), .B1(n9644), .B2(n7191), .C1(n7190), 
        .C2(n9326), .ZN(n7516) );
  AOI211_X1 U8904 ( .C1(n7193), .C2(n9822), .A(n7511), .B(n7516), .ZN(n7258)
         );
  INV_X1 U8905 ( .A(n9486), .ZN(n7626) );
  AOI22_X1 U8906 ( .A1(n7626), .A2(n6694), .B1(P1_REG1_REG_1__SCAN_IN), .B2(
        n9838), .ZN(n7194) );
  OAI21_X1 U8907 ( .B1(n7258), .B2(n9838), .A(n7194), .ZN(P1_U3524) );
  XNOR2_X1 U8908 ( .A(n7196), .B(n7195), .ZN(n7197) );
  XNOR2_X1 U8909 ( .A(n7198), .B(n7197), .ZN(n7202) );
  OAI22_X1 U8910 ( .A1(n5809), .A2(n8818), .B1(n7410), .B2(n8820), .ZN(n7282)
         );
  NAND2_X1 U8911 ( .A1(n9606), .A2(n7282), .ZN(n7199) );
  NAND2_X1 U8912 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9553) );
  OAI211_X1 U8913 ( .C1(n9616), .C2(n7277), .A(n7199), .B(n9553), .ZN(n7200)
         );
  AOI21_X1 U8914 ( .B1(n9610), .B2(n7272), .A(n7200), .ZN(n7201) );
  OAI21_X1 U8915 ( .B1(n7202), .B2(n8542), .A(n7201), .ZN(P2_U3229) );
  NAND2_X1 U8916 ( .A1(n9611), .A2(n7337), .ZN(n8505) );
  OAI22_X1 U8917 ( .A1(n8505), .A2(n7204), .B1(n7203), .B2(n8542), .ZN(n7206)
         );
  NAND2_X1 U8918 ( .A1(n7206), .A2(n7205), .ZN(n7208) );
  AOI22_X1 U8919 ( .A1(n9610), .A2(n9946), .B1(n7225), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n7207) );
  OAI211_X1 U8920 ( .C1(n5804), .C2(n8527), .A(n7208), .B(n7207), .ZN(P2_U3234) );
  NAND2_X1 U8921 ( .A1(n7210), .A2(n7209), .ZN(n7212) );
  AOI22_X1 U8922 ( .A1(n7221), .A2(n7879), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7291), .ZN(n7211) );
  NOR2_X1 U8923 ( .A1(n7212), .A2(n7211), .ZN(n7286) );
  AOI21_X1 U8924 ( .B1(n7212), .B2(n7211), .A(n7286), .ZN(n7223) );
  AOI21_X1 U8925 ( .B1(n10034), .B2(n7214), .A(n7213), .ZN(n7216) );
  AOI22_X1 U8926 ( .A1(n7221), .A2(n7290), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7291), .ZN(n7215) );
  NOR2_X1 U8927 ( .A1(n7216), .A2(n7215), .ZN(n7289) );
  AOI21_X1 U8928 ( .B1(n7216), .B2(n7215), .A(n7289), .ZN(n7219) );
  NOR2_X1 U8929 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5497), .ZN(n7217) );
  AOI21_X1 U8930 ( .B1(n9899), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n7217), .ZN(
        n7218) );
  OAI21_X1 U8931 ( .B1(n7219), .B2(n9843), .A(n7218), .ZN(n7220) );
  AOI21_X1 U8932 ( .B1(n7221), .B2(n9905), .A(n7220), .ZN(n7222) );
  OAI21_X1 U8933 ( .B1(n7223), .B2(n9841), .A(n7222), .ZN(P2_U3258) );
  AOI22_X1 U8934 ( .A1(n8750), .A2(n5805), .B1(n5807), .B2(n8751), .ZN(n7334)
         );
  OAI22_X1 U8935 ( .A1(n5785), .A2(n9952), .B1(n7334), .B2(n8481), .ZN(n7224)
         );
  AOI21_X1 U8936 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n7225), .A(n7224), .ZN(
        n7231) );
  INV_X1 U8937 ( .A(n7226), .ZN(n7228) );
  NAND3_X1 U8938 ( .A1(n7229), .A2(n7228), .A3(n7227), .ZN(n7230) );
  OAI211_X1 U8939 ( .C1(n8542), .C2(n7232), .A(n7231), .B(n7230), .ZN(P2_U3239) );
  XOR2_X1 U8940 ( .A(n7234), .B(n7233), .Z(n7237) );
  AOI22_X1 U8941 ( .A1(n7242), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n4479), .B2(
        n9095), .ZN(n7236) );
  AOI22_X1 U8942 ( .A1(n9108), .A2(n6701), .B1(n9120), .B2(n9139), .ZN(n7235)
         );
  OAI211_X1 U8943 ( .C1(n7237), .C2(n9097), .A(n7236), .B(n7235), .ZN(P1_U3235) );
  XNOR2_X1 U8944 ( .A(n7239), .B(n7238), .ZN(n7240) );
  XNOR2_X1 U8945 ( .A(n7241), .B(n7240), .ZN(n7245) );
  AOI22_X1 U8946 ( .A1(n7242), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n6694), .B2(
        n9095), .ZN(n7244) );
  AOI22_X1 U8947 ( .A1(n9108), .A2(n9138), .B1(n9120), .B2(n6696), .ZN(n7243)
         );
  OAI211_X1 U8948 ( .C1(n7245), .C2(n9097), .A(n7244), .B(n7243), .ZN(P1_U3220) );
  XOR2_X1 U8949 ( .A(n7246), .B(n7247), .Z(n7253) );
  INV_X1 U8950 ( .A(n9095), .ZN(n9123) );
  NOR2_X1 U8951 ( .A1(n9123), .A2(n9811), .ZN(n7248) );
  AOI211_X1 U8952 ( .C1(n9120), .C2(n9138), .A(n7249), .B(n7248), .ZN(n7252)
         );
  INV_X1 U8953 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7250) );
  AOI22_X1 U8954 ( .A1(n9108), .A2(n9137), .B1(n7250), .B2(n9103), .ZN(n7251)
         );
  OAI211_X1 U8955 ( .C1(n7253), .C2(n9097), .A(n7252), .B(n7251), .ZN(P1_U3216) );
  NAND2_X1 U8956 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n8560), .ZN(n7254) );
  OAI21_X1 U8957 ( .B1(n8654), .B2(n8560), .A(n7254), .ZN(P2_U3579) );
  INV_X1 U8958 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7255) );
  OAI22_X1 U8959 ( .A1(n9532), .A2(n6742), .B1(n9835), .B2(n7255), .ZN(n7256)
         );
  INV_X1 U8960 ( .A(n7256), .ZN(n7257) );
  OAI21_X1 U8961 ( .B1(n7258), .B2(n9833), .A(n7257), .ZN(P1_U3457) );
  INV_X1 U8962 ( .A(n7259), .ZN(n7261) );
  INV_X1 U8963 ( .A(n7636), .ZN(n7458) );
  OAI222_X1 U8964 ( .A1(n8980), .A2(n7260), .B1(n8968), .B2(n7261), .C1(
        P2_U3152), .C2(n7458), .ZN(P2_U3343) );
  INV_X1 U8965 ( .A(n9759), .ZN(n9153) );
  OAI222_X1 U8966 ( .A1(n9153), .A2(P1_U3084), .B1(n8089), .B2(n7261), .C1(
        n10213), .C2(n9549), .ZN(P1_U3338) );
  OR2_X1 U8967 ( .A1(n5807), .A2(n7467), .ZN(n7262) );
  NAND2_X1 U8968 ( .A1(n7263), .A2(n7262), .ZN(n7441) );
  NAND2_X1 U8969 ( .A1(n7441), .A2(n7440), .ZN(n7439) );
  NAND2_X1 U8970 ( .A1(n5809), .A2(n9958), .ZN(n7264) );
  NAND2_X1 U8971 ( .A1(n7439), .A2(n7264), .ZN(n7397) );
  XNOR2_X1 U8972 ( .A(n7397), .B(n7396), .ZN(n9968) );
  NAND3_X1 U8973 ( .A1(n7267), .A2(n7266), .A3(n7265), .ZN(n7338) );
  INV_X1 U8974 ( .A(n7268), .ZN(n7269) );
  OR2_X1 U8975 ( .A1(n7270), .A2(n8835), .ZN(n7463) );
  NAND2_X1 U8976 ( .A1(n7877), .A2(n7463), .ZN(n7271) );
  AND2_X1 U8977 ( .A1(n8839), .A2(n8835), .ZN(n8701) );
  AOI21_X1 U8978 ( .B1(n7442), .B2(n7272), .A(n10013), .ZN(n7273) );
  NAND2_X1 U8979 ( .A1(n7273), .A2(n7425), .ZN(n9964) );
  INV_X1 U8980 ( .A(n9964), .ZN(n7274) );
  AND2_X1 U8981 ( .A1(n8701), .A2(n7274), .ZN(n7279) );
  AND2_X1 U8982 ( .A1(n9947), .A2(n7275), .ZN(n7276) );
  OAI22_X1 U8983 ( .A1(n8813), .A2(n9966), .B1(n7277), .B2(n8836), .ZN(n7278)
         );
  AOI211_X1 U8984 ( .C1(n9968), .C2(n8736), .A(n7279), .B(n7278), .ZN(n7285)
         );
  NAND2_X1 U8985 ( .A1(n7436), .A2(n7280), .ZN(n7281) );
  XNOR2_X1 U8986 ( .A(n7281), .B(n7396), .ZN(n7283) );
  AOI21_X1 U8987 ( .B1(n7283), .B2(n8795), .A(n7282), .ZN(n9965) );
  MUX2_X1 U8988 ( .A(n9965), .B(n6903), .S(n9936), .Z(n7284) );
  NAND2_X1 U8989 ( .A1(n7285), .A2(n7284), .ZN(P2_U3291) );
  AOI21_X1 U8990 ( .B1(n7291), .B2(n7879), .A(n7286), .ZN(n7288) );
  AOI22_X1 U8991 ( .A1(n7448), .A2(n7926), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7454), .ZN(n7287) );
  NOR2_X1 U8992 ( .A1(n7288), .A2(n7287), .ZN(n7449) );
  AOI21_X1 U8993 ( .B1(n7288), .B2(n7287), .A(n7449), .ZN(n7300) );
  AOI21_X1 U8994 ( .B1(n7291), .B2(n7290), .A(n7289), .ZN(n7293) );
  AOI22_X1 U8995 ( .A1(n7448), .A2(n7453), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n7454), .ZN(n7292) );
  NOR2_X1 U8996 ( .A1(n7293), .A2(n7292), .ZN(n7452) );
  AOI21_X1 U8997 ( .B1(n7293), .B2(n7292), .A(n7452), .ZN(n7294) );
  NOR2_X1 U8998 ( .A1(n7294), .A2(n9843), .ZN(n7298) );
  NOR2_X1 U8999 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10318), .ZN(n7295) );
  AOI21_X1 U9000 ( .B1(n9899), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n7295), .ZN(
        n7296) );
  OAI21_X1 U9001 ( .B1(n9842), .B2(n7454), .A(n7296), .ZN(n7297) );
  NOR2_X1 U9002 ( .A1(n7298), .A2(n7297), .ZN(n7299) );
  OAI21_X1 U9003 ( .B1(n7300), .B2(n9841), .A(n7299), .ZN(P2_U3259) );
  XOR2_X1 U9004 ( .A(n7302), .B(n7301), .Z(n7306) );
  INV_X1 U9005 ( .A(n7485), .ZN(n8556) );
  AOI22_X1 U9006 ( .A1(n8556), .A2(n8751), .B1(n8750), .B2(n8558), .ZN(n7419)
         );
  NAND2_X1 U9007 ( .A1(P2_U3152), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9872) );
  OAI21_X1 U9008 ( .B1(n8481), .B2(n7419), .A(n9872), .ZN(n7304) );
  NOR2_X1 U9009 ( .A1(n9616), .A2(n7429), .ZN(n7303) );
  AOI211_X1 U9010 ( .C1(n9610), .C2(n7431), .A(n7304), .B(n7303), .ZN(n7305)
         );
  OAI21_X1 U9011 ( .B1(n7306), .B2(n8542), .A(n7305), .ZN(P2_U3241) );
  XNOR2_X1 U9012 ( .A(n7308), .B(n7307), .ZN(n7309) );
  INV_X1 U9013 ( .A(n7503), .ZN(n7310) );
  AOI22_X1 U9014 ( .A1(n9108), .A2(n9135), .B1(n7310), .B2(n9103), .ZN(n7314)
         );
  NAND2_X1 U9015 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9710) );
  INV_X1 U9016 ( .A(n9710), .ZN(n7312) );
  NOR2_X1 U9017 ( .A1(n9123), .A2(n9818), .ZN(n7311) );
  AOI211_X1 U9018 ( .C1(n9120), .C2(n9137), .A(n7312), .B(n7311), .ZN(n7313)
         );
  OAI211_X1 U9019 ( .C1(n7315), .C2(n9097), .A(n7314), .B(n7313), .ZN(P1_U3225) );
  INV_X1 U9020 ( .A(n7316), .ZN(n7357) );
  AOI22_X1 U9021 ( .A1(n9770), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9539), .ZN(n7317) );
  OAI21_X1 U9022 ( .B1(n7357), .B2(n8089), .A(n7317), .ZN(P1_U3337) );
  INV_X1 U9023 ( .A(n7319), .ZN(n7320) );
  AOI211_X1 U9024 ( .C1(n7321), .C2(n7318), .A(n9097), .B(n7320), .ZN(n7326)
         );
  INV_X1 U9025 ( .A(n9136), .ZN(n7674) );
  INV_X1 U9026 ( .A(n7322), .ZN(n7660) );
  AOI22_X1 U9027 ( .A1(n9120), .A2(n6701), .B1(n7660), .B2(n9103), .ZN(n7324)
         );
  AND2_X1 U9028 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n8110) );
  AOI21_X1 U9029 ( .B1(n9095), .B2(n7661), .A(n8110), .ZN(n7323) );
  OAI211_X1 U9030 ( .C1(n7674), .C2(n9117), .A(n7324), .B(n7323), .ZN(n7325)
         );
  OR2_X1 U9031 ( .A1(n7326), .A2(n7325), .ZN(P1_U3228) );
  OAI21_X1 U9032 ( .B1(n7329), .B2(n7328), .A(n7327), .ZN(n9956) );
  INV_X1 U9033 ( .A(n9956), .ZN(n7347) );
  OAI21_X1 U9034 ( .B1(n7332), .B2(n7331), .A(n7330), .ZN(n7333) );
  NAND2_X1 U9035 ( .A1(n7333), .A2(n8795), .ZN(n7335) );
  NAND2_X1 U9036 ( .A1(n7335), .A2(n7334), .ZN(n9954) );
  INV_X1 U9037 ( .A(n9954), .ZN(n7336) );
  MUX2_X1 U9038 ( .A(n7336), .B(n6896), .S(n9936), .Z(n7346) );
  AND2_X1 U9039 ( .A1(n7339), .A2(n7344), .ZN(n7341) );
  OR2_X1 U9040 ( .A1(n7341), .A2(n7340), .ZN(n9953) );
  INV_X1 U9041 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7342) );
  OAI22_X1 U9042 ( .A1(n8717), .A2(n9953), .B1(n7342), .B2(n8836), .ZN(n7343)
         );
  AOI21_X1 U9043 ( .B1(n9926), .B2(n7344), .A(n7343), .ZN(n7345) );
  OAI211_X1 U9044 ( .C1(n7347), .C2(n8843), .A(n7346), .B(n7345), .ZN(P2_U3294) );
  INV_X1 U9045 ( .A(n7348), .ZN(n7356) );
  OAI22_X1 U9046 ( .A1(n7139), .A2(n8836), .B1(n6898), .B2(n8839), .ZN(n7351)
         );
  NOR2_X1 U9047 ( .A1(n8717), .A2(n7349), .ZN(n7350) );
  AOI211_X1 U9048 ( .C1(n9926), .C2(n7352), .A(n7351), .B(n7350), .ZN(n7355)
         );
  NAND2_X1 U9049 ( .A1(n8736), .A2(n7353), .ZN(n7354) );
  OAI211_X1 U9050 ( .C1(n9936), .C2(n7356), .A(n7355), .B(n7354), .ZN(P2_U3295) );
  INV_X1 U9051 ( .A(n7640), .ZN(n8575) );
  OAI222_X1 U9052 ( .A1(n8980), .A2(n7358), .B1(n8575), .B2(P2_U3152), .C1(
        n8983), .C2(n7357), .ZN(P2_U3342) );
  INV_X1 U9053 ( .A(n7845), .ZN(n9832) );
  OR2_X1 U9054 ( .A1(n7359), .A2(n8342), .ZN(n7360) );
  NAND2_X1 U9055 ( .A1(n7361), .A2(n7360), .ZN(n7667) );
  NAND2_X1 U9056 ( .A1(n7697), .A2(n7661), .ZN(n7362) );
  NAND2_X1 U9057 ( .A1(n7500), .A2(n7362), .ZN(n7663) );
  OAI22_X1 U9058 ( .A1(n7663), .A2(n9827), .B1(n7363), .B2(n9826), .ZN(n7367)
         );
  XNOR2_X1 U9059 ( .A(n8287), .B(n8342), .ZN(n7366) );
  INV_X1 U9060 ( .A(n9652), .ZN(n7980) );
  NAND2_X1 U9061 ( .A1(n7667), .A2(n7980), .ZN(n7365) );
  AOI22_X1 U9062 ( .A1(n9382), .A2(n6701), .B1(n9136), .B2(n9379), .ZN(n7364)
         );
  OAI211_X1 U9063 ( .C1(n9326), .C2(n7366), .A(n7365), .B(n7364), .ZN(n7664)
         );
  AOI211_X1 U9064 ( .C1(n9832), .C2(n7667), .A(n7367), .B(n7664), .ZN(n7474)
         );
  NAND2_X1 U9065 ( .A1(n9838), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7368) );
  OAI21_X1 U9066 ( .B1(n7474), .B2(n9838), .A(n7368), .ZN(P1_U3527) );
  INV_X1 U9067 ( .A(n7369), .ZN(n7370) );
  AOI21_X1 U9068 ( .B1(n8346), .B2(n7371), .A(n7370), .ZN(n7743) );
  XNOR2_X1 U9069 ( .A(n8346), .B(n7372), .ZN(n7375) );
  AOI22_X1 U9070 ( .A1(n9382), .A2(n9139), .B1(n6701), .B2(n9379), .ZN(n7373)
         );
  OAI21_X1 U9071 ( .B1(n7743), .B2(n9652), .A(n7373), .ZN(n7374) );
  AOI21_X1 U9072 ( .B1(n9649), .B2(n7375), .A(n7374), .ZN(n7748) );
  AOI21_X1 U9073 ( .B1(n4479), .B2(n7376), .A(n7695), .ZN(n7746) );
  AOI22_X1 U9074 ( .A1(n7746), .A2(n9467), .B1(n9466), .B2(n4479), .ZN(n7378)
         );
  OAI211_X1 U9075 ( .C1(n7743), .C2(n7845), .A(n7748), .B(n7378), .ZN(n7380)
         );
  NAND2_X1 U9076 ( .A1(n7380), .A2(n9840), .ZN(n7379) );
  OAI21_X1 U9077 ( .B1(n9840), .B2(n6961), .A(n7379), .ZN(P1_U3525) );
  NAND2_X1 U9078 ( .A1(n7380), .A2(n9835), .ZN(n7381) );
  OAI21_X1 U9079 ( .B1(n9835), .B2(n6110), .A(n7381), .ZN(P1_U3460) );
  INV_X1 U9080 ( .A(n9948), .ZN(n7385) );
  AOI22_X1 U9081 ( .A1(n9948), .A2(n8795), .B1(n8751), .B2(n5805), .ZN(n9950)
         );
  INV_X1 U9082 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10394) );
  OAI22_X1 U9083 ( .A1(n9936), .A2(n9950), .B1(n10394), .B2(n8836), .ZN(n7382)
         );
  AOI21_X1 U9084 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n9936), .A(n7382), .ZN(
        n7384) );
  OAI21_X1 U9085 ( .B1(n9926), .B2(n9932), .A(n9946), .ZN(n7383) );
  OAI211_X1 U9086 ( .C1(n7385), .C2(n8843), .A(n7384), .B(n7383), .ZN(P2_U3296) );
  INV_X1 U9087 ( .A(n9781), .ZN(n9158) );
  INV_X1 U9088 ( .A(n7386), .ZN(n7476) );
  INV_X1 U9089 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10090) );
  OAI222_X1 U9090 ( .A1(P1_U3084), .A2(n9158), .B1(n8089), .B2(n7476), .C1(
        n10090), .C2(n9549), .ZN(P1_U3336) );
  INV_X1 U9091 ( .A(n7480), .ZN(n7387) );
  AOI211_X1 U9092 ( .C1(n7389), .C2(n7388), .A(n8542), .B(n7387), .ZN(n7395)
         );
  INV_X1 U9093 ( .A(n7541), .ZN(n9976) );
  INV_X1 U9094 ( .A(n8526), .ZN(n8517) );
  INV_X1 U9095 ( .A(n7548), .ZN(n8555) );
  AOI22_X1 U9096 ( .A1(n8517), .A2(n8557), .B1(n8516), .B2(n8555), .ZN(n7393)
         );
  INV_X1 U9097 ( .A(n9616), .ZN(n8479) );
  INV_X1 U9098 ( .A(n7390), .ZN(n7405) );
  AOI21_X1 U9099 ( .B1(n8479), .B2(n7405), .A(n7391), .ZN(n7392) );
  OAI211_X1 U9100 ( .C1(n9976), .C2(n5785), .A(n7393), .B(n7392), .ZN(n7394)
         );
  OR2_X1 U9101 ( .A1(n7395), .A2(n7394), .ZN(P2_U3215) );
  NAND2_X1 U9102 ( .A1(n7397), .A2(n7396), .ZN(n7400) );
  NAND2_X1 U9103 ( .A1(n9966), .A2(n7398), .ZN(n7399) );
  NAND2_X1 U9104 ( .A1(n7400), .A2(n7399), .ZN(n7423) );
  INV_X1 U9105 ( .A(n7423), .ZN(n7401) );
  NAND2_X1 U9106 ( .A1(n7401), .A2(n5999), .ZN(n7421) );
  NAND2_X1 U9107 ( .A1(n7431), .A2(n8557), .ZN(n7402) );
  OAI21_X1 U9108 ( .B1(n7404), .B2(n7403), .A(n7543), .ZN(n9980) );
  NAND2_X1 U9109 ( .A1(n7426), .A2(n9976), .ZN(n9928) );
  OAI21_X1 U9110 ( .B1(n7426), .B2(n9976), .A(n9928), .ZN(n9977) );
  INV_X1 U9111 ( .A(n8836), .ZN(n9925) );
  AOI22_X1 U9112 ( .A1(n9926), .A2(n7541), .B1(n9925), .B2(n7405), .ZN(n7406)
         );
  OAI21_X1 U9113 ( .B1(n9977), .B2(n8717), .A(n7406), .ZN(n7415) );
  OAI211_X1 U9114 ( .C1(n7409), .C2(n7408), .A(n7407), .B(n8795), .ZN(n7413)
         );
  OAI22_X1 U9115 ( .A1(n7548), .A2(n8820), .B1(n7410), .B2(n8818), .ZN(n7411)
         );
  INV_X1 U9116 ( .A(n7411), .ZN(n7412) );
  NAND2_X1 U9117 ( .A1(n7413), .A2(n7412), .ZN(n9978) );
  MUX2_X1 U9118 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9978), .S(n8839), .Z(n7414)
         );
  AOI211_X1 U9119 ( .C1(n8736), .C2(n9980), .A(n7415), .B(n7414), .ZN(n7416)
         );
  INV_X1 U9120 ( .A(n7416), .ZN(P2_U3289) );
  XNOR2_X1 U9121 ( .A(n7417), .B(n7424), .ZN(n7418) );
  NAND2_X1 U9122 ( .A1(n7418), .A2(n8795), .ZN(n7420) );
  NAND2_X1 U9123 ( .A1(n7420), .A2(n7419), .ZN(n9973) );
  INV_X1 U9124 ( .A(n9973), .ZN(n7435) );
  INV_X1 U9125 ( .A(n7421), .ZN(n7422) );
  AOI21_X1 U9126 ( .B1(n7424), .B2(n7423), .A(n7422), .ZN(n9974) );
  INV_X1 U9127 ( .A(n7431), .ZN(n9970) );
  INV_X1 U9128 ( .A(n7425), .ZN(n7428) );
  INV_X1 U9129 ( .A(n7426), .ZN(n7427) );
  OAI21_X1 U9130 ( .B1(n9970), .B2(n7428), .A(n7427), .ZN(n9971) );
  OAI22_X1 U9131 ( .A1(n8839), .A2(n6894), .B1(n7429), .B2(n8836), .ZN(n7430)
         );
  AOI21_X1 U9132 ( .B1(n9926), .B2(n7431), .A(n7430), .ZN(n7432) );
  OAI21_X1 U9133 ( .B1(n9971), .B2(n8717), .A(n7432), .ZN(n7433) );
  AOI21_X1 U9134 ( .B1(n9974), .B2(n8736), .A(n7433), .ZN(n7434) );
  OAI21_X1 U9135 ( .B1(n9936), .B2(n7435), .A(n7434), .ZN(P2_U3290) );
  OAI211_X1 U9136 ( .C1(n5103), .C2(n5810), .A(n8795), .B(n7436), .ZN(n7438)
         );
  AOI22_X1 U9137 ( .A1(n8750), .A2(n5807), .B1(n8558), .B2(n8751), .ZN(n7437)
         );
  NAND2_X1 U9138 ( .A1(n7438), .A2(n7437), .ZN(n9960) );
  INV_X1 U9139 ( .A(n9960), .ZN(n7447) );
  OAI21_X1 U9140 ( .B1(n7441), .B2(n7440), .A(n7439), .ZN(n9962) );
  OAI21_X1 U9141 ( .B1(n4512), .B2(n9958), .A(n7442), .ZN(n9959) );
  OAI22_X1 U9142 ( .A1(n8513), .A2(n8836), .B1(n6902), .B2(n8839), .ZN(n7443)
         );
  AOI21_X1 U9143 ( .B1(n9926), .B2(n8515), .A(n7443), .ZN(n7444) );
  OAI21_X1 U9144 ( .B1(n8717), .B2(n9959), .A(n7444), .ZN(n7445) );
  AOI21_X1 U9145 ( .B1(n9962), .B2(n8736), .A(n7445), .ZN(n7446) );
  OAI21_X1 U9146 ( .B1(n7447), .B2(n9936), .A(n7446), .ZN(P2_U3292) );
  NOR2_X1 U9147 ( .A1(n7448), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7450) );
  NOR2_X1 U9148 ( .A1(n7450), .A2(n7449), .ZN(n7635) );
  XNOR2_X1 U9149 ( .A(n7636), .B(n7635), .ZN(n7451) );
  NOR2_X1 U9150 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7451), .ZN(n7637) );
  AOI21_X1 U9151 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n7451), .A(n7637), .ZN(
        n7462) );
  AOI21_X1 U9152 ( .B1(n7454), .B2(n7453), .A(n7452), .ZN(n7629) );
  XOR2_X1 U9153 ( .A(n7636), .B(n7629), .Z(n7455) );
  NAND2_X1 U9154 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n7455), .ZN(n7630) );
  OAI211_X1 U9155 ( .C1(n7455), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9906), .B(
        n7630), .ZN(n7461) );
  NOR2_X1 U9156 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5540), .ZN(n7456) );
  AOI21_X1 U9157 ( .B1(n9899), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7456), .ZN(
        n7457) );
  OAI21_X1 U9158 ( .B1(n9842), .B2(n7458), .A(n7457), .ZN(n7459) );
  INV_X1 U9159 ( .A(n7459), .ZN(n7460) );
  OAI211_X1 U9160 ( .C1(n7462), .C2(n9841), .A(n7461), .B(n7460), .ZN(P2_U3260) );
  INV_X1 U9161 ( .A(n7463), .ZN(n7464) );
  AOI22_X1 U9162 ( .A1(n9932), .A2(n7466), .B1(n9925), .B2(n7465), .ZN(n7469)
         );
  NAND2_X1 U9163 ( .A1(n9926), .A2(n7467), .ZN(n7468) );
  OAI211_X1 U9164 ( .C1(n6895), .C2(n8839), .A(n7469), .B(n7468), .ZN(n7470)
         );
  AOI21_X1 U9165 ( .B1(n9933), .B2(n7471), .A(n7470), .ZN(n7472) );
  OAI21_X1 U9166 ( .B1(n7473), .B2(n9936), .A(n7472), .ZN(P2_U3293) );
  OR2_X1 U9167 ( .A1(n7474), .A2(n9833), .ZN(n7475) );
  OAI21_X1 U9168 ( .B1(n9835), .B2(n6146), .A(n7475), .ZN(P1_U3466) );
  INV_X1 U9169 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7477) );
  OAI222_X1 U9170 ( .A1(n8980), .A2(n7477), .B1(n8573), .B2(P2_U3152), .C1(
        n8983), .C2(n7476), .ZN(P2_U3341) );
  INV_X1 U9171 ( .A(n9927), .ZN(n9982) );
  INV_X1 U9172 ( .A(n7478), .ZN(n7479) );
  AOI21_X1 U9173 ( .B1(n7480), .B2(n7479), .A(n8542), .ZN(n7484) );
  NOR3_X1 U9174 ( .A1(n8505), .A2(n7481), .A3(n7485), .ZN(n7483) );
  OAI21_X1 U9175 ( .B1(n7484), .B2(n7483), .A(n7482), .ZN(n7488) );
  OAI22_X1 U9176 ( .A1(n7485), .A2(n8818), .B1(n7601), .B2(n8820), .ZN(n9921)
         );
  INV_X1 U9177 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10374) );
  NOR2_X1 U9178 ( .A1(n10374), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9885) );
  NOR2_X1 U9179 ( .A1(n9616), .A2(n9923), .ZN(n7486) );
  AOI211_X1 U9180 ( .C1(n9606), .C2(n9921), .A(n9885), .B(n7486), .ZN(n7487)
         );
  OAI211_X1 U9181 ( .C1(n9982), .C2(n5785), .A(n7488), .B(n7487), .ZN(P2_U3223) );
  INV_X1 U9182 ( .A(n7497), .ZN(n8347) );
  XNOR2_X1 U9183 ( .A(n7489), .B(n7497), .ZN(n9821) );
  INV_X1 U9184 ( .A(n9821), .ZN(n7509) );
  INV_X1 U9185 ( .A(n7490), .ZN(n9535) );
  NAND2_X1 U9186 ( .A1(n7491), .A2(n9535), .ZN(n7537) );
  AND2_X1 U9187 ( .A1(n8431), .A2(n7492), .ZN(n7493) );
  INV_X1 U9188 ( .A(n9135), .ZN(n7567) );
  INV_X1 U9189 ( .A(n9137), .ZN(n7499) );
  INV_X1 U9190 ( .A(n7494), .ZN(n7495) );
  OR2_X1 U9191 ( .A1(n8287), .A2(n7495), .ZN(n8151) );
  NAND2_X1 U9192 ( .A1(n8151), .A2(n8379), .ZN(n7496) );
  NOR2_X1 U9193 ( .A1(n7496), .A2(n7497), .ZN(n7675) );
  AOI21_X1 U9194 ( .B1(n7497), .B2(n7496), .A(n7675), .ZN(n7498) );
  OAI222_X1 U9195 ( .A1(n9646), .A2(n7567), .B1(n9644), .B2(n7499), .C1(n9326), 
        .C2(n7498), .ZN(n9819) );
  INV_X1 U9196 ( .A(n7500), .ZN(n7502) );
  INV_X1 U9197 ( .A(n7501), .ZN(n7681) );
  OAI211_X1 U9198 ( .C1(n9818), .C2(n7502), .A(n7681), .B(n9467), .ZN(n9817)
         );
  OAI22_X1 U9199 ( .A1(n9817), .A2(n9317), .B1(n9655), .B2(n7503), .ZN(n7504)
         );
  OAI21_X1 U9200 ( .B1(n9819), .B2(n7504), .A(n9660), .ZN(n7508) );
  OAI22_X1 U9201 ( .A1(n9654), .A2(n9818), .B1(n6170), .B2(n9660), .ZN(n7506)
         );
  INV_X1 U9202 ( .A(n7506), .ZN(n7507) );
  OAI211_X1 U9203 ( .C1(n7509), .C2(n9373), .A(n7508), .B(n7507), .ZN(P1_U3286) );
  NAND2_X1 U9204 ( .A1(n6070), .A2(n9317), .ZN(n7659) );
  AOI21_X1 U9205 ( .B1(n9652), .B2(n7659), .A(n7510), .ZN(n7515) );
  NAND2_X1 U9206 ( .A1(n7511), .A2(n9331), .ZN(n7512) );
  OAI21_X1 U9207 ( .B1(n9655), .B2(n7513), .A(n7512), .ZN(n7514) );
  NOR3_X1 U9208 ( .A1(n7516), .A2(n7515), .A3(n7514), .ZN(n7518) );
  AOI22_X1 U9209 ( .A1(n9334), .A2(n6694), .B1(P1_REG2_REG_1__SCAN_IN), .B2(
        n9399), .ZN(n7517) );
  OAI21_X1 U9210 ( .B1(n7518), .B2(n9399), .A(n7517), .ZN(P1_U3290) );
  INV_X1 U9211 ( .A(n7519), .ZN(n7571) );
  AOI22_X1 U9212 ( .A1(n8578), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n8965), .ZN(n7520) );
  OAI21_X1 U9213 ( .B1(n7571), .B2(n8968), .A(n7520), .ZN(P2_U3340) );
  XNOR2_X1 U9214 ( .A(n7522), .B(n7521), .ZN(n7523) );
  XNOR2_X1 U9215 ( .A(n7524), .B(n7523), .ZN(n7525) );
  NAND2_X1 U9216 ( .A1(n7525), .A2(n9115), .ZN(n7529) );
  INV_X1 U9217 ( .A(n9134), .ZN(n7755) );
  OAI22_X1 U9218 ( .A1(n9118), .A2(n7683), .B1(n9117), .B2(n7755), .ZN(n7526)
         );
  AOI211_X1 U9219 ( .C1(n9120), .C2(n9136), .A(n7527), .B(n7526), .ZN(n7528)
         );
  OAI211_X1 U9220 ( .C1(n7682), .C2(n9123), .A(n7529), .B(n7528), .ZN(P1_U3237) );
  NAND2_X1 U9221 ( .A1(n6696), .A2(n9489), .ZN(n8282) );
  INV_X1 U9222 ( .A(n8282), .ZN(n7531) );
  OR2_X1 U9223 ( .A1(n7531), .A2(n7530), .ZN(n8344) );
  INV_X1 U9224 ( .A(n8431), .ZN(n7533) );
  INV_X1 U9225 ( .A(n9488), .ZN(n7532) );
  NOR2_X1 U9226 ( .A1(n7533), .A2(n7532), .ZN(n7534) );
  AOI22_X1 U9227 ( .A1(n8344), .A2(n7534), .B1(n9379), .B2(n9139), .ZN(n9487)
         );
  INV_X2 U9228 ( .A(n9660), .ZN(n9399) );
  INV_X1 U9229 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7535) );
  OAI22_X1 U9230 ( .A1(n9660), .A2(n6084), .B1(n7535), .B2(n9655), .ZN(n7536)
         );
  INV_X1 U9231 ( .A(n7536), .ZN(n7540) );
  OAI21_X1 U9232 ( .B1(n9640), .B2(n9334), .A(n7538), .ZN(n7539) );
  OAI211_X1 U9233 ( .C1(n9487), .C2(n9399), .A(n7540), .B(n7539), .ZN(P1_U3291) );
  OR2_X1 U9234 ( .A1(n7541), .A2(n8556), .ZN(n7542) );
  INV_X1 U9235 ( .A(n7596), .ZN(n7544) );
  AOI21_X1 U9236 ( .B1(n7546), .B2(n7545), .A(n7544), .ZN(n9989) );
  INV_X1 U9237 ( .A(n9933), .ZN(n7886) );
  XNOR2_X1 U9238 ( .A(n7547), .B(n7546), .ZN(n7550) );
  OAI22_X1 U9239 ( .A1(n7548), .A2(n8818), .B1(n7772), .B2(n8820), .ZN(n7549)
         );
  AOI21_X1 U9240 ( .B1(n7550), .B2(n8795), .A(n7549), .ZN(n7551) );
  OAI21_X1 U9241 ( .B1(n9989), .B2(n7877), .A(n7551), .ZN(n9992) );
  NAND2_X1 U9242 ( .A1(n9992), .A2(n8839), .ZN(n7557) );
  OAI22_X1 U9243 ( .A1(n8839), .A2(n7552), .B1(n7577), .B2(n8836), .ZN(n7555)
         );
  AND2_X1 U9244 ( .A1(n9929), .A2(n7594), .ZN(n7553) );
  NOR2_X1 U9245 ( .A1(n9929), .A2(n7594), .ZN(n7613) );
  OR2_X1 U9246 ( .A1(n7553), .A2(n7613), .ZN(n9991) );
  NOR2_X1 U9247 ( .A1(n9991), .A2(n8717), .ZN(n7554) );
  AOI211_X1 U9248 ( .C1(n9926), .C2(n7594), .A(n7555), .B(n7554), .ZN(n7556)
         );
  OAI211_X1 U9249 ( .C1(n9989), .C2(n7886), .A(n7557), .B(n7556), .ZN(P2_U3287) );
  OAI21_X1 U9250 ( .B1(n7559), .B2(n8155), .A(n7558), .ZN(n7620) );
  INV_X1 U9251 ( .A(n7620), .ZN(n7570) );
  INV_X1 U9252 ( .A(n7680), .ZN(n7561) );
  INV_X1 U9253 ( .A(n7759), .ZN(n7560) );
  AOI211_X1 U9254 ( .C1(n7625), .C2(n7561), .A(n9827), .B(n7560), .ZN(n7619)
         );
  NOR2_X1 U9255 ( .A1(n9654), .A2(n7622), .ZN(n7564) );
  OAI22_X1 U9256 ( .A1(n9660), .A2(n7562), .B1(n7588), .B2(n9655), .ZN(n7563)
         );
  AOI211_X1 U9257 ( .C1(n7619), .C2(n9395), .A(n7564), .B(n7563), .ZN(n7569)
         );
  XOR2_X1 U9258 ( .A(n8155), .B(n7565), .Z(n7566) );
  OAI222_X1 U9259 ( .A1(n9644), .A2(n7567), .B1(n9646), .B2(n7854), .C1(n9326), 
        .C2(n7566), .ZN(n7618) );
  NAND2_X1 U9260 ( .A1(n7618), .A2(n9660), .ZN(n7568) );
  OAI211_X1 U9261 ( .C1(n7570), .C2(n9373), .A(n7569), .B(n7568), .ZN(P1_U3284) );
  INV_X1 U9262 ( .A(n9797), .ZN(n9160) );
  INV_X1 U9263 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10401) );
  OAI222_X1 U9264 ( .A1(n9160), .A2(n4476), .B1(n8089), .B2(n7571), .C1(n10401), .C2(n9549), .ZN(P1_U3335) );
  OAI21_X1 U9265 ( .B1(n7574), .B2(n7482), .A(n7572), .ZN(n7582) );
  INV_X1 U9266 ( .A(n7594), .ZN(n9990) );
  NOR3_X1 U9267 ( .A1(n7574), .A2(n7573), .A3(n8505), .ZN(n7575) );
  OAI21_X1 U9268 ( .B1(n7575), .B2(n8517), .A(n8555), .ZN(n7580) );
  INV_X1 U9269 ( .A(n7772), .ZN(n8553) );
  OAI21_X1 U9270 ( .B1(n9616), .B2(n7577), .A(n7576), .ZN(n7578) );
  AOI21_X1 U9271 ( .B1(n8516), .B2(n8553), .A(n7578), .ZN(n7579) );
  OAI211_X1 U9272 ( .C1(n9990), .C2(n5785), .A(n7580), .B(n7579), .ZN(n7581)
         );
  AOI21_X1 U9273 ( .B1(n7582), .B2(n9611), .A(n7581), .ZN(n7583) );
  INV_X1 U9274 ( .A(n7583), .ZN(P2_U3233) );
  NAND2_X1 U9275 ( .A1(n7586), .A2(n7585), .ZN(n7587) );
  XNOR2_X1 U9276 ( .A(n7584), .B(n7587), .ZN(n7593) );
  OAI22_X1 U9277 ( .A1(n9118), .A2(n7588), .B1(n9117), .B2(n7854), .ZN(n7589)
         );
  AOI211_X1 U9278 ( .C1(n9120), .C2(n9135), .A(n7590), .B(n7589), .ZN(n7592)
         );
  NAND2_X1 U9279 ( .A1(n9095), .A2(n7625), .ZN(n7591) );
  OAI211_X1 U9280 ( .C1(n7593), .C2(n9097), .A(n7592), .B(n7591), .ZN(P1_U3211) );
  OR2_X1 U9281 ( .A1(n7594), .A2(n8554), .ZN(n7595) );
  NAND2_X1 U9282 ( .A1(n7596), .A2(n7595), .ZN(n7599) );
  INV_X1 U9283 ( .A(n7599), .ZN(n7597) );
  NAND2_X1 U9284 ( .A1(n7599), .A2(n7598), .ZN(n7600) );
  NAND2_X1 U9285 ( .A1(n7648), .A2(n7600), .ZN(n9996) );
  OAI22_X1 U9286 ( .A1(n7899), .A2(n8820), .B1(n7601), .B2(n8818), .ZN(n7602)
         );
  INV_X1 U9287 ( .A(n7602), .ZN(n7610) );
  NAND2_X1 U9288 ( .A1(n7604), .A2(n7603), .ZN(n7606) );
  NAND2_X1 U9289 ( .A1(n7606), .A2(n7605), .ZN(n7608) );
  NAND3_X1 U9290 ( .A1(n7608), .A2(n7607), .A3(n8795), .ZN(n7609) );
  OAI211_X1 U9291 ( .C1(n9996), .C2(n7877), .A(n7610), .B(n7609), .ZN(n9999)
         );
  NAND2_X1 U9292 ( .A1(n9999), .A2(n8839), .ZN(n7617) );
  OAI22_X1 U9293 ( .A1(n8839), .A2(n7611), .B1(n7822), .B2(n8836), .ZN(n7615)
         );
  INV_X1 U9294 ( .A(n7829), .ZN(n9997) );
  INV_X1 U9295 ( .A(n7732), .ZN(n7612) );
  OAI21_X1 U9296 ( .B1(n9997), .B2(n7613), .A(n7612), .ZN(n9998) );
  NOR2_X1 U9297 ( .A1(n9998), .A2(n8717), .ZN(n7614) );
  AOI211_X1 U9298 ( .C1(n9926), .C2(n7829), .A(n7615), .B(n7614), .ZN(n7616)
         );
  OAI211_X1 U9299 ( .C1(n9996), .C2(n7886), .A(n7617), .B(n7616), .ZN(P2_U3286) );
  AOI211_X1 U9300 ( .C1(n9822), .C2(n7620), .A(n7619), .B(n7618), .ZN(n7628)
         );
  INV_X1 U9301 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7621) );
  OAI22_X1 U9302 ( .A1(n9532), .A2(n7622), .B1(n9835), .B2(n7621), .ZN(n7623)
         );
  INV_X1 U9303 ( .A(n7623), .ZN(n7624) );
  OAI21_X1 U9304 ( .B1(n7628), .B2(n9833), .A(n7624), .ZN(P1_U3475) );
  AOI22_X1 U9305 ( .A1(n7626), .A2(n7625), .B1(n9838), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7627) );
  OAI21_X1 U9306 ( .B1(n7628), .B2(n9838), .A(n7627), .ZN(P1_U3530) );
  NAND2_X1 U9307 ( .A1(n7636), .A2(n7629), .ZN(n7631) );
  NAND2_X1 U9308 ( .A1(n7631), .A2(n7630), .ZN(n7633) );
  XNOR2_X1 U9309 ( .A(n7640), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n7632) );
  NOR2_X1 U9310 ( .A1(n7633), .A2(n7632), .ZN(n8563) );
  AOI21_X1 U9311 ( .B1(n7633), .B2(n7632), .A(n8563), .ZN(n7646) );
  INV_X1 U9312 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n10044) );
  NAND2_X1 U9313 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8059) );
  OAI21_X1 U9314 ( .B1(n9566), .B2(n10044), .A(n8059), .ZN(n7634) );
  AOI21_X1 U9315 ( .B1(n9905), .B2(n7640), .A(n7634), .ZN(n7645) );
  NOR2_X1 U9316 ( .A1(n7636), .A2(n7635), .ZN(n7638) );
  NOR2_X1 U9317 ( .A1(n7638), .A2(n7637), .ZN(n7643) );
  NAND2_X1 U9318 ( .A1(n7640), .A2(n8576), .ZN(n7639) );
  OAI21_X1 U9319 ( .B1(n7640), .B2(n8576), .A(n7639), .ZN(n7642) );
  NAND2_X1 U9320 ( .A1(n8575), .A2(n8576), .ZN(n7641) );
  OAI211_X1 U9321 ( .C1(n8576), .C2(n8575), .A(n7643), .B(n7641), .ZN(n8574)
         );
  OAI211_X1 U9322 ( .C1(n7643), .C2(n7642), .A(n8574), .B(n9901), .ZN(n7644)
         );
  OAI211_X1 U9323 ( .C1(n7646), .C2(n9843), .A(n7645), .B(n7644), .ZN(P2_U3261) );
  NAND2_X1 U9324 ( .A1(n7829), .A2(n8553), .ZN(n7647) );
  NAND2_X1 U9325 ( .A1(n7648), .A2(n7647), .ZN(n7649) );
  OAI21_X1 U9326 ( .B1(n7649), .B2(n7652), .A(n7728), .ZN(n10004) );
  NAND2_X1 U9327 ( .A1(n7607), .A2(n7650), .ZN(n7651) );
  XOR2_X1 U9328 ( .A(n7652), .B(n7651), .Z(n7653) );
  OAI222_X1 U9329 ( .A1(n8820), .A2(n7773), .B1(n8818), .B2(n7772), .C1(n9917), 
        .C2(n7653), .ZN(n10007) );
  NAND2_X1 U9330 ( .A1(n10007), .A2(n8839), .ZN(n7658) );
  OAI22_X1 U9331 ( .A1(n8839), .A2(n7654), .B1(n7771), .B2(n8836), .ZN(n7656)
         );
  INV_X1 U9332 ( .A(n7776), .ZN(n10005) );
  XNOR2_X1 U9333 ( .A(n7732), .B(n10005), .ZN(n10006) );
  NOR2_X1 U9334 ( .A1(n10006), .A2(n8717), .ZN(n7655) );
  AOI211_X1 U9335 ( .C1(n9926), .C2(n7776), .A(n7656), .B(n7655), .ZN(n7657)
         );
  OAI211_X1 U9336 ( .C1(n8843), .C2(n10004), .A(n7658), .B(n7657), .ZN(
        P2_U3285) );
  INV_X1 U9337 ( .A(n9640), .ZN(n7986) );
  INV_X1 U9338 ( .A(n9655), .ZN(n9343) );
  AOI22_X1 U9339 ( .A1(n9334), .A2(n7661), .B1(n7660), .B2(n9343), .ZN(n7662)
         );
  OAI21_X1 U9340 ( .B1(n7986), .B2(n7663), .A(n7662), .ZN(n7666) );
  MUX2_X1 U9341 ( .A(n7664), .B(P1_REG2_REG_4__SCAN_IN), .S(n9399), .Z(n7665)
         );
  AOI211_X1 U9342 ( .C1(n9641), .C2(n7667), .A(n7666), .B(n7665), .ZN(n7668)
         );
  INV_X1 U9343 ( .A(n7668), .ZN(P1_U3287) );
  INV_X1 U9344 ( .A(n7669), .ZN(n7670) );
  OAI222_X1 U9345 ( .A1(P1_U3084), .A2(n9331), .B1(n8089), .B2(n7670), .C1(
        n10375), .C2(n9549), .ZN(P1_U3334) );
  OAI222_X1 U9346 ( .A1(n8980), .A2(n7671), .B1(n8968), .B2(n7670), .C1(n8835), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OAI21_X1 U9347 ( .B1(n7673), .B2(n8154), .A(n7672), .ZN(n7783) );
  OAI22_X1 U9348 ( .A1(n7674), .A2(n9644), .B1(n7755), .B2(n9646), .ZN(n7679)
         );
  INV_X1 U9349 ( .A(n8146), .ZN(n8150) );
  NOR2_X1 U9350 ( .A1(n7675), .A2(n8150), .ZN(n7676) );
  XOR2_X1 U9351 ( .A(n8154), .B(n7676), .Z(n7677) );
  NOR2_X1 U9352 ( .A1(n7677), .A2(n9326), .ZN(n7678) );
  AOI211_X1 U9353 ( .C1(n7980), .C2(n7783), .A(n7679), .B(n7678), .ZN(n7787)
         );
  AOI21_X1 U9354 ( .B1(n7784), .B2(n7681), .A(n7680), .ZN(n7785) );
  NOR2_X1 U9355 ( .A1(n9654), .A2(n7682), .ZN(n7686) );
  OAI22_X1 U9356 ( .A1(n9660), .A2(n7684), .B1(n7683), .B2(n9655), .ZN(n7685)
         );
  AOI211_X1 U9357 ( .C1(n7785), .C2(n9640), .A(n7686), .B(n7685), .ZN(n7688)
         );
  NAND2_X1 U9358 ( .A1(n7783), .A2(n9641), .ZN(n7687) );
  OAI211_X1 U9359 ( .C1(n7787), .C2(n9399), .A(n7688), .B(n7687), .ZN(P1_U3285) );
  XNOR2_X1 U9360 ( .A(n8343), .B(n7689), .ZN(n7694) );
  OAI21_X1 U9361 ( .B1(n7691), .B2(n8343), .A(n7690), .ZN(n9815) );
  NAND2_X1 U9362 ( .A1(n9815), .A2(n7980), .ZN(n7693) );
  AOI22_X1 U9363 ( .A1(n9382), .A2(n9138), .B1(n9137), .B2(n9379), .ZN(n7692)
         );
  OAI211_X1 U9364 ( .C1(n9326), .C2(n7694), .A(n7693), .B(n7692), .ZN(n9813)
         );
  INV_X1 U9365 ( .A(n9813), .ZN(n7703) );
  OR2_X1 U9366 ( .A1(n7695), .A2(n9811), .ZN(n7696) );
  NAND2_X1 U9367 ( .A1(n7697), .A2(n7696), .ZN(n9812) );
  NOR2_X1 U9368 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(n9655), .ZN(n7699) );
  NOR2_X1 U9369 ( .A1(n9654), .A2(n9811), .ZN(n7698) );
  AOI211_X1 U9370 ( .C1(n9399), .C2(P1_REG2_REG_3__SCAN_IN), .A(n7699), .B(
        n7698), .ZN(n7700) );
  OAI21_X1 U9371 ( .B1(n7986), .B2(n9812), .A(n7700), .ZN(n7701) );
  AOI21_X1 U9372 ( .B1(n9641), .B2(n9815), .A(n7701), .ZN(n7702) );
  OAI21_X1 U9373 ( .B1(n7703), .B2(n9399), .A(n7702), .ZN(P1_U3288) );
  INV_X1 U9374 ( .A(n9734), .ZN(n7707) );
  NOR2_X1 U9375 ( .A1(n7714), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7704) );
  NOR2_X1 U9376 ( .A1(n7705), .A2(n7704), .ZN(n9737) );
  MUX2_X1 U9377 ( .A(n7706), .B(P1_REG1_REG_12__SCAN_IN), .S(n9734), .Z(n9736)
         );
  NOR2_X1 U9378 ( .A1(n9737), .A2(n9736), .ZN(n9735) );
  AOI21_X1 U9379 ( .B1(n7707), .B2(n7706), .A(n9735), .ZN(n9749) );
  MUX2_X1 U9380 ( .A(n7708), .B(P1_REG1_REG_13__SCAN_IN), .S(n9747), .Z(n9750)
         );
  NOR2_X1 U9381 ( .A1(n9749), .A2(n9750), .ZN(n9748) );
  AOI21_X1 U9382 ( .B1(n7708), .B2(n7709), .A(n9748), .ZN(n7711) );
  AOI22_X1 U9383 ( .A1(n7720), .A2(n6349), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n9152), .ZN(n7710) );
  NOR2_X1 U9384 ( .A1(n7711), .A2(n7710), .ZN(n9151) );
  AOI21_X1 U9385 ( .B1(n7711), .B2(n7710), .A(n9151), .ZN(n7726) );
  INV_X1 U9386 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7723) );
  NAND2_X1 U9387 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n9734), .ZN(n7712) );
  OAI21_X1 U9388 ( .B1(n9734), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7712), .ZN(
        n9730) );
  OAI21_X1 U9389 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7714), .A(n7713), .ZN(
        n9731) );
  NOR2_X1 U9390 ( .A1(n9730), .A2(n9731), .ZN(n9729) );
  MUX2_X1 U9391 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n7983), .S(n9747), .Z(n7715)
         );
  INV_X1 U9392 ( .A(n7715), .ZN(n9743) );
  XNOR2_X1 U9393 ( .A(n7720), .B(n7716), .ZN(n7717) );
  NOR2_X1 U9394 ( .A1(n8014), .A2(n7717), .ZN(n9141) );
  AOI21_X1 U9395 ( .B1(n7717), .B2(n8014), .A(n9141), .ZN(n7719) );
  NAND2_X1 U9396 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9001) );
  INV_X1 U9397 ( .A(n9001), .ZN(n7718) );
  AOI21_X1 U9398 ( .B1(n9720), .B2(n7719), .A(n7718), .ZN(n7722) );
  NAND2_X1 U9399 ( .A1(n9796), .A2(n7720), .ZN(n7721) );
  OAI211_X1 U9400 ( .C1(n9806), .C2(n7723), .A(n7722), .B(n7721), .ZN(n7724)
         );
  INV_X1 U9401 ( .A(n7724), .ZN(n7725) );
  OAI21_X1 U9402 ( .B1(n7726), .B2(n9802), .A(n7725), .ZN(P1_U3255) );
  INV_X1 U9403 ( .A(n7899), .ZN(n8552) );
  NAND2_X1 U9404 ( .A1(n7776), .A2(n8552), .ZN(n7727) );
  OAI21_X1 U9405 ( .B1(n4587), .B2(n7730), .A(n7867), .ZN(n10017) );
  INV_X1 U9406 ( .A(n10017), .ZN(n7738) );
  XOR2_X1 U9407 ( .A(n7730), .B(n7729), .Z(n7731) );
  OAI222_X1 U9408 ( .A1(n8820), .A2(n7918), .B1(n8818), .B2(n7899), .C1(n7731), 
        .C2(n9917), .ZN(n10015) );
  OAI21_X1 U9409 ( .B1(n4588), .B2(n10012), .A(n7880), .ZN(n10014) );
  OAI22_X1 U9410 ( .A1(n8839), .A2(n7733), .B1(n7905), .B2(n8836), .ZN(n7734)
         );
  AOI21_X1 U9411 ( .B1(n7909), .B2(n9926), .A(n7734), .ZN(n7735) );
  OAI21_X1 U9412 ( .B1(n10014), .B2(n8717), .A(n7735), .ZN(n7736) );
  AOI21_X1 U9413 ( .B1(n10015), .B2(n8839), .A(n7736), .ZN(n7737) );
  OAI21_X1 U9414 ( .B1(n7738), .B2(n8843), .A(n7737), .ZN(P2_U3284) );
  INV_X1 U9415 ( .A(n7739), .ZN(n7779) );
  OAI222_X1 U9416 ( .A1(n8968), .A2(n7779), .B1(P2_U3152), .B2(n7741), .C1(
        n7740), .C2(n8980), .ZN(P2_U3338) );
  AOI22_X1 U9417 ( .A1(n9399), .A2(P1_REG2_REG_2__SCAN_IN), .B1(n9343), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7742) );
  OAI21_X1 U9418 ( .B1(n8281), .B2(n9654), .A(n7742), .ZN(n7745) );
  INV_X1 U9419 ( .A(n9641), .ZN(n7866) );
  NOR2_X1 U9420 ( .A1(n7743), .A2(n7866), .ZN(n7744) );
  AOI211_X1 U9421 ( .C1(n7746), .C2(n9640), .A(n7745), .B(n7744), .ZN(n7747)
         );
  OAI21_X1 U9422 ( .B1(n9399), .B2(n7748), .A(n7747), .ZN(P1_U3289) );
  NAND2_X1 U9423 ( .A1(n7750), .A2(n8351), .ZN(n7751) );
  INV_X1 U9424 ( .A(n7852), .ZN(n7754) );
  AOI21_X1 U9425 ( .B1(n7752), .B2(n8275), .A(n8351), .ZN(n7753) );
  NOR3_X1 U9426 ( .A1(n7754), .A2(n7753), .A3(n9326), .ZN(n7757) );
  OAI22_X1 U9427 ( .A1(n7799), .A2(n9646), .B1(n7755), .B2(n9644), .ZN(n7756)
         );
  AOI211_X1 U9428 ( .C1(n7839), .C2(n7980), .A(n7757), .B(n7756), .ZN(n7843)
         );
  AOI21_X1 U9429 ( .B1(n7840), .B2(n7759), .A(n7758), .ZN(n7841) );
  NOR2_X1 U9430 ( .A1(n9654), .A2(n7804), .ZN(n7762) );
  OAI22_X1 U9431 ( .A1(n9660), .A2(n7760), .B1(n7800), .B2(n9655), .ZN(n7761)
         );
  AOI211_X1 U9432 ( .C1(n7841), .C2(n9640), .A(n7762), .B(n7761), .ZN(n7764)
         );
  NAND2_X1 U9433 ( .A1(n7839), .A2(n9641), .ZN(n7763) );
  OAI211_X1 U9434 ( .C1(n7843), .C2(n9399), .A(n7764), .B(n7763), .ZN(P1_U3283) );
  INV_X1 U9435 ( .A(n7765), .ZN(n7766) );
  AOI21_X1 U9436 ( .B1(n7823), .B2(n7766), .A(n8542), .ZN(n7770) );
  NOR3_X1 U9437 ( .A1(n7767), .A2(n7772), .A3(n8505), .ZN(n7769) );
  OAI21_X1 U9438 ( .B1(n7770), .B2(n7769), .A(n7768), .ZN(n7778) );
  OAI22_X1 U9439 ( .A1(n9616), .A2(n7771), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10356), .ZN(n7775) );
  OAI22_X1 U9440 ( .A1(n8527), .A2(n7773), .B1(n7772), .B2(n8526), .ZN(n7774)
         );
  AOI211_X1 U9441 ( .C1(n9610), .C2(n7776), .A(n7775), .B(n7774), .ZN(n7777)
         );
  NAND2_X1 U9442 ( .A1(n7778), .A2(n7777), .ZN(P2_U3238) );
  OAI222_X1 U9443 ( .A1(n8339), .A2(P1_U3084), .B1(n8089), .B2(n7779), .C1(
        n10419), .C2(n9549), .ZN(P1_U3333) );
  INV_X1 U9444 ( .A(n7780), .ZN(n8088) );
  OAI222_X1 U9445 ( .A1(n8983), .A2(n8088), .B1(P2_U3152), .B2(n7782), .C1(
        n7781), .C2(n8980), .ZN(P2_U3337) );
  INV_X1 U9446 ( .A(n7783), .ZN(n7788) );
  AOI22_X1 U9447 ( .A1(n7785), .A2(n9467), .B1(n9466), .B2(n7784), .ZN(n7786)
         );
  OAI211_X1 U9448 ( .C1(n7788), .C2(n7845), .A(n7787), .B(n7786), .ZN(n7790)
         );
  NAND2_X1 U9449 ( .A1(n7790), .A2(n9840), .ZN(n7789) );
  OAI21_X1 U9450 ( .B1(n9840), .B2(n6190), .A(n7789), .ZN(P1_U3529) );
  INV_X1 U9451 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7792) );
  NAND2_X1 U9452 ( .A1(n7790), .A2(n9835), .ZN(n7791) );
  OAI21_X1 U9453 ( .B1(n9835), .B2(n7792), .A(n7791), .ZN(P1_U3472) );
  NAND2_X1 U9454 ( .A1(n7793), .A2(n7794), .ZN(n7796) );
  XNOR2_X1 U9455 ( .A(n7796), .B(n7795), .ZN(n7797) );
  NAND2_X1 U9456 ( .A1(n7797), .A2(n9115), .ZN(n7803) );
  NOR2_X1 U9457 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7798), .ZN(n9716) );
  OAI22_X1 U9458 ( .A1(n9118), .A2(n7800), .B1(n9117), .B2(n7799), .ZN(n7801)
         );
  AOI211_X1 U9459 ( .C1(n9120), .C2(n9134), .A(n9716), .B(n7801), .ZN(n7802)
         );
  OAI211_X1 U9460 ( .C1(n7804), .C2(n9123), .A(n7803), .B(n7802), .ZN(P1_U3219) );
  XNOR2_X1 U9461 ( .A(n7805), .B(n7806), .ZN(n9593) );
  INV_X1 U9462 ( .A(n9593), .ZN(n7819) );
  INV_X1 U9463 ( .A(n7806), .ZN(n8353) );
  XNOR2_X1 U9464 ( .A(n7807), .B(n8353), .ZN(n7808) );
  NAND2_X1 U9465 ( .A1(n7808), .A2(n9649), .ZN(n7810) );
  AOI22_X1 U9466 ( .A1(n9379), .A2(n9130), .B1(n9132), .B2(n9382), .ZN(n7809)
         );
  NAND2_X1 U9467 ( .A1(n7810), .A2(n7809), .ZN(n9592) );
  INV_X1 U9468 ( .A(n7895), .ZN(n9590) );
  INV_X1 U9469 ( .A(n7861), .ZN(n7812) );
  INV_X1 U9470 ( .A(n9636), .ZN(n7811) );
  OAI211_X1 U9471 ( .C1(n9590), .C2(n7812), .A(n7811), .B(n9467), .ZN(n9589)
         );
  INV_X1 U9472 ( .A(n9395), .ZN(n7816) );
  OAI22_X1 U9473 ( .A1(n9660), .A2(n7813), .B1(n7892), .B2(n9655), .ZN(n7814)
         );
  AOI21_X1 U9474 ( .B1(n7895), .B2(n9334), .A(n7814), .ZN(n7815) );
  OAI21_X1 U9475 ( .B1(n9589), .B2(n7816), .A(n7815), .ZN(n7817) );
  AOI21_X1 U9476 ( .B1(n9592), .B2(n9660), .A(n7817), .ZN(n7818) );
  OAI21_X1 U9477 ( .B1(n7819), .B2(n9373), .A(n7818), .ZN(P1_U3281) );
  AOI22_X1 U9478 ( .A1(n8517), .A2(n8554), .B1(n8516), .B2(n8552), .ZN(n7821)
         );
  OAI211_X1 U9479 ( .C1(n7822), .C2(n9616), .A(n7821), .B(n7820), .ZN(n7828)
         );
  INV_X1 U9480 ( .A(n7823), .ZN(n7824) );
  AOI211_X1 U9481 ( .C1(n7826), .C2(n7825), .A(n8542), .B(n7824), .ZN(n7827)
         );
  AOI211_X1 U9482 ( .C1(n9610), .C2(n7829), .A(n7828), .B(n7827), .ZN(n7830)
         );
  INV_X1 U9483 ( .A(n7830), .ZN(P2_U3219) );
  AOI21_X1 U9484 ( .B1(n7832), .B2(n7831), .A(n4589), .ZN(n7838) );
  INV_X1 U9485 ( .A(n7833), .ZN(n7835) );
  OAI22_X1 U9486 ( .A1(n9118), .A2(n7858), .B1(n9117), .B2(n9645), .ZN(n7834)
         );
  AOI211_X1 U9487 ( .C1(n9120), .C2(n9133), .A(n7835), .B(n7834), .ZN(n7837)
         );
  NAND2_X1 U9488 ( .A1(n9825), .A2(n9095), .ZN(n7836) );
  OAI211_X1 U9489 ( .C1(n7838), .C2(n9097), .A(n7837), .B(n7836), .ZN(P1_U3229) );
  INV_X1 U9490 ( .A(n7839), .ZN(n7844) );
  AOI22_X1 U9491 ( .A1(n7841), .A2(n9467), .B1(n9466), .B2(n7840), .ZN(n7842)
         );
  OAI211_X1 U9492 ( .C1(n7845), .C2(n7844), .A(n7843), .B(n7842), .ZN(n7848)
         );
  NAND2_X1 U9493 ( .A1(n7848), .A2(n9840), .ZN(n7846) );
  OAI21_X1 U9494 ( .B1(n9840), .B2(n7847), .A(n7846), .ZN(P1_U3531) );
  INV_X1 U9495 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7850) );
  NAND2_X1 U9496 ( .A1(n7848), .A2(n9835), .ZN(n7849) );
  OAI21_X1 U9497 ( .B1(n9835), .B2(n7850), .A(n7849), .ZN(P1_U3478) );
  XOR2_X1 U9498 ( .A(n8352), .B(n7851), .Z(n9824) );
  NAND2_X1 U9499 ( .A1(n7852), .A2(n8164), .ZN(n7853) );
  XOR2_X1 U9500 ( .A(n8352), .B(n7853), .Z(n7856) );
  OAI22_X1 U9501 ( .A1(n9645), .A2(n9646), .B1(n7854), .B2(n9644), .ZN(n7855)
         );
  AOI21_X1 U9502 ( .B1(n7856), .B2(n9649), .A(n7855), .ZN(n7857) );
  OAI21_X1 U9503 ( .B1(n9824), .B2(n9652), .A(n7857), .ZN(n9829) );
  NAND2_X1 U9504 ( .A1(n9829), .A2(n9660), .ZN(n7865) );
  OAI22_X1 U9505 ( .A1(n9660), .A2(n7859), .B1(n7858), .B2(n9655), .ZN(n7863)
         );
  NAND2_X1 U9506 ( .A1(n4759), .A2(n9825), .ZN(n7860) );
  NAND2_X1 U9507 ( .A1(n7861), .A2(n7860), .ZN(n9828) );
  NOR2_X1 U9508 ( .A1(n9828), .A2(n7986), .ZN(n7862) );
  AOI211_X1 U9509 ( .C1(n9334), .C2(n9825), .A(n7863), .B(n7862), .ZN(n7864)
         );
  OAI211_X1 U9510 ( .C1(n9824), .C2(n7866), .A(n7865), .B(n7864), .ZN(P1_U3282) );
  INV_X1 U9511 ( .A(n7869), .ZN(n7868) );
  NAND2_X1 U9512 ( .A1(n7868), .A2(n4670), .ZN(n7923) );
  NAND2_X1 U9513 ( .A1(n7869), .A2(n7871), .ZN(n7870) );
  NAND2_X1 U9514 ( .A1(n7923), .A2(n7870), .ZN(n8940) );
  XNOR2_X1 U9515 ( .A(n7872), .B(n7871), .ZN(n7875) );
  NAND2_X1 U9516 ( .A1(n8551), .A2(n8750), .ZN(n7873) );
  OAI21_X1 U9517 ( .B1(n7950), .B2(n8820), .A(n7873), .ZN(n7874) );
  AOI21_X1 U9518 ( .B1(n7875), .B2(n8795), .A(n7874), .ZN(n7876) );
  OAI21_X1 U9519 ( .B1(n8940), .B2(n7877), .A(n7876), .ZN(n8942) );
  NAND2_X1 U9520 ( .A1(n8942), .A2(n8839), .ZN(n7885) );
  OAI22_X1 U9521 ( .A1(n8839), .A2(n7879), .B1(n7878), .B2(n8836), .ZN(n7883)
         );
  AND2_X1 U9522 ( .A1(n7880), .A2(n7921), .ZN(n7881) );
  OR2_X1 U9523 ( .A1(n7881), .A2(n4571), .ZN(n8936) );
  NOR2_X1 U9524 ( .A1(n8936), .A2(n8717), .ZN(n7882) );
  AOI211_X1 U9525 ( .C1(n9926), .C2(n7921), .A(n7883), .B(n7882), .ZN(n7884)
         );
  OAI211_X1 U9526 ( .C1(n8940), .C2(n7886), .A(n7885), .B(n7884), .ZN(P2_U3283) );
  XNOR2_X1 U9527 ( .A(n7888), .B(n7887), .ZN(n7889) );
  XNOR2_X1 U9528 ( .A(n7890), .B(n7889), .ZN(n7898) );
  OAI22_X1 U9529 ( .A1(n9118), .A2(n7892), .B1(n9117), .B2(n7891), .ZN(n7893)
         );
  AOI211_X1 U9530 ( .C1(n9120), .C2(n9132), .A(n7894), .B(n7893), .ZN(n7897)
         );
  NAND2_X1 U9531 ( .A1(n7895), .A2(n9095), .ZN(n7896) );
  OAI211_X1 U9532 ( .C1(n7898), .C2(n9097), .A(n7897), .B(n7896), .ZN(P1_U3215) );
  INV_X1 U9533 ( .A(n7768), .ZN(n7902) );
  NOR3_X1 U9534 ( .A1(n7900), .A2(n7899), .A3(n8505), .ZN(n7901) );
  AOI21_X1 U9535 ( .B1(n7902), .B2(n9611), .A(n7901), .ZN(n7912) );
  INV_X1 U9536 ( .A(n7918), .ZN(n8550) );
  AOI22_X1 U9537 ( .A1(n8517), .A2(n8552), .B1(n8516), .B2(n8550), .ZN(n7904)
         );
  OAI211_X1 U9538 ( .C1(n7905), .C2(n9616), .A(n7904), .B(n7903), .ZN(n7908)
         );
  NOR2_X1 U9539 ( .A1(n7906), .A2(n8542), .ZN(n7907) );
  AOI211_X1 U9540 ( .C1(n9610), .C2(n7909), .A(n7908), .B(n7907), .ZN(n7910)
         );
  OAI21_X1 U9541 ( .B1(n7912), .B2(n7911), .A(n7910), .ZN(P2_U3226) );
  INV_X1 U9542 ( .A(n7913), .ZN(n7916) );
  OAI222_X1 U9543 ( .A1(n4476), .A2(n7915), .B1(n8089), .B2(n7916), .C1(n7914), 
        .C2(n9549), .ZN(P1_U3331) );
  OAI222_X1 U9544 ( .A1(P2_U3152), .A2(n5782), .B1(n8968), .B2(n7916), .C1(
        n8980), .C2(n5657), .ZN(P2_U3336) );
  AOI21_X1 U9545 ( .B1(n4509), .B2(n7924), .A(n9917), .ZN(n7920) );
  OAI22_X1 U9546 ( .A1(n8061), .A2(n8820), .B1(n7918), .B2(n8818), .ZN(n9596)
         );
  AOI21_X1 U9547 ( .B1(n7920), .B2(n7919), .A(n9596), .ZN(n8933) );
  NAND2_X1 U9548 ( .A1(n7921), .A2(n8550), .ZN(n7922) );
  OAI21_X1 U9549 ( .B1(n7925), .B2(n7924), .A(n7940), .ZN(n8929) );
  NAND2_X1 U9550 ( .A1(n8929), .A2(n8736), .ZN(n7930) );
  XNOR2_X1 U9551 ( .A(n4571), .B(n9600), .ZN(n8931) );
  OAI22_X1 U9552 ( .A1(n8839), .A2(n7926), .B1(n9604), .B2(n8836), .ZN(n7928)
         );
  INV_X1 U9553 ( .A(n9600), .ZN(n7942) );
  NOR2_X1 U9554 ( .A1(n7942), .A2(n8813), .ZN(n7927) );
  AOI211_X1 U9555 ( .C1(n8931), .C2(n9932), .A(n7928), .B(n7927), .ZN(n7929)
         );
  OAI211_X1 U9556 ( .C1(n9936), .C2(n8933), .A(n7930), .B(n7929), .ZN(P2_U3282) );
  XNOR2_X1 U9557 ( .A(n7932), .B(n7931), .ZN(n7938) );
  OAI22_X1 U9558 ( .A1(n9105), .A2(n9645), .B1(n9118), .B2(n9656), .ZN(n7933)
         );
  AOI211_X1 U9559 ( .C1(n9108), .C2(n9129), .A(n7934), .B(n7933), .ZN(n7937)
         );
  NAND2_X1 U9560 ( .A1(n7935), .A2(n9095), .ZN(n7936) );
  OAI211_X1 U9561 ( .C1(n7938), .C2(n9097), .A(n7937), .B(n7936), .ZN(P1_U3234) );
  OR2_X1 U9562 ( .A1(n9600), .A2(n8549), .ZN(n7939) );
  XNOR2_X1 U9563 ( .A(n8021), .B(n7941), .ZN(n8928) );
  OR2_X1 U9564 ( .A1(n9609), .A2(n7944), .ZN(n8030) );
  INV_X1 U9565 ( .A(n8030), .ZN(n7943) );
  AOI21_X1 U9566 ( .B1(n9609), .B2(n7944), .A(n7943), .ZN(n8925) );
  INV_X1 U9567 ( .A(n9609), .ZN(n7947) );
  INV_X1 U9568 ( .A(n9615), .ZN(n7945) );
  AOI22_X1 U9569 ( .A1(n9936), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n7945), .B2(
        n9925), .ZN(n7946) );
  OAI21_X1 U9570 ( .B1(n7947), .B2(n8813), .A(n7946), .ZN(n7954) );
  INV_X1 U9571 ( .A(n7948), .ZN(n7949) );
  AOI21_X1 U9572 ( .B1(n7949), .B2(n8020), .A(n9917), .ZN(n7952) );
  OAI22_X1 U9573 ( .A1(n8607), .A2(n8820), .B1(n7950), .B2(n8818), .ZN(n9605)
         );
  AOI21_X1 U9574 ( .B1(n7952), .B2(n7951), .A(n9605), .ZN(n8927) );
  NOR2_X1 U9575 ( .A1(n8927), .A2(n9936), .ZN(n7953) );
  AOI211_X1 U9576 ( .C1(n8925), .C2(n9932), .A(n7954), .B(n7953), .ZN(n7955)
         );
  OAI21_X1 U9577 ( .B1(n8928), .B2(n8843), .A(n7955), .ZN(P2_U3281) );
  NAND2_X1 U9578 ( .A1(n7958), .A2(n9545), .ZN(n7957) );
  NAND2_X1 U9579 ( .A1(n7956), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8436) );
  OAI211_X1 U9580 ( .C1(n10402), .C2(n9544), .A(n7957), .B(n8436), .ZN(
        P1_U3330) );
  NAND2_X1 U9581 ( .A1(n7958), .A2(n8972), .ZN(n7960) );
  OAI211_X1 U9582 ( .C1(n7961), .C2(n8980), .A(n7960), .B(n7959), .ZN(P2_U3335) );
  NAND2_X1 U9583 ( .A1(n7962), .A2(n8356), .ZN(n7963) );
  XNOR2_X1 U9584 ( .A(n7963), .B(n8357), .ZN(n7964) );
  NAND2_X1 U9585 ( .A1(n7964), .A2(n9649), .ZN(n7966) );
  AOI22_X1 U9586 ( .A1(n9382), .A2(n9130), .B1(n9128), .B2(n9379), .ZN(n7965)
         );
  NAND2_X1 U9587 ( .A1(n7966), .A2(n7965), .ZN(n9482) );
  INV_X1 U9588 ( .A(n9482), .ZN(n7974) );
  NOR2_X1 U9589 ( .A1(n9399), .A2(n9652), .ZN(n7968) );
  XOR2_X1 U9590 ( .A(n7967), .B(n8357), .Z(n9484) );
  OAI21_X1 U9591 ( .B1(n9641), .B2(n7968), .A(n9484), .ZN(n7973) );
  AOI211_X1 U9592 ( .C1(n7999), .C2(n9638), .A(n9827), .B(n4773), .ZN(n9483)
         );
  INV_X1 U9593 ( .A(n7999), .ZN(n9533) );
  NOR2_X1 U9594 ( .A1(n9533), .A2(n9654), .ZN(n7971) );
  OAI22_X1 U9595 ( .A1(n9660), .A2(n7969), .B1(n7997), .B2(n9655), .ZN(n7970)
         );
  AOI211_X1 U9596 ( .C1(n9483), .C2(n9395), .A(n7971), .B(n7970), .ZN(n7972)
         );
  OAI211_X1 U9597 ( .C1(n9399), .C2(n7974), .A(n7973), .B(n7972), .ZN(P1_U3279) );
  XNOR2_X1 U9598 ( .A(n7975), .B(n8361), .ZN(n9670) );
  XNOR2_X1 U9599 ( .A(n7976), .B(n4803), .ZN(n7978) );
  AOI22_X1 U9600 ( .A1(n9382), .A2(n9129), .B1(n9127), .B2(n9379), .ZN(n7977)
         );
  OAI21_X1 U9601 ( .B1(n7978), .B2(n9326), .A(n7977), .ZN(n7979) );
  AOI21_X1 U9602 ( .B1(n9670), .B2(n7980), .A(n7979), .ZN(n9672) );
  AND2_X1 U9603 ( .A1(n7981), .A2(n8167), .ZN(n7982) );
  OR2_X1 U9604 ( .A1(n7982), .A2(n8012), .ZN(n9668) );
  OAI22_X1 U9605 ( .A1(n9660), .A2(n7983), .B1(n8040), .B2(n9655), .ZN(n7984)
         );
  AOI21_X1 U9606 ( .B1(n8167), .B2(n9334), .A(n7984), .ZN(n7985) );
  OAI21_X1 U9607 ( .B1(n9668), .B2(n7986), .A(n7985), .ZN(n7987) );
  AOI21_X1 U9608 ( .B1(n9670), .B2(n9641), .A(n7987), .ZN(n7988) );
  OAI21_X1 U9609 ( .B1(n9672), .B2(n9399), .A(n7988), .ZN(P1_U3278) );
  INV_X1 U9610 ( .A(n7989), .ZN(n8004) );
  OAI222_X1 U9611 ( .A1(n8983), .A2(n8004), .B1(P2_U3152), .B2(n7991), .C1(
        n7990), .C2(n8980), .ZN(P2_U3334) );
  INV_X1 U9612 ( .A(n7993), .ZN(n7994) );
  AOI21_X1 U9613 ( .B1(n7995), .B2(n7992), .A(n7994), .ZN(n8002) );
  NOR2_X1 U9614 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7996), .ZN(n9733) );
  OAI22_X1 U9615 ( .A1(n9118), .A2(n7997), .B1(n9117), .B2(n9002), .ZN(n7998)
         );
  AOI211_X1 U9616 ( .C1(n9120), .C2(n9130), .A(n9733), .B(n7998), .ZN(n8001)
         );
  NAND2_X1 U9617 ( .A1(n7999), .A2(n9095), .ZN(n8000) );
  OAI211_X1 U9618 ( .C1(n8002), .C2(n9097), .A(n8001), .B(n8000), .ZN(P1_U3222) );
  OAI222_X1 U9619 ( .A1(n8005), .A2(n4476), .B1(n8089), .B2(n8004), .C1(n8003), 
        .C2(n9549), .ZN(P1_U3329) );
  NAND2_X1 U9620 ( .A1(n8006), .A2(n8360), .ZN(n8007) );
  NAND3_X1 U9621 ( .A1(n8008), .A2(n9649), .A3(n8007), .ZN(n8010) );
  AOI22_X1 U9622 ( .A1(n9382), .A2(n9128), .B1(n9381), .B2(n9379), .ZN(n8009)
         );
  NAND2_X1 U9623 ( .A1(n8010), .A2(n8009), .ZN(n9478) );
  INV_X1 U9624 ( .A(n9478), .ZN(n8019) );
  XNOR2_X1 U9625 ( .A(n8011), .B(n8360), .ZN(n9480) );
  INV_X1 U9626 ( .A(n9373), .ZN(n9387) );
  NAND2_X1 U9627 ( .A1(n9480), .A2(n9387), .ZN(n8018) );
  INV_X1 U9628 ( .A(n8012), .ZN(n8013) );
  AOI211_X1 U9629 ( .C1(n9007), .C2(n8013), .A(n9827), .B(n9619), .ZN(n9479)
         );
  NOR2_X1 U9630 ( .A1(n9528), .A2(n9654), .ZN(n8016) );
  OAI22_X1 U9631 ( .A1(n9660), .A2(n8014), .B1(n9004), .B2(n9655), .ZN(n8015)
         );
  AOI211_X1 U9632 ( .C1(n9479), .C2(n9395), .A(n8016), .B(n8015), .ZN(n8017)
         );
  OAI211_X1 U9633 ( .C1(n9399), .C2(n8019), .A(n8018), .B(n8017), .ZN(P1_U3277) );
  INV_X1 U9634 ( .A(n8061), .ZN(n8548) );
  NAND2_X1 U9635 ( .A1(n8022), .A2(n8026), .ZN(n8608) );
  OR2_X1 U9636 ( .A1(n8022), .A2(n8026), .ZN(n8023) );
  AOI21_X1 U9637 ( .B1(n8026), .B2(n8025), .A(n8024), .ZN(n8028) );
  AOI22_X1 U9638 ( .A1(n8548), .A2(n8750), .B1(n8546), .B2(n8751), .ZN(n8027)
         );
  OAI21_X1 U9639 ( .B1(n8028), .B2(n9917), .A(n8027), .ZN(n8029) );
  AOI21_X1 U9640 ( .B1(n8918), .B2(n9922), .A(n8029), .ZN(n8923) );
  AND2_X1 U9641 ( .A1(n8064), .A2(n8030), .ZN(n8031) );
  OR2_X1 U9642 ( .A1(n8831), .A2(n8031), .ZN(n8920) );
  OAI22_X1 U9643 ( .A1(n8839), .A2(n8576), .B1(n8060), .B2(n8836), .ZN(n8032)
         );
  AOI21_X1 U9644 ( .B1(n8064), .B2(n9926), .A(n8032), .ZN(n8033) );
  OAI21_X1 U9645 ( .B1(n8920), .B2(n8717), .A(n8033), .ZN(n8034) );
  AOI21_X1 U9646 ( .B1(n8918), .B2(n9933), .A(n8034), .ZN(n8035) );
  OAI21_X1 U9647 ( .B1(n8923), .B2(n9936), .A(n8035), .ZN(P2_U3280) );
  NOR2_X1 U9648 ( .A1(n4514), .A2(n8036), .ZN(n8037) );
  XNOR2_X1 U9649 ( .A(n8038), .B(n8037), .ZN(n8039) );
  NAND2_X1 U9650 ( .A1(n8039), .A2(n9115), .ZN(n8043) );
  AND2_X1 U9651 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9746) );
  OAI22_X1 U9652 ( .A1(n9118), .A2(n8040), .B1(n9117), .B2(n9624), .ZN(n8041)
         );
  AOI211_X1 U9653 ( .C1(n9120), .C2(n9129), .A(n9746), .B(n8041), .ZN(n8042)
         );
  OAI211_X1 U9654 ( .C1(n4777), .C2(n9123), .A(n8043), .B(n8042), .ZN(P1_U3232) );
  INV_X1 U9655 ( .A(n8914), .ZN(n8609) );
  AOI21_X1 U9656 ( .B1(n8045), .B2(n8044), .A(n8542), .ZN(n8046) );
  NAND2_X1 U9657 ( .A1(n8046), .A2(n8074), .ZN(n8051) );
  INV_X1 U9658 ( .A(n8837), .ZN(n8049) );
  INV_X1 U9659 ( .A(n8610), .ZN(n8611) );
  NOR2_X1 U9660 ( .A1(n8607), .A2(n8818), .ZN(n8047) );
  AOI21_X1 U9661 ( .B1(n8611), .B2(n8751), .A(n8047), .ZN(n8829) );
  NAND2_X1 U9662 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9897) );
  OAI21_X1 U9663 ( .B1(n8829), .B2(n8481), .A(n9897), .ZN(n8048) );
  AOI21_X1 U9664 ( .B1(n8049), .B2(n8479), .A(n8048), .ZN(n8050) );
  OAI211_X1 U9665 ( .C1(n8609), .C2(n5785), .A(n8051), .B(n8050), .ZN(P2_U3230) );
  XNOR2_X1 U9666 ( .A(n8053), .B(n8052), .ZN(n9608) );
  AOI22_X1 U9667 ( .A1(n9608), .A2(n9607), .B1(n8054), .B2(n8053), .ZN(n8058)
         );
  XNOR2_X1 U9668 ( .A(n8056), .B(n8055), .ZN(n8057) );
  XNOR2_X1 U9669 ( .A(n8058), .B(n8057), .ZN(n8066) );
  OAI21_X1 U9670 ( .B1(n9616), .B2(n8060), .A(n8059), .ZN(n8063) );
  OAI22_X1 U9671 ( .A1(n8527), .A2(n8819), .B1(n8061), .B2(n8526), .ZN(n8062)
         );
  AOI211_X1 U9672 ( .C1(n8064), .C2(n9610), .A(n8063), .B(n8062), .ZN(n8065)
         );
  OAI21_X1 U9673 ( .B1(n8066), .B2(n8542), .A(n8065), .ZN(P2_U3228) );
  INV_X1 U9674 ( .A(n8067), .ZN(n8071) );
  OAI222_X1 U9675 ( .A1(n4476), .A2(n8069), .B1(n8089), .B2(n8071), .C1(n8068), 
        .C2(n9544), .ZN(P1_U3328) );
  OAI222_X1 U9676 ( .A1(n8980), .A2(n8072), .B1(n8968), .B2(n8071), .C1(n8070), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  AOI21_X1 U9677 ( .B1(n8074), .B2(n5023), .A(n8542), .ZN(n8077) );
  NOR3_X1 U9678 ( .A1(n8075), .A2(n8819), .A3(n8505), .ZN(n8076) );
  OAI21_X1 U9679 ( .B1(n8077), .B2(n8076), .A(n8120), .ZN(n8081) );
  OAI22_X1 U9680 ( .A1(n9616), .A2(n8810), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10427), .ZN(n8079) );
  OAI22_X1 U9681 ( .A1(n8527), .A2(n8821), .B1(n8819), .B2(n8526), .ZN(n8078)
         );
  AOI211_X1 U9682 ( .C1(n8909), .C2(n9610), .A(n8079), .B(n8078), .ZN(n8080)
         );
  NAND2_X1 U9683 ( .A1(n8081), .A2(n8080), .ZN(P2_U3240) );
  INV_X1 U9684 ( .A(n8082), .ZN(n8971) );
  OAI222_X1 U9685 ( .A1(n8089), .A2(n8971), .B1(n8084), .B2(P1_U3084), .C1(
        n8083), .C2(n9544), .ZN(P1_U3324) );
  INV_X1 U9686 ( .A(n8133), .ZN(n9543) );
  OAI222_X1 U9687 ( .A1(n8980), .A2(n8086), .B1(n8968), .B2(n9543), .C1(n8085), 
        .C2(P2_U3152), .ZN(P2_U3328) );
  OAI222_X1 U9688 ( .A1(n6657), .A2(P1_U3084), .B1(n8089), .B2(n8088), .C1(
        n8087), .C2(n9549), .ZN(P1_U3332) );
  OAI21_X1 U9689 ( .B1(n8091), .B2(n8097), .A(n8090), .ZN(n9464) );
  INV_X1 U9690 ( .A(n9360), .ZN(n8092) );
  AOI211_X1 U9691 ( .C1(n9462), .C2(n8092), .A(n9827), .B(n9339), .ZN(n9461)
         );
  NOR2_X1 U9692 ( .A1(n8093), .A2(n9654), .ZN(n8095) );
  OAI22_X1 U9693 ( .A1(n9660), .A2(n9147), .B1(n9091), .B2(n9655), .ZN(n8094)
         );
  AOI211_X1 U9694 ( .C1(n9461), .C2(n9395), .A(n8095), .B(n8094), .ZN(n8101)
         );
  NAND2_X1 U9695 ( .A1(n8096), .A2(n8198), .ZN(n8098) );
  INV_X1 U9696 ( .A(n8097), .ZN(n8365) );
  XNOR2_X1 U9697 ( .A(n8098), .B(n8365), .ZN(n8099) );
  OAI222_X1 U9698 ( .A1(n9646), .A2(n9328), .B1(n9644), .B2(n9092), .C1(n9326), 
        .C2(n8099), .ZN(n9460) );
  NAND2_X1 U9699 ( .A1(n9460), .A2(n9660), .ZN(n8100) );
  OAI211_X1 U9700 ( .C1(n9464), .C2(n9373), .A(n8101), .B(n8100), .ZN(P1_U3273) );
  INV_X1 U9701 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n8114) );
  AOI21_X1 U9702 ( .B1(n8104), .B2(n8103), .A(n8102), .ZN(n8108) );
  AOI21_X1 U9703 ( .B1(n8106), .B2(n8105), .A(n9702), .ZN(n8107) );
  OAI22_X1 U9704 ( .A1(n9802), .A2(n8108), .B1(n8107), .B2(n9790), .ZN(n8109)
         );
  AOI211_X1 U9705 ( .C1(n9796), .C2(n8111), .A(n8110), .B(n8109), .ZN(n8112)
         );
  OAI211_X1 U9706 ( .C1(n9806), .C2(n8114), .A(n8113), .B(n8112), .ZN(P1_U3245) );
  NAND2_X1 U9707 ( .A1(n6615), .A2(n9545), .ZN(n8116) );
  OAI211_X1 U9708 ( .C1(n9544), .C2(n8117), .A(n8116), .B(n8115), .ZN(P1_U3325) );
  INV_X1 U9709 ( .A(n8505), .ZN(n8521) );
  NAND3_X1 U9710 ( .A1(n8118), .A2(n8521), .A3(n8611), .ZN(n8119) );
  OAI21_X1 U9711 ( .B1(n8120), .B2(n8542), .A(n8119), .ZN(n8126) );
  INV_X1 U9712 ( .A(n8121), .ZN(n8125) );
  INV_X1 U9713 ( .A(n8906), .ZN(n8802) );
  OAI22_X1 U9714 ( .A1(n8762), .A2(n8820), .B1(n8610), .B2(n8818), .ZN(n8794)
         );
  AOI22_X1 U9715 ( .A1(n8794), .A2(n9606), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3152), .ZN(n8123) );
  NAND2_X1 U9716 ( .A1(n8479), .A2(n8800), .ZN(n8122) );
  OAI211_X1 U9717 ( .C1(n8802), .C2(n5785), .A(n8123), .B(n8122), .ZN(n8124)
         );
  AOI21_X1 U9718 ( .B1(n8126), .B2(n8125), .A(n8124), .ZN(n8127) );
  OAI21_X1 U9719 ( .B1(n8128), .B2(n8542), .A(n8127), .ZN(P2_U3221) );
  NAND2_X1 U9720 ( .A1(n8133), .A2(n6244), .ZN(n8136) );
  INV_X1 U9721 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10089) );
  OR2_X1 U9722 ( .A1(n8134), .A2(n10089), .ZN(n8135) );
  INV_X1 U9723 ( .A(n9124), .ZN(n8335) );
  NAND2_X1 U9724 ( .A1(n8372), .A2(n9175), .ZN(n8137) );
  INV_X1 U9725 ( .A(n8267), .ZN(n8262) );
  INV_X1 U9726 ( .A(n8139), .ZN(n8199) );
  AND2_X1 U9727 ( .A1(n9349), .A2(n8199), .ZN(n8274) );
  MUX2_X1 U9728 ( .A(n8274), .B(n8315), .S(n8267), .Z(n8205) );
  NAND2_X1 U9729 ( .A1(n8306), .A2(n8302), .ZN(n8141) );
  INV_X1 U9730 ( .A(n8305), .ZN(n8140) );
  MUX2_X1 U9731 ( .A(n8141), .B(n8140), .S(n8267), .Z(n8203) );
  INV_X1 U9732 ( .A(n8142), .ZN(n8144) );
  AOI21_X1 U9733 ( .B1(n8145), .B2(n8144), .A(n8143), .ZN(n8153) );
  INV_X1 U9734 ( .A(n8379), .ZN(n8147) );
  NAND2_X1 U9735 ( .A1(n8147), .A2(n8146), .ZN(n8149) );
  AND2_X1 U9736 ( .A1(n8149), .A2(n8148), .ZN(n8388) );
  OAI21_X1 U9737 ( .B1(n8151), .B2(n8150), .A(n8388), .ZN(n8152) );
  MUX2_X1 U9738 ( .A(n8153), .B(n8152), .S(n8262), .Z(n8156) );
  NOR2_X1 U9739 ( .A1(n8155), .A2(n8154), .ZN(n8349) );
  NAND2_X1 U9740 ( .A1(n8156), .A2(n8349), .ZN(n8163) );
  NAND2_X1 U9741 ( .A1(n8380), .A2(n8157), .ZN(n8384) );
  NAND2_X1 U9742 ( .A1(n8384), .A2(n8275), .ZN(n8161) );
  NAND2_X1 U9743 ( .A1(n8275), .A2(n8158), .ZN(n8159) );
  NAND2_X1 U9744 ( .A1(n8159), .A2(n8380), .ZN(n8160) );
  MUX2_X1 U9745 ( .A(n8161), .B(n8160), .S(n8267), .Z(n8162) );
  NAND2_X1 U9746 ( .A1(n8163), .A2(n8162), .ZN(n8179) );
  INV_X1 U9747 ( .A(n8276), .ZN(n8165) );
  OAI21_X1 U9748 ( .B1(n8179), .B2(n8165), .A(n8164), .ZN(n8166) );
  NAND2_X1 U9749 ( .A1(n8166), .A2(n8178), .ZN(n8171) );
  OR2_X1 U9750 ( .A1(n8167), .A2(n9002), .ZN(n8168) );
  AND2_X1 U9751 ( .A1(n8173), .A2(n8168), .ZN(n8193) );
  AND4_X1 U9752 ( .A1(n8297), .A2(n8267), .A3(n8169), .A4(n8292), .ZN(n8170)
         );
  NAND3_X1 U9753 ( .A1(n8171), .A2(n8193), .A3(n8170), .ZN(n8197) );
  INV_X1 U9754 ( .A(n8299), .ZN(n8174) );
  NAND2_X1 U9755 ( .A1(n8174), .A2(n8173), .ZN(n8177) );
  INV_X1 U9756 ( .A(n8193), .ZN(n8176) );
  NAND2_X1 U9757 ( .A1(n8176), .A2(n8175), .ZN(n8300) );
  AND2_X1 U9758 ( .A1(n8185), .A2(n8178), .ZN(n8180) );
  NAND3_X1 U9759 ( .A1(n8179), .A2(n8180), .A3(n8276), .ZN(n8184) );
  NAND2_X1 U9760 ( .A1(n8187), .A2(n8262), .ZN(n8190) );
  INV_X1 U9761 ( .A(n8180), .ZN(n8278) );
  OR2_X1 U9762 ( .A1(n8181), .A2(n8278), .ZN(n8293) );
  NAND3_X1 U9763 ( .A1(n8293), .A2(n8292), .A3(n8356), .ZN(n8182) );
  NOR2_X1 U9764 ( .A1(n8190), .A2(n8182), .ZN(n8183) );
  NAND2_X1 U9765 ( .A1(n8184), .A2(n8183), .ZN(n8194) );
  AND2_X1 U9766 ( .A1(n8290), .A2(n8355), .ZN(n8291) );
  NAND2_X1 U9767 ( .A1(n8355), .A2(n8185), .ZN(n8186) );
  NAND3_X1 U9768 ( .A1(n8187), .A2(n8356), .A3(n8186), .ZN(n8188) );
  NAND3_X1 U9769 ( .A1(n8188), .A2(n8267), .A3(n8290), .ZN(n8189) );
  OAI21_X1 U9770 ( .B1(n8291), .B2(n8190), .A(n8189), .ZN(n8191) );
  INV_X1 U9771 ( .A(n8191), .ZN(n8192) );
  NAND4_X1 U9772 ( .A1(n8194), .A2(n8193), .A3(n8299), .A4(n8192), .ZN(n8195)
         );
  AND4_X1 U9773 ( .A1(n8197), .A2(n9622), .A3(n8196), .A4(n8195), .ZN(n8202)
         );
  MUX2_X1 U9774 ( .A(n8200), .B(n8306), .S(n8267), .Z(n8201) );
  OAI211_X1 U9775 ( .C1(n8203), .C2(n8202), .A(n9364), .B(n8201), .ZN(n8204)
         );
  NAND2_X1 U9776 ( .A1(n8205), .A2(n8204), .ZN(n8209) );
  NAND3_X1 U9777 ( .A1(n8209), .A2(n8208), .A3(n8206), .ZN(n8207) );
  NAND3_X1 U9778 ( .A1(n8207), .A2(n8218), .A3(n8272), .ZN(n8212) );
  AND2_X1 U9779 ( .A1(n8213), .A2(n8208), .ZN(n8312) );
  AND2_X1 U9780 ( .A1(n8272), .A2(n9349), .ZN(n8311) );
  NAND2_X1 U9781 ( .A1(n8209), .A2(n8311), .ZN(n8210) );
  NAND2_X1 U9782 ( .A1(n8312), .A2(n8210), .ZN(n8211) );
  NAND3_X1 U9783 ( .A1(n8216), .A2(n8313), .A3(n8213), .ZN(n8214) );
  INV_X1 U9784 ( .A(n9273), .ZN(n8223) );
  AOI21_X1 U9785 ( .B1(n8214), .B2(n8220), .A(n8223), .ZN(n8215) );
  NOR2_X1 U9786 ( .A1(n8215), .A2(n8341), .ZN(n8227) );
  INV_X1 U9787 ( .A(n8216), .ZN(n8217) );
  NAND2_X1 U9788 ( .A1(n8217), .A2(n8313), .ZN(n8225) );
  INV_X1 U9789 ( .A(n8218), .ZN(n8219) );
  AND2_X1 U9790 ( .A1(n8313), .A2(n8219), .ZN(n8222) );
  INV_X1 U9791 ( .A(n8220), .ZN(n8221) );
  OR3_X1 U9792 ( .A1(n8341), .A2(n8222), .A3(n8221), .ZN(n8319) );
  INV_X1 U9793 ( .A(n8319), .ZN(n8224) );
  AOI21_X1 U9794 ( .B1(n8225), .B2(n8224), .A(n8223), .ZN(n8226) );
  MUX2_X1 U9795 ( .A(n8227), .B(n8226), .S(n8267), .Z(n8240) );
  NAND3_X1 U9796 ( .A1(n8318), .A2(n8234), .A3(n9275), .ZN(n8239) );
  INV_X1 U9797 ( .A(n8228), .ZN(n8229) );
  NAND2_X1 U9798 ( .A1(n8318), .A2(n8229), .ZN(n8230) );
  AND2_X1 U9799 ( .A1(n8230), .A2(n8234), .ZN(n8231) );
  INV_X1 U9800 ( .A(n8232), .ZN(n8233) );
  NAND2_X1 U9801 ( .A1(n8234), .A2(n8233), .ZN(n8235) );
  NAND3_X1 U9802 ( .A1(n8269), .A2(n8318), .A3(n8235), .ZN(n8236) );
  MUX2_X1 U9803 ( .A(n8400), .B(n8236), .S(n8267), .Z(n8237) );
  INV_X1 U9804 ( .A(n8237), .ZN(n8238) );
  INV_X1 U9805 ( .A(n8251), .ZN(n8254) );
  NAND2_X1 U9806 ( .A1(n9236), .A2(n8269), .ZN(n8242) );
  NAND2_X1 U9807 ( .A1(n8243), .A2(n9252), .ZN(n8241) );
  MUX2_X1 U9808 ( .A(n8242), .B(n8241), .S(n8267), .Z(n8253) );
  MUX2_X1 U9809 ( .A(n9252), .B(n9236), .S(n8262), .Z(n8250) );
  NOR2_X1 U9810 ( .A1(n8243), .A2(n9252), .ZN(n8244) );
  OR2_X1 U9811 ( .A1(n9236), .A2(n8244), .ZN(n8247) );
  OAI21_X1 U9812 ( .B1(n9236), .B2(n8269), .A(n8245), .ZN(n8246) );
  MUX2_X1 U9813 ( .A(n8247), .B(n8246), .S(n8262), .Z(n8248) );
  INV_X1 U9814 ( .A(n8248), .ZN(n8249) );
  OAI211_X1 U9815 ( .C1(n8254), .C2(n8253), .A(n8252), .B(n9215), .ZN(n8256)
         );
  MUX2_X1 U9816 ( .A(n8325), .B(n8326), .S(n8262), .Z(n8255) );
  NAND3_X1 U9817 ( .A1(n8256), .A2(n9198), .A3(n8255), .ZN(n8258) );
  MUX2_X1 U9818 ( .A(n8329), .B(n8330), .S(n8267), .Z(n8257) );
  NAND2_X1 U9819 ( .A1(n8258), .A2(n8257), .ZN(n8264) );
  NAND2_X1 U9820 ( .A1(n8264), .A2(n9125), .ZN(n8259) );
  NAND2_X1 U9821 ( .A1(n9175), .A2(n9124), .ZN(n8260) );
  INV_X1 U9822 ( .A(n8265), .ZN(n8407) );
  OAI211_X1 U9823 ( .C1(n8262), .C2(n9125), .A(n8261), .B(n8407), .ZN(n8268)
         );
  NOR2_X1 U9824 ( .A1(n8264), .A2(n9125), .ZN(n8263) );
  NOR3_X1 U9825 ( .A1(n8378), .A2(n9189), .A3(n8264), .ZN(n8266) );
  OR2_X1 U9826 ( .A1(n9172), .A2(n9175), .ZN(n8374) );
  INV_X1 U9827 ( .A(n8427), .ZN(n8428) );
  AND2_X1 U9828 ( .A1(n8270), .A2(n8269), .ZN(n8271) );
  NAND2_X1 U9829 ( .A1(n8326), .A2(n8271), .ZN(n8402) );
  INV_X1 U9830 ( .A(n8272), .ZN(n8273) );
  NOR2_X1 U9831 ( .A1(n8319), .A2(n8273), .ZN(n8396) );
  INV_X1 U9832 ( .A(n8274), .ZN(n8309) );
  NAND2_X1 U9833 ( .A1(n8276), .A2(n8275), .ZN(n8277) );
  NOR2_X1 U9834 ( .A1(n8278), .A2(n8277), .ZN(n8279) );
  NAND4_X1 U9835 ( .A1(n8302), .A2(n8299), .A3(n8291), .A4(n8279), .ZN(n8280)
         );
  OR3_X1 U9836 ( .A1(n8309), .A2(n4820), .A3(n8280), .ZN(n8394) );
  AOI21_X1 U9837 ( .B1(n9138), .B2(n8281), .A(n6657), .ZN(n8285) );
  NAND2_X1 U9838 ( .A1(n9139), .A2(n6742), .ZN(n8283) );
  AND4_X1 U9839 ( .A1(n8285), .A2(n8284), .A3(n8283), .A4(n8282), .ZN(n8286)
         );
  OAI21_X1 U9840 ( .B1(n8287), .B2(n8286), .A(n8379), .ZN(n8289) );
  NAND2_X1 U9841 ( .A1(n8381), .A2(n8380), .ZN(n8288) );
  AOI21_X1 U9842 ( .B1(n8289), .B2(n8383), .A(n8288), .ZN(n8310) );
  INV_X1 U9843 ( .A(n8290), .ZN(n8296) );
  INV_X1 U9844 ( .A(n8291), .ZN(n8295) );
  AND2_X1 U9845 ( .A1(n8293), .A2(n8292), .ZN(n8294) );
  OAI22_X1 U9846 ( .A1(n8297), .A2(n8296), .B1(n8295), .B2(n8294), .ZN(n8298)
         );
  NAND2_X1 U9847 ( .A1(n8299), .A2(n8298), .ZN(n8301) );
  NAND2_X1 U9848 ( .A1(n8301), .A2(n8300), .ZN(n8303) );
  NAND2_X1 U9849 ( .A1(n8303), .A2(n8302), .ZN(n8304) );
  NAND2_X1 U9850 ( .A1(n8305), .A2(n8304), .ZN(n8307) );
  NAND2_X1 U9851 ( .A1(n8307), .A2(n8306), .ZN(n8308) );
  OR2_X1 U9852 ( .A1(n8309), .A2(n8308), .ZN(n8392) );
  OAI21_X1 U9853 ( .B1(n8394), .B2(n8310), .A(n8392), .ZN(n8321) );
  INV_X1 U9854 ( .A(n8311), .ZN(n8314) );
  OAI211_X1 U9855 ( .C1(n8315), .C2(n8314), .A(n8313), .B(n8312), .ZN(n8316)
         );
  INV_X1 U9856 ( .A(n8316), .ZN(n8320) );
  OAI211_X1 U9857 ( .C1(n8320), .C2(n8319), .A(n8318), .B(n8317), .ZN(n8398)
         );
  AOI21_X1 U9858 ( .B1(n8396), .B2(n8321), .A(n8398), .ZN(n8322) );
  NOR2_X1 U9859 ( .A1(n8322), .A2(n8400), .ZN(n8323) );
  NOR2_X1 U9860 ( .A1(n8402), .A2(n8323), .ZN(n8332) );
  NAND2_X1 U9861 ( .A1(n8325), .A2(n8324), .ZN(n8327) );
  NAND2_X1 U9862 ( .A1(n8327), .A2(n8326), .ZN(n8328) );
  NAND2_X1 U9863 ( .A1(n8329), .A2(n8328), .ZN(n8404) );
  AND2_X1 U9864 ( .A1(n8331), .A2(n8330), .ZN(n8405) );
  OAI21_X1 U9865 ( .B1(n8332), .B2(n8404), .A(n8405), .ZN(n8334) );
  INV_X1 U9866 ( .A(n8372), .ZN(n8333) );
  AOI21_X1 U9867 ( .B1(n8406), .B2(n8334), .A(n8333), .ZN(n8337) );
  INV_X1 U9868 ( .A(n8426), .ZN(n8377) );
  NAND2_X1 U9869 ( .A1(n9180), .A2(n8335), .ZN(n8336) );
  OAI21_X1 U9870 ( .B1(n8337), .B2(n8375), .A(n8374), .ZN(n8338) );
  XNOR2_X1 U9871 ( .A(n8338), .B(n9317), .ZN(n8340) );
  NAND2_X1 U9872 ( .A1(n8340), .A2(n8339), .ZN(n8423) );
  INV_X1 U9873 ( .A(n9265), .ZN(n9258) );
  NAND2_X1 U9874 ( .A1(n4795), .A2(n9273), .ZN(n9301) );
  INV_X1 U9875 ( .A(n9376), .ZN(n9385) );
  NOR3_X1 U9876 ( .A1(n8344), .A2(n8343), .A3(n8342), .ZN(n8350) );
  AND2_X1 U9877 ( .A1(n8346), .A2(n8345), .ZN(n8348) );
  AND4_X1 U9878 ( .A1(n8350), .A2(n8349), .A3(n8348), .A4(n8347), .ZN(n8354)
         );
  NAND4_X1 U9879 ( .A1(n8354), .A2(n8353), .A3(n8352), .A4(n8351), .ZN(n8358)
         );
  NAND2_X1 U9880 ( .A1(n8356), .A2(n8355), .ZN(n9642) );
  OR3_X1 U9881 ( .A1(n8358), .A2(n8357), .A3(n9642), .ZN(n8359) );
  NOR2_X1 U9882 ( .A1(n8360), .A2(n8359), .ZN(n8362) );
  NAND4_X1 U9883 ( .A1(n9385), .A2(n9622), .A3(n8362), .A4(n8361), .ZN(n8363)
         );
  NOR2_X1 U9884 ( .A1(n9359), .A2(n8363), .ZN(n8364) );
  NAND4_X1 U9885 ( .A1(n9333), .A2(n9347), .A3(n8365), .A4(n8364), .ZN(n8366)
         );
  NOR2_X1 U9886 ( .A1(n9301), .A2(n8366), .ZN(n8367) );
  NAND3_X1 U9887 ( .A1(n9275), .A2(n8367), .A3(n9308), .ZN(n8368) );
  NOR3_X1 U9888 ( .A1(n9251), .A2(n9258), .A3(n8368), .ZN(n8369) );
  NAND4_X1 U9889 ( .A1(n9198), .A2(n9215), .A3(n9229), .A4(n8369), .ZN(n8370)
         );
  NOR2_X1 U9890 ( .A1(n8371), .A2(n8370), .ZN(n8373) );
  NAND3_X1 U9891 ( .A1(n8374), .A2(n8373), .A3(n8372), .ZN(n8376) );
  NOR2_X1 U9892 ( .A1(n8376), .A2(n8375), .ZN(n8416) );
  AND2_X1 U9893 ( .A1(n8417), .A2(n9331), .ZN(n8414) );
  AND2_X1 U9894 ( .A1(n8377), .A2(n6656), .ZN(n8413) );
  INV_X1 U9895 ( .A(n8378), .ZN(n8411) );
  NAND3_X1 U9896 ( .A1(n8381), .A2(n8380), .A3(n8379), .ZN(n8390) );
  NAND2_X1 U9897 ( .A1(n8383), .A2(n8382), .ZN(n8386) );
  INV_X1 U9898 ( .A(n8384), .ZN(n8385) );
  OAI211_X1 U9899 ( .C1(n8388), .C2(n8387), .A(n8386), .B(n8385), .ZN(n8389)
         );
  OAI21_X1 U9900 ( .B1(n8391), .B2(n8390), .A(n8389), .ZN(n8393) );
  OAI21_X1 U9901 ( .B1(n8394), .B2(n8393), .A(n8392), .ZN(n8395) );
  AND2_X1 U9902 ( .A1(n8396), .A2(n8395), .ZN(n8397) );
  NOR2_X1 U9903 ( .A1(n8398), .A2(n8397), .ZN(n8399) );
  NOR2_X1 U9904 ( .A1(n8400), .A2(n8399), .ZN(n8401) );
  NOR2_X1 U9905 ( .A1(n8402), .A2(n8401), .ZN(n8403) );
  NOR2_X1 U9906 ( .A1(n8404), .A2(n8403), .ZN(n8409) );
  INV_X1 U9907 ( .A(n8405), .ZN(n8408) );
  OAI211_X1 U9908 ( .C1(n8409), .C2(n8408), .A(n8407), .B(n8406), .ZN(n8410)
         );
  NAND2_X1 U9909 ( .A1(n8411), .A2(n8410), .ZN(n8412) );
  NAND2_X1 U9910 ( .A1(n8413), .A2(n8412), .ZN(n8415) );
  NAND3_X1 U9911 ( .A1(n8416), .A2(n8414), .A3(n8415), .ZN(n8422) );
  NAND3_X1 U9912 ( .A1(n8415), .A2(n6656), .A3(n8414), .ZN(n8421) );
  INV_X1 U9913 ( .A(n8416), .ZN(n8419) );
  NAND2_X1 U9914 ( .A1(n8417), .A2(n9317), .ZN(n8424) );
  INV_X1 U9915 ( .A(n8424), .ZN(n8418) );
  NAND3_X1 U9916 ( .A1(n8419), .A2(n8418), .A3(n6657), .ZN(n8420) );
  INV_X1 U9917 ( .A(n8429), .ZN(n8437) );
  NOR4_X1 U9918 ( .A1(n8432), .A2(n8431), .A3(n4487), .A4(n8430), .ZN(n8435)
         );
  OAI21_X1 U9919 ( .B1(n8433), .B2(n8436), .A(P1_B_REG_SCAN_IN), .ZN(n8434) );
  OAI22_X1 U9920 ( .A1(n8437), .A2(n8436), .B1(n8435), .B2(n8434), .ZN(
        P1_U3240) );
  XNOR2_X1 U9921 ( .A(n8438), .B(n8439), .ZN(n8445) );
  OAI22_X1 U9922 ( .A1(n8670), .A2(n8526), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8440), .ZN(n8441) );
  AOI21_X1 U9923 ( .B1(n8662), .B2(n8479), .A(n8441), .ZN(n8442) );
  OAI21_X1 U9924 ( .B1(n8671), .B2(n8527), .A(n8442), .ZN(n8443) );
  AOI21_X1 U9925 ( .B1(n8861), .B2(n9610), .A(n8443), .ZN(n8444) );
  OAI21_X1 U9926 ( .B1(n8445), .B2(n8542), .A(n8444), .ZN(P2_U3216) );
  INV_X1 U9927 ( .A(n8446), .ZN(n8448) );
  NOR2_X1 U9928 ( .A1(n8448), .A2(n8447), .ZN(n8494) );
  INV_X1 U9929 ( .A(n8528), .ZN(n8752) );
  AOI22_X1 U9930 ( .A1(n8446), .A2(n9611), .B1(n8521), .B2(n8752), .ZN(n8454)
         );
  INV_X1 U9931 ( .A(n8730), .ZN(n8450) );
  OAI22_X1 U9932 ( .A1(n8450), .A2(n9616), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8449), .ZN(n8452) );
  OAI22_X1 U9933 ( .A1(n8619), .A2(n8527), .B1(n8763), .B2(n8526), .ZN(n8451)
         );
  AOI211_X1 U9934 ( .C1(n8883), .C2(n9610), .A(n8452), .B(n8451), .ZN(n8453)
         );
  OAI21_X1 U9935 ( .B1(n8494), .B2(n8454), .A(n8453), .ZN(P2_U3218) );
  OAI22_X1 U9936 ( .A1(n5785), .A2(n8455), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7465), .ZN(n8456) );
  AOI21_X1 U9937 ( .B1(n8479), .B2(n7465), .A(n8456), .ZN(n8463) );
  AOI22_X1 U9938 ( .A1(n8517), .A2(n5806), .B1(n8516), .B2(n8559), .ZN(n8462)
         );
  AOI21_X1 U9939 ( .B1(n8458), .B2(n8457), .A(n8542), .ZN(n8460) );
  NAND2_X1 U9940 ( .A1(n8460), .A2(n8459), .ZN(n8461) );
  NAND3_X1 U9941 ( .A1(n8463), .A2(n8462), .A3(n8461), .ZN(P2_U3220) );
  INV_X1 U9942 ( .A(n8464), .ZN(n8465) );
  AOI21_X1 U9943 ( .B1(n8466), .B2(n8465), .A(n8542), .ZN(n8470) );
  NOR3_X1 U9944 ( .A1(n8467), .A2(n8762), .A3(n8505), .ZN(n8469) );
  OAI21_X1 U9945 ( .B1(n8470), .B2(n8469), .A(n8468), .ZN(n8475) );
  NOR2_X1 U9946 ( .A1(n8471), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8473) );
  OAI22_X1 U9947 ( .A1(n8763), .A2(n8527), .B1(n8762), .B2(n8526), .ZN(n8472)
         );
  AOI211_X1 U9948 ( .C1(n8479), .C2(n8767), .A(n8473), .B(n8472), .ZN(n8474)
         );
  OAI211_X1 U9949 ( .C1(n8770), .C2(n5785), .A(n8475), .B(n8474), .ZN(P2_U3225) );
  OR2_X1 U9950 ( .A1(n8670), .A2(n8820), .ZN(n8477) );
  NAND2_X1 U9951 ( .A1(n8618), .A2(n8750), .ZN(n8476) );
  AND2_X1 U9952 ( .A1(n8477), .A2(n8476), .ZN(n8698) );
  INV_X1 U9953 ( .A(n8478), .ZN(n8702) );
  AOI22_X1 U9954 ( .A1(n8702), .A2(n8479), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8480) );
  OAI21_X1 U9955 ( .B1(n8698), .B2(n8481), .A(n8480), .ZN(n8491) );
  INV_X1 U9956 ( .A(n8486), .ZN(n8483) );
  NOR3_X1 U9957 ( .A1(n8483), .A2(n8542), .A3(n8482), .ZN(n8489) );
  INV_X1 U9958 ( .A(n8715), .ZN(n8545) );
  NAND3_X1 U9959 ( .A1(n8484), .A2(n8521), .A3(n8545), .ZN(n8485) );
  OAI21_X1 U9960 ( .B1(n8486), .B2(n8542), .A(n8485), .ZN(n8488) );
  MUX2_X1 U9961 ( .A(n8489), .B(n8488), .S(n8487), .Z(n8490) );
  AOI211_X1 U9962 ( .C1(n9610), .C2(n8873), .A(n8491), .B(n8490), .ZN(n8492)
         );
  INV_X1 U9963 ( .A(n8492), .ZN(P2_U3227) );
  NOR2_X1 U9964 ( .A1(n8494), .A2(n8493), .ZN(n8496) );
  XNOR2_X1 U9965 ( .A(n8496), .B(n8495), .ZN(n8499) );
  OAI22_X1 U9966 ( .A1(n8499), .A2(n8542), .B1(n8619), .B2(n8505), .ZN(n8497)
         );
  OAI21_X1 U9967 ( .B1(n8499), .B2(n8498), .A(n8497), .ZN(n8503) );
  OAI22_X1 U9968 ( .A1(n8718), .A2(n9616), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10361), .ZN(n8501) );
  OAI22_X1 U9969 ( .A1(n8715), .A2(n8527), .B1(n8528), .B2(n8526), .ZN(n8500)
         );
  AOI211_X1 U9970 ( .C1(n8617), .C2(n9610), .A(n8501), .B(n8500), .ZN(n8502)
         );
  NAND2_X1 U9971 ( .A1(n8503), .A2(n8502), .ZN(P2_U3231) );
  INV_X1 U9972 ( .A(n8509), .ZN(n8507) );
  NOR3_X1 U9973 ( .A1(n8505), .A2(n8504), .A3(n5809), .ZN(n8506) );
  AOI21_X1 U9974 ( .B1(n9611), .B2(n8507), .A(n8506), .ZN(n8512) );
  NAND3_X1 U9975 ( .A1(n9611), .A2(n8509), .A3(n8508), .ZN(n8511) );
  MUX2_X1 U9976 ( .A(n8512), .B(n8511), .S(n8510), .Z(n8520) );
  AND2_X1 U9977 ( .A1(P2_U3152), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n9860) );
  NOR2_X1 U9978 ( .A1(n9616), .A2(n8513), .ZN(n8514) );
  AOI211_X1 U9979 ( .C1(n9610), .C2(n8515), .A(n9860), .B(n8514), .ZN(n8519)
         );
  AOI22_X1 U9980 ( .A1(n8517), .A2(n5807), .B1(n8516), .B2(n8558), .ZN(n8518)
         );
  NAND3_X1 U9981 ( .A1(n8520), .A2(n8519), .A3(n8518), .ZN(P2_U3232) );
  NAND2_X1 U9982 ( .A1(n8616), .A2(n8521), .ZN(n8525) );
  NAND2_X1 U9983 ( .A1(n8522), .A2(n9611), .ZN(n8524) );
  MUX2_X1 U9984 ( .A(n8525), .B(n8524), .S(n8523), .Z(n8532) );
  OAI22_X1 U9985 ( .A1(n8742), .A2(n9616), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10085), .ZN(n8530) );
  OAI22_X1 U9986 ( .A1(n8528), .A2(n8527), .B1(n8784), .B2(n8526), .ZN(n8529)
         );
  AOI211_X1 U9987 ( .C1(n8889), .C2(n9610), .A(n8530), .B(n8529), .ZN(n8531)
         );
  NAND2_X1 U9988 ( .A1(n8532), .A2(n8531), .ZN(P2_U3237) );
  XNOR2_X1 U9989 ( .A(n8534), .B(n8533), .ZN(n8543) );
  OR2_X1 U9990 ( .A1(n8654), .A2(n8820), .ZN(n8536) );
  NAND2_X1 U9991 ( .A1(n8545), .A2(n8750), .ZN(n8535) );
  NAND2_X1 U9992 ( .A1(n8536), .A2(n8535), .ZN(n8690) );
  INV_X1 U9993 ( .A(n8681), .ZN(n8538) );
  OAI22_X1 U9994 ( .A1(n8538), .A2(n9616), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8537), .ZN(n8539) );
  AOI21_X1 U9995 ( .B1(n8690), .B2(n9606), .A(n8539), .ZN(n8541) );
  NAND2_X1 U9996 ( .A1(n8867), .A2(n9610), .ZN(n8540) );
  OAI211_X1 U9997 ( .C1(n8543), .C2(n8542), .A(n8541), .B(n8540), .ZN(P2_U3242) );
  MUX2_X1 U9998 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8629), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9999 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8544), .S(P2_U3966), .Z(
        P2_U3581) );
  MUX2_X1 U10000 ( .A(n8628), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8560), .Z(
        P2_U3580) );
  INV_X1 U10001 ( .A(n8670), .ZN(n8622) );
  MUX2_X1 U10002 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8622), .S(P2_U3966), .Z(
        P2_U3578) );
  MUX2_X1 U10003 ( .A(n8545), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8560), .Z(
        P2_U3577) );
  MUX2_X1 U10004 ( .A(n8618), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8560), .Z(
        P2_U3576) );
  MUX2_X1 U10005 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8752), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U10006 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8616), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U10007 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8749), .S(P2_U3966), .Z(
        P2_U3573) );
  INV_X1 U10008 ( .A(n8762), .ZN(n8614) );
  MUX2_X1 U10009 ( .A(n8614), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8560), .Z(
        P2_U3572) );
  MUX2_X1 U10010 ( .A(n8611), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8560), .Z(
        P2_U3570) );
  MUX2_X1 U10011 ( .A(n8546), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8560), .Z(
        P2_U3569) );
  MUX2_X1 U10012 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8547), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10013 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8548), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10014 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8549), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U10015 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8550), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U10016 ( .A(n8551), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8560), .Z(
        P2_U3564) );
  MUX2_X1 U10017 ( .A(n8552), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8560), .Z(
        P2_U3563) );
  MUX2_X1 U10018 ( .A(n8553), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8560), .Z(
        P2_U3562) );
  MUX2_X1 U10019 ( .A(n8554), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8560), .Z(
        P2_U3561) );
  MUX2_X1 U10020 ( .A(n8555), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8560), .Z(
        P2_U3560) );
  MUX2_X1 U10021 ( .A(n8556), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8560), .Z(
        P2_U3559) );
  MUX2_X1 U10022 ( .A(n8557), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8560), .Z(
        P2_U3558) );
  MUX2_X1 U10023 ( .A(n8558), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8560), .Z(
        P2_U3557) );
  MUX2_X1 U10024 ( .A(n8559), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8560), .Z(
        P2_U3556) );
  MUX2_X1 U10025 ( .A(n5807), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8560), .Z(
        P2_U3555) );
  MUX2_X1 U10026 ( .A(n5806), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8560), .Z(
        P2_U3554) );
  MUX2_X1 U10027 ( .A(n5805), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8560), .Z(
        P2_U3553) );
  MUX2_X1 U10028 ( .A(n8561), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8560), .Z(
        P2_U3552) );
  INV_X1 U10029 ( .A(n8578), .ZN(n8585) );
  OR2_X1 U10030 ( .A1(n8578), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8582) );
  NAND2_X1 U10031 ( .A1(n8578), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8562) );
  AND2_X1 U10032 ( .A1(n8582), .A2(n8562), .ZN(n8568) );
  INV_X1 U10033 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8565) );
  AOI21_X1 U10034 ( .B1(n8575), .B2(n8564), .A(n8563), .ZN(n9909) );
  XNOR2_X1 U10035 ( .A(n8573), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n9908) );
  NAND2_X1 U10036 ( .A1(n9909), .A2(n9908), .ZN(n9907) );
  OAI21_X1 U10037 ( .B1(n8565), .B2(n8573), .A(n9907), .ZN(n8566) );
  INV_X1 U10038 ( .A(n8566), .ZN(n8567) );
  NAND2_X1 U10039 ( .A1(n8568), .A2(n8567), .ZN(n8583) );
  OAI21_X1 U10040 ( .B1(n8568), .B2(n8567), .A(n8583), .ZN(n8572) );
  NOR2_X1 U10041 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10427), .ZN(n8571) );
  INV_X1 U10042 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8569) );
  NOR2_X1 U10043 ( .A1(n9566), .A2(n8569), .ZN(n8570) );
  AOI211_X1 U10044 ( .C1(n9906), .C2(n8572), .A(n8571), .B(n8570), .ZN(n8581)
         );
  XNOR2_X1 U10045 ( .A(n8573), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n9902) );
  OAI21_X1 U10046 ( .B1(n8576), .B2(n8575), .A(n8574), .ZN(n9903) );
  NAND2_X1 U10047 ( .A1(n9902), .A2(n9903), .ZN(n9900) );
  INV_X1 U10048 ( .A(n9900), .ZN(n8577) );
  AOI21_X1 U10049 ( .B1(n9904), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8577), .ZN(
        n8586) );
  XNOR2_X1 U10050 ( .A(n8586), .B(n8578), .ZN(n8579) );
  NAND2_X1 U10051 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8579), .ZN(n8588) );
  OAI211_X1 U10052 ( .C1(P2_REG2_REG_18__SCAN_IN), .C2(n8579), .A(n9901), .B(
        n8588), .ZN(n8580) );
  OAI211_X1 U10053 ( .C1(n9842), .C2(n8585), .A(n8581), .B(n8580), .ZN(
        P2_U3263) );
  NAND2_X1 U10054 ( .A1(n8583), .A2(n8582), .ZN(n8584) );
  XNOR2_X1 U10055 ( .A(n8584), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8591) );
  OR2_X1 U10056 ( .A1(n8586), .A2(n8585), .ZN(n8587) );
  NAND2_X1 U10057 ( .A1(n8588), .A2(n8587), .ZN(n8589) );
  XNOR2_X1 U10058 ( .A(n8589), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8593) );
  NAND2_X1 U10059 ( .A1(n8593), .A2(n9901), .ZN(n8590) );
  OAI211_X1 U10060 ( .C1(n8591), .C2(n9843), .A(n8590), .B(n9842), .ZN(n8595)
         );
  INV_X1 U10061 ( .A(n8591), .ZN(n8592) );
  OAI22_X1 U10062 ( .A1(n8593), .A2(n9841), .B1(n8592), .B2(n9843), .ZN(n8594)
         );
  MUX2_X1 U10063 ( .A(n8595), .B(n8594), .S(n8835), .Z(n8596) );
  INV_X1 U10064 ( .A(n8596), .ZN(n8598) );
  NAND2_X1 U10065 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8597) );
  OAI211_X1 U10066 ( .C1(n5108), .C2(n9566), .A(n8598), .B(n8597), .ZN(
        P2_U3264) );
  INV_X1 U10067 ( .A(n8867), .ZN(n8683) );
  INV_X1 U10068 ( .A(n8909), .ZN(n8814) );
  NAND2_X1 U10069 ( .A1(n8814), .A2(n8806), .ZN(n8807) );
  NAND2_X1 U10070 ( .A1(n8683), .A2(n8700), .ZN(n8678) );
  INV_X1 U10071 ( .A(n5817), .ZN(n8649) );
  AOI21_X1 U10072 ( .B1(n8599), .B2(P2_B_REG_SCAN_IN), .A(n8820), .ZN(n8630)
         );
  NAND2_X1 U10073 ( .A1(n8600), .A2(n8630), .ZN(n8849) );
  NOR2_X1 U10074 ( .A1(n9936), .A2(n8849), .ZN(n8604) );
  AOI21_X1 U10075 ( .B1(n9936), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8604), .ZN(
        n8602) );
  NAND2_X1 U10076 ( .A1(n8844), .A2(n9926), .ZN(n8601) );
  OAI211_X1 U10077 ( .C1(n8846), .C2(n8717), .A(n8602), .B(n8601), .ZN(
        P2_U3265) );
  INV_X1 U10078 ( .A(n8635), .ZN(n8603) );
  NAND2_X1 U10079 ( .A1(n5839), .A2(n8603), .ZN(n8847) );
  NAND3_X1 U10080 ( .A1(n8848), .A2(n9932), .A3(n8847), .ZN(n8606) );
  AOI21_X1 U10081 ( .B1(n9936), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8604), .ZN(
        n8605) );
  OAI211_X1 U10082 ( .C1(n8851), .C2(n8813), .A(n8606), .B(n8605), .ZN(
        P2_U3266) );
  NAND2_X1 U10083 ( .A1(n8608), .A2(n5095), .ZN(n8827) );
  AOI22_X1 U10084 ( .A1(n8773), .A2(n8782), .B1(n8900), .B2(n8614), .ZN(n8758)
         );
  NAND2_X1 U10085 ( .A1(n8895), .A2(n8749), .ZN(n8615) );
  NAND2_X1 U10086 ( .A1(n8710), .A2(n8709), .ZN(n8708) );
  NAND2_X1 U10087 ( .A1(n8708), .A2(n8620), .ZN(n8695) );
  INV_X1 U10088 ( .A(n8873), .ZN(n8705) );
  INV_X1 U10089 ( .A(n8861), .ZN(n8664) );
  XNOR2_X1 U10090 ( .A(n8625), .B(n8624), .ZN(n8856) );
  NAND2_X1 U10091 ( .A1(n8628), .A2(n8750), .ZN(n8632) );
  NAND2_X1 U10092 ( .A1(n8630), .A2(n8629), .ZN(n8631) );
  INV_X1 U10093 ( .A(n8855), .ZN(n8640) );
  AOI21_X1 U10094 ( .B1(n8852), .B2(n8643), .A(n8635), .ZN(n8853) );
  NAND2_X1 U10095 ( .A1(n8853), .A2(n9932), .ZN(n8638) );
  AOI22_X1 U10096 ( .A1(n8636), .A2(n9925), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n9936), .ZN(n8637) );
  OAI211_X1 U10097 ( .C1(n4785), .C2(n8813), .A(n8638), .B(n8637), .ZN(n8639)
         );
  AOI21_X1 U10098 ( .B1(n8640), .B2(n8839), .A(n8639), .ZN(n8641) );
  OAI21_X1 U10099 ( .B1(n8856), .B2(n8843), .A(n8641), .ZN(P2_U3267) );
  XNOR2_X1 U10100 ( .A(n8642), .B(n8651), .ZN(n8860) );
  INV_X1 U10101 ( .A(n8661), .ZN(n8645) );
  INV_X1 U10102 ( .A(n8643), .ZN(n8644) );
  AOI21_X1 U10103 ( .B1(n5817), .B2(n8645), .A(n8644), .ZN(n8857) );
  INV_X1 U10104 ( .A(n8646), .ZN(n8647) );
  AOI22_X1 U10105 ( .A1(n8647), .A2(n9925), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n9936), .ZN(n8648) );
  OAI21_X1 U10106 ( .B1(n8649), .B2(n8813), .A(n8648), .ZN(n8658) );
  AOI211_X1 U10107 ( .C1(n8652), .C2(n8651), .A(n9917), .B(n8650), .ZN(n8656)
         );
  OAI22_X1 U10108 ( .A1(n8654), .A2(n8818), .B1(n8653), .B2(n8820), .ZN(n8655)
         );
  NOR2_X1 U10109 ( .A1(n8656), .A2(n8655), .ZN(n8859) );
  NOR2_X1 U10110 ( .A1(n8859), .A2(n9936), .ZN(n8657) );
  AOI211_X1 U10111 ( .C1(n9932), .C2(n8857), .A(n8658), .B(n8657), .ZN(n8659)
         );
  OAI21_X1 U10112 ( .B1(n8860), .B2(n8843), .A(n8659), .ZN(P2_U3268) );
  XNOR2_X1 U10113 ( .A(n8660), .B(n8666), .ZN(n8865) );
  AOI21_X1 U10114 ( .B1(n8861), .B2(n8678), .A(n8661), .ZN(n8862) );
  AOI22_X1 U10115 ( .A1(n8662), .A2(n9925), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n9936), .ZN(n8663) );
  OAI21_X1 U10116 ( .B1(n8664), .B2(n8813), .A(n8663), .ZN(n8675) );
  INV_X1 U10117 ( .A(n8665), .ZN(n8669) );
  AOI21_X1 U10118 ( .B1(n8687), .B2(n8667), .A(n8666), .ZN(n8668) );
  NOR3_X1 U10119 ( .A1(n8669), .A2(n8668), .A3(n9917), .ZN(n8673) );
  OAI22_X1 U10120 ( .A1(n8671), .A2(n8820), .B1(n8670), .B2(n8818), .ZN(n8672)
         );
  NOR2_X1 U10121 ( .A1(n8673), .A2(n8672), .ZN(n8864) );
  NOR2_X1 U10122 ( .A1(n8864), .A2(n9936), .ZN(n8674) );
  AOI211_X1 U10123 ( .C1(n9932), .C2(n8862), .A(n8675), .B(n8674), .ZN(n8676)
         );
  OAI21_X1 U10124 ( .B1(n8865), .B2(n8843), .A(n8676), .ZN(P2_U3269) );
  XOR2_X1 U10125 ( .A(n8688), .B(n8677), .Z(n8870) );
  INV_X1 U10126 ( .A(n8700), .ZN(n8680) );
  INV_X1 U10127 ( .A(n8678), .ZN(n8679) );
  AOI211_X1 U10128 ( .C1(n8867), .C2(n8680), .A(n10013), .B(n8679), .ZN(n8866)
         );
  AOI22_X1 U10129 ( .A1(n8681), .A2(n9925), .B1(P2_REG2_REG_26__SCAN_IN), .B2(
        n9936), .ZN(n8682) );
  OAI21_X1 U10130 ( .B1(n8683), .B2(n8813), .A(n8682), .ZN(n8693) );
  INV_X1 U10131 ( .A(n8684), .ZN(n8686) );
  NOR2_X1 U10132 ( .A1(n8686), .A2(n8685), .ZN(n8689) );
  OAI21_X1 U10133 ( .B1(n8689), .B2(n8688), .A(n8687), .ZN(n8691) );
  AOI21_X1 U10134 ( .B1(n8691), .B2(n8795), .A(n8690), .ZN(n8869) );
  NOR2_X1 U10135 ( .A1(n8869), .A2(n9936), .ZN(n8692) );
  AOI211_X1 U10136 ( .C1(n8866), .C2(n8701), .A(n8693), .B(n8692), .ZN(n8694)
         );
  OAI21_X1 U10137 ( .B1(n8870), .B2(n8843), .A(n8694), .ZN(P2_U3270) );
  XNOR2_X1 U10138 ( .A(n8695), .B(n8697), .ZN(n8875) );
  OAI211_X1 U10139 ( .C1(n8697), .C2(n8696), .A(n8684), .B(n8795), .ZN(n8699)
         );
  NAND2_X1 U10140 ( .A1(n8699), .A2(n8698), .ZN(n8871) );
  AOI211_X1 U10141 ( .C1(n8873), .C2(n8716), .A(n10013), .B(n8700), .ZN(n8872)
         );
  NAND2_X1 U10142 ( .A1(n8872), .A2(n8701), .ZN(n8704) );
  AOI22_X1 U10143 ( .A1(n8702), .A2(n9925), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n9936), .ZN(n8703) );
  OAI211_X1 U10144 ( .C1(n8705), .C2(n8813), .A(n8704), .B(n8703), .ZN(n8706)
         );
  AOI21_X1 U10145 ( .B1(n8871), .B2(n8839), .A(n8706), .ZN(n8707) );
  OAI21_X1 U10146 ( .B1(n8875), .B2(n8843), .A(n8707), .ZN(P2_U3271) );
  OAI21_X1 U10147 ( .B1(n8710), .B2(n8709), .A(n8708), .ZN(n8880) );
  INV_X1 U10148 ( .A(n8880), .ZN(n8724) );
  OAI211_X1 U10149 ( .C1(n4568), .C2(n8712), .A(n8711), .B(n8795), .ZN(n8714)
         );
  NAND2_X1 U10150 ( .A1(n8752), .A2(n8750), .ZN(n8713) );
  OAI211_X1 U10151 ( .C1(n8715), .C2(n8820), .A(n8714), .B(n8713), .ZN(n8879)
         );
  OAI21_X1 U10152 ( .B1(n8876), .B2(n4572), .A(n8716), .ZN(n8877) );
  NOR2_X1 U10153 ( .A1(n8877), .A2(n8717), .ZN(n8722) );
  INV_X1 U10154 ( .A(n8718), .ZN(n8719) );
  AOI22_X1 U10155 ( .A1(n8719), .A2(n9925), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n9936), .ZN(n8720) );
  OAI21_X1 U10156 ( .B1(n8876), .B2(n8813), .A(n8720), .ZN(n8721) );
  AOI211_X1 U10157 ( .C1(n8879), .C2(n8839), .A(n8722), .B(n8721), .ZN(n8723)
         );
  OAI21_X1 U10158 ( .B1(n8724), .B2(n8843), .A(n8723), .ZN(P2_U3272) );
  AOI21_X1 U10159 ( .B1(n8727), .B2(n8726), .A(n8725), .ZN(n8728) );
  OAI222_X1 U10160 ( .A1(n8818), .A2(n8763), .B1(n8820), .B2(n8619), .C1(n9917), .C2(n8728), .ZN(n8729) );
  INV_X1 U10161 ( .A(n8729), .ZN(n8886) );
  AOI21_X1 U10162 ( .B1(n8883), .B2(n8740), .A(n4572), .ZN(n8884) );
  INV_X1 U10163 ( .A(n8883), .ZN(n8732) );
  AOI22_X1 U10164 ( .A1(n8730), .A2(n9925), .B1(P2_REG2_REG_23__SCAN_IN), .B2(
        n9936), .ZN(n8731) );
  OAI21_X1 U10165 ( .B1(n8732), .B2(n8813), .A(n8731), .ZN(n8733) );
  AOI21_X1 U10166 ( .B1(n8884), .B2(n9932), .A(n8733), .ZN(n8738) );
  NAND2_X1 U10167 ( .A1(n8735), .A2(n8734), .ZN(n8882) );
  NAND3_X1 U10168 ( .A1(n4883), .A2(n8736), .A3(n8882), .ZN(n8737) );
  OAI211_X1 U10169 ( .C1(n8886), .C2(n9936), .A(n8738), .B(n8737), .ZN(
        P2_U3273) );
  XOR2_X1 U10170 ( .A(n8747), .B(n8739), .Z(n8893) );
  INV_X1 U10171 ( .A(n8740), .ZN(n8741) );
  AOI21_X1 U10172 ( .B1(n8889), .B2(n8764), .A(n8741), .ZN(n8890) );
  INV_X1 U10173 ( .A(n8889), .ZN(n8745) );
  INV_X1 U10174 ( .A(n8742), .ZN(n8743) );
  AOI22_X1 U10175 ( .A1(n8743), .A2(n9925), .B1(n9936), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n8744) );
  OAI21_X1 U10176 ( .B1(n8745), .B2(n8813), .A(n8744), .ZN(n8756) );
  OAI211_X1 U10177 ( .C1(n8748), .C2(n8747), .A(n8746), .B(n8795), .ZN(n8754)
         );
  AOI22_X1 U10178 ( .A1(n8752), .A2(n8751), .B1(n8750), .B2(n8749), .ZN(n8753)
         );
  AND2_X1 U10179 ( .A1(n8754), .A2(n8753), .ZN(n8892) );
  NOR2_X1 U10180 ( .A1(n8892), .A2(n9936), .ZN(n8755) );
  AOI211_X1 U10181 ( .C1(n8890), .C2(n9932), .A(n8756), .B(n8755), .ZN(n8757)
         );
  OAI21_X1 U10182 ( .B1(n8893), .B2(n8843), .A(n8757), .ZN(P2_U3274) );
  XOR2_X1 U10183 ( .A(n8758), .B(n8760), .Z(n8899) );
  AOI21_X1 U10184 ( .B1(n8760), .B2(n8759), .A(n4536), .ZN(n8761) );
  OAI222_X1 U10185 ( .A1(n8820), .A2(n8763), .B1(n8818), .B2(n8762), .C1(n9917), .C2(n8761), .ZN(n8894) );
  INV_X1 U10186 ( .A(n8775), .ZN(n8766) );
  INV_X1 U10187 ( .A(n8764), .ZN(n8765) );
  AOI21_X1 U10188 ( .B1(n8895), .B2(n8766), .A(n8765), .ZN(n8896) );
  NAND2_X1 U10189 ( .A1(n8896), .A2(n9932), .ZN(n8769) );
  AOI22_X1 U10190 ( .A1(n9936), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8767), .B2(
        n9925), .ZN(n8768) );
  OAI211_X1 U10191 ( .C1(n8770), .C2(n8813), .A(n8769), .B(n8768), .ZN(n8771)
         );
  AOI21_X1 U10192 ( .B1(n8894), .B2(n8839), .A(n8771), .ZN(n8772) );
  OAI21_X1 U10193 ( .B1(n8899), .B2(n8843), .A(n8772), .ZN(P2_U3275) );
  XNOR2_X1 U10194 ( .A(n8773), .B(n8782), .ZN(n8904) );
  INV_X1 U10195 ( .A(n8774), .ZN(n8776) );
  AOI21_X1 U10196 ( .B1(n8900), .B2(n8776), .A(n8775), .ZN(n8901) );
  INV_X1 U10197 ( .A(n8777), .ZN(n8778) );
  AOI22_X1 U10198 ( .A1(n9936), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8778), .B2(
        n9925), .ZN(n8779) );
  OAI21_X1 U10199 ( .B1(n8780), .B2(n8813), .A(n8779), .ZN(n8789) );
  INV_X1 U10200 ( .A(n8781), .ZN(n8783) );
  AOI21_X1 U10201 ( .B1(n8783), .B2(n8782), .A(n9917), .ZN(n8787) );
  OAI22_X1 U10202 ( .A1(n8784), .A2(n8820), .B1(n8821), .B2(n8818), .ZN(n8785)
         );
  AOI21_X1 U10203 ( .B1(n8787), .B2(n8786), .A(n8785), .ZN(n8903) );
  NOR2_X1 U10204 ( .A1(n8903), .A2(n9936), .ZN(n8788) );
  AOI211_X1 U10205 ( .C1(n8901), .C2(n9932), .A(n8789), .B(n8788), .ZN(n8790)
         );
  OAI21_X1 U10206 ( .B1(n8843), .B2(n8904), .A(n8790), .ZN(P2_U3276) );
  XNOR2_X1 U10207 ( .A(n4577), .B(n8792), .ZN(n8908) );
  NOR2_X1 U10208 ( .A1(n8815), .A2(n8791), .ZN(n8793) );
  XNOR2_X1 U10209 ( .A(n8793), .B(n8792), .ZN(n8796) );
  AOI21_X1 U10210 ( .B1(n8796), .B2(n8795), .A(n8794), .ZN(n8798) );
  AOI21_X1 U10211 ( .B1(n8798), .B2(n8797), .A(n9936), .ZN(n8804) );
  XNOR2_X1 U10212 ( .A(n8906), .B(n8807), .ZN(n8799) );
  OAI21_X1 U10213 ( .B1(n10013), .B2(n8799), .A(n8798), .ZN(n8905) );
  AOI22_X1 U10214 ( .A1(n9936), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8800), .B2(
        n9925), .ZN(n8801) );
  OAI21_X1 U10215 ( .B1(n8802), .B2(n8813), .A(n8801), .ZN(n8803) );
  AOI21_X1 U10216 ( .B1(n8804), .B2(n8905), .A(n8803), .ZN(n8805) );
  OAI21_X1 U10217 ( .B1(n8843), .B2(n8908), .A(n8805), .ZN(P2_U3277) );
  XNOR2_X1 U10218 ( .A(n4494), .B(n8816), .ZN(n8913) );
  INV_X1 U10219 ( .A(n8806), .ZN(n8809) );
  INV_X1 U10220 ( .A(n8807), .ZN(n8808) );
  AOI21_X1 U10221 ( .B1(n8909), .B2(n8809), .A(n8808), .ZN(n8910) );
  INV_X1 U10222 ( .A(n8810), .ZN(n8811) );
  AOI22_X1 U10223 ( .A1(n9936), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8811), .B2(
        n9925), .ZN(n8812) );
  OAI21_X1 U10224 ( .B1(n8814), .B2(n8813), .A(n8812), .ZN(n8825) );
  AOI211_X1 U10225 ( .C1(n8817), .C2(n8816), .A(n9917), .B(n8815), .ZN(n8823)
         );
  OAI22_X1 U10226 ( .A1(n8821), .A2(n8820), .B1(n8819), .B2(n8818), .ZN(n8822)
         );
  NOR2_X1 U10227 ( .A1(n8823), .A2(n8822), .ZN(n8912) );
  NOR2_X1 U10228 ( .A1(n8912), .A2(n9936), .ZN(n8824) );
  AOI211_X1 U10229 ( .C1(n8910), .C2(n9932), .A(n8825), .B(n8824), .ZN(n8826)
         );
  OAI21_X1 U10230 ( .B1(n8913), .B2(n8843), .A(n8826), .ZN(P2_U3278) );
  AOI21_X1 U10231 ( .B1(n8828), .B2(n8827), .A(n4579), .ZN(n8917) );
  XNOR2_X1 U10232 ( .A(n4586), .B(n8828), .ZN(n8830) );
  OAI21_X1 U10233 ( .B1(n8830), .B2(n9917), .A(n8829), .ZN(n8834) );
  XNOR2_X1 U10234 ( .A(n8831), .B(n8914), .ZN(n8832) );
  AOI21_X1 U10235 ( .B1(n6882), .B2(n8832), .A(n8834), .ZN(n8916) );
  INV_X1 U10236 ( .A(n8916), .ZN(n8833) );
  OAI211_X1 U10237 ( .C1(n8835), .C2(n8834), .A(n8833), .B(n8839), .ZN(n8842)
         );
  INV_X1 U10238 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8838) );
  OAI22_X1 U10239 ( .A1(n8839), .A2(n8838), .B1(n8837), .B2(n8836), .ZN(n8840)
         );
  AOI21_X1 U10240 ( .B1(n8914), .B2(n9926), .A(n8840), .ZN(n8841) );
  OAI211_X1 U10241 ( .C1(n8843), .C2(n8917), .A(n8842), .B(n8841), .ZN(
        P2_U3279) );
  NAND2_X1 U10242 ( .A1(n8844), .A2(n8930), .ZN(n8845) );
  OAI211_X1 U10243 ( .C1(n8846), .C2(n10013), .A(n8845), .B(n8849), .ZN(n8943)
         );
  MUX2_X1 U10244 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8943), .S(n10036), .Z(
        P2_U3551) );
  NAND3_X1 U10245 ( .A1(n8848), .A2(n6882), .A3(n8847), .ZN(n8850) );
  OAI211_X1 U10246 ( .C1(n8851), .C2(n10011), .A(n8850), .B(n8849), .ZN(n8944)
         );
  MUX2_X1 U10247 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8944), .S(n10036), .Z(
        P2_U3550) );
  AOI22_X1 U10248 ( .A1(n8853), .A2(n6882), .B1(n8930), .B2(n8852), .ZN(n8854)
         );
  OAI211_X1 U10249 ( .C1(n8856), .C2(n8934), .A(n8855), .B(n8854), .ZN(n8945)
         );
  MUX2_X1 U10250 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8945), .S(n10036), .Z(
        P2_U3549) );
  AOI22_X1 U10251 ( .A1(n8857), .A2(n6882), .B1(n8930), .B2(n5817), .ZN(n8858)
         );
  OAI211_X1 U10252 ( .C1(n8860), .C2(n8934), .A(n8859), .B(n8858), .ZN(n8946)
         );
  MUX2_X1 U10253 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8946), .S(n10036), .Z(
        P2_U3548) );
  AOI22_X1 U10254 ( .A1(n8862), .A2(n6882), .B1(n8930), .B2(n8861), .ZN(n8863)
         );
  OAI211_X1 U10255 ( .C1(n8865), .C2(n8934), .A(n8864), .B(n8863), .ZN(n8947)
         );
  MUX2_X1 U10256 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8947), .S(n10036), .Z(
        P2_U3547) );
  AOI21_X1 U10257 ( .B1(n8930), .B2(n8867), .A(n8866), .ZN(n8868) );
  OAI211_X1 U10258 ( .C1(n8870), .C2(n8934), .A(n8869), .B(n8868), .ZN(n8948)
         );
  MUX2_X1 U10259 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8948), .S(n10036), .Z(
        P2_U3546) );
  AOI211_X1 U10260 ( .C1(n8930), .C2(n8873), .A(n8872), .B(n8871), .ZN(n8874)
         );
  OAI21_X1 U10261 ( .B1(n8875), .B2(n8934), .A(n8874), .ZN(n8949) );
  MUX2_X1 U10262 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8949), .S(n10036), .Z(
        P2_U3545) );
  OAI22_X1 U10263 ( .A1(n8877), .A2(n10013), .B1(n8876), .B2(n10011), .ZN(
        n8878) );
  AOI211_X1 U10264 ( .C1(n8880), .C2(n10018), .A(n8879), .B(n8878), .ZN(n8881)
         );
  INV_X1 U10265 ( .A(n8881), .ZN(n8950) );
  MUX2_X1 U10266 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8950), .S(n10036), .Z(
        P2_U3544) );
  NAND2_X1 U10267 ( .A1(n8882), .A2(n10018), .ZN(n8887) );
  AOI22_X1 U10268 ( .A1(n8884), .A2(n6882), .B1(n8930), .B2(n8883), .ZN(n8885)
         );
  OAI211_X1 U10269 ( .C1(n8888), .C2(n8887), .A(n8886), .B(n8885), .ZN(n8951)
         );
  MUX2_X1 U10270 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8951), .S(n10036), .Z(
        P2_U3543) );
  AOI22_X1 U10271 ( .A1(n8890), .A2(n6882), .B1(n8930), .B2(n8889), .ZN(n8891)
         );
  OAI211_X1 U10272 ( .C1(n8893), .C2(n8934), .A(n8892), .B(n8891), .ZN(n8952)
         );
  MUX2_X1 U10273 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8952), .S(n10036), .Z(
        P2_U3542) );
  INV_X1 U10274 ( .A(n8894), .ZN(n8898) );
  AOI22_X1 U10275 ( .A1(n8896), .A2(n6882), .B1(n8930), .B2(n8895), .ZN(n8897)
         );
  OAI211_X1 U10276 ( .C1(n8934), .C2(n8899), .A(n8898), .B(n8897), .ZN(n8953)
         );
  MUX2_X1 U10277 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8953), .S(n10036), .Z(
        P2_U3541) );
  AOI22_X1 U10278 ( .A1(n8901), .A2(n6882), .B1(n8930), .B2(n8900), .ZN(n8902)
         );
  OAI211_X1 U10279 ( .C1(n8904), .C2(n8934), .A(n8903), .B(n8902), .ZN(n8954)
         );
  MUX2_X1 U10280 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8954), .S(n10036), .Z(
        P2_U3540) );
  AOI21_X1 U10281 ( .B1(n8930), .B2(n8906), .A(n8905), .ZN(n8907) );
  OAI21_X1 U10282 ( .B1(n8934), .B2(n8908), .A(n8907), .ZN(n8955) );
  MUX2_X1 U10283 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8955), .S(n10036), .Z(
        P2_U3539) );
  AOI22_X1 U10284 ( .A1(n8910), .A2(n6882), .B1(n8930), .B2(n8909), .ZN(n8911)
         );
  OAI211_X1 U10285 ( .C1(n8913), .C2(n8934), .A(n8912), .B(n8911), .ZN(n8956)
         );
  MUX2_X1 U10286 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8956), .S(n10036), .Z(
        P2_U3538) );
  NAND2_X1 U10287 ( .A1(n8914), .A2(n8930), .ZN(n8915) );
  OAI211_X1 U10288 ( .C1(n8917), .C2(n8934), .A(n8916), .B(n8915), .ZN(n8957)
         );
  MUX2_X1 U10289 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8957), .S(n10036), .Z(
        P2_U3537) );
  INV_X1 U10290 ( .A(n8918), .ZN(n8924) );
  OAI22_X1 U10291 ( .A1(n8920), .A2(n10013), .B1(n8919), .B2(n10011), .ZN(
        n8921) );
  INV_X1 U10292 ( .A(n8921), .ZN(n8922) );
  OAI211_X1 U10293 ( .C1(n8939), .C2(n8924), .A(n8923), .B(n8922), .ZN(n8958)
         );
  MUX2_X1 U10294 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8958), .S(n10036), .Z(
        P2_U3536) );
  AOI22_X1 U10295 ( .A1(n8925), .A2(n6882), .B1(n8930), .B2(n9609), .ZN(n8926)
         );
  OAI211_X1 U10296 ( .C1(n8928), .C2(n8934), .A(n8927), .B(n8926), .ZN(n8959)
         );
  MUX2_X1 U10297 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8959), .S(n10036), .Z(
        P2_U3535) );
  INV_X1 U10298 ( .A(n8929), .ZN(n8935) );
  AOI22_X1 U10299 ( .A1(n8931), .A2(n6882), .B1(n8930), .B2(n9600), .ZN(n8932)
         );
  OAI211_X1 U10300 ( .C1(n8935), .C2(n8934), .A(n8933), .B(n8932), .ZN(n8960)
         );
  MUX2_X1 U10301 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8960), .S(n10036), .Z(
        P2_U3534) );
  OAI22_X1 U10302 ( .A1(n8936), .A2(n10013), .B1(n4786), .B2(n10011), .ZN(
        n8937) );
  INV_X1 U10303 ( .A(n8937), .ZN(n8938) );
  OAI21_X1 U10304 ( .B1(n8940), .B2(n8939), .A(n8938), .ZN(n8941) );
  OR2_X1 U10305 ( .A1(n8942), .A2(n8941), .ZN(n8961) );
  MUX2_X1 U10306 ( .A(n8961), .B(P2_REG1_REG_13__SCAN_IN), .S(n10033), .Z(
        P2_U3533) );
  MUX2_X1 U10307 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8943), .S(n10021), .Z(
        P2_U3519) );
  MUX2_X1 U10308 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8944), .S(n10021), .Z(
        P2_U3518) );
  MUX2_X1 U10309 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8945), .S(n10021), .Z(
        P2_U3517) );
  MUX2_X1 U10310 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8946), .S(n10021), .Z(
        P2_U3516) );
  MUX2_X1 U10311 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8947), .S(n10021), .Z(
        P2_U3515) );
  MUX2_X1 U10312 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8948), .S(n10021), .Z(
        P2_U3514) );
  MUX2_X1 U10313 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8949), .S(n10021), .Z(
        P2_U3513) );
  MUX2_X1 U10314 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8950), .S(n10021), .Z(
        P2_U3512) );
  MUX2_X1 U10315 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8951), .S(n10021), .Z(
        P2_U3511) );
  MUX2_X1 U10316 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8952), .S(n10021), .Z(
        P2_U3510) );
  MUX2_X1 U10317 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8953), .S(n10021), .Z(
        P2_U3509) );
  MUX2_X1 U10318 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8954), .S(n10021), .Z(
        P2_U3508) );
  MUX2_X1 U10319 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8955), .S(n10021), .Z(
        P2_U3507) );
  MUX2_X1 U10320 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8956), .S(n10021), .Z(
        P2_U3505) );
  MUX2_X1 U10321 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8957), .S(n10021), .Z(
        P2_U3502) );
  MUX2_X1 U10322 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8958), .S(n10021), .Z(
        P2_U3499) );
  MUX2_X1 U10323 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8959), .S(n10021), .Z(
        P2_U3496) );
  MUX2_X1 U10324 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8960), .S(n10021), .Z(
        P2_U3493) );
  MUX2_X1 U10325 ( .A(n8961), .B(P2_REG0_REG_13__SCAN_IN), .S(n10019), .Z(
        P2_U3490) );
  INV_X1 U10326 ( .A(n8962), .ZN(n9541) );
  NAND4_X1 U10327 ( .A1(n8963), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .A4(n8964), .ZN(n8967) );
  NAND2_X1 U10328 ( .A1(n8965), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8966) );
  OAI211_X1 U10329 ( .C1(n9541), .C2(n8968), .A(n8967), .B(n8966), .ZN(
        P2_U3327) );
  OAI222_X1 U10330 ( .A1(n8983), .A2(n8971), .B1(n8970), .B2(P2_U3152), .C1(
        n8969), .C2(n8980), .ZN(P2_U3329) );
  NAND2_X1 U10331 ( .A1(n6615), .A2(n8972), .ZN(n8974) );
  OAI211_X1 U10332 ( .C1(n8980), .C2(n8975), .A(n8974), .B(n8973), .ZN(
        P2_U3330) );
  INV_X1 U10333 ( .A(n6601), .ZN(n8978) );
  OAI222_X1 U10334 ( .A1(n8983), .A2(n8978), .B1(n8977), .B2(P2_U3152), .C1(
        n8976), .C2(n8980), .ZN(P2_U3331) );
  INV_X1 U10335 ( .A(n8979), .ZN(n9551) );
  OAI222_X1 U10336 ( .A1(n8983), .A2(n9551), .B1(P2_U3152), .B2(n8982), .C1(
        n8981), .C2(n8980), .ZN(P2_U3332) );
  INV_X1 U10337 ( .A(n8984), .ZN(n8985) );
  MUX2_X1 U10338 ( .A(n8985), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10339 ( .A(n8986), .ZN(n8988) );
  NOR2_X1 U10340 ( .A1(n8988), .A2(n8987), .ZN(n8989) );
  XNOR2_X1 U10341 ( .A(n8990), .B(n8989), .ZN(n8996) );
  AOI22_X1 U10342 ( .A1(n9252), .A2(n9120), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        n4476), .ZN(n8992) );
  NAND2_X1 U10343 ( .A1(n9223), .A2(n9103), .ZN(n8991) );
  OAI211_X1 U10344 ( .C1(n8993), .C2(n9117), .A(n8992), .B(n8991), .ZN(n8994)
         );
  AOI21_X1 U10345 ( .B1(n9415), .B2(n9095), .A(n8994), .ZN(n8995) );
  OAI21_X1 U10346 ( .B1(n8996), .B2(n9097), .A(n8995), .ZN(P1_U3212) );
  NAND2_X1 U10347 ( .A1(n8997), .A2(n8998), .ZN(n8999) );
  XOR2_X1 U10348 ( .A(n9000), .B(n8999), .Z(n9009) );
  OAI21_X1 U10349 ( .B1(n9105), .B2(n9002), .A(n9001), .ZN(n9006) );
  OAI22_X1 U10350 ( .A1(n9118), .A2(n9004), .B1(n9117), .B2(n9003), .ZN(n9005)
         );
  AOI211_X1 U10351 ( .C1(n9007), .C2(n9095), .A(n9006), .B(n9005), .ZN(n9008)
         );
  OAI21_X1 U10352 ( .B1(n9009), .B2(n9097), .A(n9008), .ZN(P1_U3213) );
  NAND2_X1 U10353 ( .A1(n9010), .A2(n9011), .ZN(n9012) );
  XOR2_X1 U10354 ( .A(n9013), .B(n9012), .Z(n9018) );
  OAI22_X1 U10355 ( .A1(n9313), .A2(n9105), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9014), .ZN(n9016) );
  OAI22_X1 U10356 ( .A1(n9038), .A2(n9117), .B1(n9118), .B2(n9287), .ZN(n9015)
         );
  AOI211_X1 U10357 ( .C1(n9286), .C2(n9095), .A(n9016), .B(n9015), .ZN(n9017)
         );
  OAI21_X1 U10358 ( .B1(n9018), .B2(n9097), .A(n9017), .ZN(P1_U3214) );
  INV_X1 U10359 ( .A(n9019), .ZN(n9020) );
  AOI21_X1 U10360 ( .B1(n9022), .B2(n9021), .A(n9020), .ZN(n9026) );
  AOI22_X1 U10361 ( .A1(n9120), .A2(n9367), .B1(n9344), .B2(n9103), .ZN(n9023)
         );
  NAND2_X1 U10362 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9169) );
  OAI211_X1 U10363 ( .C1(n9312), .C2(n9117), .A(n9023), .B(n9169), .ZN(n9024)
         );
  AOI21_X1 U10364 ( .B1(n9455), .B2(n9095), .A(n9024), .ZN(n9025) );
  OAI21_X1 U10365 ( .B1(n9026), .B2(n9097), .A(n9025), .ZN(P1_U3217) );
  XOR2_X1 U10366 ( .A(n9028), .B(n9027), .Z(n9033) );
  OAI22_X1 U10367 ( .A1(n9313), .A2(n9117), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9029), .ZN(n9031) );
  OAI22_X1 U10368 ( .A1(n9105), .A2(n9312), .B1(n9118), .B2(n9316), .ZN(n9030)
         );
  AOI211_X1 U10369 ( .C1(n9443), .C2(n9095), .A(n9031), .B(n9030), .ZN(n9032)
         );
  OAI21_X1 U10370 ( .B1(n9033), .B2(n9097), .A(n9032), .ZN(P1_U3221) );
  XOR2_X1 U10371 ( .A(n9035), .B(n9034), .Z(n9041) );
  NAND2_X1 U10372 ( .A1(n9252), .A2(n9108), .ZN(n9037) );
  AOI22_X1 U10373 ( .A1(n9247), .A2(n9103), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9036) );
  OAI211_X1 U10374 ( .C1(n9038), .C2(n9105), .A(n9037), .B(n9036), .ZN(n9039)
         );
  AOI21_X1 U10375 ( .B1(n9423), .B2(n9095), .A(n9039), .ZN(n9040) );
  OAI21_X1 U10376 ( .B1(n9041), .B2(n9097), .A(n9040), .ZN(P1_U3223) );
  INV_X1 U10377 ( .A(n9042), .ZN(n9043) );
  AOI21_X1 U10378 ( .B1(n9045), .B2(n9044), .A(n9043), .ZN(n9050) );
  NOR2_X1 U10379 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9046), .ZN(n9769) );
  OAI22_X1 U10380 ( .A1(n9118), .A2(n9391), .B1(n9117), .B2(n9092), .ZN(n9047)
         );
  AOI211_X1 U10381 ( .C1(n9120), .C2(n9381), .A(n9769), .B(n9047), .ZN(n9049)
         );
  NAND2_X1 U10382 ( .A1(n9390), .A2(n9095), .ZN(n9048) );
  OAI211_X1 U10383 ( .C1(n9050), .C2(n9097), .A(n9049), .B(n9048), .ZN(
        P1_U3224) );
  INV_X1 U10384 ( .A(n9465), .ZN(n9362) );
  OAI21_X1 U10385 ( .B1(n9053), .B2(n9052), .A(n9051), .ZN(n9054) );
  NAND2_X1 U10386 ( .A1(n9054), .A2(n9115), .ZN(n9057) );
  AND2_X1 U10387 ( .A1(n4476), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9780) );
  OAI22_X1 U10388 ( .A1(n9105), .A2(n9623), .B1(n9118), .B2(n9369), .ZN(n9055)
         );
  AOI211_X1 U10389 ( .C1(n9108), .C2(n9367), .A(n9780), .B(n9055), .ZN(n9056)
         );
  OAI211_X1 U10390 ( .C1(n9362), .C2(n9123), .A(n9057), .B(n9056), .ZN(
        P1_U3226) );
  INV_X1 U10391 ( .A(n9059), .ZN(n9060) );
  AOI21_X1 U10392 ( .B1(n9061), .B2(n9058), .A(n9060), .ZN(n9066) );
  NAND2_X1 U10393 ( .A1(n9267), .A2(n9108), .ZN(n9063) );
  AOI22_X1 U10394 ( .A1(n9303), .A2(n9120), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9062) );
  OAI211_X1 U10395 ( .C1(n9118), .C2(n9260), .A(n9063), .B(n9062), .ZN(n9064)
         );
  AOI21_X1 U10396 ( .B1(n9428), .B2(n9095), .A(n9064), .ZN(n9065) );
  OAI21_X1 U10397 ( .B1(n9066), .B2(n9097), .A(n9065), .ZN(P1_U3227) );
  INV_X1 U10398 ( .A(n9067), .ZN(n9072) );
  AOI21_X1 U10399 ( .B1(n9069), .B2(n9071), .A(n9068), .ZN(n9070) );
  AOI21_X1 U10400 ( .B1(n9072), .B2(n9071), .A(n9070), .ZN(n9077) );
  OAI22_X1 U10401 ( .A1(n9329), .A2(n9117), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9073), .ZN(n9075) );
  OAI22_X1 U10402 ( .A1(n9105), .A2(n9328), .B1(n9118), .B2(n9324), .ZN(n9074)
         );
  AOI211_X1 U10403 ( .C1(n9449), .C2(n9095), .A(n9075), .B(n9074), .ZN(n9076)
         );
  OAI21_X1 U10404 ( .B1(n9077), .B2(n9097), .A(n9076), .ZN(P1_U3231) );
  NAND2_X1 U10405 ( .A1(n9079), .A2(n9078), .ZN(n9080) );
  XOR2_X1 U10406 ( .A(n9081), .B(n9080), .Z(n9087) );
  OAI22_X1 U10407 ( .A1(n9105), .A2(n9329), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9082), .ZN(n9085) );
  OAI22_X1 U10408 ( .A1(n9083), .A2(n9117), .B1(n9118), .B2(n9296), .ZN(n9084)
         );
  AOI211_X1 U10409 ( .C1(n9438), .C2(n9095), .A(n9085), .B(n9084), .ZN(n9086)
         );
  OAI21_X1 U10410 ( .B1(n9087), .B2(n9097), .A(n9086), .ZN(P1_U3233) );
  NAND2_X1 U10411 ( .A1(n4504), .A2(n9088), .ZN(n9089) );
  XOR2_X1 U10412 ( .A(n9090), .B(n9089), .Z(n9098) );
  NAND2_X1 U10413 ( .A1(n4476), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9789) );
  OAI21_X1 U10414 ( .B1(n9117), .B2(n9328), .A(n9789), .ZN(n9094) );
  OAI22_X1 U10415 ( .A1(n9105), .A2(n9092), .B1(n9118), .B2(n9091), .ZN(n9093)
         );
  AOI211_X1 U10416 ( .C1(n9462), .C2(n9095), .A(n9094), .B(n9093), .ZN(n9096)
         );
  OAI21_X1 U10417 ( .B1(n9098), .B2(n9097), .A(n9096), .ZN(P1_U3236) );
  OAI211_X1 U10418 ( .C1(n9101), .C2(n9100), .A(n9099), .B(n9115), .ZN(n9110)
         );
  INV_X1 U10419 ( .A(n9102), .ZN(n9237) );
  AOI22_X1 U10420 ( .A1(n9237), .A2(n9103), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        n4476), .ZN(n9104) );
  OAI21_X1 U10421 ( .B1(n9106), .B2(n9105), .A(n9104), .ZN(n9107) );
  AOI21_X1 U10422 ( .B1(n9108), .B2(n9233), .A(n9107), .ZN(n9109) );
  OAI211_X1 U10423 ( .C1(n4765), .C2(n9123), .A(n9110), .B(n9109), .ZN(
        P1_U3238) );
  XNOR2_X1 U10424 ( .A(n9113), .B(n9112), .ZN(n9114) );
  XNOR2_X1 U10425 ( .A(n9111), .B(n9114), .ZN(n9116) );
  NAND2_X1 U10426 ( .A1(n9116), .A2(n9115), .ZN(n9122) );
  AND2_X1 U10427 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9758) );
  OAI22_X1 U10428 ( .A1(n9118), .A2(n9629), .B1(n9117), .B2(n9623), .ZN(n9119)
         );
  AOI211_X1 U10429 ( .C1(n9120), .C2(n9127), .A(n9758), .B(n9119), .ZN(n9121)
         );
  OAI211_X1 U10430 ( .C1(n9663), .C2(n9123), .A(n9122), .B(n9121), .ZN(
        P1_U3239) );
  MUX2_X1 U10431 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9124), .S(P1_U4006), .Z(
        P1_U3585) );
  INV_X1 U10432 ( .A(n9125), .ZN(n9200) );
  MUX2_X1 U10433 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9200), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10434 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9217), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10435 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9233), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10436 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9252), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10437 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9267), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10438 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9280), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10439 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9303), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10440 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9302), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10441 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9353), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10442 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9126), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10443 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9367), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10444 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9380), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10445 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9366), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10446 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9381), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10447 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9127), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10448 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9128), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10449 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9129), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10450 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9130), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10451 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9131), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10452 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9132), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10453 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9133), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10454 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9134), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10455 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9135), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10456 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9136), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10457 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9137), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10458 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n6701), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10459 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9138), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10460 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9139), .S(P1_U4006), .Z(
        P1_U3556) );
  MUX2_X1 U10461 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6696), .S(P1_U4006), .Z(
        P1_U3555) );
  NOR2_X1 U10462 ( .A1(n9140), .A2(n9152), .ZN(n9142) );
  NOR2_X1 U10463 ( .A1(n9142), .A2(n9141), .ZN(n9143) );
  NOR2_X1 U10464 ( .A1(n9143), .A2(n9153), .ZN(n9144) );
  XNOR2_X1 U10465 ( .A(n9143), .B(n9153), .ZN(n9756) );
  NOR2_X1 U10466 ( .A1(n9630), .A2(n9756), .ZN(n9755) );
  NOR2_X1 U10467 ( .A1(n9144), .A2(n9755), .ZN(n9767) );
  NAND2_X1 U10468 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9770), .ZN(n9145) );
  OAI21_X1 U10469 ( .B1(n9770), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9145), .ZN(
        n9766) );
  NOR2_X1 U10470 ( .A1(n9767), .A2(n9766), .ZN(n9765) );
  AOI21_X1 U10471 ( .B1(n9770), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9765), .ZN(
        n9778) );
  NAND2_X1 U10472 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9781), .ZN(n9146) );
  OAI21_X1 U10473 ( .B1(n9781), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9146), .ZN(
        n9777) );
  NOR2_X1 U10474 ( .A1(n9778), .A2(n9777), .ZN(n9776) );
  NOR2_X1 U10475 ( .A1(n9797), .A2(n9147), .ZN(n9148) );
  AOI21_X1 U10476 ( .B1(n9797), .B2(n9147), .A(n9148), .ZN(n9792) );
  NAND3_X1 U10477 ( .A1(n9166), .A2(n9150), .A3(n9149), .ZN(n9164) );
  XNOR2_X1 U10478 ( .A(n9797), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9800) );
  XNOR2_X1 U10479 ( .A(n9158), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9785) );
  INV_X1 U10480 ( .A(n9770), .ZN(n9156) );
  XNOR2_X1 U10481 ( .A(n9770), .B(n9476), .ZN(n9772) );
  AOI21_X1 U10482 ( .B1(n9152), .B2(n6349), .A(n9151), .ZN(n9154) );
  NAND2_X1 U10483 ( .A1(n9759), .A2(n9154), .ZN(n9155) );
  XNOR2_X1 U10484 ( .A(n9154), .B(n9153), .ZN(n9761) );
  NAND2_X1 U10485 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9761), .ZN(n9760) );
  NAND2_X1 U10486 ( .A1(n9155), .A2(n9760), .ZN(n9773) );
  NAND2_X1 U10487 ( .A1(n9772), .A2(n9773), .ZN(n9771) );
  OAI21_X1 U10488 ( .B1(n9156), .B2(n9476), .A(n9771), .ZN(n9784) );
  NAND2_X1 U10489 ( .A1(n9785), .A2(n9784), .ZN(n9782) );
  OAI21_X1 U10490 ( .B1(n9158), .B2(n9157), .A(n9782), .ZN(n9799) );
  NOR2_X1 U10491 ( .A1(n9800), .A2(n9799), .ZN(n9798) );
  AOI21_X1 U10492 ( .B1(n9160), .B2(n9159), .A(n9798), .ZN(n9162) );
  XOR2_X1 U10493 ( .A(n9162), .B(n9161), .Z(n9165) );
  AOI21_X1 U10494 ( .B1(n9165), .B2(n9783), .A(n9796), .ZN(n9163) );
  NAND2_X1 U10495 ( .A1(n9164), .A2(n9163), .ZN(n9168) );
  OAI22_X1 U10496 ( .A1(n9166), .A2(n9790), .B1(n9165), .B2(n9802), .ZN(n9167)
         );
  MUX2_X1 U10497 ( .A(n9168), .B(n9167), .S(n9331), .Z(n9171) );
  OAI21_X1 U10498 ( .B1(n9806), .B2(n4622), .A(n9169), .ZN(n9170) );
  NAND2_X1 U10499 ( .A1(n9496), .A2(n9179), .ZN(n9173) );
  XNOR2_X1 U10500 ( .A(n9172), .B(n9173), .ZN(n9400) );
  NAND2_X1 U10501 ( .A1(n9400), .A2(n9640), .ZN(n9178) );
  INV_X1 U10502 ( .A(n9403), .ZN(n9176) );
  NOR2_X1 U10503 ( .A1(n9176), .A2(n9399), .ZN(n9181) );
  AOI21_X1 U10504 ( .B1(n9399), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9181), .ZN(
        n9177) );
  OAI211_X1 U10505 ( .C1(n9654), .C2(n9172), .A(n9178), .B(n9177), .ZN(
        P1_U3261) );
  XNOR2_X1 U10506 ( .A(n9180), .B(n9179), .ZN(n9404) );
  NAND2_X1 U10507 ( .A1(n9404), .A2(n9640), .ZN(n9183) );
  AOI21_X1 U10508 ( .B1(n9399), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9181), .ZN(
        n9182) );
  OAI211_X1 U10509 ( .C1(n9496), .C2(n9654), .A(n9183), .B(n9182), .ZN(
        P1_U3262) );
  INV_X1 U10510 ( .A(n9184), .ZN(n9193) );
  NAND2_X1 U10511 ( .A1(n9185), .A2(n9395), .ZN(n9188) );
  AOI22_X1 U10512 ( .A1(n9186), .A2(n9343), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9399), .ZN(n9187) );
  OAI211_X1 U10513 ( .C1(n9189), .C2(n9654), .A(n9188), .B(n9187), .ZN(n9190)
         );
  AOI21_X1 U10514 ( .B1(n9191), .B2(n9660), .A(n9190), .ZN(n9192) );
  OAI21_X1 U10515 ( .B1(n9193), .B2(n9373), .A(n9192), .ZN(P1_U3355) );
  INV_X1 U10516 ( .A(n9410), .ZN(n9212) );
  OAI211_X1 U10517 ( .C1(n9199), .C2(n9198), .A(n9197), .B(n9649), .ZN(n9202)
         );
  AOI22_X1 U10518 ( .A1(n9200), .A2(n9379), .B1(n9233), .B2(n9382), .ZN(n9201)
         );
  NAND2_X1 U10519 ( .A1(n9202), .A2(n9201), .ZN(n9408) );
  NAND2_X1 U10520 ( .A1(n9203), .A2(n9221), .ZN(n9204) );
  NAND2_X1 U10521 ( .A1(n9204), .A2(n9467), .ZN(n9205) );
  NOR2_X1 U10522 ( .A1(n9206), .A2(n9205), .ZN(n9407) );
  NAND2_X1 U10523 ( .A1(n9407), .A2(n9395), .ZN(n9209) );
  AOI22_X1 U10524 ( .A1(n9207), .A2(n9343), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9399), .ZN(n9208) );
  OAI211_X1 U10525 ( .C1(n4761), .C2(n9654), .A(n9209), .B(n9208), .ZN(n9210)
         );
  AOI21_X1 U10526 ( .B1(n9408), .B2(n9660), .A(n9210), .ZN(n9211) );
  OAI21_X1 U10527 ( .B1(n9212), .B2(n9373), .A(n9211), .ZN(P1_U3263) );
  XOR2_X1 U10528 ( .A(n9215), .B(n9213), .Z(n9417) );
  OAI211_X1 U10529 ( .C1(n9216), .C2(n9215), .A(n9214), .B(n9649), .ZN(n9219)
         );
  AOI22_X1 U10530 ( .A1(n9217), .A2(n9379), .B1(n9382), .B2(n9252), .ZN(n9218)
         );
  NAND2_X1 U10531 ( .A1(n9219), .A2(n9218), .ZN(n9413) );
  INV_X1 U10532 ( .A(n9221), .ZN(n9222) );
  AOI211_X1 U10533 ( .C1(n9415), .C2(n4766), .A(n9827), .B(n9222), .ZN(n9414)
         );
  NAND2_X1 U10534 ( .A1(n9414), .A2(n9395), .ZN(n9225) );
  AOI22_X1 U10535 ( .A1(n9223), .A2(n9343), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9399), .ZN(n9224) );
  OAI211_X1 U10536 ( .C1(n6772), .C2(n9654), .A(n9225), .B(n9224), .ZN(n9226)
         );
  AOI21_X1 U10537 ( .B1(n9413), .B2(n9660), .A(n9226), .ZN(n9227) );
  OAI21_X1 U10538 ( .B1(n9417), .B2(n9373), .A(n9227), .ZN(P1_U3264) );
  XOR2_X1 U10539 ( .A(n9229), .B(n9228), .Z(n9420) );
  INV_X1 U10540 ( .A(n9420), .ZN(n9242) );
  INV_X1 U10541 ( .A(n9229), .ZN(n9230) );
  XNOR2_X1 U10542 ( .A(n9231), .B(n9230), .ZN(n9232) );
  NAND2_X1 U10543 ( .A1(n9232), .A2(n9649), .ZN(n9235) );
  AOI22_X1 U10544 ( .A1(n9233), .A2(n9379), .B1(n9382), .B2(n9267), .ZN(n9234)
         );
  NAND2_X1 U10545 ( .A1(n9235), .A2(n9234), .ZN(n9418) );
  AOI211_X1 U10546 ( .C1(n9236), .C2(n9244), .A(n9827), .B(n9220), .ZN(n9419)
         );
  NAND2_X1 U10547 ( .A1(n9419), .A2(n9395), .ZN(n9239) );
  AOI22_X1 U10548 ( .A1(n9237), .A2(n9343), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9399), .ZN(n9238) );
  OAI211_X1 U10549 ( .C1(n4765), .C2(n9654), .A(n9239), .B(n9238), .ZN(n9240)
         );
  AOI21_X1 U10550 ( .B1(n9660), .B2(n9418), .A(n9240), .ZN(n9241) );
  OAI21_X1 U10551 ( .B1(n9242), .B2(n9373), .A(n9241), .ZN(P1_U3265) );
  XOR2_X1 U10552 ( .A(n9243), .B(n9251), .Z(n9427) );
  INV_X1 U10553 ( .A(n9259), .ZN(n9246) );
  INV_X1 U10554 ( .A(n9244), .ZN(n9245) );
  AOI21_X1 U10555 ( .B1(n9423), .B2(n9246), .A(n9245), .ZN(n9424) );
  AOI22_X1 U10556 ( .A1(n9247), .A2(n9343), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9399), .ZN(n9248) );
  OAI21_X1 U10557 ( .B1(n9249), .B2(n9654), .A(n9248), .ZN(n9255) );
  XOR2_X1 U10558 ( .A(n9251), .B(n9250), .Z(n9253) );
  AOI222_X1 U10559 ( .A1(n9649), .A2(n9253), .B1(n9252), .B2(n9379), .C1(n9280), .C2(n9382), .ZN(n9426) );
  NOR2_X1 U10560 ( .A1(n9426), .A2(n9399), .ZN(n9254) );
  AOI211_X1 U10561 ( .C1(n9424), .C2(n9640), .A(n9255), .B(n9254), .ZN(n9256)
         );
  OAI21_X1 U10562 ( .B1(n9427), .B2(n9373), .A(n9256), .ZN(P1_U3266) );
  XNOR2_X1 U10563 ( .A(n9257), .B(n9258), .ZN(n9432) );
  AOI21_X1 U10564 ( .B1(n9428), .B2(n9283), .A(n9259), .ZN(n9429) );
  INV_X1 U10565 ( .A(n9428), .ZN(n9263) );
  INV_X1 U10566 ( .A(n9260), .ZN(n9261) );
  AOI22_X1 U10567 ( .A1(n9261), .A2(n9343), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9399), .ZN(n9262) );
  OAI21_X1 U10568 ( .B1(n9263), .B2(n9654), .A(n9262), .ZN(n9270) );
  OAI21_X1 U10569 ( .B1(n9266), .B2(n9265), .A(n9264), .ZN(n9268) );
  AOI222_X1 U10570 ( .A1(n9649), .A2(n9268), .B1(n9267), .B2(n9379), .C1(n9303), .C2(n9382), .ZN(n9431) );
  NOR2_X1 U10571 ( .A1(n9431), .A2(n9399), .ZN(n9269) );
  AOI211_X1 U10572 ( .C1(n9429), .C2(n9640), .A(n9270), .B(n9269), .ZN(n9271)
         );
  OAI21_X1 U10573 ( .B1(n9432), .B2(n9373), .A(n9271), .ZN(P1_U3267) );
  XOR2_X1 U10574 ( .A(n9275), .B(n9272), .Z(n9435) );
  INV_X1 U10575 ( .A(n9435), .ZN(n9293) );
  NAND2_X1 U10576 ( .A1(n9274), .A2(n9273), .ZN(n9277) );
  INV_X1 U10577 ( .A(n9275), .ZN(n9276) );
  XNOR2_X1 U10578 ( .A(n9277), .B(n9276), .ZN(n9278) );
  NAND2_X1 U10579 ( .A1(n9278), .A2(n9649), .ZN(n9282) );
  AOI22_X1 U10580 ( .A1(n9280), .A2(n9379), .B1(n9382), .B2(n9279), .ZN(n9281)
         );
  NAND2_X1 U10581 ( .A1(n9282), .A2(n9281), .ZN(n9433) );
  INV_X1 U10582 ( .A(n9295), .ZN(n9285) );
  INV_X1 U10583 ( .A(n9283), .ZN(n9284) );
  AOI211_X1 U10584 ( .C1(n9286), .C2(n9285), .A(n9827), .B(n9284), .ZN(n9434)
         );
  NAND2_X1 U10585 ( .A1(n9434), .A2(n9395), .ZN(n9290) );
  INV_X1 U10586 ( .A(n9287), .ZN(n9288) );
  AOI22_X1 U10587 ( .A1(n9288), .A2(n9343), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9399), .ZN(n9289) );
  OAI211_X1 U10588 ( .C1(n9509), .C2(n9654), .A(n9290), .B(n9289), .ZN(n9291)
         );
  AOI21_X1 U10589 ( .B1(n9433), .B2(n9660), .A(n9291), .ZN(n9292) );
  OAI21_X1 U10590 ( .B1(n9293), .B2(n9373), .A(n9292), .ZN(P1_U3268) );
  XNOR2_X1 U10591 ( .A(n9294), .B(n9301), .ZN(n9442) );
  AOI21_X1 U10592 ( .B1(n9438), .B2(n9314), .A(n9295), .ZN(n9439) );
  AND2_X1 U10593 ( .A1(n9438), .A2(n9334), .ZN(n9299) );
  INV_X1 U10594 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9297) );
  OAI22_X1 U10595 ( .A1(n9297), .A2(n9660), .B1(n9296), .B2(n9655), .ZN(n9298)
         );
  AOI211_X1 U10596 ( .C1(n9439), .C2(n9640), .A(n9299), .B(n9298), .ZN(n9306)
         );
  XOR2_X1 U10597 ( .A(n9301), .B(n9300), .Z(n9304) );
  AOI222_X1 U10598 ( .A1(n9649), .A2(n9304), .B1(n9303), .B2(n9379), .C1(n9302), .C2(n9382), .ZN(n9441) );
  OR2_X1 U10599 ( .A1(n9441), .A2(n9399), .ZN(n9305) );
  OAI211_X1 U10600 ( .C1(n9442), .C2(n9373), .A(n9306), .B(n9305), .ZN(
        P1_U3269) );
  XNOR2_X1 U10601 ( .A(n9307), .B(n9308), .ZN(n9446) );
  INV_X1 U10602 ( .A(n9446), .ZN(n9322) );
  AOI22_X1 U10603 ( .A1(n9443), .A2(n9334), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9399), .ZN(n9321) );
  XNOR2_X1 U10604 ( .A(n9310), .B(n9309), .ZN(n9311) );
  OAI222_X1 U10605 ( .A1(n9646), .A2(n9313), .B1(n9644), .B2(n9312), .C1(n9311), .C2(n9326), .ZN(n9444) );
  INV_X1 U10606 ( .A(n9314), .ZN(n9315) );
  AOI211_X1 U10607 ( .C1(n9443), .C2(n4573), .A(n9827), .B(n9315), .ZN(n9445)
         );
  INV_X1 U10608 ( .A(n9445), .ZN(n9318) );
  OAI22_X1 U10609 ( .A1(n9318), .A2(n9317), .B1(n9655), .B2(n9316), .ZN(n9319)
         );
  OAI21_X1 U10610 ( .B1(n9444), .B2(n9319), .A(n9660), .ZN(n9320) );
  OAI211_X1 U10611 ( .C1(n9322), .C2(n9373), .A(n9321), .B(n9320), .ZN(
        P1_U3270) );
  AOI21_X1 U10612 ( .B1(n9340), .B2(n9449), .A(n9827), .ZN(n9323) );
  AND2_X1 U10613 ( .A1(n9323), .A2(n4573), .ZN(n9451) );
  NOR2_X1 U10614 ( .A1(n9324), .A2(n9655), .ZN(n9330) );
  XOR2_X1 U10615 ( .A(n9333), .B(n9325), .Z(n9327) );
  OAI222_X1 U10616 ( .A1(n9646), .A2(n9329), .B1(n9644), .B2(n9328), .C1(n9327), .C2(n9326), .ZN(n9450) );
  AOI211_X1 U10617 ( .C1(n9451), .C2(n9331), .A(n9330), .B(n9450), .ZN(n9337)
         );
  XNOR2_X1 U10618 ( .A(n9332), .B(n9333), .ZN(n9452) );
  NAND2_X1 U10619 ( .A1(n9452), .A2(n9387), .ZN(n9336) );
  AOI22_X1 U10620 ( .A1(n9449), .A2(n9334), .B1(n9399), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n9335) );
  OAI211_X1 U10621 ( .C1(n9399), .C2(n9337), .A(n9336), .B(n9335), .ZN(
        P1_U3271) );
  XOR2_X1 U10622 ( .A(n9338), .B(n9347), .Z(n9459) );
  INV_X1 U10623 ( .A(n9339), .ZN(n9342) );
  INV_X1 U10624 ( .A(n9340), .ZN(n9341) );
  AOI21_X1 U10625 ( .B1(n9455), .B2(n9342), .A(n9341), .ZN(n9456) );
  AOI22_X1 U10626 ( .A1(n9399), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9344), .B2(
        n9343), .ZN(n9345) );
  OAI21_X1 U10627 ( .B1(n9346), .B2(n9654), .A(n9345), .ZN(n9356) );
  INV_X1 U10628 ( .A(n9347), .ZN(n9348) );
  NAND3_X1 U10629 ( .A1(n9350), .A2(n9349), .A3(n9348), .ZN(n9351) );
  NAND2_X1 U10630 ( .A1(n9352), .A2(n9351), .ZN(n9354) );
  AOI222_X1 U10631 ( .A1(n9649), .A2(n9354), .B1(n9353), .B2(n9379), .C1(n9367), .C2(n9382), .ZN(n9458) );
  NOR2_X1 U10632 ( .A1(n9458), .A2(n9399), .ZN(n9355) );
  AOI211_X1 U10633 ( .C1(n9456), .C2(n9640), .A(n9356), .B(n9355), .ZN(n9357)
         );
  OAI21_X1 U10634 ( .B1(n9459), .B2(n9373), .A(n9357), .ZN(P1_U3272) );
  XNOR2_X1 U10635 ( .A(n9358), .B(n9359), .ZN(n9472) );
  AOI21_X1 U10636 ( .B1(n9465), .B2(n9388), .A(n9360), .ZN(n9468) );
  OAI22_X1 U10637 ( .A1(n9362), .A2(n9654), .B1(n9660), .B2(n9361), .ZN(n9363)
         );
  AOI21_X1 U10638 ( .B1(n9468), .B2(n9640), .A(n9363), .ZN(n9372) );
  XNOR2_X1 U10639 ( .A(n9365), .B(n9364), .ZN(n9368) );
  AOI222_X1 U10640 ( .A1(n9649), .A2(n9368), .B1(n9367), .B2(n9379), .C1(n9366), .C2(n9382), .ZN(n9470) );
  OAI21_X1 U10641 ( .B1(n9369), .B2(n9655), .A(n9470), .ZN(n9370) );
  NAND2_X1 U10642 ( .A1(n9370), .A2(n9660), .ZN(n9371) );
  OAI211_X1 U10643 ( .C1(n9472), .C2(n9373), .A(n9372), .B(n9371), .ZN(
        P1_U3274) );
  NAND2_X1 U10644 ( .A1(n9375), .A2(n9374), .ZN(n9377) );
  XNOR2_X1 U10645 ( .A(n9377), .B(n9376), .ZN(n9378) );
  NAND2_X1 U10646 ( .A1(n9378), .A2(n9649), .ZN(n9384) );
  AOI22_X1 U10647 ( .A1(n9382), .A2(n9381), .B1(n9380), .B2(n9379), .ZN(n9383)
         );
  NAND2_X1 U10648 ( .A1(n9384), .A2(n9383), .ZN(n9473) );
  INV_X1 U10649 ( .A(n9473), .ZN(n9398) );
  XNOR2_X1 U10650 ( .A(n9386), .B(n9385), .ZN(n9475) );
  NAND2_X1 U10651 ( .A1(n9475), .A2(n9387), .ZN(n9397) );
  INV_X1 U10652 ( .A(n9388), .ZN(n9389) );
  AOI211_X1 U10653 ( .C1(n9390), .C2(n9618), .A(n9827), .B(n9389), .ZN(n9474)
         );
  INV_X1 U10654 ( .A(n9390), .ZN(n9524) );
  NOR2_X1 U10655 ( .A1(n9524), .A2(n9654), .ZN(n9394) );
  OAI22_X1 U10656 ( .A1(n9660), .A2(n9392), .B1(n9391), .B2(n9655), .ZN(n9393)
         );
  AOI211_X1 U10657 ( .C1(n9474), .C2(n9395), .A(n9394), .B(n9393), .ZN(n9396)
         );
  OAI211_X1 U10658 ( .C1(n9399), .C2(n9398), .A(n9397), .B(n9396), .ZN(
        P1_U3275) );
  AOI21_X1 U10659 ( .B1(n9400), .B2(n9467), .A(n9403), .ZN(n9490) );
  MUX2_X1 U10660 ( .A(n9401), .B(n9490), .S(n9840), .Z(n9402) );
  OAI21_X1 U10661 ( .B1(n9486), .B2(n9172), .A(n9402), .ZN(P1_U3554) );
  AOI21_X1 U10662 ( .B1(n9404), .B2(n9467), .A(n9403), .ZN(n9493) );
  MUX2_X1 U10663 ( .A(n9405), .B(n9493), .S(n9840), .Z(n9406) );
  OAI21_X1 U10664 ( .B1(n9496), .B2(n9486), .A(n9406), .ZN(P1_U3553) );
  MUX2_X1 U10665 ( .A(n9411), .B(n9497), .S(n9840), .Z(n9412) );
  OAI21_X1 U10666 ( .B1(n4761), .B2(n9486), .A(n9412), .ZN(P1_U3551) );
  AOI211_X1 U10667 ( .C1(n9466), .C2(n9415), .A(n9414), .B(n9413), .ZN(n9416)
         );
  OAI21_X1 U10668 ( .B1(n9417), .B2(n9471), .A(n9416), .ZN(n9500) );
  MUX2_X1 U10669 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9500), .S(n9840), .Z(
        P1_U3550) );
  AOI211_X1 U10670 ( .C1(n9420), .C2(n9822), .A(n9419), .B(n9418), .ZN(n9501)
         );
  MUX2_X1 U10671 ( .A(n9421), .B(n9501), .S(n9840), .Z(n9422) );
  OAI21_X1 U10672 ( .B1(n4765), .B2(n9486), .A(n9422), .ZN(P1_U3549) );
  AOI22_X1 U10673 ( .A1(n9424), .A2(n9467), .B1(n9466), .B2(n9423), .ZN(n9425)
         );
  OAI211_X1 U10674 ( .C1(n9427), .C2(n9471), .A(n9426), .B(n9425), .ZN(n9504)
         );
  MUX2_X1 U10675 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9504), .S(n9840), .Z(
        P1_U3548) );
  AOI22_X1 U10676 ( .A1(n9429), .A2(n9467), .B1(n9466), .B2(n9428), .ZN(n9430)
         );
  OAI211_X1 U10677 ( .C1(n9432), .C2(n9471), .A(n9431), .B(n9430), .ZN(n9505)
         );
  MUX2_X1 U10678 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9505), .S(n9840), .Z(
        P1_U3547) );
  AOI211_X1 U10679 ( .C1(n9435), .C2(n9822), .A(n9434), .B(n9433), .ZN(n9506)
         );
  MUX2_X1 U10680 ( .A(n9436), .B(n9506), .S(n9840), .Z(n9437) );
  OAI21_X1 U10681 ( .B1(n9509), .B2(n9486), .A(n9437), .ZN(P1_U3546) );
  AOI22_X1 U10682 ( .A1(n9439), .A2(n9467), .B1(n9466), .B2(n9438), .ZN(n9440)
         );
  OAI211_X1 U10683 ( .C1(n9442), .C2(n9471), .A(n9441), .B(n9440), .ZN(n9510)
         );
  MUX2_X1 U10684 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9510), .S(n9840), .Z(
        P1_U3545) );
  INV_X1 U10685 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9447) );
  AOI211_X1 U10686 ( .C1(n9446), .C2(n9822), .A(n9445), .B(n9444), .ZN(n9511)
         );
  MUX2_X1 U10687 ( .A(n9447), .B(n9511), .S(n9840), .Z(n9448) );
  OAI21_X1 U10688 ( .B1(n6771), .B2(n9486), .A(n9448), .ZN(P1_U3544) );
  INV_X1 U10689 ( .A(n9449), .ZN(n9517) );
  AOI211_X1 U10690 ( .C1(n9452), .C2(n9822), .A(n9451), .B(n9450), .ZN(n9514)
         );
  MUX2_X1 U10691 ( .A(n9453), .B(n9514), .S(n9840), .Z(n9454) );
  OAI21_X1 U10692 ( .B1(n9517), .B2(n9486), .A(n9454), .ZN(P1_U3543) );
  AOI22_X1 U10693 ( .A1(n9456), .A2(n9467), .B1(n9466), .B2(n9455), .ZN(n9457)
         );
  OAI211_X1 U10694 ( .C1(n9459), .C2(n9471), .A(n9458), .B(n9457), .ZN(n9518)
         );
  MUX2_X1 U10695 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9518), .S(n9840), .Z(
        P1_U3542) );
  AOI211_X1 U10696 ( .C1(n9466), .C2(n9462), .A(n9461), .B(n9460), .ZN(n9463)
         );
  OAI21_X1 U10697 ( .B1(n9464), .B2(n9471), .A(n9463), .ZN(n9519) );
  MUX2_X1 U10698 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9519), .S(n9840), .Z(
        P1_U3541) );
  AOI22_X1 U10699 ( .A1(n9468), .A2(n9467), .B1(n9466), .B2(n9465), .ZN(n9469)
         );
  OAI211_X1 U10700 ( .C1(n9472), .C2(n9471), .A(n9470), .B(n9469), .ZN(n9520)
         );
  MUX2_X1 U10701 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9520), .S(n9840), .Z(
        P1_U3540) );
  AOI211_X1 U10702 ( .C1(n9475), .C2(n9822), .A(n9474), .B(n9473), .ZN(n9521)
         );
  MUX2_X1 U10703 ( .A(n9476), .B(n9521), .S(n9840), .Z(n9477) );
  OAI21_X1 U10704 ( .B1(n9524), .B2(n9486), .A(n9477), .ZN(P1_U3539) );
  AOI211_X1 U10705 ( .C1(n9480), .C2(n9822), .A(n9479), .B(n9478), .ZN(n9525)
         );
  MUX2_X1 U10706 ( .A(n6349), .B(n9525), .S(n9840), .Z(n9481) );
  OAI21_X1 U10707 ( .B1(n9528), .B2(n9486), .A(n9481), .ZN(P1_U3537) );
  AOI211_X1 U10708 ( .C1(n9484), .C2(n9822), .A(n9483), .B(n9482), .ZN(n9529)
         );
  MUX2_X1 U10709 ( .A(n7706), .B(n9529), .S(n9840), .Z(n9485) );
  OAI21_X1 U10710 ( .B1(n9533), .B2(n9486), .A(n9485), .ZN(P1_U3535) );
  OAI21_X1 U10711 ( .B1(n9489), .B2(n9488), .A(n9487), .ZN(n9534) );
  MUX2_X1 U10712 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9534), .S(n9840), .Z(
        P1_U3523) );
  MUX2_X1 U10713 ( .A(n9491), .B(n9490), .S(n9835), .Z(n9492) );
  OAI21_X1 U10714 ( .B1(n9532), .B2(n9172), .A(n9492), .ZN(P1_U3522) );
  MUX2_X1 U10715 ( .A(n9494), .B(n9493), .S(n9835), .Z(n9495) );
  OAI21_X1 U10716 ( .B1(n9496), .B2(n9532), .A(n9495), .ZN(P1_U3521) );
  INV_X1 U10717 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9498) );
  MUX2_X1 U10718 ( .A(n9498), .B(n9497), .S(n9835), .Z(n9499) );
  OAI21_X1 U10719 ( .B1(n4761), .B2(n9532), .A(n9499), .ZN(P1_U3519) );
  MUX2_X1 U10720 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9500), .S(n9835), .Z(
        P1_U3518) );
  INV_X1 U10721 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9502) );
  MUX2_X1 U10722 ( .A(n9502), .B(n9501), .S(n9835), .Z(n9503) );
  OAI21_X1 U10723 ( .B1(n4765), .B2(n9532), .A(n9503), .ZN(P1_U3517) );
  MUX2_X1 U10724 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9504), .S(n9835), .Z(
        P1_U3516) );
  MUX2_X1 U10725 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9505), .S(n9835), .Z(
        P1_U3515) );
  INV_X1 U10726 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9507) );
  MUX2_X1 U10727 ( .A(n9507), .B(n9506), .S(n9835), .Z(n9508) );
  OAI21_X1 U10728 ( .B1(n9509), .B2(n9532), .A(n9508), .ZN(P1_U3514) );
  MUX2_X1 U10729 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9510), .S(n9835), .Z(
        P1_U3513) );
  INV_X1 U10730 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9512) );
  MUX2_X1 U10731 ( .A(n9512), .B(n9511), .S(n9835), .Z(n9513) );
  OAI21_X1 U10732 ( .B1(n6771), .B2(n9532), .A(n9513), .ZN(P1_U3512) );
  INV_X1 U10733 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9515) );
  MUX2_X1 U10734 ( .A(n9515), .B(n9514), .S(n9835), .Z(n9516) );
  OAI21_X1 U10735 ( .B1(n9517), .B2(n9532), .A(n9516), .ZN(P1_U3511) );
  MUX2_X1 U10736 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9518), .S(n9835), .Z(
        P1_U3510) );
  MUX2_X1 U10737 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9519), .S(n9835), .Z(
        P1_U3508) );
  MUX2_X1 U10738 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9520), .S(n9835), .Z(
        P1_U3505) );
  INV_X1 U10739 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9522) );
  MUX2_X1 U10740 ( .A(n9522), .B(n9521), .S(n9835), .Z(n9523) );
  OAI21_X1 U10741 ( .B1(n9524), .B2(n9532), .A(n9523), .ZN(P1_U3502) );
  INV_X1 U10742 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9526) );
  MUX2_X1 U10743 ( .A(n9526), .B(n9525), .S(n9835), .Z(n9527) );
  OAI21_X1 U10744 ( .B1(n9528), .B2(n9532), .A(n9527), .ZN(P1_U3496) );
  INV_X1 U10745 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9530) );
  MUX2_X1 U10746 ( .A(n9530), .B(n9529), .S(n9835), .Z(n9531) );
  OAI21_X1 U10747 ( .B1(n9533), .B2(n9532), .A(n9531), .ZN(P1_U3490) );
  MUX2_X1 U10748 ( .A(P1_REG0_REG_0__SCAN_IN), .B(n9534), .S(n9835), .Z(
        P1_U3454) );
  MUX2_X1 U10749 ( .A(P1_D_REG_1__SCAN_IN), .B(n9535), .S(n9808), .Z(P1_U3441)
         );
  NOR4_X1 U10750 ( .A1(n9537), .A2(P1_IR_REG_30__SCAN_IN), .A3(n4476), .A4(
        n9536), .ZN(n9538) );
  AOI21_X1 U10751 ( .B1(n9539), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9538), .ZN(
        n9540) );
  OAI21_X1 U10752 ( .B1(n9541), .B2(n8089), .A(n9540), .ZN(P1_U3322) );
  OAI222_X1 U10753 ( .A1(n9544), .A2(n10089), .B1(n8089), .B2(n9543), .C1(
        P1_U3084), .C2(n9542), .ZN(P1_U3323) );
  NAND2_X1 U10754 ( .A1(n6601), .A2(n9545), .ZN(n9547) );
  OAI211_X1 U10755 ( .C1(n9549), .C2(n9548), .A(n9547), .B(n9546), .ZN(
        P1_U3326) );
  INV_X1 U10756 ( .A(n9553), .ZN(n9554) );
  AOI21_X1 U10757 ( .B1(n9899), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n9554), .ZN(
        n9565) );
  NAND2_X1 U10758 ( .A1(n9905), .A2(n9555), .ZN(n9564) );
  OAI211_X1 U10759 ( .C1(n9558), .C2(n9557), .A(n9906), .B(n9556), .ZN(n9563)
         );
  OAI211_X1 U10760 ( .C1(n9561), .C2(n9560), .A(n9901), .B(n9559), .ZN(n9562)
         );
  NAND4_X1 U10761 ( .A1(n9565), .A2(n9564), .A3(n9563), .A4(n9562), .ZN(
        P2_U3250) );
  INV_X1 U10762 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10041) );
  OAI22_X1 U10763 ( .A1(n9566), .A2(n10041), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7139), .ZN(n9567) );
  AOI21_X1 U10764 ( .B1(n9905), .B2(n9568), .A(n9567), .ZN(n9577) );
  AND2_X1 U10765 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9571) );
  OAI211_X1 U10766 ( .C1(n9571), .C2(n9570), .A(n9901), .B(n9569), .ZN(n9576)
         );
  AND2_X1 U10767 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9574) );
  OAI211_X1 U10768 ( .C1(n9574), .C2(n9573), .A(n9906), .B(n9572), .ZN(n9575)
         );
  NAND3_X1 U10769 ( .A1(n9577), .A2(n9576), .A3(n9575), .ZN(P2_U3246) );
  AOI22_X1 U10770 ( .A1(n9899), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9588) );
  NAND2_X1 U10771 ( .A1(n9905), .A2(n9578), .ZN(n9587) );
  OAI211_X1 U10772 ( .C1(n9581), .C2(n9580), .A(n9901), .B(n9579), .ZN(n9586)
         );
  OAI211_X1 U10773 ( .C1(n9584), .C2(n9583), .A(n9906), .B(n9582), .ZN(n9585)
         );
  NAND4_X1 U10774 ( .A1(n9588), .A2(n9587), .A3(n9586), .A4(n9585), .ZN(
        P2_U3247) );
  OAI21_X1 U10775 ( .B1(n9590), .B2(n9826), .A(n9589), .ZN(n9591) );
  AOI211_X1 U10776 ( .C1(n9593), .C2(n9822), .A(n9592), .B(n9591), .ZN(n9595)
         );
  INV_X1 U10777 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9594) );
  AOI22_X1 U10778 ( .A1(n9835), .A2(n9595), .B1(n9594), .B2(n9833), .ZN(
        P1_U3484) );
  AOI22_X1 U10779 ( .A1(n9840), .A2(n9595), .B1(n6266), .B2(n9838), .ZN(
        P1_U3533) );
  AOI22_X1 U10780 ( .A1(n9606), .A2(n9596), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3152), .ZN(n9603) );
  OAI21_X1 U10781 ( .B1(n9599), .B2(n9598), .A(n9597), .ZN(n9601) );
  AOI22_X1 U10782 ( .A1(n9601), .A2(n9611), .B1(n9610), .B2(n9600), .ZN(n9602)
         );
  OAI211_X1 U10783 ( .C1(n9616), .C2(n9604), .A(n9603), .B(n9602), .ZN(
        P2_U3217) );
  AOI22_X1 U10784 ( .A1(n9606), .A2(n9605), .B1(P2_REG3_REG_15__SCAN_IN), .B2(
        P2_U3152), .ZN(n9614) );
  XNOR2_X1 U10785 ( .A(n9608), .B(n9607), .ZN(n9612) );
  AOI22_X1 U10786 ( .A1(n9612), .A2(n9611), .B1(n9610), .B2(n9609), .ZN(n9613)
         );
  OAI211_X1 U10787 ( .C1(n9616), .C2(n9615), .A(n9614), .B(n9613), .ZN(
        P2_U3243) );
  XOR2_X1 U10788 ( .A(n9617), .B(n9622), .Z(n9628) );
  INV_X1 U10789 ( .A(n9628), .ZN(n9667) );
  OAI21_X1 U10790 ( .B1(n9619), .B2(n9663), .A(n9618), .ZN(n9664) );
  INV_X1 U10791 ( .A(n9664), .ZN(n9620) );
  AOI22_X1 U10792 ( .A1(n9667), .A2(n9641), .B1(n9640), .B2(n9620), .ZN(n9634)
         );
  XOR2_X1 U10793 ( .A(n9622), .B(n9621), .Z(n9626) );
  OAI22_X1 U10794 ( .A1(n9624), .A2(n9644), .B1(n9623), .B2(n9646), .ZN(n9625)
         );
  AOI21_X1 U10795 ( .B1(n9626), .B2(n9649), .A(n9625), .ZN(n9627) );
  OAI21_X1 U10796 ( .B1(n9628), .B2(n9652), .A(n9627), .ZN(n9665) );
  NOR2_X1 U10797 ( .A1(n9663), .A2(n9654), .ZN(n9632) );
  OAI22_X1 U10798 ( .A1(n9660), .A2(n9630), .B1(n9629), .B2(n9655), .ZN(n9631)
         );
  AOI211_X1 U10799 ( .C1(n9665), .C2(n9660), .A(n9632), .B(n9631), .ZN(n9633)
         );
  NAND2_X1 U10800 ( .A1(n9634), .A2(n9633), .ZN(P1_U3276) );
  XOR2_X1 U10801 ( .A(n9635), .B(n9642), .Z(n9653) );
  INV_X1 U10802 ( .A(n9653), .ZN(n9677) );
  OR2_X1 U10803 ( .A1(n9636), .A2(n9673), .ZN(n9637) );
  NAND2_X1 U10804 ( .A1(n9638), .A2(n9637), .ZN(n9674) );
  INV_X1 U10805 ( .A(n9674), .ZN(n9639) );
  AOI22_X1 U10806 ( .A1(n9677), .A2(n9641), .B1(n9640), .B2(n9639), .ZN(n9662)
         );
  XNOR2_X1 U10807 ( .A(n9643), .B(n9642), .ZN(n9650) );
  OAI22_X1 U10808 ( .A1(n9647), .A2(n9646), .B1(n9645), .B2(n9644), .ZN(n9648)
         );
  AOI21_X1 U10809 ( .B1(n9650), .B2(n9649), .A(n9648), .ZN(n9651) );
  OAI21_X1 U10810 ( .B1(n9653), .B2(n9652), .A(n9651), .ZN(n9675) );
  NOR2_X1 U10811 ( .A1(n9673), .A2(n9654), .ZN(n9659) );
  OAI22_X1 U10812 ( .A1(n9660), .A2(n9657), .B1(n9656), .B2(n9655), .ZN(n9658)
         );
  AOI211_X1 U10813 ( .C1(n9675), .C2(n9660), .A(n9659), .B(n9658), .ZN(n9661)
         );
  NAND2_X1 U10814 ( .A1(n9662), .A2(n9661), .ZN(P1_U3280) );
  OAI22_X1 U10815 ( .A1(n9664), .A2(n9827), .B1(n9663), .B2(n9826), .ZN(n9666)
         );
  AOI211_X1 U10816 ( .C1(n9832), .C2(n9667), .A(n9666), .B(n9665), .ZN(n9679)
         );
  AOI22_X1 U10817 ( .A1(n9840), .A2(n9679), .B1(n6371), .B2(n9838), .ZN(
        P1_U3538) );
  OAI22_X1 U10818 ( .A1(n9668), .A2(n9827), .B1(n4777), .B2(n9826), .ZN(n9669)
         );
  AOI21_X1 U10819 ( .B1(n9670), .B2(n9832), .A(n9669), .ZN(n9671) );
  AND2_X1 U10820 ( .A1(n9672), .A2(n9671), .ZN(n9681) );
  AOI22_X1 U10821 ( .A1(n9840), .A2(n9681), .B1(n7708), .B2(n9838), .ZN(
        P1_U3536) );
  OAI22_X1 U10822 ( .A1(n9674), .A2(n9827), .B1(n9673), .B2(n9826), .ZN(n9676)
         );
  AOI211_X1 U10823 ( .C1(n9832), .C2(n9677), .A(n9676), .B(n9675), .ZN(n9683)
         );
  AOI22_X1 U10824 ( .A1(n9840), .A2(n9683), .B1(n6284), .B2(n9838), .ZN(
        P1_U3534) );
  INV_X1 U10825 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9678) );
  AOI22_X1 U10826 ( .A1(n9835), .A2(n9679), .B1(n9678), .B2(n9833), .ZN(
        P1_U3499) );
  INV_X1 U10827 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9680) );
  AOI22_X1 U10828 ( .A1(n9835), .A2(n9681), .B1(n9680), .B2(n9833), .ZN(
        P1_U3493) );
  INV_X1 U10829 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9682) );
  AOI22_X1 U10830 ( .A1(n9835), .A2(n9683), .B1(n9682), .B2(n9833), .ZN(
        P1_U3487) );
  XNOR2_X1 U10831 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10832 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10833 ( .A(n9684), .ZN(n9691) );
  OAI21_X1 U10834 ( .B1(n6084), .B2(n10433), .A(n9685), .ZN(n9686) );
  OAI211_X1 U10835 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9688), .A(n9687), .B(
        n9686), .ZN(n9689) );
  AND3_X1 U10836 ( .A1(n9691), .A2(n9690), .A3(n9689), .ZN(n9693) );
  NOR3_X1 U10837 ( .A1(n9802), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n10433), .ZN(
        n9692) );
  AOI211_X1 U10838 ( .C1(P1_ADDR_REG_0__SCAN_IN), .C2(n9694), .A(n9693), .B(
        n9692), .ZN(n9695) );
  OAI21_X1 U10839 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n7535), .A(n9695), .ZN(
        P1_U3241) );
  INV_X1 U10840 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9697) );
  OAI22_X1 U10841 ( .A1(n9806), .A2(n9697), .B1(n9713), .B2(n9696), .ZN(n9698)
         );
  INV_X1 U10842 ( .A(n9698), .ZN(n9711) );
  INV_X1 U10843 ( .A(n9699), .ZN(n9704) );
  NOR3_X1 U10844 ( .A1(n9702), .A2(n9701), .A3(n9700), .ZN(n9703) );
  OAI21_X1 U10845 ( .B1(n9704), .B2(n9703), .A(n9720), .ZN(n9709) );
  OAI211_X1 U10846 ( .C1(n9707), .C2(n9706), .A(n9783), .B(n9705), .ZN(n9708)
         );
  NAND4_X1 U10847 ( .A1(n9711), .A2(n9710), .A3(n9709), .A4(n9708), .ZN(
        P1_U3246) );
  INV_X1 U10848 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9714) );
  OAI22_X1 U10849 ( .A1(n9806), .A2(n9714), .B1(n9713), .B2(n9712), .ZN(n9715)
         );
  INV_X1 U10850 ( .A(n9715), .ZN(n9728) );
  INV_X1 U10851 ( .A(n9716), .ZN(n9727) );
  OAI21_X1 U10852 ( .B1(n9719), .B2(n9718), .A(n9717), .ZN(n9721) );
  NAND2_X1 U10853 ( .A1(n9721), .A2(n9720), .ZN(n9726) );
  OAI211_X1 U10854 ( .C1(n9724), .C2(n9723), .A(n9783), .B(n9722), .ZN(n9725)
         );
  NAND4_X1 U10855 ( .A1(n9728), .A2(n9727), .A3(n9726), .A4(n9725), .ZN(
        P1_U3249) );
  INV_X1 U10856 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9741) );
  AOI211_X1 U10857 ( .C1(n9731), .C2(n9730), .A(n9729), .B(n9790), .ZN(n9732)
         );
  AOI211_X1 U10858 ( .C1(n9796), .C2(n9734), .A(n9733), .B(n9732), .ZN(n9740)
         );
  AOI21_X1 U10859 ( .B1(n9737), .B2(n9736), .A(n9735), .ZN(n9738) );
  OR2_X1 U10860 ( .A1(n9738), .A2(n9802), .ZN(n9739) );
  OAI211_X1 U10861 ( .C1(n9741), .C2(n9806), .A(n9740), .B(n9739), .ZN(
        P1_U3253) );
  INV_X1 U10862 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9754) );
  AOI211_X1 U10863 ( .C1(n9744), .C2(n9743), .A(n9742), .B(n9790), .ZN(n9745)
         );
  AOI211_X1 U10864 ( .C1(n9796), .C2(n9747), .A(n9746), .B(n9745), .ZN(n9753)
         );
  AOI21_X1 U10865 ( .B1(n9750), .B2(n9749), .A(n9748), .ZN(n9751) );
  OR2_X1 U10866 ( .A1(n9802), .A2(n9751), .ZN(n9752) );
  OAI211_X1 U10867 ( .C1(n9754), .C2(n9806), .A(n9753), .B(n9752), .ZN(
        P1_U3254) );
  INV_X1 U10868 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9764) );
  AOI211_X1 U10869 ( .C1(n9756), .C2(n9630), .A(n9755), .B(n9790), .ZN(n9757)
         );
  AOI211_X1 U10870 ( .C1(n9796), .C2(n9759), .A(n9758), .B(n9757), .ZN(n9763)
         );
  OAI211_X1 U10871 ( .C1(n9761), .C2(P1_REG1_REG_15__SCAN_IN), .A(n9783), .B(
        n9760), .ZN(n9762) );
  OAI211_X1 U10872 ( .C1(n9806), .C2(n9764), .A(n9763), .B(n9762), .ZN(
        P1_U3256) );
  INV_X1 U10873 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10043) );
  AOI211_X1 U10874 ( .C1(n9767), .C2(n9766), .A(n9765), .B(n9790), .ZN(n9768)
         );
  AOI211_X1 U10875 ( .C1(n9796), .C2(n9770), .A(n9769), .B(n9768), .ZN(n9775)
         );
  OAI211_X1 U10876 ( .C1(n9773), .C2(n9772), .A(n9783), .B(n9771), .ZN(n9774)
         );
  OAI211_X1 U10877 ( .C1(n9806), .C2(n10043), .A(n9775), .B(n9774), .ZN(
        P1_U3257) );
  INV_X1 U10878 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9788) );
  AOI211_X1 U10879 ( .C1(n9778), .C2(n9777), .A(n9776), .B(n9790), .ZN(n9779)
         );
  AOI211_X1 U10880 ( .C1(n9796), .C2(n9781), .A(n9780), .B(n9779), .ZN(n9787)
         );
  OAI211_X1 U10881 ( .C1(n9785), .C2(n9784), .A(n9783), .B(n9782), .ZN(n9786)
         );
  OAI211_X1 U10882 ( .C1(n9806), .C2(n9788), .A(n9787), .B(n9786), .ZN(
        P1_U3258) );
  INV_X1 U10883 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9805) );
  INV_X1 U10884 ( .A(n9789), .ZN(n9795) );
  AOI211_X1 U10885 ( .C1(n9793), .C2(n9792), .A(n9791), .B(n9790), .ZN(n9794)
         );
  AOI211_X1 U10886 ( .C1(n9797), .C2(n9796), .A(n9795), .B(n9794), .ZN(n9804)
         );
  AOI21_X1 U10887 ( .B1(n9800), .B2(n9799), .A(n9798), .ZN(n9801) );
  OR2_X1 U10888 ( .A1(n9802), .A2(n9801), .ZN(n9803) );
  OAI211_X1 U10889 ( .C1(n9806), .C2(n9805), .A(n9804), .B(n9803), .ZN(
        P1_U3259) );
  AND2_X1 U10890 ( .A1(n9808), .A2(n9807), .ZN(n9810) );
  AND2_X1 U10891 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9809), .ZN(P1_U3292) );
  AND2_X1 U10892 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9809), .ZN(P1_U3293) );
  AND2_X1 U10893 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9809), .ZN(P1_U3294) );
  AND2_X1 U10894 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9809), .ZN(P1_U3295) );
  AND2_X1 U10895 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9809), .ZN(P1_U3296) );
  AND2_X1 U10896 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9809), .ZN(P1_U3297) );
  AND2_X1 U10897 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9809), .ZN(P1_U3298) );
  AND2_X1 U10898 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9809), .ZN(P1_U3299) );
  AND2_X1 U10899 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9809), .ZN(P1_U3300) );
  AND2_X1 U10900 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9809), .ZN(P1_U3301) );
  AND2_X1 U10901 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9809), .ZN(P1_U3302) );
  AND2_X1 U10902 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9809), .ZN(P1_U3303) );
  AND2_X1 U10903 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9809), .ZN(P1_U3304) );
  AND2_X1 U10904 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9809), .ZN(P1_U3305) );
  AND2_X1 U10905 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9809), .ZN(P1_U3306) );
  AND2_X1 U10906 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9809), .ZN(P1_U3307) );
  AND2_X1 U10907 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9809), .ZN(P1_U3308) );
  AND2_X1 U10908 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9809), .ZN(P1_U3309) );
  AND2_X1 U10909 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9809), .ZN(P1_U3310) );
  AND2_X1 U10910 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9809), .ZN(P1_U3311) );
  AND2_X1 U10911 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9809), .ZN(P1_U3312) );
  AND2_X1 U10912 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9809), .ZN(P1_U3313) );
  AND2_X1 U10913 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9809), .ZN(P1_U3314) );
  AND2_X1 U10914 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9809), .ZN(P1_U3315) );
  AND2_X1 U10915 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9809), .ZN(P1_U3316) );
  AND2_X1 U10916 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9809), .ZN(P1_U3317) );
  AND2_X1 U10917 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9809), .ZN(P1_U3318) );
  AND2_X1 U10918 ( .A1(n9809), .A2(P1_D_REG_4__SCAN_IN), .ZN(P1_U3319) );
  INV_X1 U10919 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10087) );
  NOR2_X1 U10920 ( .A1(n9810), .A2(n10087), .ZN(P1_U3320) );
  INV_X1 U10921 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10110) );
  NOR2_X1 U10922 ( .A1(n9810), .A2(n10110), .ZN(P1_U3321) );
  OAI22_X1 U10923 ( .A1(n9812), .A2(n9827), .B1(n9811), .B2(n9826), .ZN(n9814)
         );
  AOI211_X1 U10924 ( .C1(n9832), .C2(n9815), .A(n9814), .B(n9813), .ZN(n9836)
         );
  INV_X1 U10925 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9816) );
  AOI22_X1 U10926 ( .A1(n9835), .A2(n9836), .B1(n9816), .B2(n9833), .ZN(
        P1_U3463) );
  OAI21_X1 U10927 ( .B1(n9818), .B2(n9826), .A(n9817), .ZN(n9820) );
  AOI211_X1 U10928 ( .C1(n9822), .C2(n9821), .A(n9820), .B(n9819), .ZN(n9837)
         );
  INV_X1 U10929 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9823) );
  AOI22_X1 U10930 ( .A1(n9835), .A2(n9837), .B1(n9823), .B2(n9833), .ZN(
        P1_U3469) );
  INV_X1 U10931 ( .A(n9824), .ZN(n9831) );
  OAI22_X1 U10932 ( .A1(n9828), .A2(n9827), .B1(n6769), .B2(n9826), .ZN(n9830)
         );
  AOI211_X1 U10933 ( .C1(n9832), .C2(n9831), .A(n9830), .B(n9829), .ZN(n9839)
         );
  INV_X1 U10934 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9834) );
  AOI22_X1 U10935 ( .A1(n9835), .A2(n9839), .B1(n9834), .B2(n9833), .ZN(
        P1_U3481) );
  AOI22_X1 U10936 ( .A1(n9840), .A2(n9836), .B1(n7003), .B2(n9838), .ZN(
        P1_U3526) );
  AOI22_X1 U10937 ( .A1(n9840), .A2(n9837), .B1(n7007), .B2(n9838), .ZN(
        P1_U3528) );
  AOI22_X1 U10938 ( .A1(n9840), .A2(n9839), .B1(n6251), .B2(n9838), .ZN(
        P1_U3532) );
  AOI22_X1 U10939 ( .A1(n9901), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9906), .ZN(n9848) );
  AOI22_X1 U10940 ( .A1(n9899), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9847) );
  NOR2_X1 U10941 ( .A1(n9841), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9845) );
  OAI21_X1 U10942 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(n9843), .A(n9842), .ZN(
        n9844) );
  OAI21_X1 U10943 ( .B1(n9845), .B2(n9844), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n9846) );
  OAI211_X1 U10944 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n9848), .A(n9847), .B(
        n9846), .ZN(P2_U3245) );
  AOI22_X1 U10945 ( .A1(n9899), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(P2_U3152), .ZN(n9859) );
  NAND2_X1 U10946 ( .A1(n9905), .A2(n9849), .ZN(n9858) );
  OAI211_X1 U10947 ( .C1(n9852), .C2(n9851), .A(n9906), .B(n9850), .ZN(n9857)
         );
  OAI211_X1 U10948 ( .C1(n9855), .C2(n9854), .A(n9901), .B(n9853), .ZN(n9856)
         );
  NAND4_X1 U10949 ( .A1(n9859), .A2(n9858), .A3(n9857), .A4(n9856), .ZN(
        P2_U3248) );
  AOI21_X1 U10950 ( .B1(n9899), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n9860), .ZN(
        n9871) );
  NAND2_X1 U10951 ( .A1(n9905), .A2(n9861), .ZN(n9870) );
  OAI211_X1 U10952 ( .C1(n9864), .C2(n9863), .A(n9901), .B(n9862), .ZN(n9869)
         );
  OAI211_X1 U10953 ( .C1(n9867), .C2(n9866), .A(n9906), .B(n9865), .ZN(n9868)
         );
  NAND4_X1 U10954 ( .A1(n9871), .A2(n9870), .A3(n9869), .A4(n9868), .ZN(
        P2_U3249) );
  INV_X1 U10955 ( .A(n9872), .ZN(n9873) );
  AOI21_X1 U10956 ( .B1(n9899), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n9873), .ZN(
        n9884) );
  NAND2_X1 U10957 ( .A1(n9905), .A2(n9874), .ZN(n9883) );
  OAI211_X1 U10958 ( .C1(n9877), .C2(n9876), .A(n9901), .B(n9875), .ZN(n9882)
         );
  OAI211_X1 U10959 ( .C1(n9880), .C2(n9879), .A(n9906), .B(n9878), .ZN(n9881)
         );
  NAND4_X1 U10960 ( .A1(n9884), .A2(n9883), .A3(n9882), .A4(n9881), .ZN(
        P2_U3251) );
  AOI21_X1 U10961 ( .B1(n9899), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n9885), .ZN(
        n9896) );
  NAND2_X1 U10962 ( .A1(n9905), .A2(n9886), .ZN(n9895) );
  OAI211_X1 U10963 ( .C1(n9889), .C2(n9888), .A(n9887), .B(n9906), .ZN(n9894)
         );
  OAI211_X1 U10964 ( .C1(n9892), .C2(n9891), .A(n9890), .B(n9901), .ZN(n9893)
         );
  NAND4_X1 U10965 ( .A1(n9896), .A2(n9895), .A3(n9894), .A4(n9893), .ZN(
        P2_U3253) );
  INV_X1 U10966 ( .A(n9897), .ZN(n9898) );
  AOI21_X1 U10967 ( .B1(n9899), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n9898), .ZN(
        n9913) );
  OAI211_X1 U10968 ( .C1(n9903), .C2(n9902), .A(n9901), .B(n9900), .ZN(n9912)
         );
  NAND2_X1 U10969 ( .A1(n9905), .A2(n9904), .ZN(n9911) );
  OAI211_X1 U10970 ( .C1(n9909), .C2(n9908), .A(n9907), .B(n9906), .ZN(n9910)
         );
  NAND4_X1 U10971 ( .A1(n9913), .A2(n9912), .A3(n9911), .A4(n9910), .ZN(
        P2_U3262) );
  XNOR2_X1 U10972 ( .A(n9914), .B(n9915), .ZN(n9987) );
  NAND2_X1 U10973 ( .A1(n9916), .A2(n9915), .ZN(n9918) );
  AOI21_X1 U10974 ( .B1(n9919), .B2(n9918), .A(n9917), .ZN(n9920) );
  AOI211_X1 U10975 ( .C1(n9987), .C2(n9922), .A(n9921), .B(n9920), .ZN(n9984)
         );
  INV_X1 U10976 ( .A(n9923), .ZN(n9924) );
  AOI222_X1 U10977 ( .A1(n9927), .A2(n9926), .B1(P2_REG2_REG_8__SCAN_IN), .B2(
        n9936), .C1(n9925), .C2(n9924), .ZN(n9935) );
  INV_X1 U10978 ( .A(n9928), .ZN(n9930) );
  OAI21_X1 U10979 ( .B1(n9930), .B2(n9982), .A(n9929), .ZN(n9983) );
  INV_X1 U10980 ( .A(n9983), .ZN(n9931) );
  AOI22_X1 U10981 ( .A1(n9987), .A2(n9933), .B1(n9932), .B2(n9931), .ZN(n9934)
         );
  OAI211_X1 U10982 ( .C1(n9936), .C2(n9984), .A(n9935), .B(n9934), .ZN(
        P2_U3288) );
  INV_X1 U10983 ( .A(n9937), .ZN(n9939) );
  AND2_X1 U10984 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9942), .ZN(P2_U3297) );
  AND2_X1 U10985 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9942), .ZN(P2_U3298) );
  AND2_X1 U10986 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9942), .ZN(P2_U3299) );
  AND2_X1 U10987 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9942), .ZN(P2_U3300) );
  AND2_X1 U10988 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9942), .ZN(P2_U3301) );
  AND2_X1 U10989 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9942), .ZN(P2_U3302) );
  AND2_X1 U10990 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9942), .ZN(P2_U3303) );
  AND2_X1 U10991 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9942), .ZN(P2_U3304) );
  AND2_X1 U10992 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9942), .ZN(P2_U3305) );
  AND2_X1 U10993 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9942), .ZN(P2_U3306) );
  AND2_X1 U10994 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9942), .ZN(P2_U3307) );
  AND2_X1 U10995 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9942), .ZN(P2_U3308) );
  AND2_X1 U10996 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9942), .ZN(P2_U3309) );
  AND2_X1 U10997 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9942), .ZN(P2_U3310) );
  AND2_X1 U10998 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9942), .ZN(P2_U3311) );
  AND2_X1 U10999 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9942), .ZN(P2_U3312) );
  AND2_X1 U11000 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9942), .ZN(P2_U3313) );
  AND2_X1 U11001 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9942), .ZN(P2_U3314) );
  AND2_X1 U11002 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9942), .ZN(P2_U3315) );
  AND2_X1 U11003 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9942), .ZN(P2_U3316) );
  AND2_X1 U11004 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9942), .ZN(P2_U3317) );
  AND2_X1 U11005 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9942), .ZN(P2_U3318) );
  AND2_X1 U11006 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9942), .ZN(P2_U3319) );
  AND2_X1 U11007 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9942), .ZN(P2_U3320) );
  AND2_X1 U11008 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9942), .ZN(P2_U3321) );
  AND2_X1 U11009 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9942), .ZN(P2_U3322) );
  AND2_X1 U11010 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9942), .ZN(P2_U3323) );
  AND2_X1 U11011 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9942), .ZN(P2_U3324) );
  AND2_X1 U11012 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9942), .ZN(P2_U3325) );
  AND2_X1 U11013 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9942), .ZN(P2_U3326) );
  AOI22_X1 U11014 ( .A1(n9941), .A2(n9942), .B1(n9945), .B2(n9940), .ZN(
        P2_U3437) );
  AOI22_X1 U11015 ( .A1(n9945), .A2(n9944), .B1(n9943), .B2(n9942), .ZN(
        P2_U3438) );
  AOI22_X1 U11016 ( .A1(n9948), .A2(n10018), .B1(n9947), .B2(n9946), .ZN(n9949) );
  AND2_X1 U11017 ( .A1(n9950), .A2(n9949), .ZN(n10023) );
  INV_X1 U11018 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9951) );
  AOI22_X1 U11019 ( .A1(n10021), .A2(n10023), .B1(n9951), .B2(n10019), .ZN(
        P2_U3451) );
  OAI22_X1 U11020 ( .A1(n9953), .A2(n10013), .B1(n9952), .B2(n10011), .ZN(
        n9955) );
  AOI211_X1 U11021 ( .C1(n10018), .C2(n9956), .A(n9955), .B(n9954), .ZN(n10024) );
  INV_X1 U11022 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9957) );
  AOI22_X1 U11023 ( .A1(n10021), .A2(n10024), .B1(n9957), .B2(n10019), .ZN(
        P2_U3457) );
  OAI22_X1 U11024 ( .A1(n9959), .A2(n10013), .B1(n9958), .B2(n10011), .ZN(
        n9961) );
  AOI211_X1 U11025 ( .C1(n10018), .C2(n9962), .A(n9961), .B(n9960), .ZN(n10025) );
  INV_X1 U11026 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9963) );
  AOI22_X1 U11027 ( .A1(n10021), .A2(n10025), .B1(n9963), .B2(n10019), .ZN(
        P2_U3463) );
  OAI211_X1 U11028 ( .C1(n9966), .C2(n10011), .A(n9965), .B(n9964), .ZN(n9967)
         );
  AOI21_X1 U11029 ( .B1(n10018), .B2(n9968), .A(n9967), .ZN(n10026) );
  INV_X1 U11030 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9969) );
  AOI22_X1 U11031 ( .A1(n10021), .A2(n10026), .B1(n9969), .B2(n10019), .ZN(
        P2_U3466) );
  OAI22_X1 U11032 ( .A1(n9971), .A2(n10013), .B1(n9970), .B2(n10011), .ZN(
        n9972) );
  AOI211_X1 U11033 ( .C1(n9974), .C2(n10018), .A(n9973), .B(n9972), .ZN(n10027) );
  INV_X1 U11034 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9975) );
  AOI22_X1 U11035 ( .A1(n10021), .A2(n10027), .B1(n9975), .B2(n10019), .ZN(
        P2_U3469) );
  OAI22_X1 U11036 ( .A1(n9977), .A2(n10013), .B1(n9976), .B2(n10011), .ZN(
        n9979) );
  AOI211_X1 U11037 ( .C1(n9980), .C2(n10018), .A(n9979), .B(n9978), .ZN(n10028) );
  INV_X1 U11038 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9981) );
  AOI22_X1 U11039 ( .A1(n10021), .A2(n10028), .B1(n9981), .B2(n10019), .ZN(
        P2_U3472) );
  OAI22_X1 U11040 ( .A1(n9983), .A2(n10013), .B1(n9982), .B2(n10011), .ZN(
        n9986) );
  INV_X1 U11041 ( .A(n9984), .ZN(n9985) );
  AOI211_X1 U11042 ( .C1(n10002), .C2(n9987), .A(n9986), .B(n9985), .ZN(n10029) );
  INV_X1 U11043 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9988) );
  AOI22_X1 U11044 ( .A1(n10021), .A2(n10029), .B1(n9988), .B2(n10019), .ZN(
        P2_U3475) );
  INV_X1 U11045 ( .A(n9989), .ZN(n9994) );
  OAI22_X1 U11046 ( .A1(n9991), .A2(n10013), .B1(n9990), .B2(n10011), .ZN(
        n9993) );
  AOI211_X1 U11047 ( .C1(n10002), .C2(n9994), .A(n9993), .B(n9992), .ZN(n10030) );
  INV_X1 U11048 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9995) );
  AOI22_X1 U11049 ( .A1(n10021), .A2(n10030), .B1(n9995), .B2(n10019), .ZN(
        P2_U3478) );
  INV_X1 U11050 ( .A(n9996), .ZN(n10001) );
  OAI22_X1 U11051 ( .A1(n9998), .A2(n10013), .B1(n9997), .B2(n10011), .ZN(
        n10000) );
  AOI211_X1 U11052 ( .C1(n10002), .C2(n10001), .A(n10000), .B(n9999), .ZN(
        n10031) );
  INV_X1 U11053 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10003) );
  AOI22_X1 U11054 ( .A1(n10021), .A2(n10031), .B1(n10003), .B2(n10019), .ZN(
        P2_U3481) );
  INV_X1 U11055 ( .A(n10004), .ZN(n10009) );
  OAI22_X1 U11056 ( .A1(n10006), .A2(n10013), .B1(n10005), .B2(n10011), .ZN(
        n10008) );
  AOI211_X1 U11057 ( .C1(n10009), .C2(n10018), .A(n10008), .B(n10007), .ZN(
        n10032) );
  INV_X1 U11058 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10010) );
  AOI22_X1 U11059 ( .A1(n10021), .A2(n10032), .B1(n10010), .B2(n10019), .ZN(
        P2_U3484) );
  OAI22_X1 U11060 ( .A1(n10014), .A2(n10013), .B1(n10012), .B2(n10011), .ZN(
        n10016) );
  AOI211_X1 U11061 ( .C1(n10018), .C2(n10017), .A(n10016), .B(n10015), .ZN(
        n10035) );
  INV_X1 U11062 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10020) );
  AOI22_X1 U11063 ( .A1(n10021), .A2(n10035), .B1(n10020), .B2(n10019), .ZN(
        P2_U3487) );
  INV_X1 U11064 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10022) );
  AOI22_X1 U11065 ( .A1(n10036), .A2(n10023), .B1(n10022), .B2(n10033), .ZN(
        P2_U3520) );
  AOI22_X1 U11066 ( .A1(n10036), .A2(n10024), .B1(n6929), .B2(n10033), .ZN(
        P2_U3522) );
  AOI22_X1 U11067 ( .A1(n10036), .A2(n10025), .B1(n6934), .B2(n10033), .ZN(
        P2_U3524) );
  AOI22_X1 U11068 ( .A1(n10036), .A2(n10026), .B1(n6936), .B2(n10033), .ZN(
        P2_U3525) );
  AOI22_X1 U11069 ( .A1(n10036), .A2(n10027), .B1(n6927), .B2(n10033), .ZN(
        P2_U3526) );
  AOI22_X1 U11070 ( .A1(n10036), .A2(n10028), .B1(n6940), .B2(n10033), .ZN(
        P2_U3527) );
  AOI22_X1 U11071 ( .A1(n10036), .A2(n10029), .B1(n6926), .B2(n10033), .ZN(
        P2_U3528) );
  AOI22_X1 U11072 ( .A1(n10036), .A2(n10030), .B1(n6925), .B2(n10033), .ZN(
        P2_U3529) );
  AOI22_X1 U11073 ( .A1(n10036), .A2(n10031), .B1(n6924), .B2(n10033), .ZN(
        P2_U3530) );
  AOI22_X1 U11074 ( .A1(n10036), .A2(n10032), .B1(n6944), .B2(n10033), .ZN(
        P2_U3531) );
  AOI22_X1 U11075 ( .A1(n10036), .A2(n10035), .B1(n10034), .B2(n10033), .ZN(
        P2_U3532) );
  NAND3_X1 U11076 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10040) );
  NAND2_X1 U11077 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n10037) );
  NAND2_X1 U11078 ( .A1(n10038), .A2(n10037), .ZN(n10057) );
  INV_X1 U11079 ( .A(n10057), .ZN(n10039) );
  NAND2_X1 U11080 ( .A1(n10041), .A2(n10040), .ZN(n10056) );
  OAI222_X1 U11081 ( .A1(n10041), .A2(n10040), .B1(n10041), .B2(n10057), .C1(
        n10039), .C2(n10056), .ZN(ADD_1071_U5) );
  XOR2_X1 U11082 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  NOR2_X1 U11083 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(P2_ADDR_REG_17__SCAN_IN), 
        .ZN(n10042) );
  AOI21_X1 U11084 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10042), .ZN(n10062) );
  AOI22_X1 U11085 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(P2_ADDR_REG_16__SCAN_IN), 
        .B1(n10044), .B2(n10043), .ZN(n10065) );
  NOR2_X1 U11086 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(P2_ADDR_REG_15__SCAN_IN), 
        .ZN(n10045) );
  AOI21_X1 U11087 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10045), .ZN(n10068) );
  NOR2_X1 U11088 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10046) );
  AOI21_X1 U11089 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10046), .ZN(n10071) );
  NOR2_X1 U11090 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10047) );
  AOI21_X1 U11091 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10047), .ZN(n10074) );
  NOR2_X1 U11092 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10048) );
  AOI21_X1 U11093 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10048), .ZN(n10077) );
  NOR2_X1 U11094 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10049) );
  AOI21_X1 U11095 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10049), .ZN(n10080) );
  NOR2_X1 U11096 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10050) );
  AOI21_X1 U11097 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10050), .ZN(n10083) );
  NOR2_X1 U11098 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(P2_ADDR_REG_9__SCAN_IN), 
        .ZN(n10051) );
  AOI21_X1 U11099 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10051), .ZN(n10458) );
  NOR2_X1 U11100 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(P2_ADDR_REG_8__SCAN_IN), 
        .ZN(n10052) );
  AOI21_X1 U11101 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10052), .ZN(n10473) );
  NOR2_X1 U11102 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10053) );
  AOI21_X1 U11103 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n10053), .ZN(n10461) );
  NOR2_X1 U11104 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n10054) );
  AOI21_X1 U11105 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10054), .ZN(n10476) );
  NOR2_X1 U11106 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(P2_ADDR_REG_5__SCAN_IN), 
        .ZN(n10055) );
  AOI21_X1 U11107 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10055), .ZN(n10467) );
  NAND2_X1 U11108 ( .A1(n10057), .A2(n10056), .ZN(n10464) );
  NAND2_X1 U11109 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n10058) );
  OAI21_X1 U11110 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10058), .ZN(n10463) );
  NOR2_X1 U11111 ( .A1(n10464), .A2(n10463), .ZN(n10462) );
  AOI21_X1 U11112 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n10462), .ZN(n10479) );
  NAND2_X1 U11113 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10059) );
  OAI21_X1 U11114 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10059), .ZN(n10478) );
  NOR2_X1 U11115 ( .A1(n10479), .A2(n10478), .ZN(n10477) );
  AOI21_X1 U11116 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10477), .ZN(n10482) );
  NOR2_X1 U11117 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10060) );
  AOI21_X1 U11118 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n10060), .ZN(n10481) );
  NAND2_X1 U11119 ( .A1(n10482), .A2(n10481), .ZN(n10480) );
  OAI21_X1 U11120 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10480), .ZN(n10466) );
  NAND2_X1 U11121 ( .A1(n10467), .A2(n10466), .ZN(n10465) );
  OAI21_X1 U11122 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n10465), .ZN(n10475) );
  NAND2_X1 U11123 ( .A1(n10476), .A2(n10475), .ZN(n10474) );
  OAI21_X1 U11124 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n10474), .ZN(n10460) );
  NAND2_X1 U11125 ( .A1(n10461), .A2(n10460), .ZN(n10459) );
  OAI21_X1 U11126 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10459), .ZN(n10472) );
  NAND2_X1 U11127 ( .A1(n10473), .A2(n10472), .ZN(n10471) );
  OAI21_X1 U11128 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n10471), .ZN(n10457) );
  NAND2_X1 U11129 ( .A1(n10458), .A2(n10457), .ZN(n10456) );
  OAI21_X1 U11130 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n10456), .ZN(n10082) );
  NAND2_X1 U11131 ( .A1(n10083), .A2(n10082), .ZN(n10081) );
  OAI21_X1 U11132 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10081), .ZN(n10079) );
  NAND2_X1 U11133 ( .A1(n10080), .A2(n10079), .ZN(n10078) );
  OAI21_X1 U11134 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10078), .ZN(n10076) );
  NAND2_X1 U11135 ( .A1(n10077), .A2(n10076), .ZN(n10075) );
  OAI21_X1 U11136 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10075), .ZN(n10073) );
  NAND2_X1 U11137 ( .A1(n10074), .A2(n10073), .ZN(n10072) );
  OAI21_X1 U11138 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10072), .ZN(n10070) );
  NAND2_X1 U11139 ( .A1(n10071), .A2(n10070), .ZN(n10069) );
  OAI21_X1 U11140 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10069), .ZN(n10067) );
  NAND2_X1 U11141 ( .A1(n10068), .A2(n10067), .ZN(n10066) );
  OAI21_X1 U11142 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10066), .ZN(n10064) );
  NAND2_X1 U11143 ( .A1(n10065), .A2(n10064), .ZN(n10063) );
  OAI21_X1 U11144 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10063), .ZN(n10061) );
  NAND2_X1 U11145 ( .A1(n10062), .A2(n10061), .ZN(n10451) );
  OAI21_X1 U11146 ( .B1(n10062), .B2(n10061), .A(n10451), .ZN(ADD_1071_U56) );
  OAI21_X1 U11147 ( .B1(n10065), .B2(n10064), .A(n10063), .ZN(ADD_1071_U57) );
  OAI21_X1 U11148 ( .B1(n10068), .B2(n10067), .A(n10066), .ZN(ADD_1071_U58) );
  OAI21_X1 U11149 ( .B1(n10071), .B2(n10070), .A(n10069), .ZN(ADD_1071_U59) );
  OAI21_X1 U11150 ( .B1(n10074), .B2(n10073), .A(n10072), .ZN(ADD_1071_U60) );
  OAI21_X1 U11151 ( .B1(n10077), .B2(n10076), .A(n10075), .ZN(ADD_1071_U61) );
  OAI21_X1 U11152 ( .B1(n10080), .B2(n10079), .A(n10078), .ZN(ADD_1071_U62) );
  OAI21_X1 U11153 ( .B1(n10083), .B2(n10082), .A(n10081), .ZN(ADD_1071_U63) );
  INV_X1 U11154 ( .A(SI_4_), .ZN(n10255) );
  AOI22_X1 U11155 ( .A1(n10085), .A2(keyinput_f57), .B1(n6030), .B2(
        keyinput_f107), .ZN(n10084) );
  OAI221_X1 U11156 ( .B1(n10085), .B2(keyinput_f57), .C1(n6030), .C2(
        keyinput_f107), .A(n10084), .ZN(n10096) );
  AOI22_X1 U11157 ( .A1(n5572), .A2(keyinput_f50), .B1(n10087), .B2(
        keyinput_f126), .ZN(n10086) );
  OAI221_X1 U11158 ( .B1(n5572), .B2(keyinput_f50), .C1(n10087), .C2(
        keyinput_f126), .A(n10086), .ZN(n10095) );
  AOI22_X1 U11159 ( .A1(n10090), .A2(keyinput_f79), .B1(keyinput_f66), .B2(
        n10089), .ZN(n10088) );
  OAI221_X1 U11160 ( .B1(n10090), .B2(keyinput_f79), .C1(n10089), .C2(
        keyinput_f66), .A(n10088), .ZN(n10094) );
  XOR2_X1 U11161 ( .A(n5423), .B(keyinput_f53), .Z(n10092) );
  XNOR2_X1 U11162 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_f94), .ZN(n10091) );
  NAND2_X1 U11163 ( .A1(n10092), .A2(n10091), .ZN(n10093) );
  NOR4_X1 U11164 ( .A1(n10096), .A2(n10095), .A3(n10094), .A4(n10093), .ZN(
        n10250) );
  INV_X1 U11165 ( .A(SI_30_), .ZN(n10098) );
  AOI22_X1 U11166 ( .A1(n10098), .A2(keyinput_f2), .B1(n5146), .B2(
        keyinput_f21), .ZN(n10097) );
  OAI221_X1 U11167 ( .B1(n10098), .B2(keyinput_f2), .C1(n5146), .C2(
        keyinput_f21), .A(n10097), .ZN(n10108) );
  INV_X1 U11168 ( .A(SI_18_), .ZN(n10432) );
  AOI22_X1 U11169 ( .A1(n10394), .A2(keyinput_f54), .B1(n10432), .B2(
        keyinput_f14), .ZN(n10099) );
  OAI221_X1 U11170 ( .B1(n10394), .B2(keyinput_f54), .C1(n10432), .C2(
        keyinput_f14), .A(n10099), .ZN(n10107) );
  AOI22_X1 U11171 ( .A1(n10102), .A2(keyinput_f39), .B1(n10101), .B2(
        keyinput_f90), .ZN(n10100) );
  OAI221_X1 U11172 ( .B1(n10102), .B2(keyinput_f39), .C1(n10101), .C2(
        keyinput_f90), .A(n10100), .ZN(n10106) );
  XNOR2_X1 U11173 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_f117), .ZN(n10104)
         );
  XNOR2_X1 U11174 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_f36), .ZN(n10103)
         );
  NAND2_X1 U11175 ( .A1(n10104), .A2(n10103), .ZN(n10105) );
  NOR4_X1 U11176 ( .A1(n10108), .A2(n10107), .A3(n10106), .A4(n10105), .ZN(
        n10249) );
  XOR2_X1 U11177 ( .A(keyinput_f0), .B(P2_WR_REG_SCAN_IN), .Z(n10118) );
  AOI22_X1 U11178 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(keyinput_f35), .B1(SI_27_), .B2(keyinput_f5), .ZN(n10109) );
  OAI221_X1 U11179 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_f35), .C1(
        SI_27_), .C2(keyinput_f5), .A(n10109), .ZN(n10117) );
  XNOR2_X1 U11180 ( .A(n10110), .B(keyinput_f125), .ZN(n10116) );
  XNOR2_X1 U11181 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_f119), .ZN(n10114)
         );
  XNOR2_X1 U11182 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_f100), .ZN(n10113)
         );
  XNOR2_X1 U11183 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_f74), .ZN(n10112) );
  XNOR2_X1 U11184 ( .A(keyinput_f92), .B(P1_IR_REG_1__SCAN_IN), .ZN(n10111) );
  NAND4_X1 U11185 ( .A1(n10114), .A2(n10113), .A3(n10112), .A4(n10111), .ZN(
        n10115) );
  OR4_X1 U11186 ( .A1(n10118), .A2(n10117), .A3(n10116), .A4(n10115), .ZN(
        n10128) );
  OAI22_X1 U11187 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(keyinput_f101), .B1(
        keyinput_f42), .B2(P2_REG3_REG_28__SCAN_IN), .ZN(n10119) );
  AOI221_X1 U11188 ( .B1(P1_IR_REG_10__SCAN_IN), .B2(keyinput_f101), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_f42), .A(n10119), .ZN(n10126)
         );
  OAI22_X1 U11189 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput_f48), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .ZN(n10120) );
  AOI221_X1 U11190 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_f48), .C1(
        keyinput_f58), .C2(P2_REG3_REG_11__SCAN_IN), .A(n10120), .ZN(n10125)
         );
  OAI22_X1 U11191 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(keyinput_f98), .B1(
        keyinput_f12), .B2(SI_20_), .ZN(n10121) );
  AOI221_X1 U11192 ( .B1(P1_IR_REG_7__SCAN_IN), .B2(keyinput_f98), .C1(SI_20_), 
        .C2(keyinput_f12), .A(n10121), .ZN(n10124) );
  OAI22_X1 U11193 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(keyinput_f73), .B1(
        P1_IR_REG_29__SCAN_IN), .B2(keyinput_f120), .ZN(n10122) );
  AOI221_X1 U11194 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(keyinput_f73), .C1(
        keyinput_f120), .C2(P1_IR_REG_29__SCAN_IN), .A(n10122), .ZN(n10123) );
  NAND4_X1 U11195 ( .A1(n10126), .A2(n10125), .A3(n10124), .A4(n10123), .ZN(
        n10127) );
  NOR2_X1 U11196 ( .A1(n10128), .A2(n10127), .ZN(n10248) );
  OAI22_X1 U11197 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(keyinput_f105), .B1(
        keyinput_f123), .B2(P1_D_REG_0__SCAN_IN), .ZN(n10129) );
  AOI221_X1 U11198 ( .B1(P1_IR_REG_14__SCAN_IN), .B2(keyinput_f105), .C1(
        P1_D_REG_0__SCAN_IN), .C2(keyinput_f123), .A(n10129), .ZN(n10136) );
  OAI22_X1 U11199 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(keyinput_f115), .B1(
        P2_B_REG_SCAN_IN), .B2(keyinput_f64), .ZN(n10130) );
  AOI221_X1 U11200 ( .B1(P1_IR_REG_24__SCAN_IN), .B2(keyinput_f115), .C1(
        keyinput_f64), .C2(P2_B_REG_SCAN_IN), .A(n10130), .ZN(n10135) );
  OAI22_X1 U11201 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput_f87), .B1(
        keyinput_f43), .B2(P2_REG3_REG_8__SCAN_IN), .ZN(n10131) );
  AOI221_X1 U11202 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_f87), .C1(
        P2_REG3_REG_8__SCAN_IN), .C2(keyinput_f43), .A(n10131), .ZN(n10134) );
  OAI22_X1 U11203 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput_f88), .B1(
        keyinput_f46), .B2(P2_REG3_REG_12__SCAN_IN), .ZN(n10132) );
  AOI221_X1 U11204 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_f88), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput_f46), .A(n10132), .ZN(n10133)
         );
  NAND4_X1 U11205 ( .A1(n10136), .A2(n10135), .A3(n10134), .A4(n10133), .ZN(
        n10246) );
  OAI22_X1 U11206 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput_f111), .B1(
        keyinput_f59), .B2(P2_REG3_REG_2__SCAN_IN), .ZN(n10137) );
  AOI221_X1 U11207 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput_f111), .C1(
        P2_REG3_REG_2__SCAN_IN), .C2(keyinput_f59), .A(n10137), .ZN(n10162) );
  OAI22_X1 U11208 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(keyinput_f77), .B1(
        keyinput_f38), .B2(P2_REG3_REG_23__SCAN_IN), .ZN(n10138) );
  AOI221_X1 U11209 ( .B1(P2_DATAO_REG_19__SCAN_IN), .B2(keyinput_f77), .C1(
        P2_REG3_REG_23__SCAN_IN), .C2(keyinput_f38), .A(n10138), .ZN(n10141)
         );
  OAI22_X1 U11210 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(keyinput_f109), .B1(SI_16_), .B2(keyinput_f16), .ZN(n10139) );
  AOI221_X1 U11211 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(keyinput_f109), .C1(
        keyinput_f16), .C2(SI_16_), .A(n10139), .ZN(n10140) );
  OAI211_X1 U11212 ( .C1(n6063), .C2(keyinput_f118), .A(n10141), .B(n10140), 
        .ZN(n10142) );
  AOI21_X1 U11213 ( .B1(n6063), .B2(keyinput_f118), .A(n10142), .ZN(n10161) );
  AOI22_X1 U11214 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(keyinput_f121), .B1(
        P1_IR_REG_5__SCAN_IN), .B2(keyinput_f96), .ZN(n10143) );
  OAI221_X1 U11215 ( .B1(P1_IR_REG_30__SCAN_IN), .B2(keyinput_f121), .C1(
        P1_IR_REG_5__SCAN_IN), .C2(keyinput_f96), .A(n10143), .ZN(n10150) );
  AOI22_X1 U11216 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput_f41), .B1(
        P1_IR_REG_11__SCAN_IN), .B2(keyinput_f102), .ZN(n10144) );
  OAI221_X1 U11217 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .C1(
        P1_IR_REG_11__SCAN_IN), .C2(keyinput_f102), .A(n10144), .ZN(n10149) );
  AOI22_X1 U11218 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(keyinput_f78), .B1(
        P2_RD_REG_SCAN_IN), .B2(keyinput_f33), .ZN(n10145) );
  OAI221_X1 U11219 ( .B1(P2_DATAO_REG_18__SCAN_IN), .B2(keyinput_f78), .C1(
        P2_RD_REG_SCAN_IN), .C2(keyinput_f33), .A(n10145), .ZN(n10148) );
  AOI22_X1 U11220 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_f47), .B1(SI_6_), .B2(keyinput_f26), .ZN(n10146) );
  OAI221_X1 U11221 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .C1(
        SI_6_), .C2(keyinput_f26), .A(n10146), .ZN(n10147) );
  NOR4_X1 U11222 ( .A1(n10150), .A2(n10149), .A3(n10148), .A4(n10147), .ZN(
        n10160) );
  AOI22_X1 U11223 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(keyinput_f68), .B1(
        SI_0_), .B2(keyinput_f32), .ZN(n10151) );
  OAI221_X1 U11224 ( .B1(P2_DATAO_REG_28__SCAN_IN), .B2(keyinput_f68), .C1(
        SI_0_), .C2(keyinput_f32), .A(n10151), .ZN(n10158) );
  AOI22_X1 U11225 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(keyinput_f85), .B1(
        SI_19_), .B2(keyinput_f13), .ZN(n10152) );
  OAI221_X1 U11226 ( .B1(P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_f85), .C1(
        SI_19_), .C2(keyinput_f13), .A(n10152), .ZN(n10157) );
  AOI22_X1 U11227 ( .A1(SI_1_), .A2(keyinput_f31), .B1(P1_D_REG_4__SCAN_IN), 
        .B2(keyinput_f127), .ZN(n10153) );
  OAI221_X1 U11228 ( .B1(SI_1_), .B2(keyinput_f31), .C1(P1_D_REG_4__SCAN_IN), 
        .C2(keyinput_f127), .A(n10153), .ZN(n10156) );
  AOI22_X1 U11229 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_f62), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(keyinput_f70), .ZN(n10154) );
  OAI221_X1 U11230 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .C1(
        P2_DATAO_REG_26__SCAN_IN), .C2(keyinput_f70), .A(n10154), .ZN(n10155)
         );
  NOR4_X1 U11231 ( .A1(n10158), .A2(n10157), .A3(n10156), .A4(n10155), .ZN(
        n10159) );
  NAND4_X1 U11232 ( .A1(n10162), .A2(n10161), .A3(n10160), .A4(n10159), .ZN(
        n10245) );
  AOI22_X1 U11233 ( .A1(SI_31_), .A2(keyinput_f1), .B1(P1_IR_REG_0__SCAN_IN), 
        .B2(keyinput_f91), .ZN(n10163) );
  OAI221_X1 U11234 ( .B1(SI_31_), .B2(keyinput_f1), .C1(P1_IR_REG_0__SCAN_IN), 
        .C2(keyinput_f91), .A(n10163), .ZN(n10170) );
  AOI22_X1 U11235 ( .A1(SI_29_), .A2(keyinput_f3), .B1(SI_9_), .B2(
        keyinput_f23), .ZN(n10164) );
  OAI221_X1 U11236 ( .B1(SI_29_), .B2(keyinput_f3), .C1(SI_9_), .C2(
        keyinput_f23), .A(n10164), .ZN(n10169) );
  AOI22_X1 U11237 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput_f45), .B1(
        P1_IR_REG_31__SCAN_IN), .B2(keyinput_f122), .ZN(n10165) );
  OAI221_X1 U11238 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_f45), .C1(
        P1_IR_REG_31__SCAN_IN), .C2(keyinput_f122), .A(n10165), .ZN(n10168) );
  AOI22_X1 U11239 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(keyinput_f67), .B1(
        P2_REG3_REG_5__SCAN_IN), .B2(keyinput_f49), .ZN(n10166) );
  OAI221_X1 U11240 ( .B1(P2_DATAO_REG_29__SCAN_IN), .B2(keyinput_f67), .C1(
        P2_REG3_REG_5__SCAN_IN), .C2(keyinput_f49), .A(n10166), .ZN(n10167) );
  NOR4_X1 U11241 ( .A1(n10170), .A2(n10169), .A3(n10168), .A4(n10167), .ZN(
        n10198) );
  AOI22_X1 U11242 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_f51), .B1(
        P1_IR_REG_4__SCAN_IN), .B2(keyinput_f95), .ZN(n10171) );
  OAI221_X1 U11243 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .C1(
        P1_IR_REG_4__SCAN_IN), .C2(keyinput_f95), .A(n10171), .ZN(n10178) );
  AOI22_X1 U11244 ( .A1(SI_12_), .A2(keyinput_f20), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_f75), .ZN(n10172) );
  OAI221_X1 U11245 ( .B1(SI_12_), .B2(keyinput_f20), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput_f75), .A(n10172), .ZN(n10177)
         );
  AOI22_X1 U11246 ( .A1(SI_13_), .A2(keyinput_f19), .B1(P1_IR_REG_25__SCAN_IN), 
        .B2(keyinput_f116), .ZN(n10173) );
  OAI221_X1 U11247 ( .B1(SI_13_), .B2(keyinput_f19), .C1(P1_IR_REG_25__SCAN_IN), .C2(keyinput_f116), .A(n10173), .ZN(n10176) );
  AOI22_X1 U11248 ( .A1(SI_3_), .A2(keyinput_f29), .B1(P1_IR_REG_21__SCAN_IN), 
        .B2(keyinput_f112), .ZN(n10174) );
  OAI221_X1 U11249 ( .B1(SI_3_), .B2(keyinput_f29), .C1(P1_IR_REG_21__SCAN_IN), 
        .C2(keyinput_f112), .A(n10174), .ZN(n10175) );
  NOR4_X1 U11250 ( .A1(n10178), .A2(n10177), .A3(n10176), .A4(n10175), .ZN(
        n10197) );
  AOI22_X1 U11251 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(keyinput_f71), .B1(
        P1_IR_REG_12__SCAN_IN), .B2(keyinput_f103), .ZN(n10179) );
  OAI221_X1 U11252 ( .B1(P2_DATAO_REG_25__SCAN_IN), .B2(keyinput_f71), .C1(
        P1_IR_REG_12__SCAN_IN), .C2(keyinput_f103), .A(n10179), .ZN(n10186) );
  AOI22_X1 U11253 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_f34), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(keyinput_f72), .ZN(n10180) );
  OAI221_X1 U11254 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_f34), .C1(
        P2_DATAO_REG_24__SCAN_IN), .C2(keyinput_f72), .A(n10180), .ZN(n10185)
         );
  AOI22_X1 U11255 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(keyinput_f82), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(keyinput_f80), .ZN(n10181) );
  OAI221_X1 U11256 ( .B1(P2_DATAO_REG_14__SCAN_IN), .B2(keyinput_f82), .C1(
        P2_DATAO_REG_16__SCAN_IN), .C2(keyinput_f80), .A(n10181), .ZN(n10184)
         );
  AOI22_X1 U11257 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_f60), .B1(
        P1_IR_REG_17__SCAN_IN), .B2(keyinput_f108), .ZN(n10182) );
  OAI221_X1 U11258 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .C1(
        P1_IR_REG_17__SCAN_IN), .C2(keyinput_f108), .A(n10182), .ZN(n10183) );
  NOR4_X1 U11259 ( .A1(n10186), .A2(n10185), .A3(n10184), .A4(n10183), .ZN(
        n10196) );
  AOI22_X1 U11260 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_f61), .B1(SI_23_), .B2(keyinput_f9), .ZN(n10187) );
  OAI221_X1 U11261 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .C1(
        SI_23_), .C2(keyinput_f9), .A(n10187), .ZN(n10194) );
  AOI22_X1 U11262 ( .A1(SI_2_), .A2(keyinput_f30), .B1(SI_26_), .B2(
        keyinput_f6), .ZN(n10188) );
  OAI221_X1 U11263 ( .B1(SI_2_), .B2(keyinput_f30), .C1(SI_26_), .C2(
        keyinput_f6), .A(n10188), .ZN(n10193) );
  AOI22_X1 U11264 ( .A1(SI_17_), .A2(keyinput_f15), .B1(P1_IR_REG_6__SCAN_IN), 
        .B2(keyinput_f97), .ZN(n10189) );
  OAI221_X1 U11265 ( .B1(SI_17_), .B2(keyinput_f15), .C1(P1_IR_REG_6__SCAN_IN), 
        .C2(keyinput_f97), .A(n10189), .ZN(n10192) );
  AOI22_X1 U11266 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_f44), .B1(SI_25_), .B2(keyinput_f7), .ZN(n10190) );
  OAI221_X1 U11267 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .C1(
        SI_25_), .C2(keyinput_f7), .A(n10190), .ZN(n10191) );
  NOR4_X1 U11268 ( .A1(n10194), .A2(n10193), .A3(n10192), .A4(n10191), .ZN(
        n10195) );
  NAND4_X1 U11269 ( .A1(n10198), .A2(n10197), .A3(n10196), .A4(n10195), .ZN(
        n10244) );
  AOI22_X1 U11270 ( .A1(n10416), .A2(keyinput_f65), .B1(n7465), .B2(
        keyinput_f40), .ZN(n10199) );
  OAI221_X1 U11271 ( .B1(n10416), .B2(keyinput_f65), .C1(n7465), .C2(
        keyinput_f40), .A(n10199), .ZN(n10208) );
  INV_X1 U11272 ( .A(SI_24_), .ZN(n10319) );
  AOI22_X1 U11273 ( .A1(n10319), .A2(keyinput_f8), .B1(keyinput_f63), .B2(
        n5540), .ZN(n10200) );
  OAI221_X1 U11274 ( .B1(n10319), .B2(keyinput_f8), .C1(n5540), .C2(
        keyinput_f63), .A(n10200), .ZN(n10207) );
  AOI22_X1 U11275 ( .A1(n6031), .A2(keyinput_f114), .B1(keyinput_f22), .B2(
        n10202), .ZN(n10201) );
  OAI221_X1 U11276 ( .B1(n6031), .B2(keyinput_f114), .C1(n10202), .C2(
        keyinput_f22), .A(n10201), .ZN(n10206) );
  XNOR2_X1 U11277 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_f99), .ZN(n10204) );
  XNOR2_X1 U11278 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput_f69), .ZN(n10203) );
  NAND2_X1 U11279 ( .A1(n10204), .A2(n10203), .ZN(n10205) );
  NOR4_X1 U11280 ( .A1(n10208), .A2(n10207), .A3(n10206), .A4(n10205), .ZN(
        n10242) );
  AOI22_X1 U11281 ( .A1(n10347), .A2(keyinput_f55), .B1(n10419), .B2(
        keyinput_f76), .ZN(n10209) );
  OAI221_X1 U11282 ( .B1(n10347), .B2(keyinput_f55), .C1(n10419), .C2(
        keyinput_f76), .A(n10209), .ZN(n10217) );
  AOI22_X1 U11283 ( .A1(n10390), .A2(keyinput_f4), .B1(keyinput_f56), .B2(
        n5497), .ZN(n10210) );
  OAI221_X1 U11284 ( .B1(n10390), .B2(keyinput_f4), .C1(n5497), .C2(
        keyinput_f56), .A(n10210), .ZN(n10216) );
  INV_X1 U11285 ( .A(SI_7_), .ZN(n10392) );
  AOI22_X1 U11286 ( .A1(n10318), .A2(keyinput_f37), .B1(n10392), .B2(
        keyinput_f25), .ZN(n10211) );
  OAI221_X1 U11287 ( .B1(n10318), .B2(keyinput_f37), .C1(n10392), .C2(
        keyinput_f25), .A(n10211), .ZN(n10215) );
  INV_X1 U11288 ( .A(SI_14_), .ZN(n10414) );
  AOI22_X1 U11289 ( .A1(n10414), .A2(keyinput_f18), .B1(n10213), .B2(
        keyinput_f81), .ZN(n10212) );
  OAI221_X1 U11290 ( .B1(n10414), .B2(keyinput_f18), .C1(n10213), .C2(
        keyinput_f81), .A(n10212), .ZN(n10214) );
  NOR4_X1 U11291 ( .A1(n10217), .A2(n10216), .A3(n10215), .A4(n10214), .ZN(
        n10241) );
  INV_X1 U11292 ( .A(SI_21_), .ZN(n10219) );
  AOI22_X1 U11293 ( .A1(n10219), .A2(keyinput_f11), .B1(keyinput_f17), .B2(
        n10348), .ZN(n10218) );
  OAI221_X1 U11294 ( .B1(n10219), .B2(keyinput_f11), .C1(n10348), .C2(
        keyinput_f17), .A(n10218), .ZN(n10227) );
  XNOR2_X1 U11295 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_f113), .ZN(n10223)
         );
  XNOR2_X1 U11296 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_f84), .ZN(n10222) );
  XNOR2_X1 U11297 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_f104), .ZN(n10221)
         );
  XNOR2_X1 U11298 ( .A(SI_8_), .B(keyinput_f24), .ZN(n10220) );
  NAND4_X1 U11299 ( .A1(n10223), .A2(n10222), .A3(n10221), .A4(n10220), .ZN(
        n10226) );
  XNOR2_X1 U11300 ( .A(n10403), .B(keyinput_f110), .ZN(n10225) );
  XNOR2_X1 U11301 ( .A(n10343), .B(keyinput_f10), .ZN(n10224) );
  NOR4_X1 U11302 ( .A1(n10227), .A2(n10226), .A3(n10225), .A4(n10224), .ZN(
        n10240) );
  AOI22_X1 U11303 ( .A1(n10316), .A2(keyinput_f83), .B1(keyinput_f52), .B2(
        n5337), .ZN(n10228) );
  OAI221_X1 U11304 ( .B1(n10316), .B2(keyinput_f83), .C1(n5337), .C2(
        keyinput_f52), .A(n10228), .ZN(n10238) );
  INV_X1 U11305 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10429) );
  AOI22_X1 U11306 ( .A1(n10230), .A2(keyinput_f86), .B1(n10429), .B2(
        keyinput_f124), .ZN(n10229) );
  OAI221_X1 U11307 ( .B1(n10230), .B2(keyinput_f86), .C1(n10429), .C2(
        keyinput_f124), .A(n10229), .ZN(n10237) );
  AOI22_X1 U11308 ( .A1(n10232), .A2(keyinput_f89), .B1(n6020), .B2(
        keyinput_f93), .ZN(n10231) );
  OAI221_X1 U11309 ( .B1(n10232), .B2(keyinput_f89), .C1(n6020), .C2(
        keyinput_f93), .A(n10231), .ZN(n10236) );
  XNOR2_X1 U11310 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_f106), .ZN(n10234)
         );
  XNOR2_X1 U11311 ( .A(SI_5_), .B(keyinput_f27), .ZN(n10233) );
  NAND2_X1 U11312 ( .A1(n10234), .A2(n10233), .ZN(n10235) );
  NOR4_X1 U11313 ( .A1(n10238), .A2(n10237), .A3(n10236), .A4(n10235), .ZN(
        n10239) );
  NAND4_X1 U11314 ( .A1(n10242), .A2(n10241), .A3(n10240), .A4(n10239), .ZN(
        n10243) );
  NOR4_X1 U11315 ( .A1(n10246), .A2(n10245), .A3(n10244), .A4(n10243), .ZN(
        n10247) );
  NAND4_X1 U11316 ( .A1(n10250), .A2(n10249), .A3(n10248), .A4(n10247), .ZN(
        n10252) );
  AOI21_X1 U11317 ( .B1(keyinput_f28), .B2(n10252), .A(keyinput_g28), .ZN(
        n10254) );
  INV_X1 U11318 ( .A(keyinput_f28), .ZN(n10251) );
  AOI21_X1 U11319 ( .B1(n10252), .B2(n10251), .A(n10255), .ZN(n10253) );
  AOI22_X1 U11320 ( .A1(n10255), .A2(n10254), .B1(keyinput_g28), .B2(n10253), 
        .ZN(n10449) );
  XOR2_X1 U11321 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_g113), .Z(n10262) );
  AOI22_X1 U11322 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(keyinput_g66), .B1(
        P1_D_REG_2__SCAN_IN), .B2(keyinput_g125), .ZN(n10256) );
  OAI221_X1 U11323 ( .B1(P2_DATAO_REG_30__SCAN_IN), .B2(keyinput_g66), .C1(
        P1_D_REG_2__SCAN_IN), .C2(keyinput_g125), .A(n10256), .ZN(n10261) );
  AOI22_X1 U11324 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(keyinput_g67), .B1(
        SI_16_), .B2(keyinput_g16), .ZN(n10257) );
  OAI221_X1 U11325 ( .B1(P2_DATAO_REG_29__SCAN_IN), .B2(keyinput_g67), .C1(
        SI_16_), .C2(keyinput_g16), .A(n10257), .ZN(n10260) );
  AOI22_X1 U11326 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(keyinput_g84), .B1(
        P1_IR_REG_4__SCAN_IN), .B2(keyinput_g95), .ZN(n10258) );
  OAI221_X1 U11327 ( .B1(P2_DATAO_REG_12__SCAN_IN), .B2(keyinput_g84), .C1(
        P1_IR_REG_4__SCAN_IN), .C2(keyinput_g95), .A(n10258), .ZN(n10259) );
  NOR4_X1 U11328 ( .A1(n10262), .A2(n10261), .A3(n10260), .A4(n10259), .ZN(
        n10290) );
  AOI22_X1 U11329 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(keyinput_g85), .B1(
        SI_11_), .B2(keyinput_g21), .ZN(n10263) );
  OAI221_X1 U11330 ( .B1(P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_g85), .C1(
        SI_11_), .C2(keyinput_g21), .A(n10263), .ZN(n10270) );
  AOI22_X1 U11331 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(keyinput_g70), .B1(
        P1_IR_REG_26__SCAN_IN), .B2(keyinput_g117), .ZN(n10264) );
  OAI221_X1 U11332 ( .B1(P2_DATAO_REG_26__SCAN_IN), .B2(keyinput_g70), .C1(
        P1_IR_REG_26__SCAN_IN), .C2(keyinput_g117), .A(n10264), .ZN(n10269) );
  AOI22_X1 U11333 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(keyinput_g72), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(keyinput_g71), .ZN(n10265) );
  OAI221_X1 U11334 ( .B1(P2_DATAO_REG_24__SCAN_IN), .B2(keyinput_g72), .C1(
        P2_DATAO_REG_25__SCAN_IN), .C2(keyinput_g71), .A(n10265), .ZN(n10268)
         );
  AOI22_X1 U11335 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput_g87), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(keyinput_g82), .ZN(n10266) );
  OAI221_X1 U11336 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_g87), .C1(
        P2_DATAO_REG_14__SCAN_IN), .C2(keyinput_g82), .A(n10266), .ZN(n10267)
         );
  NOR4_X1 U11337 ( .A1(n10270), .A2(n10269), .A3(n10268), .A4(n10267), .ZN(
        n10289) );
  AOI22_X1 U11338 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_g46), .B1(
        P1_IR_REG_8__SCAN_IN), .B2(keyinput_g99), .ZN(n10271) );
  OAI221_X1 U11339 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .C1(
        P1_IR_REG_8__SCAN_IN), .C2(keyinput_g99), .A(n10271), .ZN(n10278) );
  AOI22_X1 U11340 ( .A1(P1_D_REG_4__SCAN_IN), .A2(keyinput_g127), .B1(
        P1_IR_REG_16__SCAN_IN), .B2(keyinput_g107), .ZN(n10272) );
  OAI221_X1 U11341 ( .B1(P1_D_REG_4__SCAN_IN), .B2(keyinput_g127), .C1(
        P1_IR_REG_16__SCAN_IN), .C2(keyinput_g107), .A(n10272), .ZN(n10277) );
  AOI22_X1 U11342 ( .A1(SI_10_), .A2(keyinput_g22), .B1(P1_IR_REG_28__SCAN_IN), 
        .B2(keyinput_g119), .ZN(n10273) );
  OAI221_X1 U11343 ( .B1(SI_10_), .B2(keyinput_g22), .C1(P1_IR_REG_28__SCAN_IN), .C2(keyinput_g119), .A(n10273), .ZN(n10276) );
  AOI22_X1 U11344 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(keyinput_g81), .B1(
        SI_21_), .B2(keyinput_g11), .ZN(n10274) );
  OAI221_X1 U11345 ( .B1(P2_DATAO_REG_15__SCAN_IN), .B2(keyinput_g81), .C1(
        SI_21_), .C2(keyinput_g11), .A(n10274), .ZN(n10275) );
  NOR4_X1 U11346 ( .A1(n10278), .A2(n10277), .A3(n10276), .A4(n10275), .ZN(
        n10288) );
  AOI22_X1 U11347 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(keyinput_g80), .B1(
        P1_IR_REG_5__SCAN_IN), .B2(keyinput_g96), .ZN(n10279) );
  OAI221_X1 U11348 ( .B1(P2_DATAO_REG_16__SCAN_IN), .B2(keyinput_g80), .C1(
        P1_IR_REG_5__SCAN_IN), .C2(keyinput_g96), .A(n10279), .ZN(n10286) );
  AOI22_X1 U11349 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(keyinput_g79), .B1(
        P1_IR_REG_2__SCAN_IN), .B2(keyinput_g93), .ZN(n10280) );
  OAI221_X1 U11350 ( .B1(P2_DATAO_REG_17__SCAN_IN), .B2(keyinput_g79), .C1(
        P1_IR_REG_2__SCAN_IN), .C2(keyinput_g93), .A(n10280), .ZN(n10285) );
  AOI22_X1 U11351 ( .A1(SI_29_), .A2(keyinput_g3), .B1(SI_17_), .B2(
        keyinput_g15), .ZN(n10281) );
  OAI221_X1 U11352 ( .B1(SI_29_), .B2(keyinput_g3), .C1(SI_17_), .C2(
        keyinput_g15), .A(n10281), .ZN(n10284) );
  AOI22_X1 U11353 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput_g88), .B1(
        SI_12_), .B2(keyinput_g20), .ZN(n10282) );
  OAI221_X1 U11354 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_g88), .C1(
        SI_12_), .C2(keyinput_g20), .A(n10282), .ZN(n10283) );
  NOR4_X1 U11355 ( .A1(n10286), .A2(n10285), .A3(n10284), .A4(n10283), .ZN(
        n10287) );
  NAND4_X1 U11356 ( .A1(n10290), .A2(n10289), .A3(n10288), .A4(n10287), .ZN(
        n10447) );
  AOI22_X1 U11357 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(keyinput_g75), .B1(
        P1_IR_REG_10__SCAN_IN), .B2(keyinput_g101), .ZN(n10291) );
  OAI221_X1 U11358 ( .B1(P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_g75), .C1(
        P1_IR_REG_10__SCAN_IN), .C2(keyinput_g101), .A(n10291), .ZN(n10298) );
  AOI22_X1 U11359 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(keyinput_g90), .B1(
        P1_D_REG_3__SCAN_IN), .B2(keyinput_g126), .ZN(n10292) );
  OAI221_X1 U11360 ( .B1(P2_DATAO_REG_6__SCAN_IN), .B2(keyinput_g90), .C1(
        P1_D_REG_3__SCAN_IN), .C2(keyinput_g126), .A(n10292), .ZN(n10297) );
  AOI22_X1 U11361 ( .A1(SI_30_), .A2(keyinput_g2), .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_g38), .ZN(n10293) );
  OAI221_X1 U11362 ( .B1(SI_30_), .B2(keyinput_g2), .C1(
        P2_REG3_REG_23__SCAN_IN), .C2(keyinput_g38), .A(n10293), .ZN(n10296)
         );
  AOI22_X1 U11363 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_g61), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(keyinput_g86), .ZN(n10294) );
  OAI221_X1 U11364 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .C1(
        P2_DATAO_REG_10__SCAN_IN), .C2(keyinput_g86), .A(n10294), .ZN(n10295)
         );
  NOR4_X1 U11365 ( .A1(n10298), .A2(n10297), .A3(n10296), .A4(n10295), .ZN(
        n10330) );
  AOI22_X1 U11366 ( .A1(SI_23_), .A2(keyinput_g9), .B1(P1_IR_REG_11__SCAN_IN), 
        .B2(keyinput_g102), .ZN(n10299) );
  OAI221_X1 U11367 ( .B1(SI_23_), .B2(keyinput_g9), .C1(P1_IR_REG_11__SCAN_IN), 
        .C2(keyinput_g102), .A(n10299), .ZN(n10306) );
  AOI22_X1 U11368 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_g57), .B1(
        P1_IR_REG_7__SCAN_IN), .B2(keyinput_g98), .ZN(n10300) );
  OAI221_X1 U11369 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .C1(
        P1_IR_REG_7__SCAN_IN), .C2(keyinput_g98), .A(n10300), .ZN(n10305) );
  AOI22_X1 U11370 ( .A1(SI_25_), .A2(keyinput_g7), .B1(P1_IR_REG_13__SCAN_IN), 
        .B2(keyinput_g104), .ZN(n10301) );
  OAI221_X1 U11371 ( .B1(SI_25_), .B2(keyinput_g7), .C1(P1_IR_REG_13__SCAN_IN), 
        .C2(keyinput_g104), .A(n10301), .ZN(n10304) );
  AOI22_X1 U11372 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_g39), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput_g34), .ZN(n10302) );
  OAI221_X1 U11373 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput_g34), .A(n10302), .ZN(n10303) );
  NOR4_X1 U11374 ( .A1(n10306), .A2(n10305), .A3(n10304), .A4(n10303), .ZN(
        n10329) );
  AOI22_X1 U11375 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(keyinput_g74), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(keyinput_g69), .ZN(n10307) );
  OAI221_X1 U11376 ( .B1(P2_DATAO_REG_22__SCAN_IN), .B2(keyinput_g74), .C1(
        P2_DATAO_REG_27__SCAN_IN), .C2(keyinput_g69), .A(n10307), .ZN(n10314)
         );
  AOI22_X1 U11377 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .ZN(n10308) );
  OAI221_X1 U11378 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput_g63), .A(n10308), .ZN(n10313)
         );
  AOI22_X1 U11379 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput_g41), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(keyinput_g68), .ZN(n10309) );
  OAI221_X1 U11380 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .C1(
        P2_DATAO_REG_28__SCAN_IN), .C2(keyinput_g68), .A(n10309), .ZN(n10312)
         );
  AOI22_X1 U11381 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(keyinput_g35), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .ZN(n10310) );
  OAI221_X1 U11382 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_g35), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_g62), .A(n10310), .ZN(n10311)
         );
  NOR4_X1 U11383 ( .A1(n10314), .A2(n10313), .A3(n10312), .A4(n10311), .ZN(
        n10328) );
  AOI22_X1 U11384 ( .A1(n8471), .A2(keyinput_g45), .B1(n10316), .B2(
        keyinput_g83), .ZN(n10315) );
  OAI221_X1 U11385 ( .B1(n8471), .B2(keyinput_g45), .C1(n10316), .C2(
        keyinput_g83), .A(n10315), .ZN(n10326) );
  AOI22_X1 U11386 ( .A1(n6055), .A2(keyinput_g115), .B1(keyinput_g37), .B2(
        n10318), .ZN(n10317) );
  OAI221_X1 U11387 ( .B1(n6055), .B2(keyinput_g115), .C1(n10318), .C2(
        keyinput_g37), .A(n10317), .ZN(n10325) );
  XOR2_X1 U11388 ( .A(n6031), .B(keyinput_g114), .Z(n10323) );
  XOR2_X1 U11389 ( .A(n10319), .B(keyinput_g8), .Z(n10322) );
  XNOR2_X1 U11390 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_g103), .ZN(n10321)
         );
  XNOR2_X1 U11391 ( .A(SI_2_), .B(keyinput_g30), .ZN(n10320) );
  NAND4_X1 U11392 ( .A1(n10323), .A2(n10322), .A3(n10321), .A4(n10320), .ZN(
        n10324) );
  NOR3_X1 U11393 ( .A1(n10326), .A2(n10325), .A3(n10324), .ZN(n10327) );
  NAND4_X1 U11394 ( .A1(n10330), .A2(n10329), .A3(n10328), .A4(n10327), .ZN(
        n10446) );
  INV_X1 U11395 ( .A(P2_B_REG_SCAN_IN), .ZN(n10332) );
  AOI22_X1 U11396 ( .A1(n10332), .A2(keyinput_g64), .B1(keyinput_g42), .B2(
        n5796), .ZN(n10331) );
  OAI221_X1 U11397 ( .B1(n10332), .B2(keyinput_g64), .C1(n5796), .C2(
        keyinput_g42), .A(n10331), .ZN(n10341) );
  INV_X1 U11398 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10334) );
  AOI22_X1 U11399 ( .A1(n5572), .A2(keyinput_g50), .B1(keyinput_g49), .B2(
        n10334), .ZN(n10333) );
  OAI221_X1 U11400 ( .B1(n5572), .B2(keyinput_g50), .C1(n10334), .C2(
        keyinput_g49), .A(n10333), .ZN(n10340) );
  XOR2_X1 U11401 ( .A(n7139), .B(keyinput_g44), .Z(n10338) );
  XNOR2_X1 U11402 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_g89), .ZN(n10337)
         );
  XNOR2_X1 U11403 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_g116), .ZN(n10336)
         );
  XNOR2_X1 U11404 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_g105), .ZN(n10335)
         );
  NAND4_X1 U11405 ( .A1(n10338), .A2(n10337), .A3(n10336), .A4(n10335), .ZN(
        n10339) );
  NOR3_X1 U11406 ( .A1(n10341), .A2(n10340), .A3(n10339), .ZN(n10385) );
  AOI22_X1 U11407 ( .A1(n10343), .A2(keyinput_g10), .B1(keyinput_g121), .B2(
        n4754), .ZN(n10342) );
  OAI221_X1 U11408 ( .B1(n10343), .B2(keyinput_g10), .C1(n4754), .C2(
        keyinput_g121), .A(n10342), .ZN(n10354) );
  AOI22_X1 U11409 ( .A1(n5497), .A2(keyinput_g56), .B1(n10345), .B2(
        keyinput_g19), .ZN(n10344) );
  OAI221_X1 U11410 ( .B1(n5497), .B2(keyinput_g56), .C1(n10345), .C2(
        keyinput_g19), .A(n10344), .ZN(n10353) );
  AOI22_X1 U11411 ( .A1(n10348), .A2(keyinput_g17), .B1(keyinput_g55), .B2(
        n10347), .ZN(n10346) );
  OAI221_X1 U11412 ( .B1(n10348), .B2(keyinput_g17), .C1(n10347), .C2(
        keyinput_g55), .A(n10346), .ZN(n10352) );
  XNOR2_X1 U11413 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_g97), .ZN(n10350) );
  XNOR2_X1 U11414 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_g36), .ZN(n10349)
         );
  NAND2_X1 U11415 ( .A1(n10350), .A2(n10349), .ZN(n10351) );
  NOR4_X1 U11416 ( .A1(n10354), .A2(n10353), .A3(n10352), .A4(n10351), .ZN(
        n10384) );
  AOI22_X1 U11417 ( .A1(n6044), .A2(keyinput_g111), .B1(keyinput_g58), .B2(
        n10356), .ZN(n10355) );
  OAI221_X1 U11418 ( .B1(n6044), .B2(keyinput_g111), .C1(n10356), .C2(
        keyinput_g58), .A(n10355), .ZN(n10367) );
  INV_X1 U11419 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10359) );
  AOI22_X1 U11420 ( .A1(n10359), .A2(keyinput_g123), .B1(keyinput_g6), .B2(
        n10358), .ZN(n10357) );
  OAI221_X1 U11421 ( .B1(n10359), .B2(keyinput_g123), .C1(n10358), .C2(
        keyinput_g6), .A(n10357), .ZN(n10366) );
  AOI22_X1 U11422 ( .A1(n6428), .A2(keyinput_g108), .B1(keyinput_g51), .B2(
        n10361), .ZN(n10360) );
  OAI221_X1 U11423 ( .B1(n6428), .B2(keyinput_g108), .C1(n10361), .C2(
        keyinput_g51), .A(n10360), .ZN(n10365) );
  XNOR2_X1 U11424 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_g106), .ZN(n10363)
         );
  XNOR2_X1 U11425 ( .A(SI_1_), .B(keyinput_g31), .ZN(n10362) );
  NAND2_X1 U11426 ( .A1(n10363), .A2(n10362), .ZN(n10364) );
  NOR4_X1 U11427 ( .A1(n10367), .A2(n10366), .A3(n10365), .A4(n10364), .ZN(
        n10383) );
  AOI22_X1 U11428 ( .A1(n5337), .A2(keyinput_g52), .B1(n10369), .B2(
        keyinput_g92), .ZN(n10368) );
  OAI221_X1 U11429 ( .B1(n5337), .B2(keyinput_g52), .C1(n10369), .C2(
        keyinput_g92), .A(n10368), .ZN(n10381) );
  INV_X1 U11430 ( .A(P2_WR_REG_SCAN_IN), .ZN(n10372) );
  AOI22_X1 U11431 ( .A1(n10372), .A2(keyinput_g0), .B1(n10371), .B2(
        keyinput_g29), .ZN(n10370) );
  OAI221_X1 U11432 ( .B1(n10372), .B2(keyinput_g0), .C1(n10371), .C2(
        keyinput_g29), .A(n10370), .ZN(n10380) );
  AOI22_X1 U11433 ( .A1(n10375), .A2(keyinput_g77), .B1(keyinput_g43), .B2(
        n10374), .ZN(n10373) );
  OAI221_X1 U11434 ( .B1(n10375), .B2(keyinput_g77), .C1(n10374), .C2(
        keyinput_g43), .A(n10373), .ZN(n10379) );
  XNOR2_X1 U11435 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_g100), .ZN(n10377)
         );
  XNOR2_X1 U11436 ( .A(SI_6_), .B(keyinput_g26), .ZN(n10376) );
  NAND2_X1 U11437 ( .A1(n10377), .A2(n10376), .ZN(n10378) );
  NOR4_X1 U11438 ( .A1(n10381), .A2(n10380), .A3(n10379), .A4(n10378), .ZN(
        n10382) );
  NAND4_X1 U11439 ( .A1(n10385), .A2(n10384), .A3(n10383), .A4(n10382), .ZN(
        n10445) );
  AOI22_X1 U11440 ( .A1(n5423), .A2(keyinput_g53), .B1(n10387), .B2(
        keyinput_g5), .ZN(n10386) );
  OAI221_X1 U11441 ( .B1(n5423), .B2(keyinput_g53), .C1(n10387), .C2(
        keyinput_g5), .A(n10386), .ZN(n10399) );
  AOI22_X1 U11442 ( .A1(n10390), .A2(keyinput_g4), .B1(n10389), .B2(
        keyinput_g12), .ZN(n10388) );
  OAI221_X1 U11443 ( .B1(n10390), .B2(keyinput_g4), .C1(n10389), .C2(
        keyinput_g12), .A(n10388), .ZN(n10398) );
  AOI22_X1 U11444 ( .A1(n7465), .A2(keyinput_g40), .B1(n10392), .B2(
        keyinput_g25), .ZN(n10391) );
  OAI221_X1 U11445 ( .B1(n7465), .B2(keyinput_g40), .C1(n10392), .C2(
        keyinput_g25), .A(n10391), .ZN(n10397) );
  INV_X1 U11446 ( .A(SI_31_), .ZN(n10395) );
  AOI22_X1 U11447 ( .A1(n10395), .A2(keyinput_g1), .B1(n10394), .B2(
        keyinput_g54), .ZN(n10393) );
  OAI221_X1 U11448 ( .B1(n10395), .B2(keyinput_g1), .C1(n10394), .C2(
        keyinput_g54), .A(n10393), .ZN(n10396) );
  NOR4_X1 U11449 ( .A1(n10399), .A2(n10398), .A3(n10397), .A4(n10396), .ZN(
        n10443) );
  AOI22_X1 U11450 ( .A1(n10402), .A2(keyinput_g73), .B1(keyinput_g78), .B2(
        n10401), .ZN(n10400) );
  OAI221_X1 U11451 ( .B1(n10402), .B2(keyinput_g73), .C1(n10401), .C2(
        keyinput_g78), .A(n10400), .ZN(n10411) );
  XNOR2_X1 U11452 ( .A(n10403), .B(keyinput_g110), .ZN(n10410) );
  XNOR2_X1 U11453 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_g94), .ZN(n10407) );
  XNOR2_X1 U11454 ( .A(SI_0_), .B(keyinput_g32), .ZN(n10406) );
  XNOR2_X1 U11455 ( .A(SI_19_), .B(keyinput_g13), .ZN(n10405) );
  XNOR2_X1 U11456 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_g112), .ZN(n10404)
         );
  NAND4_X1 U11457 ( .A1(n10407), .A2(n10406), .A3(n10405), .A4(n10404), .ZN(
        n10409) );
  XNOR2_X1 U11458 ( .A(keyinput_g47), .B(n5694), .ZN(n10408) );
  NOR4_X1 U11459 ( .A1(n10411), .A2(n10410), .A3(n10409), .A4(n10408), .ZN(
        n10442) );
  AOI22_X1 U11460 ( .A1(n10414), .A2(keyinput_g18), .B1(keyinput_g27), .B2(
        n10413), .ZN(n10412) );
  OAI221_X1 U11461 ( .B1(n10414), .B2(keyinput_g18), .C1(n10413), .C2(
        keyinput_g27), .A(n10412), .ZN(n10425) );
  AOI22_X1 U11462 ( .A1(n10416), .A2(keyinput_g65), .B1(n4620), .B2(
        keyinput_g33), .ZN(n10415) );
  OAI221_X1 U11463 ( .B1(n10416), .B2(keyinput_g65), .C1(n4620), .C2(
        keyinput_g33), .A(n10415), .ZN(n10424) );
  AOI22_X1 U11464 ( .A1(n10419), .A2(keyinput_g76), .B1(keyinput_g23), .B2(
        n10418), .ZN(n10417) );
  OAI221_X1 U11465 ( .B1(n10419), .B2(keyinput_g76), .C1(n10418), .C2(
        keyinput_g23), .A(n10417), .ZN(n10423) );
  XOR2_X1 U11466 ( .A(n6033), .B(keyinput_g120), .Z(n10421) );
  XNOR2_X1 U11467 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_g122), .ZN(n10420)
         );
  NAND2_X1 U11468 ( .A1(n10421), .A2(n10420), .ZN(n10422) );
  NOR4_X1 U11469 ( .A1(n10425), .A2(n10424), .A3(n10423), .A4(n10422), .ZN(
        n10441) );
  AOI22_X1 U11470 ( .A1(n6063), .A2(keyinput_g118), .B1(keyinput_g60), .B2(
        n10427), .ZN(n10426) );
  OAI221_X1 U11471 ( .B1(n6063), .B2(keyinput_g118), .C1(n10427), .C2(
        keyinput_g60), .A(n10426), .ZN(n10439) );
  AOI22_X1 U11472 ( .A1(n10430), .A2(keyinput_g24), .B1(n10429), .B2(
        keyinput_g124), .ZN(n10428) );
  OAI221_X1 U11473 ( .B1(n10430), .B2(keyinput_g24), .C1(n10429), .C2(
        keyinput_g124), .A(n10428), .ZN(n10438) );
  AOI22_X1 U11474 ( .A1(n10433), .A2(keyinput_g91), .B1(keyinput_g14), .B2(
        n10432), .ZN(n10431) );
  OAI221_X1 U11475 ( .B1(n10433), .B2(keyinput_g91), .C1(n10432), .C2(
        keyinput_g14), .A(n10431), .ZN(n10437) );
  AOI22_X1 U11476 ( .A1(n6043), .A2(keyinput_g109), .B1(keyinput_g48), .B2(
        n10435), .ZN(n10434) );
  OAI221_X1 U11477 ( .B1(n6043), .B2(keyinput_g109), .C1(n10435), .C2(
        keyinput_g48), .A(n10434), .ZN(n10436) );
  NOR4_X1 U11478 ( .A1(n10439), .A2(n10438), .A3(n10437), .A4(n10436), .ZN(
        n10440) );
  NAND4_X1 U11479 ( .A1(n10443), .A2(n10442), .A3(n10441), .A4(n10440), .ZN(
        n10444) );
  NOR4_X1 U11480 ( .A1(n10447), .A2(n10446), .A3(n10445), .A4(n10444), .ZN(
        n10448) );
  NOR2_X1 U11481 ( .A1(n10449), .A2(n10448), .ZN(n10455) );
  NOR2_X1 U11482 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(P2_ADDR_REG_18__SCAN_IN), 
        .ZN(n10450) );
  AOI21_X1 U11483 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(P1_ADDR_REG_18__SCAN_IN), 
        .A(n10450), .ZN(n10470) );
  OAI21_X1 U11484 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10451), .ZN(n10469) );
  NAND2_X1 U11485 ( .A1(n10470), .A2(n10469), .ZN(n10468) );
  OAI21_X1 U11486 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(P2_ADDR_REG_18__SCAN_IN), 
        .A(n10468), .ZN(n10453) );
  XNOR2_X1 U11487 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n10452) );
  XNOR2_X1 U11488 ( .A(n10453), .B(n10452), .ZN(n10454) );
  XNOR2_X1 U11489 ( .A(n10455), .B(n10454), .ZN(ADD_1071_U4) );
  OAI21_X1 U11490 ( .B1(n10458), .B2(n10457), .A(n10456), .ZN(ADD_1071_U47) );
  OAI21_X1 U11491 ( .B1(n10461), .B2(n10460), .A(n10459), .ZN(ADD_1071_U49) );
  AOI21_X1 U11492 ( .B1(n10464), .B2(n10463), .A(n10462), .ZN(ADD_1071_U54) );
  OAI21_X1 U11493 ( .B1(n10467), .B2(n10466), .A(n10465), .ZN(ADD_1071_U51) );
  OAI21_X1 U11494 ( .B1(n10470), .B2(n10469), .A(n10468), .ZN(ADD_1071_U55) );
  OAI21_X1 U11495 ( .B1(n10473), .B2(n10472), .A(n10471), .ZN(ADD_1071_U48) );
  OAI21_X1 U11496 ( .B1(n10476), .B2(n10475), .A(n10474), .ZN(ADD_1071_U50) );
  AOI21_X1 U11497 ( .B1(n10479), .B2(n10478), .A(n10477), .ZN(ADD_1071_U53) );
  OAI21_X1 U11498 ( .B1(n10482), .B2(n10481), .A(n10480), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4994 ( .A(n6118), .Z(n4484) );
  CLKBUF_X1 U4997 ( .A(n6118), .Z(n4482) );
  CLKBUF_X1 U4998 ( .A(n6118), .Z(n4486) );
  CLKBUF_X1 U4999 ( .A(n5313), .Z(n6945) );
  NAND2_X1 U5022 ( .A1(n9537), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4755) );
endmodule

