

module b20_C_SARLock_k_128_2 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, 
        ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, 
        ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, 
        ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, 
        U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, 
        P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, 
        P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, 
        P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, 
        P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, 
        P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, 
        P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, 
        P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, 
        P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, 
        P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, 
        P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, 
        P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, 
        P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, 
        P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, 
        P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, 
        P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, 
        P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, 
        P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, 
        P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, 
        P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, 
        P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, 
        P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, 
        P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, 
        P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, 
        P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, 
        P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, 
        P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, 
        P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, 
        P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, 
        P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4451, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322;

  INV_X1 U4958 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  XNOR2_X1 U4959 ( .A(n5508), .B(n5506), .ZN(n8904) );
  INV_X1 U4960 ( .A(n8077), .ZN(n8334) );
  OR2_X1 U4961 ( .A1(n10090), .A2(n7613), .ZN(n7615) );
  INV_X1 U4962 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8876) );
  NAND2_X1 U4963 ( .A1(n7433), .A2(n9294), .ZN(n6969) );
  MUX2_X1 U4964 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6004), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n6005) );
  XNOR2_X1 U4965 ( .A(n5069), .B(n5068), .ZN(n5073) );
  CLKBUF_X1 U4966 ( .A(n9032), .Z(n4451) );
  OAI21_X1 U4967 ( .B1(n5881), .B2(n7236), .A(n9893), .ZN(n9032) );
  INV_X1 U4970 ( .A(P1_STATE_REG_SCAN_IN), .ZN(n4454) );
  CLKBUF_X2 U4971 ( .A(n5286), .Z(n5631) );
  NOR2_X1 U4972 ( .A1(n10084), .A2(n10248), .ZN(n7612) );
  INV_X2 U4973 ( .A(n5781), .ZN(n5866) );
  INV_X1 U4974 ( .A(n7090), .ZN(n7091) );
  BUF_X1 U4975 ( .A(n6017), .Z(n4460) );
  OR2_X1 U4976 ( .A1(n8164), .A2(n8165), .ZN(n4962) );
  AOI21_X1 U4977 ( .B1(n4815), .B2(n4465), .A(n4477), .ZN(n8324) );
  NOR2_X1 U4978 ( .A1(n8397), .A2(n5012), .ZN(n8396) );
  XNOR2_X1 U4979 ( .A(n5199), .B(n5197), .ZN(n7103) );
  AND3_X1 U4980 ( .A1(n4596), .A2(n4592), .A3(n6679), .ZN(n6597) );
  BUF_X1 U4981 ( .A(n5144), .Z(n6585) );
  INV_X1 U4982 ( .A(n5248), .ZN(n5886) );
  AND3_X1 U4983 ( .A1(n5246), .A2(n5245), .A3(n5244), .ZN(n9953) );
  AND4_X1 U4984 ( .A1(n6023), .A2(n6022), .A3(n6021), .A4(n6020), .ZN(n7121)
         );
  NAND3_X1 U4985 ( .A1(n5833), .A2(n5834), .A3(n5830), .ZN(n6848) );
  NAND2_X1 U4986 ( .A1(n9551), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5069) );
  AND2_X1 U4987 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7222) );
  INV_X1 U4988 ( .A(n9520), .ZN(n9405) );
  INV_X1 U4989 ( .A(n5187), .ZN(n5247) );
  INV_X1 U4990 ( .A(n5286), .ZN(n5678) );
  NAND2_X2 U4991 ( .A1(n8089), .A2(n7044), .ZN(n6406) );
  NAND2_X2 U4992 ( .A1(n8156), .A2(n8174), .ZN(n8163) );
  NAND2_X1 U4993 ( .A1(n5121), .A2(n6848), .ZN(n4455) );
  XNOR2_X2 U4994 ( .A(n7665), .B(n7666), .ZN(n7616) );
  NOR2_X2 U4995 ( .A1(n10130), .A2(n4827), .ZN(n7665) );
  OAI21_X2 U4996 ( .B1(n7362), .B2(n4653), .A(n4651), .ZN(n7446) );
  AOI21_X2 U4997 ( .B1(n4854), .B2(n7103), .A(n4499), .ZN(n4853) );
  NAND2_X2 U4998 ( .A1(n4966), .A2(n4965), .ZN(n4560) );
  NAND2_X2 U4999 ( .A1(n5944), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5945) );
  INV_X2 U5000 ( .A(n7624), .ZN(n7148) );
  NAND2_X1 U5001 ( .A1(n6884), .A2(n6000), .ZN(n4456) );
  NAND2_X1 U5002 ( .A1(n6884), .A2(n6000), .ZN(n6581) );
  NAND2_X1 U5003 ( .A1(n7615), .A2(n10111), .ZN(n7614) );
  OAI21_X2 U5004 ( .B1(n7610), .B2(n10078), .A(n7609), .ZN(n10084) );
  NAND2_X2 U5005 ( .A1(n5070), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5096) );
  BUF_X2 U5006 ( .A(n10074), .Z(n4571) );
  XNOR2_X2 U5007 ( .A(n6026), .B(n6025), .ZN(n10074) );
  NAND2_X2 U5008 ( .A1(n6005), .A2(n6024), .ZN(n10057) );
  MUX2_X1 U5009 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8523), .S(n10264), .Z(n8469) );
  MUX2_X1 U5010 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8523), .S(n10240), .Z(n8524) );
  INV_X1 U5011 ( .A(n7933), .ZN(n4685) );
  NAND2_X1 U5012 ( .A1(n5788), .A2(n5787), .ZN(n5809) );
  AOI21_X1 U5013 ( .B1(n4812), .B2(n4497), .A(n4807), .ZN(n8407) );
  AND2_X1 U5014 ( .A1(n8016), .A2(n8018), .ZN(n7835) );
  OR2_X1 U5015 ( .A1(n7764), .A2(n10260), .ZN(n4572) );
  INV_X1 U5016 ( .A(n8088), .ZN(n10159) );
  NAND2_X2 U5017 ( .A1(n6042), .A2(n6409), .ZN(n10156) );
  NAND4_X1 U5018 ( .A1(n6053), .A2(n6052), .A3(n6051), .A4(n6050), .ZN(n8087)
         );
  NAND4_X1 U5019 ( .A1(n6066), .A2(n6065), .A3(n6064), .A4(n6063), .ZN(n8086)
         );
  NAND2_X1 U5020 ( .A1(n5781), .A2(n4455), .ZN(n5286) );
  BUF_X2 U5021 ( .A(n5781), .Z(n4458) );
  NAND4_X1 U5022 ( .A1(n5131), .A2(n5130), .A3(n5129), .A4(n5128), .ZN(n7274)
         );
  INV_X1 U5023 ( .A(n7092), .ZN(n10154) );
  INV_X2 U5024 ( .A(n5541), .ZN(n5529) );
  INV_X2 U5025 ( .A(n5541), .ZN(n5136) );
  INV_X2 U5026 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NAND2_X1 U5027 ( .A1(n9039), .A2(n4505), .ZN(n5876) );
  NOR2_X1 U5028 ( .A1(n9445), .A2(n4485), .ZN(n9446) );
  OAI21_X1 U5029 ( .B1(n6489), .B2(n6488), .A(n6487), .ZN(n6490) );
  XNOR2_X1 U5030 ( .A(n6752), .B(n6751), .ZN(n8265) );
  AND3_X1 U5031 ( .A1(n5040), .A2(n6378), .A3(n6377), .ZN(n6400) );
  NAND2_X1 U5032 ( .A1(n7873), .A2(n7872), .ZN(n8052) );
  OR2_X1 U5033 ( .A1(n6373), .A2(n6374), .ZN(n5040) );
  OAI21_X1 U5034 ( .B1(n9241), .B2(n9176), .A(n9175), .ZN(n9226) );
  AOI21_X1 U5035 ( .B1(n8270), .B2(n6797), .A(n8269), .ZN(n8467) );
  NAND2_X1 U5036 ( .A1(n4685), .A2(n4684), .ZN(n4683) );
  AOI21_X1 U5037 ( .B1(n4566), .B2(n6797), .A(n4563), .ZN(n8476) );
  AND2_X1 U5038 ( .A1(n4994), .A2(n4993), .ZN(n4992) );
  CLKBUF_X1 U5039 ( .A(n6444), .Z(n7822) );
  OR2_X1 U5040 ( .A1(n8295), .A2(n4802), .ZN(n4795) );
  OR2_X1 U5041 ( .A1(n4482), .A2(n8209), .ZN(n4974) );
  OR2_X1 U5042 ( .A1(n8188), .A2(n4976), .ZN(n4975) );
  XNOR2_X1 U5043 ( .A(n8207), .B(n8219), .ZN(n8188) );
  OR2_X1 U5044 ( .A1(n8295), .A2(n6440), .ZN(n4799) );
  AOI21_X1 U5045 ( .B1(n7824), .B2(n6583), .A(n6582), .ZN(n9440) );
  OR4_X1 U5046 ( .A1(n8296), .A2(n8316), .A3(n6788), .A4(n6480), .ZN(n6481) );
  XNOR2_X1 U5047 ( .A(n6380), .B(n6379), .ZN(n7824) );
  NAND2_X1 U5048 ( .A1(n4872), .A2(n4867), .ZN(n4866) );
  NOR2_X1 U5049 ( .A1(n8027), .A2(n8028), .ZN(n8026) );
  NAND2_X1 U5050 ( .A1(n4725), .A2(n9162), .ZN(n9301) );
  AND2_X1 U5051 ( .A1(n6312), .A2(n6311), .ZN(n8530) );
  AND2_X1 U5052 ( .A1(n4825), .A2(n4823), .ZN(n8347) );
  AOI21_X1 U5053 ( .B1(n8355), .B2(n8359), .A(n4988), .ZN(n8342) );
  OAI22_X2 U5054 ( .A1(n8366), .A2(n6783), .B1(n6782), .B2(n8356), .ZN(n8355)
         );
  OAI21_X1 U5055 ( .B1(n9369), .B2(n9507), .A(n9160), .ZN(n9334) );
  NAND2_X1 U5056 ( .A1(n4662), .A2(n4659), .ZN(n7963) );
  XNOR2_X1 U5057 ( .A(n5809), .B(n5808), .ZN(n8887) );
  AND2_X1 U5058 ( .A1(n4959), .A2(n8115), .ZN(n8118) );
  NAND2_X1 U5059 ( .A1(n5696), .A2(n5695), .ZN(n9304) );
  NAND2_X1 U5060 ( .A1(n8108), .A2(n8125), .ZN(n8115) );
  NAND2_X1 U5061 ( .A1(n5648), .A2(n5647), .ZN(n9500) );
  NAND2_X1 U5062 ( .A1(n5495), .A2(n5494), .ZN(n9524) );
  NAND2_X1 U5063 ( .A1(n4783), .A2(n4781), .ZN(n7521) );
  AND2_X1 U5064 ( .A1(n7479), .A2(n4484), .ZN(n5020) );
  INV_X1 U5065 ( .A(n6530), .ZN(n9988) );
  AND2_X1 U5066 ( .A1(n7711), .A2(n7715), .ZN(n6475) );
  AND2_X1 U5067 ( .A1(n7563), .A2(n7560), .ZN(n4650) );
  OAI22_X1 U5068 ( .A1(n7390), .A2(n6767), .B1(n7435), .B2(n6766), .ZN(n7403)
         );
  NAND2_X1 U5069 ( .A1(n5316), .A2(n5297), .ZN(n6875) );
  NAND2_X1 U5070 ( .A1(n6764), .A2(n6058), .ZN(n7199) );
  NOR2_X1 U5071 ( .A1(n7308), .A2(n7298), .ZN(n9875) );
  INV_X1 U5072 ( .A(n8081), .ZN(n7832) );
  INV_X1 U5073 ( .A(n7530), .ZN(n8084) );
  INV_X1 U5074 ( .A(n7558), .ZN(n8083) );
  NAND3_X1 U5075 ( .A1(n4778), .A2(n6031), .A3(n6033), .ZN(n8088) );
  AND4_X1 U5076 ( .A1(n6102), .A2(n6101), .A3(n6100), .A4(n6099), .ZN(n7530)
         );
  NAND4_X1 U5077 ( .A1(n6121), .A2(n6120), .A3(n6119), .A4(n6118), .ZN(n8082)
         );
  NAND4_X1 U5078 ( .A1(n6080), .A2(n6079), .A3(n6078), .A4(n6077), .ZN(n8085)
         );
  AND3_X1 U5079 ( .A1(n5215), .A2(n5214), .A3(n5213), .ZN(n9943) );
  AND4_X1 U5080 ( .A1(n6111), .A2(n6110), .A3(n6109), .A4(n6108), .ZN(n7558)
         );
  INV_X1 U5081 ( .A(n5136), .ZN(n5863) );
  AND2_X1 U5082 ( .A1(n5996), .A2(n5995), .ZN(n5997) );
  NAND4_X2 U5083 ( .A1(n5080), .A2(n5079), .A3(n5078), .A4(n5077), .ZN(n9065)
         );
  CLKBUF_X3 U5084 ( .A(n6019), .Z(n4461) );
  INV_X1 U5085 ( .A(n5947), .ZN(n5946) );
  CLKBUF_X1 U5086 ( .A(n5849), .Z(n6692) );
  NAND2_X2 U5087 ( .A1(n6884), .A2(n6857), .ZN(n5150) );
  XNOR2_X1 U5088 ( .A(n4562), .B(P1_IR_REG_25__SCAN_IN), .ZN(n5833) );
  NAND2_X2 U5089 ( .A1(n7054), .A2(n6509), .ZN(n6756) );
  XNOR2_X1 U5090 ( .A(n5083), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5849) );
  NAND2_X2 U5091 ( .A1(n5882), .A2(n6741), .ZN(n6884) );
  INV_X2 U5092 ( .A(n6755), .ZN(n8241) );
  NAND2_X1 U5093 ( .A1(n5085), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5083) );
  OR2_X1 U5094 ( .A1(n7544), .A2(n9394), .ZN(n6968) );
  AND2_X1 U5095 ( .A1(n5090), .A2(n5097), .ZN(n5834) );
  OAI21_X1 U5096 ( .B1(n5920), .B2(n5043), .A(n5941), .ZN(n7054) );
  NAND2_X1 U5097 ( .A1(n5094), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4562) );
  XNOR2_X1 U5098 ( .A(n5119), .B(n5118), .ZN(n7544) );
  NAND2_X1 U5099 ( .A1(n5097), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5099) );
  OAI21_X1 U5100 ( .B1(n5117), .B2(n5116), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5119) );
  XNOR2_X1 U5101 ( .A(n6055), .B(P2_IR_REG_4__SCAN_IN), .ZN(n7624) );
  INV_X2 U5102 ( .A(n4617), .ZN(n4457) );
  AND4_X1 U5103 ( .A1(n6249), .A2(n5912), .A3(n5911), .A4(n5910), .ZN(n5913)
         );
  AND2_X1 U5104 ( .A1(n4532), .A2(n5030), .ZN(n4793) );
  NAND2_X1 U5105 ( .A1(n4521), .A2(n5064), .ZN(n4941) );
  AND3_X1 U5106 ( .A1(n5909), .A2(n6220), .A3(n5908), .ZN(n6249) );
  AND2_X1 U5107 ( .A1(n5907), .A2(n5915), .ZN(n4792) );
  INV_X1 U5108 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6494) );
  INV_X1 U5109 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6220) );
  NOR2_X1 U5110 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5055) );
  INV_X1 U5111 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n8631) );
  NOR2_X1 U5112 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5905) );
  INV_X1 U5113 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6068) );
  NOR2_X1 U5114 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n4929) );
  NAND2_X1 U5115 ( .A1(n7033), .A2(n6757), .ZN(n6407) );
  OR2_X2 U5116 ( .A1(n7758), .A2(n4964), .ZN(n4963) );
  OAI21_X2 U5117 ( .B1(n8931), .B2(n5640), .A(n5639), .ZN(n8987) );
  XNOR2_X1 U5118 ( .A(n5113), .B(P1_IR_REG_19__SCAN_IN), .ZN(n9394) );
  NOR2_X2 U5119 ( .A1(n8187), .A2(n4960), .ZN(n8207) );
  NAND2_X1 U5120 ( .A1(n5123), .A2(n6848), .ZN(n5781) );
  CLKBUF_X1 U5121 ( .A(n6741), .Z(n4459) );
  XNOR2_X1 U5122 ( .A(n5099), .B(n5098), .ZN(n6741) );
  NAND2_X2 U5123 ( .A1(n7277), .A2(n6848), .ZN(n5541) );
  NOR2_X2 U5124 ( .A1(n8380), .A2(n5036), .ZN(n8366) );
  XNOR2_X2 U5125 ( .A(n5096), .B(n5095), .ZN(n5882) );
  NOR2_X1 U5126 ( .A1(n7825), .A2(n5946), .ZN(n6017) );
  INV_X2 U5127 ( .A(n4463), .ZN(n6048) );
  AND2_X4 U5129 ( .A1(n5946), .A2(n7825), .ZN(n6018) );
  XNOR2_X2 U5130 ( .A(n5945), .B(P2_IR_REG_30__SCAN_IN), .ZN(n7825) );
  INV_X1 U5131 ( .A(n6016), .ZN(n4463) );
  AND2_X1 U5132 ( .A1(n4630), .A2(n4625), .ZN(n6559) );
  AOI21_X1 U5133 ( .B1(n4627), .B2(n4626), .A(n9386), .ZN(n4625) );
  NAND3_X1 U5134 ( .A1(n7031), .A2(n4633), .A3(n7030), .ZN(n4632) );
  XNOR2_X1 U5135 ( .A(n7431), .B(n7165), .ZN(n4633) );
  NOR2_X1 U5136 ( .A1(n6792), .A2(n4999), .ZN(n4998) );
  INV_X1 U5137 ( .A(n5003), .ZN(n4999) );
  OR2_X1 U5138 ( .A1(n8304), .A2(n8313), .ZN(n6439) );
  OAI21_X1 U5139 ( .B1(n7170), .B2(n7169), .A(n6407), .ZN(n10150) );
  NOR2_X1 U5140 ( .A1(n4731), .A2(n4729), .ZN(n4728) );
  INV_X1 U5141 ( .A(n9177), .ZN(n4729) );
  NAND2_X1 U5142 ( .A1(n4761), .A2(n4764), .ZN(n9401) );
  INV_X1 U5143 ( .A(n4765), .ZN(n4764) );
  OAI21_X1 U5144 ( .B1(n4766), .B2(n4464), .A(n9153), .ZN(n4765) );
  AND4_X1 U5145 ( .A1(n5501), .A2(n5500), .A3(n5499), .A4(n5498), .ZN(n9422)
         );
  NAND2_X1 U5146 ( .A1(n4740), .A2(n4749), .ZN(n7692) );
  OR2_X1 U5147 ( .A1(n9988), .A2(n9995), .ZN(n4749) );
  NAND2_X1 U5148 ( .A1(n4610), .A2(n4609), .ZN(n4608) );
  NOR2_X1 U5149 ( .A1(n6706), .A2(n6536), .ZN(n4609) );
  AND2_X1 U5150 ( .A1(n6560), .A2(n4600), .ZN(n4599) );
  AOI21_X1 U5151 ( .B1(n4518), .B2(n6972), .A(n4601), .ZN(n4600) );
  NAND2_X1 U5152 ( .A1(n6568), .A2(n6972), .ZN(n4623) );
  NAND2_X1 U5153 ( .A1(n6456), .A2(n6457), .ZN(n4573) );
  INV_X1 U5154 ( .A(n8530), .ZN(n6322) );
  AND2_X1 U5155 ( .A1(n9998), .A2(n9844), .ZN(n6706) );
  INV_X1 U5156 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5065) );
  INV_X1 U5157 ( .A(n7868), .ZN(n4675) );
  NAND2_X1 U5158 ( .A1(n6003), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7071) );
  AND2_X1 U5159 ( .A1(n4802), .A2(n4490), .ZN(n4797) );
  AOI21_X1 U5160 ( .B1(n6429), .B2(n4823), .A(n6431), .ZN(n4822) );
  OR2_X1 U5161 ( .A1(n8034), .A2(n8368), .ZN(n6458) );
  AND2_X1 U5162 ( .A1(n8408), .A2(n8420), .ZN(n6779) );
  OR2_X1 U5163 ( .A1(n8015), .A2(n7908), .ZN(n6462) );
  AND2_X1 U5164 ( .A1(n5027), .A2(n4525), .ZN(n5026) );
  NAND2_X1 U5165 ( .A1(n7155), .A2(n10154), .ZN(n6042) );
  INV_X1 U5166 ( .A(n7033), .ZN(n7044) );
  INV_X1 U5167 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6025) );
  NAND2_X1 U5168 ( .A1(n4859), .A2(n4857), .ZN(n5338) );
  AOI21_X1 U5169 ( .B1(n4861), .B2(n4863), .A(n4858), .ZN(n4857) );
  NAND2_X1 U5170 ( .A1(n7347), .A2(n4861), .ZN(n4859) );
  INV_X1 U5171 ( .A(n7419), .ZN(n4858) );
  INV_X1 U5172 ( .A(n6577), .ZN(n6630) );
  OR2_X1 U5173 ( .A1(n9228), .A2(n9252), .ZN(n6644) );
  OR2_X1 U5174 ( .A1(n9478), .A2(n9469), .ZN(n9188) );
  NAND2_X1 U5175 ( .A1(n7586), .A2(n9845), .ZN(n4750) );
  INV_X1 U5176 ( .A(n6533), .ZN(n6702) );
  XNOR2_X1 U5177 ( .A(n6356), .B(n6355), .ZN(n6358) );
  NAND2_X1 U5178 ( .A1(n5765), .A2(n5764), .ZN(n5786) );
  NOR2_X1 U5179 ( .A1(n5063), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n4616) );
  NAND2_X1 U5180 ( .A1(n5117), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5084) );
  AOI21_X1 U5181 ( .B1(n4892), .B2(n4894), .A(n4537), .ZN(n4891) );
  INV_X1 U5182 ( .A(n5532), .ZN(n4892) );
  AOI21_X1 U5183 ( .B1(n4879), .B2(n4884), .A(n4519), .ZN(n4878) );
  XNOR2_X1 U5184 ( .A(n5340), .B(SI_8_), .ZN(n5342) );
  NAND2_X1 U5185 ( .A1(n5291), .A2(SI_7_), .ZN(n5315) );
  INV_X1 U5186 ( .A(n4666), .ZN(n7871) );
  NAND2_X1 U5187 ( .A1(n6400), .A2(n6851), .ZN(n6402) );
  INV_X2 U5188 ( .A(n6366), .ZN(n6346) );
  AND2_X1 U5189 ( .A1(n7135), .A2(n7139), .ZN(n4581) );
  NOR2_X1 U5190 ( .A1(n10063), .A2(n4839), .ZN(n7138) );
  NOR2_X1 U5191 ( .A1(n7129), .A2(n7139), .ZN(n7131) );
  NAND2_X1 U5192 ( .A1(n4585), .A2(n7794), .ZN(n8097) );
  AOI21_X1 U5193 ( .B1(n4998), .B2(n4996), .A(n4517), .ZN(n4995) );
  INV_X1 U5194 ( .A(n5001), .ZN(n4996) );
  AOI21_X1 U5195 ( .B1(n8307), .B2(n6439), .A(n6438), .ZN(n8295) );
  AOI21_X1 U5196 ( .B1(n8317), .B2(n6436), .A(n6435), .ZN(n8307) );
  AOI21_X1 U5197 ( .B1(n8324), .B2(n6434), .A(n6453), .ZN(n8317) );
  NAND2_X1 U5198 ( .A1(n5006), .A2(n5004), .ZN(n8380) );
  NAND2_X1 U5199 ( .A1(n5008), .A2(n5005), .ZN(n5004) );
  NAND2_X1 U5200 ( .A1(n8417), .A2(n4500), .ZN(n5006) );
  INV_X1 U5201 ( .A(n5011), .ZN(n5005) );
  NAND2_X1 U5202 ( .A1(n4808), .A2(n6425), .ZN(n4807) );
  NAND2_X1 U5203 ( .A1(n8415), .A2(n4809), .ZN(n4808) );
  AND2_X1 U5204 ( .A1(n6410), .A2(n6409), .ZN(n4777) );
  INV_X1 U5205 ( .A(n6038), .ZN(n6387) );
  INV_X1 U5206 ( .A(n6037), .ZN(n6332) );
  NAND2_X1 U5207 ( .A1(n7222), .A2(n5101), .ZN(n5102) );
  INV_X1 U5208 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5100) );
  AND2_X1 U5209 ( .A1(n6630), .A2(n6674), .ZN(n9195) );
  OR2_X1 U5210 ( .A1(n9244), .A2(n9174), .ZN(n9175) );
  NOR2_X1 U5211 ( .A1(n9463), .A2(n9455), .ZN(n9176) );
  BUF_X1 U5212 ( .A(n5145), .Z(n6584) );
  NAND2_X1 U5213 ( .A1(n9482), .A2(n9315), .ZN(n9168) );
  OR2_X1 U5214 ( .A1(n9304), .A2(n9163), .ZN(n9164) );
  OR2_X1 U5215 ( .A1(n9489), .A2(n9481), .ZN(n5038) );
  NAND2_X1 U5216 ( .A1(n4733), .A2(n4732), .ZN(n9160) );
  NOR2_X1 U5217 ( .A1(n4513), .A2(n9157), .ZN(n4732) );
  NAND2_X1 U5218 ( .A1(n7583), .A2(n4687), .ZN(n4689) );
  NOR2_X1 U5219 ( .A1(n6661), .A2(n4688), .ZN(n4687) );
  OR2_X1 U5220 ( .A1(n9524), .A2(n9422), .ZN(n6660) );
  NAND2_X1 U5221 ( .A1(n4767), .A2(n4772), .ZN(n4766) );
  INV_X1 U5222 ( .A(n4771), .ZN(n4767) );
  AOI21_X1 U5223 ( .B1(n7744), .B2(n4773), .A(n4510), .ZN(n4771) );
  NOR2_X1 U5224 ( .A1(n7509), .A2(n4747), .ZN(n4746) );
  INV_X1 U5225 ( .A(n6581), .ZN(n5619) );
  INV_X1 U5226 ( .A(n6884), .ZN(n5618) );
  INV_X1 U5227 ( .A(n5150), .ZN(n6583) );
  NAND2_X1 U5228 ( .A1(n4524), .A2(n4580), .ZN(n9860) );
  NAND2_X1 U5229 ( .A1(n4612), .A2(n6689), .ZN(n4611) );
  INV_X1 U5230 ( .A(n9001), .ZN(n4774) );
  XNOR2_X1 U5231 ( .A(n5853), .B(n5852), .ZN(n7823) );
  NAND2_X1 U5232 ( .A1(n4910), .A2(n5810), .ZN(n5853) );
  NAND2_X1 U5233 ( .A1(n5809), .A2(n5808), .ZN(n4910) );
  OAI21_X1 U5234 ( .B1(n5420), .B2(n4899), .A(n4897), .ZN(n5481) );
  INV_X1 U5235 ( .A(n4900), .ZN(n4899) );
  AOI21_X1 U5236 ( .B1(n4900), .B2(n4902), .A(n4898), .ZN(n4897) );
  INV_X1 U5237 ( .A(n5457), .ZN(n4898) );
  INV_X1 U5238 ( .A(n8079), .ZN(n8405) );
  NOR2_X1 U5239 ( .A1(n6538), .A2(n6589), .ZN(n4607) );
  NAND2_X1 U5240 ( .A1(n4605), .A2(n4503), .ZN(n4604) );
  NAND2_X1 U5241 ( .A1(n6540), .A2(n6704), .ZN(n4605) );
  INV_X1 U5242 ( .A(n6545), .ZN(n6546) );
  NOR2_X1 U5243 ( .A1(n6297), .A2(n8316), .ZN(n4575) );
  NAND2_X1 U5244 ( .A1(n6805), .A2(n4631), .ZN(n7031) );
  AND2_X1 U5245 ( .A1(n6804), .A2(n4634), .ZN(n4631) );
  NAND2_X1 U5246 ( .A1(n7456), .A2(n7552), .ZN(n7374) );
  NAND2_X1 U5247 ( .A1(n4678), .A2(n4681), .ZN(n4677) );
  INV_X1 U5248 ( .A(n8008), .ZN(n4678) );
  NOR2_X1 U5249 ( .A1(n7863), .A2(n4680), .ZN(n4679) );
  INV_X1 U5250 ( .A(n4682), .ZN(n4680) );
  INV_X1 U5251 ( .A(n7955), .ZN(n4669) );
  INV_X1 U5252 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5028) );
  NAND2_X1 U5253 ( .A1(n10074), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7074) );
  INV_X1 U5254 ( .A(n4844), .ZN(n4843) );
  AOI21_X1 U5255 ( .B1(n7143), .B2(n7608), .A(n4845), .ZN(n4844) );
  OR2_X1 U5256 ( .A1(n10108), .A2(n7603), .ZN(n4968) );
  NOR2_X1 U5257 ( .A1(n5921), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U5258 ( .A1(n4968), .A2(n4967), .ZN(n4966) );
  INV_X1 U5259 ( .A(n10128), .ZN(n4967) );
  NOR2_X1 U5260 ( .A1(n10140), .A2(n10254), .ZN(n4827) );
  OAI21_X1 U5261 ( .B1(n8100), .B2(n4832), .A(n4830), .ZN(n8146) );
  AOI21_X1 U5262 ( .B1(n8126), .B2(n4831), .A(n8129), .ZN(n4830) );
  NOR2_X1 U5263 ( .A1(n8195), .A2(n4584), .ZN(n8211) );
  NOR2_X1 U5264 ( .A1(n8190), .A2(n8517), .ZN(n4584) );
  NAND2_X1 U5265 ( .A1(n6439), .A2(n6437), .ZN(n6788) );
  AND2_X1 U5266 ( .A1(n8542), .A2(n8076), .ZN(n6435) );
  NAND2_X1 U5267 ( .A1(n7986), .A2(n8322), .ZN(n6436) );
  AND2_X1 U5268 ( .A1(n8325), .A2(n8334), .ZN(n6453) );
  OR2_X1 U5269 ( .A1(n8499), .A2(n8369), .ZN(n6457) );
  AND2_X1 U5270 ( .A1(n5013), .A2(n5012), .ZN(n5011) );
  NOR2_X1 U5271 ( .A1(n6779), .A2(n5016), .ZN(n5015) );
  INV_X1 U5272 ( .A(n6778), .ZN(n5016) );
  OR2_X1 U5273 ( .A1(n6225), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6238) );
  NOR2_X1 U5274 ( .A1(n6193), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n4555) );
  OR2_X1 U5275 ( .A1(n9632), .A2(n8453), .ZN(n6424) );
  INV_X1 U5276 ( .A(n4486), .ZN(n5019) );
  INV_X1 U5277 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5914) );
  INV_X1 U5278 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5904) );
  NOR2_X1 U5279 ( .A1(n9442), .A2(n9450), .ZN(n4949) );
  INV_X1 U5280 ( .A(n9234), .ZN(n4695) );
  AND2_X1 U5281 ( .A1(n5745), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5773) );
  INV_X1 U5282 ( .A(n9290), .ZN(n9184) );
  NOR2_X1 U5283 ( .A1(n9311), .A2(n9183), .ZN(n9286) );
  NAND2_X1 U5284 ( .A1(n9181), .A2(n9182), .ZN(n9183) );
  INV_X1 U5285 ( .A(n9309), .ZN(n9182) );
  NOR2_X1 U5286 ( .A1(n5622), .A2(n8722), .ZN(n5623) );
  NAND2_X1 U5287 ( .A1(n4951), .A2(n9422), .ZN(n4772) );
  NAND2_X1 U5288 ( .A1(n7654), .A2(n4956), .ZN(n4955) );
  INV_X1 U5289 ( .A(n4957), .ZN(n4956) );
  NOR2_X1 U5290 ( .A1(n5348), .A2(n8730), .ZN(n5396) );
  AND2_X1 U5291 ( .A1(n9972), .A2(n8926), .ZN(n7486) );
  OR2_X1 U5292 ( .A1(n5150), .A2(n6867), .ZN(n5112) );
  NOR2_X1 U5293 ( .A1(n4590), .A2(n4589), .ZN(n4591) );
  NAND2_X1 U5294 ( .A1(n6000), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4589) );
  NOR2_X1 U5295 ( .A1(n4935), .A2(n9299), .ZN(n4934) );
  INV_X1 U5296 ( .A(n4936), .ZN(n4935) );
  OAI21_X1 U5297 ( .B1(n6358), .B2(SI_29_), .A(n6357), .ZN(n6380) );
  INV_X1 U5298 ( .A(n4941), .ZN(n4939) );
  INV_X1 U5299 ( .A(n4925), .ZN(n4924) );
  AOI21_X1 U5300 ( .B1(n4925), .B2(n4923), .A(n4922), .ZN(n4921) );
  OAI21_X1 U5301 ( .B1(n5646), .B2(n5645), .A(n5644), .ZN(n5663) );
  NAND2_X1 U5302 ( .A1(n5153), .A2(SI_2_), .ZN(n5172) );
  INV_X1 U5303 ( .A(n6839), .ZN(n6851) );
  AOI21_X1 U5304 ( .B1(n7878), .B2(n4646), .A(n7922), .ZN(n4645) );
  INV_X1 U5305 ( .A(n7876), .ZN(n4646) );
  INV_X1 U5306 ( .A(n4645), .ZN(n4642) );
  NAND2_X1 U5307 ( .A1(n7833), .A2(n7832), .ZN(n8016) );
  AND2_X1 U5308 ( .A1(n5913), .A2(n4793), .ZN(n4794) );
  OAI21_X1 U5309 ( .B1(n10057), .B2(n7070), .A(n7071), .ZN(n10046) );
  NOR2_X1 U5310 ( .A1(n10046), .A2(n10241), .ZN(n10045) );
  NOR2_X1 U5311 ( .A1(n10066), .A2(n5048), .ZN(n7129) );
  OAI21_X1 U5312 ( .B1(n10120), .B2(n10252), .A(n7614), .ZN(n4829) );
  INV_X1 U5313 ( .A(n4966), .ZN(n10127) );
  INV_X1 U5314 ( .A(n4968), .ZN(n10129) );
  AND2_X1 U5315 ( .A1(n4829), .A2(n4828), .ZN(n10130) );
  INV_X1 U5316 ( .A(n10131), .ZN(n4828) );
  NAND2_X1 U5317 ( .A1(n7629), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4965) );
  NAND2_X1 U5318 ( .A1(n4572), .A2(n4488), .ZN(n4585) );
  NOR2_X1 U5319 ( .A1(n7678), .A2(n8638), .ZN(n4964) );
  INV_X1 U5320 ( .A(n7787), .ZN(n4558) );
  OR2_X1 U5321 ( .A1(n8108), .A2(n8125), .ZN(n4958) );
  NAND3_X1 U5322 ( .A1(n4958), .A2(n8115), .A3(P2_REG2_REG_13__SCAN_IN), .ZN(
        n4959) );
  NOR2_X1 U5323 ( .A1(n8178), .A2(n8177), .ZN(n8195) );
  XNOR2_X1 U5324 ( .A(n8211), .B(n8219), .ZN(n8198) );
  OAI21_X1 U5325 ( .B1(n10148), .B2(n10274), .A(n4569), .ZN(n4568) );
  INV_X1 U5326 ( .A(n8225), .ZN(n4569) );
  OR2_X1 U5327 ( .A1(n8209), .A2(n8836), .ZN(n4976) );
  AND2_X1 U5328 ( .A1(n6395), .A2(n6339), .ZN(n8268) );
  INV_X1 U5329 ( .A(n4998), .ZN(n4997) );
  NAND2_X1 U5330 ( .A1(n6442), .A2(n4805), .ZN(n4802) );
  NAND2_X1 U5331 ( .A1(n4801), .A2(n6442), .ZN(n4800) );
  INV_X1 U5332 ( .A(n4803), .ZN(n4801) );
  XNOR2_X1 U5333 ( .A(n8277), .B(n8281), .ZN(n8273) );
  NAND2_X1 U5334 ( .A1(n8299), .A2(n8303), .ZN(n6441) );
  NAND2_X1 U5335 ( .A1(n6442), .A2(n6340), .ZN(n8282) );
  NAND2_X1 U5336 ( .A1(n8291), .A2(n8437), .ZN(n4565) );
  OR2_X1 U5337 ( .A1(n6440), .A2(n6323), .ZN(n8296) );
  AND2_X1 U5338 ( .A1(n5977), .A2(n5976), .ZN(n8313) );
  NAND2_X1 U5339 ( .A1(n4553), .A2(n5938), .ZN(n5971) );
  AOI21_X1 U5340 ( .B1(n4981), .B2(n4985), .A(n4516), .ZN(n4978) );
  OR2_X1 U5341 ( .A1(n4818), .A2(n4817), .ZN(n4816) );
  NOR2_X1 U5342 ( .A1(n8349), .A2(n4987), .ZN(n4986) );
  INV_X1 U5343 ( .A(n8359), .ZN(n4987) );
  AOI21_X1 U5344 ( .B1(n4822), .B2(n4820), .A(n4819), .ZN(n4818) );
  INV_X1 U5345 ( .A(n4823), .ZN(n4820) );
  INV_X1 U5346 ( .A(n4822), .ZN(n4821) );
  NAND2_X1 U5347 ( .A1(n4815), .A2(n4826), .ZN(n4825) );
  NOR2_X1 U5348 ( .A1(n6780), .A2(n8405), .ZN(n5009) );
  NAND2_X1 U5349 ( .A1(n5014), .A2(n5011), .ZN(n5010) );
  AND2_X1 U5350 ( .A1(n6458), .A2(n8370), .ZN(n8385) );
  OR2_X1 U5351 ( .A1(n8401), .A2(n6779), .ZN(n5013) );
  NAND2_X1 U5352 ( .A1(n8417), .A2(n5015), .ZN(n5014) );
  INV_X1 U5353 ( .A(n6424), .ZN(n4809) );
  AND2_X1 U5354 ( .A1(n4813), .A2(n4811), .ZN(n4810) );
  INV_X1 U5355 ( .A(n4555), .ZN(n6208) );
  OR2_X1 U5356 ( .A1(n6460), .A2(n6423), .ZN(n4813) );
  NAND2_X1 U5357 ( .A1(n6169), .A2(n6168), .ZN(n7939) );
  NAND2_X1 U5358 ( .A1(n6462), .A2(n6461), .ZN(n7834) );
  NAND2_X1 U5359 ( .A1(n6134), .A2(n6133), .ZN(n7901) );
  NAND2_X1 U5360 ( .A1(n7714), .A2(n7562), .ZN(n5027) );
  AND2_X1 U5361 ( .A1(n6467), .A2(n4782), .ZN(n4781) );
  NAND2_X1 U5362 ( .A1(n7405), .A2(n6415), .ZN(n4783) );
  NAND2_X1 U5363 ( .A1(n6414), .A2(n6415), .ZN(n4782) );
  OAI211_X1 U5364 ( .C1(n6756), .C2(n10111), .A(n6105), .B(n6104), .ZN(n7447)
         );
  INV_X1 U5365 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5927) );
  INV_X1 U5366 ( .A(n6061), .ZN(n5928) );
  NAND2_X1 U5367 ( .A1(n7001), .A2(n6851), .ZN(n10158) );
  INV_X1 U5368 ( .A(n8435), .ZN(n10157) );
  INV_X1 U5369 ( .A(n10158), .ZN(n8437) );
  AND2_X1 U5370 ( .A1(n7042), .A2(n6851), .ZN(n8435) );
  NAND2_X1 U5371 ( .A1(n6390), .A2(n6389), .ZN(n6449) );
  NAND2_X1 U5372 ( .A1(n6334), .A2(n6333), .ZN(n6825) );
  NAND2_X1 U5373 ( .A1(n6805), .A2(n6804), .ZN(n6807) );
  NAND2_X1 U5374 ( .A1(n5918), .A2(n5922), .ZN(n5031) );
  NAND2_X1 U5375 ( .A1(n6496), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6500) );
  XNOR2_X1 U5376 ( .A(n5964), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7165) );
  OR2_X1 U5377 ( .A1(n6082), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U5378 ( .A1(n6003), .A2(n6025), .ZN(n6035) );
  NAND2_X1 U5379 ( .A1(n4522), .A2(n4473), .ZN(n6907) );
  AND2_X1 U5380 ( .A1(n4489), .A2(n5686), .ZN(n4847) );
  INV_X1 U5381 ( .A(n8949), .ZN(n4582) );
  NAND2_X1 U5382 ( .A1(n5120), .A2(n6968), .ZN(n5121) );
  NAND2_X1 U5383 ( .A1(n6739), .A2(n4587), .ZN(n6745) );
  AND2_X1 U5384 ( .A1(n6735), .A2(n4526), .ZN(n6737) );
  NAND2_X1 U5385 ( .A1(n4917), .A2(n4914), .ZN(n4596) );
  AND2_X1 U5386 ( .A1(n6590), .A2(n4594), .ZN(n4593) );
  OR4_X1 U5387 ( .A1(n6624), .A2(n9266), .A3(n9187), .A4(n9290), .ZN(n6625) );
  AND2_X1 U5388 ( .A1(n9692), .A2(n4716), .ZN(n9715) );
  NAND2_X1 U5389 ( .A1(n9695), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4716) );
  OR2_X1 U5390 ( .A1(n9715), .A2(n9714), .ZN(n4715) );
  NOR2_X1 U5391 ( .A1(n9570), .A2(n4708), .ZN(n9723) );
  AND2_X1 U5392 ( .A1(n9575), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4708) );
  AND2_X1 U5393 ( .A1(n4947), .A2(n4946), .ZN(n4945) );
  OR2_X1 U5394 ( .A1(n9227), .A2(n4946), .ZN(n4943) );
  NOR2_X1 U5395 ( .A1(n9148), .A2(n4948), .ZN(n4947) );
  INV_X1 U5396 ( .A(n4949), .ZN(n4948) );
  NAND2_X1 U5397 ( .A1(n9450), .A2(n9236), .ZN(n9192) );
  AND2_X1 U5398 ( .A1(n4691), .A2(n4690), .ZN(n9209) );
  AND2_X1 U5399 ( .A1(n4692), .A2(n9191), .ZN(n4690) );
  OR2_X1 U5400 ( .A1(n9251), .A2(n4693), .ZN(n4691) );
  NAND2_X1 U5401 ( .A1(n4695), .A2(n4694), .ZN(n4693) );
  INV_X1 U5402 ( .A(n9250), .ZN(n4694) );
  NAND2_X1 U5403 ( .A1(n4695), .A2(n9190), .ZN(n4692) );
  NAND2_X1 U5404 ( .A1(n6644), .A2(n9191), .ZN(n9234) );
  OR2_X1 U5405 ( .A1(n9251), .A2(n9250), .ZN(n4696) );
  AND4_X1 U5406 ( .A1(n5823), .A2(n5822), .A3(n5821), .A4(n5820), .ZN(n9252)
         );
  NAND2_X1 U5407 ( .A1(n5794), .A2(n5793), .ZN(n9244) );
  NAND2_X1 U5408 ( .A1(n8887), .A2(n6583), .ZN(n5794) );
  NAND2_X1 U5409 ( .A1(n4752), .A2(n4753), .ZN(n9241) );
  NOR2_X1 U5410 ( .A1(n4754), .A2(n4504), .ZN(n4753) );
  OR2_X1 U5411 ( .A1(n4937), .A2(n9478), .ZN(n9276) );
  NOR2_X1 U5412 ( .A1(n9167), .A2(n4501), .ZN(n4757) );
  AND2_X1 U5413 ( .A1(n9272), .A2(n9186), .ZN(n4705) );
  OR2_X1 U5414 ( .A1(n9286), .A2(n9185), .ZN(n4706) );
  AND2_X1 U5415 ( .A1(n4706), .A2(n9186), .ZN(n9273) );
  AND4_X1 U5416 ( .A1(n5727), .A2(n5726), .A3(n5725), .A4(n5724), .ZN(n9315)
         );
  INV_X1 U5417 ( .A(n6561), .ZN(n9319) );
  AOI21_X1 U5418 ( .B1(n4727), .B2(n4726), .A(n9161), .ZN(n9318) );
  NAND2_X1 U5419 ( .A1(n9339), .A2(n9324), .ZN(n4726) );
  INV_X1 U5420 ( .A(n9334), .ZN(n4727) );
  NAND2_X1 U5421 ( .A1(n6668), .A2(n6723), .ZN(n9340) );
  NOR2_X1 U5422 ( .A1(n4506), .A2(n4735), .ZN(n4734) );
  INV_X1 U5423 ( .A(n4737), .ZN(n4735) );
  NAND2_X1 U5424 ( .A1(n9406), .A2(n4699), .ZN(n4698) );
  NOR2_X1 U5425 ( .A1(n6665), .A2(n4700), .ZN(n4699) );
  INV_X1 U5426 ( .A(n6712), .ZN(n4700) );
  NAND2_X1 U5427 ( .A1(n4698), .A2(n4697), .ZN(n9366) );
  AND2_X1 U5428 ( .A1(n9368), .A2(n6666), .ZN(n4697) );
  NAND2_X1 U5429 ( .A1(n4738), .A2(n9376), .ZN(n4737) );
  AOI21_X1 U5430 ( .B1(n9401), .B2(n9400), .A(n9154), .ZN(n9384) );
  AND2_X1 U5431 ( .A1(n9520), .A2(n9388), .ZN(n9154) );
  AND2_X1 U5432 ( .A1(n6662), .A2(n6660), .ZN(n4686) );
  AND2_X1 U5433 ( .A1(n4773), .A2(n4772), .ZN(n4769) );
  AND2_X1 U5434 ( .A1(n6660), .A2(n6548), .ZN(n7749) );
  NAND2_X1 U5435 ( .A1(n4774), .A2(n8909), .ZN(n4773) );
  AOI21_X1 U5436 ( .B1(n7692), .B2(n7691), .A(n5044), .ZN(n7745) );
  AND2_X1 U5437 ( .A1(n6601), .A2(n6659), .ZN(n7744) );
  INV_X1 U5438 ( .A(n6539), .ZN(n7687) );
  INV_X1 U5439 ( .A(n4750), .ZN(n4741) );
  AND2_X1 U5440 ( .A1(n7687), .A2(n6602), .ZN(n9847) );
  INV_X1 U5441 ( .A(n4745), .ZN(n4744) );
  OAI22_X1 U5442 ( .A1(n7509), .A2(n4751), .B1(n9972), .B2(n9979), .ZN(n4745)
         );
  NAND2_X1 U5443 ( .A1(n7458), .A2(n7457), .ZN(n7485) );
  NAND2_X1 U5444 ( .A1(n7316), .A2(n4614), .ZN(n4613) );
  NAND2_X1 U5445 ( .A1(n4588), .A2(n4493), .ZN(n6525) );
  NAND2_X1 U5446 ( .A1(n7306), .A2(n7305), .ZN(n7304) );
  INV_X1 U5447 ( .A(n9881), .ZN(n9864) );
  OR2_X1 U5448 ( .A1(n7019), .A2(n5150), .ZN(n5495) );
  AND2_X1 U5449 ( .A1(n9066), .A2(n7279), .ZN(n9996) );
  AND2_X1 U5450 ( .A1(n4940), .A2(n5098), .ZN(n4938) );
  XNOR2_X1 U5451 ( .A(n6358), .B(SI_29_), .ZN(n7812) );
  NAND2_X1 U5452 ( .A1(n4909), .A2(n4907), .ZN(n6326) );
  AOI21_X1 U5453 ( .B1(n4911), .B2(n4913), .A(n4908), .ZN(n4907) );
  NAND2_X1 U5454 ( .A1(n5809), .A2(n4911), .ZN(n4909) );
  INV_X1 U5455 ( .A(n5854), .ZN(n4908) );
  XNOR2_X1 U5456 ( .A(n5786), .B(n5785), .ZN(n7755) );
  XNOR2_X1 U5457 ( .A(n5763), .B(n5762), .ZN(n7723) );
  AND2_X1 U5458 ( .A1(n5737), .A2(n5718), .ZN(n5735) );
  OR2_X1 U5459 ( .A1(n5084), .A2(n8628), .ZN(n5086) );
  INV_X1 U5460 ( .A(n9394), .ZN(n9294) );
  OAI21_X1 U5461 ( .B1(n5533), .B2(n4893), .A(n4891), .ZN(n5591) );
  NAND2_X1 U5462 ( .A1(n5511), .A2(n5510), .ZN(n5533) );
  AND2_X1 U5463 ( .A1(n5480), .A2(n5456), .ZN(n5457) );
  AOI21_X1 U5464 ( .B1(n5419), .B2(n4903), .A(n4901), .ZN(n4900) );
  INV_X1 U5465 ( .A(n5451), .ZN(n4901) );
  NAND2_X1 U5466 ( .A1(n5389), .A2(n5371), .ZN(n5420) );
  OR2_X1 U5467 ( .A1(n5420), .A2(n5419), .ZN(n4904) );
  NOR2_X1 U5468 ( .A1(n5364), .A2(SI_9_), .ZN(n5365) );
  AND2_X1 U5469 ( .A1(n5371), .A2(n5370), .ZN(n5387) );
  OAI21_X1 U5470 ( .B1(n5290), .B2(n4884), .A(n4881), .ZN(n5343) );
  AND2_X1 U5471 ( .A1(n5315), .A2(n5294), .ZN(n5295) );
  AND2_X1 U5472 ( .A1(n5289), .A2(n5278), .ZN(n5279) );
  AND4_X1 U5473 ( .A1(n6213), .A2(n6212), .A3(n6211), .A4(n6210), .ZN(n8404)
         );
  AND4_X1 U5474 ( .A1(n6159), .A2(n6158), .A3(n6157), .A4(n6156), .ZN(n7908)
         );
  AND4_X1 U5475 ( .A1(n6259), .A2(n6258), .A3(n6257), .A4(n6256), .ZN(n8368)
         );
  INV_X1 U5476 ( .A(n4660), .ZN(n4659) );
  OAI21_X1 U5477 ( .B1(n4664), .B2(n4661), .A(n7849), .ZN(n4660) );
  NAND2_X1 U5478 ( .A1(n6224), .A2(n6223), .ZN(n8408) );
  INV_X1 U5479 ( .A(n8542), .ZN(n7986) );
  AND4_X1 U5480 ( .A1(n6276), .A2(n6275), .A3(n6274), .A4(n6273), .ZN(n8383)
         );
  NAND2_X1 U5481 ( .A1(n6180), .A2(n6179), .ZN(n9636) );
  XOR2_X1 U5482 ( .A(n8344), .B(n7862), .Z(n8008) );
  INV_X1 U5483 ( .A(n8080), .ZN(n8454) );
  OR2_X1 U5484 ( .A1(n7854), .A2(n8405), .ZN(n5035) );
  AND2_X1 U5485 ( .A1(n6321), .A2(n6320), .ZN(n8267) );
  AND4_X1 U5486 ( .A1(n6230), .A2(n6229), .A3(n6228), .A4(n6227), .ZN(n8065)
         );
  OAI211_X1 U5487 ( .C1(n6349), .C2(n5959), .A(n5958), .B(n5957), .ZN(n8077)
         );
  INV_X1 U5488 ( .A(n8383), .ZN(n8356) );
  INV_X1 U5489 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10039) );
  NAND2_X1 U5490 ( .A1(n10034), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n10041) );
  XNOR2_X1 U5491 ( .A(n4560), .B(n7618), .ZN(n7605) );
  NOR2_X1 U5492 ( .A1(n7605), .A2(n7606), .ZN(n7661) );
  INV_X1 U5493 ( .A(n10139), .ZN(n10112) );
  XNOR2_X1 U5494 ( .A(n4963), .B(n7759), .ZN(n7760) );
  NOR2_X1 U5495 ( .A1(n7760), .A2(n7761), .ZN(n7784) );
  INV_X1 U5496 ( .A(n8166), .ZN(n4961) );
  OAI21_X1 U5497 ( .B1(n6867), .B2(n6857), .A(n4476), .ZN(n4787) );
  NAND2_X1 U5498 ( .A1(n5039), .A2(n4789), .ZN(n4788) );
  NOR2_X1 U5499 ( .A1(n4790), .A2(n10262), .ZN(n4789) );
  INV_X1 U5500 ( .A(n6799), .ZN(n4790) );
  AND4_X1 U5501 ( .A1(n5269), .A2(n5268), .A3(n5267), .A4(n5266), .ZN(n7424)
         );
  AND4_X1 U5502 ( .A1(n5331), .A2(n5330), .A3(n5329), .A4(n5328), .ZN(n7647)
         );
  NAND2_X1 U5503 ( .A1(n4860), .A2(n4864), .ZN(n7420) );
  NAND2_X1 U5504 ( .A1(n7347), .A2(n4865), .ZN(n4860) );
  NAND2_X1 U5505 ( .A1(n5817), .A2(n5816), .ZN(n9228) );
  NAND2_X1 U5506 ( .A1(n7823), .A2(n6583), .ZN(n5817) );
  NAND2_X1 U5507 ( .A1(n5395), .A2(n5394), .ZN(n9980) );
  NAND2_X1 U5508 ( .A1(n5261), .A2(n5260), .ZN(n7320) );
  NAND2_X1 U5509 ( .A1(n5463), .A2(n5462), .ZN(n9001) );
  OR2_X1 U5510 ( .A1(n6984), .A2(n5150), .ZN(n5463) );
  NAND2_X1 U5511 ( .A1(n5621), .A2(n5620), .ZN(n9514) );
  AND4_X1 U5512 ( .A1(n5525), .A2(n5524), .A3(n5523), .A4(n5522), .ZN(n9421)
         );
  NAND2_X1 U5513 ( .A1(n9215), .A2(n4730), .ZN(n9179) );
  NAND2_X1 U5514 ( .A1(n9450), .A2(n9198), .ZN(n4730) );
  AND4_X1 U5515 ( .A1(n5799), .A2(n5798), .A3(n5797), .A4(n5796), .ZN(n9455)
         );
  AND4_X1 U5516 ( .A1(n5778), .A2(n5777), .A3(n5776), .A4(n5775), .ZN(n9462)
         );
  AND2_X1 U5517 ( .A1(n5704), .A2(n5703), .ZN(n9481) );
  NAND2_X1 U5518 ( .A1(n5434), .A2(n5433), .ZN(n9998) );
  OR2_X1 U5519 ( .A1(n6905), .A2(n5150), .ZN(n5434) );
  NAND2_X1 U5520 ( .A1(n5067), .A2(n5066), .ZN(n9551) );
  NOR2_X1 U5521 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n5066) );
  INV_X1 U5522 ( .A(n5070), .ZN(n5067) );
  OAI21_X1 U5523 ( .B1(n7377), .B2(n7375), .A(n6687), .ZN(n6528) );
  NAND2_X1 U5524 ( .A1(n4606), .A2(n4602), .ZN(n6545) );
  NAND2_X1 U5525 ( .A1(n4604), .A2(n4603), .ZN(n4602) );
  NOR2_X1 U5526 ( .A1(n6706), .A2(n6972), .ZN(n4603) );
  NAND2_X1 U5527 ( .A1(n4629), .A2(n4628), .ZN(n4627) );
  NOR2_X1 U5528 ( .A1(n6713), .A2(n6550), .ZN(n4628) );
  NAND2_X1 U5529 ( .A1(n6551), .A2(n7749), .ZN(n4629) );
  AOI21_X1 U5530 ( .B1(n6599), .B2(n6552), .A(n6972), .ZN(n4626) );
  NOR2_X1 U5531 ( .A1(n6555), .A2(n6972), .ZN(n4601) );
  OAI21_X1 U5532 ( .B1(n6559), .B2(n6717), .A(n6558), .ZN(n6560) );
  NAND2_X1 U5533 ( .A1(n4598), .A2(n6563), .ZN(n4597) );
  NAND2_X1 U5534 ( .A1(n4621), .A2(n4474), .ZN(n4620) );
  NOR2_X1 U5535 ( .A1(n4885), .A2(n4619), .ZN(n4618) );
  NOR2_X1 U5536 ( .A1(n6647), .A2(n6972), .ZN(n4619) );
  NAND2_X1 U5537 ( .A1(n6522), .A2(n6589), .ZN(n4886) );
  NAND2_X1 U5538 ( .A1(n9192), .A2(n9191), .ZN(n6520) );
  AND2_X1 U5539 ( .A1(n7431), .A2(n8247), .ZN(n6821) );
  INV_X1 U5540 ( .A(n4864), .ZN(n4863) );
  AND2_X1 U5541 ( .A1(n4919), .A2(n4918), .ZN(n6588) );
  INV_X1 U5542 ( .A(n6579), .ZN(n4918) );
  AND2_X1 U5543 ( .A1(n9405), .A2(n9388), .ZN(n6544) );
  INV_X1 U5544 ( .A(n6884), .ZN(n4590) );
  NAND2_X1 U5545 ( .A1(n6331), .A2(n6330), .ZN(n6356) );
  NAND2_X1 U5546 ( .A1(n6326), .A2(n6325), .ZN(n6331) );
  INV_X1 U5547 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5064) );
  INV_X1 U5548 ( .A(n4927), .ZN(n4923) );
  INV_X1 U5549 ( .A(n5735), .ZN(n4922) );
  INV_X1 U5550 ( .A(n5342), .ZN(n4880) );
  AOI21_X1 U5551 ( .B1(n4650), .B2(n4648), .A(n4498), .ZN(n4647) );
  INV_X1 U5552 ( .A(n4650), .ZN(n4649) );
  NAND2_X1 U5553 ( .A1(n7955), .A2(n4684), .ZN(n4670) );
  INV_X1 U5554 ( .A(n6372), .ZN(n6378) );
  OR2_X1 U5555 ( .A1(n6825), .A2(n8268), .ZN(n6443) );
  NAND2_X1 U5556 ( .A1(n6003), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7050) );
  AND2_X1 U5557 ( .A1(n7074), .A2(n7139), .ZN(n4835) );
  INV_X1 U5558 ( .A(n10063), .ZN(n4836) );
  NAND2_X1 U5559 ( .A1(n4839), .A2(n4838), .ZN(n4837) );
  AND4_X1 U5560 ( .A1(n4834), .A2(n4837), .A3(n4833), .A4(
        P2_REG1_REG_3__SCAN_IN), .ZN(n7140) );
  NAND2_X1 U5561 ( .A1(n8098), .A2(n8097), .ZN(n8124) );
  NAND2_X1 U5562 ( .A1(n8125), .A2(n8124), .ZN(n8126) );
  NAND2_X1 U5563 ( .A1(n4557), .A2(n4541), .ZN(n8156) );
  NOR2_X1 U5564 ( .A1(n5982), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n4553) );
  AOI21_X1 U5565 ( .B1(n4984), .B2(n4983), .A(n4982), .ZN(n4981) );
  INV_X1 U5566 ( .A(n4986), .ZN(n4983) );
  NOR2_X1 U5567 ( .A1(n6279), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n4556) );
  NOR2_X1 U5568 ( .A1(n8385), .A2(n5009), .ZN(n5008) );
  NAND2_X1 U5569 ( .A1(n5936), .A2(n5935), .ZN(n6255) );
  NOR2_X1 U5570 ( .A1(n6154), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n4554) );
  NAND2_X1 U5571 ( .A1(n7573), .A2(n6475), .ZN(n4785) );
  NAND2_X1 U5572 ( .A1(n5921), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U5573 ( .A1(n8277), .A2(n8074), .ZN(n4993) );
  OR2_X1 U5574 ( .A1(n6837), .A2(n6836), .ZN(n7012) );
  INV_X1 U5575 ( .A(n6821), .ZN(n7032) );
  NAND2_X1 U5576 ( .A1(n4794), .A2(n4791), .ZN(n6493) );
  INV_X1 U5577 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5909) );
  INV_X1 U5578 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5908) );
  OR2_X1 U5579 ( .A1(n6166), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n6177) );
  INV_X1 U5580 ( .A(n8970), .ZN(n4869) );
  NAND2_X1 U5581 ( .A1(n5849), .A2(n7433), .ZN(n5114) );
  NAND2_X1 U5582 ( .A1(n9440), .A2(n6972), .ZN(n4594) );
  NAND2_X1 U5583 ( .A1(n6588), .A2(n9440), .ZN(n4917) );
  NOR2_X1 U5584 ( .A1(n6738), .A2(n4915), .ZN(n4914) );
  OAI21_X1 U5585 ( .B1(n9440), .B2(n6972), .A(n4916), .ZN(n4915) );
  NAND2_X1 U5586 ( .A1(n9140), .A2(n9196), .ZN(n4916) );
  NAND2_X1 U5587 ( .A1(n6588), .A2(n9148), .ZN(n4595) );
  NOR2_X1 U5588 ( .A1(n4467), .A2(n4755), .ZN(n4754) );
  AND2_X1 U5589 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(n5722), .ZN(n5745) );
  NOR2_X1 U5590 ( .A1(n6727), .A2(n6726), .ZN(n4701) );
  NOR2_X1 U5591 ( .A1(n9304), .A2(n9497), .ZN(n4936) );
  AND2_X1 U5592 ( .A1(n5649), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5671) );
  AND2_X1 U5593 ( .A1(n5623), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5649) );
  OR2_X1 U5594 ( .A1(n5573), .A2(n5572), .ZN(n5622) );
  NOR2_X1 U5595 ( .A1(n4763), .A2(n4464), .ZN(n4762) );
  INV_X1 U5596 ( .A(n4769), .ZN(n4763) );
  INV_X1 U5597 ( .A(n6544), .ZN(n6599) );
  OR2_X1 U5598 ( .A1(n5465), .A2(n5464), .ZN(n5497) );
  OR2_X1 U5599 ( .A1(n5326), .A2(n5325), .ZN(n5348) );
  OR2_X1 U5600 ( .A1(n7470), .A2(n7456), .ZN(n4957) );
  INV_X1 U5601 ( .A(n9899), .ZN(n4932) );
  INV_X1 U5602 ( .A(n5114), .ZN(n7277) );
  INV_X1 U5603 ( .A(n4912), .ZN(n4911) );
  OAI21_X1 U5604 ( .B1(n5808), .B2(n4913), .A(n5852), .ZN(n4912) );
  INV_X1 U5605 ( .A(n5810), .ZN(n4913) );
  NAND2_X1 U5606 ( .A1(n5786), .A2(n5785), .ZN(n5788) );
  INV_X1 U5607 ( .A(n5590), .ZN(n4890) );
  INV_X1 U5608 ( .A(n5516), .ZN(n4895) );
  AOI21_X1 U5609 ( .B1(n5295), .B2(n4883), .A(n4882), .ZN(n4881) );
  INV_X1 U5610 ( .A(n5315), .ZN(n4882) );
  INV_X1 U5611 ( .A(n5289), .ZN(n4883) );
  NAND2_X1 U5612 ( .A1(n6000), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4574) );
  NAND2_X1 U5613 ( .A1(n6314), .A2(n6313), .ZN(n6344) );
  INV_X1 U5614 ( .A(n6315), .ZN(n6314) );
  NOR2_X1 U5615 ( .A1(n6255), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U5616 ( .A1(n4556), .A2(n8649), .ZN(n5991) );
  NAND2_X1 U5617 ( .A1(n8017), .A2(n7838), .ZN(n7940) );
  INV_X1 U5618 ( .A(n4487), .ZN(n4674) );
  AOI21_X1 U5619 ( .B1(n4487), .B2(n4673), .A(n4672), .ZN(n4671) );
  INV_X1 U5620 ( .A(n4679), .ZN(n4673) );
  INV_X1 U5621 ( .A(n7867), .ZN(n4672) );
  INV_X1 U5622 ( .A(n7886), .ZN(n4661) );
  INV_X1 U5623 ( .A(n4664), .ZN(n4663) );
  INV_X1 U5624 ( .A(n7864), .ZN(n7979) );
  NAND2_X1 U5625 ( .A1(n4683), .A2(n4679), .ZN(n4676) );
  NAND2_X1 U5626 ( .A1(n5932), .A2(n5931), .ZN(n6135) );
  INV_X1 U5627 ( .A(n6116), .ZN(n5932) );
  NAND2_X1 U5628 ( .A1(n7861), .A2(n8333), .ZN(n4682) );
  OR2_X1 U5629 ( .A1(n6135), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6154) );
  OR2_X1 U5630 ( .A1(n7969), .A2(n8079), .ZN(n7853) );
  NAND2_X1 U5631 ( .A1(n8060), .A2(n4665), .ZN(n4664) );
  INV_X1 U5632 ( .A(n5049), .ZN(n4665) );
  NAND2_X1 U5633 ( .A1(n4555), .A2(n5934), .ZN(n6225) );
  AND2_X1 U5634 ( .A1(n6395), .A2(n6394), .ZN(n7814) );
  NOR2_X1 U5635 ( .A1(n10048), .A2(n10047), .ZN(n10051) );
  OR2_X1 U5636 ( .A1(n10045), .A2(n7072), .ZN(n10062) );
  NOR2_X1 U5637 ( .A1(n10067), .A2(n10068), .ZN(n10066) );
  NOR2_X1 U5638 ( .A1(n7066), .A2(n7067), .ZN(n7134) );
  OR2_X1 U5639 ( .A1(n7052), .A2(n8744), .ZN(n4972) );
  OAI21_X1 U5640 ( .B1(n7624), .B2(n7623), .A(n7622), .ZN(n10081) );
  NOR2_X1 U5641 ( .A1(n10075), .A2(n7598), .ZN(n10095) );
  NOR2_X1 U5642 ( .A1(n7612), .A2(n7611), .ZN(n10092) );
  AOI22_X1 U5643 ( .A1(n10081), .A2(n10082), .B1(n7625), .B2(n10078), .ZN(
        n10103) );
  NOR2_X1 U5644 ( .A1(n10109), .A2(n10110), .ZN(n10108) );
  INV_X1 U5645 ( .A(n5917), .ZN(n5920) );
  NOR2_X1 U5646 ( .A1(n7632), .A2(n7633), .ZN(n7674) );
  NOR2_X1 U5647 ( .A1(n7667), .A2(n7668), .ZN(n7670) );
  NOR2_X1 U5648 ( .A1(n7770), .A2(n7771), .ZN(n7801) );
  XNOR2_X1 U5649 ( .A(n8124), .B(n8099), .ZN(n8100) );
  NAND2_X1 U5650 ( .A1(n8100), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8127) );
  OAI21_X1 U5651 ( .B1(n8156), .B2(n8174), .A(n8163), .ZN(n8157) );
  AND2_X1 U5652 ( .A1(n8176), .A2(n8175), .ZN(n8178) );
  NOR2_X1 U5653 ( .A1(n8190), .A2(n8843), .ZN(n4960) );
  NOR2_X1 U5654 ( .A1(n8198), .A2(n8197), .ZN(n8212) );
  NAND2_X1 U5655 ( .A1(n4842), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4841) );
  INV_X1 U5656 ( .A(n8214), .ZN(n4842) );
  NAND2_X1 U5657 ( .A1(n4798), .A2(n4796), .ZN(n6752) );
  AOI21_X1 U5658 ( .B1(n4800), .B2(n4797), .A(n4520), .ZN(n4796) );
  NOR2_X1 U5659 ( .A1(n8282), .A2(n4804), .ZN(n4803) );
  NOR2_X1 U5660 ( .A1(n6440), .A2(n6441), .ZN(n4804) );
  NAND2_X1 U5661 ( .A1(n8299), .A2(n8075), .ZN(n5003) );
  NOR2_X1 U5662 ( .A1(n6791), .A2(n5002), .ZN(n5001) );
  INV_X1 U5663 ( .A(n6789), .ZN(n5002) );
  INV_X1 U5664 ( .A(n6788), .ZN(n8306) );
  OR2_X1 U5665 ( .A1(n6435), .A2(n5978), .ZN(n8316) );
  INV_X1 U5666 ( .A(n4553), .ZN(n5956) );
  NOR2_X1 U5667 ( .A1(n6430), .A2(n4824), .ZN(n4823) );
  INV_X1 U5668 ( .A(n6428), .ZN(n4824) );
  INV_X1 U5669 ( .A(n4556), .ZN(n6281) );
  OAI22_X1 U5670 ( .A1(n8407), .A2(n8401), .B1(n8065), .B2(n8408), .ZN(n8397)
         );
  NAND2_X1 U5671 ( .A1(n5933), .A2(n8818), .ZN(n6193) );
  INV_X1 U5672 ( .A(n6181), .ZN(n5933) );
  AND4_X1 U5673 ( .A1(n6198), .A2(n6197), .A3(n6196), .A4(n6195), .ZN(n8453)
         );
  NAND2_X1 U5674 ( .A1(n4554), .A2(n7789), .ZN(n6181) );
  INV_X1 U5675 ( .A(n4554), .ZN(n6170) );
  AOI21_X1 U5676 ( .B1(n4469), .B2(n5026), .A(n5025), .ZN(n5024) );
  NOR2_X1 U5677 ( .A1(n7719), .A2(n7832), .ZN(n5025) );
  AOI21_X1 U5678 ( .B1(n5020), .B2(n5019), .A(n4509), .ZN(n5018) );
  NAND2_X1 U5679 ( .A1(n5020), .A2(n7403), .ZN(n5017) );
  INV_X1 U5680 ( .A(n6097), .ZN(n5930) );
  OR2_X1 U5681 ( .A1(n6106), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6116) );
  NAND2_X1 U5682 ( .A1(n5022), .A2(n4486), .ZN(n5021) );
  OR2_X1 U5683 ( .A1(n6075), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6097) );
  INV_X1 U5684 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5926) );
  NAND2_X1 U5685 ( .A1(n6408), .A2(n10150), .ZN(n4779) );
  AOI21_X1 U5686 ( .B1(n7824), .B2(n6387), .A(n6362), .ZN(n6444) );
  INV_X1 U5687 ( .A(n5034), .ZN(n5033) );
  NAND2_X1 U5688 ( .A1(n5987), .A2(n5986), .ZN(n7931) );
  AND2_X1 U5689 ( .A1(n10163), .A2(n10202), .ZN(n10227) );
  OR2_X1 U5690 ( .A1(n7405), .A2(n6414), .ZN(n4780) );
  INV_X1 U5691 ( .A(n10225), .ZN(n10180) );
  OR2_X1 U5692 ( .A1(n6839), .A2(n7032), .ZN(n7183) );
  NAND2_X1 U5693 ( .A1(n7542), .A2(n6488), .ZN(n10225) );
  INV_X1 U5694 ( .A(n10227), .ZN(n10234) );
  AND2_X1 U5695 ( .A1(n7004), .A2(n7015), .ZN(n7164) );
  XNOR2_X1 U5696 ( .A(n6506), .B(P2_IR_REG_26__SCAN_IN), .ZN(n6804) );
  NAND2_X1 U5697 ( .A1(n6505), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6506) );
  CLKBUF_X1 U5698 ( .A(n6503), .Z(n6504) );
  AND2_X1 U5699 ( .A1(n5907), .A2(n5914), .ZN(n4657) );
  AND2_X1 U5700 ( .A1(n5913), .A2(n5030), .ZN(n5029) );
  OR2_X1 U5701 ( .A1(n6003), .A2(n8876), .ZN(n6026) );
  NAND2_X1 U5702 ( .A1(n7344), .A2(n7345), .ZN(n4864) );
  AND2_X1 U5703 ( .A1(n5807), .A2(n5806), .ZN(n8892) );
  NAND2_X1 U5704 ( .A1(n5133), .A2(n5286), .ZN(n5134) );
  NAND2_X1 U5705 ( .A1(n5509), .A2(n4873), .ZN(n4872) );
  INV_X1 U5706 ( .A(n5553), .ZN(n4873) );
  CLKBUF_X1 U5707 ( .A(n8921), .Z(n9015) );
  NAND2_X1 U5708 ( .A1(n5286), .A2(n7283), .ZN(n5163) );
  XNOR2_X1 U5709 ( .A(n4561), .B(n5866), .ZN(n5142) );
  NOR2_X1 U5710 ( .A1(n5264), .A2(n5263), .ZN(n5300) );
  NAND2_X1 U5711 ( .A1(n8903), .A2(n5509), .ZN(n8958) );
  AND2_X1 U5712 ( .A1(n6675), .A2(n6674), .ZN(n6735) );
  AND2_X1 U5713 ( .A1(n9596), .A2(n9597), .ZN(n9594) );
  AND2_X1 U5714 ( .A1(n4715), .A2(n4714), .ZN(n9580) );
  NAND2_X1 U5715 ( .A1(n9718), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4714) );
  NOR2_X1 U5716 ( .A1(n9579), .A2(n4711), .ZN(n9609) );
  AND2_X1 U5717 ( .A1(n6947), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4711) );
  NOR2_X1 U5718 ( .A1(n9609), .A2(n9610), .ZN(n9608) );
  NOR2_X1 U5719 ( .A1(n9723), .A2(n9724), .ZN(n9722) );
  NOR2_X1 U5720 ( .A1(n4709), .A2(n9722), .ZN(n9739) );
  AND2_X1 U5721 ( .A1(n9124), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4709) );
  NAND2_X1 U5722 ( .A1(n9739), .A2(n9740), .ZN(n9738) );
  NOR2_X1 U5723 ( .A1(n9754), .A2(n4713), .ZN(n9770) );
  AND2_X1 U5724 ( .A1(n9753), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4713) );
  NOR2_X1 U5725 ( .A1(n9770), .A2(n9771), .ZN(n9769) );
  NOR2_X1 U5726 ( .A1(n9769), .A2(n4712), .ZN(n9127) );
  AND2_X1 U5727 ( .A1(n9126), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4712) );
  AOI21_X1 U5728 ( .B1(n4705), .B2(n9185), .A(n4703), .ZN(n4702) );
  INV_X1 U5729 ( .A(n9188), .ZN(n4703) );
  NAND2_X1 U5730 ( .A1(n9335), .A2(n4936), .ZN(n9302) );
  NAND2_X1 U5731 ( .A1(n9335), .A2(n9331), .ZN(n9326) );
  NAND2_X1 U5732 ( .A1(n9331), .A2(n9488), .ZN(n9162) );
  NAND2_X1 U5733 ( .A1(n9318), .A2(n5046), .ZN(n4725) );
  NOR2_X1 U5734 ( .A1(n5497), .A2(n5496), .ZN(n5542) );
  NAND2_X1 U5735 ( .A1(n7694), .A2(n4468), .ZN(n9427) );
  NAND2_X1 U5736 ( .A1(n7694), .A2(n4774), .ZN(n7747) );
  AND2_X1 U5737 ( .A1(n5377), .A2(n5376), .ZN(n6530) );
  NAND2_X1 U5738 ( .A1(n4953), .A2(n4475), .ZN(n9856) );
  INV_X1 U5739 ( .A(n4955), .ZN(n4954) );
  NOR2_X1 U5740 ( .A1(n7382), .A2(n7456), .ZN(n7467) );
  OR2_X1 U5741 ( .A1(n7375), .A2(n7461), .ZN(n7460) );
  NAND2_X1 U5742 ( .A1(n6524), .A2(n6523), .ZN(n7278) );
  NOR2_X1 U5743 ( .A1(n7274), .A2(n9901), .ZN(n9880) );
  INV_X1 U5744 ( .A(n6969), .ZN(n6740) );
  AND2_X1 U5745 ( .A1(n9442), .A2(n9997), .ZN(n9443) );
  NAND2_X1 U5746 ( .A1(n9406), .A2(n6712), .ZN(n9387) );
  INV_X1 U5747 ( .A(n7275), .ZN(n9920) );
  XNOR2_X1 U5748 ( .A(n6386), .B(n6385), .ZN(n8875) );
  NAND2_X1 U5749 ( .A1(n6382), .A2(n6381), .ZN(n6386) );
  XNOR2_X1 U5750 ( .A(n5072), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5075) );
  INV_X1 U5751 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5098) );
  NAND2_X1 U5752 ( .A1(n4457), .A2(n4939), .ZN(n5088) );
  AND2_X1 U5753 ( .A1(n5094), .A2(n5093), .ZN(n5830) );
  NOR2_X1 U5754 ( .A1(n5712), .A2(n4928), .ZN(n4927) );
  INV_X1 U5755 ( .A(n5691), .ZN(n4928) );
  AOI21_X1 U5756 ( .B1(n4927), .B2(n4536), .A(n4926), .ZN(n4925) );
  INV_X1 U5757 ( .A(n5711), .ZN(n4926) );
  NOR2_X1 U5758 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n4874) );
  NAND2_X1 U5759 ( .A1(n5535), .A2(n5516), .ZN(n5563) );
  AND2_X1 U5760 ( .A1(n5516), .A2(n5515), .ZN(n5532) );
  AND2_X1 U5761 ( .A1(n5510), .A2(n5485), .ZN(n5486) );
  AND2_X1 U5762 ( .A1(n5273), .A2(n5235), .ZN(n5236) );
  CLKBUF_X1 U5763 ( .A(n5241), .Z(n5242) );
  NOR2_X2 U5764 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5159) );
  AND2_X1 U5765 ( .A1(n5230), .A2(n5205), .ZN(n5206) );
  INV_X1 U5766 ( .A(SI_4_), .ZN(n5203) );
  AND2_X1 U5767 ( .A1(n5200), .A2(n5177), .ZN(n5178) );
  AND2_X1 U5768 ( .A1(n4552), .A2(n5172), .ZN(n5156) );
  XNOR2_X1 U5769 ( .A(n4717), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6929) );
  NAND2_X1 U5770 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4717) );
  AOI21_X1 U5771 ( .B1(n4654), .B2(n4652), .A(n4514), .ZN(n4651) );
  INV_X1 U5772 ( .A(n4654), .ZN(n4653) );
  NAND2_X1 U5773 ( .A1(n7879), .A2(n7878), .ZN(n7923) );
  NOR2_X1 U5774 ( .A1(n7884), .A2(n7886), .ZN(n7885) );
  NAND2_X1 U5775 ( .A1(n5954), .A2(n5953), .ZN(n8325) );
  NOR2_X1 U5776 ( .A1(n4642), .A2(n7924), .ZN(n4640) );
  OAI22_X1 U5777 ( .A1(n4643), .A2(n4642), .B1(n7924), .B2(n4645), .ZN(n4641)
         );
  NOR2_X1 U5778 ( .A1(n7924), .A2(n7878), .ZN(n4643) );
  NAND2_X1 U5779 ( .A1(n7878), .A2(n7924), .ZN(n4644) );
  NAND2_X1 U5780 ( .A1(n7533), .A2(n7534), .ZN(n7561) );
  NAND2_X1 U5781 ( .A1(n7036), .A2(n7093), .ZN(n7038) );
  AND4_X1 U5782 ( .A1(n6285), .A2(n6284), .A3(n6283), .A4(n6282), .ZN(n8369)
         );
  NAND2_X1 U5783 ( .A1(n7940), .A2(n7941), .ZN(n7945) );
  AND2_X1 U5784 ( .A1(n5952), .A2(n5951), .ZN(n8322) );
  NAND2_X1 U5785 ( .A1(n4667), .A2(n4671), .ZN(n7954) );
  NAND2_X1 U5786 ( .A1(n4685), .A2(n4668), .ZN(n4667) );
  NOR2_X1 U5787 ( .A1(n4674), .A2(n7932), .ZN(n4668) );
  NOR2_X1 U5788 ( .A1(n7961), .A2(n8420), .ZN(n7850) );
  NAND2_X1 U5789 ( .A1(n7256), .A2(n7255), .ZN(n7265) );
  NAND2_X1 U5790 ( .A1(n6278), .A2(n6277), .ZN(n8499) );
  AND2_X1 U5791 ( .A1(n7117), .A2(n7642), .ZN(n8003) );
  NAND2_X1 U5792 ( .A1(n4635), .A2(n4636), .ZN(n7999) );
  INV_X1 U5793 ( .A(n4637), .ZN(n4636) );
  OAI21_X1 U5794 ( .B1(n7838), .B2(n4638), .A(n7942), .ZN(n4637) );
  NAND2_X1 U5795 ( .A1(n4683), .A2(n4682), .ZN(n8007) );
  NAND2_X1 U5796 ( .A1(n5980), .A2(n5979), .ZN(n8012) );
  NAND2_X1 U5797 ( .A1(n7903), .A2(n7835), .ZN(n8017) );
  NAND2_X1 U5798 ( .A1(n6254), .A2(n6253), .ZN(n8034) );
  OR2_X1 U5799 ( .A1(n7252), .A2(n6038), .ZN(n6254) );
  AND2_X1 U5800 ( .A1(n8042), .A2(n10180), .ZN(n8033) );
  INV_X1 U5801 ( .A(n8031), .ZN(n8062) );
  AND2_X1 U5802 ( .A1(n7043), .A2(n7001), .ZN(n8043) );
  AND2_X1 U5803 ( .A1(n7437), .A2(n7436), .ZN(n8039) );
  NOR2_X1 U5804 ( .A1(n7885), .A2(n5049), .ZN(n8061) );
  OR2_X1 U5805 ( .A1(n7885), .A2(n4664), .ZN(n8059) );
  INV_X1 U5806 ( .A(n8050), .ZN(n8058) );
  INV_X1 U5807 ( .A(n8003), .ZN(n8067) );
  XNOR2_X1 U5808 ( .A(n5962), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6833) );
  AND3_X1 U5809 ( .A1(n5985), .A2(n5984), .A3(n5983), .ZN(n8344) );
  INV_X1 U5810 ( .A(n4972), .ZN(n7130) );
  OAI21_X1 U5811 ( .B1(n7052), .B2(n4970), .A(n4969), .ZN(n7594) );
  NAND2_X1 U5812 ( .A1(n4973), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4970) );
  NAND2_X1 U5813 ( .A1(n7131), .A2(n4973), .ZN(n4969) );
  INV_X1 U5814 ( .A(n7131), .ZN(n4971) );
  AND2_X1 U5815 ( .A1(n6083), .A2(n6112), .ZN(n10100) );
  INV_X1 U5816 ( .A(n4829), .ZN(n10132) );
  AND2_X1 U5817 ( .A1(n10142), .A2(n10141), .ZN(n10145) );
  NOR2_X1 U5818 ( .A1(n7661), .A2(n7662), .ZN(n7664) );
  INV_X1 U5819 ( .A(n4560), .ZN(n7660) );
  INV_X1 U5820 ( .A(n4572), .ZN(n7793) );
  INV_X1 U5821 ( .A(n4585), .ZN(n7797) );
  NOR2_X1 U5822 ( .A1(n7784), .A2(n7785), .ZN(n7788) );
  INV_X1 U5823 ( .A(n4963), .ZN(n7783) );
  NAND2_X1 U5824 ( .A1(n4958), .A2(n8115), .ZN(n8109) );
  OR2_X1 U5825 ( .A1(n8188), .A2(n8836), .ZN(n4977) );
  NAND2_X1 U5826 ( .A1(n4975), .A2(n4974), .ZN(n8232) );
  AND2_X1 U5827 ( .A1(n4977), .A2(n4482), .ZN(n8210) );
  NAND2_X1 U5828 ( .A1(n4570), .A2(n4567), .ZN(n8228) );
  NAND2_X1 U5829 ( .A1(n8226), .A2(n8239), .ZN(n4570) );
  NOR2_X1 U5830 ( .A1(n4491), .A2(n4568), .ZN(n4567) );
  OAI21_X1 U5831 ( .B1(n6790), .B2(n4997), .A(n4995), .ZN(n8266) );
  NAND2_X1 U5832 ( .A1(n4795), .A2(n4800), .ZN(n8274) );
  AOI21_X1 U5833 ( .B1(n8295), .B2(n6441), .A(n6440), .ZN(n8283) );
  NAND2_X1 U5834 ( .A1(n4565), .A2(n4564), .ZN(n4563) );
  XNOR2_X1 U5835 ( .A(n8289), .B(n8296), .ZN(n4566) );
  NAND2_X1 U5836 ( .A1(n8290), .A2(n8435), .ZN(n4564) );
  NAND2_X1 U5837 ( .A1(n5968), .A2(n5967), .ZN(n8304) );
  NAND2_X1 U5838 ( .A1(n4980), .A2(n4984), .ZN(n8331) );
  NAND2_X1 U5839 ( .A1(n8355), .A2(n4986), .ZN(n4980) );
  OAI21_X1 U5840 ( .B1(n8372), .B2(n4821), .A(n4818), .ZN(n8336) );
  NAND2_X1 U5841 ( .A1(n4825), .A2(n6428), .ZN(n8360) );
  NAND2_X1 U5842 ( .A1(n5010), .A2(n5007), .ZN(n8381) );
  INV_X1 U5843 ( .A(n5009), .ZN(n5007) );
  NAND2_X1 U5844 ( .A1(n6237), .A2(n6236), .ZN(n8511) );
  NAND2_X1 U5845 ( .A1(n5014), .A2(n5013), .ZN(n8391) );
  NAND2_X1 U5846 ( .A1(n8417), .A2(n6778), .ZN(n8402) );
  INV_X1 U5847 ( .A(n4806), .ZN(n8416) );
  AOI21_X1 U5848 ( .B1(n4812), .B2(n4810), .A(n4809), .ZN(n4806) );
  NAND2_X1 U5849 ( .A1(n6207), .A2(n6206), .ZN(n8430) );
  NAND2_X1 U5850 ( .A1(n6192), .A2(n6191), .ZN(n9632) );
  NAND2_X1 U5851 ( .A1(n4812), .A2(n4813), .ZN(n8445) );
  NAND2_X1 U5852 ( .A1(n6422), .A2(n6421), .ZN(n8460) );
  NAND2_X1 U5853 ( .A1(n7569), .A2(n6475), .ZN(n7728) );
  OAI21_X1 U5854 ( .B1(n7572), .B2(n4469), .A(n5027), .ZN(n7712) );
  AND2_X1 U5855 ( .A1(n6115), .A2(n6114), .ZN(n7532) );
  INV_X1 U5856 ( .A(n7447), .ZN(n10201) );
  INV_X1 U5857 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7179) );
  CLKBUF_X1 U5858 ( .A(n8457), .Z(n10167) );
  INV_X1 U5859 ( .A(n6449), .ZN(n8522) );
  AND2_X1 U5860 ( .A1(n5925), .A2(n5924), .ZN(n8542) );
  AND2_X1 U5861 ( .A1(n6269), .A2(n6268), .ZN(n8864) );
  NAND2_X1 U5862 ( .A1(n6801), .A2(n6808), .ZN(n7030) );
  NAND2_X1 U5863 ( .A1(n6502), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6498) );
  INV_X1 U5864 ( .A(n10100), .ZN(n7626) );
  NAND2_X1 U5865 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n6004) );
  NAND2_X1 U5866 ( .A1(n4856), .A2(n5171), .ZN(n7104) );
  NAND2_X1 U5867 ( .A1(n5598), .A2(n5597), .ZN(n9507) );
  XNOR2_X1 U5868 ( .A(n5142), .B(n5140), .ZN(n6988) );
  INV_X1 U5869 ( .A(n4876), .ZN(n8948) );
  INV_X1 U5870 ( .A(n4583), .ZN(n8950) );
  NAND2_X1 U5871 ( .A1(n5771), .A2(n5770), .ZN(n9259) );
  NAND2_X1 U5872 ( .A1(n4870), .A2(n5558), .ZN(n8973) );
  NAND2_X1 U5873 ( .A1(n8903), .A2(n4871), .ZN(n4870) );
  INV_X1 U5874 ( .A(n4872), .ZN(n4871) );
  NAND2_X1 U5875 ( .A1(n5744), .A2(n5743), .ZN(n9478) );
  INV_X1 U5876 ( .A(n7103), .ZN(n4855) );
  AND4_X1 U5877 ( .A1(n5441), .A2(n5440), .A3(n5439), .A4(n5438), .ZN(n9844)
         );
  INV_X1 U5878 ( .A(n9005), .ZN(n4851) );
  AND4_X1 U5879 ( .A1(n5402), .A2(n5401), .A3(n5400), .A4(n5399), .ZN(n9845)
         );
  AND4_X1 U5880 ( .A1(n5305), .A2(n5304), .A3(n5303), .A4(n5302), .ZN(n7552)
         );
  NAND2_X1 U5881 ( .A1(n7320), .A2(n5262), .ZN(n7347) );
  INV_X1 U5882 ( .A(n9244), .ZN(n9463) );
  NOR2_X1 U5883 ( .A1(n9035), .A2(n9036), .ZN(n4875) );
  OR2_X1 U5884 ( .A1(n7088), .A2(n5150), .ZN(n5540) );
  OR2_X1 U5885 ( .A1(n6745), .A2(n4550), .ZN(n6746) );
  AOI21_X1 U5886 ( .B1(n6597), .B2(n6591), .A(n4512), .ZN(n6592) );
  INV_X1 U5887 ( .A(n6736), .ZN(n4586) );
  AND2_X1 U5888 ( .A1(n6683), .A2(n4722), .ZN(n4579) );
  AND4_X1 U5889 ( .A1(n5353), .A2(n5352), .A3(n5351), .A4(n5350), .ZN(n8926)
         );
  INV_X1 U5890 ( .A(n4715), .ZN(n9713) );
  NOR2_X1 U5891 ( .A1(n9608), .A2(n4710), .ZN(n6923) );
  AND2_X1 U5892 ( .A1(n6950), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4710) );
  NAND2_X1 U5893 ( .A1(n6923), .A2(n6924), .ZN(n9121) );
  XNOR2_X1 U5894 ( .A(n9127), .B(n9128), .ZN(n9790) );
  NOR2_X1 U5895 ( .A1(n9798), .A2(n4546), .ZN(n9813) );
  NAND2_X1 U5896 ( .A1(n9813), .A2(n9812), .ZN(n9811) );
  AND2_X1 U5897 ( .A1(n9811), .A2(n4707), .ZN(n9826) );
  OR2_X1 U5898 ( .A1(n9819), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4707) );
  INV_X1 U5899 ( .A(n9797), .ZN(n9825) );
  INV_X1 U5900 ( .A(n9294), .ZN(n4722) );
  NAND2_X1 U5901 ( .A1(n4470), .A2(n9829), .ZN(n4724) );
  NAND2_X1 U5902 ( .A1(n4720), .A2(n9094), .ZN(n4719) );
  NAND2_X1 U5903 ( .A1(n9803), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4720) );
  OR2_X1 U5904 ( .A1(n4947), .A2(n4946), .ZN(n4942) );
  AOI21_X1 U5905 ( .B1(n7812), .B2(n6583), .A(n6576), .ZN(n9205) );
  OAI21_X1 U5906 ( .B1(n9209), .B2(n9193), .A(n9192), .ZN(n9194) );
  NAND2_X1 U5907 ( .A1(n5856), .A2(n5855), .ZN(n9450) );
  AND2_X1 U5908 ( .A1(n9215), .A2(n9214), .ZN(n9448) );
  AND2_X1 U5909 ( .A1(n4696), .A2(n6571), .ZN(n9235) );
  NAND2_X1 U5910 ( .A1(n4691), .A2(n4692), .ZN(n9233) );
  AND4_X1 U5911 ( .A1(n5752), .A2(n5751), .A3(n5750), .A4(n5749), .ZN(n9469)
         );
  NAND2_X1 U5912 ( .A1(n4756), .A2(n4467), .ZN(n9256) );
  NAND2_X1 U5913 ( .A1(n9169), .A2(n4471), .ZN(n4756) );
  NAND2_X1 U5914 ( .A1(n4706), .A2(n4705), .ZN(n9271) );
  AND2_X1 U5915 ( .A1(n4758), .A2(n4760), .ZN(n9270) );
  NAND2_X1 U5916 ( .A1(n9169), .A2(n9168), .ZN(n4758) );
  NAND2_X1 U5917 ( .A1(n5720), .A2(n5719), .ZN(n9299) );
  NAND2_X1 U5918 ( .A1(n9340), .A2(n6669), .ZN(n9320) );
  AND2_X1 U5919 ( .A1(n4733), .A2(n4736), .ZN(n9348) );
  AND2_X1 U5920 ( .A1(n4698), .A2(n6666), .ZN(n9367) );
  NAND2_X1 U5921 ( .A1(n9155), .A2(n4737), .ZN(n9365) );
  NAND2_X1 U5922 ( .A1(n4689), .A2(n6660), .ZN(n9418) );
  NAND2_X1 U5923 ( .A1(n4768), .A2(n4766), .ZN(n9425) );
  NAND2_X1 U5924 ( .A1(n7745), .A2(n4769), .ZN(n4768) );
  NAND2_X1 U5925 ( .A1(n7583), .A2(n6659), .ZN(n7750) );
  NAND2_X1 U5926 ( .A1(n4770), .A2(n4773), .ZN(n9151) );
  OR2_X1 U5927 ( .A1(n7745), .A2(n7744), .ZN(n4770) );
  NAND2_X1 U5928 ( .A1(n4742), .A2(n4466), .ZN(n9846) );
  NAND2_X1 U5929 ( .A1(n4744), .A2(n4743), .ZN(n7588) );
  AOI21_X1 U5930 ( .B1(n7485), .B2(n7484), .A(n4748), .ZN(n7510) );
  OAI211_X1 U5931 ( .C1(n7306), .C2(n4612), .A(n4613), .B(n6689), .ZN(n9862)
         );
  OR2_X1 U5932 ( .A1(n9907), .A2(n7236), .ZN(n9896) );
  NAND2_X1 U5933 ( .A1(n7304), .A2(n6526), .ZN(n7286) );
  INV_X1 U5934 ( .A(n9896), .ZN(n9854) );
  XNOR2_X1 U5936 ( .A(n6326), .B(n6325), .ZN(n9559) );
  XNOR2_X1 U5937 ( .A(n5736), .B(n5735), .ZN(n7656) );
  NAND2_X1 U5938 ( .A1(n4920), .A2(n4925), .ZN(n5736) );
  NAND2_X1 U5939 ( .A1(n5688), .A2(n4927), .ZN(n4920) );
  NAND2_X1 U5940 ( .A1(n4896), .A2(n4900), .ZN(n5458) );
  NAND2_X1 U5941 ( .A1(n5420), .A2(n4903), .ZN(n4896) );
  NAND2_X1 U5942 ( .A1(n4904), .A2(n4903), .ZN(n5452) );
  NAND2_X1 U5943 ( .A1(n4904), .A2(n4905), .ZN(n5425) );
  OR2_X1 U5944 ( .A1(n5386), .A2(n5387), .ZN(n5388) );
  AND2_X1 U5945 ( .A1(n5393), .A2(n5427), .ZN(n9575) );
  NAND2_X1 U5946 ( .A1(n5296), .A2(n5295), .ZN(n5316) );
  OR2_X1 U5947 ( .A1(n5296), .A2(n5295), .ZN(n5297) );
  NAND2_X1 U5948 ( .A1(n5290), .A2(n5289), .ZN(n5296) );
  INV_X1 U5949 ( .A(n6929), .ZN(n9672) );
  NOR2_X2 U5950 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7223) );
  NAND2_X1 U5951 ( .A1(n10041), .A2(n4548), .ZN(n10035) );
  INV_X1 U5952 ( .A(n4557), .ZN(n8155) );
  INV_X1 U5953 ( .A(n4962), .ZN(n8167) );
  INV_X1 U5954 ( .A(n8243), .ZN(n4576) );
  OAI21_X1 U5955 ( .B1(n5034), .B2(n4788), .A(n6824), .ZN(n6826) );
  CLKBUF_X2 U5956 ( .A(n9064), .Z(P1_U3973) );
  NAND2_X1 U5957 ( .A1(n4721), .A2(n4718), .ZN(P1_U3262) );
  NAND2_X1 U5958 ( .A1(n4723), .A2(n4722), .ZN(n4721) );
  AOI21_X1 U5959 ( .B1(n9136), .B2(n9294), .A(n4719), .ZN(n4718) );
  NAND2_X1 U5960 ( .A1(n9134), .A2(n4724), .ZN(n4723) );
  INV_X1 U5961 ( .A(n8372), .ZN(n4815) );
  AND2_X1 U5962 ( .A1(n4950), .A2(n9152), .ZN(n4464) );
  NOR2_X1 U5963 ( .A1(n9450), .A2(n9236), .ZN(n9193) );
  INV_X1 U5964 ( .A(n9193), .ZN(n4887) );
  NOR2_X1 U5965 ( .A1(n4821), .A2(n4817), .ZN(n4465) );
  NOR2_X1 U5966 ( .A1(n8299), .A2(n8303), .ZN(n6440) );
  OR2_X1 U5967 ( .A1(n7587), .A2(n4741), .ZN(n4466) );
  OR2_X1 U5968 ( .A1(n4757), .A2(n9171), .ZN(n4467) );
  INV_X1 U5969 ( .A(n8082), .ZN(n7714) );
  NAND2_X1 U5970 ( .A1(n5569), .A2(n5568), .ZN(n9385) );
  AND2_X1 U5971 ( .A1(n9331), .A2(n9342), .ZN(n6727) );
  AND2_X1 U5972 ( .A1(n9514), .A2(n9506), .ZN(n9157) );
  AND2_X1 U5973 ( .A1(n4951), .A2(n4774), .ZN(n4468) );
  OR2_X1 U5974 ( .A1(n6322), .A2(n8267), .ZN(n6442) );
  NOR2_X1 U5975 ( .A1(n7714), .A2(n7562), .ZN(n4469) );
  INV_X1 U5976 ( .A(n7178), .ZN(n4776) );
  NAND2_X1 U5977 ( .A1(n6301), .A2(n6300), .ZN(n8299) );
  XOR2_X1 U5978 ( .A(n9113), .B(n9112), .Z(n4470) );
  AND2_X1 U5979 ( .A1(n4759), .A2(n9168), .ZN(n4471) );
  INV_X1 U5980 ( .A(n9213), .ZN(n4731) );
  AND2_X1 U5981 ( .A1(n4468), .A2(n4950), .ZN(n4472) );
  OR2_X1 U5982 ( .A1(n6848), .A2(n9657), .ZN(n4473) );
  INV_X1 U5983 ( .A(n4985), .ZN(n4984) );
  OAI21_X1 U5984 ( .B1(n8349), .B2(n4990), .A(n4989), .ZN(n4985) );
  AND2_X1 U5985 ( .A1(n6647), .A2(n4502), .ZN(n4474) );
  INV_X1 U5986 ( .A(n8074), .ZN(n8281) );
  NAND2_X1 U5987 ( .A1(n6352), .A2(n6351), .ZN(n8074) );
  AND2_X1 U5988 ( .A1(n4954), .A2(n7586), .ZN(n4475) );
  OAI211_X1 U5989 ( .C1(n4523), .C2(n6520), .A(n4887), .B(n4886), .ZN(n4885)
         );
  INV_X1 U5990 ( .A(n9450), .ZN(n9217) );
  NAND2_X1 U5991 ( .A1(n6857), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4476) );
  NAND2_X1 U5992 ( .A1(n4816), .A2(n6432), .ZN(n4477) );
  AND3_X1 U5993 ( .A1(n4587), .A2(n6675), .A3(n9195), .ZN(n4478) );
  OR2_X1 U5994 ( .A1(n4671), .A2(n4669), .ZN(n4479) );
  INV_X1 U5995 ( .A(n6429), .ZN(n4826) );
  AND2_X1 U5996 ( .A1(n5257), .A2(n5229), .ZN(n4480) );
  OAI21_X1 U5997 ( .B1(n4891), .B2(n4890), .A(n4538), .ZN(n4889) );
  NAND2_X1 U5998 ( .A1(n7169), .A2(n7039), .ZN(n4481) );
  NAND2_X1 U5999 ( .A1(n7561), .A2(n4650), .ZN(n7830) );
  NAND2_X1 U6000 ( .A1(n5021), .A2(n5020), .ZN(n7478) );
  INV_X1 U6001 ( .A(n7534), .ZN(n4648) );
  INV_X1 U6002 ( .A(n7363), .ZN(n4652) );
  INV_X1 U6003 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9550) );
  AND2_X1 U6004 ( .A1(n7825), .A2(n5947), .ZN(n6019) );
  INV_X1 U6005 ( .A(n7139), .ZN(n4838) );
  OR2_X1 U6006 ( .A1(n8219), .A2(n8207), .ZN(n4482) );
  NAND2_X1 U6007 ( .A1(n4676), .A2(n4677), .ZN(n7893) );
  NAND2_X1 U6008 ( .A1(n8433), .A2(n6776), .ZN(n8417) );
  AND2_X1 U6009 ( .A1(n4799), .A2(n4803), .ZN(n4483) );
  NAND2_X1 U6010 ( .A1(n7451), .A2(n8040), .ZN(n4484) );
  AND4_X1 U6011 ( .A1(n6009), .A2(n6008), .A3(n6007), .A4(n6006), .ZN(n6757)
         );
  OR2_X1 U6012 ( .A1(n9444), .A2(n9443), .ZN(n4485) );
  NAND2_X1 U6013 ( .A1(n8085), .A2(n7438), .ZN(n4486) );
  AOI21_X1 U6014 ( .B1(n8875), .B2(n6583), .A(n6515), .ZN(n9437) );
  INV_X1 U6015 ( .A(n9437), .ZN(n4946) );
  AND2_X1 U6016 ( .A1(n4677), .A2(n4675), .ZN(n4487) );
  NAND2_X1 U6017 ( .A1(n5032), .A2(n5942), .ZN(n5944) );
  INV_X1 U6018 ( .A(n6781), .ZN(n5012) );
  OR2_X1 U6019 ( .A1(n7792), .A2(n7791), .ZN(n4488) );
  XOR2_X1 U6020 ( .A(n5707), .B(n5866), .Z(n4489) );
  OR2_X1 U6021 ( .A1(n8526), .A2(n8074), .ZN(n4490) );
  AND3_X1 U6022 ( .A1(n8227), .A2(n10143), .A3(n8235), .ZN(n4491) );
  INV_X1 U6023 ( .A(n6659), .ZN(n4688) );
  INV_X1 U6024 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5030) );
  OR2_X1 U6025 ( .A1(n8277), .A2(n8074), .ZN(n4492) );
  OR2_X1 U6026 ( .A1(n9930), .A2(n9934), .ZN(n4493) );
  INV_X1 U6027 ( .A(n9524), .ZN(n4951) );
  AND2_X1 U6028 ( .A1(n5670), .A2(n5669), .ZN(n9331) );
  INV_X1 U6029 ( .A(n9331), .ZN(n9497) );
  NAND2_X1 U6030 ( .A1(n4775), .A2(n6003), .ZN(n6054) );
  INV_X1 U6031 ( .A(n8335), .ZN(n4982) );
  NAND2_X1 U6032 ( .A1(n6128), .A2(n4794), .ZN(n4494) );
  NAND2_X1 U6033 ( .A1(n6128), .A2(n5029), .ZN(n4495) );
  AND3_X1 U6034 ( .A1(n6291), .A2(n6290), .A3(n8345), .ZN(n4496) );
  AND3_X1 U6035 ( .A1(n5162), .A2(n5161), .A3(n5160), .ZN(n9930) );
  INV_X1 U6036 ( .A(n4903), .ZN(n4902) );
  NOR2_X1 U6037 ( .A1(n5424), .A2(n4906), .ZN(n4903) );
  AND2_X1 U6038 ( .A1(n4810), .A2(n8415), .ZN(n4497) );
  NAND2_X1 U6039 ( .A1(n5033), .A2(n6799), .ZN(n8258) );
  NAND2_X1 U6040 ( .A1(n6128), .A2(n5913), .ZN(n6266) );
  AND2_X1 U6041 ( .A1(n7829), .A2(n8082), .ZN(n4498) );
  INV_X1 U6042 ( .A(n8075), .ZN(n8303) );
  NAND2_X1 U6043 ( .A1(n6308), .A2(n6307), .ZN(n8075) );
  AND2_X1 U6044 ( .A1(n5199), .A2(n5198), .ZN(n4499) );
  AND2_X1 U6045 ( .A1(n5008), .A2(n5015), .ZN(n4500) );
  AND2_X1 U6046 ( .A1(n9478), .A2(n9170), .ZN(n4501) );
  AND2_X1 U6047 ( .A1(n6572), .A2(n6573), .ZN(n4502) );
  AND2_X1 U6048 ( .A1(n6603), .A2(n7687), .ZN(n4503) );
  AND2_X1 U6049 ( .A1(n9259), .A2(n9173), .ZN(n4504) );
  NOR2_X1 U6050 ( .A1(n8896), .A2(n8892), .ZN(n4505) );
  AND2_X1 U6051 ( .A1(n9156), .A2(n9358), .ZN(n4506) );
  AND2_X1 U6052 ( .A1(n6421), .A2(n4814), .ZN(n4507) );
  AND2_X1 U6053 ( .A1(n7262), .A2(n7255), .ZN(n4508) );
  AND2_X1 U6054 ( .A1(n6125), .A2(n6124), .ZN(n7562) );
  AND2_X1 U6055 ( .A1(n8084), .A2(n7447), .ZN(n4509) );
  INV_X1 U6056 ( .A(n6726), .ZN(n6669) );
  AND2_X1 U6057 ( .A1(n9524), .A2(n9150), .ZN(n4510) );
  INV_X1 U6058 ( .A(n9171), .ZN(n4759) );
  OR2_X1 U6059 ( .A1(n7597), .A2(n10078), .ZN(n4511) );
  AND2_X1 U6060 ( .A1(n6598), .A2(n6972), .ZN(n4512) );
  INV_X1 U6061 ( .A(n6440), .ZN(n4805) );
  AND2_X1 U6062 ( .A1(n4881), .A2(n4880), .ZN(n4879) );
  NOR2_X1 U6063 ( .A1(n9159), .A2(n9158), .ZN(n4513) );
  AND2_X1 U6064 ( .A1(n7440), .A2(n8085), .ZN(n4514) );
  OR2_X1 U6065 ( .A1(n8430), .A2(n8404), .ZN(n6425) );
  AND3_X1 U6066 ( .A1(n6499), .A2(n6494), .A3(n6497), .ZN(n4515) );
  AND2_X1 U6067 ( .A1(n8550), .A2(n8344), .ZN(n4516) );
  INV_X1 U6068 ( .A(n4906), .ZN(n4905) );
  NOR2_X1 U6069 ( .A1(n5418), .A2(SI_11_), .ZN(n4906) );
  INV_X1 U6070 ( .A(n7863), .ZN(n4681) );
  AND2_X1 U6071 ( .A1(n7862), .A2(n8344), .ZN(n7863) );
  INV_X1 U6072 ( .A(n4751), .ZN(n4748) );
  NAND2_X1 U6073 ( .A1(n9965), .A2(n7647), .ZN(n4751) );
  AND2_X1 U6074 ( .A1(n8530), .A2(n8267), .ZN(n4517) );
  OR2_X1 U6075 ( .A1(n6726), .A2(n6619), .ZN(n4518) );
  INV_X1 U6076 ( .A(n8277), .ZN(n8526) );
  NAND2_X1 U6077 ( .A1(n6354), .A2(n6353), .ZN(n8277) );
  AND2_X1 U6078 ( .A1(n5341), .A2(n8772), .ZN(n4519) );
  NOR2_X1 U6079 ( .A1(n8281), .A2(n8277), .ZN(n4520) );
  NAND2_X1 U6080 ( .A1(n5943), .A2(n5944), .ZN(n5947) );
  INV_X1 U6081 ( .A(n4990), .ZN(n4988) );
  NAND2_X1 U6082 ( .A1(n8363), .A2(n8369), .ZN(n4990) );
  INV_X1 U6083 ( .A(n5295), .ZN(n4884) );
  INV_X1 U6084 ( .A(n6433), .ZN(n4817) );
  AND2_X1 U6085 ( .A1(n5091), .A2(n5065), .ZN(n4521) );
  AND2_X1 U6086 ( .A1(n5134), .A2(n5135), .ZN(n4522) );
  AND2_X1 U6087 ( .A1(n6521), .A2(n6644), .ZN(n4523) );
  AND2_X1 U6088 ( .A1(n9861), .A2(n4611), .ZN(n4524) );
  NAND2_X1 U6089 ( .A1(n5347), .A2(n5346), .ZN(n9972) );
  INV_X1 U6090 ( .A(n9172), .ZN(n4755) );
  INV_X1 U6091 ( .A(n4868), .ZN(n4867) );
  NAND2_X1 U6092 ( .A1(n5558), .A2(n4869), .ZN(n4868) );
  OR2_X1 U6093 ( .A1(n7931), .A2(n8333), .ZN(n6456) );
  INV_X1 U6094 ( .A(n6456), .ZN(n4819) );
  OR2_X1 U6095 ( .A1(n7901), .A2(n8081), .ZN(n4525) );
  NAND2_X1 U6096 ( .A1(n6424), .A2(n6214), .ZN(n8444) );
  INV_X1 U6097 ( .A(n8444), .ZN(n4811) );
  OR2_X1 U6098 ( .A1(n6734), .A2(n6733), .ZN(n4526) );
  NOR2_X1 U6099 ( .A1(n8942), .A2(n4849), .ZN(n4527) );
  AND2_X1 U6100 ( .A1(n4492), .A2(n4995), .ZN(n4528) );
  INV_X1 U6101 ( .A(n6423), .ZN(n4814) );
  INV_X1 U6102 ( .A(n7941), .ZN(n4638) );
  NAND2_X1 U6103 ( .A1(n6443), .A2(n6371), .ZN(n6793) );
  AND2_X1 U6104 ( .A1(n4946), .A2(n6672), .ZN(n6598) );
  AND2_X1 U6105 ( .A1(n9437), .A2(n9140), .ZN(n6738) );
  INV_X1 U6106 ( .A(n6738), .ZN(n4587) );
  AND2_X1 U6107 ( .A1(n4800), .A2(n4490), .ZN(n4529) );
  AND2_X1 U6108 ( .A1(n6419), .A2(n4785), .ZN(n4530) );
  NAND2_X1 U6109 ( .A1(n9228), .A2(n9252), .ZN(n9191) );
  NOR2_X1 U6110 ( .A1(n4941), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n4940) );
  AND2_X1 U6111 ( .A1(n8127), .A2(n8126), .ZN(n4531) );
  AND2_X1 U6112 ( .A1(n5914), .A2(n5028), .ZN(n4532) );
  OR2_X1 U6113 ( .A1(n8012), .A2(n8344), .ZN(n6432) );
  AND2_X1 U6114 ( .A1(n4515), .A2(n4792), .ZN(n4533) );
  AND2_X1 U6115 ( .A1(n9172), .A2(n4471), .ZN(n4534) );
  NAND2_X1 U6116 ( .A1(n5521), .A2(n5520), .ZN(n9520) );
  OR2_X1 U6117 ( .A1(n4674), .A2(n4670), .ZN(n4535) );
  INV_X1 U6118 ( .A(n5699), .ZN(n5248) );
  NAND2_X1 U6119 ( .A1(n6422), .A2(n4507), .ZN(n4812) );
  AND4_X1 U6120 ( .A1(n5470), .A2(n5469), .A3(n5468), .A4(n5467), .ZN(n8909)
         );
  OR2_X1 U6121 ( .A1(n6071), .A2(n6070), .ZN(n10078) );
  INV_X1 U6122 ( .A(n10078), .ZN(n4845) );
  INV_X1 U6123 ( .A(n10140), .ZN(n7629) );
  AND2_X1 U6124 ( .A1(n5689), .A2(n5687), .ZN(n4536) );
  INV_X1 U6125 ( .A(n7932), .ZN(n4684) );
  INV_X1 U6126 ( .A(n8333), .ZN(n8357) );
  NAND2_X1 U6127 ( .A1(n7694), .A2(n4472), .ZN(n4952) );
  INV_X1 U6128 ( .A(n4894), .ZN(n4893) );
  NOR2_X1 U6129 ( .A1(n5562), .A2(n4895), .ZN(n4894) );
  AND2_X1 U6130 ( .A1(n5561), .A2(n5560), .ZN(n4537) );
  OR2_X1 U6131 ( .A1(n5589), .A2(SI_17_), .ZN(n4538) );
  AND2_X1 U6132 ( .A1(n4894), .A2(n5590), .ZN(n4539) );
  INV_X1 U6133 ( .A(n9157), .ZN(n4736) );
  INV_X1 U6134 ( .A(n9167), .ZN(n4760) );
  XNOR2_X1 U6135 ( .A(n6498), .B(n6497), .ZN(n6802) );
  INV_X1 U6136 ( .A(n9426), .ZN(n4950) );
  NAND2_X1 U6137 ( .A1(n7256), .A2(n4508), .ZN(n7361) );
  OR2_X1 U6138 ( .A1(n7570), .A2(n7573), .ZN(n7569) );
  OR2_X1 U6139 ( .A1(n7382), .A2(n4957), .ZN(n4540) );
  OR2_X1 U6140 ( .A1(n9874), .A2(n7411), .ZN(n7382) );
  INV_X1 U6141 ( .A(n7382), .ZN(n4953) );
  INV_X1 U6142 ( .A(n7484), .ZN(n4747) );
  OR2_X1 U6143 ( .A1(n8154), .A2(n8446), .ZN(n4541) );
  OAI21_X1 U6144 ( .B1(n7175), .B2(n6763), .A(n6762), .ZN(n7196) );
  NAND2_X1 U6145 ( .A1(n7437), .A2(n4654), .ZN(n8037) );
  NAND2_X1 U6146 ( .A1(n7362), .A2(n7363), .ZN(n7437) );
  OR2_X1 U6147 ( .A1(n7382), .A2(n4955), .ZN(n4542) );
  AND2_X1 U6148 ( .A1(n4780), .A2(n6415), .ZN(n4543) );
  INV_X1 U6149 ( .A(n4612), .ZN(n4614) );
  OR2_X1 U6150 ( .A1(n4615), .A2(n6607), .ZN(n4612) );
  INV_X2 U6151 ( .A(n10238), .ZN(n10240) );
  AND2_X1 U6152 ( .A1(n5021), .A2(n4484), .ZN(n4544) );
  AND2_X1 U6153 ( .A1(n7561), .A2(n7560), .ZN(n4545) );
  INV_X1 U6154 ( .A(n6509), .ZN(n6755) );
  NAND2_X1 U6155 ( .A1(n7116), .A2(n7115), .ZN(n7256) );
  AND2_X1 U6156 ( .A1(n9807), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4546) );
  OR2_X1 U6157 ( .A1(n8239), .A2(n8715), .ZN(n4547) );
  OR2_X1 U6158 ( .A1(n10034), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n4548) );
  AND2_X1 U6159 ( .A1(n4972), .A2(n4971), .ZN(n4549) );
  OR3_X1 U6160 ( .A1(n9294), .A2(n7657), .A3(n6744), .ZN(n4550) );
  INV_X1 U6161 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n4831) );
  AOI211_X1 U6162 ( .C1(n9450), .C2(n4451), .A(n5898), .B(n5897), .ZN(n5899)
         );
  OAI21_X1 U6163 ( .B1(n6000), .B2(n6859), .A(n4574), .ZN(n5104) );
  NAND2_X1 U6164 ( .A1(n4551), .A2(n6484), .ZN(n6405) );
  NAND3_X1 U6165 ( .A1(n6401), .A2(n6402), .A3(n6448), .ZN(n4551) );
  NAND2_X1 U6166 ( .A1(n5274), .A2(n5273), .ZN(n5280) );
  AOI21_X1 U6167 ( .B1(n5367), .B2(n5366), .A(n5365), .ZN(n5386) );
  AOI21_X1 U6168 ( .B1(n4888), .B2(n4539), .A(n4889), .ZN(n5607) );
  OAI21_X1 U6169 ( .B1(n5688), .B2(n4924), .A(n4921), .ZN(n5738) );
  OR2_X1 U6170 ( .A1(n5104), .A2(SI_1_), .ZN(n5105) );
  NAND2_X1 U6171 ( .A1(n4704), .A2(n4702), .ZN(n9265) );
  NOR2_X1 U6172 ( .A1(n9264), .A2(n9189), .ZN(n9251) );
  OAI21_X1 U6173 ( .B1(n5678), .B2(n7311), .A(n5193), .ZN(n5194) );
  INV_X1 U6174 ( .A(n5876), .ZN(n8894) );
  NAND2_X1 U6175 ( .A1(n5479), .A2(n5478), .ZN(n5508) );
  NAND2_X1 U6176 ( .A1(n4848), .A2(n4847), .ZN(n4852) );
  OAI21_X2 U6177 ( .B1(n9004), .B2(n9008), .A(n8914), .ZN(n8980) );
  NAND2_X1 U6178 ( .A1(n5661), .A2(n4527), .ZN(n4848) );
  NAND2_X1 U6179 ( .A1(n7518), .A2(n6768), .ZN(n6771) );
  NAND2_X1 U6180 ( .A1(n5018), .A2(n5017), .ZN(n7518) );
  NAND2_X1 U6181 ( .A1(n5155), .A2(n5154), .ZN(n4552) );
  INV_X1 U6182 ( .A(n6000), .ZN(n6860) );
  MUX2_X1 U6183 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n6000), .Z(n5153) );
  AND2_X4 U6184 ( .A1(n5103), .A2(n5102), .ZN(n6000) );
  NAND2_X1 U6185 ( .A1(n5000), .A2(n5003), .ZN(n8279) );
  OAI21_X1 U6186 ( .B1(n8320), .B2(n6785), .A(n6784), .ZN(n8311) );
  AOI22_X1 U6187 ( .A1(n7701), .A2(n6773), .B1(n7708), .B2(n8454), .ZN(n8450)
         );
  NAND2_X1 U6188 ( .A1(n5970), .A2(n5969), .ZN(n6302) );
  AOI21_X1 U6189 ( .B1(n5042), .B2(n6488), .A(n7431), .ZN(n6487) );
  NOR2_X1 U6190 ( .A1(n8157), .A2(n8427), .ZN(n8164) );
  NAND2_X1 U6191 ( .A1(n4559), .A2(n4558), .ZN(n8107) );
  NOR2_X1 U6192 ( .A1(n10077), .A2(n10076), .ZN(n10075) );
  NOR2_X1 U6193 ( .A1(n10095), .A2(n10094), .ZN(n10093) );
  OR2_X2 U6194 ( .A1(n8118), .A2(n8117), .ZN(n4557) );
  INV_X1 U6195 ( .A(n8107), .ZN(n8105) );
  INV_X1 U6196 ( .A(n7788), .ZN(n4559) );
  NAND2_X1 U6197 ( .A1(n8107), .A2(n5051), .ZN(n8108) );
  NAND2_X1 U6198 ( .A1(n5124), .A2(n5125), .ZN(n4561) );
  AOI21_X2 U6199 ( .B1(n4848), .B2(n5686), .A(n4489), .ZN(n9008) );
  NAND2_X2 U6200 ( .A1(n4876), .A2(n4875), .ZN(n9039) );
  AOI21_X1 U6201 ( .B1(n8980), .B2(n8979), .A(n8978), .ZN(n8982) );
  NAND2_X1 U6202 ( .A1(n4979), .A2(n4978), .ZN(n8320) );
  AOI21_X1 U6203 ( .B1(n7730), .B2(n7834), .A(n6772), .ZN(n7701) );
  AOI21_X1 U6204 ( .B1(n8450), .B2(n6775), .A(n6774), .ZN(n8434) );
  OAI21_X1 U6205 ( .B1(n8311), .B2(n6787), .A(n6786), .ZN(n8301) );
  MUX2_X1 U6206 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(P1_DATAO_REG_0__SCAN_IN), 
        .S(n6000), .Z(n5106) );
  NAND2_X1 U6207 ( .A1(n4511), .A2(n7596), .ZN(n10077) );
  AOI21_X1 U6208 ( .B1(n8220), .B2(n8219), .A(n8218), .ZN(n8222) );
  NOR2_X1 U6209 ( .A1(n7134), .A2(n4581), .ZN(n7137) );
  XNOR2_X1 U6210 ( .A(n4577), .B(n4576), .ZN(n8255) );
  NOR2_X1 U6211 ( .A1(n7674), .A2(n7675), .ZN(n7676) );
  OR2_X2 U6212 ( .A1(n10093), .A2(n7600), .ZN(n7602) );
  NOR2_X1 U6213 ( .A1(n10256), .A2(n7616), .ZN(n7667) );
  INV_X1 U6214 ( .A(n7607), .ZN(n4846) );
  NOR2_X2 U6215 ( .A1(n7141), .A2(n7140), .ZN(n7144) );
  NAND2_X1 U6216 ( .A1(n8213), .A2(n4842), .ZN(n4840) );
  NAND2_X1 U6217 ( .A1(n4846), .A2(n7608), .ZN(n7610) );
  NOR2_X2 U6218 ( .A1(n7670), .A2(n7669), .ZN(n7762) );
  INV_X1 U6219 ( .A(n7074), .ZN(n4839) );
  NOR2_X1 U6220 ( .A1(n8212), .A2(n8213), .ZN(n8215) );
  AOI21_X1 U6221 ( .B1(n6163), .B2(n6162), .A(n6161), .ZN(n6164) );
  NAND2_X1 U6222 ( .A1(n6149), .A2(n6150), .ZN(n6163) );
  OAI21_X1 U6223 ( .B1(n4496), .B2(n4573), .A(n6455), .ZN(n6292) );
  NAND2_X1 U6224 ( .A1(n6405), .A2(n7431), .ZN(n6491) );
  OR2_X2 U6225 ( .A1(n6400), .A2(n6399), .ZN(n6401) );
  OAI21_X1 U6226 ( .B1(n6293), .B2(n6294), .A(n4575), .ZN(n6298) );
  NAND2_X2 U6227 ( .A1(n8904), .A2(n8905), .ZN(n8903) );
  NAND3_X1 U6228 ( .A1(n4975), .A2(n4547), .A3(n4974), .ZN(n4577) );
  NAND2_X1 U6229 ( .A1(n4595), .A2(n4593), .ZN(n4592) );
  NAND3_X1 U6230 ( .A1(n6750), .A2(n5050), .A3(n4578), .ZN(P1_U3242) );
  NAND3_X1 U6231 ( .A1(n6629), .A2(n6681), .A3(n4579), .ZN(n4578) );
  NAND2_X1 U6232 ( .A1(n4608), .A2(n4607), .ZN(n4606) );
  OAI21_X1 U6233 ( .B1(n6556), .B2(n6589), .A(n4599), .ZN(n4598) );
  NAND3_X1 U6234 ( .A1(n7305), .A2(n6689), .A3(n7306), .ZN(n4580) );
  NAND2_X1 U6235 ( .A1(n6567), .A2(n6589), .ZN(n4624) );
  INV_X1 U6236 ( .A(n7278), .ZN(n4588) );
  NAND2_X1 U6237 ( .A1(n4620), .A2(n4618), .ZN(n6574) );
  AOI21_X1 U6238 ( .B1(n4597), .B2(n6564), .A(n9309), .ZN(n6566) );
  NOR2_X1 U6239 ( .A1(n7768), .A2(n7769), .ZN(n7770) );
  NOR2_X1 U6240 ( .A1(n7801), .A2(n7802), .ZN(n8092) );
  NAND2_X1 U6241 ( .A1(n4622), .A2(n6569), .ZN(n4621) );
  NAND2_X1 U6242 ( .A1(n6580), .A2(n9195), .ZN(n4919) );
  NAND2_X1 U6243 ( .A1(n6553), .A2(n6972), .ZN(n4630) );
  NAND2_X1 U6244 ( .A1(n6532), .A2(n6531), .ZN(n4610) );
  NAND2_X2 U6245 ( .A1(n4583), .A2(n4582), .ZN(n4876) );
  OR2_X2 U6246 ( .A1(n8982), .A2(n5761), .ZN(n4583) );
  INV_X1 U6247 ( .A(n5171), .ZN(n4854) );
  NAND2_X1 U6248 ( .A1(n5164), .A2(n5163), .ZN(n5165) );
  NAND2_X1 U6249 ( .A1(n4852), .A2(n4851), .ZN(n4850) );
  NAND2_X1 U6250 ( .A1(n5489), .A2(n5058), .ZN(n5492) );
  NOR2_X1 U6251 ( .A1(n7664), .A2(n7663), .ZN(n7758) );
  NAND2_X1 U6252 ( .A1(n7595), .A2(n5052), .ZN(n7597) );
  INV_X1 U6253 ( .A(n7132), .ZN(n4973) );
  NAND2_X1 U6254 ( .A1(n4836), .A2(n4835), .ZN(n4834) );
  INV_X1 U6255 ( .A(n6003), .ZN(n6024) );
  NAND2_X1 U6256 ( .A1(n5107), .A2(n5108), .ZN(n5152) );
  NAND2_X1 U6257 ( .A1(n5237), .A2(n5236), .ZN(n5274) );
  NAND2_X1 U6258 ( .A1(n4877), .A2(n4878), .ZN(n5367) );
  NAND3_X1 U6259 ( .A1(n6628), .A2(n4478), .A3(n4586), .ZN(n6681) );
  NOR2_X1 U6260 ( .A1(n4933), .A2(n4591), .ZN(n4931) );
  NAND2_X1 U6261 ( .A1(n4931), .A2(n5112), .ZN(n7275) );
  INV_X1 U6262 ( .A(n6526), .ZN(n4615) );
  NAND2_X1 U6263 ( .A1(n5489), .A2(n4616), .ZN(n4617) );
  NAND2_X1 U6264 ( .A1(n4457), .A2(n4940), .ZN(n5097) );
  NAND3_X1 U6265 ( .A1(n4624), .A2(n4623), .A3(n9272), .ZN(n4622) );
  NAND2_X4 U6266 ( .A1(n4632), .A2(n7032), .ZN(n7090) );
  INV_X1 U6267 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n4634) );
  NAND2_X1 U6268 ( .A1(n7094), .A2(n7093), .ZN(n7095) );
  NAND3_X1 U6269 ( .A1(n4481), .A2(n7036), .A3(n7093), .ZN(n7094) );
  NAND3_X1 U6270 ( .A1(n7903), .A2(n7835), .A3(n7941), .ZN(n4635) );
  NAND2_X1 U6271 ( .A1(n8052), .A2(n4640), .ZN(n4639) );
  OAI211_X1 U6272 ( .C1(n8052), .C2(n4644), .A(n4641), .B(n4639), .ZN(n7930)
         );
  NAND2_X1 U6273 ( .A1(n8052), .A2(n7876), .ZN(n7879) );
  OAI21_X2 U6274 ( .B1(n7533), .B2(n4649), .A(n4647), .ZN(n7831) );
  AND2_X1 U6275 ( .A1(n8038), .A2(n7436), .ZN(n4654) );
  NOR2_X1 U6276 ( .A1(n4655), .A2(n5906), .ZN(n6128) );
  NAND3_X1 U6277 ( .A1(n4775), .A2(n6003), .A3(n5907), .ZN(n4655) );
  NOR2_X1 U6278 ( .A1(n4656), .A2(n5906), .ZN(n4658) );
  NAND3_X1 U6279 ( .A1(n4775), .A2(n6003), .A3(n4657), .ZN(n4656) );
  NOR2_X2 U6280 ( .A1(n6054), .A2(n5906), .ZN(n6122) );
  NAND2_X1 U6281 ( .A1(n5029), .A2(n4658), .ZN(n5963) );
  NAND2_X1 U6282 ( .A1(n7884), .A2(n4663), .ZN(n4662) );
  OAI21_X1 U6283 ( .B1(n7933), .B2(n4535), .A(n4479), .ZN(n4666) );
  NAND2_X1 U6284 ( .A1(n4689), .A2(n4686), .ZN(n9416) );
  INV_X1 U6285 ( .A(n4696), .ZN(n9249) );
  NAND2_X1 U6286 ( .A1(n9340), .A2(n4701), .ZN(n9180) );
  NAND2_X1 U6287 ( .A1(n9286), .A2(n4705), .ZN(n4704) );
  INV_X1 U6288 ( .A(n4706), .ZN(n9288) );
  NAND2_X2 U6289 ( .A1(n5280), .A2(n5279), .ZN(n5290) );
  MUX2_X1 U6290 ( .A(n8753), .B(P1_REG2_REG_1__SCAN_IN), .S(n6929), .Z(n9664)
         );
  NAND2_X1 U6291 ( .A1(n9178), .A2(n9177), .ZN(n9212) );
  NAND2_X1 U6292 ( .A1(n9178), .A2(n4728), .ZN(n9215) );
  OAI21_X2 U6293 ( .B1(n6875), .B2(n5150), .A(n5299), .ZN(n7456) );
  NAND2_X1 U6294 ( .A1(n9155), .A2(n4734), .ZN(n4733) );
  INV_X1 U6295 ( .A(n9385), .ZN(n4738) );
  INV_X1 U6296 ( .A(n9847), .ZN(n4739) );
  NAND3_X1 U6297 ( .A1(n4466), .A2(n4742), .A3(n4739), .ZN(n4740) );
  NAND3_X1 U6298 ( .A1(n4744), .A2(n4750), .A3(n4743), .ZN(n4742) );
  NAND2_X1 U6299 ( .A1(n4746), .A2(n7485), .ZN(n4743) );
  NAND2_X1 U6300 ( .A1(n9169), .A2(n4534), .ZN(n4752) );
  NAND2_X1 U6301 ( .A1(n7745), .A2(n4762), .ZN(n4761) );
  NOR2_X4 U6302 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6003) );
  NOR2_X1 U6303 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4775) );
  NAND2_X1 U6304 ( .A1(n4779), .A2(n6409), .ZN(n7177) );
  AOI22_X1 U6305 ( .A1(n4777), .A2(n4779), .B1(n4776), .B2(n6410), .ZN(n7198)
         );
  XNOR2_X1 U6306 ( .A(n8088), .B(n10179), .ZN(n7178) );
  AND2_X1 U6307 ( .A1(n6032), .A2(n6034), .ZN(n4778) );
  NAND2_X1 U6308 ( .A1(n7570), .A2(n6475), .ZN(n4784) );
  NAND2_X1 U6309 ( .A1(n4784), .A2(n4530), .ZN(n6420) );
  NAND2_X1 U6310 ( .A1(n6756), .A2(n4787), .ZN(n4786) );
  NAND2_X1 U6311 ( .A1(n6756), .A2(n6000), .ZN(n6038) );
  OAI21_X1 U6312 ( .B1(n6756), .B2(n10057), .A(n4786), .ZN(n7033) );
  NAND2_X1 U6313 ( .A1(n6756), .A2(n6857), .ZN(n6037) );
  AND2_X1 U6314 ( .A1(n6122), .A2(n4792), .ZN(n4791) );
  AND4_X2 U6315 ( .A1(n6122), .A2(n5913), .A3(n4793), .A4(n4533), .ZN(n6503)
         );
  NAND2_X1 U6316 ( .A1(n8295), .A2(n4529), .ZN(n4798) );
  NOR2_X2 U6317 ( .A1(n8384), .A2(n6427), .ZN(n8372) );
  NOR2_X1 U6318 ( .A1(n8396), .A2(n6426), .ZN(n8384) );
  NAND2_X2 U6319 ( .A1(n6406), .A2(n6407), .ZN(n7170) );
  OAI21_X1 U6320 ( .B1(n8265), .B2(n10163), .A(n6800), .ZN(n5034) );
  INV_X1 U6321 ( .A(n8126), .ZN(n4832) );
  NAND2_X1 U6322 ( .A1(n10063), .A2(n4838), .ZN(n4833) );
  NAND3_X1 U6323 ( .A1(n4834), .A2(n4837), .A3(n4833), .ZN(n7075) );
  MUX2_X1 U6324 ( .A(n8891), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  MUX2_X1 U6325 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8891), .S(n6756), .Z(n7037) );
  OAI21_X1 U6326 ( .B1(n8198), .B2(n4841), .A(n4840), .ZN(n8234) );
  AOI21_X1 U6327 ( .B1(n7144), .B2(n7608), .A(n4843), .ZN(n7611) );
  NOR2_X1 U6328 ( .A1(n7144), .A2(n7143), .ZN(n7607) );
  NAND2_X1 U6329 ( .A1(n5661), .A2(n5660), .ZN(n8941) );
  INV_X1 U6330 ( .A(n5660), .ZN(n4849) );
  INV_X1 U6331 ( .A(n4852), .ZN(n9006) );
  INV_X1 U6332 ( .A(n4850), .ZN(n9004) );
  OAI21_X2 U6333 ( .B1(n4856), .B2(n4855), .A(n4853), .ZN(n7243) );
  NAND2_X1 U6334 ( .A1(n7020), .A2(n7021), .ZN(n4856) );
  INV_X1 U6335 ( .A(n4862), .ZN(n4861) );
  OAI21_X1 U6336 ( .B1(n4865), .B2(n4863), .A(n7418), .ZN(n4862) );
  OR2_X1 U6337 ( .A1(n7344), .A2(n7345), .ZN(n4865) );
  OAI211_X2 U6338 ( .C1(n8903), .C2(n4868), .A(n4866), .B(n8969), .ZN(n8931)
         );
  NAND2_X1 U6339 ( .A1(n5613), .A2(n5082), .ZN(n5616) );
  NAND2_X1 U6340 ( .A1(n5613), .A2(n4874), .ZN(n5117) );
  NAND2_X1 U6341 ( .A1(n7241), .A2(n5229), .ZN(n5261) );
  NAND2_X2 U6342 ( .A1(n5226), .A2(n5225), .ZN(n7241) );
  NAND2_X1 U6343 ( .A1(n7241), .A2(n4480), .ZN(n7319) );
  NAND2_X1 U6344 ( .A1(n5290), .A2(n4879), .ZN(n4877) );
  INV_X1 U6345 ( .A(n5533), .ZN(n4888) );
  NAND2_X1 U6346 ( .A1(n5533), .A2(n5532), .ZN(n5535) );
  OAI21_X1 U6347 ( .B1(n5688), .B2(n4536), .A(n5691), .ZN(n5713) );
  NAND4_X1 U6348 ( .A1(n5056), .A2(n5057), .A3(n5055), .A4(n4929), .ZN(n4930)
         );
  NAND3_X1 U6349 ( .A1(n5159), .A2(n5053), .A3(n5181), .ZN(n5239) );
  NAND4_X1 U6350 ( .A1(n5159), .A2(n5053), .A3(n5181), .A4(n5054), .ZN(n5241)
         );
  NOR2_X2 U6351 ( .A1(n5241), .A2(n4930), .ZN(n5489) );
  NAND2_X1 U6352 ( .A1(n4932), .A2(n9930), .ZN(n7297) );
  NAND3_X1 U6353 ( .A1(n4931), .A2(n5112), .A3(n9901), .ZN(n9899) );
  NOR2_X1 U6354 ( .A1(n6884), .A2(n9672), .ZN(n4933) );
  NAND2_X1 U6355 ( .A1(n9335), .A2(n4934), .ZN(n4937) );
  INV_X1 U6356 ( .A(n4937), .ZN(n9292) );
  NAND2_X1 U6357 ( .A1(n4457), .A2(n4938), .ZN(n5070) );
  NAND2_X1 U6358 ( .A1(n4457), .A2(n5064), .ZN(n5087) );
  AND2_X1 U6359 ( .A1(n9227), .A2(n4949), .ZN(n9201) );
  NAND2_X1 U6360 ( .A1(n9227), .A2(n9217), .ZN(n9216) );
  NAND2_X1 U6361 ( .A1(n9227), .A2(n4947), .ZN(n9144) );
  NAND3_X1 U6362 ( .A1(n4944), .A2(n4943), .A3(n4942), .ZN(n9137) );
  NAND2_X1 U6363 ( .A1(n4945), .A2(n9227), .ZN(n4944) );
  NAND3_X1 U6364 ( .A1(n9405), .A2(n4472), .A3(n7694), .ZN(n9390) );
  INV_X1 U6365 ( .A(n4952), .ZN(n9428) );
  INV_X1 U6366 ( .A(n4959), .ZN(n8116) );
  AND2_X2 U6367 ( .A1(n4962), .A2(n4961), .ZN(n8187) );
  XNOR2_X1 U6368 ( .A(n7129), .B(n7139), .ZN(n7052) );
  INV_X1 U6369 ( .A(n4977), .ZN(n8208) );
  NAND2_X1 U6370 ( .A1(n8355), .A2(n4981), .ZN(n4979) );
  OR2_X1 U6371 ( .A1(n7931), .A2(n8357), .ZN(n4989) );
  NAND2_X1 U6372 ( .A1(n6790), .A2(n4528), .ZN(n4991) );
  NAND2_X1 U6373 ( .A1(n4991), .A2(n4992), .ZN(n6794) );
  NAND2_X1 U6374 ( .A1(n6790), .A2(n5001), .ZN(n5000) );
  NAND2_X1 U6375 ( .A1(n6790), .A2(n6789), .ZN(n8289) );
  NAND3_X1 U6376 ( .A1(n4995), .A2(n4997), .A3(n4492), .ZN(n4994) );
  INV_X1 U6377 ( .A(n7403), .ZN(n5022) );
  NAND2_X1 U6378 ( .A1(n7572), .A2(n5026), .ZN(n5023) );
  NAND2_X1 U6379 ( .A1(n5023), .A2(n5024), .ZN(n7730) );
  INV_X1 U6380 ( .A(n5032), .ZN(n5941) );
  NOR2_X2 U6381 ( .A1(n5921), .A2(n5031), .ZN(n5032) );
  NAND4_X1 U6382 ( .A1(n6799), .A2(n5039), .A3(n10240), .A4(n5033), .ZN(n6844)
         );
  INV_X4 U6383 ( .A(n6000), .ZN(n6857) );
  NAND2_X1 U6384 ( .A1(n4887), .A2(n9192), .ZN(n9213) );
  INV_X2 U6385 ( .A(n5247), .ZN(n5885) );
  CLKBUF_X1 U6386 ( .A(n5492), .Z(n5536) );
  OAI21_X2 U6387 ( .B1(n8026), .B2(n7915), .A(n7914), .ZN(n7913) );
  AOI21_X2 U6388 ( .B1(n7852), .B2(n7851), .A(n7850), .ZN(n7971) );
  XNOR2_X2 U6389 ( .A(n7275), .B(n9065), .ZN(n9885) );
  AOI22_X2 U6390 ( .A1(n7989), .A2(n7860), .B1(n7859), .B2(n8369), .ZN(n7933)
         );
  NAND2_X1 U6391 ( .A1(n8434), .A2(n8444), .ZN(n8433) );
  NAND2_X1 U6392 ( .A1(n6493), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6495) );
  AND2_X1 U6393 ( .A1(n8868), .A2(n8368), .ZN(n5036) );
  OR2_X1 U6394 ( .A1(n8259), .A2(n8873), .ZN(n5037) );
  OR2_X1 U6395 ( .A1(n8265), .A2(n10202), .ZN(n5039) );
  OR2_X1 U6396 ( .A1(n8259), .A2(n8519), .ZN(n5041) );
  AND3_X1 U6397 ( .A1(n6486), .A2(n6485), .A3(n6484), .ZN(n5042) );
  AND2_X1 U6398 ( .A1(n5918), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5043) );
  AND2_X1 U6399 ( .A1(n7696), .A2(n9844), .ZN(n5044) );
  NAND3_X1 U6400 ( .A1(n8619), .A2(n5537), .A3(n5081), .ZN(n5045) );
  OR2_X1 U6401 ( .A1(n9331), .A2(n9488), .ZN(n5046) );
  AND2_X1 U6402 ( .A1(n5497), .A2(n5496), .ZN(n5047) );
  AND2_X1 U6403 ( .A1(n4571), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5048) );
  AND2_X1 U6404 ( .A1(n7846), .A2(n8453), .ZN(n5049) );
  INV_X1 U6405 ( .A(n7997), .ZN(n7842) );
  AND4_X1 U6406 ( .A1(n5547), .A2(n5546), .A3(n5545), .A4(n5544), .ZN(n9152)
         );
  INV_X1 U6407 ( .A(n8404), .ZN(n6777) );
  INV_X1 U6408 ( .A(n7908), .ZN(n7836) );
  AND4_X1 U6409 ( .A1(n6749), .A2(n6748), .A3(n6747), .A4(n6746), .ZN(n5050)
         );
  OR2_X1 U6410 ( .A1(n8106), .A2(n7786), .ZN(n5051) );
  OR2_X1 U6411 ( .A1(n7624), .A2(n8717), .ZN(n5052) );
  AND2_X1 U6412 ( .A1(n6796), .A2(n6795), .ZN(n8451) );
  INV_X1 U6413 ( .A(n8451), .ZN(n6797) );
  INV_X1 U6414 ( .A(n7165), .ZN(n6488) );
  INV_X1 U6415 ( .A(n5877), .ZN(n5872) );
  NAND2_X1 U6416 ( .A1(n6376), .A2(n6375), .ZN(n6377) );
  INV_X1 U6417 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5916) );
  INV_X1 U6418 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5907) );
  INV_X1 U6419 ( .A(n6727), .ZN(n6670) );
  INV_X1 U6420 ( .A(n8436), .ZN(n7841) );
  INV_X1 U6421 ( .A(n7445), .ZN(n7442) );
  INV_X1 U6422 ( .A(n7796), .ZN(n7794) );
  NAND2_X1 U6423 ( .A1(n9184), .A2(n9287), .ZN(n9185) );
  INV_X1 U6424 ( .A(n9424), .ZN(n6662) );
  INV_X1 U6425 ( .A(n6238), .ZN(n5936) );
  AND2_X1 U6426 ( .A1(n8418), .A2(n8419), .ZN(n6776) );
  OR2_X1 U6427 ( .A1(n6037), .A2(n6862), .ZN(n6028) );
  NOR2_X1 U6428 ( .A1(n9205), .A2(n9210), .ZN(n6578) );
  OR2_X1 U6429 ( .A1(n5436), .A2(n5435), .ZN(n5465) );
  INV_X1 U6430 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5058) );
  INV_X1 U6431 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5054) );
  INV_X1 U6432 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5101) );
  INV_X1 U6433 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U6434 ( .A1(n7837), .A2(n7836), .ZN(n7838) );
  XNOR2_X1 U6435 ( .A(n7831), .B(n7832), .ZN(n7902) );
  OR2_X1 U6436 ( .A1(n5991), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5982) );
  INV_X1 U6437 ( .A(n8146), .ZN(n8128) );
  INV_X1 U6438 ( .A(n5971), .ZN(n5970) );
  NAND2_X1 U6439 ( .A1(n6833), .A2(n7165), .ZN(n6839) );
  OAI21_X1 U6440 ( .B1(n7196), .B2(n6765), .A(n6764), .ZN(n7390) );
  OR2_X1 U6441 ( .A1(n6177), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n6251) );
  INV_X1 U6442 ( .A(n7244), .ZN(n5225) );
  INV_X1 U6443 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5263) );
  INV_X1 U6444 ( .A(n6578), .ZN(n6674) );
  AND2_X1 U6445 ( .A1(n5396), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5398) );
  INV_X1 U6446 ( .A(n7544), .ZN(n6743) );
  NAND2_X1 U6447 ( .A1(n5421), .A2(SI_12_), .ZN(n5451) );
  NAND2_X1 U6448 ( .A1(n5232), .A2(SI_5_), .ZN(n5273) );
  NAND2_X1 U6449 ( .A1(n5930), .A2(n5929), .ZN(n6106) );
  NAND2_X1 U6450 ( .A1(n6270), .A2(n5937), .ZN(n6279) );
  NAND2_X1 U6451 ( .A1(n7848), .A2(n6777), .ZN(n7849) );
  NAND2_X1 U6452 ( .A1(n5928), .A2(n5927), .ZN(n6075) );
  NAND2_X1 U6453 ( .A1(n7179), .A2(n5926), .ZN(n6061) );
  XNOR2_X1 U6454 ( .A(n8012), .B(n7090), .ZN(n7862) );
  OR2_X1 U6455 ( .A1(n6302), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6315) );
  OAI21_X1 U6456 ( .B1(n7615), .B2(n10111), .A(n7614), .ZN(n10120) );
  INV_X1 U6457 ( .A(n10121), .ZN(n10133) );
  OR2_X1 U6458 ( .A1(n6344), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n7819) );
  AND2_X1 U6459 ( .A1(n6456), .A2(n6455), .ZN(n8349) );
  NAND2_X1 U6460 ( .A1(n6761), .A2(n6760), .ZN(n7175) );
  INV_X1 U6461 ( .A(n6825), .ZN(n8259) );
  INV_X1 U6462 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n8730) );
  NOR2_X1 U6463 ( .A1(n5795), .A2(n9040), .ZN(n5818) );
  AND2_X1 U6464 ( .A1(n5857), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9202) );
  AND2_X1 U6465 ( .A1(n5671), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5697) );
  AND2_X1 U6466 ( .A1(n9708), .A2(n9709), .ZN(n9710) );
  INV_X1 U6467 ( .A(n9205), .ZN(n9442) );
  AND2_X1 U6468 ( .A1(n9299), .A2(n9166), .ZN(n9167) );
  AND2_X1 U6469 ( .A1(n9500), .A2(n9351), .ZN(n9161) );
  AND2_X1 U6470 ( .A1(n6692), .A2(n6743), .ZN(n7279) );
  OR2_X1 U6471 ( .A1(n6743), .A2(n6692), .ZN(n6977) );
  AND2_X1 U6472 ( .A1(n5596), .A2(n5595), .ZN(n5608) );
  XNOR2_X1 U6473 ( .A(n5418), .B(SI_11_), .ZN(n5419) );
  XNOR2_X1 U6474 ( .A(n5363), .B(SI_9_), .ZN(n5366) );
  INV_X1 U6475 ( .A(n6756), .ZN(n6853) );
  NAND2_X1 U6476 ( .A1(n6491), .A2(n6490), .ZN(n6492) );
  AND3_X1 U6477 ( .A1(n5994), .A2(n5993), .A3(n5992), .ZN(n8333) );
  INV_X1 U6478 ( .A(n7121), .ZN(n7155) );
  INV_X1 U6479 ( .A(n8250), .ZN(n10143) );
  INV_X1 U6480 ( .A(n8411), .ZN(n8429) );
  INV_X1 U6481 ( .A(n8447), .ZN(n8461) );
  NAND2_X1 U6482 ( .A1(n10262), .A2(n6823), .ZN(n6824) );
  NAND2_X1 U6483 ( .A1(n10238), .A2(n6842), .ZN(n6843) );
  OR2_X1 U6484 ( .A1(n6995), .A2(n6835), .ZN(n6841) );
  INV_X1 U6485 ( .A(n6804), .ZN(n6808) );
  INV_X1 U6486 ( .A(n9056), .ZN(n9038) );
  AND4_X1 U6487 ( .A1(n5862), .A2(n5861), .A3(n5860), .A4(n5859), .ZN(n9236)
         );
  AND4_X1 U6488 ( .A1(n5578), .A2(n5577), .A3(n5576), .A4(n5575), .ZN(n9376)
         );
  INV_X1 U6489 ( .A(n9784), .ZN(n9829) );
  INV_X1 U6490 ( .A(n9187), .ZN(n9272) );
  INV_X1 U6491 ( .A(n9415), .ZN(n9877) );
  INV_X1 U6492 ( .A(n9420), .ZN(n9890) );
  AND2_X1 U6493 ( .A1(n5836), .A2(n9549), .ZN(n6979) );
  INV_X1 U6494 ( .A(n9997), .ZN(n10007) );
  AND2_X1 U6495 ( .A1(n6848), .A2(n6847), .ZN(n9546) );
  AND2_X1 U6496 ( .A1(n5432), .A2(n5460), .ZN(n9737) );
  AND2_X1 U6497 ( .A1(n5322), .A2(n5344), .ZN(n6950) );
  INV_X1 U6498 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5181) );
  AND2_X1 U6499 ( .A1(n6999), .A2(n6998), .ZN(n8050) );
  OR2_X1 U6500 ( .A1(n6511), .A2(n6510), .ZN(n6512) );
  INV_X1 U6501 ( .A(n8322), .ZN(n8076) );
  INV_X1 U6502 ( .A(n8065), .ZN(n8420) );
  OR2_X1 U6503 ( .A1(n7171), .A2(n10153), .ZN(n8411) );
  INV_X1 U6504 ( .A(n10264), .ZN(n10262) );
  INV_X1 U6505 ( .A(n8299), .ZN(n8534) );
  AND2_X1 U6506 ( .A1(n6841), .A2(n6840), .ZN(n10238) );
  AND2_X1 U6507 ( .A1(n6850), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7015) );
  INV_X1 U6508 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6897) );
  AND2_X1 U6509 ( .A1(n5900), .A2(n5899), .ZN(n5901) );
  INV_X1 U6510 ( .A(n7470), .ZN(n9965) );
  INV_X1 U6511 ( .A(n9803), .ZN(n9840) );
  OR2_X1 U6512 ( .A1(n9907), .A2(n7289), .ZN(n9415) );
  AND2_X1 U6513 ( .A1(n7237), .A2(n9893), .ZN(n9851) );
  INV_X1 U6514 ( .A(n9851), .ZN(n9238) );
  INV_X1 U6515 ( .A(n10033), .ZN(n10031) );
  INV_X1 U6516 ( .A(n10013), .ZN(n10011) );
  INV_X1 U6517 ( .A(n9917), .ZN(n9918) );
  AND2_X1 U6518 ( .A1(n9547), .A2(n9546), .ZN(n9917) );
  INV_X1 U6519 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n8687) );
  INV_X1 U6520 ( .A(n8224), .ZN(P2_U3893) );
  NOR2_X2 U6521 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5053) );
  NOR2_X1 U6522 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5057) );
  NOR2_X1 U6523 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5056) );
  NOR2_X1 U6524 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5062) );
  NOR2_X1 U6525 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5061) );
  NOR2_X1 U6526 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5060) );
  NOR2_X1 U6527 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5059) );
  NAND4_X1 U6528 ( .A1(n5062), .A2(n5061), .A3(n5060), .A4(n5059), .ZN(n5063)
         );
  INV_X1 U6529 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5068) );
  INV_X1 U6530 ( .A(n5073), .ZN(n5076) );
  NAND2_X1 U6531 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n5071) );
  NAND2_X1 U6532 ( .A1(n5096), .A2(n5071), .ZN(n5072) );
  INV_X1 U6533 ( .A(n5075), .ZN(n5074) );
  AND2_X2 U6534 ( .A1(n5076), .A2(n5074), .ZN(n5699) );
  NAND2_X1 U6535 ( .A1(n5699), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5080) );
  AND2_X2 U6536 ( .A1(n5073), .A2(n5074), .ZN(n5187) );
  NAND2_X1 U6537 ( .A1(n5187), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5079) );
  AND2_X2 U6538 ( .A1(n5076), .A2(n9557), .ZN(n5145) );
  NAND2_X1 U6539 ( .A1(n5145), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5078) );
  AND2_X2 U6540 ( .A1(n5073), .A2(n9557), .ZN(n5144) );
  NAND2_X1 U6541 ( .A1(n5144), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5077) );
  INV_X1 U6542 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8619) );
  INV_X1 U6543 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5537) );
  INV_X1 U6544 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5081) );
  NOR2_X2 U6545 ( .A1(n5492), .A2(n5045), .ZN(n5613) );
  INV_X1 U6546 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5082) );
  INV_X1 U6547 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8628) );
  NAND2_X1 U6548 ( .A1(n5084), .A2(n8628), .ZN(n5085) );
  AND2_X2 U6549 ( .A1(n5086), .A2(n5085), .ZN(n6744) );
  NAND2_X1 U6551 ( .A1(n5087), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5092) );
  INV_X1 U6552 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5091) );
  NAND2_X1 U6553 ( .A1(n5092), .A2(n5091), .ZN(n5094) );
  NAND2_X1 U6554 ( .A1(n5088), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5089) );
  MUX2_X1 U6555 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5089), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n5090) );
  OR2_X1 U6556 ( .A1(n5092), .A2(n5091), .ZN(n5093) );
  NAND2_X1 U6557 ( .A1(n9065), .A2(n5529), .ZN(n5125) );
  INV_X1 U6558 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U6559 ( .A1(n7223), .A2(n5100), .ZN(n5103) );
  NAND2_X1 U6560 ( .A1(n5104), .A2(SI_1_), .ZN(n5151) );
  AND2_X1 U6561 ( .A1(n5105), .A2(n5151), .ZN(n5107) );
  AND2_X1 U6562 ( .A1(n5106), .A2(SI_0_), .ZN(n5108) );
  INV_X1 U6563 ( .A(n5107), .ZN(n5110) );
  INV_X1 U6564 ( .A(n5108), .ZN(n5109) );
  NAND2_X1 U6565 ( .A1(n5110), .A2(n5109), .ZN(n5111) );
  NAND2_X1 U6566 ( .A1(n5152), .A2(n5111), .ZN(n6867) );
  INV_X1 U6567 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6859) );
  NAND2_X1 U6568 ( .A1(n5616), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5113) );
  NAND2_X1 U6569 ( .A1(n5114), .A2(n6969), .ZN(n5120) );
  INV_X1 U6570 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5115) );
  NAND2_X1 U6571 ( .A1(n8628), .A2(n5115), .ZN(n5116) );
  INV_X1 U6572 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5118) );
  NAND2_X4 U6573 ( .A1(n5121), .A2(n6848), .ZN(n5868) );
  INV_X1 U6574 ( .A(n5849), .ZN(n7515) );
  NAND2_X1 U6575 ( .A1(n7515), .A2(n6968), .ZN(n5122) );
  NAND2_X1 U6576 ( .A1(n5849), .A2(n6744), .ZN(n6974) );
  NAND2_X1 U6577 ( .A1(n5122), .A2(n6974), .ZN(n5123) );
  NAND2_X1 U6578 ( .A1(n7275), .A2(n5286), .ZN(n5124) );
  INV_X2 U6579 ( .A(n5868), .ZN(n5708) );
  NAND2_X1 U6580 ( .A1(n9065), .A2(n5708), .ZN(n5127) );
  NAND2_X1 U6581 ( .A1(n7275), .A2(n5136), .ZN(n5126) );
  NAND2_X1 U6582 ( .A1(n5127), .A2(n5126), .ZN(n5140) );
  NAND2_X1 U6583 ( .A1(n5699), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5131) );
  NAND2_X1 U6584 ( .A1(n5187), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5130) );
  NAND2_X1 U6585 ( .A1(n5145), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5129) );
  NAND2_X1 U6586 ( .A1(n5144), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5128) );
  NAND2_X1 U6587 ( .A1(n7274), .A2(n5136), .ZN(n5135) );
  INV_X1 U6588 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9071) );
  NAND2_X1 U6589 ( .A1(n6857), .A2(SI_0_), .ZN(n5132) );
  INV_X1 U6590 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8718) );
  XNOR2_X1 U6591 ( .A(n5132), .B(n8718), .ZN(n6855) );
  MUX2_X1 U6592 ( .A(n9071), .B(n6855), .S(n6884), .Z(n9901) );
  INV_X1 U6593 ( .A(n9901), .ZN(n5133) );
  INV_X1 U6594 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9657) );
  NAND2_X1 U6595 ( .A1(n7274), .A2(n5708), .ZN(n5139) );
  INV_X1 U6596 ( .A(n6848), .ZN(n5137) );
  NAND2_X1 U6597 ( .A1(n5137), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n5138) );
  OAI211_X1 U6598 ( .C1(n9901), .C2(n5541), .A(n5139), .B(n5138), .ZN(n6906)
         );
  AOI22_X1 U6599 ( .A1(n6907), .A2(n6906), .B1(n4522), .B2(n5866), .ZN(n6987)
         );
  NAND2_X1 U6600 ( .A1(n6988), .A2(n6987), .ZN(n6986) );
  INV_X1 U6601 ( .A(n5140), .ZN(n5141) );
  NAND2_X1 U6602 ( .A1(n5142), .A2(n5141), .ZN(n5143) );
  NAND2_X1 U6603 ( .A1(n6986), .A2(n5143), .ZN(n7020) );
  NAND2_X1 U6604 ( .A1(n5187), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5149) );
  NAND2_X1 U6605 ( .A1(n5144), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5148) );
  NAND2_X1 U6606 ( .A1(n5145), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5147) );
  NAND2_X1 U6607 ( .A1(n5699), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5146) );
  NAND4_X1 U6608 ( .A1(n5149), .A2(n5148), .A3(n5147), .A4(n5146), .ZN(n9934)
         );
  NAND2_X1 U6609 ( .A1(n9934), .A2(n5136), .ZN(n5164) );
  NAND2_X1 U6610 ( .A1(n5152), .A2(n5151), .ZN(n5157) );
  INV_X1 U6611 ( .A(n5153), .ZN(n5155) );
  INV_X1 U6612 ( .A(SI_2_), .ZN(n5154) );
  NAND2_X1 U6613 ( .A1(n5157), .A2(n5156), .ZN(n5173) );
  OR2_X1 U6614 ( .A1(n5157), .A2(n5156), .ZN(n5158) );
  NAND2_X1 U6615 ( .A1(n5173), .A2(n5158), .ZN(n6861) );
  OR2_X1 U6616 ( .A1(n5150), .A2(n6861), .ZN(n5162) );
  INV_X1 U6617 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6858) );
  OR2_X1 U6618 ( .A1(n4456), .A2(n6858), .ZN(n5161) );
  OR2_X1 U6619 ( .A1(n5159), .A2(n9550), .ZN(n5210) );
  XNOR2_X1 U6620 ( .A(n5210), .B(n5181), .ZN(n9077) );
  OR2_X1 U6621 ( .A1(n6884), .A2(n9077), .ZN(n5160) );
  XNOR2_X1 U6622 ( .A(n5165), .B(n5866), .ZN(n5170) );
  OR2_X1 U6623 ( .A1(n9930), .A2(n5541), .ZN(n5167) );
  NAND2_X1 U6624 ( .A1(n9934), .A2(n5708), .ZN(n5166) );
  NAND2_X1 U6625 ( .A1(n5167), .A2(n5166), .ZN(n5168) );
  XNOR2_X1 U6626 ( .A(n5170), .B(n5168), .ZN(n7021) );
  INV_X1 U6627 ( .A(n5168), .ZN(n5169) );
  NAND2_X1 U6628 ( .A1(n5170), .A2(n5169), .ZN(n5171) );
  NAND2_X1 U6629 ( .A1(n5173), .A2(n5172), .ZN(n5179) );
  MUX2_X1 U6630 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n6860), .Z(n5174) );
  NAND2_X1 U6631 ( .A1(n5174), .A2(SI_3_), .ZN(n5200) );
  INV_X1 U6632 ( .A(n5174), .ZN(n5176) );
  INV_X1 U6633 ( .A(SI_3_), .ZN(n5175) );
  NAND2_X1 U6634 ( .A1(n5176), .A2(n5175), .ZN(n5177) );
  NAND2_X1 U6635 ( .A1(n5179), .A2(n5178), .ZN(n5201) );
  OR2_X1 U6636 ( .A1(n5179), .A2(n5178), .ZN(n5180) );
  NAND2_X1 U6637 ( .A1(n5201), .A2(n5180), .ZN(n6863) );
  OR2_X1 U6638 ( .A1(n5150), .A2(n6863), .ZN(n5186) );
  INV_X1 U6639 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n8841) );
  OR2_X1 U6640 ( .A1(n6581), .A2(n8841), .ZN(n5185) );
  NAND2_X1 U6641 ( .A1(n5210), .A2(n5181), .ZN(n5182) );
  NAND2_X1 U6642 ( .A1(n5182), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5183) );
  XNOR2_X1 U6643 ( .A(n5183), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6935) );
  INV_X1 U6644 ( .A(n6935), .ZN(n9603) );
  OR2_X1 U6645 ( .A1(n6884), .A2(n9603), .ZN(n5184) );
  AND3_X2 U6646 ( .A1(n5186), .A2(n5185), .A3(n5184), .ZN(n7311) );
  NAND2_X1 U6647 ( .A1(n5187), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U6648 ( .A1(n5145), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5191) );
  NAND2_X1 U6649 ( .A1(n5144), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5190) );
  INV_X1 U6650 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5188) );
  NAND2_X1 U6651 ( .A1(n5699), .A2(n5188), .ZN(n5189) );
  NAND4_X1 U6652 ( .A1(n5192), .A2(n5191), .A3(n5190), .A4(n5189), .ZN(n9063)
         );
  NAND2_X1 U6653 ( .A1(n9063), .A2(n5136), .ZN(n5193) );
  XNOR2_X1 U6654 ( .A(n5194), .B(n5866), .ZN(n5199) );
  OR2_X1 U6655 ( .A1(n7311), .A2(n5541), .ZN(n5196) );
  NAND2_X1 U6656 ( .A1(n9063), .A2(n5708), .ZN(n5195) );
  NAND2_X1 U6657 ( .A1(n5196), .A2(n5195), .ZN(n5197) );
  INV_X1 U6658 ( .A(n5197), .ZN(n5198) );
  INV_X1 U6659 ( .A(n7243), .ZN(n5226) );
  NAND2_X1 U6660 ( .A1(n5201), .A2(n5200), .ZN(n5207) );
  MUX2_X1 U6661 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n6860), .Z(n5202) );
  NAND2_X1 U6662 ( .A1(n5202), .A2(SI_4_), .ZN(n5230) );
  INV_X1 U6663 ( .A(n5202), .ZN(n5204) );
  NAND2_X1 U6664 ( .A1(n5204), .A2(n5203), .ZN(n5205) );
  NAND2_X1 U6665 ( .A1(n5207), .A2(n5206), .ZN(n5231) );
  OR2_X1 U6666 ( .A1(n5207), .A2(n5206), .ZN(n5208) );
  NAND2_X1 U6667 ( .A1(n5231), .A2(n5208), .ZN(n6866) );
  OR2_X1 U6668 ( .A1(n5150), .A2(n6866), .ZN(n5215) );
  INV_X1 U6669 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6865) );
  OR2_X1 U6670 ( .A1(n6581), .A2(n6865), .ZN(n5214) );
  OAI21_X1 U6671 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(P1_IR_REG_3__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5209) );
  NAND2_X1 U6672 ( .A1(n5210), .A2(n5209), .ZN(n5212) );
  INV_X1 U6673 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5211) );
  XNOR2_X1 U6674 ( .A(n5212), .B(n5211), .ZN(n6938) );
  INV_X1 U6675 ( .A(n6938), .ZN(n9687) );
  OR2_X1 U6676 ( .A1(n6884), .A2(n9687), .ZN(n5213) );
  NAND2_X1 U6677 ( .A1(n5144), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5220) );
  NAND2_X1 U6678 ( .A1(n5885), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5219) );
  AND2_X1 U6679 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5249) );
  NOR2_X1 U6680 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5216) );
  NOR2_X1 U6681 ( .A1(n5249), .A2(n5216), .ZN(n7299) );
  NAND2_X1 U6682 ( .A1(n5699), .A2(n7299), .ZN(n5218) );
  NAND2_X1 U6683 ( .A1(n5145), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5217) );
  NAND4_X1 U6684 ( .A1(n5220), .A2(n5219), .A3(n5218), .A4(n5217), .ZN(n9863)
         );
  NAND2_X1 U6685 ( .A1(n9863), .A2(n5529), .ZN(n5221) );
  OAI21_X1 U6686 ( .B1(n9943), .B2(n5678), .A(n5221), .ZN(n5222) );
  XNOR2_X1 U6687 ( .A(n5222), .B(n4458), .ZN(n5228) );
  OR2_X1 U6688 ( .A1(n9943), .A2(n5541), .ZN(n5224) );
  NAND2_X1 U6689 ( .A1(n9863), .A2(n5708), .ZN(n5223) );
  NAND2_X1 U6690 ( .A1(n5224), .A2(n5223), .ZN(n5227) );
  XNOR2_X1 U6691 ( .A(n5228), .B(n5227), .ZN(n7244) );
  NAND2_X1 U6692 ( .A1(n5228), .A2(n5227), .ZN(n5229) );
  NAND2_X1 U6693 ( .A1(n5231), .A2(n5230), .ZN(n5237) );
  MUX2_X1 U6694 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n6857), .Z(n5232) );
  INV_X1 U6695 ( .A(n5232), .ZN(n5234) );
  INV_X1 U6696 ( .A(SI_5_), .ZN(n5233) );
  NAND2_X1 U6697 ( .A1(n5234), .A2(n5233), .ZN(n5235) );
  OR2_X1 U6698 ( .A1(n5237), .A2(n5236), .ZN(n5238) );
  NAND2_X1 U6699 ( .A1(n5274), .A2(n5238), .ZN(n6870) );
  OR2_X1 U6700 ( .A1(n5150), .A2(n6870), .ZN(n5246) );
  INV_X1 U6701 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6869) );
  OR2_X1 U6702 ( .A1(n6581), .A2(n6869), .ZN(n5245) );
  NAND2_X1 U6703 ( .A1(n5239), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5240) );
  MUX2_X1 U6704 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5240), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5243) );
  NAND2_X1 U6705 ( .A1(n5243), .A2(n5242), .ZN(n6928) );
  OR2_X1 U6706 ( .A1(n6884), .A2(n6928), .ZN(n5244) );
  NAND2_X1 U6707 ( .A1(n5885), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U6708 ( .A1(n5144), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5253) );
  NAND2_X1 U6709 ( .A1(n5249), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5264) );
  OAI21_X1 U6710 ( .B1(n5249), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5264), .ZN(
        n9868) );
  INV_X1 U6711 ( .A(n9868), .ZN(n5250) );
  NAND2_X1 U6712 ( .A1(n5886), .A2(n5250), .ZN(n5252) );
  NAND2_X1 U6713 ( .A1(n5145), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5251) );
  NAND4_X1 U6714 ( .A1(n5254), .A2(n5253), .A3(n5252), .A4(n5251), .ZN(n9062)
         );
  NAND2_X1 U6715 ( .A1(n9062), .A2(n5136), .ZN(n5255) );
  OAI21_X1 U6716 ( .B1(n9953), .B2(n5678), .A(n5255), .ZN(n5256) );
  XNOR2_X1 U6717 ( .A(n5256), .B(n4458), .ZN(n5260) );
  INV_X1 U6718 ( .A(n5260), .ZN(n5257) );
  OR2_X1 U6719 ( .A1(n9953), .A2(n5863), .ZN(n5259) );
  NAND2_X1 U6720 ( .A1(n9062), .A2(n5708), .ZN(n5258) );
  NAND2_X1 U6721 ( .A1(n5259), .A2(n5258), .ZN(n7322) );
  NAND2_X1 U6722 ( .A1(n7319), .A2(n7322), .ZN(n5262) );
  NAND2_X1 U6723 ( .A1(n6585), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5269) );
  NAND2_X1 U6724 ( .A1(n5885), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5268) );
  AND2_X1 U6725 ( .A1(n5264), .A2(n5263), .ZN(n5265) );
  NOR2_X1 U6726 ( .A1(n5300), .A2(n5265), .ZN(n7353) );
  NAND2_X1 U6727 ( .A1(n5699), .A2(n7353), .ZN(n5267) );
  NAND2_X1 U6728 ( .A1(n5145), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5266) );
  OR2_X1 U6729 ( .A1(n7424), .A2(n5868), .ZN(n5285) );
  NAND2_X1 U6730 ( .A1(n5242), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5270) );
  MUX2_X1 U6731 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5270), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5272) );
  NOR2_X1 U6732 ( .A1(n5242), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5318) );
  INV_X1 U6733 ( .A(n5318), .ZN(n5271) );
  NAND2_X1 U6734 ( .A1(n5272), .A2(n5271), .ZN(n6944) );
  MUX2_X1 U6735 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6857), .Z(n5275) );
  NAND2_X1 U6736 ( .A1(n5275), .A2(SI_6_), .ZN(n5289) );
  INV_X1 U6737 ( .A(n5275), .ZN(n5277) );
  INV_X1 U6738 ( .A(SI_6_), .ZN(n5276) );
  NAND2_X1 U6739 ( .A1(n5277), .A2(n5276), .ZN(n5278) );
  OR2_X1 U6740 ( .A1(n5280), .A2(n5279), .ZN(n5281) );
  NAND2_X1 U6741 ( .A1(n5290), .A2(n5281), .ZN(n6873) );
  OR2_X1 U6742 ( .A1(n6873), .A2(n5150), .ZN(n5283) );
  INV_X1 U6743 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6874) );
  OR2_X1 U6744 ( .A1(n6581), .A2(n6874), .ZN(n5282) );
  OAI211_X1 U6745 ( .C1(n6884), .C2(n6944), .A(n5283), .B(n5282), .ZN(n7411)
         );
  NAND2_X1 U6746 ( .A1(n7411), .A2(n5529), .ZN(n5284) );
  NAND2_X1 U6747 ( .A1(n5285), .A2(n5284), .ZN(n7345) );
  NAND2_X1 U6748 ( .A1(n7411), .A2(n5631), .ZN(n5287) );
  OAI21_X1 U6749 ( .B1(n7424), .B2(n5863), .A(n5287), .ZN(n5288) );
  XNOR2_X1 U6750 ( .A(n5288), .B(n4458), .ZN(n7344) );
  MUX2_X1 U6751 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6857), .Z(n5291) );
  INV_X1 U6752 ( .A(n5291), .ZN(n5293) );
  INV_X1 U6753 ( .A(SI_7_), .ZN(n5292) );
  NAND2_X1 U6754 ( .A1(n5293), .A2(n5292), .ZN(n5294) );
  OR2_X1 U6755 ( .A1(n5318), .A2(n9550), .ZN(n5298) );
  XNOR2_X1 U6756 ( .A(n5298), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6947) );
  AOI22_X1 U6757 ( .A1(n5619), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5618), .B2(
        n6947), .ZN(n5299) );
  NAND2_X1 U6758 ( .A1(n7456), .A2(n5631), .ZN(n5307) );
  NAND2_X1 U6759 ( .A1(n6585), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5305) );
  NAND2_X1 U6760 ( .A1(n5885), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5304) );
  NAND2_X1 U6761 ( .A1(n5300), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5326) );
  OR2_X1 U6762 ( .A1(n5300), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5301) );
  AND2_X1 U6763 ( .A1(n5326), .A2(n5301), .ZN(n7427) );
  NAND2_X1 U6764 ( .A1(n5886), .A2(n7427), .ZN(n5303) );
  NAND2_X1 U6765 ( .A1(n5145), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5302) );
  OR2_X1 U6766 ( .A1(n7552), .A2(n5863), .ZN(n5306) );
  NAND2_X1 U6767 ( .A1(n5307), .A2(n5306), .ZN(n5308) );
  XNOR2_X1 U6768 ( .A(n5308), .B(n5866), .ZN(n5311) );
  NAND2_X1 U6769 ( .A1(n7456), .A2(n5136), .ZN(n5310) );
  OR2_X1 U6770 ( .A1(n7552), .A2(n5868), .ZN(n5309) );
  AND2_X1 U6771 ( .A1(n5310), .A2(n5309), .ZN(n5312) );
  NAND2_X1 U6772 ( .A1(n5311), .A2(n5312), .ZN(n7418) );
  INV_X1 U6773 ( .A(n5311), .ZN(n5314) );
  INV_X1 U6774 ( .A(n5312), .ZN(n5313) );
  NAND2_X1 U6775 ( .A1(n5314), .A2(n5313), .ZN(n7419) );
  MUX2_X1 U6776 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n6857), .Z(n5340) );
  XNOR2_X1 U6777 ( .A(n5343), .B(n5342), .ZN(n6877) );
  NAND2_X1 U6778 ( .A1(n6877), .A2(n6583), .ZN(n5324) );
  INV_X1 U6779 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5317) );
  AND2_X1 U6780 ( .A1(n5318), .A2(n5317), .ZN(n5373) );
  OR2_X1 U6781 ( .A1(n5373), .A2(n9550), .ZN(n5321) );
  INV_X1 U6782 ( .A(n5321), .ZN(n5319) );
  NAND2_X1 U6783 ( .A1(n5319), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5322) );
  INV_X1 U6784 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5320) );
  NAND2_X1 U6785 ( .A1(n5321), .A2(n5320), .ZN(n5344) );
  AOI22_X1 U6786 ( .A1(n5619), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5618), .B2(
        n6950), .ZN(n5323) );
  NAND2_X1 U6787 ( .A1(n5324), .A2(n5323), .ZN(n7470) );
  NAND2_X1 U6788 ( .A1(n7470), .A2(n5631), .ZN(n5333) );
  NAND2_X1 U6789 ( .A1(n5885), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5331) );
  NAND2_X1 U6790 ( .A1(n5145), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5330) );
  INV_X1 U6791 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5325) );
  NAND2_X1 U6792 ( .A1(n5326), .A2(n5325), .ZN(n5327) );
  AND2_X1 U6793 ( .A1(n5348), .A2(n5327), .ZN(n7466) );
  NAND2_X1 U6794 ( .A1(n5886), .A2(n7466), .ZN(n5329) );
  NAND2_X1 U6795 ( .A1(n6585), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5328) );
  OR2_X1 U6796 ( .A1(n7647), .A2(n5863), .ZN(n5332) );
  NAND2_X1 U6797 ( .A1(n5333), .A2(n5332), .ZN(n5334) );
  XNOR2_X1 U6798 ( .A(n5334), .B(n5866), .ZN(n5336) );
  XNOR2_X2 U6799 ( .A(n5338), .B(n5336), .ZN(n7549) );
  NOR2_X1 U6800 ( .A1(n7647), .A2(n5868), .ZN(n5335) );
  AOI21_X1 U6801 ( .B1(n7470), .B2(n5136), .A(n5335), .ZN(n7548) );
  NAND2_X1 U6802 ( .A1(n7549), .A2(n7548), .ZN(n7547) );
  INV_X1 U6803 ( .A(n5336), .ZN(n5337) );
  OR2_X1 U6804 ( .A1(n5338), .A2(n5337), .ZN(n5339) );
  NAND2_X1 U6805 ( .A1(n7547), .A2(n5339), .ZN(n7644) );
  INV_X1 U6806 ( .A(n5340), .ZN(n5341) );
  INV_X1 U6807 ( .A(SI_8_), .ZN(n8772) );
  MUX2_X1 U6808 ( .A(n6897), .B(n8687), .S(n6857), .Z(n5363) );
  XNOR2_X1 U6809 ( .A(n5367), .B(n5366), .ZN(n6891) );
  NAND2_X1 U6810 ( .A1(n6891), .A2(n6583), .ZN(n5347) );
  NAND2_X1 U6811 ( .A1(n5344), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5345) );
  XNOR2_X1 U6812 ( .A(n5345), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9122) );
  AOI22_X1 U6813 ( .A1(n5619), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5618), .B2(
        n9122), .ZN(n5346) );
  NAND2_X1 U6814 ( .A1(n9972), .A2(n5631), .ZN(n5355) );
  NAND2_X1 U6815 ( .A1(n5885), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U6816 ( .A1(n5145), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5352) );
  AND2_X1 U6817 ( .A1(n5348), .A2(n8730), .ZN(n5349) );
  NOR2_X1 U6818 ( .A1(n5396), .A2(n5349), .ZN(n7648) );
  NAND2_X1 U6819 ( .A1(n5886), .A2(n7648), .ZN(n5351) );
  NAND2_X1 U6820 ( .A1(n6585), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5350) );
  OR2_X1 U6821 ( .A1(n8926), .A2(n5863), .ZN(n5354) );
  NAND2_X1 U6822 ( .A1(n5355), .A2(n5354), .ZN(n5356) );
  XNOR2_X1 U6823 ( .A(n5356), .B(n4458), .ZN(n5358) );
  NOR2_X1 U6824 ( .A1(n8926), .A2(n5868), .ZN(n5357) );
  AOI21_X1 U6825 ( .B1(n9972), .B2(n5529), .A(n5357), .ZN(n5359) );
  XNOR2_X1 U6826 ( .A(n5358), .B(n5359), .ZN(n7645) );
  NAND2_X1 U6827 ( .A1(n7644), .A2(n7645), .ZN(n5362) );
  INV_X1 U6828 ( .A(n5358), .ZN(n5360) );
  NAND2_X1 U6829 ( .A1(n5360), .A2(n5359), .ZN(n5361) );
  NAND2_X1 U6830 ( .A1(n5362), .A2(n5361), .ZN(n8921) );
  INV_X1 U6831 ( .A(n5363), .ZN(n5364) );
  MUX2_X1 U6832 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6857), .Z(n5368) );
  NAND2_X1 U6833 ( .A1(n5368), .A2(SI_10_), .ZN(n5371) );
  INV_X1 U6834 ( .A(n5368), .ZN(n5369) );
  INV_X1 U6835 ( .A(SI_10_), .ZN(n8750) );
  NAND2_X1 U6836 ( .A1(n5369), .A2(n8750), .ZN(n5370) );
  NAND2_X1 U6837 ( .A1(n5386), .A2(n5387), .ZN(n5389) );
  MUX2_X1 U6838 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6857), .Z(n5418) );
  XNOR2_X1 U6839 ( .A(n5420), .B(n5419), .ZN(n6900) );
  NAND2_X1 U6840 ( .A1(n6900), .A2(n6583), .ZN(n5377) );
  NOR2_X1 U6841 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5372) );
  AND2_X1 U6842 ( .A1(n5373), .A2(n5372), .ZN(n5390) );
  INV_X1 U6843 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U6844 ( .A1(n5390), .A2(n5374), .ZN(n5427) );
  NAND2_X1 U6845 ( .A1(n5427), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5375) );
  XNOR2_X1 U6846 ( .A(n5375), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9124) );
  AOI22_X1 U6847 ( .A1(n5619), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5618), .B2(
        n9124), .ZN(n5376) );
  NAND2_X1 U6848 ( .A1(n5885), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5382) );
  NAND2_X1 U6849 ( .A1(n6584), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5381) );
  NAND2_X1 U6850 ( .A1(n5398), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5436) );
  OR2_X1 U6851 ( .A1(n5398), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5378) );
  AND2_X1 U6852 ( .A1(n5436), .A2(n5378), .ZN(n9853) );
  NAND2_X1 U6853 ( .A1(n5886), .A2(n9853), .ZN(n5380) );
  NAND2_X1 U6854 ( .A1(n6585), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5379) );
  NAND4_X1 U6855 ( .A1(n5382), .A2(n5381), .A3(n5380), .A4(n5379), .ZN(n9995)
         );
  INV_X1 U6856 ( .A(n9995), .ZN(n7740) );
  OAI22_X1 U6857 ( .A1(n6530), .A2(n5678), .B1(n7740), .B2(n5863), .ZN(n5383)
         );
  XNOR2_X1 U6858 ( .A(n5383), .B(n4458), .ZN(n9018) );
  OR2_X1 U6859 ( .A1(n6530), .A2(n5863), .ZN(n5385) );
  NAND2_X1 U6860 ( .A1(n9995), .A2(n5708), .ZN(n5384) );
  NAND2_X1 U6861 ( .A1(n5385), .A2(n5384), .ZN(n5411) );
  NAND2_X1 U6862 ( .A1(n5389), .A2(n5388), .ZN(n6890) );
  OR2_X1 U6863 ( .A1(n6890), .A2(n5150), .ZN(n5395) );
  NOR2_X1 U6864 ( .A1(n5390), .A2(n9550), .ZN(n5391) );
  MUX2_X1 U6865 ( .A(n9550), .B(n5391), .S(P1_IR_REG_10__SCAN_IN), .Z(n5392)
         );
  INV_X1 U6866 ( .A(n5392), .ZN(n5393) );
  AOI22_X1 U6867 ( .A1(n5619), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5618), .B2(
        n9575), .ZN(n5394) );
  NAND2_X1 U6868 ( .A1(n9980), .A2(n5136), .ZN(n5404) );
  NAND2_X1 U6869 ( .A1(n5885), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5402) );
  NAND2_X1 U6870 ( .A1(n5145), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5401) );
  NOR2_X1 U6871 ( .A1(n5396), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5397) );
  OR2_X1 U6872 ( .A1(n5398), .A2(n5397), .ZN(n7492) );
  INV_X1 U6873 ( .A(n7492), .ZN(n8924) );
  NAND2_X1 U6874 ( .A1(n5699), .A2(n8924), .ZN(n5400) );
  NAND2_X1 U6875 ( .A1(n6585), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5399) );
  OR2_X1 U6876 ( .A1(n9845), .A2(n5868), .ZN(n5403) );
  NAND2_X1 U6877 ( .A1(n5404), .A2(n5403), .ZN(n8922) );
  NAND2_X1 U6878 ( .A1(n9980), .A2(n5631), .ZN(n5406) );
  OR2_X1 U6879 ( .A1(n9845), .A2(n5863), .ZN(n5405) );
  NAND2_X1 U6880 ( .A1(n5406), .A2(n5405), .ZN(n5407) );
  XNOR2_X1 U6881 ( .A(n5407), .B(n4458), .ZN(n5409) );
  AOI22_X1 U6882 ( .A1(n9018), .A2(n5411), .B1(n8922), .B2(n5409), .ZN(n5408)
         );
  NAND2_X1 U6883 ( .A1(n8921), .A2(n5408), .ZN(n5417) );
  INV_X1 U6884 ( .A(n9018), .ZN(n5415) );
  INV_X1 U6885 ( .A(n5409), .ZN(n9016) );
  INV_X1 U6886 ( .A(n8922), .ZN(n5410) );
  NAND2_X1 U6887 ( .A1(n9016), .A2(n5410), .ZN(n5412) );
  NAND2_X1 U6888 ( .A1(n5412), .A2(n5411), .ZN(n5414) );
  INV_X1 U6889 ( .A(n5411), .ZN(n9017) );
  INV_X1 U6890 ( .A(n5412), .ZN(n5413) );
  AOI22_X1 U6891 ( .A1(n5415), .A2(n5414), .B1(n9017), .B2(n5413), .ZN(n5416)
         );
  NAND2_X1 U6892 ( .A1(n5417), .A2(n5416), .ZN(n7736) );
  MUX2_X1 U6893 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6857), .Z(n5421) );
  INV_X1 U6894 ( .A(n5421), .ZN(n5422) );
  INV_X1 U6895 ( .A(SI_12_), .ZN(n8752) );
  NAND2_X1 U6896 ( .A1(n5422), .A2(n8752), .ZN(n5423) );
  NAND2_X1 U6897 ( .A1(n5451), .A2(n5423), .ZN(n5424) );
  NAND2_X1 U6898 ( .A1(n5425), .A2(n5424), .ZN(n5426) );
  NAND2_X1 U6899 ( .A1(n5426), .A2(n5452), .ZN(n6905) );
  OR2_X1 U6900 ( .A1(n5427), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5428) );
  NAND2_X1 U6901 ( .A1(n5428), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5431) );
  INV_X1 U6902 ( .A(n5431), .ZN(n5429) );
  NAND2_X1 U6903 ( .A1(n5429), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5432) );
  INV_X1 U6904 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U6905 ( .A1(n5431), .A2(n5430), .ZN(n5460) );
  AOI22_X1 U6906 ( .A1(n5619), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5618), .B2(
        n9737), .ZN(n5433) );
  NAND2_X1 U6907 ( .A1(n9998), .A2(n5631), .ZN(n5443) );
  NAND2_X1 U6908 ( .A1(n5187), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U6909 ( .A1(n6584), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5440) );
  INV_X1 U6910 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U6911 ( .A1(n5436), .A2(n5435), .ZN(n5437) );
  AND2_X1 U6912 ( .A1(n5465), .A2(n5437), .ZN(n7738) );
  NAND2_X1 U6913 ( .A1(n5699), .A2(n7738), .ZN(n5439) );
  NAND2_X1 U6914 ( .A1(n6585), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5438) );
  OR2_X1 U6915 ( .A1(n9844), .A2(n5863), .ZN(n5442) );
  NAND2_X1 U6916 ( .A1(n5443), .A2(n5442), .ZN(n5444) );
  XNOR2_X1 U6917 ( .A(n5444), .B(n4458), .ZN(n5446) );
  NOR2_X1 U6918 ( .A1(n9844), .A2(n5868), .ZN(n5445) );
  AOI21_X1 U6919 ( .B1(n9998), .B2(n5529), .A(n5445), .ZN(n5447) );
  XNOR2_X1 U6920 ( .A(n5446), .B(n5447), .ZN(n7737) );
  NAND2_X1 U6921 ( .A1(n7736), .A2(n7737), .ZN(n5450) );
  INV_X1 U6922 ( .A(n5446), .ZN(n5448) );
  NAND2_X1 U6923 ( .A1(n5448), .A2(n5447), .ZN(n5449) );
  NAND2_X1 U6924 ( .A1(n5450), .A2(n5449), .ZN(n8996) );
  MUX2_X1 U6925 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6857), .Z(n5453) );
  NAND2_X1 U6926 ( .A1(n5453), .A2(SI_13_), .ZN(n5480) );
  INV_X1 U6927 ( .A(n5453), .ZN(n5455) );
  INV_X1 U6928 ( .A(SI_13_), .ZN(n5454) );
  NAND2_X1 U6929 ( .A1(n5455), .A2(n5454), .ZN(n5456) );
  OR2_X1 U6930 ( .A1(n5458), .A2(n5457), .ZN(n5459) );
  NAND2_X1 U6931 ( .A1(n5481), .A2(n5459), .ZN(n6984) );
  NAND2_X1 U6932 ( .A1(n5460), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5461) );
  XNOR2_X1 U6933 ( .A(n5461), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9753) );
  AOI22_X1 U6934 ( .A1(n5619), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5618), .B2(
        n9753), .ZN(n5462) );
  NAND2_X1 U6935 ( .A1(n9001), .A2(n5631), .ZN(n5472) );
  NAND2_X1 U6936 ( .A1(n6585), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U6937 ( .A1(n5885), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5469) );
  INV_X1 U6938 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U6939 ( .A1(n5465), .A2(n5464), .ZN(n5466) );
  AND2_X1 U6940 ( .A1(n5497), .A2(n5466), .ZN(n8998) );
  NAND2_X1 U6941 ( .A1(n5886), .A2(n8998), .ZN(n5468) );
  NAND2_X1 U6942 ( .A1(n6584), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5467) );
  OR2_X1 U6943 ( .A1(n8909), .A2(n5863), .ZN(n5471) );
  NAND2_X1 U6944 ( .A1(n5472), .A2(n5471), .ZN(n5473) );
  XNOR2_X1 U6945 ( .A(n5473), .B(n4458), .ZN(n5475) );
  NOR2_X1 U6946 ( .A1(n8909), .A2(n5868), .ZN(n5474) );
  AOI21_X1 U6947 ( .B1(n9001), .B2(n5136), .A(n5474), .ZN(n5476) );
  XNOR2_X1 U6948 ( .A(n5475), .B(n5476), .ZN(n8997) );
  NAND2_X1 U6949 ( .A1(n8996), .A2(n8997), .ZN(n5479) );
  INV_X1 U6950 ( .A(n5475), .ZN(n5477) );
  NAND2_X1 U6951 ( .A1(n5477), .A2(n5476), .ZN(n5478) );
  NAND2_X1 U6952 ( .A1(n5481), .A2(n5480), .ZN(n5487) );
  MUX2_X1 U6953 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6857), .Z(n5482) );
  NAND2_X1 U6954 ( .A1(n5482), .A2(SI_14_), .ZN(n5510) );
  INV_X1 U6955 ( .A(n5482), .ZN(n5484) );
  INV_X1 U6956 ( .A(SI_14_), .ZN(n5483) );
  NAND2_X1 U6957 ( .A1(n5484), .A2(n5483), .ZN(n5485) );
  NAND2_X1 U6958 ( .A1(n5487), .A2(n5486), .ZN(n5511) );
  OR2_X1 U6959 ( .A1(n5487), .A2(n5486), .ZN(n5488) );
  NAND2_X1 U6960 ( .A1(n5511), .A2(n5488), .ZN(n7019) );
  NOR2_X1 U6961 ( .A1(n5489), .A2(n9550), .ZN(n5490) );
  MUX2_X1 U6962 ( .A(n9550), .B(n5490), .S(P1_IR_REG_14__SCAN_IN), .Z(n5491)
         );
  INV_X1 U6963 ( .A(n5491), .ZN(n5493) );
  AND2_X1 U6964 ( .A1(n5493), .A2(n5536), .ZN(n9126) );
  AOI22_X1 U6965 ( .A1(n5619), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5618), .B2(
        n9126), .ZN(n5494) );
  NAND2_X1 U6966 ( .A1(n9524), .A2(n5631), .ZN(n5503) );
  NAND2_X1 U6967 ( .A1(n5885), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5501) );
  NAND2_X1 U6968 ( .A1(n6585), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5500) );
  INV_X1 U6969 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5496) );
  NOR2_X1 U6970 ( .A1(n5542), .A2(n5047), .ZN(n8907) );
  NAND2_X1 U6971 ( .A1(n5699), .A2(n8907), .ZN(n5499) );
  NAND2_X1 U6972 ( .A1(n6584), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5498) );
  OR2_X1 U6973 ( .A1(n9422), .A2(n5863), .ZN(n5502) );
  NAND2_X1 U6974 ( .A1(n5503), .A2(n5502), .ZN(n5504) );
  XNOR2_X1 U6975 ( .A(n5504), .B(n4458), .ZN(n5506) );
  NOR2_X1 U6976 ( .A1(n9422), .A2(n5868), .ZN(n5505) );
  AOI21_X1 U6977 ( .B1(n9524), .B2(n5136), .A(n5505), .ZN(n8905) );
  INV_X1 U6978 ( .A(n5506), .ZN(n5507) );
  NAND2_X1 U6979 ( .A1(n5508), .A2(n5507), .ZN(n5509) );
  MUX2_X1 U6980 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6857), .Z(n5512) );
  NAND2_X1 U6981 ( .A1(n5512), .A2(SI_15_), .ZN(n5516) );
  INV_X1 U6982 ( .A(n5512), .ZN(n5514) );
  INV_X1 U6983 ( .A(SI_15_), .ZN(n5513) );
  NAND2_X1 U6984 ( .A1(n5514), .A2(n5513), .ZN(n5515) );
  MUX2_X1 U6985 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n6857), .Z(n5559) );
  XNOR2_X1 U6986 ( .A(n5559), .B(SI_16_), .ZN(n5562) );
  XNOR2_X1 U6987 ( .A(n5563), .B(n5562), .ZN(n7125) );
  NAND2_X1 U6988 ( .A1(n7125), .A2(n6583), .ZN(n5521) );
  OR2_X1 U6989 ( .A1(n5536), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n5517) );
  NAND2_X1 U6990 ( .A1(n5517), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5518) );
  OR2_X1 U6991 ( .A1(n5518), .A2(n8619), .ZN(n5519) );
  NAND2_X1 U6992 ( .A1(n5518), .A2(n8619), .ZN(n5566) );
  AND2_X1 U6993 ( .A1(n5519), .A2(n5566), .ZN(n9807) );
  AOI22_X1 U6994 ( .A1(n5619), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5618), .B2(
        n9807), .ZN(n5520) );
  NAND2_X1 U6995 ( .A1(n9520), .A2(n5631), .ZN(n5527) );
  NAND2_X1 U6996 ( .A1(n5542), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5573) );
  XNOR2_X1 U6997 ( .A(n5573), .B(P1_REG3_REG_16__SCAN_IN), .ZN(n9403) );
  NAND2_X1 U6998 ( .A1(n5886), .A2(n9403), .ZN(n5525) );
  NAND2_X1 U6999 ( .A1(n5187), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U7000 ( .A1(n6584), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5523) );
  NAND2_X1 U7001 ( .A1(n6585), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5522) );
  OR2_X1 U7002 ( .A1(n9421), .A2(n5863), .ZN(n5526) );
  NAND2_X1 U7003 ( .A1(n5527), .A2(n5526), .ZN(n5528) );
  XNOR2_X1 U7004 ( .A(n5528), .B(n4458), .ZN(n8961) );
  NAND2_X1 U7005 ( .A1(n9520), .A2(n5136), .ZN(n5531) );
  OR2_X1 U7006 ( .A1(n9421), .A2(n5868), .ZN(n5530) );
  NAND2_X1 U7007 ( .A1(n5531), .A2(n5530), .ZN(n8960) );
  OR2_X1 U7008 ( .A1(n5533), .A2(n5532), .ZN(n5534) );
  NAND2_X1 U7009 ( .A1(n5535), .A2(n5534), .ZN(n7088) );
  NAND2_X1 U7010 ( .A1(n5536), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5538) );
  XNOR2_X1 U7011 ( .A(n5538), .B(n5537), .ZN(n9128) );
  INV_X1 U7012 ( .A(n9128), .ZN(n9793) );
  AOI22_X1 U7013 ( .A1(n5619), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5618), .B2(
        n9793), .ZN(n5539) );
  NAND2_X2 U7014 ( .A1(n5540), .A2(n5539), .ZN(n9426) );
  NAND2_X1 U7015 ( .A1(n9426), .A2(n5529), .ZN(n5549) );
  NAND2_X1 U7016 ( .A1(n5885), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5547) );
  NAND2_X1 U7017 ( .A1(n5145), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5546) );
  OR2_X1 U7018 ( .A1(n5542), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5543) );
  AND2_X1 U7019 ( .A1(n5543), .A2(n5573), .ZN(n9423) );
  NAND2_X1 U7020 ( .A1(n5886), .A2(n9423), .ZN(n5545) );
  NAND2_X1 U7021 ( .A1(n6585), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5544) );
  OR2_X1 U7022 ( .A1(n9152), .A2(n5868), .ZN(n5548) );
  NAND2_X1 U7023 ( .A1(n5549), .A2(n5548), .ZN(n9048) );
  NAND2_X1 U7024 ( .A1(n9426), .A2(n5631), .ZN(n5551) );
  OR2_X1 U7025 ( .A1(n9152), .A2(n5863), .ZN(n5550) );
  NAND2_X1 U7026 ( .A1(n5551), .A2(n5550), .ZN(n5552) );
  XNOR2_X1 U7027 ( .A(n5552), .B(n4458), .ZN(n8957) );
  OAI22_X1 U7028 ( .A1(n8961), .A2(n8960), .B1(n9048), .B2(n8957), .ZN(n5553)
         );
  NAND2_X1 U7029 ( .A1(n8957), .A2(n9048), .ZN(n5555) );
  INV_X1 U7030 ( .A(n8960), .ZN(n5554) );
  NAND2_X1 U7031 ( .A1(n5555), .A2(n5554), .ZN(n5557) );
  INV_X1 U7032 ( .A(n5555), .ZN(n5556) );
  AOI22_X1 U7033 ( .A1(n8961), .A2(n5557), .B1(n5556), .B2(n8960), .ZN(n5558)
         );
  INV_X1 U7034 ( .A(n5559), .ZN(n5561) );
  INV_X1 U7035 ( .A(SI_16_), .ZN(n5560) );
  INV_X1 U7036 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n5565) );
  INV_X1 U7037 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5564) );
  MUX2_X1 U7038 ( .A(n5565), .B(n5564), .S(n6857), .Z(n5588) );
  XNOR2_X1 U7039 ( .A(n5588), .B(SI_17_), .ZN(n5590) );
  XNOR2_X1 U7040 ( .A(n5591), .B(n5590), .ZN(n7192) );
  NAND2_X1 U7041 ( .A1(n7192), .A2(n6583), .ZN(n5569) );
  NAND2_X1 U7042 ( .A1(n5566), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5567) );
  XNOR2_X1 U7043 ( .A(n5567), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9819) );
  AOI22_X1 U7044 ( .A1(n5619), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5618), .B2(
        n9819), .ZN(n5568) );
  NAND2_X1 U7045 ( .A1(n9385), .A2(n5631), .ZN(n5580) );
  NAND2_X1 U7046 ( .A1(n5885), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U7047 ( .A1(n6585), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5577) );
  INV_X1 U7048 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5571) );
  INV_X1 U7049 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5570) );
  OAI21_X1 U7050 ( .B1(n5573), .B2(n5571), .A(n5570), .ZN(n5574) );
  NAND2_X1 U7051 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_REG3_REG_16__SCAN_IN), 
        .ZN(n5572) );
  AND2_X1 U7052 ( .A1(n5574), .A2(n5622), .ZN(n9392) );
  NAND2_X1 U7053 ( .A1(n5886), .A2(n9392), .ZN(n5576) );
  NAND2_X1 U7054 ( .A1(n6584), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5575) );
  OR2_X1 U7055 ( .A1(n9376), .A2(n5863), .ZN(n5579) );
  NAND2_X1 U7056 ( .A1(n5580), .A2(n5579), .ZN(n5581) );
  XNOR2_X1 U7057 ( .A(n5581), .B(n4458), .ZN(n5584) );
  NAND2_X1 U7058 ( .A1(n9385), .A2(n5529), .ZN(n5583) );
  OR2_X1 U7059 ( .A1(n9376), .A2(n5868), .ZN(n5582) );
  NAND2_X1 U7060 ( .A1(n5583), .A2(n5582), .ZN(n5585) );
  AND2_X1 U7061 ( .A1(n5584), .A2(n5585), .ZN(n8970) );
  INV_X1 U7062 ( .A(n5584), .ZN(n5587) );
  INV_X1 U7063 ( .A(n5585), .ZN(n5586) );
  NAND2_X1 U7064 ( .A1(n5587), .A2(n5586), .ZN(n8969) );
  INV_X1 U7065 ( .A(n5588), .ZN(n5589) );
  MUX2_X1 U7066 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6857), .Z(n5592) );
  NAND2_X1 U7067 ( .A1(n5592), .A2(SI_18_), .ZN(n5596) );
  INV_X1 U7068 ( .A(n5592), .ZN(n5594) );
  INV_X1 U7069 ( .A(SI_18_), .ZN(n5593) );
  NAND2_X1 U7070 ( .A1(n5594), .A2(n5593), .ZN(n5595) );
  NAND2_X1 U7071 ( .A1(n5607), .A2(n5608), .ZN(n5612) );
  NAND2_X1 U7072 ( .A1(n5612), .A2(n5596), .ZN(n5646) );
  MUX2_X1 U7073 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n6857), .Z(n5641) );
  XNOR2_X1 U7074 ( .A(n5641), .B(SI_19_), .ZN(n5645) );
  XNOR2_X1 U7075 ( .A(n5646), .B(n5645), .ZN(n7356) );
  NAND2_X1 U7076 ( .A1(n7356), .A2(n6583), .ZN(n5598) );
  AOI22_X1 U7077 ( .A1(n5619), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n4722), .B2(
        n5618), .ZN(n5597) );
  NAND2_X1 U7078 ( .A1(n9507), .A2(n5631), .ZN(n5603) );
  INV_X1 U7079 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8722) );
  NOR2_X1 U7080 ( .A1(n5623), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5599) );
  OR2_X1 U7081 ( .A1(n5649), .A2(n5599), .ZN(n9355) );
  AOI22_X1 U7082 ( .A1(n5885), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n5144), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n5601) );
  NAND2_X1 U7083 ( .A1(n6584), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5600) );
  OAI211_X1 U7084 ( .C1(n9355), .C2(n5248), .A(n5601), .B(n5600), .ZN(n9369)
         );
  NAND2_X1 U7085 ( .A1(n9369), .A2(n5529), .ZN(n5602) );
  NAND2_X1 U7086 ( .A1(n5603), .A2(n5602), .ZN(n5604) );
  XNOR2_X1 U7087 ( .A(n5604), .B(n4458), .ZN(n8934) );
  NAND2_X1 U7088 ( .A1(n9507), .A2(n5529), .ZN(n5606) );
  NAND2_X1 U7089 ( .A1(n9369), .A2(n5708), .ZN(n5605) );
  NAND2_X1 U7090 ( .A1(n5606), .A2(n5605), .ZN(n5636) );
  INV_X1 U7091 ( .A(n5607), .ZN(n5610) );
  INV_X1 U7092 ( .A(n5608), .ZN(n5609) );
  NAND2_X1 U7093 ( .A1(n5610), .A2(n5609), .ZN(n5611) );
  NAND2_X1 U7094 ( .A1(n5612), .A2(n5611), .ZN(n7252) );
  OR2_X1 U7095 ( .A1(n7252), .A2(n5150), .ZN(n5621) );
  INV_X1 U7096 ( .A(n5613), .ZN(n5614) );
  NAND2_X1 U7097 ( .A1(n5614), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5615) );
  MUX2_X1 U7098 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5615), .S(
        P1_IR_REG_18__SCAN_IN), .Z(n5617) );
  NAND2_X1 U7099 ( .A1(n5617), .A2(n5616), .ZN(n9834) );
  INV_X1 U7100 ( .A(n9834), .ZN(n9114) );
  AOI22_X1 U7101 ( .A1(n5619), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5618), .B2(
        n9114), .ZN(n5620) );
  NAND2_X1 U7102 ( .A1(n9514), .A2(n5529), .ZN(n5630) );
  AND2_X1 U7103 ( .A1(n5622), .A2(n8722), .ZN(n5624) );
  OR2_X1 U7104 ( .A1(n5624), .A2(n5623), .ZN(n9373) );
  NAND2_X1 U7105 ( .A1(n6585), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U7106 ( .A1(n5885), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5625) );
  AND2_X1 U7107 ( .A1(n5626), .A2(n5625), .ZN(n5628) );
  NAND2_X1 U7108 ( .A1(n6584), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5627) );
  OAI211_X1 U7109 ( .C1(n9373), .C2(n5248), .A(n5628), .B(n5627), .ZN(n9506)
         );
  NAND2_X1 U7110 ( .A1(n9506), .A2(n5708), .ZN(n5629) );
  NAND2_X1 U7111 ( .A1(n5630), .A2(n5629), .ZN(n9027) );
  NAND2_X1 U7112 ( .A1(n9514), .A2(n5631), .ZN(n5633) );
  NAND2_X1 U7113 ( .A1(n9506), .A2(n5136), .ZN(n5632) );
  NAND2_X1 U7114 ( .A1(n5633), .A2(n5632), .ZN(n5634) );
  XNOR2_X1 U7115 ( .A(n5634), .B(n4458), .ZN(n8930) );
  OAI22_X1 U7116 ( .A1(n8934), .A2(n5636), .B1(n9027), .B2(n8930), .ZN(n5640)
         );
  NAND2_X1 U7117 ( .A1(n8930), .A2(n9027), .ZN(n5635) );
  INV_X1 U7118 ( .A(n5636), .ZN(n8933) );
  NAND2_X1 U7119 ( .A1(n5635), .A2(n8933), .ZN(n5638) );
  INV_X1 U7120 ( .A(n5635), .ZN(n5637) );
  AOI22_X1 U7121 ( .A1(n8934), .A2(n5638), .B1(n5637), .B2(n5636), .ZN(n5639)
         );
  INV_X1 U7122 ( .A(n5641), .ZN(n5643) );
  INV_X1 U7123 ( .A(SI_19_), .ZN(n5642) );
  NAND2_X1 U7124 ( .A1(n5643), .A2(n5642), .ZN(n5644) );
  INV_X1 U7125 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8625) );
  INV_X1 U7126 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8776) );
  MUX2_X1 U7127 ( .A(n8625), .B(n8776), .S(n6857), .Z(n5665) );
  XNOR2_X1 U7128 ( .A(n5665), .B(SI_20_), .ZN(n5662) );
  XNOR2_X1 U7129 ( .A(n5663), .B(n5662), .ZN(n7430) );
  NAND2_X1 U7130 ( .A1(n7430), .A2(n6583), .ZN(n5648) );
  OR2_X1 U7131 ( .A1(n6581), .A2(n8776), .ZN(n5647) );
  NAND2_X1 U7132 ( .A1(n9500), .A2(n5631), .ZN(n5654) );
  NOR2_X1 U7133 ( .A1(n5649), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5650) );
  OR2_X1 U7134 ( .A1(n5671), .A2(n5650), .ZN(n9336) );
  AOI22_X1 U7135 ( .A1(n5885), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n5144), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n5652) );
  NAND2_X1 U7136 ( .A1(n6584), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5651) );
  OAI211_X1 U7137 ( .C1(n9336), .C2(n5248), .A(n5652), .B(n5651), .ZN(n9351)
         );
  NAND2_X1 U7138 ( .A1(n9351), .A2(n5529), .ZN(n5653) );
  NAND2_X1 U7139 ( .A1(n5654), .A2(n5653), .ZN(n5655) );
  XNOR2_X1 U7140 ( .A(n5655), .B(n5866), .ZN(n8989) );
  AND2_X1 U7141 ( .A1(n9351), .A2(n5708), .ZN(n5656) );
  AOI21_X1 U7142 ( .B1(n9500), .B2(n5529), .A(n5656), .ZN(n5658) );
  NAND2_X1 U7143 ( .A1(n8989), .A2(n5658), .ZN(n5657) );
  NAND2_X1 U7144 ( .A1(n8987), .A2(n5657), .ZN(n5661) );
  INV_X1 U7145 ( .A(n8989), .ZN(n5659) );
  INV_X1 U7146 ( .A(n5658), .ZN(n8988) );
  NAND2_X1 U7147 ( .A1(n5659), .A2(n8988), .ZN(n5660) );
  NAND2_X1 U7148 ( .A1(n5663), .A2(n5662), .ZN(n5667) );
  INV_X1 U7149 ( .A(SI_20_), .ZN(n5664) );
  NAND2_X1 U7150 ( .A1(n5665), .A2(n5664), .ZN(n5666) );
  NAND2_X1 U7151 ( .A1(n5667), .A2(n5666), .ZN(n5688) );
  INV_X1 U7152 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7514) );
  INV_X1 U7153 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7517) );
  MUX2_X1 U7154 ( .A(n7514), .B(n7517), .S(n6857), .Z(n5689) );
  XNOR2_X1 U7155 ( .A(n5689), .B(SI_21_), .ZN(n5668) );
  XNOR2_X1 U7156 ( .A(n5688), .B(n5668), .ZN(n7513) );
  NAND2_X1 U7157 ( .A1(n7513), .A2(n6583), .ZN(n5670) );
  OR2_X1 U7158 ( .A1(n6581), .A2(n7517), .ZN(n5669) );
  NOR2_X1 U7159 ( .A1(n5671), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5672) );
  OR2_X1 U7160 ( .A1(n5697), .A2(n5672), .ZN(n9327) );
  INV_X1 U7161 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5675) );
  NAND2_X1 U7162 ( .A1(n6585), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5674) );
  NAND2_X1 U7163 ( .A1(n6584), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5673) );
  OAI211_X1 U7164 ( .C1(n5247), .C2(n5675), .A(n5674), .B(n5673), .ZN(n5676)
         );
  INV_X1 U7165 ( .A(n5676), .ZN(n5677) );
  OAI21_X1 U7166 ( .B1(n9327), .B2(n5248), .A(n5677), .ZN(n9342) );
  INV_X1 U7167 ( .A(n9342), .ZN(n9488) );
  OAI22_X1 U7168 ( .A1(n9331), .A2(n5678), .B1(n9488), .B2(n5863), .ZN(n5679)
         );
  XNOR2_X1 U7169 ( .A(n5679), .B(n4458), .ZN(n5682) );
  OR2_X1 U7170 ( .A1(n9331), .A2(n5863), .ZN(n5681) );
  NAND2_X1 U7171 ( .A1(n9342), .A2(n5708), .ZN(n5680) );
  NAND2_X1 U7172 ( .A1(n5681), .A2(n5680), .ZN(n5683) );
  XNOR2_X1 U7173 ( .A(n5682), .B(n5683), .ZN(n8942) );
  INV_X1 U7174 ( .A(n5682), .ZN(n5685) );
  INV_X1 U7175 ( .A(n5683), .ZN(n5684) );
  NAND2_X1 U7176 ( .A1(n5685), .A2(n5684), .ZN(n5686) );
  INV_X1 U7177 ( .A(SI_21_), .ZN(n5687) );
  INV_X1 U7178 ( .A(n5689), .ZN(n5690) );
  NAND2_X1 U7179 ( .A1(n5690), .A2(SI_21_), .ZN(n5691) );
  INV_X1 U7180 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7543) );
  INV_X1 U7181 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7546) );
  MUX2_X1 U7182 ( .A(n7543), .B(n7546), .S(n6857), .Z(n5692) );
  NAND2_X1 U7183 ( .A1(n5692), .A2(n8749), .ZN(n5711) );
  INV_X1 U7184 ( .A(n5692), .ZN(n5693) );
  NAND2_X1 U7185 ( .A1(n5693), .A2(SI_22_), .ZN(n5694) );
  NAND2_X1 U7186 ( .A1(n5711), .A2(n5694), .ZN(n5712) );
  XNOR2_X1 U7187 ( .A(n5713), .B(n5712), .ZN(n7541) );
  NAND2_X1 U7188 ( .A1(n7541), .A2(n6583), .ZN(n5696) );
  OR2_X1 U7189 ( .A1(n6581), .A2(n7546), .ZN(n5695) );
  NAND2_X1 U7190 ( .A1(n9304), .A2(n5631), .ZN(n5706) );
  OR2_X1 U7191 ( .A1(n5697), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5698) );
  NAND2_X1 U7192 ( .A1(n5697), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5721) );
  AND2_X1 U7193 ( .A1(n5698), .A2(n5721), .ZN(n9305) );
  NAND2_X1 U7194 ( .A1(n9305), .A2(n5699), .ZN(n5704) );
  INV_X1 U7195 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n8720) );
  NAND2_X1 U7196 ( .A1(n6585), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5701) );
  NAND2_X1 U7197 ( .A1(n6584), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5700) );
  OAI211_X1 U7198 ( .C1(n5247), .C2(n8720), .A(n5701), .B(n5700), .ZN(n5702)
         );
  INV_X1 U7199 ( .A(n5702), .ZN(n5703) );
  INV_X1 U7200 ( .A(n9481), .ZN(n9163) );
  NAND2_X1 U7201 ( .A1(n9163), .A2(n5136), .ZN(n5705) );
  NAND2_X1 U7202 ( .A1(n5706), .A2(n5705), .ZN(n5707) );
  NAND2_X1 U7203 ( .A1(n9304), .A2(n5529), .ZN(n5710) );
  NAND2_X1 U7204 ( .A1(n9163), .A2(n5708), .ZN(n5709) );
  NAND2_X1 U7205 ( .A1(n5710), .A2(n5709), .ZN(n9005) );
  INV_X1 U7206 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5714) );
  INV_X1 U7207 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7659) );
  MUX2_X1 U7208 ( .A(n5714), .B(n7659), .S(n6857), .Z(n5716) );
  INV_X1 U7209 ( .A(SI_23_), .ZN(n5715) );
  NAND2_X1 U7210 ( .A1(n5716), .A2(n5715), .ZN(n5737) );
  INV_X1 U7211 ( .A(n5716), .ZN(n5717) );
  NAND2_X1 U7212 ( .A1(n5717), .A2(SI_23_), .ZN(n5718) );
  NAND2_X1 U7213 ( .A1(n7656), .A2(n6583), .ZN(n5720) );
  OR2_X1 U7214 ( .A1(n6581), .A2(n7659), .ZN(n5719) );
  NAND2_X1 U7215 ( .A1(n9299), .A2(n5631), .ZN(n5729) );
  NAND2_X1 U7216 ( .A1(n6585), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5727) );
  NAND2_X1 U7217 ( .A1(n5885), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5726) );
  INV_X1 U7218 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8779) );
  NAND2_X1 U7219 ( .A1(n8779), .A2(n5721), .ZN(n5723) );
  INV_X1 U7220 ( .A(n5721), .ZN(n5722) );
  INV_X1 U7221 ( .A(n5745), .ZN(n5747) );
  AND2_X1 U7222 ( .A1(n5723), .A2(n5747), .ZN(n9293) );
  NAND2_X1 U7223 ( .A1(n5886), .A2(n9293), .ZN(n5725) );
  NAND2_X1 U7224 ( .A1(n6584), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5724) );
  OR2_X1 U7225 ( .A1(n9315), .A2(n5863), .ZN(n5728) );
  NAND2_X1 U7226 ( .A1(n5729), .A2(n5728), .ZN(n5730) );
  XNOR2_X1 U7227 ( .A(n5730), .B(n5866), .ZN(n5733) );
  NOR2_X1 U7228 ( .A1(n9315), .A2(n5868), .ZN(n5731) );
  AOI21_X1 U7229 ( .B1(n9299), .B2(n5136), .A(n5731), .ZN(n5732) );
  NAND2_X1 U7230 ( .A1(n5733), .A2(n5732), .ZN(n8979) );
  OR2_X1 U7231 ( .A1(n5733), .A2(n5732), .ZN(n5734) );
  AND2_X1 U7232 ( .A1(n8979), .A2(n5734), .ZN(n8914) );
  NAND2_X1 U7233 ( .A1(n5738), .A2(n5737), .ZN(n5763) );
  INV_X1 U7234 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8647) );
  INV_X1 U7235 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7724) );
  MUX2_X1 U7236 ( .A(n8647), .B(n7724), .S(n6857), .Z(n5740) );
  INV_X1 U7237 ( .A(SI_24_), .ZN(n5739) );
  NAND2_X1 U7238 ( .A1(n5740), .A2(n5739), .ZN(n5764) );
  INV_X1 U7239 ( .A(n5740), .ZN(n5741) );
  NAND2_X1 U7240 ( .A1(n5741), .A2(SI_24_), .ZN(n5742) );
  AND2_X1 U7241 ( .A1(n5764), .A2(n5742), .ZN(n5762) );
  NAND2_X1 U7242 ( .A1(n7723), .A2(n6583), .ZN(n5744) );
  OR2_X1 U7243 ( .A1(n6581), .A2(n7724), .ZN(n5743) );
  NAND2_X1 U7244 ( .A1(n9478), .A2(n5631), .ZN(n5754) );
  NAND2_X1 U7245 ( .A1(n6585), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5752) );
  NAND2_X1 U7246 ( .A1(n5187), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5751) );
  INV_X1 U7247 ( .A(n5773), .ZN(n5772) );
  INV_X1 U7248 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5746) );
  NAND2_X1 U7249 ( .A1(n5747), .A2(n5746), .ZN(n5748) );
  AND2_X1 U7250 ( .A1(n5772), .A2(n5748), .ZN(n9278) );
  NAND2_X1 U7251 ( .A1(n5886), .A2(n9278), .ZN(n5750) );
  NAND2_X1 U7252 ( .A1(n6584), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5749) );
  OR2_X1 U7253 ( .A1(n9469), .A2(n5863), .ZN(n5753) );
  NAND2_X1 U7254 ( .A1(n5754), .A2(n5753), .ZN(n5755) );
  XNOR2_X1 U7255 ( .A(n5755), .B(n5866), .ZN(n5758) );
  NOR2_X1 U7256 ( .A1(n9469), .A2(n5868), .ZN(n5756) );
  AOI21_X1 U7257 ( .B1(n9478), .B2(n5136), .A(n5756), .ZN(n5757) );
  NAND2_X1 U7258 ( .A1(n5758), .A2(n5757), .ZN(n5760) );
  OR2_X1 U7259 ( .A1(n5758), .A2(n5757), .ZN(n5759) );
  NAND2_X1 U7260 ( .A1(n5760), .A2(n5759), .ZN(n8978) );
  INV_X1 U7261 ( .A(n5760), .ZN(n5761) );
  NAND2_X1 U7262 ( .A1(n5763), .A2(n5762), .ZN(n5765) );
  INV_X1 U7263 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7756) );
  INV_X1 U7264 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7779) );
  MUX2_X1 U7265 ( .A(n7756), .B(n7779), .S(n6857), .Z(n5767) );
  INV_X1 U7266 ( .A(SI_25_), .ZN(n5766) );
  NAND2_X1 U7267 ( .A1(n5767), .A2(n5766), .ZN(n5787) );
  INV_X1 U7268 ( .A(n5767), .ZN(n5768) );
  NAND2_X1 U7269 ( .A1(n5768), .A2(SI_25_), .ZN(n5769) );
  AND2_X1 U7270 ( .A1(n5787), .A2(n5769), .ZN(n5785) );
  NAND2_X1 U7271 ( .A1(n7755), .A2(n6583), .ZN(n5771) );
  OR2_X1 U7272 ( .A1(n6581), .A2(n7779), .ZN(n5770) );
  NAND2_X1 U7273 ( .A1(n9259), .A2(n5631), .ZN(n5780) );
  NAND2_X1 U7274 ( .A1(n5187), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5778) );
  NAND2_X1 U7275 ( .A1(n6585), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5777) );
  INV_X1 U7276 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8951) );
  NAND2_X1 U7277 ( .A1(n5772), .A2(n8951), .ZN(n5774) );
  NAND2_X1 U7278 ( .A1(n5773), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5795) );
  AND2_X1 U7279 ( .A1(n5774), .A2(n5795), .ZN(n9260) );
  NAND2_X1 U7280 ( .A1(n5886), .A2(n9260), .ZN(n5776) );
  NAND2_X1 U7281 ( .A1(n6584), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5775) );
  OR2_X1 U7282 ( .A1(n9462), .A2(n5863), .ZN(n5779) );
  NAND2_X1 U7283 ( .A1(n5780), .A2(n5779), .ZN(n5782) );
  XNOR2_X1 U7284 ( .A(n5782), .B(n4458), .ZN(n5784) );
  INV_X1 U7285 ( .A(n9259), .ZN(n9470) );
  OAI22_X1 U7286 ( .A1(n9470), .A2(n5863), .B1(n9462), .B2(n5868), .ZN(n5783)
         );
  XNOR2_X1 U7287 ( .A(n5784), .B(n5783), .ZN(n8949) );
  NOR2_X1 U7288 ( .A1(n5784), .A2(n5783), .ZN(n9036) );
  INV_X1 U7289 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8889) );
  INV_X1 U7290 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9563) );
  MUX2_X1 U7291 ( .A(n8889), .B(n9563), .S(n6857), .Z(n5790) );
  INV_X1 U7292 ( .A(SI_26_), .ZN(n5789) );
  NAND2_X1 U7293 ( .A1(n5790), .A2(n5789), .ZN(n5810) );
  INV_X1 U7294 ( .A(n5790), .ZN(n5791) );
  NAND2_X1 U7295 ( .A1(n5791), .A2(SI_26_), .ZN(n5792) );
  AND2_X1 U7296 ( .A1(n5810), .A2(n5792), .ZN(n5808) );
  OR2_X1 U7297 ( .A1(n6581), .A2(n9563), .ZN(n5793) );
  NAND2_X1 U7298 ( .A1(n9244), .A2(n5631), .ZN(n5801) );
  NAND2_X1 U7299 ( .A1(n6585), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5799) );
  NAND2_X1 U7300 ( .A1(n5187), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5798) );
  INV_X1 U7301 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9040) );
  AOI21_X1 U7302 ( .B1(n5795), .B2(n9040), .A(n5818), .ZN(n9245) );
  NAND2_X1 U7303 ( .A1(n5886), .A2(n9245), .ZN(n5797) );
  NAND2_X1 U7304 ( .A1(n6584), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5796) );
  OR2_X1 U7305 ( .A1(n9455), .A2(n5863), .ZN(n5800) );
  NAND2_X1 U7306 ( .A1(n5801), .A2(n5800), .ZN(n5802) );
  XNOR2_X1 U7307 ( .A(n5802), .B(n5866), .ZN(n5804) );
  NOR2_X1 U7308 ( .A1(n9455), .A2(n5868), .ZN(n5803) );
  AOI21_X1 U7309 ( .B1(n9244), .B2(n5136), .A(n5803), .ZN(n5805) );
  XNOR2_X1 U7310 ( .A(n5804), .B(n5805), .ZN(n9035) );
  INV_X1 U7311 ( .A(n5804), .ZN(n5807) );
  INV_X1 U7312 ( .A(n5805), .ZN(n5806) );
  INV_X1 U7313 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5811) );
  INV_X1 U7314 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8735) );
  MUX2_X1 U7315 ( .A(n5811), .B(n8735), .S(n6857), .Z(n5813) );
  INV_X1 U7316 ( .A(SI_27_), .ZN(n5812) );
  NAND2_X1 U7317 ( .A1(n5813), .A2(n5812), .ZN(n5854) );
  INV_X1 U7318 ( .A(n5813), .ZN(n5814) );
  NAND2_X1 U7319 ( .A1(n5814), .A2(SI_27_), .ZN(n5815) );
  AND2_X1 U7320 ( .A1(n5854), .A2(n5815), .ZN(n5852) );
  OR2_X1 U7321 ( .A1(n6581), .A2(n8735), .ZN(n5816) );
  NAND2_X1 U7322 ( .A1(n9228), .A2(n5631), .ZN(n5825) );
  NAND2_X1 U7323 ( .A1(n6585), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5823) );
  NAND2_X1 U7324 ( .A1(n5885), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5822) );
  INV_X1 U7325 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8897) );
  INV_X1 U7326 ( .A(n5818), .ZN(n5819) );
  NAND2_X1 U7327 ( .A1(n5818), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5858) );
  INV_X1 U7328 ( .A(n5858), .ZN(n5857) );
  AOI21_X1 U7329 ( .B1(n8897), .B2(n5819), .A(n5857), .ZN(n9229) );
  NAND2_X1 U7330 ( .A1(n5886), .A2(n9229), .ZN(n5821) );
  NAND2_X1 U7331 ( .A1(n6584), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5820) );
  OR2_X1 U7332 ( .A1(n9252), .A2(n5863), .ZN(n5824) );
  NAND2_X1 U7333 ( .A1(n5825), .A2(n5824), .ZN(n5826) );
  XNOR2_X1 U7334 ( .A(n5826), .B(n5866), .ZN(n5829) );
  NOR2_X1 U7335 ( .A1(n9252), .A2(n5868), .ZN(n5827) );
  AOI21_X1 U7336 ( .B1(n9228), .B2(n5529), .A(n5827), .ZN(n5828) );
  NAND2_X1 U7337 ( .A1(n5829), .A2(n5828), .ZN(n5877) );
  OAI21_X1 U7338 ( .B1(n5829), .B2(n5828), .A(n5877), .ZN(n8896) );
  INV_X1 U7339 ( .A(P1_B_REG_SCAN_IN), .ZN(n9138) );
  OR2_X1 U7340 ( .A1(n5833), .A2(n9138), .ZN(n5831) );
  INV_X1 U7341 ( .A(n5830), .ZN(n7726) );
  MUX2_X1 U7342 ( .A(P1_B_REG_SCAN_IN), .B(n5831), .S(n7726), .Z(n5832) );
  NAND2_X1 U7343 ( .A1(n5832), .A2(n5834), .ZN(n9547) );
  OR2_X1 U7344 ( .A1(n9547), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5835) );
  INV_X1 U7345 ( .A(n5833), .ZN(n7782) );
  INV_X1 U7346 ( .A(n5834), .ZN(n9566) );
  NAND2_X1 U7347 ( .A1(n7782), .A2(n9566), .ZN(n9548) );
  NAND2_X1 U7348 ( .A1(n5835), .A2(n9548), .ZN(n6963) );
  INV_X1 U7349 ( .A(n6963), .ZN(n7228) );
  OR2_X1 U7350 ( .A1(n9547), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5836) );
  NAND2_X1 U7351 ( .A1(n9566), .A2(n7726), .ZN(n9549) );
  NOR4_X1 U7352 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5840) );
  NOR4_X1 U7353 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n5839) );
  NOR4_X1 U7354 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n5838) );
  NOR4_X1 U7355 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5837) );
  NAND4_X1 U7356 ( .A1(n5840), .A2(n5839), .A3(n5838), .A4(n5837), .ZN(n5846)
         );
  NOR2_X1 U7357 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .ZN(
        n5844) );
  NOR4_X1 U7358 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_31__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5843) );
  NOR4_X1 U7359 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5842) );
  NOR4_X1 U7360 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n5841) );
  NAND4_X1 U7361 ( .A1(n5844), .A2(n5843), .A3(n5842), .A4(n5841), .ZN(n5845)
         );
  NOR2_X1 U7362 ( .A1(n5846), .A2(n5845), .ZN(n5847) );
  OR2_X1 U7363 ( .A1(n9547), .A2(n5847), .ZN(n6965) );
  NAND3_X1 U7364 ( .A1(n7228), .A2(n6979), .A3(n6965), .ZN(n5891) );
  NAND2_X1 U7365 ( .A1(n4617), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5848) );
  XNOR2_X1 U7366 ( .A(n5848), .B(P1_IR_REG_23__SCAN_IN), .ZN(n6593) );
  INV_X1 U7367 ( .A(n6593), .ZN(n6882) );
  AND2_X1 U7368 ( .A1(n6882), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6847) );
  INV_X1 U7369 ( .A(n9546), .ZN(n6885) );
  OR2_X1 U7370 ( .A1(n5891), .A2(n6885), .ZN(n5881) );
  INV_X1 U7371 ( .A(n5881), .ZN(n5851) );
  NOR2_X2 U7372 ( .A1(n6977), .A2(n6740), .ZN(n9997) );
  NOR2_X1 U7373 ( .A1(n9997), .A2(n7279), .ZN(n5850) );
  NAND2_X1 U7374 ( .A1(n5851), .A2(n5850), .ZN(n9056) );
  MUX2_X1 U7375 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n6857), .Z(n6327) );
  INV_X1 U7376 ( .A(SI_28_), .ZN(n6328) );
  XNOR2_X1 U7377 ( .A(n6327), .B(n6328), .ZN(n6325) );
  NAND2_X1 U7378 ( .A1(n9559), .A2(n6583), .ZN(n5856) );
  INV_X1 U7379 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9561) );
  OR2_X1 U7380 ( .A1(n6581), .A2(n9561), .ZN(n5855) );
  NAND2_X1 U7381 ( .A1(n9450), .A2(n5631), .ZN(n5865) );
  NAND2_X1 U7382 ( .A1(n6585), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U7383 ( .A1(n5187), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5861) );
  INV_X1 U7384 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5883) );
  AOI21_X1 U7385 ( .B1(n5883), .B2(n5858), .A(n9202), .ZN(n5895) );
  NAND2_X1 U7386 ( .A1(n5886), .A2(n5895), .ZN(n5860) );
  NAND2_X1 U7387 ( .A1(n6584), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5859) );
  OR2_X1 U7388 ( .A1(n9236), .A2(n5863), .ZN(n5864) );
  NAND2_X1 U7389 ( .A1(n5865), .A2(n5864), .ZN(n5867) );
  XNOR2_X1 U7390 ( .A(n5867), .B(n5866), .ZN(n5871) );
  NOR2_X1 U7391 ( .A1(n9236), .A2(n5868), .ZN(n5869) );
  AOI21_X1 U7392 ( .B1(n9450), .B2(n5136), .A(n5869), .ZN(n5870) );
  XNOR2_X1 U7393 ( .A(n5871), .B(n5870), .ZN(n5874) );
  INV_X1 U7394 ( .A(n5874), .ZN(n5878) );
  NAND3_X1 U7395 ( .A1(n8894), .A2(n9038), .A3(n5878), .ZN(n5903) );
  NOR2_X1 U7396 ( .A1(n5872), .A2(n9056), .ZN(n5873) );
  AND2_X1 U7397 ( .A1(n5874), .A2(n5873), .ZN(n5875) );
  NAND2_X1 U7398 ( .A1(n5876), .A2(n5875), .ZN(n5902) );
  NAND3_X1 U7399 ( .A1(n5878), .A2(n5872), .A3(n9038), .ZN(n5900) );
  INV_X1 U7400 ( .A(n6977), .ZN(n7230) );
  NAND2_X1 U7401 ( .A1(n7230), .A2(n6744), .ZN(n7236) );
  NOR2_X2 U7402 ( .A1(n6977), .A2(n6744), .ZN(n9900) );
  AND2_X1 U7403 ( .A1(n9546), .A2(n4722), .ZN(n5879) );
  NAND2_X1 U7404 ( .A1(n9900), .A2(n5879), .ZN(n9893) );
  AND2_X1 U7405 ( .A1(n7279), .A2(n6740), .ZN(n7231) );
  INV_X1 U7406 ( .A(n7231), .ZN(n5880) );
  NOR2_X1 U7407 ( .A1(n5881), .A2(n5880), .ZN(n5884) );
  INV_X1 U7408 ( .A(n5882), .ZN(n9066) );
  NAND2_X1 U7409 ( .A1(n5884), .A2(n9066), .ZN(n9041) );
  OAI22_X1 U7410 ( .A1(n9041), .A2(n9252), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5883), .ZN(n5898) );
  NAND2_X1 U7411 ( .A1(n5884), .A2(n5882), .ZN(n9053) );
  NAND2_X1 U7412 ( .A1(n5885), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U7413 ( .A1(n6585), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5889) );
  NAND2_X1 U7414 ( .A1(n6584), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5888) );
  NAND2_X1 U7415 ( .A1(n5886), .A2(n9202), .ZN(n5887) );
  NAND4_X1 U7416 ( .A1(n5890), .A2(n5889), .A3(n5888), .A4(n5887), .ZN(n9210)
         );
  INV_X1 U7417 ( .A(n9210), .ZN(n5896) );
  NAND2_X1 U7418 ( .A1(n9900), .A2(n4722), .ZN(n6962) );
  NAND2_X1 U7419 ( .A1(n5891), .A2(n6962), .ZN(n5893) );
  NAND2_X1 U7420 ( .A1(n7279), .A2(n6969), .ZN(n6964) );
  AND2_X1 U7421 ( .A1(n6964), .A2(n6848), .ZN(n5892) );
  NAND2_X1 U7422 ( .A1(n5893), .A2(n5892), .ZN(n6909) );
  OR2_X1 U7423 ( .A1(n6909), .A2(n6593), .ZN(n5894) );
  NAND2_X1 U7424 ( .A1(n5894), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9029) );
  INV_X1 U7425 ( .A(n5895), .ZN(n9218) );
  OAI22_X1 U7426 ( .A1(n9053), .A2(n5896), .B1(n9029), .B2(n9218), .ZN(n5897)
         );
  NAND3_X1 U7427 ( .A1(n5903), .A2(n5902), .A3(n5901), .ZN(P1_U3220) );
  NAND4_X1 U7428 ( .A1(n5905), .A2(n6068), .A3(n5904), .A4(n8631), .ZN(n5906)
         );
  NOR2_X1 U7429 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5912) );
  NOR2_X1 U7430 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5911) );
  NOR2_X1 U7431 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5910) );
  INV_X1 U7432 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5915) );
  INV_X1 U7433 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6499) );
  INV_X1 U7434 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6497) );
  NAND2_X1 U7435 ( .A1(n6503), .A2(n5916), .ZN(n5921) );
  OAI21_X1 U7436 ( .B1(n5919), .B2(n8876), .A(P2_IR_REG_28__SCAN_IN), .ZN(
        n5917) );
  INV_X1 U7437 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5918) );
  INV_X1 U7438 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5922) );
  XNOR2_X2 U7439 ( .A(n5923), .B(n5922), .ZN(n6509) );
  NAND2_X1 U7440 ( .A1(n7723), .A2(n6387), .ZN(n5925) );
  OR2_X1 U7441 ( .A1(n6037), .A2(n8647), .ZN(n5924) );
  INV_X1 U7442 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5931) );
  INV_X1 U7443 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7789) );
  INV_X1 U7444 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5934) );
  INV_X1 U7445 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5935) );
  INV_X1 U7446 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8676) );
  INV_X1 U7447 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5937) );
  INV_X1 U7448 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8649) );
  INV_X1 U7449 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5938) );
  NAND2_X1 U7450 ( .A1(n5956), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5939) );
  NAND2_X1 U7451 ( .A1(n5971), .A2(n5939), .ZN(n8315) );
  NAND2_X1 U7452 ( .A1(n5941), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5940) );
  MUX2_X1 U7453 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5940), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5943) );
  INV_X1 U7454 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5942) );
  NAND2_X1 U7455 ( .A1(n8315), .A2(n6018), .ZN(n5952) );
  NOR2_X1 U7456 ( .A1(n7825), .A2(n5947), .ZN(n6016) );
  INV_X1 U7457 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8661) );
  NAND2_X1 U7458 ( .A1(n4460), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5949) );
  NAND2_X1 U7459 ( .A1(n4461), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5948) );
  OAI211_X1 U7460 ( .C1(n4463), .C2(n8661), .A(n5949), .B(n5948), .ZN(n5950)
         );
  INV_X1 U7461 ( .A(n5950), .ZN(n5951) );
  NAND2_X1 U7462 ( .A1(n7656), .A2(n6387), .ZN(n5954) );
  NAND2_X1 U7463 ( .A1(n6332), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5953) );
  INV_X1 U7464 ( .A(n4461), .ZN(n6349) );
  INV_X1 U7465 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U7466 ( .A1(n5982), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5955) );
  NAND2_X1 U7467 ( .A1(n5956), .A2(n5955), .ZN(n8326) );
  NAND2_X1 U7468 ( .A1(n8326), .A2(n6018), .ZN(n5958) );
  INV_X1 U7469 ( .A(n4460), .ZN(n6366) );
  AOI22_X1 U7470 ( .A1(n6346), .A2(P2_REG0_REG_23__SCAN_IN), .B1(n6048), .B2(
        P2_REG1_REG_23__SCAN_IN), .ZN(n5957) );
  INV_X1 U7471 ( .A(n6453), .ZN(n5960) );
  AND2_X1 U7472 ( .A1(n6436), .A2(n5960), .ZN(n5961) );
  OR2_X1 U7473 ( .A1(n5961), .A2(n6435), .ZN(n5966) );
  OR2_X1 U7474 ( .A1(n8325), .A2(n8334), .ZN(n6434) );
  INV_X1 U7475 ( .A(n6434), .ZN(n6454) );
  OAI21_X1 U7476 ( .B1(n6435), .B2(n6454), .A(n6436), .ZN(n5965) );
  NAND2_X1 U7477 ( .A1(n4494), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U7478 ( .A1(n5963), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5964) );
  MUX2_X1 U7479 ( .A(n5966), .B(n5965), .S(n6839), .Z(n6299) );
  NAND2_X1 U7480 ( .A1(n7755), .A2(n6387), .ZN(n5968) );
  NAND2_X1 U7481 ( .A1(n6332), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5967) );
  INV_X1 U7482 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U7483 ( .A1(n5971), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U7484 ( .A1(n6302), .A2(n5972), .ZN(n8305) );
  NAND2_X1 U7485 ( .A1(n8305), .A2(n6018), .ZN(n5977) );
  INV_X1 U7486 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8536) );
  NAND2_X1 U7487 ( .A1(n4461), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5974) );
  NAND2_X1 U7488 ( .A1(n6048), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5973) );
  OAI211_X1 U7489 ( .C1(n6366), .C2(n8536), .A(n5974), .B(n5973), .ZN(n5975)
         );
  INV_X1 U7490 ( .A(n5975), .ZN(n5976) );
  NAND2_X1 U7491 ( .A1(n8304), .A2(n8313), .ZN(n6437) );
  INV_X1 U7492 ( .A(n6436), .ZN(n5978) );
  NAND2_X1 U7493 ( .A1(n7541), .A2(n6387), .ZN(n5980) );
  NAND2_X1 U7494 ( .A1(n6332), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5979) );
  NAND2_X1 U7495 ( .A1(n5991), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7496 ( .A1(n5982), .A2(n5981), .ZN(n8337) );
  NAND2_X1 U7497 ( .A1(n8337), .A2(n6018), .ZN(n5985) );
  AOI22_X1 U7498 ( .A1(n6346), .A2(P2_REG0_REG_22__SCAN_IN), .B1(n6048), .B2(
        P2_REG1_REG_22__SCAN_IN), .ZN(n5984) );
  NAND2_X1 U7499 ( .A1(n4461), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5983) );
  NAND2_X1 U7500 ( .A1(n8012), .A2(n8344), .ZN(n6433) );
  NAND2_X1 U7501 ( .A1(n6432), .A2(n6433), .ZN(n8335) );
  NAND2_X1 U7502 ( .A1(n7513), .A2(n6387), .ZN(n5987) );
  NAND2_X1 U7503 ( .A1(n6332), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7504 ( .A1(n6048), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5989) );
  NAND2_X1 U7505 ( .A1(n6346), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5988) );
  AND2_X1 U7506 ( .A1(n5989), .A2(n5988), .ZN(n5994) );
  NAND2_X1 U7507 ( .A1(n6281), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7508 ( .A1(n5991), .A2(n5990), .ZN(n8350) );
  NAND2_X1 U7509 ( .A1(n8350), .A2(n6018), .ZN(n5993) );
  NAND2_X1 U7510 ( .A1(n4462), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5992) );
  NAND2_X1 U7511 ( .A1(n7931), .A2(n8333), .ZN(n6455) );
  NAND2_X1 U7512 ( .A1(n6016), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5999) );
  NAND2_X1 U7513 ( .A1(n4460), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U7514 ( .A1(n6018), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5996) );
  NAND2_X1 U7515 ( .A1(n4462), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5995) );
  NAND3_X2 U7516 ( .A1(n5999), .A2(n5998), .A3(n5997), .ZN(n6010) );
  INV_X1 U7517 ( .A(n6010), .ZN(n6002) );
  NAND2_X1 U7518 ( .A1(n6000), .A2(SI_0_), .ZN(n6001) );
  XNOR2_X1 U7519 ( .A(n6001), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8891) );
  NAND2_X1 U7520 ( .A1(n6002), .A2(n7037), .ZN(n7169) );
  INV_X1 U7521 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6868) );
  NAND2_X1 U7522 ( .A1(n6016), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6009) );
  NAND2_X1 U7523 ( .A1(n6017), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6008) );
  NAND2_X1 U7524 ( .A1(n6018), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7525 ( .A1(n6019), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6006) );
  INV_X1 U7526 ( .A(n7037), .ZN(n7189) );
  NAND2_X1 U7527 ( .A1(n6010), .A2(n7189), .ZN(n6463) );
  NAND2_X1 U7528 ( .A1(n6463), .A2(n7165), .ZN(n6011) );
  NAND2_X1 U7529 ( .A1(n6407), .A2(n6011), .ZN(n6012) );
  NAND2_X1 U7530 ( .A1(n6012), .A2(n6839), .ZN(n6013) );
  OAI21_X1 U7531 ( .B1(n7165), .B2(n7169), .A(n6013), .ZN(n6015) );
  INV_X2 U7532 ( .A(n6757), .ZN(n8089) );
  AOI21_X1 U7533 ( .B1(n6406), .B2(n6463), .A(n6839), .ZN(n6014) );
  AOI21_X1 U7534 ( .B1(n6015), .B2(n6406), .A(n6014), .ZN(n6030) );
  NOR2_X1 U7535 ( .A1(n6407), .A2(n6839), .ZN(n6029) );
  NAND2_X1 U7536 ( .A1(n6016), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U7537 ( .A1(n4460), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6022) );
  NAND2_X1 U7538 ( .A1(n6018), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6021) );
  NAND2_X1 U7539 ( .A1(n4461), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6020) );
  INV_X1 U7540 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6862) );
  OR2_X1 U7541 ( .A1(n6038), .A2(n6861), .ZN(n6027) );
  OAI211_X1 U7542 ( .C1(n6756), .C2(n4571), .A(n6028), .B(n6027), .ZN(n7092)
         );
  NAND2_X1 U7543 ( .A1(n7121), .A2(n7092), .ZN(n6409) );
  OR3_X1 U7544 ( .A1(n6030), .A2(n6029), .A3(n10156), .ZN(n6047) );
  NAND2_X1 U7545 ( .A1(n6018), .A2(n7179), .ZN(n6034) );
  NAND2_X1 U7546 ( .A1(n4460), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6033) );
  NAND2_X1 U7547 ( .A1(n6016), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6032) );
  NAND2_X1 U7548 ( .A1(n4461), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7549 ( .A1(n6035), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6036) );
  XNOR2_X1 U7550 ( .A(n6036), .B(P2_IR_REG_3__SCAN_IN), .ZN(n7139) );
  INV_X1 U7551 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6864) );
  OR2_X1 U7552 ( .A1(n6037), .A2(n6864), .ZN(n6040) );
  OR2_X1 U7553 ( .A1(n6038), .A2(n6863), .ZN(n6039) );
  OAI211_X1 U7554 ( .C1(n6756), .C2(n4838), .A(n6040), .B(n6039), .ZN(n10179)
         );
  INV_X1 U7555 ( .A(n10179), .ZN(n6041) );
  NAND2_X1 U7556 ( .A1(n8088), .A2(n6041), .ZN(n6060) );
  NAND2_X1 U7557 ( .A1(n6060), .A2(n6042), .ZN(n6044) );
  NAND2_X1 U7558 ( .A1(n10159), .A2(n10179), .ZN(n6410) );
  NAND2_X1 U7559 ( .A1(n6409), .A2(n6410), .ZN(n6043) );
  MUX2_X1 U7560 ( .A(n6044), .B(n6043), .S(n6839), .Z(n6045) );
  INV_X1 U7561 ( .A(n6045), .ZN(n6046) );
  NAND2_X1 U7562 ( .A1(n6047), .A2(n6046), .ZN(n6059) );
  NAND2_X1 U7563 ( .A1(n6016), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7564 ( .A1(n4461), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U7565 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6049) );
  NAND2_X1 U7566 ( .A1(n6061), .A2(n6049), .ZN(n7271) );
  NAND2_X1 U7567 ( .A1(n6018), .A2(n7271), .ZN(n6051) );
  NAND2_X1 U7568 ( .A1(n4460), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6050) );
  INV_X1 U7569 ( .A(n8087), .ZN(n7258) );
  NAND2_X1 U7570 ( .A1(n6054), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6055) );
  INV_X1 U7571 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n8672) );
  OR2_X1 U7572 ( .A1(n6037), .A2(n8672), .ZN(n6057) );
  OR2_X1 U7573 ( .A1(n6038), .A2(n6866), .ZN(n6056) );
  OAI211_X1 U7574 ( .C1(n6756), .C2(n7148), .A(n6057), .B(n6056), .ZN(n7257)
         );
  INV_X1 U7575 ( .A(n7257), .ZN(n7266) );
  NAND2_X1 U7576 ( .A1(n7258), .A2(n7266), .ZN(n6764) );
  AND2_X1 U7577 ( .A1(n8087), .A2(n7257), .ZN(n6765) );
  INV_X1 U7578 ( .A(n6765), .ZN(n6058) );
  NAND2_X1 U7579 ( .A1(n6059), .A2(n7199), .ZN(n6090) );
  INV_X1 U7580 ( .A(n6060), .ZN(n6074) );
  NAND2_X1 U7581 ( .A1(n4460), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6066) );
  NAND2_X1 U7582 ( .A1(n6016), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7583 ( .A1(n6061), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7584 ( .A1(n6075), .A2(n6062), .ZN(n7396) );
  NAND2_X1 U7585 ( .A1(n6018), .A2(n7396), .ZN(n6064) );
  NAND2_X1 U7586 ( .A1(n4461), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6063) );
  INV_X1 U7587 ( .A(n8086), .ZN(n7435) );
  NOR2_X1 U7588 ( .A1(n6054), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n6069) );
  NOR2_X1 U7589 ( .A1(n6069), .A2(n8876), .ZN(n6067) );
  MUX2_X1 U7590 ( .A(n8876), .B(n6067), .S(P2_IR_REG_5__SCAN_IN), .Z(n6071) );
  NAND2_X1 U7591 ( .A1(n6069), .A2(n6068), .ZN(n6082) );
  INV_X1 U7592 ( .A(n6082), .ZN(n6070) );
  INV_X1 U7593 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6871) );
  OR2_X1 U7594 ( .A1(n6037), .A2(n6871), .ZN(n6073) );
  OR2_X1 U7595 ( .A1(n6038), .A2(n6870), .ZN(n6072) );
  OAI211_X1 U7596 ( .C1(n6756), .C2(n10078), .A(n6073), .B(n6072), .ZN(n7397)
         );
  NAND2_X1 U7597 ( .A1(n7435), .A2(n7397), .ZN(n6465) );
  NAND2_X1 U7598 ( .A1(n7258), .A2(n7257), .ZN(n6411) );
  OAI211_X1 U7599 ( .C1(n6090), .C2(n6074), .A(n6465), .B(n6411), .ZN(n6087)
         );
  INV_X1 U7600 ( .A(n7397), .ZN(n6766) );
  NAND2_X1 U7601 ( .A1(n8086), .A2(n6766), .ZN(n6464) );
  NAND2_X1 U7602 ( .A1(n6346), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7603 ( .A1(n6048), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U7604 ( .A1(n6075), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7605 ( .A1(n6097), .A2(n6076), .ZN(n8044) );
  NAND2_X1 U7606 ( .A1(n6018), .A2(n8044), .ZN(n6078) );
  NAND2_X1 U7607 ( .A1(n4461), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U7608 ( .A1(n6082), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6081) );
  MUX2_X1 U7609 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6081), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n6083) );
  OR2_X1 U7610 ( .A1(n6038), .A2(n6873), .ZN(n6085) );
  INV_X1 U7611 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6872) );
  OR2_X1 U7612 ( .A1(n6037), .A2(n6872), .ZN(n6084) );
  OAI211_X1 U7613 ( .C1(n6756), .C2(n7626), .A(n6085), .B(n6084), .ZN(n7438)
         );
  INV_X1 U7614 ( .A(n7438), .ZN(n8040) );
  NAND2_X1 U7615 ( .A1(n8085), .A2(n8040), .ZN(n6415) );
  AND2_X1 U7616 ( .A1(n6464), .A2(n6415), .ZN(n6086) );
  NOR2_X1 U7617 ( .A1(n8085), .A2(n8040), .ZN(n6414) );
  AOI21_X1 U7618 ( .B1(n6087), .B2(n6086), .A(n6414), .ZN(n6096) );
  INV_X1 U7619 ( .A(n6410), .ZN(n6089) );
  NAND2_X1 U7620 ( .A1(n8087), .A2(n7266), .ZN(n6088) );
  OAI211_X1 U7621 ( .C1(n6090), .C2(n6089), .A(n6088), .B(n6464), .ZN(n6094)
         );
  INV_X1 U7622 ( .A(n6465), .ZN(n6091) );
  NOR2_X1 U7623 ( .A1(n6091), .A2(n6414), .ZN(n6093) );
  INV_X1 U7624 ( .A(n6415), .ZN(n6092) );
  AOI21_X1 U7625 ( .B1(n6094), .B2(n6093), .A(n6092), .ZN(n6095) );
  MUX2_X1 U7626 ( .A(n6096), .B(n6095), .S(n6851), .Z(n6127) );
  NAND2_X1 U7627 ( .A1(n6346), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6102) );
  NAND2_X1 U7628 ( .A1(n6048), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U7629 ( .A1(n6097), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7630 ( .A1(n6106), .A2(n6098), .ZN(n7475) );
  NAND2_X1 U7631 ( .A1(n6018), .A2(n7475), .ZN(n6100) );
  NAND2_X1 U7632 ( .A1(n4462), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6099) );
  NAND2_X1 U7633 ( .A1(n6112), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6103) );
  XNOR2_X1 U7634 ( .A(n6103), .B(n8631), .ZN(n10111) );
  OR2_X1 U7635 ( .A1(n6038), .A2(n6875), .ZN(n6105) );
  INV_X1 U7636 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n8780) );
  OR2_X1 U7637 ( .A1(n6037), .A2(n8780), .ZN(n6104) );
  NAND2_X1 U7638 ( .A1(n7530), .A2(n7447), .ZN(n6142) );
  NAND2_X1 U7639 ( .A1(n8084), .A2(n10201), .ZN(n7520) );
  NAND2_X1 U7640 ( .A1(n6142), .A2(n7520), .ZN(n7479) );
  INV_X1 U7641 ( .A(n7479), .ZN(n6467) );
  NAND2_X1 U7642 ( .A1(n6346), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U7643 ( .A1(n6048), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6110) );
  NAND2_X1 U7644 ( .A1(n6106), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6107) );
  NAND2_X1 U7645 ( .A1(n6116), .A2(n6107), .ZN(n7539) );
  NAND2_X1 U7646 ( .A1(n6018), .A2(n7539), .ZN(n6109) );
  NAND2_X1 U7647 ( .A1(n4461), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U7648 ( .A1(n6877), .A2(n6387), .ZN(n6115) );
  OAI21_X1 U7649 ( .B1(n6112), .B2(P2_IR_REG_7__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6113) );
  XNOR2_X1 U7650 ( .A(n6113), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10140) );
  AOI22_X1 U7651 ( .A1(n6332), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6853), .B2(
        n10140), .ZN(n6114) );
  INV_X1 U7652 ( .A(n7532), .ZN(n6769) );
  NAND2_X1 U7653 ( .A1(n7558), .A2(n6769), .ZN(n6470) );
  NAND2_X1 U7654 ( .A1(n6346), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6121) );
  NAND2_X1 U7655 ( .A1(n6048), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U7656 ( .A1(n6116), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6117) );
  NAND2_X1 U7657 ( .A1(n6135), .A2(n6117), .ZN(n7577) );
  NAND2_X1 U7658 ( .A1(n6018), .A2(n7577), .ZN(n6119) );
  NAND2_X1 U7659 ( .A1(n4462), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6118) );
  NAND2_X1 U7660 ( .A1(n6891), .A2(n6387), .ZN(n6125) );
  OR2_X1 U7661 ( .A1(n6122), .A2(n8876), .ZN(n6123) );
  XNOR2_X1 U7662 ( .A(n6123), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7666) );
  AOI22_X1 U7663 ( .A1(n6332), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6853), .B2(
        n7666), .ZN(n6124) );
  INV_X1 U7664 ( .A(n7562), .ZN(n7580) );
  NAND2_X1 U7665 ( .A1(n7714), .A2(n7580), .ZN(n6418) );
  NAND3_X1 U7666 ( .A1(n6470), .A2(n6418), .A3(n6839), .ZN(n6141) );
  NAND2_X1 U7667 ( .A1(n7562), .A2(n8082), .ZN(n7715) );
  NAND2_X1 U7668 ( .A1(n8083), .A2(n7532), .ZN(n6469) );
  NAND3_X1 U7669 ( .A1(n7715), .A2(n6851), .A3(n6469), .ZN(n6126) );
  NAND2_X1 U7670 ( .A1(n6141), .A2(n6126), .ZN(n6144) );
  NAND3_X1 U7671 ( .A1(n6127), .A2(n6467), .A3(n6144), .ZN(n6150) );
  AND2_X1 U7672 ( .A1(n7520), .A2(n6469), .ZN(n6416) );
  OR2_X1 U7673 ( .A1(n6890), .A2(n6038), .ZN(n6134) );
  NOR2_X1 U7674 ( .A1(n6128), .A2(n8876), .ZN(n6129) );
  MUX2_X1 U7675 ( .A(n8876), .B(n6129), .S(P2_IR_REG_10__SCAN_IN), .Z(n6132)
         );
  INV_X1 U7676 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6130) );
  NAND2_X1 U7677 ( .A1(n6128), .A2(n6130), .ZN(n6166) );
  INV_X1 U7678 ( .A(n6166), .ZN(n6131) );
  OR2_X1 U7679 ( .A1(n6132), .A2(n6131), .ZN(n7763) );
  INV_X1 U7680 ( .A(n7763), .ZN(n7678) );
  AOI22_X1 U7681 ( .A1(n6332), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6853), .B2(
        n7678), .ZN(n6133) );
  NAND2_X1 U7682 ( .A1(n6346), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7683 ( .A1(n6048), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6139) );
  NAND2_X1 U7684 ( .A1(n6135), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6136) );
  NAND2_X1 U7685 ( .A1(n6154), .A2(n6136), .ZN(n7910) );
  NAND2_X1 U7686 ( .A1(n6018), .A2(n7910), .ZN(n6138) );
  NAND2_X1 U7687 ( .A1(n4461), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6137) );
  NAND4_X1 U7688 ( .A1(n6140), .A2(n6139), .A3(n6138), .A4(n6137), .ZN(n8081)
         );
  OR2_X1 U7689 ( .A1(n7901), .A2(n7832), .ZN(n7711) );
  OAI21_X1 U7690 ( .B1(n6416), .B2(n6141), .A(n6475), .ZN(n6147) );
  NAND2_X1 U7691 ( .A1(n6470), .A2(n6142), .ZN(n6143) );
  NAND2_X1 U7692 ( .A1(n6144), .A2(n6143), .ZN(n6145) );
  NAND2_X1 U7693 ( .A1(n7901), .A2(n7832), .ZN(n7727) );
  AND2_X1 U7694 ( .A1(n7727), .A2(n6418), .ZN(n6474) );
  NAND2_X1 U7695 ( .A1(n6145), .A2(n6474), .ZN(n6146) );
  MUX2_X1 U7696 ( .A(n6147), .B(n6146), .S(n6851), .Z(n6148) );
  INV_X1 U7697 ( .A(n6148), .ZN(n6149) );
  NAND2_X1 U7698 ( .A1(n6900), .A2(n6387), .ZN(n6153) );
  NAND2_X1 U7699 ( .A1(n6166), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6151) );
  XNOR2_X1 U7700 ( .A(n6151), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7792) );
  AOI22_X1 U7701 ( .A1(n6332), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6853), .B2(
        n7792), .ZN(n6152) );
  NAND2_X1 U7702 ( .A1(n6153), .A2(n6152), .ZN(n8015) );
  NAND2_X1 U7703 ( .A1(n6346), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6159) );
  NAND2_X1 U7704 ( .A1(n6048), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U7705 ( .A1(n6154), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6155) );
  NAND2_X1 U7706 ( .A1(n6170), .A2(n6155), .ZN(n8023) );
  NAND2_X1 U7707 ( .A1(n6018), .A2(n8023), .ZN(n6157) );
  NAND2_X1 U7708 ( .A1(n4461), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6156) );
  NAND2_X1 U7709 ( .A1(n8015), .A2(n7908), .ZN(n6461) );
  AND2_X1 U7710 ( .A1(n6461), .A2(n7727), .ZN(n6419) );
  INV_X1 U7711 ( .A(n6462), .ZN(n6160) );
  AOI21_X1 U7712 ( .B1(n6163), .B2(n6419), .A(n6160), .ZN(n6165) );
  AND2_X1 U7713 ( .A1(n6462), .A2(n7711), .ZN(n6162) );
  INV_X1 U7714 ( .A(n6461), .ZN(n6161) );
  MUX2_X1 U7715 ( .A(n6165), .B(n6164), .S(n6851), .Z(n6176) );
  OR2_X1 U7716 ( .A1(n6905), .A2(n6038), .ZN(n6169) );
  NAND2_X1 U7717 ( .A1(n6177), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6167) );
  XNOR2_X1 U7718 ( .A(n6167), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8106) );
  AOI22_X1 U7719 ( .A1(n6332), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6853), .B2(
        n8106), .ZN(n6168) );
  NAND2_X1 U7720 ( .A1(n6346), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U7721 ( .A1(n6048), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6174) );
  NAND2_X1 U7722 ( .A1(n6170), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U7723 ( .A1(n6181), .A2(n6171), .ZN(n7950) );
  NAND2_X1 U7724 ( .A1(n6018), .A2(n7950), .ZN(n6173) );
  NAND2_X1 U7725 ( .A1(n4462), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6172) );
  NAND4_X1 U7726 ( .A1(n6175), .A2(n6174), .A3(n6173), .A4(n6172), .ZN(n8080)
         );
  XNOR2_X1 U7727 ( .A(n7939), .B(n8080), .ZN(n6459) );
  NAND2_X1 U7728 ( .A1(n6176), .A2(n6459), .ZN(n6190) );
  OR2_X1 U7729 ( .A1(n6984), .A2(n6038), .ZN(n6180) );
  NAND2_X1 U7730 ( .A1(n6251), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6178) );
  XNOR2_X1 U7731 ( .A(n6178), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8099) );
  AOI22_X1 U7732 ( .A1(n6332), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6853), .B2(
        n8099), .ZN(n6179) );
  NAND2_X1 U7733 ( .A1(n6048), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6186) );
  NAND2_X1 U7734 ( .A1(n6346), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6185) );
  NAND2_X1 U7735 ( .A1(n6181), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6182) );
  NAND2_X1 U7736 ( .A1(n6193), .A2(n6182), .ZN(n8000) );
  NAND2_X1 U7737 ( .A1(n6018), .A2(n8000), .ZN(n6184) );
  NAND2_X1 U7738 ( .A1(n4461), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6183) );
  NAND4_X1 U7739 ( .A1(n6186), .A2(n6185), .A3(n6184), .A4(n6183), .ZN(n8436)
         );
  OR2_X1 U7740 ( .A1(n9636), .A2(n8436), .ZN(n6775) );
  AND2_X1 U7741 ( .A1(n9636), .A2(n8436), .ZN(n6774) );
  INV_X1 U7742 ( .A(n6774), .ZN(n6200) );
  NAND2_X1 U7743 ( .A1(n6775), .A2(n6200), .ZN(n6460) );
  OR2_X1 U7744 ( .A1(n7939), .A2(n6839), .ZN(n6188) );
  NAND2_X1 U7745 ( .A1(n7939), .A2(n6839), .ZN(n6187) );
  MUX2_X1 U7746 ( .A(n6188), .B(n6187), .S(n8454), .Z(n6189) );
  NAND3_X1 U7747 ( .A1(n6190), .A2(n6460), .A3(n6189), .ZN(n6202) );
  OR2_X1 U7748 ( .A1(n7019), .A2(n6038), .ZN(n6192) );
  OAI21_X1 U7749 ( .B1(n6251), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6204) );
  XNOR2_X1 U7750 ( .A(n6204), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8154) );
  AOI22_X1 U7751 ( .A1(n6332), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6853), .B2(
        n8154), .ZN(n6191) );
  NAND2_X1 U7752 ( .A1(n6048), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6198) );
  NAND2_X1 U7753 ( .A1(n6193), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7754 ( .A1(n6208), .A2(n6194), .ZN(n8439) );
  NAND2_X1 U7755 ( .A1(n6018), .A2(n8439), .ZN(n6197) );
  NAND2_X1 U7756 ( .A1(n4461), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6196) );
  NAND2_X1 U7757 ( .A1(n6346), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U7758 ( .A1(n9632), .A2(n8453), .ZN(n6214) );
  MUX2_X1 U7759 ( .A(n8436), .B(n9636), .S(n6851), .Z(n6199) );
  NAND2_X1 U7760 ( .A1(n6200), .A2(n6199), .ZN(n6201) );
  NAND3_X1 U7761 ( .A1(n6202), .A2(n4811), .A3(n6201), .ZN(n6216) );
  OR2_X1 U7762 ( .A1(n7088), .A2(n6038), .ZN(n6207) );
  INV_X1 U7763 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6203) );
  NAND2_X1 U7764 ( .A1(n6204), .A2(n6203), .ZN(n6205) );
  NAND2_X1 U7765 ( .A1(n6205), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6218) );
  XNOR2_X1 U7766 ( .A(n6218), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8148) );
  AOI22_X1 U7767 ( .A1(n6332), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6853), .B2(
        n8148), .ZN(n6206) );
  NAND2_X1 U7768 ( .A1(n4460), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6213) );
  NAND2_X1 U7769 ( .A1(n6048), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U7770 ( .A1(n6208), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U7771 ( .A1(n6225), .A2(n6209), .ZN(n8425) );
  NAND2_X1 U7772 ( .A1(n6018), .A2(n8425), .ZN(n6211) );
  NAND2_X1 U7773 ( .A1(n4461), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U7774 ( .A1(n8430), .A2(n8404), .ZN(n6231) );
  NAND2_X1 U7775 ( .A1(n6425), .A2(n6231), .ZN(n8418) );
  INV_X1 U7776 ( .A(n8418), .ZN(n8415) );
  MUX2_X1 U7777 ( .A(n6214), .B(n6424), .S(n6851), .Z(n6215) );
  NAND3_X1 U7778 ( .A1(n6216), .A2(n8415), .A3(n6215), .ZN(n6233) );
  NAND2_X1 U7779 ( .A1(n7125), .A2(n6387), .ZN(n6224) );
  INV_X1 U7780 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7781 ( .A1(n6218), .A2(n6217), .ZN(n6219) );
  NAND2_X1 U7782 ( .A1(n6219), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6221) );
  NAND2_X1 U7783 ( .A1(n6221), .A2(n6220), .ZN(n6234) );
  OR2_X1 U7784 ( .A1(n6221), .A2(n6220), .ZN(n6222) );
  AND2_X1 U7785 ( .A1(n6234), .A2(n6222), .ZN(n8190) );
  AOI22_X1 U7786 ( .A1(n6332), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6853), .B2(
        n8190), .ZN(n6223) );
  NAND2_X1 U7787 ( .A1(n6346), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6230) );
  NAND2_X1 U7788 ( .A1(n6048), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6229) );
  NAND2_X1 U7789 ( .A1(n6225), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6226) );
  NAND2_X1 U7790 ( .A1(n6238), .A2(n6226), .ZN(n8409) );
  NAND2_X1 U7791 ( .A1(n6018), .A2(n8409), .ZN(n6228) );
  NAND2_X1 U7792 ( .A1(n4461), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6227) );
  XNOR2_X1 U7793 ( .A(n8408), .B(n8065), .ZN(n8401) );
  INV_X1 U7794 ( .A(n8401), .ZN(n8406) );
  MUX2_X1 U7795 ( .A(n6231), .B(n6425), .S(n6839), .Z(n6232) );
  NAND3_X1 U7796 ( .A1(n6233), .A2(n8406), .A3(n6232), .ZN(n6247) );
  NAND2_X1 U7797 ( .A1(n7192), .A2(n6387), .ZN(n6237) );
  NAND2_X1 U7798 ( .A1(n6234), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6235) );
  XNOR2_X1 U7799 ( .A(n6235), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8219) );
  AOI22_X1 U7800 ( .A1(n6332), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6853), .B2(
        n8219), .ZN(n6236) );
  NAND2_X1 U7801 ( .A1(n6346), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6243) );
  NAND2_X1 U7802 ( .A1(n6048), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6242) );
  NAND2_X1 U7803 ( .A1(n6238), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6239) );
  NAND2_X1 U7804 ( .A1(n6255), .A2(n6239), .ZN(n8394) );
  NAND2_X1 U7805 ( .A1(n6018), .A2(n8394), .ZN(n6241) );
  NAND2_X1 U7806 ( .A1(n4461), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6240) );
  NAND4_X1 U7807 ( .A1(n6243), .A2(n6242), .A3(n6241), .A4(n6240), .ZN(n8079)
         );
  XNOR2_X1 U7808 ( .A(n8511), .B(n8079), .ZN(n6781) );
  NAND2_X1 U7809 ( .A1(n8408), .A2(n6839), .ZN(n6245) );
  OR2_X1 U7810 ( .A1(n8408), .A2(n6839), .ZN(n6244) );
  MUX2_X1 U7811 ( .A(n6245), .B(n6244), .S(n8420), .Z(n6246) );
  NAND3_X1 U7812 ( .A1(n6247), .A2(n6781), .A3(n6246), .ZN(n6265) );
  NOR2_X1 U7813 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n6248) );
  NAND2_X1 U7814 ( .A1(n6249), .A2(n6248), .ZN(n6250) );
  OAI21_X1 U7815 ( .B1(n6251), .B2(n6250), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6252) );
  XNOR2_X1 U7816 ( .A(n6252), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8239) );
  AOI22_X1 U7817 ( .A1(n6332), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6853), .B2(
        n8239), .ZN(n6253) );
  NAND2_X1 U7818 ( .A1(n6048), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6259) );
  NAND2_X1 U7819 ( .A1(n4460), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6258) );
  XNOR2_X1 U7820 ( .A(n6255), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n8386) );
  NAND2_X1 U7821 ( .A1(n6018), .A2(n8386), .ZN(n6257) );
  NAND2_X1 U7822 ( .A1(n4461), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6256) );
  NAND2_X1 U7823 ( .A1(n8034), .A2(n8368), .ZN(n8370) );
  AND2_X1 U7824 ( .A1(n8511), .A2(n8405), .ZN(n6426) );
  INV_X1 U7825 ( .A(n6426), .ZN(n6260) );
  NAND2_X1 U7826 ( .A1(n8370), .A2(n6260), .ZN(n6262) );
  OAI21_X1 U7827 ( .B1(n8405), .B2(n8511), .A(n6458), .ZN(n6261) );
  MUX2_X1 U7828 ( .A(n6262), .B(n6261), .S(n6839), .Z(n6263) );
  INV_X1 U7829 ( .A(n6263), .ZN(n6264) );
  NAND2_X1 U7830 ( .A1(n6265), .A2(n6264), .ZN(n6289) );
  NAND2_X1 U7831 ( .A1(n7356), .A2(n6387), .ZN(n6269) );
  NAND2_X1 U7832 ( .A1(n6266), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6267) );
  XNOR2_X1 U7833 ( .A(n6267), .B(n5030), .ZN(n8247) );
  INV_X1 U7834 ( .A(n8247), .ZN(n6830) );
  AOI22_X1 U7835 ( .A1(n6332), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6830), .B2(
        n6853), .ZN(n6268) );
  INV_X1 U7836 ( .A(n8864), .ZN(n6782) );
  NAND2_X1 U7837 ( .A1(n6346), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6276) );
  NAND2_X1 U7838 ( .A1(n6048), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6275) );
  INV_X1 U7839 ( .A(n6270), .ZN(n6271) );
  NAND2_X1 U7840 ( .A1(n6271), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6272) );
  NAND2_X1 U7841 ( .A1(n6279), .A2(n6272), .ZN(n8375) );
  NAND2_X1 U7842 ( .A1(n6018), .A2(n8375), .ZN(n6274) );
  NAND2_X1 U7843 ( .A1(n4462), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6273) );
  NAND2_X1 U7844 ( .A1(n6782), .A2(n8383), .ZN(n6290) );
  NAND2_X1 U7845 ( .A1(n6290), .A2(n8370), .ZN(n6429) );
  NAND2_X1 U7846 ( .A1(n6289), .A2(n4826), .ZN(n6286) );
  NAND2_X1 U7847 ( .A1(n7430), .A2(n6387), .ZN(n6278) );
  OR2_X1 U7848 ( .A1(n6037), .A2(n8625), .ZN(n6277) );
  NAND2_X1 U7849 ( .A1(n4460), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U7850 ( .A1(n6048), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6284) );
  NAND2_X1 U7851 ( .A1(n6279), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6280) );
  NAND2_X1 U7852 ( .A1(n6281), .A2(n6280), .ZN(n8361) );
  NAND2_X1 U7853 ( .A1(n6018), .A2(n8361), .ZN(n6283) );
  NAND2_X1 U7854 ( .A1(n4462), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6282) );
  OR2_X1 U7855 ( .A1(n6782), .A2(n8383), .ZN(n6428) );
  NAND3_X1 U7856 ( .A1(n6286), .A2(n6457), .A3(n6428), .ZN(n6287) );
  NAND2_X1 U7857 ( .A1(n8499), .A2(n8369), .ZN(n8345) );
  AND4_X1 U7858 ( .A1(n6455), .A2(n6287), .A3(n6839), .A4(n8345), .ZN(n6288)
         );
  OR2_X1 U7859 ( .A1(n8335), .A2(n6288), .ZN(n6294) );
  NAND3_X1 U7860 ( .A1(n6289), .A2(n6458), .A3(n6428), .ZN(n6291) );
  MUX2_X1 U7861 ( .A(n4819), .B(n6292), .S(n6851), .Z(n6293) );
  NAND2_X1 U7862 ( .A1(n6434), .A2(n6432), .ZN(n6296) );
  OR2_X1 U7863 ( .A1(n6453), .A2(n4817), .ZN(n6295) );
  MUX2_X1 U7864 ( .A(n6296), .B(n6295), .S(n6839), .Z(n6297) );
  NAND3_X1 U7865 ( .A1(n6299), .A2(n8306), .A3(n6298), .ZN(n6310) );
  MUX2_X1 U7866 ( .A(n6437), .B(n6439), .S(n6851), .Z(n6309) );
  NAND2_X1 U7867 ( .A1(n8887), .A2(n6387), .ZN(n6301) );
  NAND2_X1 U7868 ( .A1(n6332), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6300) );
  NAND2_X1 U7869 ( .A1(n6302), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6303) );
  NAND2_X1 U7870 ( .A1(n6315), .A2(n6303), .ZN(n8292) );
  NAND2_X1 U7871 ( .A1(n8292), .A2(n6018), .ZN(n6308) );
  INV_X1 U7872 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8293) );
  NAND2_X1 U7873 ( .A1(n6048), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6305) );
  NAND2_X1 U7874 ( .A1(n6346), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6304) );
  OAI211_X1 U7875 ( .C1(n6349), .C2(n8293), .A(n6305), .B(n6304), .ZN(n6306)
         );
  INV_X1 U7876 ( .A(n6306), .ZN(n6307) );
  INV_X1 U7877 ( .A(n6441), .ZN(n6323) );
  AOI21_X1 U7878 ( .B1(n6310), .B2(n6309), .A(n8296), .ZN(n6343) );
  NAND2_X1 U7879 ( .A1(n7823), .A2(n6387), .ZN(n6312) );
  NAND2_X1 U7880 ( .A1(n6332), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6311) );
  INV_X1 U7881 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6313) );
  NAND2_X1 U7882 ( .A1(n6315), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6316) );
  NAND2_X1 U7883 ( .A1(n6344), .A2(n6316), .ZN(n8284) );
  NAND2_X1 U7884 ( .A1(n8284), .A2(n6018), .ZN(n6321) );
  INV_X1 U7885 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8528) );
  NAND2_X1 U7886 ( .A1(n4461), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6318) );
  NAND2_X1 U7887 ( .A1(n6048), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6317) );
  OAI211_X1 U7888 ( .C1(n6366), .C2(n8528), .A(n6318), .B(n6317), .ZN(n6319)
         );
  INV_X1 U7889 ( .A(n6319), .ZN(n6320) );
  NAND2_X1 U7890 ( .A1(n6322), .A2(n8267), .ZN(n6340) );
  MUX2_X1 U7891 ( .A(n6323), .B(n6440), .S(n6851), .Z(n6324) );
  OR2_X1 U7892 ( .A1(n8282), .A2(n6324), .ZN(n6342) );
  INV_X1 U7893 ( .A(n6327), .ZN(n6329) );
  NAND2_X1 U7894 ( .A1(n6329), .A2(n6328), .ZN(n6330) );
  INV_X1 U7895 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7813) );
  INV_X1 U7896 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9558) );
  MUX2_X1 U7897 ( .A(n7813), .B(n9558), .S(n6857), .Z(n6355) );
  NAND2_X1 U7898 ( .A1(n7812), .A2(n6387), .ZN(n6334) );
  NAND2_X1 U7899 ( .A1(n6332), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6333) );
  INV_X1 U7900 ( .A(n7819), .ZN(n6335) );
  NAND2_X1 U7901 ( .A1(n6335), .A2(n6018), .ZN(n6395) );
  INV_X1 U7902 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8733) );
  NAND2_X1 U7903 ( .A1(n6048), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6337) );
  NAND2_X1 U7904 ( .A1(n4460), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6336) );
  OAI211_X1 U7905 ( .C1(n8733), .C2(n6349), .A(n6337), .B(n6336), .ZN(n6338)
         );
  INV_X1 U7906 ( .A(n6338), .ZN(n6339) );
  NAND2_X1 U7907 ( .A1(n6825), .A2(n8268), .ZN(n6371) );
  INV_X2 U7908 ( .A(n6793), .ZN(n6751) );
  MUX2_X1 U7909 ( .A(n6340), .B(n6442), .S(n6839), .Z(n6341) );
  OAI211_X1 U7910 ( .C1(n6343), .C2(n6342), .A(n6751), .B(n6341), .ZN(n6373)
         );
  NAND2_X1 U7911 ( .A1(n6344), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6345) );
  NAND2_X1 U7912 ( .A1(n7819), .A2(n6345), .ZN(n7925) );
  NAND2_X1 U7913 ( .A1(n7925), .A2(n6018), .ZN(n6352) );
  INV_X1 U7914 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8271) );
  NAND2_X1 U7915 ( .A1(n6048), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6348) );
  NAND2_X1 U7916 ( .A1(n6346), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6347) );
  OAI211_X1 U7917 ( .C1(n6349), .C2(n8271), .A(n6348), .B(n6347), .ZN(n6350)
         );
  INV_X1 U7918 ( .A(n6350), .ZN(n6351) );
  NAND2_X1 U7919 ( .A1(n9559), .A2(n6387), .ZN(n6354) );
  INV_X1 U7920 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8882) );
  OR2_X1 U7921 ( .A1(n6037), .A2(n8882), .ZN(n6353) );
  MUX2_X1 U7922 ( .A(n8281), .B(n8526), .S(n6839), .Z(n6374) );
  NAND2_X1 U7923 ( .A1(n6356), .A2(n6355), .ZN(n6357) );
  INV_X1 U7924 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7826) );
  INV_X1 U7925 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8690) );
  MUX2_X1 U7926 ( .A(n7826), .B(n8690), .S(n6857), .Z(n6359) );
  INV_X1 U7927 ( .A(SI_30_), .ZN(n8816) );
  NAND2_X1 U7928 ( .A1(n6359), .A2(n8816), .ZN(n6381) );
  INV_X1 U7929 ( .A(n6359), .ZN(n6360) );
  NAND2_X1 U7930 ( .A1(n6360), .A2(SI_30_), .ZN(n6361) );
  AND2_X1 U7931 ( .A1(n6381), .A2(n6361), .ZN(n6379) );
  NOR2_X1 U7932 ( .A1(n6037), .A2(n7826), .ZN(n6362) );
  INV_X1 U7933 ( .A(n6444), .ZN(n6370) );
  INV_X1 U7934 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6365) );
  NAND2_X1 U7935 ( .A1(n6048), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6364) );
  NAND2_X1 U7936 ( .A1(n4461), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6363) );
  OAI211_X1 U7937 ( .C1(n6366), .C2(n6365), .A(n6364), .B(n6363), .ZN(n6367)
         );
  INV_X1 U7938 ( .A(n6367), .ZN(n6368) );
  NAND2_X1 U7939 ( .A1(n6395), .A2(n6368), .ZN(n8072) );
  INV_X1 U7940 ( .A(n8072), .ZN(n6369) );
  NAND2_X1 U7941 ( .A1(n6370), .A2(n6369), .ZN(n6396) );
  NAND2_X1 U7942 ( .A1(n6396), .A2(n6371), .ZN(n6446) );
  AND2_X1 U7943 ( .A1(n6444), .A2(n8072), .ZN(n6450) );
  INV_X1 U7944 ( .A(n6450), .ZN(n6398) );
  NAND2_X1 U7945 ( .A1(n6398), .A2(n6443), .ZN(n6482) );
  MUX2_X1 U7946 ( .A(n6446), .B(n6482), .S(n6851), .Z(n6372) );
  OAI21_X1 U7947 ( .B1(n6374), .B2(n6793), .A(n6373), .ZN(n6376) );
  MUX2_X1 U7948 ( .A(n8281), .B(n8526), .S(n6851), .Z(n6375) );
  NAND2_X1 U7949 ( .A1(n6380), .A2(n6379), .ZN(n6382) );
  MUX2_X1 U7950 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n6857), .Z(n6384) );
  INV_X1 U7951 ( .A(SI_31_), .ZN(n6383) );
  XNOR2_X1 U7952 ( .A(n6384), .B(n6383), .ZN(n6385) );
  NAND2_X1 U7953 ( .A1(n8875), .A2(n6387), .ZN(n6390) );
  INV_X1 U7954 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6388) );
  OR2_X1 U7955 ( .A1(n6037), .A2(n6388), .ZN(n6389) );
  NAND2_X1 U7956 ( .A1(n4460), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6393) );
  NAND2_X1 U7957 ( .A1(n6048), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6392) );
  NAND2_X1 U7958 ( .A1(n4462), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6391) );
  AND3_X1 U7959 ( .A1(n6393), .A2(n6392), .A3(n6391), .ZN(n6394) );
  OR2_X1 U7960 ( .A1(n6449), .A2(n7814), .ZN(n6448) );
  INV_X1 U7961 ( .A(n6396), .ZN(n6397) );
  AOI21_X1 U7962 ( .B1(n6839), .B2(n6398), .A(n6397), .ZN(n6399) );
  NAND2_X1 U7963 ( .A1(n6449), .A2(n7814), .ZN(n6484) );
  NAND2_X1 U7964 ( .A1(n4495), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6403) );
  MUX2_X1 U7965 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6403), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n6404) );
  NAND2_X1 U7966 ( .A1(n6404), .A2(n5963), .ZN(n7431) );
  INV_X1 U7967 ( .A(n7431), .ZN(n6831) );
  INV_X1 U7968 ( .A(n10156), .ZN(n6408) );
  NAND2_X1 U7969 ( .A1(n7198), .A2(n7199), .ZN(n6412) );
  NAND2_X1 U7970 ( .A1(n6412), .A2(n6411), .ZN(n7391) );
  NAND2_X1 U7971 ( .A1(n7391), .A2(n6464), .ZN(n6413) );
  NAND2_X1 U7972 ( .A1(n6413), .A2(n6465), .ZN(n7405) );
  NAND2_X1 U7973 ( .A1(n7521), .A2(n6416), .ZN(n6417) );
  NAND2_X1 U7974 ( .A1(n6417), .A2(n6470), .ZN(n7570) );
  NAND2_X1 U7975 ( .A1(n7715), .A2(n6418), .ZN(n7573) );
  NAND2_X1 U7976 ( .A1(n6420), .A2(n6462), .ZN(n7705) );
  NAND2_X1 U7977 ( .A1(n7705), .A2(n6459), .ZN(n6422) );
  OR2_X1 U7978 ( .A1(n7939), .A2(n8454), .ZN(n6421) );
  NOR2_X1 U7979 ( .A1(n9636), .A2(n7841), .ZN(n6423) );
  INV_X1 U7980 ( .A(n6458), .ZN(n6427) );
  INV_X1 U7981 ( .A(n6457), .ZN(n6430) );
  NAND2_X1 U7982 ( .A1(n6455), .A2(n8345), .ZN(n6431) );
  INV_X1 U7983 ( .A(n6437), .ZN(n6438) );
  INV_X1 U7984 ( .A(n6443), .ZN(n6445) );
  OAI22_X1 U7985 ( .A1(n6752), .A2(n6445), .B1(n7822), .B2(n6449), .ZN(n6452)
         );
  INV_X1 U7986 ( .A(n6446), .ZN(n6447) );
  NAND2_X1 U7987 ( .A1(n6448), .A2(n6447), .ZN(n6483) );
  NOR2_X1 U7988 ( .A1(n6450), .A2(n7814), .ZN(n6451) );
  OAI22_X1 U7989 ( .A1(n6452), .A2(n6483), .B1(n8522), .B2(n6451), .ZN(n6489)
         );
  NOR2_X1 U7990 ( .A1(n6454), .A2(n6453), .ZN(n8323) );
  NAND2_X1 U7991 ( .A1(n6457), .A2(n8345), .ZN(n8359) );
  XNOR2_X1 U7992 ( .A(n8864), .B(n8356), .ZN(n8373) );
  INV_X1 U7993 ( .A(n6459), .ZN(n7706) );
  INV_X1 U7994 ( .A(n6460), .ZN(n8459) );
  INV_X1 U7995 ( .A(n7834), .ZN(n6473) );
  XNOR2_X1 U7996 ( .A(n8085), .B(n8040), .ZN(n7406) );
  AND2_X1 U7997 ( .A1(n7169), .A2(n6463), .ZN(n7186) );
  INV_X1 U7998 ( .A(n7199), .ZN(n6466) );
  NAND2_X1 U7999 ( .A1(n6465), .A2(n6464), .ZN(n7389) );
  NOR4_X1 U8000 ( .A1(n6466), .A2(n10156), .A3(n7170), .A4(n7389), .ZN(n6468)
         );
  NAND3_X1 U8001 ( .A1(n7186), .A2(n6468), .A3(n6467), .ZN(n6471) );
  NAND2_X1 U8002 ( .A1(n6470), .A2(n6469), .ZN(n7522) );
  NOR4_X1 U8003 ( .A1(n4776), .A2(n7406), .A3(n6471), .A4(n7522), .ZN(n6472)
         );
  NAND4_X1 U8004 ( .A1(n6475), .A2(n6474), .A3(n6473), .A4(n6472), .ZN(n6476)
         );
  NOR4_X1 U8005 ( .A1(n8444), .A2(n7706), .A3(n8459), .A4(n6476), .ZN(n6477)
         );
  NAND4_X1 U8006 ( .A1(n8385), .A2(n8415), .A3(n6477), .A4(n8406), .ZN(n6478)
         );
  NOR4_X1 U8007 ( .A1(n8359), .A2(n5012), .A3(n8373), .A4(n6478), .ZN(n6479)
         );
  NAND4_X1 U8008 ( .A1(n8323), .A2(n4982), .A3(n8349), .A4(n6479), .ZN(n6480)
         );
  NOR4_X1 U8009 ( .A1(n6482), .A2(n8273), .A3(n8282), .A4(n6481), .ZN(n6486)
         );
  INV_X1 U8010 ( .A(n6483), .ZN(n6485) );
  XNOR2_X1 U8011 ( .A(n6492), .B(n8247), .ZN(n6513) );
  XNOR2_X1 U8012 ( .A(n6495), .B(n6494), .ZN(n6850) );
  OR2_X1 U8013 ( .A1(n6850), .A2(P2_U3151), .ZN(n7642) );
  NAND2_X1 U8014 ( .A1(n6495), .A2(n6494), .ZN(n6496) );
  NAND2_X1 U8015 ( .A1(n6500), .A2(n6499), .ZN(n6502) );
  INV_X1 U8016 ( .A(n6802), .ZN(n6508) );
  OR2_X1 U8017 ( .A1(n6500), .A2(n6499), .ZN(n6501) );
  NAND2_X1 U8018 ( .A1(n6502), .A2(n6501), .ZN(n6801) );
  INV_X1 U8019 ( .A(n6504), .ZN(n6505) );
  NOR2_X1 U8020 ( .A1(n6801), .A2(n6808), .ZN(n6507) );
  NAND2_X1 U8021 ( .A1(n6508), .A2(n6507), .ZN(n7004) );
  INV_X1 U8022 ( .A(n7164), .ZN(n6838) );
  NOR4_X1 U8023 ( .A1(n6838), .A2(n6755), .A3(n7054), .A4(n7183), .ZN(n6511)
         );
  OAI21_X1 U8024 ( .B1(n7642), .B2(n6833), .A(P2_B_REG_SCAN_IN), .ZN(n6510) );
  OAI21_X1 U8025 ( .B1(n6513), .B2(n7642), .A(n6512), .ZN(P2_U3296) );
  INV_X1 U8026 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6514) );
  NOR2_X1 U8027 ( .A1(n4456), .A2(n6514), .ZN(n6515) );
  INV_X1 U8028 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n6518) );
  NAND2_X1 U8029 ( .A1(n6584), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6517) );
  NAND2_X1 U8030 ( .A1(n6585), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6516) );
  OAI211_X1 U8031 ( .C1(n5247), .C2(n6518), .A(n6517), .B(n6516), .ZN(n9196)
         );
  INV_X1 U8032 ( .A(n9196), .ZN(n6627) );
  NOR2_X1 U8033 ( .A1(n9437), .A2(n6627), .ZN(n6590) );
  AND2_X1 U8034 ( .A1(n7544), .A2(n4722), .ZN(n6972) );
  INV_X1 U8035 ( .A(n6520), .ZN(n6647) );
  INV_X1 U8036 ( .A(n6644), .ZN(n6519) );
  INV_X1 U8037 ( .A(n9236), .ZN(n9198) );
  AOI21_X1 U8038 ( .B1(n6647), .B2(n6519), .A(n9193), .ZN(n6575) );
  INV_X1 U8039 ( .A(n6972), .ZN(n6589) );
  OR2_X1 U8040 ( .A1(n9244), .A2(n9455), .ZN(n6643) );
  OR2_X1 U8041 ( .A1(n9259), .A2(n9462), .ZN(n6635) );
  NAND2_X1 U8042 ( .A1(n6643), .A2(n6635), .ZN(n6570) );
  NAND2_X1 U8043 ( .A1(n9259), .A2(n9462), .ZN(n6641) );
  NAND2_X1 U8044 ( .A1(n9244), .A2(n9455), .ZN(n6571) );
  OAI21_X1 U8045 ( .B1(n6570), .B2(n6641), .A(n6571), .ZN(n6522) );
  NAND3_X1 U8046 ( .A1(n6570), .A2(n6972), .A3(n6571), .ZN(n6521) );
  INV_X1 U8047 ( .A(n9500), .ZN(n9339) );
  AND2_X1 U8048 ( .A1(n9339), .A2(n9351), .ZN(n6726) );
  INV_X1 U8049 ( .A(n9507), .ZN(n9159) );
  AND2_X1 U8050 ( .A1(n9159), .A2(n9369), .ZN(n6619) );
  NOR2_X1 U8051 ( .A1(n9426), .A2(n9152), .ZN(n6549) );
  NAND2_X1 U8052 ( .A1(n9520), .A2(n9421), .ZN(n6712) );
  INV_X1 U8053 ( .A(n9421), .ZN(n9388) );
  NAND2_X1 U8054 ( .A1(n9880), .A2(n9885), .ZN(n6524) );
  OR2_X1 U8055 ( .A1(n9920), .A2(n9065), .ZN(n6523) );
  NAND2_X1 U8056 ( .A1(n9930), .A2(n9934), .ZN(n6690) );
  AND2_X1 U8057 ( .A1(n6525), .A2(n6690), .ZN(n7306) );
  XNOR2_X1 U8058 ( .A(n7311), .B(n9063), .ZN(n7316) );
  OR2_X1 U8059 ( .A1(n7311), .A2(n9063), .ZN(n6526) );
  NOR2_X1 U8060 ( .A1(n9943), .A2(n9863), .ZN(n6607) );
  NAND2_X1 U8061 ( .A1(n9943), .A2(n9863), .ZN(n6689) );
  NAND2_X1 U8062 ( .A1(n9953), .A2(n9062), .ZN(n6691) );
  OR2_X1 U8063 ( .A1(n9953), .A2(n9062), .ZN(n6527) );
  AND2_X1 U8064 ( .A1(n6691), .A2(n6527), .ZN(n9861) );
  NAND2_X1 U8065 ( .A1(n9860), .A2(n6691), .ZN(n7331) );
  NAND2_X1 U8066 ( .A1(n7424), .A2(n7411), .ZN(n7329) );
  NAND2_X1 U8067 ( .A1(n7331), .A2(n7329), .ZN(n6650) );
  INV_X1 U8068 ( .A(n7411), .ZN(n7371) );
  INV_X1 U8069 ( .A(n7424), .ZN(n9865) );
  NAND2_X1 U8070 ( .A1(n7371), .A2(n9865), .ZN(n7330) );
  NAND2_X1 U8071 ( .A1(n6650), .A2(n7330), .ZN(n7377) );
  NOR2_X1 U8072 ( .A1(n7456), .A2(n7552), .ZN(n7375) );
  NAND2_X1 U8073 ( .A1(n7470), .A2(n7647), .ZN(n7459) );
  AND2_X1 U8074 ( .A1(n7459), .A2(n7374), .ZN(n6687) );
  OR2_X1 U8075 ( .A1(n7470), .A2(n7647), .ZN(n7500) );
  AOI21_X1 U8076 ( .B1(n6528), .B2(n7500), .A(n7486), .ZN(n6529) );
  MUX2_X1 U8077 ( .A(n6529), .B(n6528), .S(n6589), .Z(n6535) );
  INV_X1 U8078 ( .A(n9972), .ZN(n7654) );
  INV_X1 U8079 ( .A(n8926), .ZN(n9979) );
  AND2_X1 U8080 ( .A1(n7654), .A2(n9979), .ZN(n7487) );
  NAND2_X1 U8081 ( .A1(n9980), .A2(n9845), .ZN(n9841) );
  OAI21_X1 U8082 ( .B1(n6535), .B2(n7487), .A(n9841), .ZN(n6532) );
  AND2_X1 U8083 ( .A1(n6530), .A2(n9995), .ZN(n6539) );
  INV_X1 U8084 ( .A(n9980), .ZN(n7586) );
  INV_X1 U8085 ( .A(n9845), .ZN(n9060) );
  AND2_X1 U8086 ( .A1(n7586), .A2(n9060), .ZN(n6533) );
  NOR2_X1 U8087 ( .A1(n6539), .A2(n6533), .ZN(n6531) );
  AND2_X1 U8088 ( .A1(n9988), .A2(n7740), .ZN(n6536) );
  NOR2_X1 U8089 ( .A1(n9998), .A2(n9844), .ZN(n6538) );
  INV_X1 U8090 ( .A(n7487), .ZN(n6606) );
  NAND2_X1 U8091 ( .A1(n6606), .A2(n7500), .ZN(n6534) );
  INV_X1 U8092 ( .A(n7486), .ZN(n6651) );
  NAND2_X1 U8093 ( .A1(n6534), .A2(n6651), .ZN(n6699) );
  NAND3_X1 U8094 ( .A1(n6535), .A2(n6702), .A3(n6699), .ZN(n6540) );
  INV_X1 U8095 ( .A(n6536), .ZN(n6602) );
  NAND2_X1 U8096 ( .A1(n6602), .A2(n9841), .ZN(n6655) );
  AND2_X1 U8097 ( .A1(n6702), .A2(n7486), .ZN(n6537) );
  NOR2_X1 U8098 ( .A1(n6655), .A2(n6537), .ZN(n6704) );
  INV_X1 U8099 ( .A(n6538), .ZN(n6603) );
  OR2_X1 U8100 ( .A1(n9001), .A2(n8909), .ZN(n6601) );
  NAND2_X1 U8101 ( .A1(n6660), .A2(n6601), .ZN(n6709) );
  INV_X1 U8102 ( .A(n6709), .ZN(n6542) );
  NAND2_X1 U8103 ( .A1(n9426), .A2(n9152), .ZN(n6663) );
  NAND2_X1 U8104 ( .A1(n6712), .A2(n6663), .ZN(n6552) );
  AND2_X1 U8105 ( .A1(n9524), .A2(n9422), .ZN(n6547) );
  NAND2_X1 U8106 ( .A1(n9001), .A2(n8909), .ZN(n6659) );
  NOR2_X1 U8107 ( .A1(n6709), .A2(n6659), .ZN(n6541) );
  OR3_X1 U8108 ( .A1(n6552), .A2(n6547), .A3(n6541), .ZN(n6711) );
  AOI21_X1 U8109 ( .B1(n6545), .B2(n6542), .A(n6711), .ZN(n6543) );
  AOI211_X1 U8110 ( .C1(n6549), .C2(n6712), .A(n6544), .B(n6543), .ZN(n6553)
         );
  OAI21_X1 U8111 ( .B1(n6546), .B2(n4688), .A(n6601), .ZN(n6551) );
  INV_X1 U8112 ( .A(n6547), .ZN(n6548) );
  INV_X1 U8113 ( .A(n6660), .ZN(n6550) );
  INV_X1 U8114 ( .A(n6549), .ZN(n6600) );
  NAND2_X1 U8115 ( .A1(n6599), .A2(n6600), .ZN(n6713) );
  XNOR2_X1 U8116 ( .A(n9385), .B(n9376), .ZN(n9386) );
  INV_X1 U8117 ( .A(n9506), .ZN(n9358) );
  OR2_X1 U8118 ( .A1(n9514), .A2(n9358), .ZN(n6721) );
  OR2_X1 U8119 ( .A1(n9385), .A2(n9376), .ZN(n6666) );
  NAND2_X1 U8120 ( .A1(n6721), .A2(n6666), .ZN(n6716) );
  INV_X1 U8121 ( .A(n9369), .ZN(n9158) );
  NAND2_X1 U8122 ( .A1(n9507), .A2(n9158), .ZN(n6723) );
  NAND2_X1 U8123 ( .A1(n9514), .A2(n9358), .ZN(n6667) );
  OAI211_X1 U8124 ( .C1(n6559), .C2(n6716), .A(n6723), .B(n6667), .ZN(n6556)
         );
  INV_X1 U8125 ( .A(n9351), .ZN(n9324) );
  AND2_X1 U8126 ( .A1(n9500), .A2(n9324), .ZN(n6561) );
  INV_X1 U8127 ( .A(n6723), .ZN(n6554) );
  NOR2_X1 U8128 ( .A1(n6561), .A2(n6554), .ZN(n6555) );
  NAND2_X1 U8129 ( .A1(n9385), .A2(n9376), .ZN(n6664) );
  NAND2_X1 U8130 ( .A1(n6667), .A2(n6664), .ZN(n6717) );
  INV_X1 U8131 ( .A(n6721), .ZN(n6557) );
  NOR3_X1 U8132 ( .A1(n6619), .A2(n6972), .A3(n6557), .ZN(n6558) );
  NAND2_X1 U8133 ( .A1(n9497), .A2(n9488), .ZN(n6621) );
  AND2_X1 U8134 ( .A1(n6621), .A2(n9319), .ZN(n6637) );
  NOR2_X1 U8135 ( .A1(n6727), .A2(n6726), .ZN(n6562) );
  MUX2_X1 U8136 ( .A(n6637), .B(n6562), .S(n6589), .Z(n6563) );
  MUX2_X1 U8137 ( .A(n6670), .B(n6621), .S(n6589), .Z(n6564) );
  OR2_X1 U8138 ( .A1(n9304), .A2(n9481), .ZN(n9287) );
  NAND2_X1 U8139 ( .A1(n9304), .A2(n9481), .ZN(n6565) );
  NAND2_X1 U8140 ( .A1(n9287), .A2(n6565), .ZN(n9309) );
  OR2_X1 U8141 ( .A1(n9299), .A2(n9315), .ZN(n6623) );
  NAND2_X1 U8142 ( .A1(n6623), .A2(n9287), .ZN(n6631) );
  NAND2_X1 U8143 ( .A1(n9299), .A2(n9315), .ZN(n9186) );
  OAI21_X1 U8144 ( .B1(n6566), .B2(n6631), .A(n9186), .ZN(n6568) );
  NAND2_X1 U8145 ( .A1(n9186), .A2(n6565), .ZN(n6636) );
  OAI21_X1 U8146 ( .B1(n6566), .B2(n6636), .A(n6623), .ZN(n6567) );
  NAND2_X1 U8147 ( .A1(n9478), .A2(n9469), .ZN(n6640) );
  NAND2_X1 U8148 ( .A1(n9188), .A2(n6640), .ZN(n9187) );
  MUX2_X1 U8149 ( .A(n6640), .B(n9188), .S(n6972), .Z(n6569) );
  INV_X1 U8150 ( .A(n6570), .ZN(n6573) );
  INV_X1 U8151 ( .A(n6571), .ZN(n9190) );
  INV_X1 U8152 ( .A(n6641), .ZN(n9189) );
  NOR2_X1 U8153 ( .A1(n9190), .A2(n9189), .ZN(n6572) );
  OAI21_X1 U8154 ( .B1(n6972), .B2(n6575), .A(n6574), .ZN(n6580) );
  NOR2_X1 U8155 ( .A1(n6581), .A2(n9558), .ZN(n6576) );
  AND2_X1 U8156 ( .A1(n9205), .A2(n9210), .ZN(n6577) );
  MUX2_X1 U8157 ( .A(n6578), .B(n6577), .S(n6589), .Z(n6579) );
  NOR2_X1 U8158 ( .A1(n6581), .A2(n8690), .ZN(n6582) );
  INV_X1 U8159 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n8669) );
  NAND2_X1 U8160 ( .A1(n6584), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6587) );
  NAND2_X1 U8161 ( .A1(n6585), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6586) );
  OAI211_X1 U8162 ( .C1(n5247), .C2(n8669), .A(n6587), .B(n6586), .ZN(n9140)
         );
  INV_X1 U8163 ( .A(n9140), .ZN(n6672) );
  AOI21_X1 U8164 ( .B1(n6738), .B2(n4722), .A(n6743), .ZN(n6591) );
  INV_X1 U8165 ( .A(n6592), .ZN(n6596) );
  NAND2_X1 U8166 ( .A1(n6593), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7657) );
  INV_X1 U8167 ( .A(n7657), .ZN(n6595) );
  INV_X1 U8168 ( .A(n6974), .ZN(n6594) );
  NAND3_X1 U8169 ( .A1(n6596), .A2(n6595), .A3(n6594), .ZN(n6750) );
  OAI21_X1 U8170 ( .B1(n6597), .B2(n7544), .A(n6692), .ZN(n6629) );
  INV_X1 U8171 ( .A(n6598), .ZN(n6679) );
  INV_X1 U8172 ( .A(n9440), .ZN(n9148) );
  OR2_X1 U8173 ( .A1(n9148), .A2(n6627), .ZN(n6676) );
  NAND2_X1 U8174 ( .A1(n6679), .A2(n6676), .ZN(n6736) );
  NAND2_X1 U8175 ( .A1(n6721), .A2(n6667), .ZN(n9364) );
  NAND2_X1 U8176 ( .A1(n6599), .A2(n6712), .ZN(n9400) );
  NAND2_X1 U8177 ( .A1(n6600), .A2(n6663), .ZN(n9424) );
  INV_X1 U8178 ( .A(n6706), .ZN(n6657) );
  NAND2_X1 U8179 ( .A1(n6603), .A2(n6657), .ZN(n7691) );
  NAND2_X1 U8180 ( .A1(n6702), .A2(n9841), .ZN(n7587) );
  INV_X1 U8181 ( .A(n7375), .ZN(n6604) );
  AND3_X1 U8182 ( .A1(n7500), .A2(n6604), .A3(n7330), .ZN(n6605) );
  NAND2_X1 U8183 ( .A1(n6606), .A2(n6605), .ZN(n6649) );
  NAND2_X1 U8184 ( .A1(n4493), .A2(n6690), .ZN(n7291) );
  INV_X1 U8185 ( .A(n6607), .ZN(n6608) );
  NAND2_X1 U8186 ( .A1(n6608), .A2(n6689), .ZN(n7334) );
  NOR2_X1 U8187 ( .A1(n7291), .A2(n7334), .ZN(n6611) );
  INV_X1 U8188 ( .A(n9880), .ZN(n6609) );
  NAND2_X1 U8189 ( .A1(n7274), .A2(n9901), .ZN(n6694) );
  AND2_X1 U8190 ( .A1(n6609), .A2(n6694), .ZN(n7232) );
  INV_X1 U8191 ( .A(n9861), .ZN(n9873) );
  NOR2_X1 U8192 ( .A1(n9873), .A2(n6692), .ZN(n6610) );
  NAND4_X1 U8193 ( .A1(n6611), .A2(n7232), .A3(n6610), .A4(n7329), .ZN(n6613)
         );
  INV_X1 U8194 ( .A(n7316), .ZN(n7305) );
  NAND2_X1 U8195 ( .A1(n7305), .A2(n9885), .ZN(n6612) );
  NOR2_X1 U8196 ( .A1(n6613), .A2(n6612), .ZN(n6614) );
  NAND3_X1 U8197 ( .A1(n6651), .A2(n6687), .A3(n6614), .ZN(n6615) );
  OR3_X1 U8198 ( .A1(n7587), .A2(n6649), .A3(n6615), .ZN(n6616) );
  NOR2_X1 U8199 ( .A1(n7691), .A2(n6616), .ZN(n6617) );
  NAND4_X1 U8200 ( .A1(n7749), .A2(n7744), .A3(n9847), .A4(n6617), .ZN(n6618)
         );
  OR4_X1 U8201 ( .A1(n9364), .A2(n9400), .A3(n9424), .A4(n6618), .ZN(n6620) );
  NAND2_X1 U8202 ( .A1(n6669), .A2(n9319), .ZN(n9341) );
  INV_X1 U8203 ( .A(n6619), .ZN(n6720) );
  NAND2_X1 U8204 ( .A1(n6720), .A2(n6723), .ZN(n9347) );
  OR4_X1 U8205 ( .A1(n6620), .A2(n9386), .A3(n9341), .A4(n9347), .ZN(n6622) );
  NAND2_X1 U8206 ( .A1(n6670), .A2(n6621), .ZN(n9321) );
  OR3_X1 U8207 ( .A1(n9309), .A2(n6622), .A3(n9321), .ZN(n6624) );
  NAND2_X1 U8208 ( .A1(n6635), .A2(n6641), .ZN(n9266) );
  NAND2_X1 U8209 ( .A1(n6623), .A2(n9186), .ZN(n9290) );
  XNOR2_X1 U8210 ( .A(n9244), .B(n9455), .ZN(n9250) );
  OR3_X1 U8211 ( .A1(n6625), .A2(n9234), .A3(n9250), .ZN(n6626) );
  NOR2_X1 U8212 ( .A1(n9213), .A2(n6626), .ZN(n6628) );
  NAND2_X1 U8213 ( .A1(n9148), .A2(n6627), .ZN(n6675) );
  NOR2_X1 U8214 ( .A1(n7433), .A2(n7657), .ZN(n6683) );
  AND2_X1 U8215 ( .A1(n6630), .A2(n4887), .ZN(n6685) );
  NAND2_X1 U8216 ( .A1(n6631), .A2(n9186), .ZN(n6632) );
  NAND2_X1 U8217 ( .A1(n9188), .A2(n6632), .ZN(n6633) );
  NAND2_X1 U8218 ( .A1(n6633), .A2(n6640), .ZN(n6634) );
  NAND2_X1 U8219 ( .A1(n6635), .A2(n6634), .ZN(n6728) );
  INV_X1 U8220 ( .A(n6636), .ZN(n6639) );
  INV_X1 U8221 ( .A(n6637), .ZN(n6638) );
  NAND2_X1 U8222 ( .A1(n6638), .A2(n6670), .ZN(n9181) );
  AND3_X1 U8223 ( .A1(n6640), .A2(n6639), .A3(n9181), .ZN(n6642) );
  OAI21_X1 U8224 ( .B1(n6728), .B2(n6642), .A(n6641), .ZN(n6645) );
  AND2_X1 U8225 ( .A1(n6644), .A2(n6643), .ZN(n6648) );
  OAI21_X1 U8226 ( .B1(n9190), .B2(n6645), .A(n6648), .ZN(n6646) );
  AND2_X1 U8227 ( .A1(n6647), .A2(n6646), .ZN(n6686) );
  INV_X1 U8228 ( .A(n6648), .ZN(n6730) );
  INV_X1 U8229 ( .A(n6649), .ZN(n6698) );
  NAND2_X1 U8230 ( .A1(n6650), .A2(n6698), .ZN(n6701) );
  NAND3_X1 U8231 ( .A1(n6701), .A2(n6687), .A3(n6651), .ZN(n6652) );
  NAND2_X1 U8232 ( .A1(n6652), .A2(n6699), .ZN(n7489) );
  INV_X1 U8233 ( .A(n7489), .ZN(n6654) );
  INV_X1 U8234 ( .A(n7587), .ZN(n6653) );
  NAND2_X1 U8235 ( .A1(n6654), .A2(n6653), .ZN(n9842) );
  INV_X1 U8236 ( .A(n6655), .ZN(n6656) );
  NAND2_X1 U8237 ( .A1(n9842), .A2(n6656), .ZN(n7688) );
  NAND2_X1 U8238 ( .A1(n7688), .A2(n4503), .ZN(n6658) );
  NAND2_X1 U8239 ( .A1(n6658), .A2(n6657), .ZN(n7584) );
  NAND2_X1 U8240 ( .A1(n7584), .A2(n7744), .ZN(n7583) );
  INV_X1 U8241 ( .A(n7749), .ZN(n6661) );
  NAND2_X1 U8242 ( .A1(n9416), .A2(n6663), .ZN(n9407) );
  INV_X1 U8243 ( .A(n9400), .ZN(n9408) );
  NAND2_X1 U8244 ( .A1(n9407), .A2(n9408), .ZN(n9406) );
  INV_X1 U8245 ( .A(n6664), .ZN(n6665) );
  INV_X1 U8246 ( .A(n9364), .ZN(n9368) );
  NAND2_X1 U8247 ( .A1(n9366), .A2(n6667), .ZN(n9350) );
  INV_X1 U8248 ( .A(n9347), .ZN(n9349) );
  NAND2_X1 U8249 ( .A1(n9350), .A2(n9349), .ZN(n6668) );
  OR3_X1 U8250 ( .A1(n6730), .A2(n6728), .A3(n9180), .ZN(n6671) );
  NAND2_X1 U8251 ( .A1(n6686), .A2(n6671), .ZN(n6673) );
  AOI22_X1 U8252 ( .A1(n6685), .A2(n6673), .B1(n6672), .B2(n9148), .ZN(n6678)
         );
  INV_X1 U8253 ( .A(n6676), .ZN(n6677) );
  AOI22_X1 U8254 ( .A1(n6678), .A2(n6735), .B1(n6677), .B2(n9140), .ZN(n6680)
         );
  OAI211_X1 U8255 ( .C1(n6680), .C2(n6738), .A(n7279), .B(n6679), .ZN(n6682)
         );
  NAND2_X1 U8256 ( .A1(n6682), .A2(n6681), .ZN(n6684) );
  NAND3_X1 U8257 ( .A1(n6684), .A2(n6683), .A3(n9294), .ZN(n6749) );
  INV_X1 U8258 ( .A(n6685), .ZN(n6734) );
  INV_X1 U8259 ( .A(n6686), .ZN(n6732) );
  INV_X1 U8260 ( .A(n6687), .ZN(n7501) );
  NAND2_X1 U8261 ( .A1(n7311), .A2(n9063), .ZN(n6688) );
  NAND4_X1 U8262 ( .A1(n6691), .A2(n6690), .A3(n6689), .A4(n6688), .ZN(n6696)
         );
  NAND2_X1 U8263 ( .A1(n9920), .A2(n9065), .ZN(n6693) );
  NAND3_X1 U8264 ( .A1(n6694), .A2(n6693), .A3(n6692), .ZN(n6695) );
  NOR2_X1 U8265 ( .A1(n6696), .A2(n6695), .ZN(n6697) );
  AOI22_X1 U8266 ( .A1(n7501), .A2(n6699), .B1(n6698), .B2(n6697), .ZN(n6700)
         );
  NAND2_X1 U8267 ( .A1(n6701), .A2(n6700), .ZN(n6703) );
  NAND2_X1 U8268 ( .A1(n6703), .A2(n6702), .ZN(n6705) );
  NAND2_X1 U8269 ( .A1(n6705), .A2(n6704), .ZN(n6707) );
  AOI21_X1 U8270 ( .B1(n6707), .B2(n4503), .A(n6706), .ZN(n6708) );
  NOR2_X1 U8271 ( .A1(n6709), .A2(n6708), .ZN(n6710) );
  NOR2_X1 U8272 ( .A1(n6711), .A2(n6710), .ZN(n6715) );
  AND2_X1 U8273 ( .A1(n6713), .A2(n6712), .ZN(n6714) );
  OR3_X1 U8274 ( .A1(n6716), .A2(n6715), .A3(n6714), .ZN(n6719) );
  INV_X1 U8275 ( .A(n6717), .ZN(n6718) );
  NAND2_X1 U8276 ( .A1(n6719), .A2(n6718), .ZN(n6722) );
  NAND3_X1 U8277 ( .A1(n6722), .A2(n6721), .A3(n6720), .ZN(n6724) );
  AND2_X1 U8278 ( .A1(n6724), .A2(n6723), .ZN(n6725) );
  OR4_X1 U8279 ( .A1(n6728), .A2(n6727), .A3(n6726), .A4(n6725), .ZN(n6729) );
  NOR2_X1 U8280 ( .A1(n6730), .A2(n6729), .ZN(n6731) );
  NOR2_X1 U8281 ( .A1(n6732), .A2(n6731), .ZN(n6733) );
  OR2_X1 U8282 ( .A1(n6737), .A2(n6736), .ZN(n6739) );
  NAND3_X1 U8283 ( .A1(n6745), .A2(n6595), .A3(n6740), .ZN(n6748) );
  INV_X1 U8284 ( .A(n4459), .ZN(n6953) );
  AND2_X1 U8285 ( .A1(n9066), .A2(n6953), .ZN(n9069) );
  NAND3_X1 U8286 ( .A1(n7231), .A2(n9546), .A3(n9069), .ZN(n6742) );
  OAI211_X1 U8287 ( .C1(n6743), .C2(n7657), .A(n6742), .B(P1_B_REG_SCAN_IN), 
        .ZN(n6747) );
  INV_X1 U8288 ( .A(n6833), .ZN(n7542) );
  OAI211_X1 U8289 ( .C1(n6833), .C2(n7431), .A(n10225), .B(n8247), .ZN(n6753)
         );
  INV_X1 U8290 ( .A(n6753), .ZN(n6754) );
  NAND2_X1 U8291 ( .A1(n6754), .A2(n7183), .ZN(n10163) );
  XNOR2_X1 U8292 ( .A(n7054), .B(n8241), .ZN(n7001) );
  INV_X1 U8293 ( .A(n7001), .ZN(n7042) );
  AOI21_X1 U8294 ( .B1(P2_B_REG_SCAN_IN), .B2(n6756), .A(n10158), .ZN(n7815)
         );
  AOI22_X1 U8295 ( .A1(n8435), .A2(n8074), .B1(n8072), .B2(n7815), .ZN(n6800)
         );
  NAND2_X1 U8296 ( .A1(n6010), .A2(n7037), .ZN(n7154) );
  NAND2_X1 U8297 ( .A1(n7154), .A2(n7170), .ZN(n6759) );
  NAND2_X1 U8298 ( .A1(n6757), .A2(n7044), .ZN(n6758) );
  NAND2_X1 U8299 ( .A1(n6759), .A2(n6758), .ZN(n10155) );
  NAND2_X1 U8300 ( .A1(n10155), .A2(n10156), .ZN(n6761) );
  NAND2_X1 U8301 ( .A1(n7121), .A2(n10154), .ZN(n6760) );
  NOR2_X1 U8302 ( .A1(n8088), .A2(n10179), .ZN(n6763) );
  NAND2_X1 U8303 ( .A1(n8088), .A2(n10179), .ZN(n6762) );
  NOR2_X1 U8304 ( .A1(n8086), .A2(n7397), .ZN(n6767) );
  INV_X1 U8305 ( .A(n8085), .ZN(n7451) );
  NAND2_X1 U8306 ( .A1(n7558), .A2(n7532), .ZN(n6768) );
  NAND2_X1 U8307 ( .A1(n8083), .A2(n6769), .ZN(n6770) );
  NAND2_X1 U8308 ( .A1(n6771), .A2(n6770), .ZN(n7572) );
  INV_X1 U8309 ( .A(n7901), .ZN(n7719) );
  AND2_X1 U8310 ( .A1(n8015), .A2(n7836), .ZN(n6772) );
  NAND2_X1 U8311 ( .A1(n7939), .A2(n8080), .ZN(n6773) );
  INV_X1 U8312 ( .A(n7939), .ZN(n7708) );
  INV_X1 U8313 ( .A(n8453), .ZN(n8421) );
  OR2_X1 U8314 ( .A1(n9632), .A2(n8421), .ZN(n8419) );
  INV_X1 U8315 ( .A(n8430), .ZN(n9623) );
  NAND2_X1 U8316 ( .A1(n8430), .A2(n6777), .ZN(n6778) );
  INV_X1 U8317 ( .A(n8511), .ZN(n6780) );
  INV_X1 U8318 ( .A(n8034), .ZN(n8868) );
  NOR2_X1 U8319 ( .A1(n8864), .A2(n8383), .ZN(n6783) );
  INV_X1 U8320 ( .A(n8499), .ZN(n8363) );
  INV_X1 U8321 ( .A(n8012), .ZN(n8550) );
  NOR2_X1 U8322 ( .A1(n8325), .A2(n8077), .ZN(n6785) );
  NAND2_X1 U8323 ( .A1(n8325), .A2(n8077), .ZN(n6784) );
  NOR2_X1 U8324 ( .A1(n8542), .A2(n8322), .ZN(n6787) );
  NAND2_X1 U8325 ( .A1(n8542), .A2(n8322), .ZN(n6786) );
  NAND2_X1 U8326 ( .A1(n8301), .A2(n6788), .ZN(n6790) );
  INV_X1 U8327 ( .A(n8304), .ZN(n8538) );
  NAND2_X1 U8328 ( .A1(n8538), .A2(n8313), .ZN(n6789) );
  NOR2_X1 U8329 ( .A1(n8299), .A2(n8075), .ZN(n6791) );
  NOR2_X1 U8330 ( .A1(n8530), .A2(n8267), .ZN(n6792) );
  XNOR2_X1 U8331 ( .A(n6794), .B(n6751), .ZN(n6798) );
  NAND2_X1 U8332 ( .A1(n6833), .A2(n6830), .ZN(n6796) );
  NAND2_X1 U8333 ( .A1(n7165), .A2(n6831), .ZN(n6795) );
  NAND2_X1 U8334 ( .A1(n6798), .A2(n6797), .ZN(n6799) );
  AND2_X1 U8335 ( .A1(n7431), .A2(n6830), .ZN(n7166) );
  NAND2_X1 U8336 ( .A1(n7542), .A2(n7166), .ZN(n10202) );
  XNOR2_X1 U8337 ( .A(n6801), .B(P2_B_REG_SCAN_IN), .ZN(n6803) );
  NAND2_X1 U8338 ( .A1(n6803), .A2(n6802), .ZN(n6805) );
  OR2_X1 U8339 ( .A1(n6807), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6806) );
  NAND2_X1 U8340 ( .A1(n6802), .A2(n6808), .ZN(n6888) );
  NAND2_X1 U8341 ( .A1(n6806), .A2(n6888), .ZN(n6827) );
  NAND2_X1 U8342 ( .A1(n7031), .A2(n7030), .ZN(n6828) );
  NAND3_X1 U8343 ( .A1(n6833), .A2(n6831), .A3(n8247), .ZN(n6809) );
  NAND2_X1 U8344 ( .A1(n6839), .A2(n6809), .ZN(n6810) );
  MUX2_X1 U8345 ( .A(n6827), .B(n6828), .S(n6810), .Z(n7157) );
  NOR4_X1 U8346 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_31__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6819) );
  INV_X1 U8347 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n8760) );
  INV_X1 U8348 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n8835) );
  INV_X1 U8349 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n8764) );
  INV_X1 U8350 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n8731) );
  NAND4_X1 U8351 ( .A1(n8760), .A2(n8835), .A3(n8764), .A4(n8731), .ZN(n6816)
         );
  NOR4_X1 U8352 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6814) );
  NOR4_X1 U8353 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6813) );
  NOR4_X1 U8354 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6812) );
  NOR4_X1 U8355 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n6811) );
  NAND4_X1 U8356 ( .A1(n6814), .A2(n6813), .A3(n6812), .A4(n6811), .ZN(n6815)
         );
  NOR4_X1 U8357 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        n6816), .A4(n6815), .ZN(n6818) );
  NOR4_X1 U8358 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n6817) );
  AND3_X1 U8359 ( .A1(n6819), .A2(n6818), .A3(n6817), .ZN(n6820) );
  OR2_X1 U8360 ( .A1(n6807), .A2(n6820), .ZN(n6829) );
  OR2_X1 U8361 ( .A1(n6839), .A2(n6821), .ZN(n7003) );
  AND3_X1 U8362 ( .A1(n6829), .A2(n7164), .A3(n7003), .ZN(n7158) );
  NAND2_X1 U8363 ( .A1(n6828), .A2(n6827), .ZN(n6837) );
  OR2_X1 U8364 ( .A1(n10202), .A2(n7165), .ZN(n7162) );
  AND3_X1 U8365 ( .A1(n7158), .A2(n6837), .A3(n7162), .ZN(n6822) );
  AND2_X2 U8366 ( .A1(n7157), .A2(n6822), .ZN(n10264) );
  INV_X1 U8367 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6823) );
  NAND2_X1 U8368 ( .A1(n10264), .A2(n10180), .ZN(n8519) );
  NAND2_X1 U8369 ( .A1(n6826), .A2(n5041), .ZN(P2_U3488) );
  OR2_X1 U8370 ( .A1(n6828), .A2(n6827), .ZN(n7159) );
  INV_X1 U8371 ( .A(n6829), .ZN(n6836) );
  NOR2_X1 U8372 ( .A1(n7159), .A2(n6836), .ZN(n7009) );
  NAND2_X1 U8373 ( .A1(n7009), .A2(n7164), .ZN(n6995) );
  NAND2_X1 U8374 ( .A1(n6831), .A2(n6830), .ZN(n6832) );
  NOR2_X1 U8375 ( .A1(n6832), .A2(n7165), .ZN(n6834) );
  NAND2_X1 U8376 ( .A1(n6834), .A2(n6833), .ZN(n6996) );
  AND2_X1 U8377 ( .A1(n7183), .A2(n6996), .ZN(n6835) );
  NOR2_X1 U8378 ( .A1(n7012), .A2(n6838), .ZN(n6997) );
  NAND3_X1 U8379 ( .A1(n6996), .A2(n6839), .A3(n10225), .ZN(n6994) );
  OR2_X1 U8380 ( .A1(n10225), .A2(n7166), .ZN(n10153) );
  NAND2_X1 U8381 ( .A1(n6994), .A2(n10153), .ZN(n7002) );
  NAND2_X1 U8382 ( .A1(n6997), .A2(n7002), .ZN(n6840) );
  INV_X1 U8383 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6842) );
  NAND2_X1 U8384 ( .A1(n6844), .A2(n6843), .ZN(n6845) );
  NAND2_X1 U8385 ( .A1(n10240), .A2(n10180), .ZN(n8873) );
  NAND2_X1 U8386 ( .A1(n6845), .A2(n5037), .ZN(P2_U3456) );
  INV_X1 U8387 ( .A(n7015), .ZN(n6846) );
  OR2_X2 U8388 ( .A1(n7004), .A2(n6846), .ZN(n8224) );
  INV_X1 U8389 ( .A(n6847), .ZN(n6908) );
  NOR2_X1 U8390 ( .A1(n6848), .A2(n6908), .ZN(n9064) );
  INV_X1 U8391 ( .A(n6850), .ZN(n6849) );
  OR2_X1 U8392 ( .A1(n7004), .A2(n6849), .ZN(n7057) );
  NAND2_X1 U8393 ( .A1(n6851), .A2(n6850), .ZN(n6852) );
  NAND2_X1 U8394 ( .A1(n7057), .A2(n6852), .ZN(n7056) );
  OR2_X1 U8395 ( .A1(n7056), .A2(n6853), .ZN(n6854) );
  NAND2_X1 U8396 ( .A1(n6854), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  XNOR2_X1 U8397 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  MUX2_X1 U8398 ( .A(n6855), .B(n9071), .S(P1_STATE_REG_SCAN_IN), .Z(n6856) );
  INV_X1 U8399 ( .A(n6856), .ZN(P1_U3355) );
  OR2_X2 U8400 ( .A1(n6860), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9562) );
  NAND2_X1 U8401 ( .A1(n6857), .A2(P1_U3086), .ZN(n9565) );
  INV_X1 U8402 ( .A(n9565), .ZN(n7655) );
  INV_X1 U8403 ( .A(n7655), .ZN(n7781) );
  OAI222_X1 U8404 ( .A1(n9562), .A2(n6858), .B1(n7781), .B2(n6861), .C1(n9077), 
        .C2(P1_U3086), .ZN(P1_U3353) );
  OAI222_X1 U8405 ( .A1(n9562), .A2(n6859), .B1(n7781), .B2(n6867), .C1(n9672), 
        .C2(n4454), .ZN(P1_U3354) );
  AND2_X1 U8406 ( .A1(n6857), .A2(P2_U3151), .ZN(n8884) );
  INV_X2 U8407 ( .A(n8884), .ZN(n8888) );
  OR2_X1 U8408 ( .A1(n6860), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7757) );
  OAI222_X1 U8409 ( .A1(n8888), .A2(n6862), .B1(n4571), .B2(P2_U3151), .C1(
        n7757), .C2(n6861), .ZN(P2_U3293) );
  OAI222_X1 U8410 ( .A1(n9562), .A2(n8841), .B1(n7781), .B2(n6863), .C1(n9603), 
        .C2(P1_U3086), .ZN(P1_U3352) );
  OAI222_X1 U8411 ( .A1(n8888), .A2(n6864), .B1(n4838), .B2(P2_U3151), .C1(
        n7757), .C2(n6863), .ZN(P2_U3292) );
  OAI222_X1 U8412 ( .A1(n9562), .A2(n6865), .B1(P1_U3086), .B2(n9687), .C1(
        n6866), .C2(n7781), .ZN(P1_U3351) );
  OAI222_X1 U8413 ( .A1(n8888), .A2(n8672), .B1(n7148), .B2(P2_U3151), .C1(
        n7757), .C2(n6866), .ZN(P2_U3291) );
  INV_X1 U8414 ( .A(n7757), .ZN(n8879) );
  INV_X1 U8415 ( .A(n8879), .ZN(n8890) );
  OAI222_X1 U8416 ( .A1(n8888), .A2(n6868), .B1(n10057), .B2(P2_U3151), .C1(
        n8890), .C2(n6867), .ZN(P2_U3294) );
  OAI222_X1 U8417 ( .A1(n9562), .A2(n6869), .B1(n7781), .B2(n6870), .C1(n6928), 
        .C2(n4454), .ZN(P1_U3350) );
  OAI222_X1 U8418 ( .A1(n8888), .A2(n6871), .B1(n10078), .B2(P2_U3151), .C1(
        n7757), .C2(n6870), .ZN(P2_U3290) );
  OAI222_X1 U8419 ( .A1(n7757), .A2(n6873), .B1(n7626), .B2(P2_U3151), .C1(
        n6872), .C2(n8888), .ZN(P2_U3289) );
  OAI222_X1 U8420 ( .A1(n9562), .A2(n6874), .B1(n9565), .B2(n6873), .C1(n6944), 
        .C2(P1_U3086), .ZN(P1_U3349) );
  OAI222_X1 U8421 ( .A1(n7757), .A2(n6875), .B1(n10111), .B2(P2_U3151), .C1(
        n8780), .C2(n8888), .ZN(P2_U3288) );
  INV_X1 U8422 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6876) );
  INV_X1 U8423 ( .A(n6947), .ZN(n9589) );
  OAI222_X1 U8424 ( .A1(n9562), .A2(n6876), .B1(n9565), .B2(n6875), .C1(n9589), 
        .C2(n4454), .ZN(P1_U3348) );
  INV_X1 U8425 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6878) );
  INV_X1 U8426 ( .A(n6877), .ZN(n6879) );
  OAI222_X1 U8427 ( .A1(n8888), .A2(n6878), .B1(n8890), .B2(n6879), .C1(
        P2_U3151), .C2(n7629), .ZN(P2_U3287) );
  INV_X1 U8428 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6880) );
  INV_X1 U8429 ( .A(n6950), .ZN(n9618) );
  OAI222_X1 U8430 ( .A1(n9562), .A2(n6880), .B1(n7781), .B2(n6879), .C1(n4454), 
        .C2(n9618), .ZN(P1_U3347) );
  INV_X1 U8431 ( .A(n9562), .ZN(n9553) );
  AOI22_X1 U8432 ( .A1(n9575), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9553), .ZN(n6881) );
  OAI21_X1 U8433 ( .B1(n6890), .B2(n9565), .A(n6881), .ZN(P1_U3345) );
  NAND2_X1 U8434 ( .A1(n7279), .A2(n6882), .ZN(n6883) );
  AND2_X1 U8435 ( .A1(n6884), .A2(n6883), .ZN(n6926) );
  INV_X1 U8436 ( .A(n6926), .ZN(n6886) );
  NAND2_X1 U8437 ( .A1(n6885), .A2(n7657), .ZN(n6925) );
  AND2_X1 U8438 ( .A1(n6886), .A2(n6925), .ZN(n9803) );
  NOR2_X1 U8439 ( .A1(n9803), .A2(P1_U3973), .ZN(P1_U3085) );
  NAND2_X1 U8440 ( .A1(n7164), .A2(n6807), .ZN(n6895) );
  INV_X1 U8441 ( .A(n7030), .ZN(n6887) );
  AOI22_X1 U8442 ( .A1(n6895), .A2(n4634), .B1(n7015), .B2(n6887), .ZN(
        P2_U3376) );
  INV_X1 U8443 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n8763) );
  INV_X1 U8444 ( .A(n6888), .ZN(n6889) );
  AOI22_X1 U8445 ( .A1(n6895), .A2(n8763), .B1(n7015), .B2(n6889), .ZN(
        P2_U3377) );
  INV_X1 U8446 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n8759) );
  OAI222_X1 U8447 ( .A1(n8890), .A2(n6890), .B1(n7763), .B2(P2_U3151), .C1(
        n8759), .C2(n8888), .ZN(P2_U3285) );
  INV_X1 U8448 ( .A(n6891), .ZN(n6894) );
  INV_X1 U8449 ( .A(n7666), .ZN(n7618) );
  OAI222_X1 U8450 ( .A1(n7757), .A2(n6894), .B1(n7618), .B2(P2_U3151), .C1(
        n6897), .C2(n8888), .ZN(P2_U3286) );
  AND2_X1 U8451 ( .A1(n6895), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8452 ( .A1(n6895), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8453 ( .A1(n6895), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8454 ( .A1(n6895), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8455 ( .A1(n6895), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8456 ( .A1(n6895), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8457 ( .A1(n6895), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8458 ( .A1(n6895), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8459 ( .A1(n6895), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8460 ( .A1(n6895), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8461 ( .A1(n6895), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8462 ( .A1(n6895), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8463 ( .A1(n6895), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8464 ( .A1(n6895), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8465 ( .A1(n6895), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8466 ( .A1(n6895), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8467 ( .A1(n6895), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8468 ( .A1(n6895), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8469 ( .A1(n6895), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8470 ( .A1(n6895), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8471 ( .A1(n6895), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8472 ( .A1(n6895), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8473 ( .A1(n6895), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  INV_X1 U8474 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6893) );
  NAND2_X1 U8475 ( .A1(n7274), .A2(n9064), .ZN(n6892) );
  OAI21_X1 U8476 ( .B1(P1_U3973), .B2(n6893), .A(n6892), .ZN(P1_U3554) );
  INV_X1 U8477 ( .A(n9122), .ZN(n6957) );
  OAI222_X1 U8478 ( .A1(n9562), .A2(n8687), .B1(n7781), .B2(n6894), .C1(n6957), 
        .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U8479 ( .A(n6895), .ZN(n6896) );
  INV_X1 U8480 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n8828) );
  NOR2_X1 U8481 ( .A1(n6896), .A2(n8828), .ZN(P2_U3254) );
  INV_X1 U8482 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n8827) );
  NOR2_X1 U8483 ( .A1(n6896), .A2(n8827), .ZN(P2_U3258) );
  INV_X1 U8484 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n8714) );
  NOR2_X1 U8485 ( .A1(n6896), .A2(n8714), .ZN(P2_U3253) );
  NOR2_X1 U8486 ( .A1(n6896), .A2(n8835), .ZN(P2_U3259) );
  NOR2_X1 U8487 ( .A1(n6896), .A2(n8760), .ZN(P2_U3244) );
  NOR2_X1 U8488 ( .A1(n6896), .A2(n8764), .ZN(P2_U3237) );
  NOR2_X1 U8489 ( .A1(n6896), .A2(n8731), .ZN(P2_U3241) );
  MUX2_X1 U8490 ( .A(n6897), .B(n8926), .S(n9064), .Z(n6898) );
  INV_X1 U8491 ( .A(n6898), .ZN(P1_U3563) );
  AOI22_X1 U8492 ( .A1(n9737), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9553), .ZN(n6899) );
  OAI21_X1 U8493 ( .B1(n6905), .B2(n9565), .A(n6899), .ZN(P1_U3343) );
  INV_X1 U8494 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6901) );
  INV_X1 U8495 ( .A(n6900), .ZN(n6902) );
  INV_X1 U8496 ( .A(n7792), .ZN(n7759) );
  OAI222_X1 U8497 ( .A1(n8888), .A2(n6901), .B1(n8890), .B2(n6902), .C1(
        P2_U3151), .C2(n7759), .ZN(P2_U3284) );
  INV_X1 U8498 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6903) );
  INV_X1 U8499 ( .A(n9124), .ZN(n9732) );
  OAI222_X1 U8500 ( .A1(n9562), .A2(n6903), .B1(n7781), .B2(n6902), .C1(
        P1_U3086), .C2(n9732), .ZN(P1_U3344) );
  INV_X1 U8501 ( .A(n8106), .ZN(n7803) );
  INV_X1 U8502 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6904) );
  OAI222_X1 U8503 ( .A1(n7757), .A2(n6905), .B1(n7803), .B2(P2_U3151), .C1(
        n6904), .C2(n8888), .ZN(P2_U3283) );
  XNOR2_X1 U8504 ( .A(n6907), .B(n6906), .ZN(n9067) );
  NOR2_X1 U8505 ( .A1(n6909), .A2(n6908), .ZN(n7022) );
  INV_X1 U8506 ( .A(n7022), .ZN(n6910) );
  AOI22_X1 U8507 ( .A1(n6910), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n5133), .B2(
        n4451), .ZN(n6912) );
  INV_X1 U8508 ( .A(n9053), .ZN(n9021) );
  NAND2_X1 U8509 ( .A1(n9021), .A2(n9065), .ZN(n6911) );
  OAI211_X1 U8510 ( .C1(n9067), .C2(n9056), .A(n6912), .B(n6911), .ZN(P1_U3232) );
  NOR2_X1 U8511 ( .A1(n9122), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6913) );
  AOI21_X1 U8512 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n9122), .A(n6913), .ZN(
        n6924) );
  INV_X1 U8513 ( .A(n6944), .ZN(n9718) );
  INV_X1 U8514 ( .A(n6928), .ZN(n9695) );
  XNOR2_X1 U8515 ( .A(n6928), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n9694) );
  XNOR2_X1 U8516 ( .A(n9077), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n9079) );
  NAND2_X1 U8517 ( .A1(n6929), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6915) );
  INV_X1 U8518 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n8753) );
  INV_X1 U8519 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7240) );
  NOR2_X1 U8520 ( .A1(n9071), .A2(n7240), .ZN(n9068) );
  INV_X1 U8521 ( .A(n9068), .ZN(n9663) );
  NOR2_X1 U8522 ( .A1(n9664), .A2(n9663), .ZN(n9662) );
  INV_X1 U8523 ( .A(n9662), .ZN(n6914) );
  NAND2_X1 U8524 ( .A1(n6915), .A2(n6914), .ZN(n9080) );
  NAND2_X1 U8525 ( .A1(n9079), .A2(n9080), .ZN(n9084) );
  INV_X1 U8526 ( .A(n9077), .ZN(n6933) );
  NAND2_X1 U8527 ( .A1(n6933), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6916) );
  NAND2_X1 U8528 ( .A1(n9084), .A2(n6916), .ZN(n9596) );
  OR2_X1 U8529 ( .A1(n6935), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6918) );
  NAND2_X1 U8530 ( .A1(n6935), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6917) );
  AND2_X1 U8531 ( .A1(n6918), .A2(n6917), .ZN(n9597) );
  AOI21_X1 U8532 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n6935), .A(n9594), .ZN(
        n9678) );
  INV_X1 U8533 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6919) );
  AOI22_X1 U8534 ( .A1(n6938), .A2(n6919), .B1(P1_REG2_REG_4__SCAN_IN), .B2(
        n9687), .ZN(n9679) );
  NOR2_X1 U8535 ( .A1(n9678), .A2(n9679), .ZN(n9677) );
  AOI21_X1 U8536 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n6938), .A(n9677), .ZN(
        n6920) );
  INV_X1 U8537 ( .A(n6920), .ZN(n9693) );
  NAND2_X1 U8538 ( .A1(n9694), .A2(n9693), .ZN(n9692) );
  NAND2_X1 U8539 ( .A1(n9718), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6921) );
  OAI21_X1 U8540 ( .B1(n9718), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6921), .ZN(
        n9714) );
  INV_X1 U8541 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6922) );
  AOI22_X1 U8542 ( .A1(n6947), .A2(n6922), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n9589), .ZN(n9581) );
  NOR2_X1 U8543 ( .A1(n9580), .A2(n9581), .ZN(n9579) );
  INV_X1 U8544 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n8788) );
  AOI22_X1 U8545 ( .A1(n6950), .A2(n8788), .B1(P1_REG2_REG_8__SCAN_IN), .B2(
        n9618), .ZN(n9610) );
  OAI21_X1 U8546 ( .B1(n6924), .B2(n6923), .A(n9121), .ZN(n6959) );
  NAND2_X1 U8547 ( .A1(n6926), .A2(n6925), .ZN(n9660) );
  INV_X1 U8548 ( .A(n9069), .ZN(n6927) );
  OR2_X1 U8549 ( .A1(n9660), .A2(n6927), .ZN(n9797) );
  OR2_X1 U8550 ( .A1(n9660), .A2(n9066), .ZN(n9835) );
  INV_X1 U8551 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10026) );
  AOI22_X1 U8552 ( .A1(n9122), .A2(P1_REG1_REG_9__SCAN_IN), .B1(n10026), .B2(
        n6957), .ZN(n6952) );
  XNOR2_X1 U8553 ( .A(n6928), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n9696) );
  NAND2_X1 U8554 ( .A1(n6938), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6941) );
  XNOR2_X1 U8555 ( .A(n9077), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9085) );
  NAND2_X1 U8556 ( .A1(n6929), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6932) );
  OR2_X1 U8557 ( .A1(n6929), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6930) );
  NAND2_X1 U8558 ( .A1(n6930), .A2(n6932), .ZN(n9668) );
  NOR3_X1 U8559 ( .A1(n9071), .A2(n9657), .A3(n9668), .ZN(n9666) );
  INV_X1 U8560 ( .A(n9666), .ZN(n6931) );
  NAND2_X1 U8561 ( .A1(n6932), .A2(n6931), .ZN(n9086) );
  NAND2_X1 U8562 ( .A1(n9085), .A2(n9086), .ZN(n9090) );
  NAND2_X1 U8563 ( .A1(n6933), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6934) );
  NAND2_X1 U8564 ( .A1(n9090), .A2(n6934), .ZN(n9599) );
  OR2_X1 U8565 ( .A1(n6935), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6936) );
  NAND2_X1 U8566 ( .A1(n6935), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6937) );
  AND2_X1 U8567 ( .A1(n6936), .A2(n6937), .ZN(n9600) );
  NAND2_X1 U8568 ( .A1(n9599), .A2(n9600), .ZN(n9598) );
  AND2_X1 U8569 ( .A1(n9598), .A2(n6937), .ZN(n9683) );
  INV_X1 U8570 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6939) );
  MUX2_X1 U8571 ( .A(n6939), .B(P1_REG1_REG_4__SCAN_IN), .S(n6938), .Z(n9682)
         );
  NOR2_X1 U8572 ( .A1(n9683), .A2(n9682), .ZN(n9681) );
  INV_X1 U8573 ( .A(n9681), .ZN(n6940) );
  NAND2_X1 U8574 ( .A1(n6941), .A2(n6940), .ZN(n9697) );
  NAND2_X1 U8575 ( .A1(n9696), .A2(n9697), .ZN(n9701) );
  NAND2_X1 U8576 ( .A1(n9695), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6942) );
  NAND2_X1 U8577 ( .A1(n9701), .A2(n6942), .ZN(n9708) );
  INV_X1 U8578 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6943) );
  NOR2_X1 U8579 ( .A1(n6944), .A2(n6943), .ZN(n6945) );
  AOI21_X1 U8580 ( .B1(n6944), .B2(n6943), .A(n6945), .ZN(n9709) );
  NOR2_X1 U8581 ( .A1(n9710), .A2(n6945), .ZN(n9585) );
  INV_X1 U8582 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6946) );
  MUX2_X1 U8583 ( .A(n6946), .B(P1_REG1_REG_7__SCAN_IN), .S(n6947), .Z(n9584)
         );
  NOR2_X1 U8584 ( .A1(n9585), .A2(n9584), .ZN(n9583) );
  AOI21_X1 U8585 ( .B1(n6947), .B2(P1_REG1_REG_7__SCAN_IN), .A(n9583), .ZN(
        n9613) );
  OR2_X1 U8586 ( .A1(n6950), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6949) );
  NAND2_X1 U8587 ( .A1(n6950), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6948) );
  NAND2_X1 U8588 ( .A1(n6949), .A2(n6948), .ZN(n9614) );
  NOR2_X1 U8589 ( .A1(n9613), .A2(n9614), .ZN(n9612) );
  AOI21_X1 U8590 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n6950), .A(n9612), .ZN(
        n6951) );
  NAND2_X1 U8591 ( .A1(n6952), .A2(n6951), .ZN(n9099) );
  OAI21_X1 U8592 ( .B1(n6952), .B2(n6951), .A(n9099), .ZN(n6954) );
  OR2_X1 U8593 ( .A1(n9660), .A2(n6953), .ZN(n9784) );
  NAND2_X1 U8594 ( .A1(n6954), .A2(n9829), .ZN(n6956) );
  NOR2_X1 U8595 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8730), .ZN(n7651) );
  AOI21_X1 U8596 ( .B1(n9803), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7651), .ZN(
        n6955) );
  OAI211_X1 U8597 ( .C1(n9835), .C2(n6957), .A(n6956), .B(n6955), .ZN(n6958)
         );
  AOI21_X1 U8598 ( .B1(n6959), .B2(n9825), .A(n6958), .ZN(n6960) );
  INV_X1 U8599 ( .A(n6960), .ZN(P1_U3252) );
  AOI22_X1 U8600 ( .A1(n9753), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9553), .ZN(n6961) );
  OAI21_X1 U8601 ( .B1(n6984), .B2(n9565), .A(n6961), .ZN(P1_U3342) );
  NAND2_X1 U8602 ( .A1(n6963), .A2(n6962), .ZN(n6967) );
  AND2_X1 U8603 ( .A1(n6964), .A2(n9546), .ZN(n6966) );
  NAND2_X1 U8604 ( .A1(n6966), .A2(n6965), .ZN(n7226) );
  NOR2_X1 U8605 ( .A1(n6967), .A2(n7226), .ZN(n6980) );
  INV_X1 U8606 ( .A(n6979), .ZN(n7229) );
  AND2_X2 U8607 ( .A1(n6980), .A2(n7229), .ZN(n10013) );
  INV_X1 U8608 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n8637) );
  NAND2_X1 U8609 ( .A1(n6969), .A2(n6968), .ZN(n6970) );
  NAND2_X1 U8610 ( .A1(n6970), .A2(n6977), .ZN(n6971) );
  OR2_X1 U8611 ( .A1(n6971), .A2(n7231), .ZN(n9887) );
  NAND2_X1 U8612 ( .A1(n6972), .A2(n7433), .ZN(n9991) );
  NAND2_X1 U8613 ( .A1(n9887), .A2(n9991), .ZN(n10009) );
  OR2_X1 U8614 ( .A1(n7544), .A2(n9294), .ZN(n6973) );
  AND2_X1 U8615 ( .A1(n6974), .A2(n6973), .ZN(n9420) );
  INV_X1 U8616 ( .A(n7232), .ZN(n6975) );
  OAI21_X1 U8617 ( .B1(n10009), .B2(n9890), .A(n6975), .ZN(n6976) );
  NAND2_X1 U8618 ( .A1(n7279), .A2(n5882), .ZN(n9881) );
  NAND2_X1 U8619 ( .A1(n9065), .A2(n9864), .ZN(n7233) );
  OAI211_X1 U8620 ( .C1(n6977), .C2(n9901), .A(n6976), .B(n7233), .ZN(n6981)
         );
  NAND2_X1 U8621 ( .A1(n6981), .A2(n10013), .ZN(n6978) );
  OAI21_X1 U8622 ( .B1(n10013), .B2(n8637), .A(n6978), .ZN(P1_U3453) );
  AND2_X2 U8623 ( .A1(n6980), .A2(n6979), .ZN(n10033) );
  NAND2_X1 U8624 ( .A1(n6981), .A2(n10033), .ZN(n6982) );
  OAI21_X1 U8625 ( .B1(n10033), .B2(n9657), .A(n6982), .ZN(P1_U3522) );
  INV_X1 U8626 ( .A(n8099), .ZN(n8125) );
  INV_X1 U8627 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6983) );
  OAI222_X1 U8628 ( .A1(n7757), .A2(n6984), .B1(n8125), .B2(P2_U3151), .C1(
        n6983), .C2(n8888), .ZN(P2_U3282) );
  NAND2_X1 U8629 ( .A1(n8224), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6985) );
  OAI21_X1 U8630 ( .B1(n8344), .B2(n8224), .A(n6985), .ZN(P2_U3513) );
  OAI21_X1 U8631 ( .B1(n6988), .B2(n6987), .A(n6986), .ZN(n6991) );
  INV_X1 U8632 ( .A(n4451), .ZN(n9046) );
  INV_X1 U8633 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9892) );
  OAI22_X1 U8634 ( .A1(n9046), .A2(n9920), .B1(n7022), .B2(n9892), .ZN(n6990)
         );
  INV_X1 U8635 ( .A(n7274), .ZN(n9884) );
  INV_X1 U8636 ( .A(n9934), .ZN(n9882) );
  OAI22_X1 U8637 ( .A1(n9884), .A2(n9041), .B1(n9053), .B2(n9882), .ZN(n6989)
         );
  AOI211_X1 U8638 ( .C1(n6991), .C2(n9038), .A(n6990), .B(n6989), .ZN(n6992)
         );
  INV_X1 U8639 ( .A(n6992), .ZN(P1_U3222) );
  NAND2_X1 U8640 ( .A1(n7164), .A2(n7166), .ZN(n6993) );
  NAND2_X1 U8641 ( .A1(n6995), .A2(n6993), .ZN(n8042) );
  INV_X1 U8642 ( .A(n8033), .ZN(n8070) );
  INV_X1 U8643 ( .A(n7186), .ZN(n7027) );
  OR2_X1 U8644 ( .A1(n6995), .A2(n6994), .ZN(n6999) );
  INV_X1 U8645 ( .A(n6996), .ZN(n7005) );
  NAND2_X1 U8646 ( .A1(n6997), .A2(n7005), .ZN(n6998) );
  INV_X1 U8647 ( .A(n7183), .ZN(n7000) );
  NAND2_X1 U8648 ( .A1(n7164), .A2(n7000), .ZN(n7010) );
  NOR2_X1 U8649 ( .A1(n7012), .A2(n7010), .ZN(n7043) );
  AOI22_X1 U8650 ( .A1(n7027), .A2(n8058), .B1(n8043), .B2(n8089), .ZN(n7017)
         );
  INV_X1 U8651 ( .A(n7002), .ZN(n7008) );
  AND2_X1 U8652 ( .A1(n7004), .A2(n7003), .ZN(n7007) );
  NAND2_X1 U8653 ( .A1(n7012), .A2(n7005), .ZN(n7006) );
  OAI211_X1 U8654 ( .C1(n7009), .C2(n7008), .A(n7007), .B(n7006), .ZN(n7014)
         );
  INV_X1 U8655 ( .A(n7010), .ZN(n7011) );
  AND2_X1 U8656 ( .A1(n7012), .A2(n7011), .ZN(n7013) );
  AOI21_X1 U8657 ( .B1(n7014), .B2(P2_STATE_REG_SCAN_IN), .A(n7013), .ZN(n7117) );
  NAND2_X1 U8658 ( .A1(n7117), .A2(n7015), .ZN(n7097) );
  NAND2_X1 U8659 ( .A1(n7097), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7016) );
  OAI211_X1 U8660 ( .C1(n8070), .C2(n7189), .A(n7017), .B(n7016), .ZN(P2_U3172) );
  INV_X1 U8661 ( .A(n8154), .ZN(n8138) );
  INV_X1 U8662 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7018) );
  OAI222_X1 U8663 ( .A1(n7757), .A2(n7019), .B1(n8138), .B2(P2_U3151), .C1(
        n7018), .C2(n8888), .ZN(P2_U3281) );
  INV_X1 U8664 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n8678) );
  INV_X1 U8665 ( .A(n9126), .ZN(n9779) );
  OAI222_X1 U8666 ( .A1(n9562), .A2(n8678), .B1(n7781), .B2(n7019), .C1(n9779), 
        .C2(n4454), .ZN(P1_U3341) );
  XOR2_X1 U8667 ( .A(n7020), .B(n7021), .Z(n7026) );
  INV_X1 U8668 ( .A(n9041), .ZN(n9051) );
  INV_X1 U8669 ( .A(n9063), .ZN(n7294) );
  NOR2_X1 U8670 ( .A1(n9053), .A2(n7294), .ZN(n7024) );
  INV_X1 U8671 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n8684) );
  OAI22_X1 U8672 ( .A1(n9046), .A2(n9930), .B1(n7022), .B2(n8684), .ZN(n7023)
         );
  AOI211_X1 U8673 ( .C1(n9051), .C2(n9065), .A(n7024), .B(n7023), .ZN(n7025)
         );
  OAI21_X1 U8674 ( .B1(n7026), .B2(n9056), .A(n7025), .ZN(P1_U3237) );
  INV_X1 U8675 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n8685) );
  OAI21_X1 U8676 ( .B1(n6797), .B2(n10234), .A(n7027), .ZN(n7028) );
  OR2_X1 U8677 ( .A1(n6757), .A2(n10158), .ZN(n7184) );
  OAI211_X1 U8678 ( .C1(n10225), .C2(n7189), .A(n7028), .B(n7184), .ZN(n7085)
         );
  NAND2_X1 U8679 ( .A1(n7085), .A2(n10264), .ZN(n7029) );
  OAI21_X1 U8680 ( .B1(n10264), .B2(n8685), .A(n7029), .ZN(P2_U3459) );
  XNOR2_X1 U8681 ( .A(n7033), .B(n7090), .ZN(n7034) );
  NAND2_X1 U8682 ( .A1(n6757), .A2(n7034), .ZN(n7093) );
  INV_X1 U8683 ( .A(n7034), .ZN(n7035) );
  NAND2_X1 U8684 ( .A1(n7035), .A2(n8089), .ZN(n7036) );
  OAI21_X1 U8685 ( .B1(n7037), .B2(n7091), .A(n7154), .ZN(n7041) );
  NAND2_X1 U8686 ( .A1(n7189), .A2(n7091), .ZN(n7039) );
  INV_X1 U8687 ( .A(n7094), .ZN(n7040) );
  AOI21_X1 U8688 ( .B1(n7038), .B2(n7041), .A(n7040), .ZN(n7048) );
  INV_X1 U8689 ( .A(n8043), .ZN(n8064) );
  NAND2_X1 U8690 ( .A1(n7043), .A2(n7042), .ZN(n8031) );
  NOR2_X1 U8691 ( .A1(n7044), .A2(n10225), .ZN(n10172) );
  AOI22_X1 U8692 ( .A1(n8062), .A2(n6010), .B1(n10172), .B2(n8042), .ZN(n7045)
         );
  OAI21_X1 U8693 ( .B1(n7121), .B2(n8064), .A(n7045), .ZN(n7046) );
  AOI21_X1 U8694 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7097), .A(n7046), .ZN(
        n7047) );
  OAI21_X1 U8695 ( .B1(n7048), .B2(n8050), .A(n7047), .ZN(P2_U3162) );
  INV_X1 U8696 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n8744) );
  AND2_X1 U8697 ( .A1(n10039), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7049) );
  OAI21_X1 U8698 ( .B1(n10057), .B2(n7049), .A(n7050), .ZN(n10048) );
  INV_X1 U8699 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10047) );
  INV_X1 U8700 ( .A(n7050), .ZN(n7051) );
  NOR2_X1 U8701 ( .A1(n10051), .A2(n7051), .ZN(n10067) );
  XNOR2_X1 U8702 ( .A(n10074), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n10068) );
  AOI21_X1 U8703 ( .B1(n8744), .B2(n7052), .A(n7130), .ZN(n7083) );
  INV_X1 U8704 ( .A(n7054), .ZN(n7068) );
  NAND2_X1 U8705 ( .A1(n7068), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8880) );
  OR2_X1 U8706 ( .A1(n7056), .A2(n8880), .ZN(n7076) );
  INV_X1 U8707 ( .A(n7076), .ZN(n10036) );
  NAND2_X1 U8708 ( .A1(n10036), .A2(n6755), .ZN(n10135) );
  INV_X1 U8709 ( .A(n7057), .ZN(n7053) );
  NOR2_X2 U8710 ( .A1(P2_U3150), .A2(n7053), .ZN(n10115) );
  NAND2_X1 U8711 ( .A1(n10115), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n7082) );
  AND2_X1 U8712 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7118) );
  NOR2_X1 U8713 ( .A1(n8241), .A2(P2_U3151), .ZN(n8883) );
  NAND2_X1 U8714 ( .A1(n8883), .A2(n7054), .ZN(n7055) );
  OR2_X1 U8715 ( .A1(n7056), .A2(n7055), .ZN(n7059) );
  OR2_X1 U8716 ( .A1(n8880), .A2(n7057), .ZN(n7058) );
  NAND2_X1 U8717 ( .A1(n7059), .A2(n7058), .ZN(n10139) );
  MUX2_X1 U8718 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8241), .Z(n7133) );
  XNOR2_X1 U8719 ( .A(n7133), .B(n4838), .ZN(n7067) );
  INV_X1 U8720 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10241) );
  MUX2_X1 U8721 ( .A(n10047), .B(n10241), .S(n6509), .Z(n7061) );
  XNOR2_X1 U8722 ( .A(n7061), .B(n10057), .ZN(n10040) );
  INV_X1 U8723 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7060) );
  MUX2_X1 U8724 ( .A(n7060), .B(n8685), .S(n6509), .Z(n10034) );
  INV_X1 U8725 ( .A(n7061), .ZN(n7062) );
  AOI22_X1 U8726 ( .A1(n10040), .A2(n10041), .B1(n10057), .B2(n7062), .ZN(
        n10058) );
  MUX2_X1 U8727 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n6509), .Z(n7063) );
  XNOR2_X1 U8728 ( .A(n7063), .B(n4571), .ZN(n10059) );
  INV_X1 U8729 ( .A(n4571), .ZN(n7065) );
  INV_X1 U8730 ( .A(n7063), .ZN(n7064) );
  OAI22_X1 U8731 ( .A1(n10058), .A2(n10059), .B1(n7065), .B2(n7064), .ZN(n7066) );
  AOI21_X1 U8732 ( .B1(n7067), .B2(n7066), .A(n7134), .ZN(n7069) );
  OR2_X1 U8733 ( .A1(n8224), .A2(n7068), .ZN(n8250) );
  OR2_X1 U8734 ( .A1(n7069), .A2(n8250), .ZN(n7079) );
  INV_X1 U8735 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10245) );
  AND2_X1 U8736 ( .A1(n10039), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7070) );
  INV_X1 U8737 ( .A(n7071), .ZN(n7072) );
  OAI21_X1 U8738 ( .B1(n4571), .B2(P2_REG1_REG_2__SCAN_IN), .A(n7074), .ZN(
        n10064) );
  INV_X1 U8739 ( .A(n10064), .ZN(n7073) );
  AND2_X2 U8740 ( .A1(n10062), .A2(n7073), .ZN(n10063) );
  AOI21_X1 U8741 ( .B1(n10245), .B2(n7075), .A(n7140), .ZN(n7077) );
  NOR2_X1 U8742 ( .A1(n7076), .A2(n6755), .ZN(n10121) );
  OR2_X1 U8743 ( .A1(n7077), .A2(n10133), .ZN(n7078) );
  OAI211_X1 U8744 ( .C1(n10112), .C2(n4838), .A(n7079), .B(n7078), .ZN(n7080)
         );
  NOR2_X1 U8745 ( .A1(n7118), .A2(n7080), .ZN(n7081) );
  OAI211_X1 U8746 ( .C1(n7083), .C2(n10135), .A(n7082), .B(n7081), .ZN(
        P2_U3185) );
  INV_X1 U8747 ( .A(n8148), .ZN(n8174) );
  INV_X1 U8748 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7084) );
  OAI222_X1 U8749 ( .A1(n7757), .A2(n7088), .B1(n8174), .B2(P2_U3151), .C1(
        n7084), .C2(n8888), .ZN(P2_U3280) );
  INV_X1 U8750 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7087) );
  NAND2_X1 U8751 ( .A1(n7085), .A2(n10240), .ZN(n7086) );
  OAI21_X1 U8752 ( .B1(n7087), .B2(n10240), .A(n7086), .ZN(P2_U3390) );
  INV_X1 U8753 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7089) );
  OAI222_X1 U8754 ( .A1(n9562), .A2(n7089), .B1(n7781), .B2(n7088), .C1(n9128), 
        .C2(P1_U3086), .ZN(P1_U3340) );
  XNOR2_X1 U8755 ( .A(n7092), .B(n7091), .ZN(n7111) );
  XNOR2_X1 U8756 ( .A(n7121), .B(n7111), .ZN(n7096) );
  NAND2_X1 U8757 ( .A1(n7095), .A2(n7096), .ZN(n7114) );
  OAI21_X1 U8758 ( .B1(n7096), .B2(n7095), .A(n7114), .ZN(n7101) );
  NAND2_X1 U8759 ( .A1(n7097), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7099) );
  NOR2_X1 U8760 ( .A1(n10154), .A2(n10225), .ZN(n10176) );
  AOI22_X1 U8761 ( .A1(n8062), .A2(n8089), .B1(n10176), .B2(n8042), .ZN(n7098)
         );
  OAI211_X1 U8762 ( .C1(n10159), .C2(n8064), .A(n7099), .B(n7098), .ZN(n7100)
         );
  AOI21_X1 U8763 ( .B1(n7101), .B2(n8058), .A(n7100), .ZN(n7102) );
  INV_X1 U8764 ( .A(n7102), .ZN(P2_U3177) );
  XNOR2_X1 U8765 ( .A(n7103), .B(n7104), .ZN(n7109) );
  INV_X1 U8766 ( .A(n9863), .ZN(n7336) );
  OAI22_X1 U8767 ( .A1(n9882), .A2(n9041), .B1(n9053), .B2(n7336), .ZN(n7108)
         );
  INV_X1 U8768 ( .A(n7311), .ZN(n9935) );
  NAND2_X1 U8769 ( .A1(n4454), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9605) );
  INV_X1 U8770 ( .A(n9605), .ZN(n7105) );
  AOI21_X1 U8771 ( .B1(n4451), .B2(n9935), .A(n7105), .ZN(n7106) );
  OAI21_X1 U8772 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(n9029), .A(n7106), .ZN(
        n7107) );
  AOI211_X1 U8773 ( .C1(n7109), .C2(n9038), .A(n7108), .B(n7107), .ZN(n7110)
         );
  INV_X1 U8774 ( .A(n7110), .ZN(P1_U3218) );
  INV_X1 U8775 ( .A(n7111), .ZN(n7112) );
  NAND2_X1 U8776 ( .A1(n7121), .A2(n7112), .ZN(n7113) );
  AND2_X1 U8777 ( .A1(n7114), .A2(n7113), .ZN(n7116) );
  XNOR2_X1 U8778 ( .A(n10179), .B(n7090), .ZN(n7253) );
  XNOR2_X1 U8779 ( .A(n8088), .B(n7253), .ZN(n7115) );
  OAI211_X1 U8780 ( .C1(n7116), .C2(n7115), .A(n7256), .B(n8058), .ZN(n7124)
         );
  NAND2_X1 U8781 ( .A1(n8033), .A2(n10179), .ZN(n7120) );
  AOI21_X1 U8782 ( .B1(n8043), .B2(n8087), .A(n7118), .ZN(n7119) );
  OAI211_X1 U8783 ( .C1(n7121), .C2(n8031), .A(n7120), .B(n7119), .ZN(n7122)
         );
  AOI21_X1 U8784 ( .B1(n8067), .B2(n7179), .A(n7122), .ZN(n7123) );
  NAND2_X1 U8785 ( .A1(n7124), .A2(n7123), .ZN(P2_U3158) );
  INV_X1 U8786 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7126) );
  INV_X1 U8787 ( .A(n7125), .ZN(n7127) );
  INV_X1 U8788 ( .A(n8190), .ZN(n8196) );
  OAI222_X1 U8789 ( .A1(n8888), .A2(n7126), .B1(n8890), .B2(n7127), .C1(
        P2_U3151), .C2(n8196), .ZN(P2_U3279) );
  INV_X1 U8790 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7128) );
  INV_X1 U8791 ( .A(n9807), .ZN(n9130) );
  OAI222_X1 U8792 ( .A1(n9562), .A2(n7128), .B1(n7781), .B2(n7127), .C1(n4454), 
        .C2(n9130), .ZN(P1_U3339) );
  INV_X1 U8793 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n8717) );
  AOI22_X1 U8794 ( .A1(n7624), .A2(P2_REG2_REG_4__SCAN_IN), .B1(n8717), .B2(
        n7148), .ZN(n7132) );
  AOI21_X1 U8795 ( .B1(n4549), .B2(n7132), .A(n7594), .ZN(n7153) );
  NAND2_X1 U8796 ( .A1(n10115), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n7152) );
  NAND2_X1 U8797 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7267) );
  INV_X1 U8798 ( .A(n7267), .ZN(n7150) );
  INV_X1 U8799 ( .A(n7133), .ZN(n7135) );
  MUX2_X1 U8800 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8241), .Z(n7621) );
  XNOR2_X1 U8801 ( .A(n7621), .B(n7624), .ZN(n7136) );
  NAND2_X1 U8802 ( .A1(n7137), .A2(n7136), .ZN(n7622) );
  OAI211_X1 U8803 ( .C1(n7137), .C2(n7136), .A(n10143), .B(n7622), .ZN(n7147)
         );
  NOR2_X1 U8804 ( .A1(n7139), .A2(n7138), .ZN(n7141) );
  INV_X1 U8805 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7142) );
  OR2_X1 U8806 ( .A1(n7624), .A2(n7142), .ZN(n7608) );
  OAI21_X1 U8807 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n7148), .A(n7608), .ZN(
        n7143) );
  AOI21_X1 U8808 ( .B1(n7144), .B2(n7143), .A(n7607), .ZN(n7145) );
  OR2_X1 U8809 ( .A1(n7145), .A2(n10133), .ZN(n7146) );
  OAI211_X1 U8810 ( .C1(n10112), .C2(n7148), .A(n7147), .B(n7146), .ZN(n7149)
         );
  NOR2_X1 U8811 ( .A1(n7150), .A2(n7149), .ZN(n7151) );
  OAI211_X1 U8812 ( .C1(n7153), .C2(n10135), .A(n7152), .B(n7151), .ZN(
        P2_U3186) );
  XNOR2_X1 U8813 ( .A(n7170), .B(n7154), .ZN(n7156) );
  AOI222_X1 U8814 ( .A1(n6797), .A2(n7156), .B1(n7155), .B2(n8437), .C1(n6010), 
        .C2(n8435), .ZN(n10170) );
  INV_X1 U8815 ( .A(n7157), .ZN(n7161) );
  AND2_X1 U8816 ( .A1(n7159), .A2(n7158), .ZN(n7160) );
  NAND2_X1 U8817 ( .A1(n7161), .A2(n7160), .ZN(n7171) );
  INV_X1 U8818 ( .A(n7162), .ZN(n7163) );
  NAND2_X1 U8819 ( .A1(n7164), .A2(n7163), .ZN(n10151) );
  NAND2_X1 U8820 ( .A1(n7171), .A2(n10151), .ZN(n8457) );
  INV_X2 U8821 ( .A(n8457), .ZN(n8442) );
  AND2_X1 U8822 ( .A1(n7166), .A2(n7165), .ZN(n10166) );
  INV_X1 U8823 ( .A(n10166), .ZN(n7167) );
  NAND2_X1 U8824 ( .A1(n10163), .A2(n7167), .ZN(n7168) );
  NAND2_X1 U8825 ( .A1(n10167), .A2(n7168), .ZN(n8447) );
  XNOR2_X1 U8826 ( .A(n7170), .B(n7169), .ZN(n10173) );
  INV_X1 U8827 ( .A(n10151), .ZN(n8440) );
  AOI22_X1 U8828 ( .A1(n8429), .A2(n7033), .B1(n8440), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n7172) );
  OAI21_X1 U8829 ( .B1(n10047), .B2(n10167), .A(n7172), .ZN(n7173) );
  AOI21_X1 U8830 ( .B1(n8461), .B2(n10173), .A(n7173), .ZN(n7174) );
  OAI21_X1 U8831 ( .B1(n10170), .B2(n8442), .A(n7174), .ZN(P2_U3232) );
  XNOR2_X1 U8832 ( .A(n7175), .B(n4776), .ZN(n7176) );
  AOI222_X1 U8833 ( .A1(n6797), .A2(n7176), .B1(n8087), .B2(n8437), .C1(n7155), 
        .C2(n8435), .ZN(n10183) );
  XNOR2_X1 U8834 ( .A(n7178), .B(n7177), .ZN(n10181) );
  AOI22_X1 U8835 ( .A1(n8429), .A2(n10179), .B1(n8440), .B2(n7179), .ZN(n7180)
         );
  OAI21_X1 U8836 ( .B1(n8744), .B2(n10167), .A(n7180), .ZN(n7181) );
  AOI21_X1 U8837 ( .B1(n10181), .B2(n8461), .A(n7181), .ZN(n7182) );
  OAI21_X1 U8838 ( .B1(n10183), .B2(n8442), .A(n7182), .ZN(P2_U3230) );
  NAND2_X1 U8839 ( .A1(n7183), .A2(n10225), .ZN(n7185) );
  OAI21_X1 U8840 ( .B1(n7186), .B2(n7185), .A(n7184), .ZN(n7187) );
  MUX2_X1 U8841 ( .A(n7187), .B(P2_REG2_REG_0__SCAN_IN), .S(n8442), .Z(n7191)
         );
  INV_X1 U8842 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7188) );
  OAI22_X1 U8843 ( .A1(n8411), .A2(n7189), .B1(n7188), .B2(n10151), .ZN(n7190)
         );
  OR2_X1 U8844 ( .A1(n7191), .A2(n7190), .ZN(P2_U3233) );
  INV_X1 U8845 ( .A(n7192), .ZN(n7195) );
  AOI22_X1 U8846 ( .A1(n9819), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9553), .ZN(n7193) );
  OAI21_X1 U8847 ( .B1(n7195), .B2(n9565), .A(n7193), .ZN(P1_U3338) );
  AOI22_X1 U8848 ( .A1(n8219), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n8884), .ZN(n7194) );
  OAI21_X1 U8849 ( .B1(n7195), .B2(n8890), .A(n7194), .ZN(P2_U3278) );
  XNOR2_X1 U8850 ( .A(n7199), .B(n7196), .ZN(n7197) );
  AOI222_X1 U8851 ( .A1(n6797), .A2(n7197), .B1(n8088), .B2(n8435), .C1(n8086), 
        .C2(n8437), .ZN(n10185) );
  XNOR2_X1 U8852 ( .A(n7199), .B(n7198), .ZN(n10188) );
  AOI22_X1 U8853 ( .A1(n8429), .A2(n7257), .B1(n8440), .B2(n7271), .ZN(n7200)
         );
  OAI21_X1 U8854 ( .B1(n8717), .B2(n10167), .A(n7200), .ZN(n7201) );
  AOI21_X1 U8855 ( .B1(n10188), .B2(n8461), .A(n7201), .ZN(n7202) );
  OAI21_X1 U8856 ( .B1(n10185), .B2(n8442), .A(n7202), .ZN(P2_U3229) );
  INV_X1 U8857 ( .A(n8239), .ZN(n8235) );
  INV_X1 U8858 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n8747) );
  OAI222_X1 U8859 ( .A1(n7757), .A2(n7252), .B1(n8235), .B2(P2_U3151), .C1(
        n8747), .C2(n8888), .ZN(P2_U3277) );
  INV_X1 U8860 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10274) );
  INV_X1 U8861 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9839) );
  INV_X1 U8862 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9823) );
  INV_X1 U8863 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n7203) );
  AOI22_X1 U8864 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .B1(n9823), .B2(n7203), .ZN(n10277) );
  INV_X1 U8865 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7205) );
  INV_X1 U8866 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7204) );
  AOI22_X1 U8867 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(P2_ADDR_REG_16__SCAN_IN), 
        .B1(n7205), .B2(n7204), .ZN(n10280) );
  NOR2_X1 U8868 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7206) );
  AOI21_X1 U8869 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7206), .ZN(n10283) );
  NOR2_X1 U8870 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7207) );
  AOI21_X1 U8871 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7207), .ZN(n10286) );
  INV_X1 U8872 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7208) );
  INV_X1 U8873 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9768) );
  AOI22_X1 U8874 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), 
        .B1(n7208), .B2(n9768), .ZN(n10289) );
  NOR2_X1 U8875 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7209) );
  AOI21_X1 U8876 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7209), .ZN(n10292) );
  NOR2_X1 U8877 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7210) );
  AOI21_X1 U8878 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7210), .ZN(n10295) );
  NOR2_X1 U8879 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7211) );
  AOI21_X1 U8880 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7211), .ZN(n10298) );
  NOR2_X1 U8881 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7212) );
  AOI21_X1 U8882 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7212), .ZN(n10307) );
  NOR2_X1 U8883 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7213) );
  AOI21_X1 U8884 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7213), .ZN(n10313) );
  NOR2_X1 U8885 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7214) );
  AOI21_X1 U8886 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7214), .ZN(n10310) );
  NOR2_X1 U8887 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7215) );
  AOI21_X1 U8888 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7215), .ZN(n10301) );
  NOR2_X1 U8889 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7216) );
  AOI21_X1 U8890 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7216), .ZN(n10304) );
  AND2_X1 U8891 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7217) );
  NOR2_X1 U8892 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7217), .ZN(n10266) );
  INV_X1 U8893 ( .A(n10266), .ZN(n10267) );
  INV_X1 U8894 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10269) );
  NAND3_X1 U8895 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10268) );
  NAND2_X1 U8896 ( .A1(n10269), .A2(n10268), .ZN(n10265) );
  NAND2_X1 U8897 ( .A1(n10267), .A2(n10265), .ZN(n10316) );
  NAND2_X1 U8898 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7218) );
  OAI21_X1 U8899 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7218), .ZN(n10315) );
  NOR2_X1 U8900 ( .A1(n10316), .A2(n10315), .ZN(n10314) );
  AOI21_X1 U8901 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10314), .ZN(n10319) );
  NAND2_X1 U8902 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7219) );
  OAI21_X1 U8903 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7219), .ZN(n10318) );
  NOR2_X1 U8904 ( .A1(n10319), .A2(n10318), .ZN(n10317) );
  AOI21_X1 U8905 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10317), .ZN(n10322) );
  NOR2_X1 U8906 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7220) );
  AOI21_X1 U8907 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7220), .ZN(n10321) );
  NAND2_X1 U8908 ( .A1(n10322), .A2(n10321), .ZN(n10320) );
  OAI21_X1 U8909 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10320), .ZN(n10303) );
  NAND2_X1 U8910 ( .A1(n10304), .A2(n10303), .ZN(n10302) );
  OAI21_X1 U8911 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10302), .ZN(n10300) );
  NAND2_X1 U8912 ( .A1(n10301), .A2(n10300), .ZN(n10299) );
  OAI21_X1 U8913 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10299), .ZN(n10309) );
  NAND2_X1 U8914 ( .A1(n10310), .A2(n10309), .ZN(n10308) );
  OAI21_X1 U8915 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10308), .ZN(n10312) );
  NAND2_X1 U8916 ( .A1(n10313), .A2(n10312), .ZN(n10311) );
  OAI21_X1 U8917 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10311), .ZN(n10306) );
  NAND2_X1 U8918 ( .A1(n10307), .A2(n10306), .ZN(n10305) );
  OAI21_X1 U8919 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10305), .ZN(n10297) );
  NAND2_X1 U8920 ( .A1(n10298), .A2(n10297), .ZN(n10296) );
  OAI21_X1 U8921 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10296), .ZN(n10294) );
  NAND2_X1 U8922 ( .A1(n10295), .A2(n10294), .ZN(n10293) );
  OAI21_X1 U8923 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10293), .ZN(n10291) );
  NAND2_X1 U8924 ( .A1(n10292), .A2(n10291), .ZN(n10290) );
  OAI21_X1 U8925 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10290), .ZN(n10288) );
  NAND2_X1 U8926 ( .A1(n10289), .A2(n10288), .ZN(n10287) );
  OAI21_X1 U8927 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10287), .ZN(n10285) );
  NAND2_X1 U8928 ( .A1(n10286), .A2(n10285), .ZN(n10284) );
  OAI21_X1 U8929 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10284), .ZN(n10282) );
  NAND2_X1 U8930 ( .A1(n10283), .A2(n10282), .ZN(n10281) );
  OAI21_X1 U8931 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10281), .ZN(n10279) );
  NAND2_X1 U8932 ( .A1(n10280), .A2(n10279), .ZN(n10278) );
  OAI21_X1 U8933 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10278), .ZN(n10276) );
  NAND2_X1 U8934 ( .A1(n10277), .A2(n10276), .ZN(n10275) );
  OAI21_X1 U8935 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10275), .ZN(n7221) );
  OR2_X1 U8936 ( .A1(n9839), .A2(n7221), .ZN(n10273) );
  NAND2_X1 U8937 ( .A1(n10274), .A2(n10273), .ZN(n10270) );
  NAND2_X1 U8938 ( .A1(n9839), .A2(n7221), .ZN(n10272) );
  NAND2_X1 U8939 ( .A1(n10270), .A2(n10272), .ZN(n7225) );
  NOR2_X1 U8940 ( .A1(n7223), .A2(n7222), .ZN(n7224) );
  XNOR2_X1 U8941 ( .A(n7225), .B(n7224), .ZN(ADD_1068_U4) );
  INV_X1 U8942 ( .A(n7226), .ZN(n7227) );
  NAND3_X1 U8943 ( .A1(n7229), .A2(n7228), .A3(n7227), .ZN(n7237) );
  NOR3_X1 U8944 ( .A1(n7232), .A2(n7231), .A3(n7230), .ZN(n7235) );
  INV_X1 U8945 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n8707) );
  OAI21_X1 U8946 ( .B1(n8707), .B2(n9893), .A(n7233), .ZN(n7234) );
  OAI21_X1 U8947 ( .B1(n7235), .B2(n7234), .A(n9238), .ZN(n7239) );
  INV_X2 U8948 ( .A(n9238), .ZN(n9907) );
  OR2_X1 U8949 ( .A1(n7237), .A2(n4722), .ZN(n9380) );
  INV_X1 U8950 ( .A(n9900), .ZN(n9944) );
  NOR2_X1 U8951 ( .A1(n9380), .A2(n9944), .ZN(n9431) );
  OAI21_X1 U8952 ( .B1(n9854), .B2(n9431), .A(n5133), .ZN(n7238) );
  OAI211_X1 U8953 ( .C1(n7240), .C2(n9238), .A(n7239), .B(n7238), .ZN(P1_U3293) );
  INV_X1 U8954 ( .A(n7241), .ZN(n7242) );
  AOI211_X1 U8955 ( .C1(n7244), .C2(n7243), .A(n9056), .B(n7242), .ZN(n7250)
         );
  INV_X1 U8956 ( .A(n9062), .ZN(n7350) );
  OAI22_X1 U8957 ( .A1(n7294), .A2(n9041), .B1(n9053), .B2(n7350), .ZN(n7249)
         );
  INV_X1 U8958 ( .A(n7299), .ZN(n7247) );
  INV_X1 U8959 ( .A(n9943), .ZN(n7298) );
  INV_X1 U8960 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n7245) );
  NOR2_X1 U8961 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7245), .ZN(n9676) );
  AOI21_X1 U8962 ( .B1(n4451), .B2(n7298), .A(n9676), .ZN(n7246) );
  OAI21_X1 U8963 ( .B1(n7247), .B2(n9029), .A(n7246), .ZN(n7248) );
  OR3_X1 U8964 ( .A1(n7250), .A2(n7249), .A3(n7248), .ZN(P1_U3230) );
  INV_X1 U8965 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7251) );
  OAI222_X1 U8966 ( .A1(n4454), .A2(n9834), .B1(n7781), .B2(n7252), .C1(n7251), 
        .C2(n9562), .ZN(P1_U3337) );
  INV_X1 U8967 ( .A(n7253), .ZN(n7254) );
  NAND2_X1 U8968 ( .A1(n7254), .A2(n8088), .ZN(n7255) );
  XNOR2_X1 U8969 ( .A(n7257), .B(n7090), .ZN(n7259) );
  NAND2_X1 U8970 ( .A1(n7258), .A2(n7259), .ZN(n7364) );
  INV_X1 U8971 ( .A(n7259), .ZN(n7260) );
  NAND2_X1 U8972 ( .A1(n7260), .A2(n8087), .ZN(n7261) );
  NAND2_X1 U8973 ( .A1(n7364), .A2(n7261), .ZN(n7264) );
  INV_X1 U8974 ( .A(n7264), .ZN(n7262) );
  INV_X1 U8975 ( .A(n7361), .ZN(n7263) );
  AOI21_X1 U8976 ( .B1(n7265), .B2(n7264), .A(n7263), .ZN(n7273) );
  INV_X1 U8977 ( .A(n8042), .ZN(n7953) );
  NOR2_X1 U8978 ( .A1(n7266), .A2(n10225), .ZN(n10187) );
  INV_X1 U8979 ( .A(n10187), .ZN(n7269) );
  AOI22_X1 U8980 ( .A1(n8062), .A2(n8088), .B1(n8043), .B2(n8086), .ZN(n7268)
         );
  OAI211_X1 U8981 ( .C1(n7953), .C2(n7269), .A(n7268), .B(n7267), .ZN(n7270)
         );
  AOI21_X1 U8982 ( .B1(n7271), .B2(n8067), .A(n7270), .ZN(n7272) );
  OAI21_X1 U8983 ( .B1(n7273), .B2(n8050), .A(n7272), .ZN(P2_U3170) );
  AND2_X1 U8984 ( .A1(n5133), .A2(n7274), .ZN(n9886) );
  OR2_X1 U8985 ( .A1(n9065), .A2(n7275), .ZN(n7276) );
  OAI21_X1 U8986 ( .B1(n9886), .B2(n9885), .A(n7276), .ZN(n7290) );
  XOR2_X1 U8987 ( .A(n7290), .B(n7291), .Z(n9926) );
  NAND2_X1 U8988 ( .A1(n7277), .A2(n4722), .ZN(n7288) );
  NOR2_X1 U8989 ( .A1(n9851), .A2(n7288), .ZN(n9904) );
  INV_X1 U8990 ( .A(n9904), .ZN(n7473) );
  XOR2_X1 U8991 ( .A(n7278), .B(n7291), .Z(n7280) );
  AOI222_X1 U8992 ( .A1(n9890), .A2(n7280), .B1(n9063), .B2(n9864), .C1(n9065), 
        .C2(n9996), .ZN(n9929) );
  INV_X1 U8993 ( .A(n9930), .ZN(n7283) );
  INV_X1 U8994 ( .A(n7297), .ZN(n7309) );
  AOI211_X1 U8995 ( .C1(n7283), .C2(n9899), .A(n9944), .B(n7309), .ZN(n9927)
         );
  INV_X1 U8996 ( .A(n9893), .ZN(n9852) );
  AOI22_X1 U8997 ( .A1(n9927), .A2(n9294), .B1(n9852), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7281) );
  OAI211_X1 U8998 ( .C1(n9926), .C2(n9887), .A(n9929), .B(n7281), .ZN(n7282)
         );
  NAND2_X1 U8999 ( .A1(n7282), .A2(n9238), .ZN(n7285) );
  AOI22_X1 U9000 ( .A1(n9854), .A2(n7283), .B1(P1_REG2_REG_2__SCAN_IN), .B2(
        n9851), .ZN(n7284) );
  OAI211_X1 U9001 ( .C1(n9926), .C2(n7473), .A(n7285), .B(n7284), .ZN(P1_U3291) );
  XOR2_X1 U9002 ( .A(n7286), .B(n7334), .Z(n7287) );
  AOI222_X1 U9003 ( .A1(n9890), .A2(n7287), .B1(n9062), .B2(n9864), .C1(n9063), 
        .C2(n9996), .ZN(n9946) );
  AND2_X1 U9004 ( .A1(n9887), .A2(n7288), .ZN(n7289) );
  NAND2_X1 U9005 ( .A1(n7291), .A2(n7290), .ZN(n7293) );
  NAND2_X1 U9006 ( .A1(n9882), .A2(n9930), .ZN(n7292) );
  NAND2_X1 U9007 ( .A1(n7293), .A2(n7292), .ZN(n7315) );
  NAND2_X1 U9008 ( .A1(n7315), .A2(n7316), .ZN(n7296) );
  NAND2_X1 U9009 ( .A1(n7294), .A2(n7311), .ZN(n7295) );
  NAND2_X1 U9010 ( .A1(n7296), .A2(n7295), .ZN(n7335) );
  XNOR2_X1 U9011 ( .A(n7335), .B(n7334), .ZN(n9949) );
  OR2_X1 U9012 ( .A1(n7297), .A2(n9935), .ZN(n7308) );
  AOI21_X1 U9013 ( .B1(n7298), .B2(n7308), .A(n9875), .ZN(n9942) );
  NAND2_X1 U9014 ( .A1(n9942), .A2(n9431), .ZN(n7301) );
  AOI22_X1 U9015 ( .A1(n9851), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7299), .B2(
        n9852), .ZN(n7300) );
  OAI211_X1 U9016 ( .C1(n9943), .C2(n9896), .A(n7301), .B(n7300), .ZN(n7302)
         );
  AOI21_X1 U9017 ( .B1(n9877), .B2(n9949), .A(n7302), .ZN(n7303) );
  OAI21_X1 U9018 ( .B1(n9946), .B2(n9851), .A(n7303), .ZN(P1_U3289) );
  OAI21_X1 U9019 ( .B1(n7306), .B2(n7305), .A(n7304), .ZN(n7307) );
  AOI22_X1 U9020 ( .A1(n7307), .A2(n9890), .B1(n9864), .B2(n9863), .ZN(n9938)
         );
  INV_X1 U9021 ( .A(n9380), .ZN(n9903) );
  OAI211_X1 U9022 ( .C1(n7309), .C2(n7311), .A(n9900), .B(n7308), .ZN(n9936)
         );
  INV_X1 U9023 ( .A(n9936), .ZN(n7314) );
  INV_X1 U9024 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7310) );
  OAI22_X1 U9025 ( .A1(n9238), .A2(n7310), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9893), .ZN(n7313) );
  INV_X1 U9026 ( .A(n9996), .ZN(n9883) );
  OR2_X1 U9027 ( .A1(n9907), .A2(n9883), .ZN(n9377) );
  OAI22_X1 U9028 ( .A1(n9882), .A2(n9377), .B1(n9896), .B2(n7311), .ZN(n7312)
         );
  AOI211_X1 U9029 ( .C1(n9903), .C2(n7314), .A(n7313), .B(n7312), .ZN(n7318)
         );
  XNOR2_X1 U9030 ( .A(n7316), .B(n7315), .ZN(n9940) );
  NAND2_X1 U9031 ( .A1(n9940), .A2(n9877), .ZN(n7317) );
  OAI211_X1 U9032 ( .C1(n9938), .C2(n9851), .A(n7318), .B(n7317), .ZN(P1_U3290) );
  NAND2_X1 U9033 ( .A1(n7319), .A2(n7320), .ZN(n7321) );
  XOR2_X1 U9034 ( .A(n7322), .B(n7321), .Z(n7328) );
  OAI22_X1 U9035 ( .A1(n7424), .A2(n9053), .B1(n9041), .B2(n7336), .ZN(n7326)
         );
  NOR2_X1 U9036 ( .A1(n9046), .A2(n9953), .ZN(n7325) );
  NOR2_X1 U9037 ( .A1(n9029), .A2(n9868), .ZN(n7324) );
  NAND2_X1 U9038 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9705) );
  INV_X1 U9039 ( .A(n9705), .ZN(n7323) );
  NOR4_X1 U9040 ( .A1(n7326), .A2(n7325), .A3(n7324), .A4(n7323), .ZN(n7327)
         );
  OAI21_X1 U9041 ( .B1(n7328), .B2(n9056), .A(n7327), .ZN(P1_U3227) );
  NAND2_X1 U9042 ( .A1(n7330), .A2(n7329), .ZN(n7369) );
  XNOR2_X1 U9043 ( .A(n7331), .B(n7369), .ZN(n7332) );
  INV_X1 U9044 ( .A(n7552), .ZN(n9061) );
  AOI222_X1 U9045 ( .A1(n9890), .A2(n7332), .B1(n9061), .B2(n9864), .C1(n9062), 
        .C2(n9996), .ZN(n7413) );
  NAND2_X1 U9046 ( .A1(n9875), .A2(n9953), .ZN(n9874) );
  AOI211_X1 U9047 ( .C1(n7411), .C2(n9874), .A(n9944), .B(n4953), .ZN(n7410)
         );
  AOI22_X1 U9048 ( .A1(n9851), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7353), .B2(
        n9852), .ZN(n7333) );
  OAI21_X1 U9049 ( .B1(n9896), .B2(n7371), .A(n7333), .ZN(n7342) );
  NAND2_X1 U9050 ( .A1(n7335), .A2(n7334), .ZN(n7338) );
  NAND2_X1 U9051 ( .A1(n7336), .A2(n9943), .ZN(n7337) );
  NAND2_X1 U9052 ( .A1(n7338), .A2(n7337), .ZN(n9872) );
  NAND2_X1 U9053 ( .A1(n9872), .A2(n9873), .ZN(n7340) );
  NAND2_X1 U9054 ( .A1(n7350), .A2(n9953), .ZN(n7339) );
  NAND2_X1 U9055 ( .A1(n7340), .A2(n7339), .ZN(n7370) );
  XOR2_X1 U9056 ( .A(n7370), .B(n7369), .Z(n7414) );
  NOR2_X1 U9057 ( .A1(n7414), .A2(n9415), .ZN(n7341) );
  AOI211_X1 U9058 ( .C1(n7410), .C2(n9903), .A(n7342), .B(n7341), .ZN(n7343)
         );
  OAI21_X1 U9059 ( .B1(n9907), .B2(n7413), .A(n7343), .ZN(P1_U3287) );
  XOR2_X1 U9060 ( .A(n7345), .B(n7344), .Z(n7346) );
  XNOR2_X1 U9061 ( .A(n7347), .B(n7346), .ZN(n7355) );
  INV_X1 U9062 ( .A(n9029), .ZN(n9050) );
  NAND2_X1 U9063 ( .A1(n4454), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9719) );
  INV_X1 U9064 ( .A(n9719), .ZN(n7348) );
  AOI21_X1 U9065 ( .B1(n4451), .B2(n7411), .A(n7348), .ZN(n7349) );
  INV_X1 U9066 ( .A(n7349), .ZN(n7352) );
  OAI22_X1 U9067 ( .A1(n7350), .A2(n9041), .B1(n9053), .B2(n7552), .ZN(n7351)
         );
  AOI211_X1 U9068 ( .C1(n7353), .C2(n9050), .A(n7352), .B(n7351), .ZN(n7354)
         );
  OAI21_X1 U9069 ( .B1(n7355), .B2(n9056), .A(n7354), .ZN(P1_U3239) );
  INV_X1 U9070 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7357) );
  INV_X1 U9071 ( .A(n7356), .ZN(n7358) );
  OAI222_X1 U9072 ( .A1(n9562), .A2(n7357), .B1(n7781), .B2(n7358), .C1(
        P1_U3086), .C2(n9294), .ZN(P1_U3336) );
  INV_X1 U9073 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7359) );
  OAI222_X1 U9074 ( .A1(n8888), .A2(n7359), .B1(n8890), .B2(n7358), .C1(
        P2_U3151), .C2(n8247), .ZN(P2_U3276) );
  NAND2_X1 U9075 ( .A1(n7397), .A2(n10180), .ZN(n10191) );
  AOI22_X1 U9076 ( .A1(n8062), .A2(n8087), .B1(n8043), .B2(n8085), .ZN(n7360)
         );
  NAND2_X1 U9077 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10088) );
  OAI211_X1 U9078 ( .C1(n7953), .C2(n10191), .A(n7360), .B(n10088), .ZN(n7367)
         );
  NAND2_X1 U9079 ( .A1(n7361), .A2(n7364), .ZN(n7362) );
  XNOR2_X1 U9080 ( .A(n7397), .B(n7090), .ZN(n7434) );
  XNOR2_X1 U9081 ( .A(n7434), .B(n8086), .ZN(n7363) );
  NAND3_X1 U9082 ( .A1(n7361), .A2(n4652), .A3(n7364), .ZN(n7365) );
  AOI21_X1 U9083 ( .B1(n7437), .B2(n7365), .A(n8050), .ZN(n7366) );
  AOI211_X1 U9084 ( .C1(n7396), .C2(n8067), .A(n7367), .B(n7366), .ZN(n7368)
         );
  INV_X1 U9085 ( .A(n7368), .ZN(P2_U3167) );
  NAND2_X1 U9086 ( .A1(n7370), .A2(n7369), .ZN(n7373) );
  NAND2_X1 U9087 ( .A1(n7371), .A2(n7424), .ZN(n7372) );
  NAND2_X1 U9088 ( .A1(n7373), .A2(n7372), .ZN(n7455) );
  INV_X1 U9089 ( .A(n7374), .ZN(n7461) );
  INV_X1 U9090 ( .A(n7460), .ZN(n7376) );
  XNOR2_X1 U9091 ( .A(n7455), .B(n7376), .ZN(n7381) );
  XNOR2_X1 U9092 ( .A(n7377), .B(n7460), .ZN(n7379) );
  OAI22_X1 U9093 ( .A1(n7424), .A2(n9883), .B1(n7647), .B2(n9881), .ZN(n7378)
         );
  AOI21_X1 U9094 ( .B1(n7379), .B2(n9890), .A(n7378), .ZN(n7380) );
  OAI21_X1 U9095 ( .B1(n7381), .B2(n9887), .A(n7380), .ZN(n9959) );
  INV_X1 U9096 ( .A(n9959), .ZN(n7388) );
  INV_X1 U9097 ( .A(n7381), .ZN(n9961) );
  INV_X1 U9098 ( .A(n7456), .ZN(n9958) );
  INV_X1 U9099 ( .A(n7467), .ZN(n7383) );
  OAI211_X1 U9100 ( .C1(n9958), .C2(n4953), .A(n7383), .B(n9900), .ZN(n9957)
         );
  OR2_X1 U9101 ( .A1(n9907), .A2(n4722), .ZN(n9223) );
  AOI22_X1 U9102 ( .A1(n9851), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7427), .B2(
        n9852), .ZN(n7385) );
  NAND2_X1 U9103 ( .A1(n9854), .A2(n7456), .ZN(n7384) );
  OAI211_X1 U9104 ( .C1(n9957), .C2(n9223), .A(n7385), .B(n7384), .ZN(n7386)
         );
  AOI21_X1 U9105 ( .B1(n9961), .B2(n9904), .A(n7386), .ZN(n7387) );
  OAI21_X1 U9106 ( .B1(n7388), .B2(n9851), .A(n7387), .ZN(P1_U3286) );
  INV_X1 U9107 ( .A(n7389), .ZN(n7392) );
  XNOR2_X1 U9108 ( .A(n7390), .B(n7392), .ZN(n7395) );
  XNOR2_X1 U9109 ( .A(n7391), .B(n7392), .ZN(n10190) );
  INV_X1 U9110 ( .A(n10163), .ZN(n10207) );
  NAND2_X1 U9111 ( .A1(n10190), .A2(n10207), .ZN(n7394) );
  AOI22_X1 U9112 ( .A1(n8435), .A2(n8087), .B1(n8085), .B2(n8437), .ZN(n7393)
         );
  OAI211_X1 U9113 ( .C1(n7395), .C2(n8451), .A(n7394), .B(n7393), .ZN(n10194)
         );
  INV_X1 U9114 ( .A(n10194), .ZN(n7402) );
  NAND2_X1 U9115 ( .A1(n10167), .A2(n10166), .ZN(n8264) );
  INV_X1 U9116 ( .A(n8264), .ZN(n7400) );
  INV_X1 U9117 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10076) );
  AOI22_X1 U9118 ( .A1(n8429), .A2(n7397), .B1(n8440), .B2(n7396), .ZN(n7398)
         );
  OAI21_X1 U9119 ( .B1(n10076), .B2(n10167), .A(n7398), .ZN(n7399) );
  AOI21_X1 U9120 ( .B1(n10190), .B2(n7400), .A(n7399), .ZN(n7401) );
  OAI21_X1 U9121 ( .B1(n7402), .B2(n8442), .A(n7401), .ZN(P2_U3228) );
  XOR2_X1 U9122 ( .A(n7403), .B(n7406), .Z(n7404) );
  AOI222_X1 U9123 ( .A1(n6797), .A2(n7404), .B1(n8084), .B2(n8437), .C1(n8086), 
        .C2(n8435), .ZN(n10196) );
  XOR2_X1 U9124 ( .A(n7405), .B(n7406), .Z(n10199) );
  INV_X1 U9125 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7599) );
  AOI22_X1 U9126 ( .A1(n8429), .A2(n7438), .B1(n8440), .B2(n8044), .ZN(n7407)
         );
  OAI21_X1 U9127 ( .B1(n7599), .B2(n10167), .A(n7407), .ZN(n7408) );
  AOI21_X1 U9128 ( .B1(n10199), .B2(n8461), .A(n7408), .ZN(n7409) );
  OAI21_X1 U9129 ( .B1(n10196), .B2(n8442), .A(n7409), .ZN(P2_U3227) );
  INV_X1 U9130 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n8770) );
  INV_X1 U9131 ( .A(n10009), .ZN(n9528) );
  AOI21_X1 U9132 ( .B1(n9997), .B2(n7411), .A(n7410), .ZN(n7412) );
  OAI211_X1 U9133 ( .C1(n9528), .C2(n7414), .A(n7413), .B(n7412), .ZN(n7416)
         );
  NAND2_X1 U9134 ( .A1(n7416), .A2(n10013), .ZN(n7415) );
  OAI21_X1 U9135 ( .B1(n10013), .B2(n8770), .A(n7415), .ZN(P1_U3471) );
  NAND2_X1 U9136 ( .A1(n7416), .A2(n10033), .ZN(n7417) );
  OAI21_X1 U9137 ( .B1(n10033), .B2(n6943), .A(n7417), .ZN(P1_U3528) );
  NAND2_X1 U9138 ( .A1(n7419), .A2(n7418), .ZN(n7421) );
  XOR2_X1 U9139 ( .A(n7421), .B(n7420), .Z(n7429) );
  NAND2_X1 U9140 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9591) );
  INV_X1 U9141 ( .A(n9591), .ZN(n7422) );
  AOI21_X1 U9142 ( .B1(n4451), .B2(n7456), .A(n7422), .ZN(n7423) );
  INV_X1 U9143 ( .A(n7423), .ZN(n7426) );
  OAI22_X1 U9144 ( .A1(n7424), .A2(n9041), .B1(n9053), .B2(n7647), .ZN(n7425)
         );
  AOI211_X1 U9145 ( .C1(n7427), .C2(n9050), .A(n7426), .B(n7425), .ZN(n7428)
         );
  OAI21_X1 U9146 ( .B1(n7429), .B2(n9056), .A(n7428), .ZN(P1_U3213) );
  INV_X1 U9147 ( .A(n7430), .ZN(n7432) );
  OAI222_X1 U9148 ( .A1(n8890), .A2(n7432), .B1(n7431), .B2(P2_U3151), .C1(
        n8625), .C2(n8888), .ZN(P2_U3275) );
  OAI222_X1 U9149 ( .A1(P1_U3086), .A2(n7433), .B1(n7781), .B2(n7432), .C1(
        n8776), .C2(n9562), .ZN(P1_U3335) );
  NAND2_X1 U9150 ( .A1(n7435), .A2(n7434), .ZN(n7436) );
  XNOR2_X1 U9151 ( .A(n7438), .B(n7090), .ZN(n7439) );
  XNOR2_X1 U9152 ( .A(n7439), .B(n8085), .ZN(n8038) );
  INV_X1 U9153 ( .A(n7439), .ZN(n7440) );
  XNOR2_X1 U9154 ( .A(n7447), .B(n7090), .ZN(n7441) );
  NAND2_X1 U9155 ( .A1(n7530), .A2(n7441), .ZN(n7535) );
  OAI21_X1 U9156 ( .B1(n7530), .B2(n7441), .A(n7535), .ZN(n7445) );
  INV_X1 U9157 ( .A(n7446), .ZN(n7443) );
  NAND2_X1 U9158 ( .A1(n7443), .A2(n7442), .ZN(n7531) );
  INV_X1 U9159 ( .A(n7531), .ZN(n7444) );
  AOI21_X1 U9160 ( .B1(n7446), .B2(n7445), .A(n7444), .ZN(n7454) );
  NAND2_X1 U9161 ( .A1(n8033), .A2(n7447), .ZN(n7450) );
  NAND2_X1 U9162 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10125) );
  INV_X1 U9163 ( .A(n10125), .ZN(n7448) );
  AOI21_X1 U9164 ( .B1(n8043), .B2(n8083), .A(n7448), .ZN(n7449) );
  OAI211_X1 U9165 ( .C1(n7451), .C2(n8031), .A(n7450), .B(n7449), .ZN(n7452)
         );
  AOI21_X1 U9166 ( .B1(n8067), .B2(n7475), .A(n7452), .ZN(n7453) );
  OAI21_X1 U9167 ( .B1(n7454), .B2(n8050), .A(n7453), .ZN(P2_U3153) );
  NAND2_X1 U9168 ( .A1(n7455), .A2(n7460), .ZN(n7458) );
  OR2_X1 U9169 ( .A1(n7456), .A2(n9061), .ZN(n7457) );
  NAND2_X1 U9170 ( .A1(n7500), .A2(n7459), .ZN(n7484) );
  XNOR2_X1 U9171 ( .A(n7485), .B(n4747), .ZN(n9963) );
  NOR2_X1 U9172 ( .A1(n7377), .A2(n7460), .ZN(n7502) );
  NOR2_X1 U9173 ( .A1(n7502), .A2(n7461), .ZN(n7462) );
  XNOR2_X1 U9174 ( .A(n7462), .B(n7484), .ZN(n7464) );
  OAI22_X1 U9175 ( .A1(n7552), .A2(n9883), .B1(n8926), .B2(n9881), .ZN(n7463)
         );
  AOI21_X1 U9176 ( .B1(n7464), .B2(n9890), .A(n7463), .ZN(n7465) );
  OAI21_X1 U9177 ( .B1(n9963), .B2(n9887), .A(n7465), .ZN(n9966) );
  NAND2_X1 U9178 ( .A1(n9966), .A2(n9238), .ZN(n7472) );
  INV_X1 U9179 ( .A(n7466), .ZN(n7551) );
  OAI22_X1 U9180 ( .A1(n9238), .A2(n8788), .B1(n7551), .B2(n9893), .ZN(n7469)
         );
  OAI211_X1 U9181 ( .C1(n9965), .C2(n7467), .A(n4540), .B(n9900), .ZN(n9964)
         );
  NOR2_X1 U9182 ( .A1(n9964), .A2(n9380), .ZN(n7468) );
  AOI211_X1 U9183 ( .C1(n9854), .C2(n7470), .A(n7469), .B(n7468), .ZN(n7471)
         );
  OAI211_X1 U9184 ( .C1(n9963), .C2(n7473), .A(n7472), .B(n7471), .ZN(P1_U3285) );
  INV_X1 U9185 ( .A(n7521), .ZN(n7474) );
  AOI21_X1 U9186 ( .B1(n4543), .B2(n7479), .A(n7474), .ZN(n10206) );
  INV_X1 U9187 ( .A(n10206), .ZN(n10203) );
  INV_X1 U9188 ( .A(n7475), .ZN(n7476) );
  OAI22_X1 U9189 ( .A1(n8411), .A2(n10201), .B1(n7476), .B2(n10151), .ZN(n7477) );
  AOI21_X1 U9190 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n8442), .A(n7477), .ZN(
        n7483) );
  OAI211_X1 U9191 ( .C1(n4544), .C2(n7479), .A(n7478), .B(n6797), .ZN(n7481)
         );
  AOI22_X1 U9192 ( .A1(n8083), .A2(n8437), .B1(n8435), .B2(n8085), .ZN(n7480)
         );
  NAND2_X1 U9193 ( .A1(n7481), .A2(n7480), .ZN(n10204) );
  NAND2_X1 U9194 ( .A1(n10204), .A2(n10167), .ZN(n7482) );
  OAI211_X1 U9195 ( .C1(n10203), .C2(n8447), .A(n7483), .B(n7482), .ZN(
        P2_U3226) );
  NOR2_X1 U9196 ( .A1(n7487), .A2(n7486), .ZN(n7509) );
  XNOR2_X1 U9197 ( .A(n7588), .B(n7587), .ZN(n9985) );
  INV_X1 U9198 ( .A(n9985), .ZN(n7499) );
  INV_X1 U9199 ( .A(n9842), .ZN(n7488) );
  AOI21_X1 U9200 ( .B1(n7587), .B2(n7489), .A(n7488), .ZN(n7490) );
  OAI22_X1 U9201 ( .A1(n7490), .A2(n9420), .B1(n7740), .B2(n9881), .ZN(n9983)
         );
  AOI21_X1 U9202 ( .B1(n4542), .B2(n9980), .A(n9944), .ZN(n7491) );
  NAND2_X1 U9203 ( .A1(n7491), .A2(n9856), .ZN(n9982) );
  NOR2_X1 U9204 ( .A1(n9893), .A2(n7492), .ZN(n7493) );
  AOI21_X1 U9205 ( .B1(n9907), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7493), .ZN(
        n7494) );
  OAI21_X1 U9206 ( .B1(n9377), .B2(n8926), .A(n7494), .ZN(n7495) );
  AOI21_X1 U9207 ( .B1(n9980), .B2(n9854), .A(n7495), .ZN(n7496) );
  OAI21_X1 U9208 ( .B1(n9982), .B2(n9380), .A(n7496), .ZN(n7497) );
  AOI21_X1 U9209 ( .B1(n9983), .B2(n9238), .A(n7497), .ZN(n7498) );
  OAI21_X1 U9210 ( .B1(n7499), .B2(n9415), .A(n7498), .ZN(P1_U3283) );
  OAI21_X1 U9211 ( .B1(n7502), .B2(n7501), .A(n7500), .ZN(n7503) );
  XOR2_X1 U9212 ( .A(n7509), .B(n7503), .Z(n7504) );
  NAND2_X1 U9213 ( .A1(n7504), .A2(n9890), .ZN(n9975) );
  AOI22_X1 U9214 ( .A1(n9907), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7648), .B2(
        n9852), .ZN(n7505) );
  OAI21_X1 U9215 ( .B1(n9377), .B2(n7647), .A(n7505), .ZN(n7508) );
  AOI21_X1 U9216 ( .B1(n4540), .B2(n9972), .A(n9944), .ZN(n7506) );
  AOI22_X1 U9217 ( .A1(n7506), .A2(n4542), .B1(n9864), .B2(n9060), .ZN(n9974)
         );
  NOR2_X1 U9218 ( .A1(n9974), .A2(n9380), .ZN(n7507) );
  AOI211_X1 U9219 ( .C1(n9854), .C2(n9972), .A(n7508), .B(n7507), .ZN(n7512)
         );
  XNOR2_X1 U9220 ( .A(n7510), .B(n7509), .ZN(n9977) );
  NAND2_X1 U9221 ( .A1(n9977), .A2(n9877), .ZN(n7511) );
  OAI211_X1 U9222 ( .C1(n9975), .C2(n9851), .A(n7512), .B(n7511), .ZN(P1_U3284) );
  INV_X1 U9223 ( .A(n7513), .ZN(n7516) );
  OAI222_X1 U9224 ( .A1(n8890), .A2(n7516), .B1(n6488), .B2(P2_U3151), .C1(
        n7514), .C2(n8888), .ZN(P2_U3274) );
  OAI222_X1 U9225 ( .A1(n9562), .A2(n7517), .B1(n7781), .B2(n7516), .C1(n7515), 
        .C2(n4454), .ZN(P1_U3334) );
  XOR2_X1 U9226 ( .A(n7518), .B(n7522), .Z(n7519) );
  AOI222_X1 U9227 ( .A1(n6797), .A2(n7519), .B1(n8082), .B2(n8437), .C1(n8084), 
        .C2(n8435), .ZN(n10209) );
  NAND2_X1 U9228 ( .A1(n7521), .A2(n7520), .ZN(n7523) );
  XNOR2_X1 U9229 ( .A(n7523), .B(n7522), .ZN(n10212) );
  AOI22_X1 U9230 ( .A1(n8442), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n8440), .B2(
        n7539), .ZN(n7524) );
  OAI21_X1 U9231 ( .B1(n7532), .B2(n8411), .A(n7524), .ZN(n7525) );
  AOI21_X1 U9232 ( .B1(n10212), .B2(n8461), .A(n7525), .ZN(n7526) );
  OAI21_X1 U9233 ( .B1(n10209), .B2(n8442), .A(n7526), .ZN(P2_U3225) );
  INV_X1 U9234 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7527) );
  NOR2_X1 U9235 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7527), .ZN(n10138) );
  AOI21_X1 U9236 ( .B1(n8043), .B2(n8082), .A(n10138), .ZN(n7529) );
  NOR2_X1 U9237 ( .A1(n7532), .A2(n10225), .ZN(n10211) );
  NAND2_X1 U9238 ( .A1(n8042), .A2(n10211), .ZN(n7528) );
  OAI211_X1 U9239 ( .C1(n7530), .C2(n8031), .A(n7529), .B(n7528), .ZN(n7538)
         );
  NAND2_X1 U9240 ( .A1(n7531), .A2(n7535), .ZN(n7533) );
  XNOR2_X1 U9241 ( .A(n7532), .B(n7090), .ZN(n7557) );
  XNOR2_X1 U9242 ( .A(n7557), .B(n7558), .ZN(n7534) );
  NAND3_X1 U9243 ( .A1(n7531), .A2(n4648), .A3(n7535), .ZN(n7536) );
  AOI21_X1 U9244 ( .B1(n7561), .B2(n7536), .A(n8050), .ZN(n7537) );
  AOI211_X1 U9245 ( .C1(n7539), .C2(n8067), .A(n7538), .B(n7537), .ZN(n7540)
         );
  INV_X1 U9246 ( .A(n7540), .ZN(P2_U3161) );
  INV_X1 U9247 ( .A(n7541), .ZN(n7545) );
  OAI222_X1 U9248 ( .A1(n8888), .A2(n7543), .B1(n8890), .B2(n7545), .C1(
        P2_U3151), .C2(n7542), .ZN(P2_U3273) );
  OAI222_X1 U9249 ( .A1(n9562), .A2(n7546), .B1(n7781), .B2(n7545), .C1(
        P1_U3086), .C2(n7544), .ZN(P1_U3333) );
  OAI21_X1 U9250 ( .B1(n7549), .B2(n7548), .A(n7547), .ZN(n7550) );
  NAND2_X1 U9251 ( .A1(n7550), .A2(n9038), .ZN(n7556) );
  NAND2_X1 U9252 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9620) );
  INV_X1 U9253 ( .A(n9620), .ZN(n7554) );
  OAI22_X1 U9254 ( .A1(n9041), .A2(n7552), .B1(n9029), .B2(n7551), .ZN(n7553)
         );
  AOI211_X1 U9255 ( .C1(n9021), .C2(n9979), .A(n7554), .B(n7553), .ZN(n7555)
         );
  OAI211_X1 U9256 ( .C1(n9965), .C2(n9046), .A(n7556), .B(n7555), .ZN(P1_U3221) );
  NOR2_X1 U9257 ( .A1(n7562), .A2(n10225), .ZN(n10216) );
  INV_X1 U9258 ( .A(n10216), .ZN(n7568) );
  INV_X1 U9259 ( .A(n7557), .ZN(n7559) );
  NAND2_X1 U9260 ( .A1(n7559), .A2(n7558), .ZN(n7560) );
  XNOR2_X1 U9261 ( .A(n7562), .B(n7090), .ZN(n7829) );
  XNOR2_X1 U9262 ( .A(n7829), .B(n7714), .ZN(n7563) );
  OAI211_X1 U9263 ( .C1(n4545), .C2(n7563), .A(n7830), .B(n8058), .ZN(n7567)
         );
  AND2_X1 U9264 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7637) );
  AOI21_X1 U9265 ( .B1(n8062), .B2(n8083), .A(n7637), .ZN(n7564) );
  OAI21_X1 U9266 ( .B1(n7832), .B2(n8064), .A(n7564), .ZN(n7565) );
  AOI21_X1 U9267 ( .B1(n8067), .B2(n7577), .A(n7565), .ZN(n7566) );
  OAI211_X1 U9268 ( .C1(n7953), .C2(n7568), .A(n7567), .B(n7566), .ZN(P2_U3171) );
  NAND2_X1 U9269 ( .A1(n7570), .A2(n7573), .ZN(n7571) );
  NAND2_X1 U9270 ( .A1(n7569), .A2(n7571), .ZN(n10214) );
  XOR2_X1 U9271 ( .A(n7572), .B(n7573), .Z(n7574) );
  NAND2_X1 U9272 ( .A1(n7574), .A2(n6797), .ZN(n7576) );
  AOI22_X1 U9273 ( .A1(n8083), .A2(n8435), .B1(n8437), .B2(n8081), .ZN(n7575)
         );
  OAI211_X1 U9274 ( .C1(n10163), .C2(n10214), .A(n7576), .B(n7575), .ZN(n10215) );
  NAND2_X1 U9275 ( .A1(n10215), .A2(n10167), .ZN(n7582) );
  INV_X1 U9276 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7606) );
  INV_X1 U9277 ( .A(n7577), .ZN(n7578) );
  OAI22_X1 U9278 ( .A1(n10167), .A2(n7606), .B1(n7578), .B2(n10151), .ZN(n7579) );
  AOI21_X1 U9279 ( .B1(n8429), .B2(n7580), .A(n7579), .ZN(n7581) );
  OAI211_X1 U9280 ( .C1(n10214), .C2(n8264), .A(n7582), .B(n7581), .ZN(
        P2_U3224) );
  OAI21_X1 U9281 ( .B1(n7744), .B2(n7584), .A(n7583), .ZN(n7585) );
  INV_X1 U9282 ( .A(n9422), .ZN(n9150) );
  INV_X1 U9283 ( .A(n9844), .ZN(n9059) );
  AOI222_X1 U9284 ( .A1(n9890), .A2(n7585), .B1(n9150), .B2(n9864), .C1(n9059), 
        .C2(n9996), .ZN(n10006) );
  INV_X1 U9285 ( .A(n9998), .ZN(n7696) );
  XNOR2_X1 U9286 ( .A(n7745), .B(n7744), .ZN(n10010) );
  NAND2_X1 U9287 ( .A1(n10010), .A2(n9877), .ZN(n7593) );
  NOR2_X2 U9288 ( .A1(n9856), .A2(n9988), .ZN(n9855) );
  AND2_X2 U9289 ( .A1(n9855), .A2(n7696), .ZN(n7694) );
  OAI211_X1 U9290 ( .C1(n7694), .C2(n4774), .A(n9900), .B(n7747), .ZN(n10005)
         );
  INV_X1 U9291 ( .A(n10005), .ZN(n7591) );
  INV_X1 U9292 ( .A(n9223), .ZN(n9413) );
  AOI22_X1 U9293 ( .A1(n9851), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8998), .B2(
        n9852), .ZN(n7589) );
  OAI21_X1 U9294 ( .B1(n4774), .B2(n9896), .A(n7589), .ZN(n7590) );
  AOI21_X1 U9295 ( .B1(n7591), .B2(n9413), .A(n7590), .ZN(n7592) );
  OAI211_X1 U9296 ( .C1(n9907), .C2(n10006), .A(n7593), .B(n7592), .ZN(
        P1_U3280) );
  INV_X1 U9297 ( .A(n7594), .ZN(n7595) );
  NAND2_X1 U9298 ( .A1(n7597), .A2(n10078), .ZN(n7596) );
  INV_X1 U9299 ( .A(n7596), .ZN(n7598) );
  AOI22_X1 U9300 ( .A1(n10100), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n7599), .B2(
        n7626), .ZN(n10094) );
  NOR2_X1 U9301 ( .A1(n10100), .A2(n7599), .ZN(n7600) );
  NAND2_X1 U9302 ( .A1(n7602), .A2(n10111), .ZN(n7601) );
  INV_X1 U9303 ( .A(n7601), .ZN(n7603) );
  INV_X1 U9304 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10109) );
  OAI21_X1 U9305 ( .B1(n7602), .B2(n10111), .A(n7601), .ZN(n10110) );
  INV_X1 U9306 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7604) );
  AOI22_X1 U9307 ( .A1(n10140), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n7604), .B2(
        n7629), .ZN(n10128) );
  AOI21_X1 U9308 ( .B1(n7606), .B2(n7605), .A(n7661), .ZN(n7640) );
  INV_X1 U9309 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10256) );
  INV_X1 U9310 ( .A(n7611), .ZN(n7609) );
  INV_X1 U9311 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10248) );
  INV_X1 U9312 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10250) );
  AOI22_X1 U9313 ( .A1(n10100), .A2(P2_REG1_REG_6__SCAN_IN), .B1(n10250), .B2(
        n7626), .ZN(n10091) );
  NOR2_X1 U9314 ( .A1(n10092), .A2(n10091), .ZN(n10090) );
  NOR2_X1 U9315 ( .A1(n10100), .A2(n10250), .ZN(n7613) );
  INV_X1 U9316 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10252) );
  INV_X1 U9317 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10254) );
  AOI22_X1 U9318 ( .A1(n10140), .A2(P2_REG1_REG_8__SCAN_IN), .B1(n10254), .B2(
        n7629), .ZN(n10131) );
  AOI21_X1 U9319 ( .B1(n10256), .B2(n7616), .A(n7667), .ZN(n7617) );
  NOR2_X1 U9320 ( .A1(n7617), .A2(n10133), .ZN(n7638) );
  INV_X1 U9321 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n8644) );
  INV_X1 U9322 ( .A(n10115), .ZN(n10148) );
  OAI22_X1 U9323 ( .A1(n10112), .A2(n7618), .B1(n8644), .B2(n10148), .ZN(n7636) );
  MUX2_X1 U9324 ( .A(n7606), .B(n10256), .S(n8241), .Z(n7620) );
  AND2_X1 U9325 ( .A1(n7620), .A2(n7666), .ZN(n7675) );
  INV_X1 U9326 ( .A(n7675), .ZN(n7619) );
  OAI21_X1 U9327 ( .B1(n7666), .B2(n7620), .A(n7619), .ZN(n7633) );
  MUX2_X1 U9328 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n6509), .Z(n7630) );
  NOR2_X1 U9329 ( .A1(n7630), .A2(n7629), .ZN(n7631) );
  MUX2_X1 U9330 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8241), .Z(n7628) );
  MUX2_X1 U9331 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8241), .Z(n7627) );
  INV_X1 U9332 ( .A(n7621), .ZN(n7623) );
  MUX2_X1 U9333 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8241), .Z(n7625) );
  XNOR2_X1 U9334 ( .A(n7625), .B(n4845), .ZN(n10082) );
  XNOR2_X1 U9335 ( .A(n7627), .B(n10100), .ZN(n10102) );
  NAND2_X1 U9336 ( .A1(n10103), .A2(n10102), .ZN(n10101) );
  OAI21_X1 U9337 ( .B1(n7627), .B2(n7626), .A(n10101), .ZN(n10118) );
  XOR2_X1 U9338 ( .A(n10111), .B(n7628), .Z(n10117) );
  NAND2_X1 U9339 ( .A1(n10118), .A2(n10117), .ZN(n10116) );
  OAI21_X1 U9340 ( .B1(n7628), .B2(n10111), .A(n10116), .ZN(n10142) );
  AOI21_X1 U9341 ( .B1(n7630), .B2(n7629), .A(n7631), .ZN(n10141) );
  NOR2_X1 U9342 ( .A1(n7631), .A2(n10145), .ZN(n7632) );
  AOI21_X1 U9343 ( .B1(n7633), .B2(n7632), .A(n7674), .ZN(n7634) );
  NOR2_X1 U9344 ( .A1(n7634), .A2(n8250), .ZN(n7635) );
  NOR4_X1 U9345 ( .A1(n7638), .A2(n7637), .A3(n7636), .A4(n7635), .ZN(n7639)
         );
  OAI21_X1 U9346 ( .B1(n7640), .B2(n10135), .A(n7639), .ZN(P2_U3191) );
  INV_X1 U9347 ( .A(n7656), .ZN(n7643) );
  NAND2_X1 U9348 ( .A1(n8884), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7641) );
  OAI211_X1 U9349 ( .C1(n7643), .C2(n8890), .A(n7642), .B(n7641), .ZN(P2_U3272) );
  XNOR2_X1 U9350 ( .A(n7644), .B(n7645), .ZN(n7646) );
  NAND2_X1 U9351 ( .A1(n7646), .A2(n9038), .ZN(n7653) );
  INV_X1 U9352 ( .A(n7647), .ZN(n9971) );
  INV_X1 U9353 ( .A(n7648), .ZN(n7649) );
  OAI22_X1 U9354 ( .A1(n9053), .A2(n9845), .B1(n9029), .B2(n7649), .ZN(n7650)
         );
  AOI211_X1 U9355 ( .C1(n9051), .C2(n9971), .A(n7651), .B(n7650), .ZN(n7652)
         );
  OAI211_X1 U9356 ( .C1(n7654), .C2(n9046), .A(n7653), .B(n7652), .ZN(P1_U3231) );
  NAND2_X1 U9357 ( .A1(n7656), .A2(n7655), .ZN(n7658) );
  OAI211_X1 U9358 ( .C1(n7659), .C2(n9562), .A(n7658), .B(n7657), .ZN(P1_U3332) );
  NOR2_X1 U9359 ( .A1(n7666), .A2(n7660), .ZN(n7662) );
  INV_X1 U9360 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8638) );
  AOI22_X1 U9361 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7678), .B1(n7763), .B2(
        n8638), .ZN(n7663) );
  AOI21_X1 U9362 ( .B1(n7664), .B2(n7663), .A(n7758), .ZN(n7686) );
  NOR2_X1 U9363 ( .A1(n7666), .A2(n7665), .ZN(n7668) );
  INV_X1 U9364 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10258) );
  AOI22_X1 U9365 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7678), .B1(n7763), .B2(
        n10258), .ZN(n7669) );
  AOI21_X1 U9366 ( .B1(n7670), .B2(n7669), .A(n7762), .ZN(n7671) );
  NOR2_X1 U9367 ( .A1(n7671), .A2(n10133), .ZN(n7684) );
  MUX2_X1 U9368 ( .A(n8638), .B(n10258), .S(n6509), .Z(n7673) );
  AND2_X1 U9369 ( .A1(n7673), .A2(n7678), .ZN(n7769) );
  INV_X1 U9370 ( .A(n7769), .ZN(n7672) );
  OAI21_X1 U9371 ( .B1(n7678), .B2(n7673), .A(n7672), .ZN(n7677) );
  NOR2_X1 U9372 ( .A1(n7676), .A2(n7677), .ZN(n7768) );
  AOI21_X1 U9373 ( .B1(n7677), .B2(n7676), .A(n7768), .ZN(n7682) );
  AOI22_X1 U9374 ( .A1(n10139), .A2(n7678), .B1(n10115), .B2(
        P2_ADDR_REG_10__SCAN_IN), .ZN(n7681) );
  INV_X1 U9375 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7679) );
  NOR2_X1 U9376 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7679), .ZN(n7906) );
  INV_X1 U9377 ( .A(n7906), .ZN(n7680) );
  OAI211_X1 U9378 ( .C1(n7682), .C2(n8250), .A(n7681), .B(n7680), .ZN(n7683)
         );
  NOR2_X1 U9379 ( .A1(n7684), .A2(n7683), .ZN(n7685) );
  OAI21_X1 U9380 ( .B1(n7686), .B2(n10135), .A(n7685), .ZN(P2_U3192) );
  NAND2_X1 U9381 ( .A1(n7688), .A2(n7687), .ZN(n7689) );
  XNOR2_X1 U9382 ( .A(n7689), .B(n7691), .ZN(n7690) );
  INV_X1 U9383 ( .A(n8909), .ZN(n9058) );
  AOI22_X1 U9384 ( .A1(n7690), .A2(n9890), .B1(n9864), .B2(n9058), .ZN(n10001)
         );
  XNOR2_X1 U9385 ( .A(n7692), .B(n7691), .ZN(n10003) );
  NAND2_X1 U9386 ( .A1(n10003), .A2(n9877), .ZN(n7700) );
  AOI22_X1 U9387 ( .A1(n9907), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7738), .B2(
        n9852), .ZN(n7693) );
  OAI21_X1 U9388 ( .B1(n9377), .B2(n7740), .A(n7693), .ZN(n7698) );
  INV_X1 U9389 ( .A(n7694), .ZN(n7695) );
  OAI211_X1 U9390 ( .C1(n7696), .C2(n9855), .A(n7695), .B(n9900), .ZN(n9999)
         );
  NOR2_X1 U9391 ( .A1(n9999), .A2(n9380), .ZN(n7697) );
  AOI211_X1 U9392 ( .C1(n9854), .C2(n9998), .A(n7698), .B(n7697), .ZN(n7699)
         );
  OAI211_X1 U9393 ( .C1(n9907), .C2(n10001), .A(n7700), .B(n7699), .ZN(
        P1_U3281) );
  XNOR2_X1 U9394 ( .A(n7701), .B(n7706), .ZN(n7704) );
  NAND2_X1 U9395 ( .A1(n8436), .A2(n8437), .ZN(n7702) );
  OAI21_X1 U9396 ( .B1(n7908), .B2(n10157), .A(n7702), .ZN(n7703) );
  AOI21_X1 U9397 ( .B1(n7704), .B2(n6797), .A(n7703), .ZN(n10237) );
  XNOR2_X1 U9398 ( .A(n7705), .B(n7706), .ZN(n10235) );
  AOI22_X1 U9399 ( .A1(n8442), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n8440), .B2(
        n7950), .ZN(n7707) );
  OAI21_X1 U9400 ( .B1(n7708), .B2(n8411), .A(n7707), .ZN(n7709) );
  AOI21_X1 U9401 ( .B1(n10235), .B2(n8461), .A(n7709), .ZN(n7710) );
  OAI21_X1 U9402 ( .B1(n10237), .B2(n8442), .A(n7710), .ZN(P2_U3221) );
  NAND2_X1 U9403 ( .A1(n7711), .A2(n7727), .ZN(n7716) );
  XOR2_X1 U9404 ( .A(n7716), .B(n7712), .Z(n7713) );
  OAI222_X1 U9405 ( .A1(n10158), .A2(n7908), .B1(n10157), .B2(n7714), .C1(
        n8451), .C2(n7713), .ZN(n10221) );
  INV_X1 U9406 ( .A(n10221), .ZN(n7722) );
  NAND2_X1 U9407 ( .A1(n7569), .A2(n7715), .ZN(n7717) );
  XNOR2_X1 U9408 ( .A(n7717), .B(n7716), .ZN(n10223) );
  AOI22_X1 U9409 ( .A1(n8442), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n8440), .B2(
        n7910), .ZN(n7718) );
  OAI21_X1 U9410 ( .B1(n7719), .B2(n8411), .A(n7718), .ZN(n7720) );
  AOI21_X1 U9411 ( .B1(n10223), .B2(n8461), .A(n7720), .ZN(n7721) );
  OAI21_X1 U9412 ( .B1(n7722), .B2(n8442), .A(n7721), .ZN(P2_U3223) );
  INV_X1 U9413 ( .A(n7723), .ZN(n7725) );
  OAI222_X1 U9414 ( .A1(n7757), .A2(n7725), .B1(P2_U3151), .B2(n6801), .C1(
        n8647), .C2(n8888), .ZN(P2_U3271) );
  OAI222_X1 U9415 ( .A1(n7726), .A2(n4454), .B1(n7781), .B2(n7725), .C1(n7724), 
        .C2(n9562), .ZN(P1_U3331) );
  NAND2_X1 U9416 ( .A1(n7728), .A2(n7727), .ZN(n7729) );
  XNOR2_X1 U9417 ( .A(n7729), .B(n7834), .ZN(n10228) );
  XNOR2_X1 U9418 ( .A(n7730), .B(n7834), .ZN(n7731) );
  OAI222_X1 U9419 ( .A1(n10158), .A2(n8454), .B1(n10157), .B2(n7832), .C1(
        n7731), .C2(n8451), .ZN(n10230) );
  NAND2_X1 U9420 ( .A1(n10230), .A2(n10167), .ZN(n7735) );
  INV_X1 U9421 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7761) );
  INV_X1 U9422 ( .A(n8023), .ZN(n7732) );
  OAI22_X1 U9423 ( .A1(n10167), .A2(n7761), .B1(n7732), .B2(n10151), .ZN(n7733) );
  AOI21_X1 U9424 ( .B1(n8015), .B2(n8429), .A(n7733), .ZN(n7734) );
  OAI211_X1 U9425 ( .C1(n8447), .C2(n10228), .A(n7735), .B(n7734), .ZN(
        P2_U3222) );
  XOR2_X1 U9426 ( .A(n7736), .B(n7737), .Z(n7743) );
  AOI22_X1 U9427 ( .A1(n9021), .A2(n9058), .B1(n9050), .B2(n7738), .ZN(n7739)
         );
  NAND2_X1 U9428 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(n4454), .ZN(n9750) );
  OAI211_X1 U9429 ( .C1(n7740), .C2(n9041), .A(n7739), .B(n9750), .ZN(n7741)
         );
  AOI21_X1 U9430 ( .B1(n9998), .B2(n4451), .A(n7741), .ZN(n7742) );
  OAI21_X1 U9431 ( .B1(n7743), .B2(n9056), .A(n7742), .ZN(P1_U3224) );
  XNOR2_X1 U9432 ( .A(n9151), .B(n7749), .ZN(n9529) );
  INV_X1 U9433 ( .A(n9427), .ZN(n7746) );
  AOI21_X1 U9434 ( .B1(n9524), .B2(n7747), .A(n7746), .ZN(n9525) );
  AOI22_X1 U9435 ( .A1(n9851), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8907), .B2(
        n9852), .ZN(n7748) );
  OAI21_X1 U9436 ( .B1(n4951), .B2(n9896), .A(n7748), .ZN(n7753) );
  XNOR2_X1 U9437 ( .A(n7750), .B(n7749), .ZN(n7751) );
  INV_X1 U9438 ( .A(n9152), .ZN(n9409) );
  AOI222_X1 U9439 ( .A1(n9890), .A2(n7751), .B1(n9058), .B2(n9996), .C1(n9409), 
        .C2(n9864), .ZN(n9527) );
  NOR2_X1 U9440 ( .A1(n9527), .A2(n9851), .ZN(n7752) );
  AOI211_X1 U9441 ( .C1(n9525), .C2(n9431), .A(n7753), .B(n7752), .ZN(n7754)
         );
  OAI21_X1 U9442 ( .B1(n9529), .B2(n9415), .A(n7754), .ZN(P1_U3279) );
  INV_X1 U9443 ( .A(n7755), .ZN(n7780) );
  OAI222_X1 U9444 ( .A1(n7757), .A2(n7780), .B1(P2_U3151), .B2(n6802), .C1(
        n7756), .C2(n8888), .ZN(P2_U3270) );
  AOI21_X1 U9445 ( .B1(n7761), .B2(n7760), .A(n7784), .ZN(n7778) );
  INV_X1 U9446 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10260) );
  AOI21_X2 U9447 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n7763), .A(n7762), .ZN(
        n7791) );
  XNOR2_X1 U9448 ( .A(n7791), .B(n7792), .ZN(n7764) );
  AOI21_X1 U9449 ( .B1(n10260), .B2(n7764), .A(n7793), .ZN(n7765) );
  NOR2_X1 U9450 ( .A1(n7765), .A2(n10133), .ZN(n7776) );
  MUX2_X1 U9451 ( .A(n7761), .B(n10260), .S(n6509), .Z(n7767) );
  AND2_X1 U9452 ( .A1(n7767), .A2(n7792), .ZN(n7802) );
  INV_X1 U9453 ( .A(n7802), .ZN(n7766) );
  OAI21_X1 U9454 ( .B1(n7792), .B2(n7767), .A(n7766), .ZN(n7771) );
  AOI21_X1 U9455 ( .B1(n7771), .B2(n7770), .A(n7801), .ZN(n7774) );
  AOI22_X1 U9456 ( .A1(n10139), .A2(n7792), .B1(n10115), .B2(
        P2_ADDR_REG_11__SCAN_IN), .ZN(n7773) );
  INV_X1 U9457 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8793) );
  NOR2_X1 U9458 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8793), .ZN(n8020) );
  INV_X1 U9459 ( .A(n8020), .ZN(n7772) );
  OAI211_X1 U9460 ( .C1(n7774), .C2(n8250), .A(n7773), .B(n7772), .ZN(n7775)
         );
  NOR2_X1 U9461 ( .A1(n7776), .A2(n7775), .ZN(n7777) );
  OAI21_X1 U9462 ( .B1(n7778), .B2(n10135), .A(n7777), .ZN(P2_U3193) );
  OAI222_X1 U9463 ( .A1(n7782), .A2(P1_U3086), .B1(n7781), .B2(n7780), .C1(
        n7779), .C2(n9562), .ZN(P1_U3330) );
  NOR2_X1 U9464 ( .A1(n7792), .A2(n7783), .ZN(n7785) );
  INV_X1 U9465 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7786) );
  AOI22_X1 U9466 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n8106), .B1(n7803), .B2(
        n7786), .ZN(n7787) );
  AOI21_X1 U9467 ( .B1(n7788), .B2(n7787), .A(n8105), .ZN(n7811) );
  NOR2_X1 U9468 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7789), .ZN(n7947) );
  INV_X1 U9469 ( .A(n7947), .ZN(n7790) );
  OAI21_X1 U9470 ( .B1(n10112), .B2(n7803), .A(n7790), .ZN(n7800) );
  INV_X1 U9471 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8096) );
  MUX2_X1 U9472 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n8096), .S(n8106), .Z(n7796)
         );
  INV_X1 U9473 ( .A(n8097), .ZN(n7795) );
  AOI21_X1 U9474 ( .B1(n7797), .B2(n7796), .A(n7795), .ZN(n7798) );
  NOR2_X1 U9475 ( .A1(n7798), .A2(n10133), .ZN(n7799) );
  AOI211_X1 U9476 ( .C1(n10115), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n7800), .B(
        n7799), .ZN(n7810) );
  MUX2_X1 U9477 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8241), .Z(n7804) );
  AND2_X1 U9478 ( .A1(n7804), .A2(n7803), .ZN(n8090) );
  INV_X1 U9479 ( .A(n8090), .ZN(n7806) );
  MUX2_X1 U9480 ( .A(n7786), .B(n8096), .S(n8241), .Z(n7805) );
  NAND2_X1 U9481 ( .A1(n7805), .A2(n8106), .ZN(n8091) );
  NAND2_X1 U9482 ( .A1(n7806), .A2(n8091), .ZN(n7807) );
  XNOR2_X1 U9483 ( .A(n8092), .B(n7807), .ZN(n7808) );
  NAND2_X1 U9484 ( .A1(n7808), .A2(n10143), .ZN(n7809) );
  OAI211_X1 U9485 ( .C1(n7811), .C2(n10135), .A(n7810), .B(n7809), .ZN(
        P2_U3194) );
  INV_X1 U9486 ( .A(n7812), .ZN(n9556) );
  OAI222_X1 U9487 ( .A1(n8890), .A2(n9556), .B1(n5947), .B2(P2_U3151), .C1(
        n7813), .C2(n8888), .ZN(P2_U3266) );
  INV_X1 U9488 ( .A(n7814), .ZN(n8071) );
  NAND2_X1 U9489 ( .A1(n8071), .A2(n7815), .ZN(n7818) );
  NOR2_X1 U9490 ( .A1(n7818), .A2(n10238), .ZN(n8520) );
  AOI21_X1 U9491 ( .B1(n10238), .B2(P2_REG0_REG_30__SCAN_IN), .A(n8520), .ZN(
        n7816) );
  OAI21_X1 U9492 ( .B1(n7822), .B2(n8873), .A(n7816), .ZN(P2_U3457) );
  NOR2_X1 U9493 ( .A1(n7818), .A2(n10262), .ZN(n8465) );
  AOI21_X1 U9494 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n10262), .A(n8465), .ZN(
        n7817) );
  OAI21_X1 U9495 ( .B1(n7822), .B2(n8519), .A(n7817), .ZN(P2_U3489) );
  INV_X1 U9496 ( .A(n7818), .ZN(n7820) );
  NOR2_X1 U9497 ( .A1(n7819), .A2(n10151), .ZN(n8261) );
  AOI21_X1 U9498 ( .B1(n7820), .B2(n10167), .A(n8261), .ZN(n8257) );
  NAND2_X1 U9499 ( .A1(n8442), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7821) );
  OAI211_X1 U9500 ( .C1(n7822), .C2(n8411), .A(n8257), .B(n7821), .ZN(P2_U3203) );
  INV_X1 U9501 ( .A(n7823), .ZN(n8886) );
  OAI222_X1 U9502 ( .A1(n9562), .A2(n8735), .B1(n9565), .B2(n8886), .C1(n4459), 
        .C2(P1_U3086), .ZN(P1_U3328) );
  INV_X1 U9503 ( .A(n7824), .ZN(n7828) );
  OAI222_X1 U9504 ( .A1(n9562), .A2(n8690), .B1(n9565), .B2(n7828), .C1(n5073), 
        .C2(n4454), .ZN(P1_U3325) );
  INV_X1 U9505 ( .A(n7825), .ZN(n7827) );
  OAI222_X1 U9506 ( .A1(n8890), .A2(n7828), .B1(n7827), .B2(P2_U3151), .C1(
        n7826), .C2(n8888), .ZN(P2_U3265) );
  XNOR2_X1 U9507 ( .A(n8864), .B(n7090), .ZN(n7858) );
  XNOR2_X1 U9508 ( .A(n7901), .B(n7090), .ZN(n7904) );
  NAND2_X1 U9509 ( .A1(n7902), .A2(n7904), .ZN(n7903) );
  INV_X1 U9510 ( .A(n7831), .ZN(n7833) );
  XNOR2_X1 U9511 ( .A(n7834), .B(n7091), .ZN(n8018) );
  INV_X1 U9512 ( .A(n8018), .ZN(n7837) );
  XNOR2_X1 U9513 ( .A(n7939), .B(n7090), .ZN(n7839) );
  NAND2_X1 U9514 ( .A1(n7839), .A2(n8454), .ZN(n7941) );
  INV_X1 U9515 ( .A(n7839), .ZN(n7840) );
  NAND2_X1 U9516 ( .A1(n7840), .A2(n8080), .ZN(n7942) );
  XNOR2_X1 U9517 ( .A(n9636), .B(n7091), .ZN(n7997) );
  NAND2_X1 U9518 ( .A1(n7842), .A2(n7841), .ZN(n7843) );
  NAND2_X1 U9519 ( .A1(n7999), .A2(n7843), .ZN(n7845) );
  NAND2_X1 U9520 ( .A1(n7997), .A2(n8436), .ZN(n7844) );
  NAND2_X1 U9521 ( .A1(n7845), .A2(n7844), .ZN(n7884) );
  XNOR2_X1 U9522 ( .A(n9632), .B(n7090), .ZN(n7846) );
  XNOR2_X1 U9523 ( .A(n7846), .B(n8453), .ZN(n7886) );
  XNOR2_X1 U9524 ( .A(n8430), .B(n7090), .ZN(n7847) );
  XOR2_X1 U9525 ( .A(n8404), .B(n7847), .Z(n8060) );
  INV_X1 U9526 ( .A(n7847), .ZN(n7848) );
  INV_X1 U9527 ( .A(n7963), .ZN(n7852) );
  XOR2_X1 U9528 ( .A(n7090), .B(n8408), .Z(n7961) );
  NAND2_X1 U9529 ( .A1(n7961), .A2(n8420), .ZN(n7851) );
  XNOR2_X1 U9530 ( .A(n8511), .B(n7091), .ZN(n7969) );
  NAND2_X1 U9531 ( .A1(n7971), .A2(n7853), .ZN(n7855) );
  INV_X1 U9532 ( .A(n7969), .ZN(n7854) );
  NAND2_X1 U9533 ( .A1(n7855), .A2(n5035), .ZN(n8027) );
  XNOR2_X1 U9534 ( .A(n8034), .B(n7090), .ZN(n7856) );
  NAND2_X1 U9535 ( .A1(n7856), .A2(n8368), .ZN(n7857) );
  OAI21_X1 U9536 ( .B1(n7856), .B2(n8368), .A(n7857), .ZN(n8028) );
  INV_X1 U9537 ( .A(n7857), .ZN(n7915) );
  XNOR2_X1 U9538 ( .A(n7858), .B(n8383), .ZN(n7914) );
  OAI21_X1 U9539 ( .B1(n7858), .B2(n8356), .A(n7913), .ZN(n7989) );
  XNOR2_X1 U9540 ( .A(n8499), .B(n7091), .ZN(n7990) );
  INV_X1 U9541 ( .A(n8369), .ZN(n8078) );
  NAND2_X1 U9542 ( .A1(n7990), .A2(n8078), .ZN(n7860) );
  INV_X1 U9543 ( .A(n7990), .ZN(n7859) );
  XNOR2_X1 U9544 ( .A(n7931), .B(n7090), .ZN(n7861) );
  XNOR2_X1 U9545 ( .A(n7861), .B(n8333), .ZN(n7932) );
  XNOR2_X1 U9546 ( .A(n8542), .B(n7091), .ZN(n7980) );
  XNOR2_X1 U9547 ( .A(n8325), .B(n7091), .ZN(n7864) );
  OAI22_X1 U9548 ( .A1(n7980), .A2(n8322), .B1(n8334), .B2(n7979), .ZN(n7868)
         );
  OAI21_X1 U9549 ( .B1(n7864), .B2(n8077), .A(n8076), .ZN(n7866) );
  NOR2_X1 U9550 ( .A1(n8076), .A2(n8077), .ZN(n7865) );
  AOI22_X1 U9551 ( .A1(n7980), .A2(n7866), .B1(n7865), .B2(n7979), .ZN(n7867)
         );
  XNOR2_X1 U9552 ( .A(n8304), .B(n7090), .ZN(n7869) );
  XOR2_X1 U9553 ( .A(n8313), .B(n7869), .Z(n7955) );
  NAND2_X1 U9554 ( .A1(n7869), .A2(n8313), .ZN(n7870) );
  NAND2_X1 U9555 ( .A1(n7871), .A2(n7870), .ZN(n8049) );
  INV_X1 U9556 ( .A(n8049), .ZN(n7873) );
  XNOR2_X1 U9557 ( .A(n8299), .B(n7090), .ZN(n7874) );
  XNOR2_X1 U9558 ( .A(n7874), .B(n8303), .ZN(n8051) );
  INV_X1 U9559 ( .A(n8051), .ZN(n7872) );
  INV_X1 U9560 ( .A(n7874), .ZN(n7875) );
  NAND2_X1 U9561 ( .A1(n7875), .A2(n8075), .ZN(n7876) );
  XNOR2_X1 U9562 ( .A(n8530), .B(n7091), .ZN(n7877) );
  NOR2_X1 U9563 ( .A1(n7877), .A2(n8267), .ZN(n7922) );
  AOI21_X1 U9564 ( .B1(n8267), .B2(n7877), .A(n7922), .ZN(n7878) );
  OAI211_X1 U9565 ( .C1(n7879), .C2(n7878), .A(n7923), .B(n8058), .ZN(n7883)
         );
  AOI22_X1 U9566 ( .A1(n8075), .A2(n8062), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n7880) );
  OAI21_X1 U9567 ( .B1(n8281), .B2(n8064), .A(n7880), .ZN(n7881) );
  AOI21_X1 U9568 ( .B1(n8284), .B2(n8067), .A(n7881), .ZN(n7882) );
  OAI211_X1 U9569 ( .C1(n8530), .C2(n8070), .A(n7883), .B(n7882), .ZN(P2_U3154) );
  AOI21_X1 U9570 ( .B1(n7886), .B2(n7884), .A(n7885), .ZN(n7892) );
  NAND2_X1 U9571 ( .A1(n8067), .A2(n8439), .ZN(n7889) );
  INV_X1 U9572 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7887) );
  NOR2_X1 U9573 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7887), .ZN(n8130) );
  AOI21_X1 U9574 ( .B1(n8062), .B2(n8436), .A(n8130), .ZN(n7888) );
  OAI211_X1 U9575 ( .C1(n8404), .C2(n8064), .A(n7889), .B(n7888), .ZN(n7890)
         );
  AOI21_X1 U9576 ( .B1(n9632), .B2(n8033), .A(n7890), .ZN(n7891) );
  OAI21_X1 U9577 ( .B1(n7892), .B2(n8050), .A(n7891), .ZN(P2_U3155) );
  XNOR2_X1 U9578 ( .A(n7893), .B(n7979), .ZN(n7894) );
  NAND2_X1 U9579 ( .A1(n7894), .A2(n8077), .ZN(n7977) );
  OAI211_X1 U9580 ( .C1(n7894), .C2(n8077), .A(n7977), .B(n8058), .ZN(n7900)
         );
  INV_X1 U9581 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8673) );
  OAI22_X1 U9582 ( .A1(n8344), .A2(n8031), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8673), .ZN(n7895) );
  AOI21_X1 U9583 ( .B1(n8076), .B2(n8043), .A(n7895), .ZN(n7899) );
  NAND2_X1 U9584 ( .A1(n8325), .A2(n8033), .ZN(n7898) );
  INV_X1 U9585 ( .A(n8326), .ZN(n7896) );
  OR2_X1 U9586 ( .A1(n8003), .A2(n7896), .ZN(n7897) );
  NAND4_X1 U9587 ( .A1(n7900), .A2(n7899), .A3(n7898), .A4(n7897), .ZN(
        P2_U3156) );
  NAND2_X1 U9588 ( .A1(n7901), .A2(n10180), .ZN(n10220) );
  OAI21_X1 U9589 ( .B1(n7902), .B2(n7904), .A(n7903), .ZN(n7905) );
  NAND2_X1 U9590 ( .A1(n7905), .A2(n8058), .ZN(n7912) );
  AOI21_X1 U9591 ( .B1(n8062), .B2(n8082), .A(n7906), .ZN(n7907) );
  OAI21_X1 U9592 ( .B1(n7908), .B2(n8064), .A(n7907), .ZN(n7909) );
  AOI21_X1 U9593 ( .B1(n8067), .B2(n7910), .A(n7909), .ZN(n7911) );
  OAI211_X1 U9594 ( .C1(n7953), .C2(n10220), .A(n7912), .B(n7911), .ZN(
        P2_U3157) );
  INV_X1 U9595 ( .A(n7913), .ZN(n7917) );
  NOR3_X1 U9596 ( .A1(n8026), .A2(n7915), .A3(n7914), .ZN(n7916) );
  OAI21_X1 U9597 ( .B1(n7917), .B2(n7916), .A(n8058), .ZN(n7921) );
  NAND2_X1 U9598 ( .A1(n8043), .A2(n8078), .ZN(n7918) );
  NAND2_X1 U9599 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8246) );
  OAI211_X1 U9600 ( .C1(n8368), .C2(n8031), .A(n7918), .B(n8246), .ZN(n7919)
         );
  AOI21_X1 U9601 ( .B1(n8067), .B2(n8375), .A(n7919), .ZN(n7920) );
  OAI211_X1 U9602 ( .C1(n8864), .C2(n8070), .A(n7921), .B(n7920), .ZN(P2_U3159) );
  XOR2_X1 U9603 ( .A(n7090), .B(n8273), .Z(n7924) );
  INV_X1 U9604 ( .A(n7925), .ZN(n8272) );
  INV_X1 U9605 ( .A(n8268), .ZN(n8073) );
  INV_X1 U9606 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8659) );
  OAI22_X1 U9607 ( .A1(n8267), .A2(n8031), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8659), .ZN(n7926) );
  AOI21_X1 U9608 ( .B1(n8043), .B2(n8073), .A(n7926), .ZN(n7927) );
  OAI21_X1 U9609 ( .B1(n8272), .B2(n8003), .A(n7927), .ZN(n7928) );
  AOI21_X1 U9610 ( .B1(n8277), .B2(n8033), .A(n7928), .ZN(n7929) );
  OAI21_X1 U9611 ( .B1(n7930), .B2(n8050), .A(n7929), .ZN(P2_U3160) );
  INV_X1 U9612 ( .A(n7931), .ZN(n8554) );
  XNOR2_X1 U9613 ( .A(n7933), .B(n7932), .ZN(n7934) );
  NAND2_X1 U9614 ( .A1(n7934), .A2(n8058), .ZN(n7938) );
  NOR2_X1 U9615 ( .A1(n8031), .A2(n8369), .ZN(n7936) );
  OAI22_X1 U9616 ( .A1(n8064), .A2(n8344), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8649), .ZN(n7935) );
  AOI211_X1 U9617 ( .C1(n8067), .C2(n8350), .A(n7936), .B(n7935), .ZN(n7937)
         );
  OAI211_X1 U9618 ( .C1(n8554), .C2(n8070), .A(n7938), .B(n7937), .ZN(P2_U3163) );
  NAND2_X1 U9619 ( .A1(n7939), .A2(n10180), .ZN(n10232) );
  INV_X1 U9620 ( .A(n7942), .ZN(n7946) );
  AOI21_X1 U9621 ( .B1(n7942), .B2(n7941), .A(n7940), .ZN(n7943) );
  NOR2_X1 U9622 ( .A1(n7943), .A2(n8050), .ZN(n7944) );
  OAI21_X1 U9623 ( .B1(n7946), .B2(n7945), .A(n7944), .ZN(n7952) );
  AOI21_X1 U9624 ( .B1(n8062), .B2(n7836), .A(n7947), .ZN(n7948) );
  OAI21_X1 U9625 ( .B1(n7841), .B2(n8064), .A(n7948), .ZN(n7949) );
  AOI21_X1 U9626 ( .B1(n8067), .B2(n7950), .A(n7949), .ZN(n7951) );
  OAI211_X1 U9627 ( .C1(n7953), .C2(n10232), .A(n7952), .B(n7951), .ZN(
        P2_U3164) );
  XOR2_X1 U9628 ( .A(n7955), .B(n7954), .Z(n7960) );
  AOI22_X1 U9629 ( .A1(n8075), .A2(n8043), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n7957) );
  NAND2_X1 U9630 ( .A1(n8067), .A2(n8305), .ZN(n7956) );
  OAI211_X1 U9631 ( .C1(n8322), .C2(n8031), .A(n7957), .B(n7956), .ZN(n7958)
         );
  AOI21_X1 U9632 ( .B1(n8304), .B2(n8033), .A(n7958), .ZN(n7959) );
  OAI21_X1 U9633 ( .B1(n7960), .B2(n8050), .A(n7959), .ZN(P2_U3165) );
  XNOR2_X1 U9634 ( .A(n7961), .B(n8065), .ZN(n7962) );
  XNOR2_X1 U9635 ( .A(n7963), .B(n7962), .ZN(n7968) );
  NAND2_X1 U9636 ( .A1(n8067), .A2(n8409), .ZN(n7965) );
  AND2_X1 U9637 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8179) );
  AOI21_X1 U9638 ( .B1(n8062), .B2(n6777), .A(n8179), .ZN(n7964) );
  OAI211_X1 U9639 ( .C1(n8405), .C2(n8064), .A(n7965), .B(n7964), .ZN(n7966)
         );
  AOI21_X1 U9640 ( .B1(n8408), .B2(n8033), .A(n7966), .ZN(n7967) );
  OAI21_X1 U9641 ( .B1(n7968), .B2(n8050), .A(n7967), .ZN(P2_U3166) );
  XNOR2_X1 U9642 ( .A(n7969), .B(n8405), .ZN(n7970) );
  XNOR2_X1 U9643 ( .A(n7971), .B(n7970), .ZN(n7976) );
  NAND2_X1 U9644 ( .A1(n8067), .A2(n8394), .ZN(n7973) );
  INV_X1 U9645 ( .A(n8368), .ZN(n8392) );
  AND2_X1 U9646 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8199) );
  AOI21_X1 U9647 ( .B1(n8043), .B2(n8392), .A(n8199), .ZN(n7972) );
  OAI211_X1 U9648 ( .C1(n8065), .C2(n8031), .A(n7973), .B(n7972), .ZN(n7974)
         );
  AOI21_X1 U9649 ( .B1(n8511), .B2(n8033), .A(n7974), .ZN(n7975) );
  OAI21_X1 U9650 ( .B1(n7976), .B2(n8050), .A(n7975), .ZN(P2_U3168) );
  INV_X1 U9651 ( .A(n7893), .ZN(n7978) );
  OAI21_X1 U9652 ( .B1(n7979), .B2(n7978), .A(n7977), .ZN(n7982) );
  XNOR2_X1 U9653 ( .A(n7980), .B(n8076), .ZN(n7981) );
  XNOR2_X1 U9654 ( .A(n7982), .B(n7981), .ZN(n7988) );
  INV_X1 U9655 ( .A(n8313), .ZN(n8290) );
  AOI22_X1 U9656 ( .A1(n8290), .A2(n8043), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n7984) );
  NAND2_X1 U9657 ( .A1(n8067), .A2(n8315), .ZN(n7983) );
  OAI211_X1 U9658 ( .C1(n8334), .C2(n8031), .A(n7984), .B(n7983), .ZN(n7985)
         );
  AOI21_X1 U9659 ( .B1(n7986), .B2(n8033), .A(n7985), .ZN(n7987) );
  OAI21_X1 U9660 ( .B1(n7988), .B2(n8050), .A(n7987), .ZN(P2_U3169) );
  XNOR2_X1 U9661 ( .A(n7990), .B(n8078), .ZN(n7991) );
  XNOR2_X1 U9662 ( .A(n7989), .B(n7991), .ZN(n7996) );
  NAND2_X1 U9663 ( .A1(n8067), .A2(n8361), .ZN(n7993) );
  AOI22_X1 U9664 ( .A1(n8357), .A2(n8043), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n7992) );
  OAI211_X1 U9665 ( .C1(n8383), .C2(n8031), .A(n7993), .B(n7992), .ZN(n7994)
         );
  AOI21_X1 U9666 ( .B1(n8499), .B2(n8033), .A(n7994), .ZN(n7995) );
  OAI21_X1 U9667 ( .B1(n7996), .B2(n8050), .A(n7995), .ZN(P2_U3173) );
  XNOR2_X1 U9668 ( .A(n7997), .B(n7841), .ZN(n7998) );
  XNOR2_X1 U9669 ( .A(n7999), .B(n7998), .ZN(n8006) );
  INV_X1 U9670 ( .A(n8000), .ZN(n8455) );
  INV_X1 U9671 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8818) );
  NOR2_X1 U9672 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8818), .ZN(n8095) );
  NOR2_X1 U9673 ( .A1(n8031), .A2(n8454), .ZN(n8001) );
  AOI211_X1 U9674 ( .C1(n8043), .C2(n8421), .A(n8095), .B(n8001), .ZN(n8002)
         );
  OAI21_X1 U9675 ( .B1(n8455), .B2(n8003), .A(n8002), .ZN(n8004) );
  AOI21_X1 U9676 ( .B1(n8033), .B2(n9636), .A(n8004), .ZN(n8005) );
  OAI21_X1 U9677 ( .B1(n8006), .B2(n8050), .A(n8005), .ZN(P2_U3174) );
  XOR2_X1 U9678 ( .A(n8008), .B(n8007), .Z(n8014) );
  NAND2_X1 U9679 ( .A1(n8067), .A2(n8337), .ZN(n8010) );
  AOI22_X1 U9680 ( .A1(n8062), .A2(n8357), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8009) );
  OAI211_X1 U9681 ( .C1(n8334), .C2(n8064), .A(n8010), .B(n8009), .ZN(n8011)
         );
  AOI21_X1 U9682 ( .B1(n8012), .B2(n8033), .A(n8011), .ZN(n8013) );
  OAI21_X1 U9683 ( .B1(n8014), .B2(n8050), .A(n8013), .ZN(P2_U3175) );
  INV_X1 U9684 ( .A(n8015), .ZN(n10226) );
  AND2_X1 U9685 ( .A1(n7903), .A2(n8016), .ZN(n8019) );
  OAI211_X1 U9686 ( .C1(n8019), .C2(n8018), .A(n8058), .B(n8017), .ZN(n8025)
         );
  AOI21_X1 U9687 ( .B1(n8062), .B2(n8081), .A(n8020), .ZN(n8021) );
  OAI21_X1 U9688 ( .B1(n8454), .B2(n8064), .A(n8021), .ZN(n8022) );
  AOI21_X1 U9689 ( .B1(n8067), .B2(n8023), .A(n8022), .ZN(n8024) );
  OAI211_X1 U9690 ( .C1(n10226), .C2(n8070), .A(n8025), .B(n8024), .ZN(
        P2_U3176) );
  AOI21_X1 U9691 ( .B1(n8028), .B2(n8027), .A(n8026), .ZN(n8036) );
  NAND2_X1 U9692 ( .A1(n8067), .A2(n8386), .ZN(n8030) );
  NOR2_X1 U9693 ( .A1(n8676), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8225) );
  AOI21_X1 U9694 ( .B1(n8043), .B2(n8356), .A(n8225), .ZN(n8029) );
  OAI211_X1 U9695 ( .C1(n8405), .C2(n8031), .A(n8030), .B(n8029), .ZN(n8032)
         );
  AOI21_X1 U9696 ( .B1(n8034), .B2(n8033), .A(n8032), .ZN(n8035) );
  OAI21_X1 U9697 ( .B1(n8036), .B2(n8050), .A(n8035), .ZN(P2_U3178) );
  OAI211_X1 U9698 ( .C1(n8039), .C2(n8038), .A(n8037), .B(n8058), .ZN(n8048)
         );
  NOR2_X1 U9699 ( .A1(n8040), .A2(n10225), .ZN(n10198) );
  INV_X1 U9700 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8041) );
  NOR2_X1 U9701 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8041), .ZN(n10099) );
  AOI21_X1 U9702 ( .B1(n8042), .B2(n10198), .A(n10099), .ZN(n8047) );
  AOI22_X1 U9703 ( .A1(n8062), .A2(n8086), .B1(n8043), .B2(n8084), .ZN(n8046)
         );
  NAND2_X1 U9704 ( .A1(n8067), .A2(n8044), .ZN(n8045) );
  NAND4_X1 U9705 ( .A1(n8048), .A2(n8047), .A3(n8046), .A4(n8045), .ZN(
        P2_U3179) );
  AOI21_X1 U9706 ( .B1(n8049), .B2(n8051), .A(n8050), .ZN(n8053) );
  NAND2_X1 U9707 ( .A1(n8053), .A2(n8052), .ZN(n8057) );
  AOI22_X1 U9708 ( .A1(n8290), .A2(n8062), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8054) );
  OAI21_X1 U9709 ( .B1(n8267), .B2(n8064), .A(n8054), .ZN(n8055) );
  AOI21_X1 U9710 ( .B1(n8292), .B2(n8067), .A(n8055), .ZN(n8056) );
  OAI211_X1 U9711 ( .C1(n8534), .C2(n8070), .A(n8057), .B(n8056), .ZN(P2_U3180) );
  OAI211_X1 U9712 ( .C1(n8061), .C2(n8060), .A(n8059), .B(n8058), .ZN(n8069)
         );
  AND2_X1 U9713 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8144) );
  AOI21_X1 U9714 ( .B1(n8062), .B2(n8421), .A(n8144), .ZN(n8063) );
  OAI21_X1 U9715 ( .B1(n8065), .B2(n8064), .A(n8063), .ZN(n8066) );
  AOI21_X1 U9716 ( .B1(n8067), .B2(n8425), .A(n8066), .ZN(n8068) );
  OAI211_X1 U9717 ( .C1(n9623), .C2(n8070), .A(n8069), .B(n8068), .ZN(P2_U3181) );
  MUX2_X1 U9718 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8071), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9719 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8072), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9720 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8073), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U9721 ( .A(n8074), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8224), .Z(
        P2_U3519) );
  INV_X1 U9722 ( .A(n8267), .ZN(n8291) );
  MUX2_X1 U9723 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8291), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9724 ( .A(n8075), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8224), .Z(
        P2_U3517) );
  MUX2_X1 U9725 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8290), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9726 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8076), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9727 ( .A(n8077), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8224), .Z(
        P2_U3514) );
  MUX2_X1 U9728 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8357), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9729 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8078), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9730 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8356), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9731 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8392), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9732 ( .A(n8079), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8224), .Z(
        P2_U3508) );
  MUX2_X1 U9733 ( .A(n8420), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8224), .Z(
        P2_U3507) );
  MUX2_X1 U9734 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n6777), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9735 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8421), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U9736 ( .A(n8436), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8224), .Z(
        P2_U3504) );
  MUX2_X1 U9737 ( .A(n8080), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8224), .Z(
        P2_U3503) );
  MUX2_X1 U9738 ( .A(n7836), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8224), .Z(
        P2_U3502) );
  MUX2_X1 U9739 ( .A(n8081), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8224), .Z(
        P2_U3501) );
  MUX2_X1 U9740 ( .A(n8082), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8224), .Z(
        P2_U3500) );
  MUX2_X1 U9741 ( .A(n8083), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8224), .Z(
        P2_U3499) );
  MUX2_X1 U9742 ( .A(n8084), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8224), .Z(
        P2_U3498) );
  MUX2_X1 U9743 ( .A(n8085), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8224), .Z(
        P2_U3497) );
  MUX2_X1 U9744 ( .A(n8086), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8224), .Z(
        P2_U3496) );
  MUX2_X1 U9745 ( .A(n8087), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8224), .Z(
        P2_U3495) );
  MUX2_X1 U9746 ( .A(n8088), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8224), .Z(
        P2_U3494) );
  MUX2_X1 U9747 ( .A(n7155), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8224), .Z(
        P2_U3493) );
  MUX2_X1 U9748 ( .A(n8089), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8224), .Z(
        P2_U3492) );
  MUX2_X1 U9749 ( .A(n6010), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8224), .Z(
        P2_U3491) );
  AOI21_X1 U9750 ( .B1(n8092), .B2(n8091), .A(n8090), .ZN(n8094) );
  MUX2_X1 U9751 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8241), .Z(n8119) );
  XNOR2_X1 U9752 ( .A(n8119), .B(n8099), .ZN(n8093) );
  NAND2_X1 U9753 ( .A1(n8094), .A2(n8093), .ZN(n8120) );
  OAI21_X1 U9754 ( .B1(n8094), .B2(n8093), .A(n8120), .ZN(n8113) );
  NAND2_X1 U9755 ( .A1(n10115), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n8104) );
  AOI21_X1 U9756 ( .B1(n10139), .B2(n8099), .A(n8095), .ZN(n8103) );
  OR2_X1 U9757 ( .A1(n8106), .A2(n8096), .ZN(n8098) );
  OAI21_X1 U9758 ( .B1(n8100), .B2(P2_REG1_REG_13__SCAN_IN), .A(n8127), .ZN(
        n8101) );
  NAND2_X1 U9759 ( .A1(n10121), .A2(n8101), .ZN(n8102) );
  NAND3_X1 U9760 ( .A1(n8104), .A2(n8103), .A3(n8102), .ZN(n8112) );
  INV_X1 U9761 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8464) );
  AOI21_X1 U9762 ( .B1(n8109), .B2(n8464), .A(n8116), .ZN(n8110) );
  NOR2_X1 U9763 ( .A1(n8110), .A2(n10135), .ZN(n8111) );
  AOI211_X1 U9764 ( .C1(n10143), .C2(n8113), .A(n8112), .B(n8111), .ZN(n8114)
         );
  INV_X1 U9765 ( .A(n8114), .ZN(P2_U3195) );
  INV_X1 U9766 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8446) );
  AOI22_X1 U9767 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8154), .B1(n8138), .B2(
        n8446), .ZN(n8117) );
  AOI21_X1 U9768 ( .B1(n8118), .B2(n8117), .A(n8155), .ZN(n8137) );
  MUX2_X1 U9769 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n6509), .Z(n8139) );
  XNOR2_X1 U9770 ( .A(n8139), .B(n8154), .ZN(n8123) );
  OR2_X1 U9771 ( .A1(n8119), .A2(n8125), .ZN(n8121) );
  NAND2_X1 U9772 ( .A1(n8121), .A2(n8120), .ZN(n8122) );
  NAND2_X1 U9773 ( .A1(n8123), .A2(n8122), .ZN(n8140) );
  OAI21_X1 U9774 ( .B1(n8123), .B2(n8122), .A(n8140), .ZN(n8135) );
  INV_X1 U9775 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8145) );
  MUX2_X1 U9776 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8145), .S(n8154), .Z(n8129)
         );
  AOI21_X1 U9777 ( .B1(n4531), .B2(n8129), .A(n8128), .ZN(n8133) );
  NAND2_X1 U9778 ( .A1(n10115), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n8132) );
  AOI21_X1 U9779 ( .B1(n10139), .B2(n8154), .A(n8130), .ZN(n8131) );
  OAI211_X1 U9780 ( .C1(n10133), .C2(n8133), .A(n8132), .B(n8131), .ZN(n8134)
         );
  AOI21_X1 U9781 ( .B1(n10143), .B2(n8135), .A(n8134), .ZN(n8136) );
  OAI21_X1 U9782 ( .B1(n8137), .B2(n10135), .A(n8136), .ZN(P2_U3196) );
  MUX2_X1 U9783 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8241), .Z(n8168) );
  XNOR2_X1 U9784 ( .A(n8168), .B(n8148), .ZN(n8143) );
  OR2_X1 U9785 ( .A1(n8139), .A2(n8138), .ZN(n8141) );
  NAND2_X1 U9786 ( .A1(n8141), .A2(n8140), .ZN(n8142) );
  NAND2_X1 U9787 ( .A1(n8143), .A2(n8142), .ZN(n8169) );
  OAI21_X1 U9788 ( .B1(n8143), .B2(n8142), .A(n8169), .ZN(n8161) );
  NAND2_X1 U9789 ( .A1(n10115), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n8153) );
  AOI21_X1 U9790 ( .B1(n10139), .B2(n8148), .A(n8144), .ZN(n8152) );
  OR2_X1 U9791 ( .A1(n8154), .A2(n8145), .ZN(n8147) );
  NAND2_X1 U9792 ( .A1(n8147), .A2(n8146), .ZN(n8173) );
  XNOR2_X1 U9793 ( .A(n8173), .B(n8148), .ZN(n8149) );
  NAND2_X1 U9794 ( .A1(n8149), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8176) );
  OAI21_X1 U9795 ( .B1(n8149), .B2(P2_REG1_REG_15__SCAN_IN), .A(n8176), .ZN(
        n8150) );
  NAND2_X1 U9796 ( .A1(n10121), .A2(n8150), .ZN(n8151) );
  NAND3_X1 U9797 ( .A1(n8153), .A2(n8152), .A3(n8151), .ZN(n8160) );
  INV_X1 U9798 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8427) );
  AOI21_X1 U9799 ( .B1(n8157), .B2(n8427), .A(n8164), .ZN(n8158) );
  NOR2_X1 U9800 ( .A1(n8158), .A2(n10135), .ZN(n8159) );
  AOI211_X1 U9801 ( .C1(n10143), .C2(n8161), .A(n8160), .B(n8159), .ZN(n8162)
         );
  INV_X1 U9802 ( .A(n8162), .ZN(P2_U3197) );
  INV_X1 U9803 ( .A(n8163), .ZN(n8165) );
  INV_X1 U9804 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8843) );
  AOI22_X1 U9805 ( .A1(n8190), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8843), .B2(
        n8196), .ZN(n8166) );
  AOI21_X1 U9806 ( .B1(n8167), .B2(n8166), .A(n8187), .ZN(n8186) );
  INV_X1 U9807 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8517) );
  MUX2_X1 U9808 ( .A(n8843), .B(n8517), .S(n8241), .Z(n8189) );
  XNOR2_X1 U9809 ( .A(n8189), .B(n8196), .ZN(n8172) );
  OR2_X1 U9810 ( .A1(n8168), .A2(n8174), .ZN(n8170) );
  NAND2_X1 U9811 ( .A1(n8170), .A2(n8169), .ZN(n8171) );
  NAND2_X1 U9812 ( .A1(n8172), .A2(n8171), .ZN(n8191) );
  OAI21_X1 U9813 ( .B1(n8172), .B2(n8171), .A(n8191), .ZN(n8184) );
  NAND2_X1 U9814 ( .A1(n8174), .A2(n8173), .ZN(n8175) );
  MUX2_X1 U9815 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8517), .S(n8190), .Z(n8177)
         );
  AOI21_X1 U9816 ( .B1(n8178), .B2(n8177), .A(n8195), .ZN(n8182) );
  NAND2_X1 U9817 ( .A1(n10115), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n8181) );
  AOI21_X1 U9818 ( .B1(n10139), .B2(n8190), .A(n8179), .ZN(n8180) );
  OAI211_X1 U9819 ( .C1(n10133), .C2(n8182), .A(n8181), .B(n8180), .ZN(n8183)
         );
  AOI21_X1 U9820 ( .B1(n10143), .B2(n8184), .A(n8183), .ZN(n8185) );
  OAI21_X1 U9821 ( .B1(n8186), .B2(n10135), .A(n8185), .ZN(P2_U3198) );
  INV_X1 U9822 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8836) );
  AOI21_X1 U9823 ( .B1(n8836), .B2(n8188), .A(n8208), .ZN(n8206) );
  INV_X1 U9824 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8197) );
  MUX2_X1 U9825 ( .A(n8836), .B(n8197), .S(n6509), .Z(n8220) );
  XOR2_X1 U9826 ( .A(n8219), .B(n8220), .Z(n8194) );
  NAND2_X1 U9827 ( .A1(n8190), .A2(n8189), .ZN(n8192) );
  NAND2_X1 U9828 ( .A1(n8192), .A2(n8191), .ZN(n8193) );
  NAND2_X1 U9829 ( .A1(n8194), .A2(n8193), .ZN(n8217) );
  OAI21_X1 U9830 ( .B1(n8194), .B2(n8193), .A(n8217), .ZN(n8204) );
  AOI21_X1 U9831 ( .B1(n8198), .B2(n8197), .A(n8212), .ZN(n8202) );
  AOI21_X1 U9832 ( .B1(n10139), .B2(n8219), .A(n8199), .ZN(n8201) );
  NAND2_X1 U9833 ( .A1(n10115), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n8200) );
  OAI211_X1 U9834 ( .C1(n10133), .C2(n8202), .A(n8201), .B(n8200), .ZN(n8203)
         );
  AOI21_X1 U9835 ( .B1(n10143), .B2(n8204), .A(n8203), .ZN(n8205) );
  OAI21_X1 U9836 ( .B1(n8206), .B2(n10135), .A(n8205), .ZN(P2_U3199) );
  INV_X1 U9837 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8715) );
  AOI22_X1 U9838 ( .A1(n8239), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8715), .B2(
        n8235), .ZN(n8209) );
  AOI21_X1 U9839 ( .B1(n8210), .B2(n8209), .A(n8232), .ZN(n8231) );
  NOR2_X1 U9840 ( .A1(n8219), .A2(n8211), .ZN(n8213) );
  INV_X1 U9841 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8509) );
  AOI22_X1 U9842 ( .A1(n8239), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n8509), .B2(
        n8235), .ZN(n8214) );
  AOI21_X1 U9843 ( .B1(n8215), .B2(n8214), .A(n8234), .ZN(n8216) );
  INV_X1 U9844 ( .A(n8216), .ZN(n8229) );
  INV_X1 U9845 ( .A(n8217), .ZN(n8218) );
  MUX2_X1 U9846 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8241), .Z(n8221) );
  NOR2_X1 U9847 ( .A1(n8222), .A2(n8221), .ZN(n8237) );
  INV_X1 U9848 ( .A(n8237), .ZN(n8223) );
  NAND2_X1 U9849 ( .A1(n8222), .A2(n8221), .ZN(n8238) );
  NAND2_X1 U9850 ( .A1(n8223), .A2(n8238), .ZN(n8227) );
  OAI21_X1 U9851 ( .B1(n8224), .B2(n8227), .A(n10112), .ZN(n8226) );
  AOI21_X1 U9852 ( .B1(n8229), .B2(n10121), .A(n8228), .ZN(n8230) );
  OAI21_X1 U9853 ( .B1(n8231), .B2(n10135), .A(n8230), .ZN(P2_U3200) );
  INV_X1 U9854 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8233) );
  MUX2_X1 U9855 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8233), .S(n8247), .Z(n8243)
         );
  AOI21_X1 U9856 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n8235), .A(n8234), .ZN(
        n8236) );
  XNOR2_X1 U9857 ( .A(n8247), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8240) );
  XNOR2_X1 U9858 ( .A(n8236), .B(n8240), .ZN(n8253) );
  AOI21_X1 U9859 ( .B1(n8239), .B2(n8238), .A(n8237), .ZN(n8245) );
  INV_X1 U9860 ( .A(n8240), .ZN(n8242) );
  MUX2_X1 U9861 ( .A(n8243), .B(n8242), .S(n8241), .Z(n8244) );
  XNOR2_X1 U9862 ( .A(n8245), .B(n8244), .ZN(n8251) );
  OAI21_X1 U9863 ( .B1(n10112), .B2(n8247), .A(n8246), .ZN(n8248) );
  AOI21_X1 U9864 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(n10115), .A(n8248), .ZN(
        n8249) );
  OAI21_X1 U9865 ( .B1(n8251), .B2(n8250), .A(n8249), .ZN(n8252) );
  AOI21_X1 U9866 ( .B1(n8253), .B2(n10121), .A(n8252), .ZN(n8254) );
  OAI21_X1 U9867 ( .B1(n8255), .B2(n10135), .A(n8254), .ZN(P2_U3201) );
  NAND2_X1 U9868 ( .A1(n8442), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8256) );
  OAI211_X1 U9869 ( .C1(n8522), .C2(n8411), .A(n8257), .B(n8256), .ZN(P2_U3202) );
  NAND2_X1 U9870 ( .A1(n8258), .A2(n8457), .ZN(n8263) );
  NOR2_X1 U9871 ( .A1(n8259), .A2(n8411), .ZN(n8260) );
  AOI211_X1 U9872 ( .C1(n8442), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8261), .B(
        n8260), .ZN(n8262) );
  OAI211_X1 U9873 ( .C1(n8265), .C2(n8264), .A(n8263), .B(n8262), .ZN(P2_U3204) );
  XNOR2_X1 U9874 ( .A(n8266), .B(n8273), .ZN(n8270) );
  OAI22_X1 U9875 ( .A1(n8268), .A2(n10158), .B1(n8267), .B2(n10157), .ZN(n8269) );
  OAI22_X1 U9876 ( .A1(n8272), .A2(n10151), .B1(n10167), .B2(n8271), .ZN(n8276) );
  XNOR2_X1 U9877 ( .A(n8274), .B(n8273), .ZN(n8468) );
  NOR2_X1 U9878 ( .A1(n8468), .A2(n8447), .ZN(n8275) );
  AOI211_X1 U9879 ( .C1(n8429), .C2(n8277), .A(n8276), .B(n8275), .ZN(n8278)
         );
  OAI21_X1 U9880 ( .B1(n8467), .B2(n8442), .A(n8278), .ZN(P2_U3205) );
  XNOR2_X1 U9881 ( .A(n8279), .B(n8282), .ZN(n8280) );
  OAI222_X1 U9882 ( .A1(n10158), .A2(n8281), .B1(n10157), .B2(n8303), .C1(
        n8280), .C2(n8451), .ZN(n8473) );
  AND2_X1 U9883 ( .A1(n8283), .A2(n8282), .ZN(n8471) );
  NOR3_X1 U9884 ( .A1(n4483), .A2(n8471), .A3(n8447), .ZN(n8287) );
  AOI22_X1 U9885 ( .A1(n8284), .A2(n8440), .B1(n8442), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8285) );
  OAI21_X1 U9886 ( .B1(n8530), .B2(n8411), .A(n8285), .ZN(n8286) );
  AOI211_X1 U9887 ( .C1(n8473), .C2(n10167), .A(n8287), .B(n8286), .ZN(n8288)
         );
  INV_X1 U9888 ( .A(n8288), .ZN(P2_U3206) );
  INV_X1 U9889 ( .A(n8292), .ZN(n8294) );
  OAI22_X1 U9890 ( .A1(n8294), .A2(n10151), .B1(n10167), .B2(n8293), .ZN(n8298) );
  XOR2_X1 U9891 ( .A(n8296), .B(n8295), .Z(n8477) );
  NOR2_X1 U9892 ( .A1(n8477), .A2(n8447), .ZN(n8297) );
  AOI211_X1 U9893 ( .C1(n8429), .C2(n8299), .A(n8298), .B(n8297), .ZN(n8300)
         );
  OAI21_X1 U9894 ( .B1(n8476), .B2(n8442), .A(n8300), .ZN(P2_U3207) );
  INV_X1 U9895 ( .A(n10153), .ZN(n8441) );
  XNOR2_X1 U9896 ( .A(n8301), .B(n8306), .ZN(n8302) );
  OAI222_X1 U9897 ( .A1(n10157), .A2(n8322), .B1(n10158), .B2(n8303), .C1(
        n8451), .C2(n8302), .ZN(n8480) );
  AOI21_X1 U9898 ( .B1(n8441), .B2(n8304), .A(n8480), .ZN(n8310) );
  AOI22_X1 U9899 ( .A1(n8305), .A2(n8440), .B1(n8442), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8309) );
  XNOR2_X1 U9900 ( .A(n8307), .B(n8306), .ZN(n8481) );
  NAND2_X1 U9901 ( .A1(n8481), .A2(n8461), .ZN(n8308) );
  OAI211_X1 U9902 ( .C1(n8310), .C2(n8442), .A(n8309), .B(n8308), .ZN(P2_U3208) );
  NOR2_X1 U9903 ( .A1(n8542), .A2(n10153), .ZN(n8314) );
  XNOR2_X1 U9904 ( .A(n8311), .B(n8316), .ZN(n8312) );
  OAI222_X1 U9905 ( .A1(n10157), .A2(n8334), .B1(n10158), .B2(n8313), .C1(
        n8312), .C2(n8451), .ZN(n8484) );
  AOI211_X1 U9906 ( .C1(n8440), .C2(n8315), .A(n8314), .B(n8484), .ZN(n8319)
         );
  XNOR2_X1 U9907 ( .A(n8317), .B(n8316), .ZN(n8485) );
  AOI22_X1 U9908 ( .A1(n8485), .A2(n8461), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n8442), .ZN(n8318) );
  OAI21_X1 U9909 ( .B1(n8319), .B2(n8442), .A(n8318), .ZN(P2_U3209) );
  XNOR2_X1 U9910 ( .A(n8320), .B(n8323), .ZN(n8321) );
  OAI222_X1 U9911 ( .A1(n10158), .A2(n8322), .B1(n10157), .B2(n8344), .C1(
        n8451), .C2(n8321), .ZN(n8487) );
  INV_X1 U9912 ( .A(n8487), .ZN(n8330) );
  XNOR2_X1 U9913 ( .A(n8324), .B(n8323), .ZN(n8488) );
  INV_X1 U9914 ( .A(n8325), .ZN(n8546) );
  AOI22_X1 U9915 ( .A1(n8442), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8440), .B2(
        n8326), .ZN(n8327) );
  OAI21_X1 U9916 ( .B1(n8546), .B2(n8411), .A(n8327), .ZN(n8328) );
  AOI21_X1 U9917 ( .B1(n8488), .B2(n8461), .A(n8328), .ZN(n8329) );
  OAI21_X1 U9918 ( .B1(n8330), .B2(n8442), .A(n8329), .ZN(P2_U3210) );
  XNOR2_X1 U9919 ( .A(n8331), .B(n4982), .ZN(n8332) );
  OAI222_X1 U9920 ( .A1(n10158), .A2(n8334), .B1(n10157), .B2(n8333), .C1(
        n8451), .C2(n8332), .ZN(n8491) );
  INV_X1 U9921 ( .A(n8491), .ZN(n8341) );
  XNOR2_X1 U9922 ( .A(n8336), .B(n8335), .ZN(n8492) );
  AOI22_X1 U9923 ( .A1(n8442), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8440), .B2(
        n8337), .ZN(n8338) );
  OAI21_X1 U9924 ( .B1(n8550), .B2(n8411), .A(n8338), .ZN(n8339) );
  AOI21_X1 U9925 ( .B1(n8492), .B2(n8461), .A(n8339), .ZN(n8340) );
  OAI21_X1 U9926 ( .B1(n8341), .B2(n8442), .A(n8340), .ZN(P2_U3211) );
  XOR2_X1 U9927 ( .A(n8349), .B(n8342), .Z(n8343) );
  OAI22_X1 U9928 ( .A1(n8343), .A2(n8451), .B1(n8369), .B2(n10157), .ZN(n8495)
         );
  NOR2_X1 U9929 ( .A1(n8344), .A2(n10158), .ZN(n8496) );
  OAI21_X1 U9930 ( .B1(n8495), .B2(n8496), .A(n10167), .ZN(n8354) );
  INV_X1 U9931 ( .A(n8345), .ZN(n8346) );
  NOR2_X1 U9932 ( .A1(n8347), .A2(n8346), .ZN(n8348) );
  XOR2_X1 U9933 ( .A(n8349), .B(n8348), .Z(n8497) );
  AOI22_X1 U9934 ( .A1(n8442), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8440), .B2(
        n8350), .ZN(n8351) );
  OAI21_X1 U9935 ( .B1(n8554), .B2(n8411), .A(n8351), .ZN(n8352) );
  AOI21_X1 U9936 ( .B1(n8497), .B2(n8461), .A(n8352), .ZN(n8353) );
  NAND2_X1 U9937 ( .A1(n8354), .A2(n8353), .ZN(P2_U3212) );
  XNOR2_X1 U9938 ( .A(n8355), .B(n8359), .ZN(n8358) );
  AOI222_X1 U9939 ( .A1(n6797), .A2(n8358), .B1(n8357), .B2(n8437), .C1(n8356), 
        .C2(n8435), .ZN(n8502) );
  XNOR2_X1 U9940 ( .A(n8360), .B(n8359), .ZN(n8500) );
  AOI22_X1 U9941 ( .A1(n8442), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8440), .B2(
        n8361), .ZN(n8362) );
  OAI21_X1 U9942 ( .B1(n8363), .B2(n8411), .A(n8362), .ZN(n8364) );
  AOI21_X1 U9943 ( .B1(n8500), .B2(n8461), .A(n8364), .ZN(n8365) );
  OAI21_X1 U9944 ( .B1(n8502), .B2(n8442), .A(n8365), .ZN(P2_U3213) );
  XNOR2_X1 U9945 ( .A(n8366), .B(n8373), .ZN(n8367) );
  OAI222_X1 U9946 ( .A1(n10158), .A2(n8369), .B1(n10157), .B2(n8368), .C1(
        n8367), .C2(n8451), .ZN(n8503) );
  INV_X1 U9947 ( .A(n8503), .ZN(n8379) );
  INV_X1 U9948 ( .A(n8370), .ZN(n8371) );
  NOR2_X1 U9949 ( .A1(n8372), .A2(n8371), .ZN(n8374) );
  XNOR2_X1 U9950 ( .A(n8374), .B(n8373), .ZN(n8504) );
  AOI22_X1 U9951 ( .A1(n8442), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8440), .B2(
        n8375), .ZN(n8376) );
  OAI21_X1 U9952 ( .B1(n8864), .B2(n8411), .A(n8376), .ZN(n8377) );
  AOI21_X1 U9953 ( .B1(n8504), .B2(n8461), .A(n8377), .ZN(n8378) );
  OAI21_X1 U9954 ( .B1(n8379), .B2(n8442), .A(n8378), .ZN(P2_U3214) );
  AOI21_X1 U9955 ( .B1(n8385), .B2(n8381), .A(n8380), .ZN(n8382) );
  OAI222_X1 U9956 ( .A1(n10157), .A2(n8405), .B1(n10158), .B2(n8383), .C1(
        n8451), .C2(n8382), .ZN(n8507) );
  INV_X1 U9957 ( .A(n8507), .ZN(n8390) );
  XOR2_X1 U9958 ( .A(n8385), .B(n8384), .Z(n8508) );
  AOI22_X1 U9959 ( .A1(n8442), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8386), .B2(
        n8440), .ZN(n8387) );
  OAI21_X1 U9960 ( .B1(n8868), .B2(n8411), .A(n8387), .ZN(n8388) );
  AOI21_X1 U9961 ( .B1(n8508), .B2(n8461), .A(n8388), .ZN(n8389) );
  OAI21_X1 U9962 ( .B1(n8390), .B2(n8442), .A(n8389), .ZN(P2_U3215) );
  XNOR2_X1 U9963 ( .A(n8391), .B(n5012), .ZN(n8393) );
  AOI222_X1 U9964 ( .A1(n6797), .A2(n8393), .B1(n8392), .B2(n8437), .C1(n8420), 
        .C2(n8435), .ZN(n8513) );
  INV_X1 U9965 ( .A(n8394), .ZN(n8395) );
  OAI22_X1 U9966 ( .A1(n10167), .A2(n8836), .B1(n8395), .B2(n10151), .ZN(n8399) );
  AOI21_X1 U9967 ( .B1(n5012), .B2(n8397), .A(n8396), .ZN(n8514) );
  NOR2_X1 U9968 ( .A1(n8514), .A2(n8447), .ZN(n8398) );
  AOI211_X1 U9969 ( .C1(n8429), .C2(n8511), .A(n8399), .B(n8398), .ZN(n8400)
         );
  OAI21_X1 U9970 ( .B1(n8513), .B2(n8442), .A(n8400), .ZN(P2_U3216) );
  XNOR2_X1 U9971 ( .A(n8402), .B(n8401), .ZN(n8403) );
  OAI222_X1 U9972 ( .A1(n10158), .A2(n8405), .B1(n10157), .B2(n8404), .C1(
        n8451), .C2(n8403), .ZN(n8515) );
  INV_X1 U9973 ( .A(n8515), .ZN(n8414) );
  XNOR2_X1 U9974 ( .A(n8407), .B(n8406), .ZN(n8516) );
  INV_X1 U9975 ( .A(n8408), .ZN(n8874) );
  AOI22_X1 U9976 ( .A1(n8442), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8440), .B2(
        n8409), .ZN(n8410) );
  OAI21_X1 U9977 ( .B1(n8874), .B2(n8411), .A(n8410), .ZN(n8412) );
  AOI21_X1 U9978 ( .B1(n8516), .B2(n8461), .A(n8412), .ZN(n8413) );
  OAI21_X1 U9979 ( .B1(n8414), .B2(n8442), .A(n8413), .ZN(P2_U3217) );
  XNOR2_X1 U9980 ( .A(n8416), .B(n8415), .ZN(n9624) );
  NAND2_X1 U9981 ( .A1(n8417), .A2(n6797), .ZN(n8424) );
  AOI21_X1 U9982 ( .B1(n8433), .B2(n8419), .A(n8418), .ZN(n8423) );
  AOI22_X1 U9983 ( .A1(n8435), .A2(n8421), .B1(n8420), .B2(n8437), .ZN(n8422)
         );
  OAI21_X1 U9984 ( .B1(n8424), .B2(n8423), .A(n8422), .ZN(n9626) );
  NAND2_X1 U9985 ( .A1(n9626), .A2(n8457), .ZN(n8432) );
  INV_X1 U9986 ( .A(n8425), .ZN(n8426) );
  OAI22_X1 U9987 ( .A1(n10167), .A2(n8427), .B1(n8426), .B2(n10151), .ZN(n8428) );
  AOI21_X1 U9988 ( .B1(n8430), .B2(n8429), .A(n8428), .ZN(n8431) );
  OAI211_X1 U9989 ( .C1(n9624), .C2(n8447), .A(n8432), .B(n8431), .ZN(P2_U3218) );
  OAI21_X1 U9990 ( .B1(n8434), .B2(n8444), .A(n8433), .ZN(n8438) );
  AOI222_X1 U9991 ( .A1(n6797), .A2(n8438), .B1(n6777), .B2(n8437), .C1(n8436), 
        .C2(n8435), .ZN(n9629) );
  AOI22_X1 U9992 ( .A1(n9632), .A2(n8441), .B1(n8440), .B2(n8439), .ZN(n8443)
         );
  AOI21_X1 U9993 ( .B1(n9629), .B2(n8443), .A(n8442), .ZN(n8449) );
  XNOR2_X1 U9994 ( .A(n8445), .B(n8444), .ZN(n9628) );
  OAI22_X1 U9995 ( .A1(n9628), .A2(n8447), .B1(n8446), .B2(n10167), .ZN(n8448)
         );
  OR2_X1 U9996 ( .A1(n8449), .A2(n8448), .ZN(P2_U3219) );
  XNOR2_X1 U9997 ( .A(n8450), .B(n8459), .ZN(n8452) );
  OAI222_X1 U9998 ( .A1(n10157), .A2(n8454), .B1(n10158), .B2(n8453), .C1(
        n8452), .C2(n8451), .ZN(n9634) );
  INV_X1 U9999 ( .A(n9636), .ZN(n8456) );
  OAI22_X1 U10000 ( .A1(n8456), .A2(n10153), .B1(n8455), .B2(n10151), .ZN(
        n8458) );
  OAI21_X1 U10001 ( .B1(n9634), .B2(n8458), .A(n8457), .ZN(n8463) );
  XNOR2_X1 U10002 ( .A(n8460), .B(n8459), .ZN(n9633) );
  NAND2_X1 U10003 ( .A1(n9633), .A2(n8461), .ZN(n8462) );
  OAI211_X1 U10004 ( .C1(n8464), .C2(n10167), .A(n8463), .B(n8462), .ZN(
        P2_U3220) );
  AOI21_X1 U10005 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n10262), .A(n8465), .ZN(
        n8466) );
  OAI21_X1 U10006 ( .B1(n8522), .B2(n8519), .A(n8466), .ZN(P2_U3490) );
  OAI21_X1 U10007 ( .B1(n10227), .B2(n8468), .A(n8467), .ZN(n8523) );
  INV_X1 U10008 ( .A(n8469), .ZN(n8470) );
  OAI21_X1 U10009 ( .B1(n8526), .B2(n8519), .A(n8470), .ZN(P2_U3487) );
  INV_X1 U10010 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8474) );
  NOR3_X1 U10011 ( .A1(n4483), .A2(n8471), .A3(n10227), .ZN(n8472) );
  NOR2_X1 U10012 ( .A1(n8473), .A2(n8472), .ZN(n8527) );
  MUX2_X1 U10013 ( .A(n8474), .B(n8527), .S(n10264), .Z(n8475) );
  OAI21_X1 U10014 ( .B1(n8530), .B2(n8519), .A(n8475), .ZN(P2_U3486) );
  OAI21_X1 U10015 ( .B1(n10227), .B2(n8477), .A(n8476), .ZN(n8531) );
  MUX2_X1 U10016 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8531), .S(n10264), .Z(
        n8478) );
  INV_X1 U10017 ( .A(n8478), .ZN(n8479) );
  OAI21_X1 U10018 ( .B1(n8534), .B2(n8519), .A(n8479), .ZN(P2_U3485) );
  INV_X1 U10019 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8482) );
  AOI21_X1 U10020 ( .B1(n10234), .B2(n8481), .A(n8480), .ZN(n8535) );
  MUX2_X1 U10021 ( .A(n8482), .B(n8535), .S(n10264), .Z(n8483) );
  OAI21_X1 U10022 ( .B1(n8538), .B2(n8519), .A(n8483), .ZN(P2_U3484) );
  AOI21_X1 U10023 ( .B1(n8485), .B2(n10234), .A(n8484), .ZN(n8539) );
  MUX2_X1 U10024 ( .A(n8661), .B(n8539), .S(n10264), .Z(n8486) );
  OAI21_X1 U10025 ( .B1(n8542), .B2(n8519), .A(n8486), .ZN(P2_U3483) );
  INV_X1 U10026 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8489) );
  AOI21_X1 U10027 ( .B1(n10234), .B2(n8488), .A(n8487), .ZN(n8543) );
  MUX2_X1 U10028 ( .A(n8489), .B(n8543), .S(n10264), .Z(n8490) );
  OAI21_X1 U10029 ( .B1(n8546), .B2(n8519), .A(n8490), .ZN(P2_U3482) );
  INV_X1 U10030 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8493) );
  AOI21_X1 U10031 ( .B1(n10234), .B2(n8492), .A(n8491), .ZN(n8547) );
  MUX2_X1 U10032 ( .A(n8493), .B(n8547), .S(n10264), .Z(n8494) );
  OAI21_X1 U10033 ( .B1(n8550), .B2(n8519), .A(n8494), .ZN(P2_U3481) );
  INV_X1 U10034 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8624) );
  AOI211_X1 U10035 ( .C1(n8497), .C2(n10234), .A(n8496), .B(n8495), .ZN(n8551)
         );
  MUX2_X1 U10036 ( .A(n8624), .B(n8551), .S(n10264), .Z(n8498) );
  OAI21_X1 U10037 ( .B1(n8554), .B2(n8519), .A(n8498), .ZN(P2_U3480) );
  AOI22_X1 U10038 ( .A1(n8500), .A2(n10234), .B1(n10180), .B2(n8499), .ZN(
        n8501) );
  NAND2_X1 U10039 ( .A1(n8502), .A2(n8501), .ZN(n8555) );
  MUX2_X1 U10040 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8555), .S(n10264), .Z(
        P2_U3479) );
  INV_X1 U10041 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8505) );
  AOI21_X1 U10042 ( .B1(n10234), .B2(n8504), .A(n8503), .ZN(n8861) );
  MUX2_X1 U10043 ( .A(n8505), .B(n8861), .S(n10264), .Z(n8506) );
  OAI21_X1 U10044 ( .B1(n8864), .B2(n8519), .A(n8506), .ZN(P2_U3478) );
  AOI21_X1 U10045 ( .B1(n8508), .B2(n10234), .A(n8507), .ZN(n8865) );
  MUX2_X1 U10046 ( .A(n8509), .B(n8865), .S(n10264), .Z(n8510) );
  OAI21_X1 U10047 ( .B1(n8868), .B2(n8519), .A(n8510), .ZN(P2_U3477) );
  NAND2_X1 U10048 ( .A1(n8511), .A2(n10180), .ZN(n8512) );
  OAI211_X1 U10049 ( .C1(n10227), .C2(n8514), .A(n8513), .B(n8512), .ZN(n8869)
         );
  MUX2_X1 U10050 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8869), .S(n10264), .Z(
        P2_U3476) );
  AOI21_X1 U10051 ( .B1(n8516), .B2(n10234), .A(n8515), .ZN(n8870) );
  MUX2_X1 U10052 ( .A(n8517), .B(n8870), .S(n10264), .Z(n8518) );
  OAI21_X1 U10053 ( .B1(n8874), .B2(n8519), .A(n8518), .ZN(P2_U3475) );
  AOI21_X1 U10054 ( .B1(n10238), .B2(P2_REG0_REG_31__SCAN_IN), .A(n8520), .ZN(
        n8521) );
  OAI21_X1 U10055 ( .B1(n8522), .B2(n8873), .A(n8521), .ZN(P2_U3458) );
  INV_X1 U10056 ( .A(n8524), .ZN(n8525) );
  OAI21_X1 U10057 ( .B1(n8526), .B2(n8873), .A(n8525), .ZN(P2_U3455) );
  MUX2_X1 U10058 ( .A(n8528), .B(n8527), .S(n10240), .Z(n8529) );
  OAI21_X1 U10059 ( .B1(n8530), .B2(n8873), .A(n8529), .ZN(P2_U3454) );
  MUX2_X1 U10060 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8531), .S(n10240), .Z(
        n8532) );
  INV_X1 U10061 ( .A(n8532), .ZN(n8533) );
  OAI21_X1 U10062 ( .B1(n8534), .B2(n8873), .A(n8533), .ZN(P2_U3453) );
  MUX2_X1 U10063 ( .A(n8536), .B(n8535), .S(n10240), .Z(n8537) );
  OAI21_X1 U10064 ( .B1(n8538), .B2(n8873), .A(n8537), .ZN(P2_U3452) );
  INV_X1 U10065 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8540) );
  MUX2_X1 U10066 ( .A(n8540), .B(n8539), .S(n10240), .Z(n8541) );
  OAI21_X1 U10067 ( .B1(n8542), .B2(n8873), .A(n8541), .ZN(P2_U3451) );
  INV_X1 U10068 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8544) );
  MUX2_X1 U10069 ( .A(n8544), .B(n8543), .S(n10240), .Z(n8545) );
  OAI21_X1 U10070 ( .B1(n8546), .B2(n8873), .A(n8545), .ZN(P2_U3450) );
  INV_X1 U10071 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8548) );
  MUX2_X1 U10072 ( .A(n8548), .B(n8547), .S(n10240), .Z(n8549) );
  OAI21_X1 U10073 ( .B1(n8550), .B2(n8873), .A(n8549), .ZN(P2_U3449) );
  INV_X1 U10074 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8552) );
  MUX2_X1 U10075 ( .A(n8552), .B(n8551), .S(n10240), .Z(n8553) );
  OAI21_X1 U10076 ( .B1(n8554), .B2(n8873), .A(n8553), .ZN(P2_U3448) );
  MUX2_X1 U10077 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8555), .S(n10240), .Z(
        n8860) );
  INV_X1 U10078 ( .A(keyinput75), .ZN(n8556) );
  NAND4_X1 U10079 ( .A1(keyinput74), .A2(keyinput50), .A3(keyinput76), .A4(
        n8556), .ZN(n8616) );
  NOR2_X1 U10080 ( .A1(keyinput20), .A2(keyinput125), .ZN(n8557) );
  NAND3_X1 U10081 ( .A1(keyinput117), .A2(keyinput115), .A3(n8557), .ZN(n8615)
         );
  NAND4_X1 U10082 ( .A1(keyinput103), .A2(keyinput48), .A3(keyinput19), .A4(
        keyinput59), .ZN(n8558) );
  NOR3_X1 U10083 ( .A1(keyinput86), .A2(keyinput69), .A3(n8558), .ZN(n8567) );
  NAND2_X1 U10084 ( .A1(keyinput34), .A2(keyinput51), .ZN(n8559) );
  NOR3_X1 U10085 ( .A1(keyinput32), .A2(keyinput6), .A3(n8559), .ZN(n8564) );
  INV_X1 U10086 ( .A(keyinput78), .ZN(n8560) );
  NOR4_X1 U10087 ( .A1(keyinput113), .A2(keyinput43), .A3(keyinput41), .A4(
        n8560), .ZN(n8563) );
  NOR4_X1 U10088 ( .A1(keyinput39), .A2(keyinput98), .A3(keyinput58), .A4(
        keyinput95), .ZN(n8562) );
  NOR4_X1 U10089 ( .A1(keyinput49), .A2(keyinput118), .A3(keyinput54), .A4(
        keyinput122), .ZN(n8561) );
  NAND4_X1 U10090 ( .A1(n8564), .A2(n8563), .A3(n8562), .A4(n8561), .ZN(n8565)
         );
  NOR2_X1 U10091 ( .A1(n8565), .A2(keyinput61), .ZN(n8566) );
  NAND3_X1 U10092 ( .A1(keyinput100), .A2(n8567), .A3(n8566), .ZN(n8614) );
  NOR4_X1 U10093 ( .A1(keyinput56), .A2(keyinput46), .A3(keyinput36), .A4(
        keyinput0), .ZN(n8568) );
  NAND4_X1 U10094 ( .A1(keyinput38), .A2(keyinput96), .A3(keyinput112), .A4(
        n8568), .ZN(n8580) );
  NOR2_X1 U10095 ( .A1(keyinput108), .A2(keyinput55), .ZN(n8569) );
  NAND3_X1 U10096 ( .A1(keyinput21), .A2(keyinput33), .A3(n8569), .ZN(n8579)
         );
  NOR2_X1 U10097 ( .A1(keyinput102), .A2(keyinput89), .ZN(n8570) );
  NAND3_X1 U10098 ( .A1(keyinput10), .A2(keyinput124), .A3(n8570), .ZN(n8578)
         );
  NOR4_X1 U10099 ( .A1(keyinput12), .A2(keyinput52), .A3(keyinput127), .A4(
        keyinput111), .ZN(n8576) );
  NAND2_X1 U10100 ( .A1(keyinput5), .A2(keyinput64), .ZN(n8571) );
  NOR3_X1 U10101 ( .A1(keyinput71), .A2(keyinput11), .A3(n8571), .ZN(n8575) );
  NAND3_X1 U10102 ( .A1(keyinput24), .A2(keyinput99), .A3(keyinput101), .ZN(
        n8572) );
  NOR2_X1 U10103 ( .A1(keyinput22), .A2(n8572), .ZN(n8574) );
  NOR4_X1 U10104 ( .A1(keyinput31), .A2(keyinput105), .A3(keyinput13), .A4(
        keyinput42), .ZN(n8573) );
  NAND4_X1 U10105 ( .A1(n8576), .A2(n8575), .A3(n8574), .A4(n8573), .ZN(n8577)
         );
  NOR4_X1 U10106 ( .A1(n8580), .A2(n8579), .A3(n8578), .A4(n8577), .ZN(n8612)
         );
  INV_X1 U10107 ( .A(keyinput121), .ZN(n8581) );
  NAND4_X1 U10108 ( .A1(keyinput14), .A2(keyinput1), .A3(keyinput84), .A4(
        n8581), .ZN(n8588) );
  NOR2_X1 U10109 ( .A1(keyinput35), .A2(keyinput30), .ZN(n8582) );
  NAND3_X1 U10110 ( .A1(keyinput94), .A2(keyinput17), .A3(n8582), .ZN(n8587)
         );
  NOR2_X1 U10111 ( .A1(keyinput57), .A2(keyinput66), .ZN(n8583) );
  NAND3_X1 U10112 ( .A1(keyinput3), .A2(keyinput27), .A3(n8583), .ZN(n8586) );
  INV_X1 U10113 ( .A(keyinput85), .ZN(n8584) );
  NAND4_X1 U10114 ( .A1(keyinput53), .A2(keyinput70), .A3(keyinput29), .A4(
        n8584), .ZN(n8585) );
  NOR4_X1 U10115 ( .A1(n8588), .A2(n8587), .A3(n8586), .A4(n8585), .ZN(n8611)
         );
  INV_X1 U10116 ( .A(keyinput28), .ZN(n8589) );
  NOR4_X1 U10117 ( .A1(keyinput15), .A2(keyinput67), .A3(keyinput104), .A4(
        n8589), .ZN(n8590) );
  NAND3_X1 U10118 ( .A1(keyinput126), .A2(keyinput120), .A3(n8590), .ZN(n8594)
         );
  NOR2_X1 U10119 ( .A1(keyinput60), .A2(keyinput114), .ZN(n8592) );
  NOR4_X1 U10120 ( .A1(keyinput83), .A2(keyinput107), .A3(keyinput23), .A4(
        keyinput90), .ZN(n8591) );
  NAND4_X1 U10121 ( .A1(n8592), .A2(keyinput72), .A3(keyinput9), .A4(n8591), 
        .ZN(n8593) );
  NOR4_X1 U10122 ( .A1(keyinput62), .A2(keyinput45), .A3(n8594), .A4(n8593), 
        .ZN(n8610) );
  NAND4_X1 U10123 ( .A1(keyinput44), .A2(keyinput26), .A3(keyinput93), .A4(
        keyinput82), .ZN(n8608) );
  NOR2_X1 U10124 ( .A1(keyinput40), .A2(keyinput81), .ZN(n8595) );
  NAND3_X1 U10125 ( .A1(keyinput109), .A2(keyinput73), .A3(n8595), .ZN(n8607)
         );
  NAND4_X1 U10126 ( .A1(keyinput106), .A2(keyinput7), .A3(keyinput77), .A4(
        keyinput8), .ZN(n8596) );
  NOR3_X1 U10127 ( .A1(keyinput37), .A2(keyinput116), .A3(n8596), .ZN(n8597)
         );
  NAND3_X1 U10128 ( .A1(keyinput65), .A2(keyinput91), .A3(n8597), .ZN(n8606)
         );
  INV_X1 U10129 ( .A(keyinput79), .ZN(n8598) );
  NOR4_X1 U10130 ( .A1(keyinput110), .A2(keyinput47), .A3(keyinput123), .A4(
        n8598), .ZN(n8604) );
  NAND2_X1 U10131 ( .A1(keyinput2), .A2(keyinput87), .ZN(n8599) );
  NOR3_X1 U10132 ( .A1(keyinput63), .A2(keyinput97), .A3(n8599), .ZN(n8603) );
  NOR4_X1 U10133 ( .A1(keyinput4), .A2(keyinput68), .A3(keyinput88), .A4(
        keyinput18), .ZN(n8602) );
  NAND2_X1 U10134 ( .A1(keyinput80), .A2(keyinput119), .ZN(n8600) );
  NOR3_X1 U10135 ( .A1(keyinput16), .A2(keyinput25), .A3(n8600), .ZN(n8601) );
  NAND4_X1 U10136 ( .A1(n8604), .A2(n8603), .A3(n8602), .A4(n8601), .ZN(n8605)
         );
  NOR4_X1 U10137 ( .A1(n8608), .A2(n8607), .A3(n8606), .A4(n8605), .ZN(n8609)
         );
  NAND4_X1 U10138 ( .A1(n8612), .A2(n8611), .A3(n8610), .A4(n8609), .ZN(n8613)
         );
  NOR4_X1 U10139 ( .A1(n8616), .A2(n8615), .A3(n8614), .A4(n8613), .ZN(n8617)
         );
  OAI21_X1 U10140 ( .B1(keyinput92), .B2(n8617), .A(n8644), .ZN(n8858) );
  AOI22_X1 U10141 ( .A1(n8619), .A2(keyinput112), .B1(keyinput71), .B2(n8145), 
        .ZN(n8618) );
  OAI221_X1 U10142 ( .B1(n8619), .B2(keyinput112), .C1(n8145), .C2(keyinput71), 
        .A(n8618), .ZN(n8702) );
  INV_X1 U10143 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8622) );
  INV_X1 U10144 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n8621) );
  AOI22_X1 U10145 ( .A1(n8622), .A2(keyinput0), .B1(n8621), .B2(keyinput96), 
        .ZN(n8620) );
  OAI221_X1 U10146 ( .B1(n8622), .B2(keyinput0), .C1(n8621), .C2(keyinput96), 
        .A(n8620), .ZN(n8701) );
  INV_X1 U10147 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9607) );
  INV_X1 U10148 ( .A(keyinput36), .ZN(n8627) );
  AOI22_X1 U10149 ( .A1(n8625), .A2(keyinput56), .B1(keyinput46), .B2(n8624), 
        .ZN(n8623) );
  OAI221_X1 U10150 ( .B1(n8625), .B2(keyinput56), .C1(n8624), .C2(keyinput46), 
        .A(n8623), .ZN(n8626) );
  AOI221_X1 U10151 ( .B1(keyinput36), .B2(n9607), .C1(n8627), .C2(
        P1_ADDR_REG_3__SCAN_IN), .A(n8626), .ZN(n8643) );
  XNOR2_X1 U10152 ( .A(n8628), .B(keyinput5), .ZN(n8635) );
  XNOR2_X1 U10153 ( .A(P1_REG3_REG_11__SCAN_IN), .B(keyinput10), .ZN(n8630) );
  XNOR2_X1 U10154 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput12), .ZN(n8629) );
  NAND2_X1 U10155 ( .A1(n8630), .A2(n8629), .ZN(n8634) );
  XNOR2_X1 U10156 ( .A(n8631), .B(keyinput11), .ZN(n8633) );
  XNOR2_X1 U10157 ( .A(keyinput64), .B(n5916), .ZN(n8632) );
  OR4_X1 U10158 ( .A1(n8635), .A2(n8634), .A3(n8633), .A4(n8632), .ZN(n8641)
         );
  AOI22_X1 U10159 ( .A1(n8638), .A2(keyinput52), .B1(n8637), .B2(keyinput127), 
        .ZN(n8636) );
  OAI221_X1 U10160 ( .B1(n8638), .B2(keyinput52), .C1(n8637), .C2(keyinput127), 
        .A(n8636), .ZN(n8640) );
  INV_X1 U10161 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n9911) );
  XNOR2_X1 U10162 ( .A(n9911), .B(keyinput111), .ZN(n8639) );
  NOR3_X1 U10163 ( .A1(n8641), .A2(n8640), .A3(n8639), .ZN(n8642) );
  OAI211_X1 U10164 ( .C1(keyinput92), .C2(n8644), .A(n8643), .B(n8642), .ZN(
        n8700) );
  INV_X1 U10165 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n9915) );
  INV_X1 U10166 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9131) );
  AOI22_X1 U10167 ( .A1(n9915), .A2(keyinput94), .B1(keyinput17), .B2(n9131), 
        .ZN(n8645) );
  OAI221_X1 U10168 ( .B1(n9915), .B2(keyinput94), .C1(n9131), .C2(keyinput17), 
        .A(n8645), .ZN(n8655) );
  INV_X1 U10169 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9627) );
  AOI22_X1 U10170 ( .A1(n9627), .A2(keyinput14), .B1(n8647), .B2(keyinput1), 
        .ZN(n8646) );
  OAI221_X1 U10171 ( .B1(n9627), .B2(keyinput14), .C1(n8647), .C2(keyinput1), 
        .A(n8646), .ZN(n8654) );
  AOI22_X1 U10172 ( .A1(n8649), .A2(keyinput30), .B1(n8882), .B2(keyinput121), 
        .ZN(n8648) );
  OAI221_X1 U10173 ( .B1(n8649), .B2(keyinput30), .C1(n8882), .C2(keyinput121), 
        .A(n8648), .ZN(n8653) );
  XNOR2_X1 U10174 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput60), .ZN(n8651) );
  XNOR2_X1 U10175 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(keyinput84), .ZN(n8650)
         );
  NAND2_X1 U10176 ( .A1(n8651), .A2(n8650), .ZN(n8652) );
  NOR4_X1 U10177 ( .A1(n8655), .A2(n8654), .A3(n8653), .A4(n8652), .ZN(n8698)
         );
  INV_X1 U10178 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8657) );
  INV_X1 U10179 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9994) );
  AOI22_X1 U10180 ( .A1(n8657), .A2(keyinput120), .B1(n9994), .B2(keyinput35), 
        .ZN(n8656) );
  OAI221_X1 U10181 ( .B1(n8657), .B2(keyinput120), .C1(n9994), .C2(keyinput35), 
        .A(n8656), .ZN(n8667) );
  INV_X1 U10182 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10231) );
  AOI22_X1 U10183 ( .A1(n8659), .A2(keyinput28), .B1(keyinput67), .B2(n10231), 
        .ZN(n8658) );
  OAI221_X1 U10184 ( .B1(n8659), .B2(keyinput28), .C1(n10231), .C2(keyinput67), 
        .A(n8658), .ZN(n8666) );
  INV_X1 U10185 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n9908) );
  AOI22_X1 U10186 ( .A1(n9908), .A2(keyinput104), .B1(keyinput126), .B2(n8661), 
        .ZN(n8660) );
  OAI221_X1 U10187 ( .B1(n9908), .B2(keyinput104), .C1(n8661), .C2(keyinput126), .A(n8660), .ZN(n8665) );
  XNOR2_X1 U10188 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput15), .ZN(n8663) );
  XNOR2_X1 U10189 ( .A(SI_29_), .B(keyinput45), .ZN(n8662) );
  NAND2_X1 U10190 ( .A1(n8663), .A2(n8662), .ZN(n8664) );
  NOR4_X1 U10191 ( .A1(n8667), .A2(n8666), .A3(n8665), .A4(n8664), .ZN(n8697)
         );
  INV_X1 U10192 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n8670) );
  AOI22_X1 U10193 ( .A1(n8670), .A2(keyinput85), .B1(keyinput57), .B2(n8669), 
        .ZN(n8668) );
  OAI221_X1 U10194 ( .B1(n8670), .B2(keyinput85), .C1(n8669), .C2(keyinput57), 
        .A(n8668), .ZN(n8682) );
  AOI22_X1 U10195 ( .A1(n8673), .A2(keyinput53), .B1(n8672), .B2(keyinput29), 
        .ZN(n8671) );
  OAI221_X1 U10196 ( .B1(n8673), .B2(keyinput53), .C1(n8672), .C2(keyinput29), 
        .A(n8671), .ZN(n8681) );
  INV_X1 U10197 ( .A(keyinput86), .ZN(n8675) );
  AOI22_X1 U10198 ( .A1(n8676), .A2(keyinput27), .B1(P2_ADDR_REG_18__SCAN_IN), 
        .B2(n8675), .ZN(n8674) );
  OAI221_X1 U10199 ( .B1(n8676), .B2(keyinput27), .C1(n8675), .C2(
        P2_ADDR_REG_18__SCAN_IN), .A(n8674), .ZN(n8680) );
  AOI22_X1 U10200 ( .A1(n6939), .A2(keyinput3), .B1(n8678), .B2(keyinput66), 
        .ZN(n8677) );
  OAI221_X1 U10201 ( .B1(n6939), .B2(keyinput3), .C1(n8678), .C2(keyinput66), 
        .A(n8677), .ZN(n8679) );
  NOR4_X1 U10202 ( .A1(n8682), .A2(n8681), .A3(n8680), .A4(n8679), .ZN(n8696)
         );
  AOI22_X1 U10203 ( .A1(n8685), .A2(keyinput107), .B1(n8684), .B2(keyinput23), 
        .ZN(n8683) );
  OAI221_X1 U10204 ( .B1(n8685), .B2(keyinput107), .C1(n8684), .C2(keyinput23), 
        .A(n8683), .ZN(n8694) );
  INV_X1 U10205 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10219) );
  AOI22_X1 U10206 ( .A1(n8687), .A2(keyinput114), .B1(keyinput83), .B2(n10219), 
        .ZN(n8686) );
  OAI221_X1 U10207 ( .B1(n8687), .B2(keyinput114), .C1(n10219), .C2(keyinput83), .A(n8686), .ZN(n8693) );
  AOI22_X1 U10208 ( .A1(n10076), .A2(keyinput9), .B1(keyinput70), .B2(n10241), 
        .ZN(n8688) );
  OAI221_X1 U10209 ( .B1(n10076), .B2(keyinput9), .C1(n10241), .C2(keyinput70), 
        .A(n8688), .ZN(n8692) );
  INV_X1 U10210 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9986) );
  AOI22_X1 U10211 ( .A1(n8690), .A2(keyinput90), .B1(n9986), .B2(keyinput72), 
        .ZN(n8689) );
  OAI221_X1 U10212 ( .B1(n8690), .B2(keyinput90), .C1(n9986), .C2(keyinput72), 
        .A(n8689), .ZN(n8691) );
  NOR4_X1 U10213 ( .A1(n8694), .A2(n8693), .A3(n8692), .A4(n8691), .ZN(n8695)
         );
  NAND4_X1 U10214 ( .A1(n8698), .A2(n8697), .A3(n8696), .A4(n8695), .ZN(n8699)
         );
  NOR4_X1 U10215 ( .A1(n8702), .A2(n8701), .A3(n8700), .A4(n8699), .ZN(n8857)
         );
  INV_X1 U10216 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10169) );
  AOI22_X1 U10217 ( .A1(n9563), .A2(keyinput118), .B1(keyinput54), .B2(n10169), 
        .ZN(n8703) );
  OAI221_X1 U10218 ( .B1(n9563), .B2(keyinput118), .C1(n10169), .C2(keyinput54), .A(n8703), .ZN(n8712) );
  INV_X1 U10219 ( .A(P2_B_REG_SCAN_IN), .ZN(n8705) );
  AOI22_X1 U10220 ( .A1(n8951), .A2(keyinput122), .B1(keyinput39), .B2(n8705), 
        .ZN(n8704) );
  OAI221_X1 U10221 ( .B1(n8951), .B2(keyinput122), .C1(n8705), .C2(keyinput39), 
        .A(n8704), .ZN(n8711) );
  AOI22_X1 U10222 ( .A1(n8707), .A2(keyinput98), .B1(keyinput58), .B2(n8293), 
        .ZN(n8706) );
  OAI221_X1 U10223 ( .B1(n8707), .B2(keyinput98), .C1(n8293), .C2(keyinput58), 
        .A(n8706), .ZN(n8710) );
  INV_X1 U10224 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10044) );
  INV_X1 U10225 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9933) );
  AOI22_X1 U10226 ( .A1(n10044), .A2(keyinput95), .B1(n9933), .B2(keyinput20), 
        .ZN(n8708) );
  OAI221_X1 U10227 ( .B1(n10044), .B2(keyinput95), .C1(n9933), .C2(keyinput20), 
        .A(n8708), .ZN(n8709) );
  NOR4_X1 U10228 ( .A1(n8712), .A2(n8711), .A3(n8710), .A4(n8709), .ZN(n8728)
         );
  AOI22_X1 U10229 ( .A1(n8715), .A2(keyinput40), .B1(n8714), .B2(keyinput73), 
        .ZN(n8713) );
  OAI221_X1 U10230 ( .B1(n8715), .B2(keyinput40), .C1(n8714), .C2(keyinput73), 
        .A(n8713), .ZN(n8726) );
  AOI22_X1 U10231 ( .A1(n8718), .A2(keyinput81), .B1(keyinput44), .B2(n8717), 
        .ZN(n8716) );
  OAI221_X1 U10232 ( .B1(n8718), .B2(keyinput81), .C1(n8717), .C2(keyinput44), 
        .A(n8716), .ZN(n8725) );
  INV_X1 U10233 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n9916) );
  AOI22_X1 U10234 ( .A1(n8720), .A2(keyinput26), .B1(n9916), .B2(keyinput93), 
        .ZN(n8719) );
  OAI221_X1 U10235 ( .B1(n8720), .B2(keyinput26), .C1(n9916), .C2(keyinput93), 
        .A(n8719), .ZN(n8724) );
  INV_X1 U10236 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10213) );
  AOI22_X1 U10237 ( .A1(n10213), .A2(keyinput82), .B1(n8722), .B2(keyinput87), 
        .ZN(n8721) );
  OAI221_X1 U10238 ( .B1(n10213), .B2(keyinput82), .C1(n8722), .C2(keyinput87), 
        .A(n8721), .ZN(n8723) );
  NOR4_X1 U10239 ( .A1(n8726), .A2(n8725), .A3(n8724), .A4(n8723), .ZN(n8727)
         );
  AND2_X1 U10240 ( .A1(n8728), .A2(n8727), .ZN(n8855) );
  AOI22_X1 U10241 ( .A1(n8731), .A2(keyinput117), .B1(n8730), .B2(keyinput125), 
        .ZN(n8729) );
  OAI221_X1 U10242 ( .B1(n8731), .B2(keyinput117), .C1(n8730), .C2(keyinput125), .A(n8729), .ZN(n8741) );
  INV_X1 U10243 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9123) );
  AOI22_X1 U10244 ( .A1(n8733), .A2(keyinput115), .B1(n9123), .B2(keyinput74), 
        .ZN(n8732) );
  OAI221_X1 U10245 ( .B1(n8733), .B2(keyinput115), .C1(n9123), .C2(keyinput74), 
        .A(n8732), .ZN(n8740) );
  INV_X1 U10246 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n9909) );
  AOI22_X1 U10247 ( .A1(n8735), .A2(keyinput75), .B1(n9909), .B2(keyinput50), 
        .ZN(n8734) );
  OAI221_X1 U10248 ( .B1(n8735), .B2(keyinput75), .C1(n9909), .C2(keyinput50), 
        .A(n8734), .ZN(n8739) );
  INV_X1 U10249 ( .A(keyinput109), .ZN(n8737) );
  AOI22_X1 U10250 ( .A1(n9561), .A2(keyinput76), .B1(P2_ADDR_REG_15__SCAN_IN), 
        .B2(n8737), .ZN(n8736) );
  OAI221_X1 U10251 ( .B1(n9561), .B2(keyinput76), .C1(n8737), .C2(
        P2_ADDR_REG_15__SCAN_IN), .A(n8736), .ZN(n8738) );
  NOR4_X1 U10252 ( .A1(n8741), .A2(n8740), .A3(n8739), .A4(n8738), .ZN(n8854)
         );
  INV_X1 U10253 ( .A(keyinput4), .ZN(n8743) );
  AOI22_X1 U10254 ( .A1(n8744), .A2(keyinput16), .B1(P1_ADDR_REG_13__SCAN_IN), 
        .B2(n8743), .ZN(n8742) );
  OAI221_X1 U10255 ( .B1(n8744), .B2(keyinput16), .C1(n8743), .C2(
        P1_ADDR_REG_13__SCAN_IN), .A(n8742), .ZN(n8757) );
  INV_X1 U10256 ( .A(keyinput68), .ZN(n8746) );
  AOI22_X1 U10257 ( .A1(n8747), .A2(keyinput80), .B1(P1_ADDR_REG_16__SCAN_IN), 
        .B2(n8746), .ZN(n8745) );
  OAI221_X1 U10258 ( .B1(n8747), .B2(keyinput80), .C1(n8746), .C2(
        P1_ADDR_REG_16__SCAN_IN), .A(n8745), .ZN(n8756) );
  INV_X1 U10259 ( .A(SI_22_), .ZN(n8749) );
  AOI22_X1 U10260 ( .A1(n8750), .A2(keyinput25), .B1(n8749), .B2(keyinput88), 
        .ZN(n8748) );
  OAI221_X1 U10261 ( .B1(n8750), .B2(keyinput25), .C1(n8749), .C2(keyinput88), 
        .A(n8748), .ZN(n8755) );
  AOI22_X1 U10262 ( .A1(n8753), .A2(keyinput18), .B1(n8752), .B2(keyinput65), 
        .ZN(n8751) );
  OAI221_X1 U10263 ( .B1(n8753), .B2(keyinput18), .C1(n8752), .C2(keyinput65), 
        .A(n8751), .ZN(n8754) );
  NOR4_X1 U10264 ( .A1(n8757), .A2(n8756), .A3(n8755), .A4(n8754), .ZN(n8853)
         );
  AOI22_X1 U10265 ( .A1(n8760), .A2(keyinput48), .B1(n8759), .B2(keyinput100), 
        .ZN(n8758) );
  OAI221_X1 U10266 ( .B1(n8760), .B2(keyinput48), .C1(n8759), .C2(keyinput100), 
        .A(n8758), .ZN(n8767) );
  INV_X1 U10267 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n8762) );
  AOI22_X1 U10268 ( .A1(n8763), .A2(keyinput105), .B1(n8762), .B2(keyinput99), 
        .ZN(n8761) );
  OAI221_X1 U10269 ( .B1(n8763), .B2(keyinput105), .C1(n8762), .C2(keyinput99), 
        .A(n8761), .ZN(n8766) );
  XNOR2_X1 U10270 ( .A(n8764), .B(keyinput49), .ZN(n8765) );
  NOR3_X1 U10271 ( .A1(n8767), .A2(n8766), .A3(n8765), .ZN(n8814) );
  INV_X1 U10272 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n8769) );
  AOI22_X1 U10273 ( .A1(n8770), .A2(keyinput41), .B1(n8769), .B2(keyinput32), 
        .ZN(n8768) );
  OAI221_X1 U10274 ( .B1(n8770), .B2(keyinput41), .C1(n8769), .C2(keyinput32), 
        .A(n8768), .ZN(n8774) );
  AOI22_X1 U10275 ( .A1(n8271), .A2(keyinput97), .B1(n8772), .B2(keyinput63), 
        .ZN(n8771) );
  OAI221_X1 U10276 ( .B1(n8271), .B2(keyinput97), .C1(n8772), .C2(keyinput63), 
        .A(n8771), .ZN(n8773) );
  NOR2_X1 U10277 ( .A1(n8774), .A2(n8773), .ZN(n8784) );
  INV_X1 U10278 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n8777) );
  AOI22_X1 U10279 ( .A1(n8777), .A2(keyinput51), .B1(n8776), .B2(keyinput34), 
        .ZN(n8775) );
  OAI221_X1 U10280 ( .B1(n8777), .B2(keyinput51), .C1(n8776), .C2(keyinput34), 
        .A(n8775), .ZN(n8782) );
  AOI22_X1 U10281 ( .A1(n8780), .A2(keyinput116), .B1(keyinput106), .B2(n8779), 
        .ZN(n8778) );
  OAI221_X1 U10282 ( .B1(n8780), .B2(keyinput116), .C1(n8779), .C2(keyinput106), .A(n8778), .ZN(n8781) );
  NOR2_X1 U10283 ( .A1(n8782), .A2(n8781), .ZN(n8783) );
  AND2_X1 U10284 ( .A1(n8784), .A2(n8783), .ZN(n8813) );
  INV_X1 U10285 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n8786) );
  INV_X1 U10286 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9647) );
  AOI22_X1 U10287 ( .A1(n8786), .A2(keyinput89), .B1(keyinput21), .B2(n9647), 
        .ZN(n8785) );
  OAI221_X1 U10288 ( .B1(n8786), .B2(keyinput89), .C1(n9647), .C2(keyinput21), 
        .A(n8785), .ZN(n8790) );
  INV_X1 U10289 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n9910) );
  AOI22_X1 U10290 ( .A1(n9910), .A2(keyinput47), .B1(keyinput110), .B2(n8788), 
        .ZN(n8787) );
  OAI221_X1 U10291 ( .B1(n9910), .B2(keyinput47), .C1(n8788), .C2(keyinput110), 
        .A(n8787), .ZN(n8789) );
  NOR2_X1 U10292 ( .A1(n8790), .A2(n8789), .ZN(n8812) );
  INV_X1 U10293 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8792) );
  AOI22_X1 U10294 ( .A1(n8793), .A2(keyinput69), .B1(n8792), .B2(keyinput103), 
        .ZN(n8791) );
  OAI221_X1 U10295 ( .B1(n8793), .B2(keyinput69), .C1(n8792), .C2(keyinput103), 
        .A(n8791), .ZN(n8798) );
  XNOR2_X1 U10296 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput62), .ZN(n8796) );
  XNOR2_X1 U10297 ( .A(P2_IR_REG_13__SCAN_IN), .B(keyinput55), .ZN(n8795) );
  XNOR2_X1 U10298 ( .A(keyinput42), .B(P2_REG0_REG_13__SCAN_IN), .ZN(n8794) );
  NAND3_X1 U10299 ( .A1(n8796), .A2(n8795), .A3(n8794), .ZN(n8797) );
  NOR2_X1 U10300 ( .A1(n8798), .A2(n8797), .ZN(n8810) );
  XNOR2_X1 U10301 ( .A(P1_REG1_REG_27__SCAN_IN), .B(keyinput31), .ZN(n8802) );
  XNOR2_X1 U10302 ( .A(P2_IR_REG_20__SCAN_IN), .B(keyinput119), .ZN(n8801) );
  XNOR2_X1 U10303 ( .A(P1_REG3_REG_15__SCAN_IN), .B(keyinput123), .ZN(n8800)
         );
  XNOR2_X1 U10304 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(keyinput91), .ZN(n8799) );
  NAND4_X1 U10305 ( .A1(n8802), .A2(n8801), .A3(n8800), .A4(n8799), .ZN(n8808)
         );
  XNOR2_X1 U10306 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput37), .ZN(n8806) );
  XNOR2_X1 U10307 ( .A(P2_IR_REG_5__SCAN_IN), .B(keyinput19), .ZN(n8805) );
  XNOR2_X1 U10308 ( .A(P2_IR_REG_15__SCAN_IN), .B(keyinput6), .ZN(n8804) );
  XNOR2_X1 U10309 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput59), .ZN(n8803) );
  NAND4_X1 U10310 ( .A1(n8806), .A2(n8805), .A3(n8804), .A4(n8803), .ZN(n8807)
         );
  NOR2_X1 U10311 ( .A1(n8808), .A2(n8807), .ZN(n8809) );
  AND2_X1 U10312 ( .A1(n8810), .A2(n8809), .ZN(n8811) );
  NAND4_X1 U10313 ( .A1(n8814), .A2(n8813), .A3(n8812), .A4(n8811), .ZN(n8851)
         );
  AOI22_X1 U10314 ( .A1(n8816), .A2(keyinput101), .B1(n9071), .B2(keyinput24), 
        .ZN(n8815) );
  OAI221_X1 U10315 ( .B1(n8816), .B2(keyinput101), .C1(n9071), .C2(keyinput24), 
        .A(n8815), .ZN(n8817) );
  INV_X1 U10316 ( .A(n8817), .ZN(n8822) );
  INV_X1 U10317 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10200) );
  XNOR2_X1 U10318 ( .A(keyinput113), .B(n10200), .ZN(n8820) );
  XNOR2_X1 U10319 ( .A(keyinput61), .B(n8818), .ZN(n8819) );
  NOR2_X1 U10320 ( .A1(n8820), .A2(n8819), .ZN(n8821) );
  NAND2_X1 U10321 ( .A1(n8822), .A2(n8821), .ZN(n8825) );
  INV_X1 U10322 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n9912) );
  INV_X1 U10323 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10239) );
  AOI22_X1 U10324 ( .A1(n9912), .A2(keyinput22), .B1(keyinput13), .B2(n10239), 
        .ZN(n8823) );
  OAI221_X1 U10325 ( .B1(n9912), .B2(keyinput22), .C1(n10239), .C2(keyinput13), 
        .A(n8823), .ZN(n8824) );
  NOR2_X1 U10326 ( .A1(n8825), .A2(n8824), .ZN(n8849) );
  AOI22_X1 U10327 ( .A1(n8828), .A2(keyinput2), .B1(keyinput79), .B2(n8827), 
        .ZN(n8826) );
  OAI221_X1 U10328 ( .B1(n8828), .B2(keyinput2), .C1(n8827), .C2(keyinput79), 
        .A(n8826), .ZN(n8831) );
  INV_X1 U10329 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n9913) );
  INV_X1 U10330 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n9914) );
  AOI22_X1 U10331 ( .A1(n9913), .A2(keyinput7), .B1(keyinput77), .B2(n9914), 
        .ZN(n8829) );
  OAI221_X1 U10332 ( .B1(n9913), .B2(keyinput7), .C1(n9914), .C2(keyinput77), 
        .A(n8829), .ZN(n8830) );
  NOR2_X1 U10333 ( .A1(n8831), .A2(n8830), .ZN(n8848) );
  INV_X1 U10334 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n8833) );
  AOI22_X1 U10335 ( .A1(n8833), .A2(keyinput38), .B1(keyinput8), .B2(n5929), 
        .ZN(n8832) );
  OAI221_X1 U10336 ( .B1(n8833), .B2(keyinput38), .C1(n5929), .C2(keyinput8), 
        .A(n8832), .ZN(n8838) );
  AOI22_X1 U10337 ( .A1(n8836), .A2(keyinput43), .B1(n8835), .B2(keyinput78), 
        .ZN(n8834) );
  OAI221_X1 U10338 ( .B1(n8836), .B2(keyinput43), .C1(n8835), .C2(keyinput78), 
        .A(n8834), .ZN(n8837) );
  NOR2_X1 U10339 ( .A1(n8838), .A2(n8837), .ZN(n8847) );
  INV_X1 U10340 ( .A(keyinput108), .ZN(n8840) );
  AOI22_X1 U10341 ( .A1(n8841), .A2(keyinput33), .B1(SI_31_), .B2(n8840), .ZN(
        n8839) );
  OAI221_X1 U10342 ( .B1(n8841), .B2(keyinput33), .C1(n8840), .C2(SI_31_), .A(
        n8839), .ZN(n8845) );
  AOI22_X1 U10343 ( .A1(n8843), .A2(keyinput102), .B1(n6328), .B2(keyinput124), 
        .ZN(n8842) );
  OAI221_X1 U10344 ( .B1(n8843), .B2(keyinput102), .C1(n6328), .C2(keyinput124), .A(n8842), .ZN(n8844) );
  NOR2_X1 U10345 ( .A1(n8845), .A2(n8844), .ZN(n8846) );
  NAND4_X1 U10346 ( .A1(n8849), .A2(n8848), .A3(n8847), .A4(n8846), .ZN(n8850)
         );
  NOR2_X1 U10347 ( .A1(n8851), .A2(n8850), .ZN(n8852) );
  AND4_X1 U10348 ( .A1(n8855), .A2(n8854), .A3(n8853), .A4(n8852), .ZN(n8856)
         );
  NAND3_X1 U10349 ( .A1(n8858), .A2(n8857), .A3(n8856), .ZN(n8859) );
  XNOR2_X1 U10350 ( .A(n8860), .B(n8859), .ZN(P2_U3447) );
  INV_X1 U10351 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8862) );
  MUX2_X1 U10352 ( .A(n8862), .B(n8861), .S(n10240), .Z(n8863) );
  OAI21_X1 U10353 ( .B1(n8864), .B2(n8873), .A(n8863), .ZN(P2_U3446) );
  INV_X1 U10354 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8866) );
  MUX2_X1 U10355 ( .A(n8866), .B(n8865), .S(n10240), .Z(n8867) );
  OAI21_X1 U10356 ( .B1(n8868), .B2(n8873), .A(n8867), .ZN(P2_U3444) );
  MUX2_X1 U10357 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8869), .S(n10240), .Z(
        P2_U3441) );
  INV_X1 U10358 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8871) );
  MUX2_X1 U10359 ( .A(n8871), .B(n8870), .S(n10240), .Z(n8872) );
  OAI21_X1 U10360 ( .B1(n8874), .B2(n8873), .A(n8872), .ZN(P2_U3438) );
  INV_X1 U10361 ( .A(n8875), .ZN(n9555) );
  NOR4_X1 U10362 ( .A1(n5944), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n8876), .ZN(n8877) );
  AOI21_X1 U10363 ( .B1(n8884), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8877), .ZN(
        n8878) );
  OAI21_X1 U10364 ( .B1(n9555), .B2(n8890), .A(n8878), .ZN(P2_U3264) );
  NAND2_X1 U10365 ( .A1(n9559), .A2(n8879), .ZN(n8881) );
  OAI211_X1 U10366 ( .C1(n8882), .C2(n8888), .A(n8881), .B(n8880), .ZN(
        P2_U3267) );
  AOI21_X1 U10367 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n8884), .A(n8883), .ZN(
        n8885) );
  OAI21_X1 U10368 ( .B1(n8886), .B2(n8890), .A(n8885), .ZN(P2_U3268) );
  INV_X1 U10369 ( .A(n8887), .ZN(n9564) );
  OAI222_X1 U10370 ( .A1(n8890), .A2(n9564), .B1(P2_U3151), .B2(n6808), .C1(
        n8889), .C2(n8888), .ZN(P2_U3269) );
  INV_X1 U10371 ( .A(n8892), .ZN(n8893) );
  NAND2_X1 U10372 ( .A1(n9039), .A2(n8893), .ZN(n8895) );
  AOI21_X1 U10373 ( .B1(n8896), .B2(n8895), .A(n8894), .ZN(n8902) );
  OAI22_X1 U10374 ( .A1(n9041), .A2(n9455), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8897), .ZN(n8900) );
  INV_X1 U10375 ( .A(n9229), .ZN(n8898) );
  OAI22_X1 U10376 ( .A1(n9029), .A2(n8898), .B1(n9236), .B2(n9053), .ZN(n8899)
         );
  AOI211_X1 U10377 ( .C1(n9228), .C2(n4451), .A(n8900), .B(n8899), .ZN(n8901)
         );
  OAI21_X1 U10378 ( .B1(n8902), .B2(n9056), .A(n8901), .ZN(P1_U3214) );
  OAI21_X1 U10379 ( .B1(n8905), .B2(n8904), .A(n8903), .ZN(n8906) );
  NAND2_X1 U10380 ( .A1(n8906), .A2(n9038), .ZN(n8913) );
  NAND2_X1 U10381 ( .A1(n4454), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9781) );
  INV_X1 U10382 ( .A(n9781), .ZN(n8911) );
  INV_X1 U10383 ( .A(n8907), .ZN(n8908) );
  OAI22_X1 U10384 ( .A1(n9041), .A2(n8909), .B1(n9029), .B2(n8908), .ZN(n8910)
         );
  AOI211_X1 U10385 ( .C1(n9021), .C2(n9409), .A(n8911), .B(n8910), .ZN(n8912)
         );
  OAI211_X1 U10386 ( .C1(n4951), .C2(n9046), .A(n8913), .B(n8912), .ZN(
        P1_U3215) );
  INV_X1 U10387 ( .A(n8980), .ZN(n8916) );
  NOR3_X1 U10388 ( .A1(n9004), .A2(n9008), .A3(n8914), .ZN(n8915) );
  OAI21_X1 U10389 ( .B1(n8916), .B2(n8915), .A(n9038), .ZN(n8920) );
  INV_X1 U10390 ( .A(n9469), .ZN(n9170) );
  AOI22_X1 U10391 ( .A1(n9021), .A2(n9170), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        n4454), .ZN(n8919) );
  AOI22_X1 U10392 ( .A1(n9163), .A2(n9051), .B1(n9293), .B2(n9050), .ZN(n8918)
         );
  NAND2_X1 U10393 ( .A1(n9299), .A2(n4451), .ZN(n8917) );
  NAND4_X1 U10394 ( .A1(n8920), .A2(n8919), .A3(n8918), .A4(n8917), .ZN(
        P1_U3216) );
  XNOR2_X1 U10395 ( .A(n9015), .B(n9016), .ZN(n8923) );
  NOR2_X1 U10396 ( .A1(n8923), .A2(n8922), .ZN(n9014) );
  AOI21_X1 U10397 ( .B1(n8923), .B2(n8922), .A(n9014), .ZN(n8929) );
  AOI22_X1 U10398 ( .A1(n9021), .A2(n9995), .B1(n9050), .B2(n8924), .ZN(n8925)
         );
  NAND2_X1 U10399 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n9576) );
  OAI211_X1 U10400 ( .C1(n8926), .C2(n9041), .A(n8925), .B(n9576), .ZN(n8927)
         );
  AOI21_X1 U10401 ( .B1(n9980), .B2(n4451), .A(n8927), .ZN(n8928) );
  OAI21_X1 U10402 ( .B1(n8929), .B2(n9056), .A(n8928), .ZN(P1_U3217) );
  INV_X1 U10403 ( .A(n8930), .ZN(n8932) );
  XOR2_X1 U10404 ( .A(n8930), .B(n8931), .Z(n9028) );
  NOR2_X1 U10405 ( .A1(n9028), .A2(n9027), .ZN(n9026) );
  AOI21_X1 U10406 ( .B1(n8932), .B2(n8931), .A(n9026), .ZN(n8936) );
  XNOR2_X1 U10407 ( .A(n8934), .B(n8933), .ZN(n8935) );
  XNOR2_X1 U10408 ( .A(n8936), .B(n8935), .ZN(n8940) );
  NAND2_X1 U10409 ( .A1(n4454), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9094) );
  OAI21_X1 U10410 ( .B1(n9324), .B2(n9053), .A(n9094), .ZN(n8938) );
  OAI22_X1 U10411 ( .A1(n9041), .A2(n9358), .B1(n9029), .B2(n9355), .ZN(n8937)
         );
  AOI211_X1 U10412 ( .C1(n9507), .C2(n4451), .A(n8938), .B(n8937), .ZN(n8939)
         );
  OAI21_X1 U10413 ( .B1(n8940), .B2(n9056), .A(n8939), .ZN(P1_U3219) );
  XOR2_X1 U10414 ( .A(n8942), .B(n8941), .Z(n8947) );
  INV_X1 U10415 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8943) );
  OAI22_X1 U10416 ( .A1(n9481), .A2(n9053), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8943), .ZN(n8945) );
  OAI22_X1 U10417 ( .A1(n9324), .A2(n9041), .B1(n9029), .B2(n9327), .ZN(n8944)
         );
  AOI211_X1 U10418 ( .C1(n9497), .C2(n4451), .A(n8945), .B(n8944), .ZN(n8946)
         );
  OAI21_X1 U10419 ( .B1(n8947), .B2(n9056), .A(n8946), .ZN(P1_U3223) );
  AOI21_X1 U10420 ( .B1(n8950), .B2(n8949), .A(n8948), .ZN(n8956) );
  OAI22_X1 U10421 ( .A1(n9053), .A2(n9455), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8951), .ZN(n8954) );
  INV_X1 U10422 ( .A(n9260), .ZN(n8952) );
  OAI22_X1 U10423 ( .A1(n9041), .A2(n9469), .B1(n9029), .B2(n8952), .ZN(n8953)
         );
  AOI211_X1 U10424 ( .C1(n9259), .C2(n4451), .A(n8954), .B(n8953), .ZN(n8955)
         );
  OAI21_X1 U10425 ( .B1(n8956), .B2(n9056), .A(n8955), .ZN(P1_U3225) );
  INV_X1 U10426 ( .A(n8957), .ZN(n8959) );
  XOR2_X1 U10427 ( .A(n8957), .B(n8958), .Z(n9049) );
  NOR2_X1 U10428 ( .A1(n9049), .A2(n9048), .ZN(n9047) );
  AOI21_X1 U10429 ( .B1(n8959), .B2(n8958), .A(n9047), .ZN(n8963) );
  XNOR2_X1 U10430 ( .A(n8961), .B(n8960), .ZN(n8962) );
  XNOR2_X1 U10431 ( .A(n8963), .B(n8962), .ZN(n8964) );
  NAND2_X1 U10432 ( .A1(n8964), .A2(n9038), .ZN(n8968) );
  INV_X1 U10433 ( .A(n9376), .ZN(n9513) );
  AND2_X1 U10434 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9802) );
  INV_X1 U10435 ( .A(n9403), .ZN(n8965) );
  OAI22_X1 U10436 ( .A1(n9041), .A2(n9152), .B1(n9029), .B2(n8965), .ZN(n8966)
         );
  AOI211_X1 U10437 ( .C1(n9021), .C2(n9513), .A(n9802), .B(n8966), .ZN(n8967)
         );
  OAI211_X1 U10438 ( .C1(n9405), .C2(n9046), .A(n8968), .B(n8967), .ZN(
        P1_U3226) );
  INV_X1 U10439 ( .A(n8969), .ZN(n8971) );
  NOR2_X1 U10440 ( .A1(n8971), .A2(n8970), .ZN(n8972) );
  XNOR2_X1 U10441 ( .A(n8973), .B(n8972), .ZN(n8977) );
  AOI22_X1 U10442 ( .A1(n9051), .A2(n9388), .B1(n9050), .B2(n9392), .ZN(n8974)
         );
  NAND2_X1 U10443 ( .A1(n4454), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9821) );
  OAI211_X1 U10444 ( .C1(n9358), .C2(n9053), .A(n8974), .B(n9821), .ZN(n8975)
         );
  AOI21_X1 U10445 ( .B1(n9385), .B2(n4451), .A(n8975), .ZN(n8976) );
  OAI21_X1 U10446 ( .B1(n8977), .B2(n9056), .A(n8976), .ZN(P1_U3228) );
  AND3_X1 U10447 ( .A1(n8980), .A2(n8979), .A3(n8978), .ZN(n8981) );
  OAI21_X1 U10448 ( .B1(n8982), .B2(n8981), .A(n9038), .ZN(n8986) );
  INV_X1 U10449 ( .A(n9462), .ZN(n9173) );
  AOI22_X1 U10450 ( .A1(n9021), .A2(n9173), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n8985) );
  INV_X1 U10451 ( .A(n9315), .ZN(n9166) );
  AOI22_X1 U10452 ( .A1(n9050), .A2(n9278), .B1(n9051), .B2(n9166), .ZN(n8984)
         );
  NAND2_X1 U10453 ( .A1(n9478), .A2(n4451), .ZN(n8983) );
  NAND4_X1 U10454 ( .A1(n8986), .A2(n8985), .A3(n8984), .A4(n8983), .ZN(
        P1_U3229) );
  XNOR2_X1 U10455 ( .A(n8989), .B(n8988), .ZN(n8990) );
  XNOR2_X1 U10456 ( .A(n8987), .B(n8990), .ZN(n8995) );
  INV_X1 U10457 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8991) );
  OAI22_X1 U10458 ( .A1(n9488), .A2(n9053), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8991), .ZN(n8993) );
  OAI22_X1 U10459 ( .A1(n9041), .A2(n9158), .B1(n9029), .B2(n9336), .ZN(n8992)
         );
  AOI211_X1 U10460 ( .C1(n9500), .C2(n4451), .A(n8993), .B(n8992), .ZN(n8994)
         );
  OAI21_X1 U10461 ( .B1(n8995), .B2(n9056), .A(n8994), .ZN(P1_U3233) );
  XOR2_X1 U10462 ( .A(n8996), .B(n8997), .Z(n9003) );
  AOI22_X1 U10463 ( .A1(n9021), .A2(n9150), .B1(n9050), .B2(n8998), .ZN(n8999)
         );
  NAND2_X1 U10464 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(n4454), .ZN(n9766) );
  OAI211_X1 U10465 ( .C1(n9844), .C2(n9041), .A(n8999), .B(n9766), .ZN(n9000)
         );
  AOI21_X1 U10466 ( .B1(n9001), .B2(n4451), .A(n9000), .ZN(n9002) );
  OAI21_X1 U10467 ( .B1(n9003), .B2(n9056), .A(n9002), .ZN(P1_U3234) );
  OAI21_X1 U10468 ( .B1(n9006), .B2(n9008), .A(n9005), .ZN(n9007) );
  OAI21_X1 U10469 ( .B1(n4850), .B2(n9008), .A(n9007), .ZN(n9012) );
  INV_X1 U10470 ( .A(n9304), .ZN(n9489) );
  AOI22_X1 U10471 ( .A1(n9021), .A2(n9166), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        n4454), .ZN(n9010) );
  AOI22_X1 U10472 ( .A1(n9051), .A2(n9342), .B1(n9050), .B2(n9305), .ZN(n9009)
         );
  OAI211_X1 U10473 ( .C1(n9489), .C2(n9046), .A(n9010), .B(n9009), .ZN(n9011)
         );
  AOI21_X1 U10474 ( .B1(n9012), .B2(n9038), .A(n9011), .ZN(n9013) );
  INV_X1 U10475 ( .A(n9013), .ZN(P1_U3235) );
  AOI21_X1 U10476 ( .B1(n9016), .B2(n9015), .A(n9014), .ZN(n9020) );
  XNOR2_X1 U10477 ( .A(n9018), .B(n9017), .ZN(n9019) );
  XNOR2_X1 U10478 ( .A(n9020), .B(n9019), .ZN(n9025) );
  AOI22_X1 U10479 ( .A1(n9021), .A2(n9059), .B1(n9050), .B2(n9853), .ZN(n9022)
         );
  NAND2_X1 U10480 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9734) );
  OAI211_X1 U10481 ( .C1(n9845), .C2(n9041), .A(n9022), .B(n9734), .ZN(n9023)
         );
  AOI21_X1 U10482 ( .B1(n9988), .B2(n4451), .A(n9023), .ZN(n9024) );
  OAI21_X1 U10483 ( .B1(n9025), .B2(n9056), .A(n9024), .ZN(P1_U3236) );
  AOI21_X1 U10484 ( .B1(n9028), .B2(n9027), .A(n9026), .ZN(n9034) );
  NAND2_X1 U10485 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9837) );
  OAI21_X1 U10486 ( .B1(n9041), .B2(n9376), .A(n9837), .ZN(n9031) );
  OAI22_X1 U10487 ( .A1(n9053), .A2(n9158), .B1(n9029), .B2(n9373), .ZN(n9030)
         );
  AOI211_X1 U10488 ( .C1(n9514), .C2(n4451), .A(n9031), .B(n9030), .ZN(n9033)
         );
  OAI21_X1 U10489 ( .B1(n9034), .B2(n9056), .A(n9033), .ZN(P1_U3238) );
  OAI21_X1 U10490 ( .B1(n8948), .B2(n9036), .A(n9035), .ZN(n9037) );
  NAND3_X1 U10491 ( .A1(n9039), .A2(n9038), .A3(n9037), .ZN(n9045) );
  NOR2_X1 U10492 ( .A1(n9053), .A2(n9252), .ZN(n9043) );
  OAI22_X1 U10493 ( .A1(n9041), .A2(n9462), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9040), .ZN(n9042) );
  AOI211_X1 U10494 ( .C1(n9050), .C2(n9245), .A(n9043), .B(n9042), .ZN(n9044)
         );
  OAI211_X1 U10495 ( .C1(n9463), .C2(n9046), .A(n9045), .B(n9044), .ZN(
        P1_U3240) );
  AOI21_X1 U10496 ( .B1(n9049), .B2(n9048), .A(n9047), .ZN(n9057) );
  AOI22_X1 U10497 ( .A1(n9051), .A2(n9150), .B1(n9050), .B2(n9423), .ZN(n9052)
         );
  NAND2_X1 U10498 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9794) );
  OAI211_X1 U10499 ( .C1(n9421), .C2(n9053), .A(n9052), .B(n9794), .ZN(n9054)
         );
  AOI21_X1 U10500 ( .B1(n9426), .B2(n4451), .A(n9054), .ZN(n9055) );
  OAI21_X1 U10501 ( .B1(n9057), .B2(n9056), .A(n9055), .ZN(P1_U3241) );
  MUX2_X1 U10502 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9140), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U10503 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9196), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10504 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9210), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10505 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9198), .S(P1_U3973), .Z(
        P1_U3582) );
  INV_X1 U10506 ( .A(n9252), .ZN(n9449) );
  MUX2_X1 U10507 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9449), .S(P1_U3973), .Z(
        P1_U3581) );
  INV_X1 U10508 ( .A(n9455), .ZN(n9174) );
  MUX2_X1 U10509 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9174), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10510 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9173), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10511 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9170), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10512 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9166), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10513 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9163), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10514 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9342), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10515 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9351), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10516 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9369), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10517 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9506), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10518 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9513), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10519 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9388), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10520 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9409), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10521 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9150), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10522 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9058), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10523 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9059), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10524 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9995), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10525 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9060), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10526 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9971), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10527 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9061), .S(n9064), .Z(
        P1_U3561) );
  MUX2_X1 U10528 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9865), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10529 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9062), .S(n9064), .Z(
        P1_U3559) );
  MUX2_X1 U10530 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9863), .S(n9064), .Z(
        P1_U3558) );
  MUX2_X1 U10531 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9063), .S(n9064), .Z(
        P1_U3557) );
  MUX2_X1 U10532 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9934), .S(n9064), .Z(
        P1_U3556) );
  MUX2_X1 U10533 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9065), .S(n9064), .Z(
        P1_U3555) );
  NAND3_X1 U10534 ( .A1(n9067), .A2(n9066), .A3(n4459), .ZN(n9074) );
  NAND2_X1 U10535 ( .A1(n9069), .A2(n9068), .ZN(n9073) );
  NOR2_X1 U10536 ( .A1(n4459), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9070) );
  OR2_X1 U10537 ( .A1(n5882), .A2(n9070), .ZN(n9656) );
  NAND2_X1 U10538 ( .A1(n9656), .A2(n9071), .ZN(n9072) );
  NAND4_X1 U10539 ( .A1(n9074), .A2(P1_U3973), .A3(n9073), .A4(n9072), .ZN(
        n9689) );
  NAND2_X1 U10540 ( .A1(n9803), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n9076) );
  NAND2_X1 U10541 ( .A1(P1_U3086), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9075) );
  OAI211_X1 U10542 ( .C1(n9835), .C2(n9077), .A(n9076), .B(n9075), .ZN(n9078)
         );
  INV_X1 U10543 ( .A(n9078), .ZN(n9093) );
  INV_X1 U10544 ( .A(n9079), .ZN(n9082) );
  INV_X1 U10545 ( .A(n9080), .ZN(n9081) );
  NAND2_X1 U10546 ( .A1(n9082), .A2(n9081), .ZN(n9083) );
  NAND3_X1 U10547 ( .A1(n9825), .A2(n9084), .A3(n9083), .ZN(n9092) );
  INV_X1 U10548 ( .A(n9085), .ZN(n9088) );
  INV_X1 U10549 ( .A(n9086), .ZN(n9087) );
  NAND2_X1 U10550 ( .A1(n9088), .A2(n9087), .ZN(n9089) );
  NAND3_X1 U10551 ( .A1(n9829), .A2(n9090), .A3(n9089), .ZN(n9091) );
  NAND4_X1 U10552 ( .A1(n9689), .A2(n9093), .A3(n9092), .A4(n9091), .ZN(
        P1_U3245) );
  OR2_X1 U10553 ( .A1(n9819), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9108) );
  NOR2_X1 U10554 ( .A1(n9819), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9095) );
  AOI21_X1 U10555 ( .B1(n9819), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9095), .ZN(
        n9815) );
  INV_X1 U10556 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9096) );
  AOI22_X1 U10557 ( .A1(n9807), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9096), .B2(
        n9130), .ZN(n9806) );
  INV_X1 U10558 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9097) );
  MUX2_X1 U10559 ( .A(n9097), .B(P1_REG1_REG_13__SCAN_IN), .S(n9753), .Z(n9760) );
  OR2_X1 U10560 ( .A1(n9737), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9102) );
  INV_X1 U10561 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9098) );
  MUX2_X1 U10562 ( .A(n9098), .B(P1_REG1_REG_10__SCAN_IN), .S(n9575), .Z(n9568) );
  OAI21_X1 U10563 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9122), .A(n9099), .ZN(
        n9569) );
  NOR2_X1 U10564 ( .A1(n9568), .A2(n9569), .ZN(n9567) );
  AOI21_X1 U10565 ( .B1(n9575), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9567), .ZN(
        n9727) );
  INV_X1 U10566 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9100) );
  MUX2_X1 U10567 ( .A(n9100), .B(P1_REG1_REG_11__SCAN_IN), .S(n9124), .Z(n9728) );
  NOR2_X1 U10568 ( .A1(n9727), .A2(n9728), .ZN(n9726) );
  AOI21_X1 U10569 ( .B1(n9124), .B2(P1_REG1_REG_11__SCAN_IN), .A(n9726), .ZN(
        n9743) );
  INV_X1 U10570 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9101) );
  MUX2_X1 U10571 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9101), .S(n9737), .Z(n9744) );
  NAND2_X1 U10572 ( .A1(n9743), .A2(n9744), .ZN(n9742) );
  NAND2_X1 U10573 ( .A1(n9102), .A2(n9742), .ZN(n9759) );
  NOR2_X1 U10574 ( .A1(n9760), .A2(n9759), .ZN(n9758) );
  AOI21_X1 U10575 ( .B1(n9753), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9758), .ZN(
        n9775) );
  INV_X1 U10576 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9103) );
  OR2_X1 U10577 ( .A1(n9126), .A2(n9103), .ZN(n9105) );
  NAND2_X1 U10578 ( .A1(n9126), .A2(n9103), .ZN(n9104) );
  AND2_X1 U10579 ( .A1(n9105), .A2(n9104), .ZN(n9774) );
  NOR2_X1 U10580 ( .A1(n9775), .A2(n9774), .ZN(n9773) );
  AOI21_X1 U10581 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9126), .A(n9773), .ZN(
        n9106) );
  NOR2_X1 U10582 ( .A1(n9106), .A2(n9128), .ZN(n9107) );
  INV_X1 U10583 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9786) );
  XNOR2_X1 U10584 ( .A(n9128), .B(n9106), .ZN(n9787) );
  NOR2_X1 U10585 ( .A1(n9786), .A2(n9787), .ZN(n9785) );
  NOR2_X1 U10586 ( .A1(n9107), .A2(n9785), .ZN(n9805) );
  NAND2_X1 U10587 ( .A1(n9806), .A2(n9805), .ZN(n9804) );
  OAI21_X1 U10588 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n9807), .A(n9804), .ZN(
        n9816) );
  NAND2_X1 U10589 ( .A1(n9815), .A2(n9816), .ZN(n9814) );
  AND2_X1 U10590 ( .A1(n9108), .A2(n9814), .ZN(n9831) );
  NAND2_X1 U10591 ( .A1(n9114), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9111) );
  INV_X1 U10592 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9109) );
  NAND2_X1 U10593 ( .A1(n9834), .A2(n9109), .ZN(n9110) );
  AND2_X1 U10594 ( .A1(n9111), .A2(n9110), .ZN(n9830) );
  NAND2_X1 U10595 ( .A1(n9831), .A2(n9830), .ZN(n9828) );
  NAND2_X1 U10596 ( .A1(n9828), .A2(n9111), .ZN(n9113) );
  INV_X1 U10597 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9112) );
  NAND2_X1 U10598 ( .A1(n9114), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9132) );
  INV_X1 U10599 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9115) );
  NAND2_X1 U10600 ( .A1(n9834), .A2(n9115), .ZN(n9116) );
  AND2_X1 U10601 ( .A1(n9132), .A2(n9116), .ZN(n9827) );
  NOR2_X1 U10602 ( .A1(n9819), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9117) );
  AOI21_X1 U10603 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n9819), .A(n9117), .ZN(
        n9812) );
  NAND2_X1 U10604 ( .A1(n9753), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9118) );
  OAI21_X1 U10605 ( .B1(n9753), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9118), .ZN(
        n9756) );
  NOR2_X1 U10606 ( .A1(n9737), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n9119) );
  AOI21_X1 U10607 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9737), .A(n9119), .ZN(
        n9740) );
  NAND2_X1 U10608 ( .A1(n9575), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9120) );
  OAI21_X1 U10609 ( .B1(n9575), .B2(P1_REG2_REG_10__SCAN_IN), .A(n9120), .ZN(
        n9571) );
  OAI21_X1 U10610 ( .B1(n9122), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9121), .ZN(
        n9572) );
  NOR2_X1 U10611 ( .A1(n9571), .A2(n9572), .ZN(n9570) );
  AOI22_X1 U10612 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n9732), .B1(n9124), .B2(
        n9123), .ZN(n9724) );
  OAI21_X1 U10613 ( .B1(n9737), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9738), .ZN(
        n9755) );
  NOR2_X1 U10614 ( .A1(n9756), .A2(n9755), .ZN(n9754) );
  NAND2_X1 U10615 ( .A1(n9126), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9125) );
  OAI21_X1 U10616 ( .B1(n9126), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9125), .ZN(
        n9771) );
  NOR2_X1 U10617 ( .A1(n9127), .A2(n9128), .ZN(n9129) );
  INV_X1 U10618 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9789) );
  NOR2_X1 U10619 ( .A1(n9789), .A2(n9790), .ZN(n9788) );
  NOR2_X1 U10620 ( .A1(n9129), .A2(n9788), .ZN(n9800) );
  AOI22_X1 U10621 ( .A1(n9807), .A2(n9131), .B1(P1_REG2_REG_16__SCAN_IN), .B2(
        n9130), .ZN(n9799) );
  NOR2_X1 U10622 ( .A1(n9800), .A2(n9799), .ZN(n9798) );
  NAND2_X1 U10623 ( .A1(n9827), .A2(n9826), .ZN(n9824) );
  NAND2_X1 U10624 ( .A1(n9824), .A2(n9132), .ZN(n9133) );
  XNOR2_X1 U10625 ( .A(n9133), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9135) );
  INV_X1 U10626 ( .A(n9835), .ZN(n9818) );
  AOI21_X1 U10627 ( .B1(n9825), .B2(n9135), .A(n9818), .ZN(n9134) );
  OAI22_X1 U10628 ( .A1(n9135), .A2(n9797), .B1(n9784), .B2(n4470), .ZN(n9136)
         );
  INV_X1 U10629 ( .A(n9478), .ZN(n9281) );
  OR2_X2 U10630 ( .A1(n9390), .A2(n9385), .ZN(n9391) );
  OR2_X2 U10631 ( .A1(n9391), .A2(n9514), .ZN(n9372) );
  OR2_X2 U10632 ( .A1(n9372), .A2(n9507), .ZN(n9353) );
  NOR2_X2 U10633 ( .A1(n9500), .A2(n9353), .ZN(n9335) );
  OR2_X2 U10634 ( .A1(n9276), .A2(n9259), .ZN(n9257) );
  OR2_X2 U10635 ( .A1(n9244), .A2(n9257), .ZN(n9242) );
  NOR2_X2 U10636 ( .A1(n9228), .A2(n9242), .ZN(n9227) );
  NAND2_X1 U10637 ( .A1(n9137), .A2(n9900), .ZN(n9436) );
  NAND2_X1 U10638 ( .A1(n9907), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9141) );
  NOR2_X1 U10639 ( .A1(n4459), .A2(n9138), .ZN(n9139) );
  NOR2_X1 U10640 ( .A1(n9881), .A2(n9139), .ZN(n9197) );
  NAND2_X1 U10641 ( .A1(n9140), .A2(n9197), .ZN(n9438) );
  OR2_X1 U10642 ( .A1(n9907), .A2(n9438), .ZN(n9145) );
  OAI211_X1 U10643 ( .C1(n9437), .C2(n9896), .A(n9141), .B(n9145), .ZN(n9142)
         );
  INV_X1 U10644 ( .A(n9142), .ZN(n9143) );
  OAI21_X1 U10645 ( .B1(n9436), .B2(n9380), .A(n9143), .ZN(P1_U3263) );
  OAI211_X1 U10646 ( .C1(n9201), .C2(n9440), .A(n9900), .B(n9144), .ZN(n9439)
         );
  INV_X1 U10647 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9146) );
  OAI21_X1 U10648 ( .B1(n9238), .B2(n9146), .A(n9145), .ZN(n9147) );
  AOI21_X1 U10649 ( .B1(n9148), .B2(n9854), .A(n9147), .ZN(n9149) );
  OAI21_X1 U10650 ( .B1(n9439), .B2(n9380), .A(n9149), .ZN(P1_U3264) );
  NAND2_X1 U10651 ( .A1(n9426), .A2(n9409), .ZN(n9153) );
  OAI21_X1 U10652 ( .B1(n9376), .B2(n4738), .A(n9384), .ZN(n9155) );
  INV_X1 U10653 ( .A(n9514), .ZN(n9156) );
  NAND2_X1 U10654 ( .A1(n9301), .A2(n5038), .ZN(n9165) );
  NAND2_X1 U10655 ( .A1(n9165), .A2(n9164), .ZN(n9284) );
  INV_X1 U10656 ( .A(n9284), .ZN(n9169) );
  INV_X1 U10657 ( .A(n9299), .ZN(n9482) );
  NOR2_X1 U10658 ( .A1(n9478), .A2(n9170), .ZN(n9171) );
  NAND2_X1 U10659 ( .A1(n9470), .A2(n9462), .ZN(n9172) );
  NAND2_X1 U10660 ( .A1(n9226), .A2(n9234), .ZN(n9178) );
  INV_X1 U10661 ( .A(n9228), .ZN(n9456) );
  NAND2_X1 U10662 ( .A1(n9456), .A2(n9252), .ZN(n9177) );
  XNOR2_X1 U10663 ( .A(n9179), .B(n9195), .ZN(n9441) );
  INV_X1 U10664 ( .A(n9441), .ZN(n9208) );
  INV_X1 U10665 ( .A(n9180), .ZN(n9311) );
  INV_X1 U10666 ( .A(n9181), .ZN(n9310) );
  NOR2_X1 U10667 ( .A1(n9265), .A2(n9266), .ZN(n9264) );
  XOR2_X1 U10668 ( .A(n9195), .B(n9194), .Z(n9200) );
  AOI22_X1 U10669 ( .A1(n9198), .A2(n9996), .B1(n9197), .B2(n9196), .ZN(n9199)
         );
  OAI21_X1 U10670 ( .B1(n9200), .B2(n9420), .A(n9199), .ZN(n9445) );
  AOI211_X1 U10671 ( .C1(n9442), .C2(n9216), .A(n9944), .B(n9201), .ZN(n9444)
         );
  NAND2_X1 U10672 ( .A1(n9444), .A2(n9903), .ZN(n9204) );
  AOI22_X1 U10673 ( .A1(n9907), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9852), .B2(
        n9202), .ZN(n9203) );
  OAI211_X1 U10674 ( .C1(n9205), .C2(n9896), .A(n9204), .B(n9203), .ZN(n9206)
         );
  AOI21_X1 U10675 ( .B1(n9445), .B2(n9238), .A(n9206), .ZN(n9207) );
  OAI21_X1 U10676 ( .B1(n9208), .B2(n9415), .A(n9207), .ZN(P1_U3356) );
  XNOR2_X1 U10677 ( .A(n9209), .B(n9213), .ZN(n9211) );
  AOI22_X1 U10678 ( .A1(n9211), .A2(n9890), .B1(n9864), .B2(n9210), .ZN(n9453)
         );
  NAND2_X1 U10679 ( .A1(n9212), .A2(n4731), .ZN(n9214) );
  OAI211_X1 U10680 ( .C1(n9217), .C2(n9227), .A(n9900), .B(n9216), .ZN(n9451)
         );
  NOR2_X1 U10681 ( .A1(n9893), .A2(n9218), .ZN(n9219) );
  AOI21_X1 U10682 ( .B1(n9907), .B2(P1_REG2_REG_28__SCAN_IN), .A(n9219), .ZN(
        n9220) );
  OAI21_X1 U10683 ( .B1(n9377), .B2(n9252), .A(n9220), .ZN(n9221) );
  AOI21_X1 U10684 ( .B1(n9450), .B2(n9854), .A(n9221), .ZN(n9222) );
  OAI21_X1 U10685 ( .B1(n9451), .B2(n9223), .A(n9222), .ZN(n9224) );
  AOI21_X1 U10686 ( .B1(n9448), .B2(n9877), .A(n9224), .ZN(n9225) );
  OAI21_X1 U10687 ( .B1(n9907), .B2(n9453), .A(n9225), .ZN(P1_U3265) );
  XOR2_X1 U10688 ( .A(n9234), .B(n9226), .Z(n9461) );
  AOI211_X1 U10689 ( .C1(n9228), .C2(n9242), .A(n9944), .B(n9227), .ZN(n9458)
         );
  NAND2_X1 U10690 ( .A1(n9228), .A2(n9854), .ZN(n9231) );
  AOI22_X1 U10691 ( .A1(n9907), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9229), .B2(
        n9852), .ZN(n9230) );
  OAI211_X1 U10692 ( .C1(n9455), .C2(n9377), .A(n9231), .B(n9230), .ZN(n9232)
         );
  AOI21_X1 U10693 ( .B1(n9458), .B2(n9903), .A(n9232), .ZN(n9240) );
  AOI21_X1 U10694 ( .B1(n9235), .B2(n9234), .A(n9233), .ZN(n9237) );
  OAI22_X1 U10695 ( .A1(n9237), .A2(n9420), .B1(n9236), .B2(n9881), .ZN(n9459)
         );
  NAND2_X1 U10696 ( .A1(n9459), .A2(n9238), .ZN(n9239) );
  OAI211_X1 U10697 ( .C1(n9461), .C2(n9415), .A(n9240), .B(n9239), .ZN(
        P1_U3266) );
  XNOR2_X1 U10698 ( .A(n9241), .B(n9250), .ZN(n9468) );
  INV_X1 U10699 ( .A(n9242), .ZN(n9243) );
  AOI211_X1 U10700 ( .C1(n9244), .C2(n9257), .A(n9944), .B(n9243), .ZN(n9465)
         );
  NAND2_X1 U10701 ( .A1(n9244), .A2(n9854), .ZN(n9247) );
  AOI22_X1 U10702 ( .A1(n9907), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9245), .B2(
        n9852), .ZN(n9246) );
  OAI211_X1 U10703 ( .C1(n9462), .C2(n9377), .A(n9247), .B(n9246), .ZN(n9248)
         );
  AOI21_X1 U10704 ( .B1(n9465), .B2(n9413), .A(n9248), .ZN(n9255) );
  AOI21_X1 U10705 ( .B1(n9251), .B2(n9250), .A(n9249), .ZN(n9253) );
  OAI22_X1 U10706 ( .A1(n9253), .A2(n9420), .B1(n9252), .B2(n9881), .ZN(n9466)
         );
  NAND2_X1 U10707 ( .A1(n9466), .A2(n9238), .ZN(n9254) );
  OAI211_X1 U10708 ( .C1(n9468), .C2(n9415), .A(n9255), .B(n9254), .ZN(
        P1_U3267) );
  XNOR2_X1 U10709 ( .A(n9256), .B(n9266), .ZN(n9475) );
  INV_X1 U10710 ( .A(n9257), .ZN(n9258) );
  AOI211_X1 U10711 ( .C1(n9259), .C2(n9276), .A(n9944), .B(n9258), .ZN(n9472)
         );
  NAND2_X1 U10712 ( .A1(n9259), .A2(n9854), .ZN(n9262) );
  AOI22_X1 U10713 ( .A1(n9907), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9260), .B2(
        n9852), .ZN(n9261) );
  OAI211_X1 U10714 ( .C1(n9469), .C2(n9377), .A(n9262), .B(n9261), .ZN(n9263)
         );
  AOI21_X1 U10715 ( .B1(n9472), .B2(n9903), .A(n9263), .ZN(n9269) );
  AOI21_X1 U10716 ( .B1(n9266), .B2(n9265), .A(n9264), .ZN(n9267) );
  OAI22_X1 U10717 ( .A1(n9267), .A2(n9420), .B1(n9455), .B2(n9881), .ZN(n9473)
         );
  NAND2_X1 U10718 ( .A1(n9473), .A2(n9238), .ZN(n9268) );
  OAI211_X1 U10719 ( .C1(n9475), .C2(n9415), .A(n9269), .B(n9268), .ZN(
        P1_U3268) );
  XNOR2_X1 U10720 ( .A(n9270), .B(n9272), .ZN(n9480) );
  OAI211_X1 U10721 ( .C1(n9273), .C2(n9272), .A(n9271), .B(n9890), .ZN(n9275)
         );
  OR2_X1 U10722 ( .A1(n9462), .A2(n9881), .ZN(n9274) );
  OAI211_X1 U10723 ( .C1(n9315), .C2(n9883), .A(n9275), .B(n9274), .ZN(n9476)
         );
  INV_X1 U10724 ( .A(n9276), .ZN(n9277) );
  AOI211_X1 U10725 ( .C1(n9478), .C2(n4937), .A(n9944), .B(n9277), .ZN(n9477)
         );
  NAND2_X1 U10726 ( .A1(n9477), .A2(n9903), .ZN(n9280) );
  AOI22_X1 U10727 ( .A1(n9907), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9278), .B2(
        n9852), .ZN(n9279) );
  OAI211_X1 U10728 ( .C1(n9281), .C2(n9896), .A(n9280), .B(n9279), .ZN(n9282)
         );
  AOI21_X1 U10729 ( .B1(n9476), .B2(n9238), .A(n9282), .ZN(n9283) );
  OAI21_X1 U10730 ( .B1(n9480), .B2(n9415), .A(n9283), .ZN(P1_U3269) );
  XOR2_X1 U10731 ( .A(n9284), .B(n9290), .Z(n9487) );
  INV_X1 U10732 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9285) );
  OAI22_X1 U10733 ( .A1(n9481), .A2(n9377), .B1(n9285), .B2(n9238), .ZN(n9298)
         );
  INV_X1 U10734 ( .A(n9286), .ZN(n9313) );
  NAND2_X1 U10735 ( .A1(n9313), .A2(n9287), .ZN(n9289) );
  AOI21_X1 U10736 ( .B1(n9290), .B2(n9289), .A(n9288), .ZN(n9291) );
  OAI22_X1 U10737 ( .A1(n9291), .A2(n9420), .B1(n9469), .B2(n9881), .ZN(n9485)
         );
  INV_X1 U10738 ( .A(n9485), .ZN(n9296) );
  AOI211_X1 U10739 ( .C1(n9299), .C2(n9302), .A(n9944), .B(n9292), .ZN(n9484)
         );
  AOI22_X1 U10740 ( .A1(n9484), .A2(n9294), .B1(n9852), .B2(n9293), .ZN(n9295)
         );
  AOI21_X1 U10741 ( .B1(n9296), .B2(n9295), .A(n9851), .ZN(n9297) );
  AOI211_X1 U10742 ( .C1(n9854), .C2(n9299), .A(n9298), .B(n9297), .ZN(n9300)
         );
  OAI21_X1 U10743 ( .B1(n9487), .B2(n9415), .A(n9300), .ZN(P1_U3270) );
  XOR2_X1 U10744 ( .A(n9301), .B(n9309), .Z(n9494) );
  INV_X1 U10745 ( .A(n9302), .ZN(n9303) );
  AOI211_X1 U10746 ( .C1(n9304), .C2(n9326), .A(n9944), .B(n9303), .ZN(n9491)
         );
  NAND2_X1 U10747 ( .A1(n9304), .A2(n9854), .ZN(n9307) );
  AOI22_X1 U10748 ( .A1(n9305), .A2(n9852), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9851), .ZN(n9306) );
  OAI211_X1 U10749 ( .C1(n9488), .C2(n9377), .A(n9307), .B(n9306), .ZN(n9308)
         );
  AOI21_X1 U10750 ( .B1(n9491), .B2(n9903), .A(n9308), .ZN(n9317) );
  OAI21_X1 U10751 ( .B1(n9311), .B2(n9310), .A(n9309), .ZN(n9312) );
  NAND3_X1 U10752 ( .A1(n9313), .A2(n9890), .A3(n9312), .ZN(n9314) );
  OAI21_X1 U10753 ( .B1(n9315), .B2(n9881), .A(n9314), .ZN(n9492) );
  NAND2_X1 U10754 ( .A1(n9492), .A2(n9238), .ZN(n9316) );
  OAI211_X1 U10755 ( .C1(n9494), .C2(n9415), .A(n9317), .B(n9316), .ZN(
        P1_U3271) );
  XOR2_X1 U10756 ( .A(n9321), .B(n9318), .Z(n9499) );
  NAND2_X1 U10757 ( .A1(n9320), .A2(n9319), .ZN(n9322) );
  XNOR2_X1 U10758 ( .A(n9322), .B(n9321), .ZN(n9323) );
  OAI222_X1 U10759 ( .A1(n9881), .A2(n9481), .B1(n9883), .B2(n9324), .C1(n9323), .C2(n9420), .ZN(n9495) );
  OR2_X1 U10760 ( .A1(n9331), .A2(n9335), .ZN(n9325) );
  AND3_X1 U10761 ( .A1(n9326), .A2(n9325), .A3(n9900), .ZN(n9496) );
  NAND2_X1 U10762 ( .A1(n9496), .A2(n9903), .ZN(n9330) );
  INV_X1 U10763 ( .A(n9327), .ZN(n9328) );
  AOI22_X1 U10764 ( .A1(n9328), .A2(n9852), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9851), .ZN(n9329) );
  OAI211_X1 U10765 ( .C1(n9331), .C2(n9896), .A(n9330), .B(n9329), .ZN(n9332)
         );
  AOI21_X1 U10766 ( .B1(n9495), .B2(n9238), .A(n9332), .ZN(n9333) );
  OAI21_X1 U10767 ( .B1(n9499), .B2(n9415), .A(n9333), .ZN(P1_U3272) );
  XOR2_X1 U10768 ( .A(n9341), .B(n9334), .Z(n9504) );
  AOI21_X1 U10769 ( .B1(n9500), .B2(n9353), .A(n9335), .ZN(n9501) );
  INV_X1 U10770 ( .A(n9336), .ZN(n9337) );
  AOI22_X1 U10771 ( .A1(n9851), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9337), .B2(
        n9852), .ZN(n9338) );
  OAI21_X1 U10772 ( .B1(n9339), .B2(n9896), .A(n9338), .ZN(n9345) );
  XOR2_X1 U10773 ( .A(n9341), .B(n9340), .Z(n9343) );
  AOI222_X1 U10774 ( .A1(n9890), .A2(n9343), .B1(n9342), .B2(n9864), .C1(n9369), .C2(n9996), .ZN(n9503) );
  NOR2_X1 U10775 ( .A1(n9503), .A2(n9851), .ZN(n9344) );
  AOI211_X1 U10776 ( .C1(n9501), .C2(n9431), .A(n9345), .B(n9344), .ZN(n9346)
         );
  OAI21_X1 U10777 ( .B1(n9504), .B2(n9415), .A(n9346), .ZN(P1_U3273) );
  XNOR2_X1 U10778 ( .A(n9348), .B(n9347), .ZN(n9505) );
  XNOR2_X1 U10779 ( .A(n9350), .B(n9349), .ZN(n9352) );
  AOI22_X1 U10780 ( .A1(n9352), .A2(n9890), .B1(n9864), .B2(n9351), .ZN(n9510)
         );
  NOR2_X1 U10781 ( .A1(n9510), .A2(n9851), .ZN(n9362) );
  AOI21_X1 U10782 ( .B1(n9507), .B2(n9372), .A(n9944), .ZN(n9354) );
  NAND2_X1 U10783 ( .A1(n9354), .A2(n9353), .ZN(n9508) );
  NOR2_X1 U10784 ( .A1(n9355), .A2(n9893), .ZN(n9356) );
  AOI21_X1 U10785 ( .B1(n9907), .B2(P1_REG2_REG_19__SCAN_IN), .A(n9356), .ZN(
        n9357) );
  OAI21_X1 U10786 ( .B1(n9377), .B2(n9358), .A(n9357), .ZN(n9359) );
  AOI21_X1 U10787 ( .B1(n9507), .B2(n9854), .A(n9359), .ZN(n9360) );
  OAI21_X1 U10788 ( .B1(n9508), .B2(n9380), .A(n9360), .ZN(n9361) );
  AOI211_X1 U10789 ( .C1(n9505), .C2(n9877), .A(n9362), .B(n9361), .ZN(n9363)
         );
  INV_X1 U10790 ( .A(n9363), .ZN(P1_U3274) );
  XNOR2_X1 U10791 ( .A(n9365), .B(n9364), .ZN(n9512) );
  OAI21_X1 U10792 ( .B1(n9368), .B2(n9367), .A(n9366), .ZN(n9370) );
  AOI22_X1 U10793 ( .A1(n9370), .A2(n9890), .B1(n9864), .B2(n9369), .ZN(n9517)
         );
  NOR2_X1 U10794 ( .A1(n9517), .A2(n9907), .ZN(n9382) );
  NAND2_X1 U10795 ( .A1(n9391), .A2(n9514), .ZN(n9371) );
  NAND3_X1 U10796 ( .A1(n9372), .A2(n9900), .A3(n9371), .ZN(n9515) );
  NOR2_X1 U10797 ( .A1(n9893), .A2(n9373), .ZN(n9374) );
  AOI21_X1 U10798 ( .B1(n9907), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9374), .ZN(
        n9375) );
  OAI21_X1 U10799 ( .B1(n9377), .B2(n9376), .A(n9375), .ZN(n9378) );
  AOI21_X1 U10800 ( .B1(n9514), .B2(n9854), .A(n9378), .ZN(n9379) );
  OAI21_X1 U10801 ( .B1(n9515), .B2(n9380), .A(n9379), .ZN(n9381) );
  AOI211_X1 U10802 ( .C1(n9512), .C2(n9877), .A(n9382), .B(n9381), .ZN(n9383)
         );
  INV_X1 U10803 ( .A(n9383), .ZN(P1_U3275) );
  XNOR2_X1 U10804 ( .A(n9384), .B(n9386), .ZN(n9646) );
  INV_X1 U10805 ( .A(n9646), .ZN(n9399) );
  AOI22_X1 U10806 ( .A1(n9385), .A2(n9854), .B1(P1_REG2_REG_17__SCAN_IN), .B2(
        n9851), .ZN(n9398) );
  XOR2_X1 U10807 ( .A(n9387), .B(n9386), .Z(n9389) );
  AOI222_X1 U10808 ( .A1(n9890), .A2(n9389), .B1(n9506), .B2(n9864), .C1(n9388), .C2(n9996), .ZN(n9644) );
  INV_X1 U10809 ( .A(n9644), .ZN(n9396) );
  INV_X1 U10810 ( .A(n9390), .ZN(n9402) );
  OAI211_X1 U10811 ( .C1(n9402), .C2(n4738), .A(n9900), .B(n9391), .ZN(n9643)
         );
  INV_X1 U10812 ( .A(n9392), .ZN(n9393) );
  OAI22_X1 U10813 ( .A1(n9643), .A2(n4722), .B1(n9893), .B2(n9393), .ZN(n9395)
         );
  OAI21_X1 U10814 ( .B1(n9396), .B2(n9395), .A(n9238), .ZN(n9397) );
  OAI211_X1 U10815 ( .C1(n9399), .C2(n9415), .A(n9398), .B(n9397), .ZN(
        P1_U3276) );
  XNOR2_X1 U10816 ( .A(n9401), .B(n9400), .ZN(n9523) );
  AOI211_X1 U10817 ( .C1(n9520), .C2(n4952), .A(n9944), .B(n9402), .ZN(n9519)
         );
  AOI22_X1 U10818 ( .A1(n9851), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9403), .B2(
        n9852), .ZN(n9404) );
  OAI21_X1 U10819 ( .B1(n9405), .B2(n9896), .A(n9404), .ZN(n9412) );
  OAI21_X1 U10820 ( .B1(n9408), .B2(n9407), .A(n9406), .ZN(n9410) );
  AOI222_X1 U10821 ( .A1(n9890), .A2(n9410), .B1(n9513), .B2(n9864), .C1(n9409), .C2(n9996), .ZN(n9522) );
  NOR2_X1 U10822 ( .A1(n9522), .A2(n9851), .ZN(n9411) );
  AOI211_X1 U10823 ( .C1(n9519), .C2(n9413), .A(n9412), .B(n9411), .ZN(n9414)
         );
  OAI21_X1 U10824 ( .B1(n9415), .B2(n9523), .A(n9414), .ZN(P1_U3277) );
  INV_X1 U10825 ( .A(n9416), .ZN(n9417) );
  AOI21_X1 U10826 ( .B1(n9424), .B2(n9418), .A(n9417), .ZN(n9419) );
  OAI222_X1 U10827 ( .A1(n9883), .A2(n9422), .B1(n9881), .B2(n9421), .C1(n9420), .C2(n9419), .ZN(n9650) );
  AOI21_X1 U10828 ( .B1(n9423), .B2(n9852), .A(n9650), .ZN(n9435) );
  XOR2_X1 U10829 ( .A(n9425), .B(n9424), .Z(n9651) );
  NAND2_X1 U10830 ( .A1(n9651), .A2(n9877), .ZN(n9434) );
  AND2_X1 U10831 ( .A1(n9427), .A2(n9426), .ZN(n9429) );
  OR2_X1 U10832 ( .A1(n9429), .A2(n9428), .ZN(n9648) );
  INV_X1 U10833 ( .A(n9648), .ZN(n9432) );
  OAI22_X1 U10834 ( .A1(n4950), .A2(n9896), .B1(n9789), .B2(n9238), .ZN(n9430)
         );
  AOI21_X1 U10835 ( .B1(n9432), .B2(n9431), .A(n9430), .ZN(n9433) );
  OAI211_X1 U10836 ( .C1(n9907), .C2(n9435), .A(n9434), .B(n9433), .ZN(
        P1_U3278) );
  OAI211_X1 U10837 ( .C1(n9437), .C2(n10007), .A(n9436), .B(n9438), .ZN(n9530)
         );
  MUX2_X1 U10838 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9530), .S(n10033), .Z(
        P1_U3553) );
  OAI211_X1 U10839 ( .C1(n9440), .C2(n10007), .A(n9439), .B(n9438), .ZN(n9531)
         );
  MUX2_X1 U10840 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9531), .S(n10033), .Z(
        P1_U3552) );
  NAND2_X1 U10841 ( .A1(n9441), .A2(n10009), .ZN(n9447) );
  NAND2_X1 U10842 ( .A1(n9447), .A2(n9446), .ZN(n9532) );
  MUX2_X1 U10843 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9532), .S(n10033), .Z(
        P1_U3551) );
  NAND2_X1 U10844 ( .A1(n9448), .A2(n10009), .ZN(n9454) );
  AOI22_X1 U10845 ( .A1(n9450), .A2(n9997), .B1(n9996), .B2(n9449), .ZN(n9452)
         );
  NAND4_X1 U10846 ( .A1(n9454), .A2(n9453), .A3(n9452), .A4(n9451), .ZN(n9533)
         );
  MUX2_X1 U10847 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9533), .S(n10033), .Z(
        P1_U3550) );
  OAI22_X1 U10848 ( .A1(n9456), .A2(n10007), .B1(n9455), .B2(n9883), .ZN(n9457) );
  NOR3_X1 U10849 ( .A1(n9459), .A2(n9458), .A3(n9457), .ZN(n9460) );
  OAI21_X1 U10850 ( .B1(n9461), .B2(n9528), .A(n9460), .ZN(n9534) );
  MUX2_X1 U10851 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9534), .S(n10033), .Z(
        P1_U3549) );
  OAI22_X1 U10852 ( .A1(n9463), .A2(n10007), .B1(n9462), .B2(n9883), .ZN(n9464) );
  NOR3_X1 U10853 ( .A1(n9466), .A2(n9465), .A3(n9464), .ZN(n9467) );
  OAI21_X1 U10854 ( .B1(n9468), .B2(n9528), .A(n9467), .ZN(n9535) );
  MUX2_X1 U10855 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9535), .S(n10033), .Z(
        P1_U3548) );
  OAI22_X1 U10856 ( .A1(n9470), .A2(n10007), .B1(n9469), .B2(n9883), .ZN(n9471) );
  NOR3_X1 U10857 ( .A1(n9473), .A2(n9472), .A3(n9471), .ZN(n9474) );
  OAI21_X1 U10858 ( .B1(n9475), .B2(n9528), .A(n9474), .ZN(n9536) );
  MUX2_X1 U10859 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9536), .S(n10033), .Z(
        P1_U3547) );
  AOI211_X1 U10860 ( .C1(n9997), .C2(n9478), .A(n9477), .B(n9476), .ZN(n9479)
         );
  OAI21_X1 U10861 ( .B1(n9480), .B2(n9528), .A(n9479), .ZN(n9537) );
  MUX2_X1 U10862 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9537), .S(n10033), .Z(
        P1_U3546) );
  OAI22_X1 U10863 ( .A1(n9482), .A2(n10007), .B1(n9481), .B2(n9883), .ZN(n9483) );
  NOR3_X1 U10864 ( .A1(n9485), .A2(n9484), .A3(n9483), .ZN(n9486) );
  OAI21_X1 U10865 ( .B1(n9487), .B2(n9528), .A(n9486), .ZN(n9538) );
  MUX2_X1 U10866 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9538), .S(n10033), .Z(
        P1_U3545) );
  OAI22_X1 U10867 ( .A1(n9489), .A2(n10007), .B1(n9488), .B2(n9883), .ZN(n9490) );
  NOR3_X1 U10868 ( .A1(n9492), .A2(n9491), .A3(n9490), .ZN(n9493) );
  OAI21_X1 U10869 ( .B1(n9494), .B2(n9528), .A(n9493), .ZN(n9539) );
  MUX2_X1 U10870 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9539), .S(n10033), .Z(
        P1_U3544) );
  AOI211_X1 U10871 ( .C1(n9997), .C2(n9497), .A(n9496), .B(n9495), .ZN(n9498)
         );
  OAI21_X1 U10872 ( .B1(n9499), .B2(n9528), .A(n9498), .ZN(n9540) );
  MUX2_X1 U10873 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9540), .S(n10033), .Z(
        P1_U3543) );
  AOI22_X1 U10874 ( .A1(n9501), .A2(n9900), .B1(n9997), .B2(n9500), .ZN(n9502)
         );
  OAI211_X1 U10875 ( .C1(n9504), .C2(n9528), .A(n9503), .B(n9502), .ZN(n9541)
         );
  MUX2_X1 U10876 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9541), .S(n10033), .Z(
        P1_U3542) );
  NAND2_X1 U10877 ( .A1(n9505), .A2(n10009), .ZN(n9511) );
  AOI22_X1 U10878 ( .A1(n9507), .A2(n9997), .B1(n9996), .B2(n9506), .ZN(n9509)
         );
  NAND4_X1 U10879 ( .A1(n9511), .A2(n9510), .A3(n9509), .A4(n9508), .ZN(n9542)
         );
  MUX2_X1 U10880 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9542), .S(n10033), .Z(
        P1_U3541) );
  NAND2_X1 U10881 ( .A1(n9512), .A2(n10009), .ZN(n9518) );
  AOI22_X1 U10882 ( .A1(n9514), .A2(n9997), .B1(n9996), .B2(n9513), .ZN(n9516)
         );
  NAND4_X1 U10883 ( .A1(n9518), .A2(n9517), .A3(n9516), .A4(n9515), .ZN(n9543)
         );
  MUX2_X1 U10884 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9543), .S(n10033), .Z(
        P1_U3540) );
  AOI21_X1 U10885 ( .B1(n9997), .B2(n9520), .A(n9519), .ZN(n9521) );
  OAI211_X1 U10886 ( .C1(n9523), .C2(n9528), .A(n9522), .B(n9521), .ZN(n9544)
         );
  MUX2_X1 U10887 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9544), .S(n10033), .Z(
        P1_U3538) );
  AOI22_X1 U10888 ( .A1(n9525), .A2(n9900), .B1(n9997), .B2(n9524), .ZN(n9526)
         );
  OAI211_X1 U10889 ( .C1(n9529), .C2(n9528), .A(n9527), .B(n9526), .ZN(n9545)
         );
  MUX2_X1 U10890 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9545), .S(n10033), .Z(
        P1_U3536) );
  MUX2_X1 U10891 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9530), .S(n10013), .Z(
        P1_U3521) );
  MUX2_X1 U10892 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9531), .S(n10013), .Z(
        P1_U3520) );
  MUX2_X1 U10893 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9532), .S(n10013), .Z(
        P1_U3519) );
  MUX2_X1 U10894 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9533), .S(n10013), .Z(
        P1_U3518) );
  MUX2_X1 U10895 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9534), .S(n10013), .Z(
        P1_U3517) );
  MUX2_X1 U10896 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9535), .S(n10013), .Z(
        P1_U3516) );
  MUX2_X1 U10897 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9536), .S(n10013), .Z(
        P1_U3515) );
  MUX2_X1 U10898 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9537), .S(n10013), .Z(
        P1_U3514) );
  MUX2_X1 U10899 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9538), .S(n10013), .Z(
        P1_U3513) );
  MUX2_X1 U10900 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9539), .S(n10013), .Z(
        P1_U3512) );
  MUX2_X1 U10901 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9540), .S(n10013), .Z(
        P1_U3511) );
  MUX2_X1 U10902 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9541), .S(n10013), .Z(
        P1_U3510) );
  MUX2_X1 U10903 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9542), .S(n10013), .Z(
        P1_U3509) );
  MUX2_X1 U10904 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9543), .S(n10013), .Z(
        P1_U3507) );
  MUX2_X1 U10905 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9544), .S(n10013), .Z(
        P1_U3501) );
  MUX2_X1 U10906 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9545), .S(n10013), .Z(
        P1_U3495) );
  MUX2_X1 U10907 ( .A(P1_D_REG_1__SCAN_IN), .B(n9548), .S(n9917), .Z(P1_U3440)
         );
  MUX2_X1 U10908 ( .A(P1_D_REG_0__SCAN_IN), .B(n9549), .S(n9917), .Z(P1_U3439)
         );
  NOR4_X1 U10909 ( .A1(n9551), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9550), .A4(
        n4454), .ZN(n9552) );
  AOI21_X1 U10910 ( .B1(n9553), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9552), .ZN(
        n9554) );
  OAI21_X1 U10911 ( .B1(n9555), .B2(n9565), .A(n9554), .ZN(P1_U3324) );
  OAI222_X1 U10912 ( .A1(n9562), .A2(n9558), .B1(n4454), .B2(n9557), .C1(n9556), .C2(n9565), .ZN(P1_U3326) );
  INV_X1 U10913 ( .A(n9559), .ZN(n9560) );
  OAI222_X1 U10914 ( .A1(n9562), .A2(n9561), .B1(n9565), .B2(n9560), .C1(n5882), .C2(n4454), .ZN(P1_U3327) );
  OAI222_X1 U10915 ( .A1(n9566), .A2(n4454), .B1(n9565), .B2(n9564), .C1(n9563), .C2(n9562), .ZN(P1_U3329) );
  INV_X1 U10916 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9578) );
  AOI211_X1 U10917 ( .C1(n9569), .C2(n9568), .A(n9567), .B(n9784), .ZN(n9574)
         );
  AOI211_X1 U10918 ( .C1(n9572), .C2(n9571), .A(n9570), .B(n9797), .ZN(n9573)
         );
  AOI211_X1 U10919 ( .C1(n9818), .C2(n9575), .A(n9574), .B(n9573), .ZN(n9577)
         );
  OAI211_X1 U10920 ( .C1(n9840), .C2(n9578), .A(n9577), .B(n9576), .ZN(
        P1_U3253) );
  INV_X1 U10921 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9593) );
  AOI21_X1 U10922 ( .B1(n9581), .B2(n9580), .A(n9579), .ZN(n9582) );
  NAND2_X1 U10923 ( .A1(n9825), .A2(n9582), .ZN(n9588) );
  AOI21_X1 U10924 ( .B1(n9585), .B2(n9584), .A(n9583), .ZN(n9586) );
  NAND2_X1 U10925 ( .A1(n9829), .A2(n9586), .ZN(n9587) );
  OAI211_X1 U10926 ( .C1(n9835), .C2(n9589), .A(n9588), .B(n9587), .ZN(n9590)
         );
  INV_X1 U10927 ( .A(n9590), .ZN(n9592) );
  OAI211_X1 U10928 ( .C1(n9840), .C2(n9593), .A(n9592), .B(n9591), .ZN(
        P1_U3250) );
  INV_X1 U10929 ( .A(n9594), .ZN(n9595) );
  OAI211_X1 U10930 ( .C1(n9597), .C2(n9596), .A(n9825), .B(n9595), .ZN(n9602)
         );
  OAI211_X1 U10931 ( .C1(n9600), .C2(n9599), .A(n9829), .B(n9598), .ZN(n9601)
         );
  OAI211_X1 U10932 ( .C1(n9835), .C2(n9603), .A(n9602), .B(n9601), .ZN(n9604)
         );
  INV_X1 U10933 ( .A(n9604), .ZN(n9606) );
  OAI211_X1 U10934 ( .C1(n9840), .C2(n9607), .A(n9606), .B(n9605), .ZN(
        P1_U3246) );
  INV_X1 U10935 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9622) );
  AOI21_X1 U10936 ( .B1(n9610), .B2(n9609), .A(n9608), .ZN(n9611) );
  NAND2_X1 U10937 ( .A1(n9825), .A2(n9611), .ZN(n9617) );
  AOI21_X1 U10938 ( .B1(n9614), .B2(n9613), .A(n9612), .ZN(n9615) );
  NAND2_X1 U10939 ( .A1(n9829), .A2(n9615), .ZN(n9616) );
  OAI211_X1 U10940 ( .C1(n9835), .C2(n9618), .A(n9617), .B(n9616), .ZN(n9619)
         );
  INV_X1 U10941 ( .A(n9619), .ZN(n9621) );
  OAI211_X1 U10942 ( .C1(n9840), .C2(n9622), .A(n9621), .B(n9620), .ZN(
        P1_U3251) );
  OAI22_X1 U10943 ( .A1(n9624), .A2(n10227), .B1(n9623), .B2(n10225), .ZN(
        n9625) );
  NOR2_X1 U10944 ( .A1(n9626), .A2(n9625), .ZN(n9638) );
  AOI22_X1 U10945 ( .A1(n10264), .A2(n9638), .B1(n9627), .B2(n10262), .ZN(
        P2_U3474) );
  NOR2_X1 U10946 ( .A1(n9628), .A2(n10227), .ZN(n9631) );
  INV_X1 U10947 ( .A(n9629), .ZN(n9630) );
  AOI211_X1 U10948 ( .C1(n10180), .C2(n9632), .A(n9631), .B(n9630), .ZN(n9640)
         );
  AOI22_X1 U10949 ( .A1(n10264), .A2(n9640), .B1(n8145), .B2(n10262), .ZN(
        P2_U3473) );
  AND2_X1 U10950 ( .A1(n9633), .A2(n10234), .ZN(n9635) );
  AOI211_X1 U10951 ( .C1(n10180), .C2(n9636), .A(n9635), .B(n9634), .ZN(n9642)
         );
  AOI22_X1 U10952 ( .A1(n10264), .A2(n9642), .B1(n4831), .B2(n10262), .ZN(
        P2_U3472) );
  INV_X1 U10953 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9637) );
  AOI22_X1 U10954 ( .A1(n10240), .A2(n9638), .B1(n9637), .B2(n10238), .ZN(
        P2_U3435) );
  INV_X1 U10955 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9639) );
  AOI22_X1 U10956 ( .A1(n10240), .A2(n9640), .B1(n9639), .B2(n10238), .ZN(
        P2_U3432) );
  INV_X1 U10957 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9641) );
  AOI22_X1 U10958 ( .A1(n10240), .A2(n9642), .B1(n9641), .B2(n10238), .ZN(
        P2_U3429) );
  OAI211_X1 U10959 ( .C1(n4738), .C2(n10007), .A(n9644), .B(n9643), .ZN(n9645)
         );
  AOI21_X1 U10960 ( .B1(n9646), .B2(n10009), .A(n9645), .ZN(n9653) );
  AOI22_X1 U10961 ( .A1(n10033), .A2(n9653), .B1(n9647), .B2(n10031), .ZN(
        P1_U3539) );
  OAI22_X1 U10962 ( .A1(n9648), .A2(n9944), .B1(n4950), .B2(n10007), .ZN(n9649) );
  AOI211_X1 U10963 ( .C1(n9651), .C2(n10009), .A(n9650), .B(n9649), .ZN(n9655)
         );
  AOI22_X1 U10964 ( .A1(n10033), .A2(n9655), .B1(n9786), .B2(n10031), .ZN(
        P1_U3537) );
  INV_X1 U10965 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9652) );
  AOI22_X1 U10966 ( .A1(n10013), .A2(n9653), .B1(n9652), .B2(n10011), .ZN(
        P1_U3504) );
  INV_X1 U10967 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9654) );
  AOI22_X1 U10968 ( .A1(n10013), .A2(n9655), .B1(n9654), .B2(n10011), .ZN(
        P1_U3498) );
  XNOR2_X1 U10969 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  AOI21_X1 U10970 ( .B1(n4459), .B2(n9657), .A(n9656), .ZN(n9658) );
  XNOR2_X1 U10971 ( .A(n9658), .B(P1_IR_REG_0__SCAN_IN), .ZN(n9661) );
  AOI22_X1 U10972 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9803), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n4454), .ZN(n9659) );
  OAI21_X1 U10973 ( .B1(n9661), .B2(n9660), .A(n9659), .ZN(P1_U3243) );
  AOI22_X1 U10974 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n9803), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9675) );
  AOI21_X1 U10975 ( .B1(n9664), .B2(n9663), .A(n9662), .ZN(n9665) );
  NAND2_X1 U10976 ( .A1(n9825), .A2(n9665), .ZN(n9671) );
  NAND2_X1 U10977 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9667) );
  AOI21_X1 U10978 ( .B1(n9668), .B2(n9667), .A(n9666), .ZN(n9669) );
  NAND2_X1 U10979 ( .A1(n9829), .A2(n9669), .ZN(n9670) );
  OAI211_X1 U10980 ( .C1(n9835), .C2(n9672), .A(n9671), .B(n9670), .ZN(n9673)
         );
  INV_X1 U10981 ( .A(n9673), .ZN(n9674) );
  NAND2_X1 U10982 ( .A1(n9675), .A2(n9674), .ZN(P1_U3244) );
  AOI21_X1 U10983 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(n9803), .A(n9676), .ZN(
        n9691) );
  AOI21_X1 U10984 ( .B1(n9679), .B2(n9678), .A(n9677), .ZN(n9680) );
  NAND2_X1 U10985 ( .A1(n9825), .A2(n9680), .ZN(n9686) );
  AOI21_X1 U10986 ( .B1(n9683), .B2(n9682), .A(n9681), .ZN(n9684) );
  NAND2_X1 U10987 ( .A1(n9829), .A2(n9684), .ZN(n9685) );
  OAI211_X1 U10988 ( .C1(n9687), .C2(n9835), .A(n9686), .B(n9685), .ZN(n9688)
         );
  INV_X1 U10989 ( .A(n9688), .ZN(n9690) );
  NAND3_X1 U10990 ( .A1(n9691), .A2(n9690), .A3(n9689), .ZN(P1_U3247) );
  INV_X1 U10991 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9707) );
  OAI211_X1 U10992 ( .C1(n9694), .C2(n9693), .A(n9825), .B(n9692), .ZN(n9704)
         );
  NAND2_X1 U10993 ( .A1(n9818), .A2(n9695), .ZN(n9703) );
  INV_X1 U10994 ( .A(n9696), .ZN(n9699) );
  INV_X1 U10995 ( .A(n9697), .ZN(n9698) );
  NAND2_X1 U10996 ( .A1(n9699), .A2(n9698), .ZN(n9700) );
  NAND3_X1 U10997 ( .A1(n9829), .A2(n9701), .A3(n9700), .ZN(n9702) );
  AND3_X1 U10998 ( .A1(n9704), .A2(n9703), .A3(n9702), .ZN(n9706) );
  OAI211_X1 U10999 ( .C1(n9840), .C2(n9707), .A(n9706), .B(n9705), .ZN(
        P1_U3248) );
  INV_X1 U11000 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9721) );
  INV_X1 U11001 ( .A(n9708), .ZN(n9712) );
  INV_X1 U11002 ( .A(n9709), .ZN(n9711) );
  AOI211_X1 U11003 ( .C1(n9712), .C2(n9711), .A(n9710), .B(n9784), .ZN(n9717)
         );
  AOI211_X1 U11004 ( .C1(n9715), .C2(n9714), .A(n9713), .B(n9797), .ZN(n9716)
         );
  AOI211_X1 U11005 ( .C1(n9818), .C2(n9718), .A(n9717), .B(n9716), .ZN(n9720)
         );
  OAI211_X1 U11006 ( .C1(n9840), .C2(n9721), .A(n9720), .B(n9719), .ZN(
        P1_U3249) );
  INV_X1 U11007 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9736) );
  AOI21_X1 U11008 ( .B1(n9724), .B2(n9723), .A(n9722), .ZN(n9725) );
  NAND2_X1 U11009 ( .A1(n9825), .A2(n9725), .ZN(n9731) );
  AOI21_X1 U11010 ( .B1(n9728), .B2(n9727), .A(n9726), .ZN(n9729) );
  NAND2_X1 U11011 ( .A1(n9829), .A2(n9729), .ZN(n9730) );
  OAI211_X1 U11012 ( .C1(n9835), .C2(n9732), .A(n9731), .B(n9730), .ZN(n9733)
         );
  INV_X1 U11013 ( .A(n9733), .ZN(n9735) );
  OAI211_X1 U11014 ( .C1(n9840), .C2(n9736), .A(n9735), .B(n9734), .ZN(
        P1_U3254) );
  INV_X1 U11015 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9752) );
  INV_X1 U11016 ( .A(n9737), .ZN(n9748) );
  OAI21_X1 U11017 ( .B1(n9740), .B2(n9739), .A(n9738), .ZN(n9741) );
  NAND2_X1 U11018 ( .A1(n9825), .A2(n9741), .ZN(n9747) );
  OAI21_X1 U11019 ( .B1(n9744), .B2(n9743), .A(n9742), .ZN(n9745) );
  NAND2_X1 U11020 ( .A1(n9829), .A2(n9745), .ZN(n9746) );
  OAI211_X1 U11021 ( .C1(n9835), .C2(n9748), .A(n9747), .B(n9746), .ZN(n9749)
         );
  INV_X1 U11022 ( .A(n9749), .ZN(n9751) );
  OAI211_X1 U11023 ( .C1(n9840), .C2(n9752), .A(n9751), .B(n9750), .ZN(
        P1_U3255) );
  INV_X1 U11024 ( .A(n9753), .ZN(n9764) );
  AOI21_X1 U11025 ( .B1(n9756), .B2(n9755), .A(n9754), .ZN(n9757) );
  NAND2_X1 U11026 ( .A1(n9825), .A2(n9757), .ZN(n9763) );
  AOI21_X1 U11027 ( .B1(n9760), .B2(n9759), .A(n9758), .ZN(n9761) );
  NAND2_X1 U11028 ( .A1(n9829), .A2(n9761), .ZN(n9762) );
  OAI211_X1 U11029 ( .C1(n9835), .C2(n9764), .A(n9763), .B(n9762), .ZN(n9765)
         );
  INV_X1 U11030 ( .A(n9765), .ZN(n9767) );
  OAI211_X1 U11031 ( .C1(n9768), .C2(n9840), .A(n9767), .B(n9766), .ZN(
        P1_U3256) );
  INV_X1 U11032 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9783) );
  AOI21_X1 U11033 ( .B1(n9771), .B2(n9770), .A(n9769), .ZN(n9772) );
  NAND2_X1 U11034 ( .A1(n9825), .A2(n9772), .ZN(n9778) );
  AOI21_X1 U11035 ( .B1(n9775), .B2(n9774), .A(n9773), .ZN(n9776) );
  NAND2_X1 U11036 ( .A1(n9829), .A2(n9776), .ZN(n9777) );
  OAI211_X1 U11037 ( .C1(n9835), .C2(n9779), .A(n9778), .B(n9777), .ZN(n9780)
         );
  INV_X1 U11038 ( .A(n9780), .ZN(n9782) );
  OAI211_X1 U11039 ( .C1(n9840), .C2(n9783), .A(n9782), .B(n9781), .ZN(
        P1_U3257) );
  INV_X1 U11040 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9796) );
  AOI211_X1 U11041 ( .C1(n9787), .C2(n9786), .A(n9785), .B(n9784), .ZN(n9792)
         );
  AOI211_X1 U11042 ( .C1(n9790), .C2(n9789), .A(n9788), .B(n9797), .ZN(n9791)
         );
  AOI211_X1 U11043 ( .C1(n9818), .C2(n9793), .A(n9792), .B(n9791), .ZN(n9795)
         );
  OAI211_X1 U11044 ( .C1(n9840), .C2(n9796), .A(n9795), .B(n9794), .ZN(
        P1_U3258) );
  AOI211_X1 U11045 ( .C1(n9800), .C2(n9799), .A(n9798), .B(n9797), .ZN(n9801)
         );
  AOI211_X1 U11046 ( .C1(P1_ADDR_REG_16__SCAN_IN), .C2(n9803), .A(n9802), .B(
        n9801), .ZN(n9810) );
  OAI21_X1 U11047 ( .B1(n9806), .B2(n9805), .A(n9804), .ZN(n9808) );
  AOI22_X1 U11048 ( .A1(n9808), .A2(n9829), .B1(n9807), .B2(n9818), .ZN(n9809)
         );
  NAND2_X1 U11049 ( .A1(n9810), .A2(n9809), .ZN(P1_U3259) );
  OAI21_X1 U11050 ( .B1(n9813), .B2(n9812), .A(n9811), .ZN(n9820) );
  OAI21_X1 U11051 ( .B1(n9816), .B2(n9815), .A(n9814), .ZN(n9817) );
  AOI222_X1 U11052 ( .A1(n9820), .A2(n9825), .B1(n9819), .B2(n9818), .C1(n9817), .C2(n9829), .ZN(n9822) );
  OAI211_X1 U11053 ( .C1(n9840), .C2(n9823), .A(n9822), .B(n9821), .ZN(
        P1_U3260) );
  OAI211_X1 U11054 ( .C1(n9827), .C2(n9826), .A(n9825), .B(n9824), .ZN(n9833)
         );
  OAI211_X1 U11055 ( .C1(n9831), .C2(n9830), .A(n9829), .B(n9828), .ZN(n9832)
         );
  OAI211_X1 U11056 ( .C1(n9835), .C2(n9834), .A(n9833), .B(n9832), .ZN(n9836)
         );
  INV_X1 U11057 ( .A(n9836), .ZN(n9838) );
  OAI211_X1 U11058 ( .C1(n9840), .C2(n9839), .A(n9838), .B(n9837), .ZN(
        P1_U3261) );
  NAND2_X1 U11059 ( .A1(n9842), .A2(n9841), .ZN(n9843) );
  XNOR2_X1 U11060 ( .A(n9843), .B(n9847), .ZN(n9850) );
  OAI22_X1 U11061 ( .A1(n9845), .A2(n9883), .B1(n9844), .B2(n9881), .ZN(n9849)
         );
  XOR2_X1 U11062 ( .A(n9847), .B(n9846), .Z(n9992) );
  NOR2_X1 U11063 ( .A1(n9992), .A2(n9887), .ZN(n9848) );
  AOI211_X1 U11064 ( .C1(n9850), .C2(n9890), .A(n9849), .B(n9848), .ZN(n9990)
         );
  AOI222_X1 U11065 ( .A1(n9988), .A2(n9854), .B1(n9853), .B2(n9852), .C1(
        P1_REG2_REG_11__SCAN_IN), .C2(n9851), .ZN(n9859) );
  INV_X1 U11066 ( .A(n9992), .ZN(n9857) );
  AOI211_X1 U11067 ( .C1(n9988), .C2(n9856), .A(n9944), .B(n9855), .ZN(n9987)
         );
  AOI22_X1 U11068 ( .A1(n9857), .A2(n9904), .B1(n9903), .B2(n9987), .ZN(n9858)
         );
  OAI211_X1 U11069 ( .C1(n9907), .C2(n9990), .A(n9859), .B(n9858), .ZN(
        P1_U3282) );
  OAI211_X1 U11070 ( .C1(n9862), .C2(n9861), .A(n9860), .B(n9890), .ZN(n9867)
         );
  AOI22_X1 U11071 ( .A1(n9865), .A2(n9864), .B1(n9996), .B2(n9863), .ZN(n9866)
         );
  AND2_X1 U11072 ( .A1(n9867), .A2(n9866), .ZN(n9952) );
  NOR2_X1 U11073 ( .A1(n9893), .A2(n9868), .ZN(n9869) );
  AOI21_X1 U11074 ( .B1(n9907), .B2(P1_REG2_REG_5__SCAN_IN), .A(n9869), .ZN(
        n9870) );
  OAI21_X1 U11075 ( .B1(n9896), .B2(n9953), .A(n9870), .ZN(n9871) );
  INV_X1 U11076 ( .A(n9871), .ZN(n9879) );
  XNOR2_X1 U11077 ( .A(n9872), .B(n9873), .ZN(n9955) );
  OAI211_X1 U11078 ( .C1(n9875), .C2(n9953), .A(n9874), .B(n9900), .ZN(n9951)
         );
  INV_X1 U11079 ( .A(n9951), .ZN(n9876) );
  AOI22_X1 U11080 ( .A1(n9955), .A2(n9877), .B1(n9903), .B2(n9876), .ZN(n9878)
         );
  OAI211_X1 U11081 ( .C1(n9907), .C2(n9952), .A(n9879), .B(n9878), .ZN(
        P1_U3288) );
  XNOR2_X1 U11082 ( .A(n9880), .B(n9885), .ZN(n9891) );
  OAI22_X1 U11083 ( .A1(n9884), .A2(n9883), .B1(n9882), .B2(n9881), .ZN(n9889)
         );
  XOR2_X1 U11084 ( .A(n9886), .B(n9885), .Z(n9898) );
  NOR2_X1 U11085 ( .A1(n9898), .A2(n9887), .ZN(n9888) );
  AOI211_X1 U11086 ( .C1(n9891), .C2(n9890), .A(n9889), .B(n9888), .ZN(n9921)
         );
  NOR2_X1 U11087 ( .A1(n9893), .A2(n9892), .ZN(n9894) );
  AOI21_X1 U11088 ( .B1(n9907), .B2(P1_REG2_REG_1__SCAN_IN), .A(n9894), .ZN(
        n9895) );
  OAI21_X1 U11089 ( .B1(n9896), .B2(n9920), .A(n9895), .ZN(n9897) );
  INV_X1 U11090 ( .A(n9897), .ZN(n9906) );
  INV_X1 U11091 ( .A(n9898), .ZN(n9924) );
  OAI211_X1 U11092 ( .C1(n9920), .C2(n9901), .A(n9900), .B(n9899), .ZN(n9919)
         );
  INV_X1 U11093 ( .A(n9919), .ZN(n9902) );
  AOI22_X1 U11094 ( .A1(n9924), .A2(n9904), .B1(n9903), .B2(n9902), .ZN(n9905)
         );
  OAI211_X1 U11095 ( .C1(n9907), .C2(n9921), .A(n9906), .B(n9905), .ZN(
        P1_U3292) );
  NOR2_X1 U11096 ( .A1(n9917), .A2(n9908), .ZN(P1_U3294) );
  AND2_X1 U11097 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9918), .ZN(P1_U3295) );
  AND2_X1 U11098 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9918), .ZN(P1_U3296) );
  AND2_X1 U11099 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9918), .ZN(P1_U3297) );
  AND2_X1 U11100 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9918), .ZN(P1_U3298) );
  AND2_X1 U11101 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9918), .ZN(P1_U3299) );
  NOR2_X1 U11102 ( .A1(n9917), .A2(n9909), .ZN(P1_U3300) );
  AND2_X1 U11103 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9918), .ZN(P1_U3301) );
  AND2_X1 U11104 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9918), .ZN(P1_U3302) );
  NOR2_X1 U11105 ( .A1(n9917), .A2(n9910), .ZN(P1_U3303) );
  AND2_X1 U11106 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9918), .ZN(P1_U3304) );
  NOR2_X1 U11107 ( .A1(n9917), .A2(n9911), .ZN(P1_U3305) );
  AND2_X1 U11108 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9918), .ZN(P1_U3306) );
  AND2_X1 U11109 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9918), .ZN(P1_U3307) );
  AND2_X1 U11110 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9918), .ZN(P1_U3308) );
  AND2_X1 U11111 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9918), .ZN(P1_U3309) );
  NOR2_X1 U11112 ( .A1(n9917), .A2(n9912), .ZN(P1_U3310) );
  NOR2_X1 U11113 ( .A1(n9917), .A2(n9913), .ZN(P1_U3311) );
  AND2_X1 U11114 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9918), .ZN(P1_U3312) );
  AND2_X1 U11115 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9918), .ZN(P1_U3313) );
  AND2_X1 U11116 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9918), .ZN(P1_U3314) );
  AND2_X1 U11117 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9918), .ZN(P1_U3315) );
  NOR2_X1 U11118 ( .A1(n9917), .A2(n9914), .ZN(P1_U3316) );
  AND2_X1 U11119 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9918), .ZN(P1_U3317) );
  NOR2_X1 U11120 ( .A1(n9917), .A2(n9915), .ZN(P1_U3318) );
  AND2_X1 U11121 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9918), .ZN(P1_U3319) );
  AND2_X1 U11122 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9918), .ZN(P1_U3320) );
  AND2_X1 U11123 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9918), .ZN(P1_U3321) );
  NOR2_X1 U11124 ( .A1(n9917), .A2(n9916), .ZN(P1_U3322) );
  AND2_X1 U11125 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9918), .ZN(P1_U3323) );
  INV_X1 U11126 ( .A(n9991), .ZN(n9969) );
  OAI21_X1 U11127 ( .B1(n9920), .B2(n10007), .A(n9919), .ZN(n9923) );
  INV_X1 U11128 ( .A(n9921), .ZN(n9922) );
  AOI211_X1 U11129 ( .C1(n9969), .C2(n9924), .A(n9923), .B(n9922), .ZN(n10015)
         );
  INV_X1 U11130 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9925) );
  AOI22_X1 U11131 ( .A1(n10013), .A2(n10015), .B1(n9925), .B2(n10011), .ZN(
        P1_U3456) );
  INV_X1 U11132 ( .A(n9926), .ZN(n9932) );
  INV_X1 U11133 ( .A(n9927), .ZN(n9928) );
  OAI211_X1 U11134 ( .C1(n9930), .C2(n10007), .A(n9929), .B(n9928), .ZN(n9931)
         );
  AOI21_X1 U11135 ( .B1(n10009), .B2(n9932), .A(n9931), .ZN(n10017) );
  AOI22_X1 U11136 ( .A1(n10013), .A2(n10017), .B1(n9933), .B2(n10011), .ZN(
        P1_U3459) );
  AOI22_X1 U11137 ( .A1(n9935), .A2(n9997), .B1(n9996), .B2(n9934), .ZN(n9937)
         );
  NAND3_X1 U11138 ( .A1(n9938), .A2(n9937), .A3(n9936), .ZN(n9939) );
  AOI21_X1 U11139 ( .B1(n9940), .B2(n10009), .A(n9939), .ZN(n10019) );
  INV_X1 U11140 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9941) );
  AOI22_X1 U11141 ( .A1(n10013), .A2(n10019), .B1(n9941), .B2(n10011), .ZN(
        P1_U3462) );
  INV_X1 U11142 ( .A(n9942), .ZN(n9945) );
  OAI22_X1 U11143 ( .A1(n9945), .A2(n9944), .B1(n9943), .B2(n10007), .ZN(n9948) );
  INV_X1 U11144 ( .A(n9946), .ZN(n9947) );
  AOI211_X1 U11145 ( .C1(n10009), .C2(n9949), .A(n9948), .B(n9947), .ZN(n10020) );
  INV_X1 U11146 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9950) );
  AOI22_X1 U11147 ( .A1(n10013), .A2(n10020), .B1(n9950), .B2(n10011), .ZN(
        P1_U3465) );
  OAI211_X1 U11148 ( .C1(n9953), .C2(n10007), .A(n9952), .B(n9951), .ZN(n9954)
         );
  AOI21_X1 U11149 ( .B1(n10009), .B2(n9955), .A(n9954), .ZN(n10022) );
  INV_X1 U11150 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9956) );
  AOI22_X1 U11151 ( .A1(n10013), .A2(n10022), .B1(n9956), .B2(n10011), .ZN(
        P1_U3468) );
  OAI21_X1 U11152 ( .B1(n9958), .B2(n10007), .A(n9957), .ZN(n9960) );
  AOI211_X1 U11153 ( .C1(n9969), .C2(n9961), .A(n9960), .B(n9959), .ZN(n10023)
         );
  INV_X1 U11154 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9962) );
  AOI22_X1 U11155 ( .A1(n10013), .A2(n10023), .B1(n9962), .B2(n10011), .ZN(
        P1_U3474) );
  INV_X1 U11156 ( .A(n9963), .ZN(n9968) );
  OAI21_X1 U11157 ( .B1(n9965), .B2(n10007), .A(n9964), .ZN(n9967) );
  AOI211_X1 U11158 ( .C1(n9969), .C2(n9968), .A(n9967), .B(n9966), .ZN(n10025)
         );
  INV_X1 U11159 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9970) );
  AOI22_X1 U11160 ( .A1(n10013), .A2(n10025), .B1(n9970), .B2(n10011), .ZN(
        P1_U3477) );
  AOI22_X1 U11161 ( .A1(n9972), .A2(n9997), .B1(n9996), .B2(n9971), .ZN(n9973)
         );
  NAND3_X1 U11162 ( .A1(n9975), .A2(n9974), .A3(n9973), .ZN(n9976) );
  AOI21_X1 U11163 ( .B1(n10009), .B2(n9977), .A(n9976), .ZN(n10027) );
  INV_X1 U11164 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9978) );
  AOI22_X1 U11165 ( .A1(n10013), .A2(n10027), .B1(n9978), .B2(n10011), .ZN(
        P1_U3480) );
  AOI22_X1 U11166 ( .A1(n9980), .A2(n9997), .B1(n9996), .B2(n9979), .ZN(n9981)
         );
  NAND2_X1 U11167 ( .A1(n9982), .A2(n9981), .ZN(n9984) );
  AOI211_X1 U11168 ( .C1(n10009), .C2(n9985), .A(n9984), .B(n9983), .ZN(n10028) );
  AOI22_X1 U11169 ( .A1(n10013), .A2(n10028), .B1(n9986), .B2(n10011), .ZN(
        P1_U3483) );
  AOI21_X1 U11170 ( .B1(n9997), .B2(n9988), .A(n9987), .ZN(n9989) );
  OAI211_X1 U11171 ( .C1(n9992), .C2(n9991), .A(n9990), .B(n9989), .ZN(n9993)
         );
  INV_X1 U11172 ( .A(n9993), .ZN(n10029) );
  AOI22_X1 U11173 ( .A1(n10013), .A2(n10029), .B1(n9994), .B2(n10011), .ZN(
        P1_U3486) );
  AOI22_X1 U11174 ( .A1(n9998), .A2(n9997), .B1(n9996), .B2(n9995), .ZN(n10000) );
  NAND3_X1 U11175 ( .A1(n10001), .A2(n10000), .A3(n9999), .ZN(n10002) );
  AOI21_X1 U11176 ( .B1(n10003), .B2(n10009), .A(n10002), .ZN(n10030) );
  INV_X1 U11177 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10004) );
  AOI22_X1 U11178 ( .A1(n10013), .A2(n10030), .B1(n10004), .B2(n10011), .ZN(
        P1_U3489) );
  OAI211_X1 U11179 ( .C1(n4774), .C2(n10007), .A(n10006), .B(n10005), .ZN(
        n10008) );
  AOI21_X1 U11180 ( .B1(n10010), .B2(n10009), .A(n10008), .ZN(n10032) );
  INV_X1 U11181 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10012) );
  AOI22_X1 U11182 ( .A1(n10013), .A2(n10032), .B1(n10012), .B2(n10011), .ZN(
        P1_U3492) );
  INV_X1 U11183 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10014) );
  AOI22_X1 U11184 ( .A1(n10033), .A2(n10015), .B1(n10014), .B2(n10031), .ZN(
        P1_U3523) );
  INV_X1 U11185 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10016) );
  AOI22_X1 U11186 ( .A1(n10033), .A2(n10017), .B1(n10016), .B2(n10031), .ZN(
        P1_U3524) );
  INV_X1 U11187 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10018) );
  AOI22_X1 U11188 ( .A1(n10033), .A2(n10019), .B1(n10018), .B2(n10031), .ZN(
        P1_U3525) );
  AOI22_X1 U11189 ( .A1(n10033), .A2(n10020), .B1(n6939), .B2(n10031), .ZN(
        P1_U3526) );
  INV_X1 U11190 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10021) );
  AOI22_X1 U11191 ( .A1(n10033), .A2(n10022), .B1(n10021), .B2(n10031), .ZN(
        P1_U3527) );
  AOI22_X1 U11192 ( .A1(n10033), .A2(n10023), .B1(n6946), .B2(n10031), .ZN(
        P1_U3529) );
  INV_X1 U11193 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10024) );
  AOI22_X1 U11194 ( .A1(n10033), .A2(n10025), .B1(n10024), .B2(n10031), .ZN(
        P1_U3530) );
  AOI22_X1 U11195 ( .A1(n10033), .A2(n10027), .B1(n10026), .B2(n10031), .ZN(
        P1_U3531) );
  AOI22_X1 U11196 ( .A1(n10033), .A2(n10028), .B1(n9098), .B2(n10031), .ZN(
        P1_U3532) );
  AOI22_X1 U11197 ( .A1(n10033), .A2(n10029), .B1(n9100), .B2(n10031), .ZN(
        P1_U3533) );
  AOI22_X1 U11198 ( .A1(n10033), .A2(n10030), .B1(n9101), .B2(n10031), .ZN(
        P1_U3534) );
  AOI22_X1 U11199 ( .A1(n10033), .A2(n10032), .B1(n9097), .B2(n10031), .ZN(
        P1_U3535) );
  AOI22_X1 U11200 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n10115), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n10038) );
  OAI21_X1 U11201 ( .B1(n10036), .B2(n10143), .A(n10035), .ZN(n10037) );
  OAI211_X1 U11202 ( .C1(n10112), .C2(n10039), .A(n10038), .B(n10037), .ZN(
        P2_U3182) );
  XOR2_X1 U11203 ( .A(n10040), .B(n10041), .Z(n10042) );
  NAND2_X1 U11204 ( .A1(n10042), .A2(n10143), .ZN(n10043) );
  OAI21_X1 U11205 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n10044), .A(n10043), .ZN(
        n10055) );
  AOI21_X1 U11206 ( .B1(n10241), .B2(n10046), .A(n10045), .ZN(n10053) );
  AND2_X1 U11207 ( .A1(n10048), .A2(n10047), .ZN(n10050) );
  INV_X1 U11208 ( .A(n10135), .ZN(n10049) );
  OAI21_X1 U11209 ( .B1(n10051), .B2(n10050), .A(n10049), .ZN(n10052) );
  OAI21_X1 U11210 ( .B1(n10133), .B2(n10053), .A(n10052), .ZN(n10054) );
  AOI211_X1 U11211 ( .C1(n10115), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n10055), .B(
        n10054), .ZN(n10056) );
  OAI21_X1 U11212 ( .B1(n10057), .B2(n10112), .A(n10056), .ZN(P2_U3183) );
  INV_X1 U11213 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10152) );
  XOR2_X1 U11214 ( .A(n10059), .B(n10058), .Z(n10060) );
  NAND2_X1 U11215 ( .A1(n10060), .A2(n10143), .ZN(n10061) );
  OAI21_X1 U11216 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n10152), .A(n10061), .ZN(
        n10072) );
  INV_X1 U11217 ( .A(n10062), .ZN(n10065) );
  AOI21_X1 U11218 ( .B1(n10065), .B2(n10064), .A(n10063), .ZN(n10070) );
  AOI21_X1 U11219 ( .B1(n10068), .B2(n10067), .A(n10066), .ZN(n10069) );
  OAI22_X1 U11220 ( .A1(n10133), .A2(n10070), .B1(n10069), .B2(n10135), .ZN(
        n10071) );
  AOI211_X1 U11221 ( .C1(n10115), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n10072), .B(
        n10071), .ZN(n10073) );
  OAI21_X1 U11222 ( .B1(n10112), .B2(n4571), .A(n10073), .ZN(P2_U3184) );
  AOI21_X1 U11223 ( .B1(n10077), .B2(n10076), .A(n10075), .ZN(n10079) );
  OAI22_X1 U11224 ( .A1(n10079), .A2(n10135), .B1(n10112), .B2(n10078), .ZN(
        n10080) );
  AOI21_X1 U11225 ( .B1(n10115), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n10080), .ZN(
        n10089) );
  XOR2_X1 U11226 ( .A(n10082), .B(n10081), .Z(n10083) );
  NAND2_X1 U11227 ( .A1(n10083), .A2(n10143), .ZN(n10087) );
  XNOR2_X1 U11228 ( .A(n10084), .B(n10248), .ZN(n10085) );
  NAND2_X1 U11229 ( .A1(n10121), .A2(n10085), .ZN(n10086) );
  NAND4_X1 U11230 ( .A1(n10089), .A2(n10088), .A3(n10087), .A4(n10086), .ZN(
        P2_U3187) );
  INV_X1 U11231 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10107) );
  AOI21_X1 U11232 ( .B1(n10092), .B2(n10091), .A(n10090), .ZN(n10097) );
  AOI21_X1 U11233 ( .B1(n10095), .B2(n10094), .A(n10093), .ZN(n10096) );
  OAI22_X1 U11234 ( .A1(n10097), .A2(n10133), .B1(n10096), .B2(n10135), .ZN(
        n10098) );
  AOI211_X1 U11235 ( .C1(n10100), .C2(n10139), .A(n10099), .B(n10098), .ZN(
        n10106) );
  OAI21_X1 U11236 ( .B1(n10103), .B2(n10102), .A(n10101), .ZN(n10104) );
  NAND2_X1 U11237 ( .A1(n10104), .A2(n10143), .ZN(n10105) );
  OAI211_X1 U11238 ( .C1(n10107), .C2(n10148), .A(n10106), .B(n10105), .ZN(
        P2_U3188) );
  AOI21_X1 U11239 ( .B1(n10110), .B2(n10109), .A(n10108), .ZN(n10113) );
  OAI22_X1 U11240 ( .A1(n10113), .A2(n10135), .B1(n10112), .B2(n10111), .ZN(
        n10114) );
  AOI21_X1 U11241 ( .B1(n10115), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n10114), .ZN(
        n10126) );
  OAI21_X1 U11242 ( .B1(n10118), .B2(n10117), .A(n10116), .ZN(n10119) );
  NAND2_X1 U11243 ( .A1(n10119), .A2(n10143), .ZN(n10124) );
  XNOR2_X1 U11244 ( .A(n10120), .B(n10252), .ZN(n10122) );
  NAND2_X1 U11245 ( .A1(n10122), .A2(n10121), .ZN(n10123) );
  NAND4_X1 U11246 ( .A1(n10126), .A2(n10125), .A3(n10124), .A4(n10123), .ZN(
        P2_U3189) );
  INV_X1 U11247 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10149) );
  AOI21_X1 U11248 ( .B1(n10129), .B2(n10128), .A(n10127), .ZN(n10136) );
  AOI21_X1 U11249 ( .B1(n10132), .B2(n10131), .A(n10130), .ZN(n10134) );
  OAI22_X1 U11250 ( .A1(n10136), .A2(n10135), .B1(n10134), .B2(n10133), .ZN(
        n10137) );
  AOI211_X1 U11251 ( .C1(n10140), .C2(n10139), .A(n10138), .B(n10137), .ZN(
        n10147) );
  NOR2_X1 U11252 ( .A1(n10142), .A2(n10141), .ZN(n10144) );
  OAI21_X1 U11253 ( .B1(n10145), .B2(n10144), .A(n10143), .ZN(n10146) );
  OAI211_X1 U11254 ( .C1(n10149), .C2(n10148), .A(n10147), .B(n10146), .ZN(
        P2_U3190) );
  XNOR2_X1 U11255 ( .A(n10150), .B(n10156), .ZN(n10164) );
  INV_X1 U11256 ( .A(n10164), .ZN(n10177) );
  OAI22_X1 U11257 ( .A1(n10154), .A2(n10153), .B1(n10152), .B2(n10151), .ZN(
        n10165) );
  XNOR2_X1 U11258 ( .A(n10155), .B(n10156), .ZN(n10161) );
  OAI22_X1 U11259 ( .A1(n10159), .A2(n10158), .B1(n6757), .B2(n10157), .ZN(
        n10160) );
  AOI21_X1 U11260 ( .B1(n10161), .B2(n6797), .A(n10160), .ZN(n10162) );
  OAI21_X1 U11261 ( .B1(n10164), .B2(n10163), .A(n10162), .ZN(n10175) );
  AOI211_X1 U11262 ( .C1(n10166), .C2(n10177), .A(n10165), .B(n10175), .ZN(
        n10168) );
  AOI22_X1 U11263 ( .A1(n8442), .A2(n10169), .B1(n10168), .B2(n10167), .ZN(
        P2_U3231) );
  INV_X1 U11264 ( .A(n10170), .ZN(n10171) );
  AOI211_X1 U11265 ( .C1(n10234), .C2(n10173), .A(n10172), .B(n10171), .ZN(
        n10242) );
  INV_X1 U11266 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10174) );
  AOI22_X1 U11267 ( .A1(n10240), .A2(n10242), .B1(n10174), .B2(n10238), .ZN(
        P2_U3393) );
  INV_X1 U11268 ( .A(n10202), .ZN(n10218) );
  AOI211_X1 U11269 ( .C1(n10218), .C2(n10177), .A(n10176), .B(n10175), .ZN(
        n10244) );
  INV_X1 U11270 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10178) );
  AOI22_X1 U11271 ( .A1(n10240), .A2(n10244), .B1(n10178), .B2(n10238), .ZN(
        P2_U3396) );
  AOI22_X1 U11272 ( .A1(n10181), .A2(n10234), .B1(n10180), .B2(n10179), .ZN(
        n10182) );
  AND2_X1 U11273 ( .A1(n10183), .A2(n10182), .ZN(n10246) );
  INV_X1 U11274 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10184) );
  AOI22_X1 U11275 ( .A1(n10240), .A2(n10246), .B1(n10184), .B2(n10238), .ZN(
        P2_U3399) );
  INV_X1 U11276 ( .A(n10185), .ZN(n10186) );
  AOI211_X1 U11277 ( .C1(n10234), .C2(n10188), .A(n10187), .B(n10186), .ZN(
        n10247) );
  INV_X1 U11278 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10189) );
  AOI22_X1 U11279 ( .A1(n10240), .A2(n10247), .B1(n10189), .B2(n10238), .ZN(
        P2_U3402) );
  INV_X1 U11280 ( .A(n10190), .ZN(n10192) );
  OAI21_X1 U11281 ( .B1(n10192), .B2(n10202), .A(n10191), .ZN(n10193) );
  NOR2_X1 U11282 ( .A1(n10194), .A2(n10193), .ZN(n10249) );
  INV_X1 U11283 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10195) );
  AOI22_X1 U11284 ( .A1(n10240), .A2(n10249), .B1(n10195), .B2(n10238), .ZN(
        P2_U3405) );
  INV_X1 U11285 ( .A(n10196), .ZN(n10197) );
  AOI211_X1 U11286 ( .C1(n10234), .C2(n10199), .A(n10198), .B(n10197), .ZN(
        n10251) );
  AOI22_X1 U11287 ( .A1(n10240), .A2(n10251), .B1(n10200), .B2(n10238), .ZN(
        P2_U3408) );
  OAI22_X1 U11288 ( .A1(n10203), .A2(n10202), .B1(n10201), .B2(n10225), .ZN(
        n10205) );
  AOI211_X1 U11289 ( .C1(n10207), .C2(n10206), .A(n10205), .B(n10204), .ZN(
        n10253) );
  INV_X1 U11290 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10208) );
  AOI22_X1 U11291 ( .A1(n10240), .A2(n10253), .B1(n10208), .B2(n10238), .ZN(
        P2_U3411) );
  INV_X1 U11292 ( .A(n10209), .ZN(n10210) );
  AOI211_X1 U11293 ( .C1(n10234), .C2(n10212), .A(n10211), .B(n10210), .ZN(
        n10255) );
  AOI22_X1 U11294 ( .A1(n10240), .A2(n10255), .B1(n10213), .B2(n10238), .ZN(
        P2_U3414) );
  INV_X1 U11295 ( .A(n10214), .ZN(n10217) );
  AOI211_X1 U11296 ( .C1(n10218), .C2(n10217), .A(n10216), .B(n10215), .ZN(
        n10257) );
  AOI22_X1 U11297 ( .A1(n10240), .A2(n10257), .B1(n10219), .B2(n10238), .ZN(
        P2_U3417) );
  INV_X1 U11298 ( .A(n10220), .ZN(n10222) );
  AOI211_X1 U11299 ( .C1(n10234), .C2(n10223), .A(n10222), .B(n10221), .ZN(
        n10259) );
  INV_X1 U11300 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10224) );
  AOI22_X1 U11301 ( .A1(n10240), .A2(n10259), .B1(n10224), .B2(n10238), .ZN(
        P2_U3420) );
  OAI22_X1 U11302 ( .A1(n10228), .A2(n10227), .B1(n10226), .B2(n10225), .ZN(
        n10229) );
  NOR2_X1 U11303 ( .A1(n10230), .A2(n10229), .ZN(n10261) );
  AOI22_X1 U11304 ( .A1(n10240), .A2(n10261), .B1(n10231), .B2(n10238), .ZN(
        P2_U3423) );
  INV_X1 U11305 ( .A(n10232), .ZN(n10233) );
  AOI21_X1 U11306 ( .B1(n10235), .B2(n10234), .A(n10233), .ZN(n10236) );
  AND2_X1 U11307 ( .A1(n10237), .A2(n10236), .ZN(n10263) );
  AOI22_X1 U11308 ( .A1(n10240), .A2(n10263), .B1(n10239), .B2(n10238), .ZN(
        P2_U3426) );
  AOI22_X1 U11309 ( .A1(n10264), .A2(n10242), .B1(n10241), .B2(n10262), .ZN(
        P2_U3460) );
  INV_X1 U11310 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10243) );
  AOI22_X1 U11311 ( .A1(n10264), .A2(n10244), .B1(n10243), .B2(n10262), .ZN(
        P2_U3461) );
  AOI22_X1 U11312 ( .A1(n10264), .A2(n10246), .B1(n10245), .B2(n10262), .ZN(
        P2_U3462) );
  AOI22_X1 U11313 ( .A1(n10264), .A2(n10247), .B1(n7142), .B2(n10262), .ZN(
        P2_U3463) );
  AOI22_X1 U11314 ( .A1(n10264), .A2(n10249), .B1(n10248), .B2(n10262), .ZN(
        P2_U3464) );
  AOI22_X1 U11315 ( .A1(n10264), .A2(n10251), .B1(n10250), .B2(n10262), .ZN(
        P2_U3465) );
  AOI22_X1 U11316 ( .A1(n10264), .A2(n10253), .B1(n10252), .B2(n10262), .ZN(
        P2_U3466) );
  AOI22_X1 U11317 ( .A1(n10264), .A2(n10255), .B1(n10254), .B2(n10262), .ZN(
        P2_U3467) );
  AOI22_X1 U11318 ( .A1(n10264), .A2(n10257), .B1(n10256), .B2(n10262), .ZN(
        P2_U3468) );
  AOI22_X1 U11319 ( .A1(n10264), .A2(n10259), .B1(n10258), .B2(n10262), .ZN(
        P2_U3469) );
  AOI22_X1 U11320 ( .A1(n10264), .A2(n10261), .B1(n10260), .B2(n10262), .ZN(
        P2_U3470) );
  AOI22_X1 U11321 ( .A1(n10264), .A2(n10263), .B1(n8096), .B2(n10262), .ZN(
        P2_U3471) );
  OAI222_X1 U11322 ( .A1(n10269), .A2(n10268), .B1(n10269), .B2(n10267), .C1(
        n10266), .C2(n10265), .ZN(ADD_1068_U5) );
  XOR2_X1 U11323 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  INV_X1 U11324 ( .A(n10272), .ZN(n10271) );
  OAI222_X1 U11325 ( .A1(n10274), .A2(n10273), .B1(n10274), .B2(n10272), .C1(
        n10271), .C2(n10270), .ZN(ADD_1068_U55) );
  OAI21_X1 U11326 ( .B1(n10277), .B2(n10276), .A(n10275), .ZN(ADD_1068_U56) );
  OAI21_X1 U11327 ( .B1(n10280), .B2(n10279), .A(n10278), .ZN(ADD_1068_U57) );
  OAI21_X1 U11328 ( .B1(n10283), .B2(n10282), .A(n10281), .ZN(ADD_1068_U58) );
  OAI21_X1 U11329 ( .B1(n10286), .B2(n10285), .A(n10284), .ZN(ADD_1068_U59) );
  OAI21_X1 U11330 ( .B1(n10289), .B2(n10288), .A(n10287), .ZN(ADD_1068_U60) );
  OAI21_X1 U11331 ( .B1(n10292), .B2(n10291), .A(n10290), .ZN(ADD_1068_U61) );
  OAI21_X1 U11332 ( .B1(n10295), .B2(n10294), .A(n10293), .ZN(ADD_1068_U62) );
  OAI21_X1 U11333 ( .B1(n10298), .B2(n10297), .A(n10296), .ZN(ADD_1068_U63) );
  OAI21_X1 U11334 ( .B1(n10301), .B2(n10300), .A(n10299), .ZN(ADD_1068_U50) );
  OAI21_X1 U11335 ( .B1(n10304), .B2(n10303), .A(n10302), .ZN(ADD_1068_U51) );
  OAI21_X1 U11336 ( .B1(n10307), .B2(n10306), .A(n10305), .ZN(ADD_1068_U47) );
  OAI21_X1 U11337 ( .B1(n10310), .B2(n10309), .A(n10308), .ZN(ADD_1068_U49) );
  OAI21_X1 U11338 ( .B1(n10313), .B2(n10312), .A(n10311), .ZN(ADD_1068_U48) );
  AOI21_X1 U11339 ( .B1(n10316), .B2(n10315), .A(n10314), .ZN(ADD_1068_U54) );
  AOI21_X1 U11340 ( .B1(n10319), .B2(n10318), .A(n10317), .ZN(ADD_1068_U53) );
  OAI21_X1 U11341 ( .B1(n10322), .B2(n10321), .A(n10320), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U4968 ( .A(n6019), .Z(n4462) );
  CLKBUF_X1 U4969 ( .A(n5075), .Z(n9557) );
  INV_X1 U5128 ( .A(n6744), .ZN(n7433) );
endmodule

