

module b14_C_AntiSAT_k_256_9 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990;

  CLKBUF_X2 U2474 ( .A(n2508), .Z(n3040) );
  INV_X1 U2475 ( .A(n3295), .ZN(n3291) );
  INV_X4 U2476 ( .A(n2232), .ZN(n2233) );
  CLKBUF_X2 U2477 ( .A(n2482), .Z(n3489) );
  INV_X1 U2478 ( .A(n3172), .ZN(n3246) );
  BUF_X2 U2479 ( .A(n2466), .Z(n2950) );
  NAND2_X1 U2480 ( .A1(n2408), .A2(IR_REG_31__SCAN_IN), .ZN(n2410) );
  XNOR2_X1 U2481 ( .A(n2430), .B(IR_REG_1__SCAN_IN), .ZN(n4682) );
  INV_X1 U2483 ( .A(n3038), .ZN(n2846) );
  INV_X1 U2484 ( .A(n2943), .ZN(n2232) );
  INV_X1 U2486 ( .A(IR_REG_31__SCAN_IN), .ZN(n2681) );
  NAND2_X1 U2487 ( .A1(n3500), .A2(n2565), .ZN(n3347) );
  AND2_X1 U2488 ( .A1(n2872), .A2(n4111), .ZN(n4971) );
  INV_X1 U2489 ( .A(n4134), .ZN(U4043) );
  AND2_X2 U2491 ( .A1(n2398), .A2(REG1_REG_2__SCAN_IN), .ZN(n2469) );
  NOR2_X2 U2492 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2320)
         );
  NOR2_X2 U2493 ( .A1(n2276), .A2(n2521), .ZN(n2275) );
  AND2_X4 U2494 ( .A1(n3070), .A2(n2399), .ZN(n2465) );
  NAND2_X2 U2495 ( .A1(n3485), .A2(n2395), .ZN(n2399) );
  AOI21_X2 U2496 ( .B1(n4714), .B2(n4716), .A(n4715), .ZN(n3870) );
  AOI22_X2 U2497 ( .A1(n3908), .A2(n2741), .B1(n2740), .B2(n3905), .ZN(n4714)
         );
  NAND3_X2 U2498 ( .A1(n2402), .A2(n2401), .A3(n2400), .ZN(n2899) );
  AND2_X1 U2499 ( .A1(n2397), .A2(n2396), .ZN(n2402) );
  NAND2_X2 U2500 ( .A1(n2334), .A2(n2484), .ZN(n4132) );
  OR2_X2 U2501 ( .A1(n2392), .A2(n2681), .ZN(n2391) );
  XNOR2_X2 U2502 ( .A(n2410), .B(n2409), .ZN(n2852) );
  NAND2_X1 U2503 ( .A1(n4508), .A2(n2918), .ZN(n4468) );
  NAND2_X1 U2504 ( .A1(n4054), .A2(n4057), .ZN(n4023) );
  CLKBUF_X1 U2505 ( .A(n2900), .Z(n2234) );
  NAND4_X1 U2506 ( .A1(n2501), .A2(n2500), .A3(n2499), .A4(n2498), .ZN(n3200)
         );
  INV_X1 U2507 ( .A(n3141), .ZN(n3156) );
  CLKBUF_X2 U2508 ( .A(n2447), .Z(n2496) );
  AOI21_X1 U2509 ( .B1(n3857), .B2(n2356), .A(n2353), .ZN(n2352) );
  AOI22_X2 U2510 ( .A1(n4296), .A2(n2938), .B1(n4283), .B2(n4308), .ZN(n4278)
         );
  NAND2_X1 U2511 ( .A1(n4421), .A2(n2926), .ZN(n4392) );
  NAND2_X1 U2512 ( .A1(n4450), .A2(n2375), .ZN(n4433) );
  NAND2_X1 U2513 ( .A1(n3446), .A2(n3444), .ZN(n2639) );
  NAND2_X1 U2514 ( .A1(n2325), .A2(n2246), .ZN(n3500) );
  CLKBUF_X1 U2515 ( .A(n2452), .Z(n3059) );
  NAND2_X2 U2516 ( .A1(n4117), .A2(n3162), .ZN(n3038) );
  CLKBUF_X3 U2517 ( .A(n2950), .Z(n2996) );
  NAND2_X1 U2518 ( .A1(n2446), .A2(n2445), .ZN(n3136) );
  NAND2_X1 U2519 ( .A1(n4111), .A2(n4046), .ZN(n3162) );
  BUF_X2 U2520 ( .A(n2496), .Z(n2949) );
  XNOR2_X1 U2521 ( .A(n2416), .B(n2415), .ZN(n4111) );
  NAND2_X1 U2522 ( .A1(n3070), .A2(n3065), .ZN(n2482) );
  INV_X1 U2523 ( .A(n2399), .ZN(n3065) );
  NAND2_X1 U2524 ( .A1(n2242), .A2(IR_REG_31__SCAN_IN), .ZN(n2869) );
  XNOR2_X1 U2525 ( .A(n2419), .B(IR_REG_21__SCAN_IN), .ZN(n4046) );
  NAND2_X1 U2526 ( .A1(n2438), .A2(n2437), .ZN(n2440) );
  MUX2_X1 U2527 ( .A(IR_REG_31__SCAN_IN), .B(n2394), .S(IR_REG_29__SCAN_IN), 
        .Z(n2395) );
  NAND2_X1 U2528 ( .A1(n2414), .A2(IR_REG_31__SCAN_IN), .ZN(n2438) );
  AND2_X1 U2529 ( .A1(n2298), .A2(n2413), .ZN(n2422) );
  NOR2_X1 U2530 ( .A1(n2297), .A2(IR_REG_29__SCAN_IN), .ZN(n2296) );
  NOR2_X1 U2531 ( .A1(n2350), .A2(n2348), .ZN(n2347) );
  NAND2_X1 U2532 ( .A1(n2251), .A2(n2351), .ZN(n2350) );
  AND2_X1 U2533 ( .A1(n2389), .A2(n2387), .ZN(n2295) );
  AND3_X1 U2534 ( .A1(n2424), .A2(n2421), .A3(n2427), .ZN(n2389) );
  NOR2_X1 U2535 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2387)
         );
  INV_X1 U2536 ( .A(IR_REG_21__SCAN_IN), .ZN(n2388) );
  INV_X1 U2537 ( .A(IR_REG_23__SCAN_IN), .ZN(n2868) );
  INV_X1 U2538 ( .A(IR_REG_24__SCAN_IN), .ZN(n2409) );
  NOR2_X1 U2539 ( .A1(IR_REG_2__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2321)
         );
  NOR3_X1 U2540 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .A3(
        IR_REG_15__SCAN_IN), .ZN(n2386) );
  NAND2_X1 U2541 ( .A1(n4332), .A2(n2933), .ZN(n4313) );
  NAND2_X1 U2542 ( .A1(n4334), .A2(n4333), .ZN(n4332) );
  INV_X1 U2543 ( .A(n2915), .ZN(n4855) );
  OAI21_X1 U2544 ( .B1(n3435), .B2(n2249), .A(n2372), .ZN(n2915) );
  NAND4_X1 U2545 ( .A1(n2451), .A2(n2450), .A3(n2449), .A4(n2448), .ZN(n2900)
         );
  NAND2_X1 U2546 ( .A1(n4048), .A2(n4051), .ZN(n3237) );
  NOR2_X2 U2547 ( .A1(n4444), .A2(n4713), .ZN(n4425) );
  AOI21_X2 U2548 ( .B1(n4278), .B2(n2940), .A(n2939), .ZN(n4257) );
  AND2_X4 U2549 ( .A1(n2452), .A2(n2420), .ZN(n2714) );
  AOI21_X2 U2550 ( .B1(n4433), .B2(n2924), .A(n2923), .ZN(n4423) );
  AOI21_X2 U2551 ( .B1(n4468), .B2(n2922), .A(n2921), .ZN(n4452) );
  NAND2_X1 U2552 ( .A1(n2912), .A2(n2911), .ZN(n3361) );
  INV_X4 U2553 ( .A(n2634), .ZN(n4119) );
  OAI21_X2 U2554 ( .B1(n3378), .B2(n2914), .A(n2374), .ZN(n3435) );
  AOI21_X2 U2555 ( .B1(n4392), .B2(n2927), .A(n2369), .ZN(n4371) );
  OAI21_X2 U2556 ( .B1(n4221), .B2(n4220), .A(n4219), .ZN(n4223) );
  OAI22_X2 U2557 ( .A1(n3176), .A2(n2904), .B1(n3297), .B2(n2961), .ZN(n3293)
         );
  OAI22_X2 U2558 ( .A1(n3361), .A2(n2913), .B1(n2967), .B2(n3502), .ZN(n3378)
         );
  AOI21_X2 U2559 ( .B1(n4313), .B2(n2936), .A(n2935), .ZN(n4296) );
  INV_X1 U2560 ( .A(IR_REG_18__SCAN_IN), .ZN(n2335) );
  INV_X1 U2561 ( .A(IR_REG_22__SCAN_IN), .ZN(n2351) );
  INV_X1 U2562 ( .A(n2329), .ZN(n2328) );
  INV_X1 U2563 ( .A(IR_REG_17__SCAN_IN), .ZN(n2336) );
  AOI21_X1 U2564 ( .B1(n2362), .B2(n2357), .A(n2258), .ZN(n2356) );
  INV_X1 U2565 ( .A(n2367), .ZN(n2357) );
  NAND2_X1 U2566 ( .A1(n2356), .A2(n2363), .ZN(n2354) );
  XNOR2_X1 U2567 ( .A(n2441), .B(n3038), .ZN(n2460) );
  INV_X1 U2568 ( .A(n4874), .ZN(n2872) );
  NOR2_X1 U2569 ( .A1(n4845), .A2(n4846), .ZN(n4844) );
  NOR2_X1 U2570 ( .A1(n2811), .A2(n3917), .ZN(n2837) );
  OR2_X1 U2571 ( .A1(n4874), .A2(n4111), .ZN(n4858) );
  INV_X1 U2572 ( .A(n4157), .ZN(n2263) );
  NOR2_X1 U2573 ( .A1(n4239), .A2(n4103), .ZN(n2287) );
  NAND2_X1 U2574 ( .A1(n2492), .A2(n2634), .ZN(n2326) );
  AND2_X1 U2575 ( .A1(n2674), .A2(n2236), .ZN(n2343) );
  INV_X1 U2576 ( .A(n2287), .ZN(n2284) );
  AOI21_X1 U2577 ( .B1(n2292), .B2(n2290), .A(n2289), .ZN(n2288) );
  INV_X1 U2578 ( .A(n2292), .ZN(n2291) );
  INV_X1 U2579 ( .A(n4076), .ZN(n2289) );
  NAND2_X1 U2580 ( .A1(n3179), .A2(n3172), .ZN(n4048) );
  NOR2_X1 U2581 ( .A1(n3073), .A2(n2866), .ZN(n3006) );
  NOR2_X1 U2582 ( .A1(n2978), .A2(n4377), .ZN(n2272) );
  NAND2_X1 U2583 ( .A1(n2347), .A2(n2295), .ZN(n2297) );
  INV_X1 U2584 ( .A(n2297), .ZN(n2294) );
  INV_X1 U2585 ( .A(IR_REG_13__SCAN_IN), .ZN(n2385) );
  NAND2_X1 U2586 ( .A1(n3020), .A2(n2368), .ZN(n2359) );
  NOR2_X1 U2587 ( .A1(n2675), .A2(n2346), .ZN(n2345) );
  INV_X1 U2588 ( .A(n3445), .ZN(n2346) );
  INV_X1 U2589 ( .A(n3422), .ZN(n2324) );
  NAND2_X1 U2590 ( .A1(n3136), .A2(n3035), .ZN(n2457) );
  NAND2_X1 U2591 ( .A1(n2823), .A2(n2822), .ZN(n2364) );
  OR2_X1 U2592 ( .A1(n3915), .A2(n2366), .ZN(n2365) );
  INV_X1 U2593 ( .A(n2820), .ZN(n2366) );
  XNOR2_X1 U2594 ( .A(n2526), .B(n3038), .ZN(n2527) );
  OR2_X1 U2595 ( .A1(n3083), .A2(n3005), .ZN(n3133) );
  AND2_X1 U2596 ( .A1(n2871), .A2(n3074), .ZN(n2891) );
  AND2_X1 U2597 ( .A1(n4675), .A2(n4046), .ZN(n3080) );
  INV_X1 U2598 ( .A(n2949), .ZN(n3001) );
  NAND2_X1 U2599 ( .A1(n2485), .A2(n2486), .ZN(n2329) );
  NAND2_X1 U2600 ( .A1(n2996), .A2(REG2_REG_3__SCAN_IN), .ZN(n2484) );
  INV_X1 U2601 ( .A(n2311), .ZN(n3121) );
  NAND2_X1 U2602 ( .A1(n3219), .A2(n3218), .ZN(n3220) );
  OR2_X1 U2603 ( .A1(n3217), .A2(n3114), .ZN(n3218) );
  NAND2_X1 U2604 ( .A1(n4760), .A2(n3211), .ZN(n3212) );
  INV_X1 U2605 ( .A(n3391), .ZN(n2307) );
  OR2_X1 U2606 ( .A1(n3228), .A2(n3227), .ZN(n3392) );
  NAND2_X1 U2607 ( .A1(n3384), .A2(n3385), .ZN(n3386) );
  NAND2_X1 U2608 ( .A1(n2300), .A2(n2299), .ZN(n4790) );
  NAND2_X1 U2609 ( .A1(n4176), .A2(n2301), .ZN(n2299) );
  OR2_X1 U2610 ( .A1(n4782), .A2(n2259), .ZN(n2300) );
  INV_X1 U2611 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3944) );
  NAND2_X1 U2612 ( .A1(n4189), .A2(n4188), .ZN(n4191) );
  NAND2_X1 U2613 ( .A1(n4677), .A2(REG2_REG_11__SCAN_IN), .ZN(n4188) );
  OAI21_X1 U2614 ( .B1(n4797), .B2(n4794), .A(n2314), .ZN(n4194) );
  OR2_X1 U2615 ( .A1(n4193), .A2(REG2_REG_13__SCAN_IN), .ZN(n2314) );
  NAND2_X1 U2616 ( .A1(n4829), .A2(n4198), .ZN(n4689) );
  NAND2_X1 U2617 ( .A1(n4826), .A2(n4181), .ZN(n4182) );
  AND2_X1 U2618 ( .A1(n4035), .A2(n4034), .ZN(n4222) );
  INV_X1 U2619 ( .A(n4266), .ZN(n4042) );
  NAND2_X1 U2620 ( .A1(n4358), .A2(n4336), .ZN(n2933) );
  OR2_X1 U2621 ( .A1(n4126), .A2(n4377), .ZN(n2928) );
  AND2_X1 U2622 ( .A1(n2699), .A2(REG3_REG_16__SCAN_IN), .ZN(n2725) );
  OR2_X1 U2623 ( .A1(n3357), .A2(n3423), .ZN(n2374) );
  OAI21_X1 U2624 ( .B1(n3306), .B2(n2966), .A(n4067), .ZN(n3356) );
  AND3_X1 U2625 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2531) );
  OAI21_X1 U2626 ( .B1(n3271), .B2(n3263), .A(n4071), .ZN(n3325) );
  INV_X1 U2627 ( .A(n3199), .ZN(n3179) );
  NAND2_X1 U2628 ( .A1(n2956), .A2(n4695), .ZN(n4523) );
  NOR2_X1 U2629 ( .A1(n3006), .A2(n3133), .ZN(n3148) );
  NAND2_X1 U2630 ( .A1(n2443), .A2(n2442), .ZN(n4874) );
  NOR2_X1 U2631 ( .A1(n4272), .A2(n4249), .ZN(n4248) );
  NAND2_X1 U2632 ( .A1(n4248), .A2(n4217), .ZN(n4224) );
  NOR2_X1 U2633 ( .A1(n4361), .A2(n4336), .ZN(n4335) );
  AND2_X1 U2634 ( .A1(n2347), .A2(n2387), .ZN(n2298) );
  INV_X1 U2635 ( .A(IR_REG_20__SCAN_IN), .ZN(n2415) );
  NAND2_X1 U2636 ( .A1(n2440), .A2(IR_REG_31__SCAN_IN), .ZN(n2416) );
  INV_X1 U2637 ( .A(IR_REG_9__SCAN_IN), .ZN(n2595) );
  CLKBUF_X1 U2638 ( .A(n2521), .Z(n2522) );
  AND2_X1 U2639 ( .A1(n2879), .A2(n2947), .ZN(n4252) );
  INV_X1 U2640 ( .A(n4682), .ZN(n2432) );
  NAND2_X1 U2641 ( .A1(n2955), .A2(n2954), .ZN(n4243) );
  NAND2_X1 U2642 ( .A1(n4142), .A2(n4150), .ZN(n4141) );
  NAND2_X1 U2643 ( .A1(n4702), .A2(REG1_REG_3__SCAN_IN), .ZN(n4701) );
  NAND2_X1 U2644 ( .A1(n4761), .A2(n4762), .ZN(n4760) );
  XNOR2_X1 U2645 ( .A(n3212), .B(n4920), .ZN(n4770) );
  NAND2_X1 U2646 ( .A1(n4770), .A2(REG2_REG_8__SCAN_IN), .ZN(n4769) );
  XNOR2_X1 U2647 ( .A(n4191), .B(n4916), .ZN(n4787) );
  NAND2_X1 U2648 ( .A1(n4787), .A2(REG2_REG_12__SCAN_IN), .ZN(n4786) );
  NAND2_X1 U2649 ( .A1(n4684), .A2(n2310), .ZN(n4841) );
  NAND2_X1 U2650 ( .A1(n2268), .A2(n4597), .ZN(n2310) );
  NOR2_X1 U2651 ( .A1(n4841), .A2(n4840), .ZN(n4842) );
  OAI21_X1 U2652 ( .B1(n2316), .B2(n4844), .A(n2373), .ZN(n2315) );
  NAND2_X1 U2653 ( .A1(n2317), .A2(n4833), .ZN(n2316) );
  NAND2_X1 U2654 ( .A1(n4845), .A2(n4846), .ZN(n2317) );
  INV_X1 U2655 ( .A(n4835), .ZN(n4839) );
  NOR2_X1 U2656 ( .A1(n4842), .A2(n2309), .ZN(n2308) );
  AND2_X1 U2657 ( .A1(n4847), .A2(REG1_REG_18__SCAN_IN), .ZN(n2309) );
  INV_X1 U2658 ( .A(n4695), .ZN(n4685) );
  NAND2_X1 U2659 ( .A1(n2440), .A2(n2439), .ZN(n4695) );
  OR2_X1 U2660 ( .A1(n2438), .A2(n2437), .ZN(n2439) );
  AOI21_X1 U2661 ( .B1(n2341), .B2(n2236), .A(n2340), .ZN(n2339) );
  INV_X1 U2662 ( .A(n2345), .ZN(n2340) );
  INV_X1 U2663 ( .A(n2342), .ZN(n2341) );
  OAI21_X1 U2664 ( .B1(n2674), .B2(n2236), .A(n3511), .ZN(n2342) );
  INV_X1 U2665 ( .A(n4079), .ZN(n2293) );
  INV_X1 U2666 ( .A(n4063), .ZN(n2290) );
  NAND2_X1 U2667 ( .A1(n2265), .A2(n2264), .ZN(n3103) );
  NAND2_X1 U2668 ( .A1(n4141), .A2(n2248), .ZN(n2264) );
  NAND2_X1 U2669 ( .A1(n2263), .A2(n2318), .ZN(n2265) );
  NAND2_X1 U2670 ( .A1(n4703), .A2(n3104), .ZN(n3105) );
  OR2_X1 U2671 ( .A1(n3103), .A2(n3120), .ZN(n3104) );
  AND2_X1 U2672 ( .A1(n4174), .A2(n4173), .ZN(n4175) );
  NOR2_X1 U2673 ( .A1(n4816), .A2(n2319), .ZN(n4197) );
  AND2_X1 U2674 ( .A1(n4910), .A2(REG2_REG_15__SCAN_IN), .ZN(n2319) );
  NOR2_X1 U2675 ( .A1(n4091), .A2(n2278), .ZN(n2277) );
  NOR2_X1 U2676 ( .A1(n4307), .A2(n3011), .ZN(n2273) );
  NOR2_X1 U2677 ( .A1(n3475), .A2(n4515), .ZN(n2270) );
  OAI21_X1 U2678 ( .B1(n4024), .B2(n4043), .A(n2959), .ZN(n3238) );
  NAND2_X1 U2679 ( .A1(n2349), .A2(n2388), .ZN(n2348) );
  INV_X1 U2680 ( .A(IR_REG_25__SCAN_IN), .ZN(n2349) );
  INV_X1 U2681 ( .A(IR_REG_10__SCAN_IN), .ZN(n2380) );
  INV_X1 U2682 ( .A(IR_REG_7__SCAN_IN), .ZN(n2590) );
  INV_X1 U2683 ( .A(IR_REG_5__SCAN_IN), .ZN(n2378) );
  AND2_X1 U2684 ( .A1(n2837), .A2(n2836), .ZN(n2878) );
  INV_X1 U2685 ( .A(IR_REG_4__SCAN_IN), .ZN(n3781) );
  INV_X1 U2686 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3863) );
  INV_X1 U2687 ( .A(REG3_REG_19__SCAN_IN), .ZN(n3872) );
  NAND2_X1 U2688 ( .A1(n3915), .A2(n2818), .ZN(n2367) );
  INV_X1 U2689 ( .A(n3035), .ZN(n2843) );
  XNOR2_X1 U2690 ( .A(n2330), .B(n3038), .ZN(n2493) );
  NAND2_X1 U2691 ( .A1(n2332), .A2(n2331), .ZN(n2330) );
  CLKBUF_X1 U2692 ( .A(n3410), .Z(n3411) );
  INV_X1 U2693 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2582) );
  OR2_X1 U2694 ( .A1(n2583), .A2(n2582), .ZN(n2602) );
  OR2_X1 U2695 ( .A1(n3059), .A2(n4979), .ZN(n2370) );
  INV_X1 U2696 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3952) );
  NAND2_X2 U2697 ( .A1(n2429), .A2(n2428), .ZN(n2504) );
  NAND2_X1 U2698 ( .A1(n2426), .A2(n2425), .ZN(n2429) );
  OR2_X1 U2699 ( .A1(n2874), .A2(n2424), .ZN(n2426) );
  INV_X1 U2700 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2742) );
  OR2_X1 U2701 ( .A1(n2743), .A2(n2742), .ZN(n2753) );
  AND3_X1 U2702 ( .A1(n3492), .A2(n3491), .A3(n3490), .ZN(n4009) );
  NAND2_X1 U2703 ( .A1(n4152), .A2(n2247), .ZN(n2311) );
  XNOR2_X1 U2704 ( .A(n3103), .B(n4705), .ZN(n4704) );
  NAND2_X1 U2705 ( .A1(n4704), .A2(REG2_REG_3__SCAN_IN), .ZN(n4703) );
  NAND2_X1 U2706 ( .A1(n2262), .A2(n2261), .ZN(n3209) );
  OAI21_X1 U2707 ( .B1(n3208), .B2(REG2_REG_5__SCAN_IN), .A(n4679), .ZN(n2262)
         );
  NAND2_X1 U2708 ( .A1(n3208), .A2(REG2_REG_5__SCAN_IN), .ZN(n2261) );
  NAND2_X1 U2709 ( .A1(n2303), .A2(n2302), .ZN(n3223) );
  NAND2_X1 U2710 ( .A1(n4922), .A2(n2550), .ZN(n2302) );
  NAND2_X1 U2711 ( .A1(n4747), .A2(n2238), .ZN(n2303) );
  NOR2_X1 U2712 ( .A1(n4773), .A2(n3394), .ZN(n3398) );
  OR2_X1 U2713 ( .A1(n3398), .A2(n3397), .ZN(n4174) );
  XNOR2_X1 U2714 ( .A(n4175), .B(n4916), .ZN(n4782) );
  NOR2_X1 U2715 ( .A1(n4782), .A2(n2642), .ZN(n4781) );
  NOR2_X1 U2716 ( .A1(n4790), .A2(n2371), .ZN(n4177) );
  NOR2_X1 U2717 ( .A1(n4813), .A2(n2312), .ZN(n4180) );
  AND2_X1 U2718 ( .A1(n4910), .A2(REG1_REG_15__SCAN_IN), .ZN(n2312) );
  XNOR2_X1 U2719 ( .A(n4197), .B(n2710), .ZN(n4831) );
  NAND2_X1 U2720 ( .A1(n2267), .A2(n2266), .ZN(n4845) );
  NAND2_X1 U2721 ( .A1(n4689), .A2(n4688), .ZN(n2266) );
  OAI21_X1 U2722 ( .B1(n4689), .B2(n4688), .A(n2268), .ZN(n2267) );
  NOR2_X1 U2723 ( .A1(n4224), .A2(n4225), .ZN(n4539) );
  NAND2_X1 U2724 ( .A1(n2282), .A2(n2285), .ZN(n4210) );
  AOI21_X1 U2725 ( .B1(n4206), .B2(n3993), .A(n3994), .ZN(n2285) );
  NOR2_X1 U2726 ( .A1(n2284), .A2(n4208), .ZN(n2283) );
  INV_X1 U2727 ( .A(n3990), .ZN(n4225) );
  OR2_X1 U2728 ( .A1(n2947), .A2(n2946), .ZN(n4205) );
  INV_X1 U2729 ( .A(n2286), .ZN(n4241) );
  NOR2_X1 U2730 ( .A1(n4357), .A2(n4378), .ZN(n2930) );
  NAND2_X1 U2731 ( .A1(n2982), .A2(n4093), .ZN(n4355) );
  NAND2_X1 U2732 ( .A1(n4374), .A2(n4090), .ZN(n2982) );
  AND2_X1 U2733 ( .A1(n2764), .A2(REG3_REG_20__SCAN_IN), .ZN(n2776) );
  NOR2_X1 U2734 ( .A1(n2753), .A2(n3872), .ZN(n2764) );
  OR2_X1 U2735 ( .A1(n4402), .A2(n4713), .ZN(n2926) );
  NAND2_X1 U2736 ( .A1(n4459), .A2(n4088), .ZN(n4434) );
  NAND2_X1 U2737 ( .A1(n2281), .A2(n2279), .ZN(n4479) );
  NOR2_X1 U2738 ( .A1(n4481), .A2(n2280), .ZN(n2279) );
  INV_X1 U2739 ( .A(n3976), .ZN(n2280) );
  NAND2_X1 U2740 ( .A1(n2281), .A2(n3976), .ZN(n4482) );
  NOR2_X1 U2741 ( .A1(n2688), .A2(n2687), .ZN(n2699) );
  OR2_X1 U2742 ( .A1(n2654), .A2(n3944), .ZN(n2688) );
  INV_X1 U2743 ( .A(n4477), .ZN(n4474) );
  NOR2_X1 U2744 ( .A1(n4500), .A2(n4474), .ZN(n4473) );
  AND2_X1 U2745 ( .A1(n3976), .A2(n3972), .ZN(n4491) );
  OR2_X1 U2746 ( .A1(n2602), .A2(n3414), .ZN(n2620) );
  AND2_X1 U2747 ( .A1(n3470), .A2(n2970), .ZN(n4856) );
  NAND2_X1 U2748 ( .A1(n3356), .A2(n4064), .ZN(n2968) );
  INV_X1 U2749 ( .A(n4876), .ZN(n4865) );
  INV_X1 U2750 ( .A(n4519), .ZN(n4863) );
  NAND2_X1 U2751 ( .A1(n2964), .A2(n4059), .ZN(n3306) );
  OAI21_X1 U2752 ( .B1(n3294), .B2(n2963), .A(n4057), .ZN(n3271) );
  NAND2_X1 U2753 ( .A1(n3059), .A2(n2870), .ZN(n3083) );
  INV_X1 U2754 ( .A(n4904), .ZN(n2870) );
  AND2_X1 U2755 ( .A1(n4053), .A2(n4050), .ZN(n4022) );
  NAND2_X1 U2756 ( .A1(n4673), .A2(n3080), .ZN(n4519) );
  NOR2_X1 U2757 ( .A1(n3183), .A2(n3202), .ZN(n3292) );
  INV_X1 U2758 ( .A(n3237), .ZN(n4020) );
  CLKBUF_X1 U2759 ( .A(n2957), .Z(n4024) );
  AND2_X1 U2760 ( .A1(n3156), .A2(n4875), .ZN(n3247) );
  INV_X1 U2761 ( .A(n2899), .ZN(n4879) );
  INV_X1 U2762 ( .A(n4516), .ZN(n4878) );
  INV_X1 U2763 ( .A(n3136), .ZN(n4875) );
  INV_X1 U2764 ( .A(n4858), .ZN(n4543) );
  NAND2_X1 U2765 ( .A1(n2273), .A2(n4264), .ZN(n4272) );
  INV_X1 U2766 ( .A(n2273), .ZN(n4288) );
  AND2_X1 U2767 ( .A1(n4335), .A2(n2934), .ZN(n4326) );
  NAND2_X1 U2768 ( .A1(n4425), .A2(n2241), .ZN(n4361) );
  NAND2_X1 U2769 ( .A1(n4425), .A2(n2272), .ZN(n4384) );
  AND2_X1 U2770 ( .A1(n4425), .A2(n4407), .ZN(n4405) );
  NAND2_X1 U2771 ( .A1(n4473), .A2(n4453), .ZN(n4454) );
  OR2_X1 U2772 ( .A1(n4454), .A2(n4442), .ZN(n4444) );
  NAND2_X1 U2773 ( .A1(n2270), .A2(n3513), .ZN(n4500) );
  INV_X1 U2774 ( .A(n4515), .ZN(n4525) );
  INV_X1 U2775 ( .A(n2270), .ZN(n4524) );
  AND2_X1 U2776 ( .A1(n3364), .A2(n2252), .ZN(n4869) );
  NAND2_X1 U2777 ( .A1(n3364), .A2(n2235), .ZN(n3436) );
  INV_X1 U2778 ( .A(n2967), .ZN(n3363) );
  NOR2_X1 U2779 ( .A1(n3331), .A2(n3312), .ZN(n3364) );
  NAND2_X1 U2780 ( .A1(n4523), .A2(n4941), .ZN(n4968) );
  NOR2_X1 U2781 ( .A1(n3266), .A2(n3273), .ZN(n3332) );
  NAND2_X1 U2782 ( .A1(n3332), .A2(n2271), .ZN(n3331) );
  INV_X1 U2783 ( .A(n4968), .ZN(n4952) );
  INV_X1 U2784 ( .A(n4971), .ZN(n4965) );
  OR2_X1 U2785 ( .A1(n4881), .A2(n4675), .ZN(n4941) );
  AND2_X1 U2786 ( .A1(n3148), .A2(n3008), .ZN(n3014) );
  INV_X1 U2787 ( .A(n3083), .ZN(n3074) );
  XNOR2_X1 U2788 ( .A(n2876), .B(IR_REG_28__SCAN_IN), .ZN(n3108) );
  NAND2_X1 U2789 ( .A1(n2407), .A2(n2406), .ZN(n2856) );
  INV_X1 U2790 ( .A(n2405), .ZN(n2407) );
  XNOR2_X1 U2791 ( .A(n2869), .B(n2868), .ZN(n3082) );
  INV_X1 U2792 ( .A(IR_REG_19__SCAN_IN), .ZN(n2437) );
  AND2_X1 U2793 ( .A1(n2386), .A2(n2385), .ZN(n2337) );
  NOR2_X1 U2794 ( .A1(n2521), .A2(n2384), .ZN(n2660) );
  NOR2_X1 U2795 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2487)
         );
  NAND2_X1 U2796 ( .A1(n2325), .A2(n3281), .ZN(n3499) );
  NAND2_X1 U2797 ( .A1(n2354), .A2(n2358), .ZN(n2353) );
  NAND2_X1 U2798 ( .A1(n2360), .A2(n2359), .ZN(n2358) );
  NAND2_X1 U2799 ( .A1(n2639), .A2(n2345), .ZN(n2344) );
  CLKBUF_X1 U2800 ( .A(n3877), .Z(n3881) );
  NAND2_X1 U2801 ( .A1(n2581), .A2(n2580), .ZN(n3421) );
  INV_X1 U2802 ( .A(n3515), .ZN(n3963) );
  OAI22_X1 U2803 ( .A1(n3877), .A2(n2789), .B1(n2788), .B2(n2787), .ZN(n3950)
         );
  NAND2_X1 U2804 ( .A1(n2616), .A2(n2618), .ZN(n2619) );
  NAND2_X1 U2805 ( .A1(n2460), .A2(n2462), .ZN(n2463) );
  INV_X1 U2806 ( .A(n3514), .ZN(n4724) );
  INV_X1 U2807 ( .A(n4711), .ZN(n3515) );
  OR2_X1 U2808 ( .A1(n2877), .A2(n3108), .ZN(n3514) );
  CLKBUF_X1 U2809 ( .A(n3279), .Z(n3280) );
  INV_X1 U2810 ( .A(n4728), .ZN(n3955) );
  NAND2_X1 U2811 ( .A1(n2891), .A2(n2873), .ZN(n4719) );
  INV_X1 U2812 ( .A(n4719), .ZN(n3968) );
  NAND2_X1 U2813 ( .A1(n2884), .A2(n2883), .ZN(n4266) );
  NAND2_X1 U2814 ( .A1(n2828), .A2(n2827), .ZN(n4302) );
  OAI211_X1 U2815 ( .C1(n4305), .C2(n3001), .A(n2815), .B(n2814), .ZN(n4321)
         );
  NAND4_X1 U2816 ( .A1(n2518), .A2(n2517), .A3(n2516), .A4(n2515), .ZN(n4131)
         );
  NOR2_X1 U2817 ( .A1(n2243), .A2(n2329), .ZN(n2334) );
  NAND2_X1 U2818 ( .A1(n2496), .A2(REG3_REG_2__SCAN_IN), .ZN(n2471) );
  OR2_X2 U2819 ( .A1(n3059), .A2(n4904), .ZN(n4134) );
  AND2_X1 U2820 ( .A1(n3097), .A2(n3096), .ZN(n4739) );
  OAI21_X1 U2821 ( .B1(n4682), .B2(n3116), .A(n3115), .ZN(n4139) );
  NAND2_X1 U2822 ( .A1(n4682), .A2(n3116), .ZN(n3115) );
  NAND2_X1 U2823 ( .A1(n4156), .A2(n4157), .ZN(n4155) );
  NAND2_X1 U2824 ( .A1(n4141), .A2(n3102), .ZN(n4156) );
  XNOR2_X1 U2825 ( .A(n2311), .B(n3120), .ZN(n4702) );
  OAI22_X1 U2826 ( .A1(n4167), .A2(n3125), .B1(n3124), .B2(n3123), .ZN(n3126)
         );
  NAND2_X1 U2827 ( .A1(n3126), .A2(n3127), .ZN(n3219) );
  XNOR2_X1 U2828 ( .A(n3209), .B(n4924), .ZN(n4750) );
  NAND2_X1 U2829 ( .A1(n4750), .A2(REG2_REG_6__SCAN_IN), .ZN(n4749) );
  XNOR2_X1 U2830 ( .A(n3220), .B(n4924), .ZN(n4748) );
  NAND2_X1 U2831 ( .A1(n4747), .A2(n3221), .ZN(n4756) );
  XNOR2_X1 U2832 ( .A(n3223), .B(n4920), .ZN(n4766) );
  NOR2_X1 U2833 ( .A1(n4766), .A2(n2568), .ZN(n4765) );
  NAND2_X1 U2834 ( .A1(n4769), .A2(n3213), .ZN(n3216) );
  NAND2_X1 U2835 ( .A1(n3216), .A2(n3215), .ZN(n3384) );
  NAND2_X1 U2836 ( .A1(n2307), .A2(n4917), .ZN(n2306) );
  NOR2_X1 U2837 ( .A1(n4917), .A2(n2307), .ZN(n2305) );
  NOR2_X1 U2838 ( .A1(n4774), .A2(n2604), .ZN(n4773) );
  NAND2_X1 U2839 ( .A1(n4786), .A2(n4192), .ZN(n4797) );
  XNOR2_X1 U2840 ( .A(n4194), .B(n2313), .ZN(n4805) );
  XNOR2_X1 U2841 ( .A(n4180), .B(n2710), .ZN(n4828) );
  NAND2_X1 U2842 ( .A1(n4828), .A2(n4827), .ZN(n4826) );
  AND2_X1 U2843 ( .A1(n4739), .A2(n4149), .ZN(n4835) );
  OR2_X1 U2844 ( .A1(n4218), .A2(n4217), .ZN(n4219) );
  AND2_X1 U2845 ( .A1(n4530), .A2(n3265), .ZN(n4431) );
  OR2_X1 U2846 ( .A1(n3083), .A2(n3007), .ZN(n4528) );
  AND2_X1 U2847 ( .A1(n3315), .A2(n4971), .ZN(n4871) );
  INV_X1 U2848 ( .A(n4528), .ZN(n4883) );
  INV_X1 U2849 ( .A(n4990), .ZN(n4988) );
  XNOR2_X1 U2850 ( .A(n3494), .B(n4540), .ZN(n4730) );
  AND2_X2 U2851 ( .A1(n3014), .A2(n3146), .ZN(n4978) );
  NAND2_X1 U2852 ( .A1(n3074), .A2(n3073), .ZN(n4903) );
  OR2_X1 U2853 ( .A1(n2422), .A2(n2681), .ZN(n2411) );
  NAND2_X1 U2854 ( .A1(n3082), .A2(STATE_REG_SCAN_IN), .ZN(n4904) );
  XNOR2_X1 U2855 ( .A(n2436), .B(IR_REG_22__SCAN_IN), .ZN(n4675) );
  NAND2_X1 U2856 ( .A1(n2418), .A2(IR_REG_31__SCAN_IN), .ZN(n2419) );
  INV_X1 U2857 ( .A(IR_REG_16__SCAN_IN), .ZN(n2708) );
  NOR2_X1 U2858 ( .A1(n2598), .A2(n2597), .ZN(n4678) );
  INV_X2 U2859 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  AOI21_X1 U2860 ( .B1(n4849), .B2(n4850), .A(n2315), .ZN(n4852) );
  XNOR2_X1 U2861 ( .A(n2308), .B(n4686), .ZN(n4699) );
  OR2_X1 U2862 ( .A1(n4232), .A2(n4618), .ZN(n3012) );
  OR2_X1 U2863 ( .A1(n4232), .A2(n4671), .ZN(n3017) );
  AND2_X1 U2864 ( .A1(n3363), .A2(n3423), .ZN(n2235) );
  XOR2_X1 U2865 ( .A(n2685), .B(n2846), .Z(n2236) );
  AND2_X1 U2866 ( .A1(n2286), .A2(n3985), .ZN(n2237) );
  INV_X1 U2867 ( .A(n3010), .ZN(n3437) );
  AND2_X1 U2868 ( .A1(n3221), .A2(n2257), .ZN(n2238) );
  AND2_X1 U2869 ( .A1(n2235), .A2(n3437), .ZN(n2239) );
  NAND2_X1 U2870 ( .A1(n2244), .A2(n2660), .ZN(n2240) );
  AND2_X1 U2871 ( .A1(n2272), .A2(n4362), .ZN(n2241) );
  OR2_X1 U2872 ( .A1(n2435), .A2(IR_REG_22__SCAN_IN), .ZN(n2242) );
  AND2_X1 U2873 ( .A1(n2413), .A2(n2387), .ZN(n2417) );
  NOR2_X1 U2874 ( .A1(n2482), .A2(n2483), .ZN(n2243) );
  AND2_X1 U2875 ( .A1(n2337), .A2(n2336), .ZN(n2244) );
  AND2_X1 U2876 ( .A1(n2502), .A2(n2491), .ZN(n4705) );
  NOR2_X1 U2877 ( .A1(n2435), .A2(n2350), .ZN(n2403) );
  AND2_X1 U2878 ( .A1(n3392), .A2(n3391), .ZN(n2245) );
  AND2_X1 U2879 ( .A1(n2560), .A2(n3281), .ZN(n2246) );
  NAND2_X1 U2880 ( .A1(n4681), .A2(REG1_REG_2__SCAN_IN), .ZN(n2247) );
  AND2_X1 U2881 ( .A1(n2318), .A2(n3102), .ZN(n2248) );
  INV_X1 U2882 ( .A(n4870), .ZN(n4859) );
  NAND2_X1 U2883 ( .A1(n4681), .A2(REG2_REG_2__SCAN_IN), .ZN(n2318) );
  AND2_X1 U2884 ( .A1(n4862), .A2(n3010), .ZN(n2249) );
  OR2_X1 U2885 ( .A1(n3857), .A2(n2820), .ZN(n2250) );
  AND2_X1 U2886 ( .A1(n2409), .A2(n2868), .ZN(n2251) );
  INV_X1 U2887 ( .A(IR_REG_3__SCAN_IN), .ZN(n2322) );
  AND2_X1 U2888 ( .A1(n2239), .A2(n4859), .ZN(n2252) );
  OR2_X1 U2889 ( .A1(n2341), .A2(n2343), .ZN(n2253) );
  INV_X1 U2890 ( .A(IR_REG_27__SCAN_IN), .ZN(n2424) );
  INV_X1 U2891 ( .A(n2714), .ZN(n2634) );
  NAND2_X1 U2892 ( .A1(n2639), .A2(n3445), .ZN(n3460) );
  OR2_X1 U2893 ( .A1(n3860), .A2(n3859), .ZN(n2254) );
  INV_X1 U2894 ( .A(n2714), .ZN(n2832) );
  AND2_X1 U2895 ( .A1(n2660), .A2(n2385), .ZN(n2680) );
  INV_X1 U2896 ( .A(n3326), .ZN(n2271) );
  INV_X1 U2897 ( .A(n2363), .ZN(n2362) );
  NAND2_X1 U2898 ( .A1(n2365), .A2(n2364), .ZN(n2363) );
  NAND2_X1 U2899 ( .A1(n2344), .A2(n2674), .ZN(n3510) );
  AND3_X1 U2900 ( .A1(n3048), .A2(n3047), .A3(n3968), .ZN(n2255) );
  INV_X1 U2901 ( .A(n3888), .ZN(n2361) );
  NOR2_X1 U2902 ( .A1(n4781), .A2(n4176), .ZN(n2256) );
  NAND2_X1 U2903 ( .A1(n4754), .A2(REG1_REG_7__SCAN_IN), .ZN(n2257) );
  INV_X1 U2904 ( .A(n3019), .ZN(n2360) );
  OR2_X1 U2905 ( .A1(n3019), .A2(n2361), .ZN(n2258) );
  INV_X1 U2906 ( .A(n3889), .ZN(n2368) );
  INV_X1 U2907 ( .A(n4348), .ZN(n4125) );
  AND3_X1 U2908 ( .A1(n2806), .A2(n2805), .A3(n2804), .ZN(n4348) );
  AND2_X2 U2909 ( .A1(n3149), .A2(n4528), .ZN(n4888) );
  INV_X1 U2910 ( .A(n4888), .ZN(n4457) );
  XNOR2_X1 U2911 ( .A(n2411), .B(IR_REG_26__SCAN_IN), .ZN(n2854) );
  INV_X1 U2912 ( .A(n4345), .ZN(n4336) );
  NAND2_X1 U2913 ( .A1(n3364), .A2(n3363), .ZN(n3362) );
  INV_X1 U2914 ( .A(n4088), .ZN(n2278) );
  NAND2_X1 U2915 ( .A1(n2233), .A2(DATAI_20_), .ZN(n4385) );
  NAND2_X1 U2916 ( .A1(n3364), .A2(n2239), .ZN(n2269) );
  INV_X1 U2917 ( .A(n4791), .ZN(n2301) );
  OR2_X1 U2918 ( .A1(n4791), .A2(n2642), .ZN(n2259) );
  NAND2_X1 U2919 ( .A1(n2660), .A2(n2337), .ZN(n2731) );
  INV_X1 U2920 ( .A(n4362), .ZN(n4357) );
  NAND2_X1 U2921 ( .A1(n2233), .A2(DATAI_21_), .ZN(n4362) );
  INV_X1 U2922 ( .A(n4809), .ZN(n2313) );
  OAI22_X1 U2923 ( .A1(n4166), .A2(n3107), .B1(n3106), .B2(n3123), .ZN(n3208)
         );
  AND2_X1 U2924 ( .A1(n4739), .A2(n3109), .ZN(n4833) );
  NOR2_X1 U2925 ( .A1(n4117), .A2(n3162), .ZN(n2260) );
  INV_X1 U2926 ( .A(n4690), .ZN(n2268) );
  INV_X1 U2927 ( .A(IR_REG_30__SCAN_IN), .ZN(n2390) );
  OAI21_X1 U2928 ( .B1(n3870), .B2(n3871), .A(n2763), .ZN(n3924) );
  AOI22_X2 U2929 ( .A1(n2724), .A2(n2723), .B1(n2722), .B2(n2721), .ZN(n3908)
         );
  NOR2_X4 U2930 ( .A1(n3858), .A2(n2254), .ZN(n3857) );
  OAI21_X1 U2931 ( .B1(n2327), .B2(n2243), .A(n2326), .ZN(n2331) );
  NOR2_X1 U2932 ( .A1(n2856), .A2(n2852), .ZN(n2412) );
  NAND2_X1 U2933 ( .A1(n3279), .A2(n3282), .ZN(n2325) );
  INV_X1 U2934 ( .A(n2355), .ZN(n3887) );
  AOI21_X1 U2935 ( .B1(n3253), .B2(n3252), .A(n2530), .ZN(n3279) );
  AOI21_X1 U2936 ( .B1(n3887), .B2(n3888), .A(n3889), .ZN(n3021) );
  NAND2_X2 U2937 ( .A1(n2412), .A2(n2854), .ZN(n2452) );
  NAND2_X1 U2938 ( .A1(n4831), .A2(n4830), .ZN(n4829) );
  INV_X1 U2939 ( .A(n2384), .ZN(n2274) );
  NAND2_X1 U2940 ( .A1(n2274), .A2(n2335), .ZN(n2276) );
  AND2_X2 U2941 ( .A1(n2244), .A2(n2275), .ZN(n2413) );
  NAND2_X1 U2942 ( .A1(n4459), .A2(n2277), .ZN(n4374) );
  NAND2_X1 U2943 ( .A1(n4492), .A2(n4491), .ZN(n2281) );
  NAND2_X1 U2944 ( .A1(n2993), .A2(n2287), .ZN(n2286) );
  NAND2_X1 U2945 ( .A1(n2993), .A2(n2283), .ZN(n2282) );
  NAND2_X1 U2946 ( .A1(n2993), .A2(n2992), .ZN(n4240) );
  NAND2_X1 U2947 ( .A1(n2962), .A2(n4053), .ZN(n3294) );
  OAI21_X1 U2948 ( .B1(n3372), .B2(n2291), .A(n2288), .ZN(n3468) );
  OAI21_X1 U2949 ( .B1(n3372), .B2(n4077), .A(n4063), .ZN(n3430) );
  AOI21_X1 U2950 ( .B1(n4077), .B2(n4063), .A(n2293), .ZN(n2292) );
  NAND2_X1 U2951 ( .A1(n2413), .A2(n2294), .ZN(n2393) );
  MUX2_X1 U2953 ( .A(REG2_REG_1__SCAN_IN), .B(n3101), .S(n4682), .Z(n4142) );
  NAND2_X1 U2954 ( .A1(n3392), .A2(n2305), .ZN(n2304) );
  OAI211_X1 U2955 ( .C1(n3392), .C2(n3393), .A(n2304), .B(n2306), .ZN(n4774)
         );
  INV_X1 U2956 ( .A(n2519), .ZN(n2379) );
  NAND3_X1 U2957 ( .A1(n2321), .A2(n2320), .A3(n2322), .ZN(n2519) );
  NAND2_X1 U2958 ( .A1(n3410), .A2(n2615), .ZN(n3409) );
  NAND2_X1 U2959 ( .A1(n2581), .A2(n2323), .ZN(n3410) );
  AND2_X1 U2960 ( .A1(n2580), .A2(n2324), .ZN(n2323) );
  INV_X1 U2961 ( .A(n2484), .ZN(n2333) );
  NAND2_X1 U2962 ( .A1(n2492), .A2(n2328), .ZN(n2327) );
  NAND2_X1 U2963 ( .A1(n2333), .A2(n2714), .ZN(n2332) );
  NAND2_X1 U2964 ( .A1(n2639), .A2(n2339), .ZN(n2338) );
  NAND2_X1 U2965 ( .A1(n2338), .A2(n2253), .ZN(n2716) );
  NAND2_X1 U2966 ( .A1(n2417), .A2(n2388), .ZN(n2435) );
  INV_X1 U2967 ( .A(n2352), .ZN(n3034) );
  AOI21_X1 U2968 ( .B1(n3857), .B2(n2367), .A(n2363), .ZN(n2355) );
  OAI21_X1 U2969 ( .B1(n3857), .B2(n2823), .A(n2822), .ZN(n3914) );
  MUX2_X2 U2970 ( .A(n3016), .B(n3015), .S(n4978), .Z(n3018) );
  NAND2_X1 U2971 ( .A1(n2957), .A2(n3151), .ZN(n3153) );
  NAND2_X1 U2972 ( .A1(n2959), .A2(n4044), .ZN(n2957) );
  MUX2_X2 U2973 ( .A(n3835), .B(n3015), .S(n4990), .Z(n3013) );
  INV_X1 U2974 ( .A(n2422), .ZN(n2406) );
  NAND2_X1 U2975 ( .A1(n4326), .A2(n4308), .ZN(n4307) );
  CLKBUF_X1 U2976 ( .A(n3233), .Z(n3236) );
  AND2_X1 U2977 ( .A1(n4043), .A2(n4045), .ZN(n4882) );
  NAND2_X1 U2978 ( .A1(n2504), .A2(DATAI_0_), .ZN(n2445) );
  OR2_X1 U2979 ( .A1(n2504), .A2(n2444), .ZN(n2446) );
  NAND2_X1 U2980 ( .A1(n2504), .A2(DATAI_1_), .ZN(n2431) );
  AND2_X1 U2981 ( .A1(n2233), .A2(DATAI_30_), .ZN(n4544) );
  AND2_X1 U2982 ( .A1(n2233), .A2(DATAI_31_), .ZN(n4008) );
  NAND2_X1 U2983 ( .A1(n2233), .A2(DATAI_28_), .ZN(n4217) );
  NAND2_X1 U2984 ( .A1(n2233), .A2(DATAI_26_), .ZN(n4264) );
  NAND2_X1 U2985 ( .A1(n2233), .A2(DATAI_25_), .ZN(n4289) );
  NAND2_X1 U2986 ( .A1(n2233), .A2(DATAI_24_), .ZN(n4308) );
  NAND2_X1 U2987 ( .A1(n2233), .A2(DATAI_22_), .ZN(n4345) );
  AOI21_X2 U2988 ( .B1(n4257), .B2(n2942), .A(n2941), .ZN(n4238) );
  OAI21_X2 U2989 ( .B1(n4855), .B2(n4856), .A(n2916), .ZN(n3474) );
  AND2_X1 U2990 ( .A1(n4380), .A2(n4407), .ZN(n2369) );
  AND2_X1 U2991 ( .A1(n4193), .A2(REG1_REG_13__SCAN_IN), .ZN(n2371) );
  INV_X1 U2992 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3119) );
  AND2_X1 U2993 ( .A1(n2233), .A2(DATAI_23_), .ZN(n4320) );
  NAND2_X1 U2994 ( .A1(n2969), .A2(n3437), .ZN(n2372) );
  NAND2_X1 U2995 ( .A1(n4848), .A2(n4847), .ZN(n2373) );
  INV_X1 U2996 ( .A(REG1_REG_1__SCAN_IN), .ZN(n3116) );
  OR2_X1 U2997 ( .A1(n4478), .A2(n4453), .ZN(n2375) );
  NAND2_X1 U2998 ( .A1(n2819), .A2(n2818), .ZN(n2820) );
  OR2_X1 U2999 ( .A1(n2983), .A2(n4362), .ZN(n2376) );
  INV_X1 U3000 ( .A(IR_REG_0__SCAN_IN), .ZN(n2444) );
  OR2_X1 U3001 ( .A1(n4400), .A2(n4385), .ZN(n2377) );
  INV_X1 U3002 ( .A(n4358), .ZN(n2932) );
  INV_X1 U3003 ( .A(n3498), .ZN(n2560) );
  OR2_X1 U3004 ( .A1(n4280), .A2(n4098), .ZN(n2993) );
  INV_X1 U3005 ( .A(IR_REG_26__SCAN_IN), .ZN(n2421) );
  NAND2_X1 U3006 ( .A1(n2466), .A2(REG2_REG_2__SCAN_IN), .ZN(n2467) );
  INV_X1 U3007 ( .A(n4320), .ZN(n2934) );
  INV_X1 U3008 ( .A(IR_REG_28__SCAN_IN), .ZN(n2427) );
  OR2_X1 U3009 ( .A1(n2667), .A2(n2668), .ZN(n2675) );
  OR2_X1 U3010 ( .A1(n2762), .A2(n2761), .ZN(n2763) );
  INV_X1 U3011 ( .A(n2617), .ZN(n2618) );
  OR2_X1 U3012 ( .A1(n2802), .A2(n3863), .ZN(n2811) );
  NAND2_X1 U3013 ( .A1(n4681), .A2(n3119), .ZN(n3118) );
  INV_X1 U3014 ( .A(n4917), .ZN(n3393) );
  OR2_X1 U3015 ( .A1(n4243), .A2(n4217), .ZN(n4207) );
  NOR2_X1 U3016 ( .A1(n4348), .A2(n2934), .ZN(n2935) );
  AND2_X1 U3017 ( .A1(n4723), .A2(n4442), .ZN(n2923) );
  OR2_X1 U3018 ( .A1(n4127), .A2(n4515), .ZN(n2918) );
  OR2_X1 U3019 ( .A1(n4129), .A2(n4870), .ZN(n2916) );
  AND2_X1 U3020 ( .A1(n2233), .A2(DATAI_27_), .ZN(n4249) );
  AND2_X1 U3021 ( .A1(n3108), .A2(n3080), .ZN(n4516) );
  INV_X1 U3022 ( .A(n3857), .ZN(n3862) );
  XNOR2_X1 U3023 ( .A(n2493), .B(n2494), .ZN(n3198) );
  NAND2_X1 U3024 ( .A1(n2776), .A2(REG3_REG_21__SCAN_IN), .ZN(n2790) );
  INV_X1 U3025 ( .A(n4462), .ZN(n4453) );
  INV_X1 U3026 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3917) );
  OR2_X1 U3027 ( .A1(n2790), .A2(n3952), .ZN(n2802) );
  AND2_X1 U3028 ( .A1(n2892), .A2(n4528), .ZN(n3953) );
  AND2_X1 U3029 ( .A1(n4205), .A2(n2948), .ZN(n4230) );
  AND2_X1 U3030 ( .A1(n2233), .A2(n3081), .ZN(n3096) );
  OAI21_X1 U3031 ( .B1(n4681), .B2(n3119), .A(n3118), .ZN(n4154) );
  INV_X1 U3032 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3414) );
  INV_X1 U3033 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3695) );
  INV_X1 U3034 ( .A(n4737), .ZN(n4149) );
  NOR2_X1 U3035 ( .A1(n2620), .A2(n3695), .ZN(n2640) );
  INV_X1 U3036 ( .A(n4264), .ZN(n4270) );
  INV_X1 U3037 ( .A(n2971), .ZN(n3476) );
  INV_X1 U3038 ( .A(IR_REG_11__SCAN_IN), .ZN(n2628) );
  INV_X1 U3040 ( .A(n3953), .ZN(n4712) );
  OR2_X1 U3041 ( .A1(n2878), .A2(n2838), .ZN(n2885) );
  AND2_X1 U3042 ( .A1(n4739), .A2(n3108), .ZN(n4848) );
  AOI21_X1 U3043 ( .B1(n2931), .B2(n2376), .A(n2930), .ZN(n4334) );
  OR2_X1 U3044 ( .A1(n4007), .A2(n4006), .ZN(n4513) );
  NAND2_X1 U3045 ( .A1(n2994), .A2(n4001), .ZN(n4876) );
  AND2_X1 U3046 ( .A1(n4056), .A2(n4071), .ZN(n4021) );
  OAI22_X1 U3047 ( .A1(n3073), .A2(D_REG_0__SCAN_IN), .B1(n2854), .B2(n3077), 
        .ZN(n3146) );
  NAND2_X1 U3048 ( .A1(n2855), .A2(n2854), .ZN(n3073) );
  AND2_X1 U3049 ( .A1(n2573), .A2(n2556), .ZN(n4754) );
  AND2_X1 U3050 ( .A1(n3084), .A2(n3097), .ZN(n4825) );
  AND2_X1 U3051 ( .A1(n2896), .A2(n2895), .ZN(n2897) );
  INV_X1 U3052 ( .A(n4009), .ZN(n4124) );
  INV_X1 U3053 ( .A(n4848), .ZN(n4838) );
  INV_X1 U3054 ( .A(n4825), .ZN(n4853) );
  INV_X1 U3055 ( .A(n4431), .ZN(n4506) );
  INV_X1 U3056 ( .A(n4871), .ZN(n4503) );
  NAND2_X1 U3057 ( .A1(n4990), .A2(n4971), .ZN(n4618) );
  AND2_X2 U3058 ( .A1(n3014), .A2(n3009), .ZN(n4990) );
  NAND2_X1 U3059 ( .A1(n4978), .A2(n4971), .ZN(n4671) );
  INV_X1 U3060 ( .A(n4978), .ZN(n4976) );
  INV_X1 U3061 ( .A(n4903), .ZN(n4902) );
  INV_X1 U3062 ( .A(n3108), .ZN(n4673) );
  AND2_X1 U3063 ( .A1(n2630), .A2(n2647), .ZN(n4677) );
  NAND2_X1 U3064 ( .A1(n2379), .A2(n2378), .ZN(n2521) );
  NOR2_X1 U3065 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2383)
         );
  NOR2_X1 U3066 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2382)
         );
  NOR2_X1 U3067 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2381)
         );
  NAND4_X1 U3068 ( .A1(n2383), .A2(n2382), .A3(n2381), .A4(n2380), .ZN(n2384)
         );
  XNOR2_X2 U3069 ( .A(n2391), .B(n2390), .ZN(n3070) );
  INV_X1 U3070 ( .A(n2392), .ZN(n3485) );
  NAND2_X1 U3071 ( .A1(n2393), .A2(IR_REG_31__SCAN_IN), .ZN(n2394) );
  NOR2_X2 U3072 ( .A1(n3070), .A2(n3065), .ZN(n2466) );
  NAND2_X1 U3073 ( .A1(n2466), .A2(REG2_REG_1__SCAN_IN), .ZN(n2397) );
  NOR2_X1 U3074 ( .A1(n3070), .A2(n2399), .ZN(n2447) );
  NAND2_X1 U3075 ( .A1(n2447), .A2(REG3_REG_1__SCAN_IN), .ZN(n2396) );
  INV_X1 U3076 ( .A(n2482), .ZN(n2398) );
  NAND2_X1 U3077 ( .A1(n2398), .A2(REG1_REG_1__SCAN_IN), .ZN(n2401) );
  NAND2_X1 U3078 ( .A1(n2465), .A2(REG0_REG_1__SCAN_IN), .ZN(n2400) );
  NOR2_X1 U3079 ( .A1(n2403), .A2(n2681), .ZN(n2404) );
  MUX2_X1 U3080 ( .A(n2681), .B(n2404), .S(IR_REG_25__SCAN_IN), .Z(n2405) );
  NAND2_X1 U3081 ( .A1(n2869), .A2(n2868), .ZN(n2408) );
  INV_X1 U3082 ( .A(n2413), .ZN(n2414) );
  INV_X1 U3083 ( .A(n2417), .ZN(n2418) );
  INV_X1 U3084 ( .A(n3162), .ZN(n2420) );
  NAND2_X1 U3085 ( .A1(n2899), .A2(n2714), .ZN(n2434) );
  NAND2_X1 U3086 ( .A1(n2422), .A2(n2421), .ZN(n2423) );
  NAND2_X2 U3087 ( .A1(n2423), .A2(IR_REG_31__SCAN_IN), .ZN(n2874) );
  NAND2_X1 U3088 ( .A1(n2874), .A2(n2427), .ZN(n2425) );
  NAND2_X1 U3089 ( .A1(n2427), .A2(IR_REG_27__SCAN_IN), .ZN(n2428) );
  NAND2_X1 U3090 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2430)
         );
  OAI21_X2 U3091 ( .B1(n2504), .B2(n2432), .A(n2431), .ZN(n3141) );
  AND2_X4 U3092 ( .A1(n2452), .A2(n3162), .ZN(n3035) );
  NAND2_X1 U3093 ( .A1(n3141), .A2(n3035), .ZN(n2433) );
  NAND2_X1 U3094 ( .A1(n2434), .A2(n2433), .ZN(n2441) );
  NAND2_X1 U3095 ( .A1(n2435), .A2(IR_REG_31__SCAN_IN), .ZN(n2436) );
  NAND2_X1 U3096 ( .A1(n4675), .A2(n4695), .ZN(n4117) );
  INV_X1 U3097 ( .A(n4675), .ZN(n2443) );
  INV_X1 U3098 ( .A(n4046), .ZN(n2442) );
  AND2_X2 U3099 ( .A1(n3035), .A2(n4965), .ZN(n2508) );
  AOI22_X1 U3100 ( .A1(n2899), .A2(n2508), .B1(n3141), .B2(n2714), .ZN(n2461)
         );
  XNOR2_X1 U3101 ( .A(n2460), .B(n2461), .ZN(n3140) );
  NAND2_X1 U3102 ( .A1(n2950), .A2(REG2_REG_0__SCAN_IN), .ZN(n2451) );
  NAND2_X1 U3103 ( .A1(n2465), .A2(REG0_REG_0__SCAN_IN), .ZN(n2450) );
  NAND2_X1 U3104 ( .A1(n2496), .A2(REG3_REG_0__SCAN_IN), .ZN(n2449) );
  INV_X1 U3105 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4979) );
  OR2_X1 U3106 ( .A1(n2482), .A2(n4979), .ZN(n2448) );
  NAND2_X1 U3107 ( .A1(n2234), .A2(n2714), .ZN(n2453) );
  NAND3_X1 U3108 ( .A1(n2457), .A2(n2453), .A3(n2370), .ZN(n3131) );
  NOR2_X1 U3109 ( .A1(n3059), .A2(n2444), .ZN(n2454) );
  AOI21_X1 U3110 ( .B1(n3136), .B2(n2714), .A(n2454), .ZN(n2456) );
  NAND2_X1 U3111 ( .A1(n2234), .A2(n2508), .ZN(n2455) );
  NAND2_X1 U3112 ( .A1(n2456), .A2(n2455), .ZN(n3132) );
  NAND2_X1 U3113 ( .A1(n3131), .A2(n3132), .ZN(n2459) );
  NAND2_X1 U3114 ( .A1(n2457), .A2(n2846), .ZN(n2458) );
  NAND2_X1 U3115 ( .A1(n2459), .A2(n2458), .ZN(n3139) );
  NAND2_X1 U3116 ( .A1(n3140), .A2(n3139), .ZN(n2464) );
  INV_X1 U3117 ( .A(n2461), .ZN(n2462) );
  NAND2_X1 U3118 ( .A1(n2464), .A2(n2463), .ZN(n3167) );
  INV_X1 U3119 ( .A(n3167), .ZN(n2480) );
  NAND2_X1 U3120 ( .A1(n2465), .A2(REG0_REG_2__SCAN_IN), .ZN(n2468) );
  NAND2_X1 U3121 ( .A1(n2468), .A2(n2467), .ZN(n2470) );
  NAND2_X2 U3122 ( .A1(n2472), .A2(n2471), .ZN(n3199) );
  OR2_X1 U3123 ( .A1(n2487), .A2(n2681), .ZN(n2473) );
  XNOR2_X2 U3124 ( .A(n2473), .B(IR_REG_2__SCAN_IN), .ZN(n4681) );
  MUX2_X1 U3125 ( .A(n4681), .B(DATAI_2_), .S(n2504), .Z(n3172) );
  AOI22_X1 U3126 ( .A1(n3199), .A2(n2508), .B1(n3172), .B2(n4119), .ZN(n2478)
         );
  NAND2_X1 U3127 ( .A1(n3199), .A2(n2714), .ZN(n2475) );
  NAND2_X1 U3128 ( .A1(n3172), .A2(n3035), .ZN(n2474) );
  NAND2_X1 U3129 ( .A1(n2475), .A2(n2474), .ZN(n2476) );
  XNOR2_X1 U3130 ( .A(n2476), .B(n2846), .ZN(n2477) );
  NAND2_X1 U3131 ( .A1(n2477), .A2(n2478), .ZN(n2481) );
  OAI21_X1 U3132 ( .B1(n2478), .B2(n2477), .A(n2481), .ZN(n3168) );
  INV_X1 U3133 ( .A(n3168), .ZN(n2479) );
  NAND2_X1 U3134 ( .A1(n2480), .A2(n2479), .ZN(n3169) );
  NAND2_X1 U3135 ( .A1(n3169), .A2(n2481), .ZN(n3197) );
  NAND2_X1 U3136 ( .A1(n2496), .A2(n3201), .ZN(n2486) );
  NAND2_X1 U3137 ( .A1(n2465), .A2(REG0_REG_3__SCAN_IN), .ZN(n2485) );
  INV_X1 U3138 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2483) );
  INV_X1 U3139 ( .A(IR_REG_2__SCAN_IN), .ZN(n2488) );
  NAND2_X1 U3140 ( .A1(n2487), .A2(n2488), .ZN(n2489) );
  NAND2_X1 U3141 ( .A1(n2489), .A2(IR_REG_31__SCAN_IN), .ZN(n2490) );
  NAND2_X1 U3142 ( .A1(n2490), .A2(n2322), .ZN(n2502) );
  OR2_X1 U3143 ( .A1(n2490), .A2(n2322), .ZN(n2491) );
  MUX2_X1 U3144 ( .A(n4705), .B(DATAI_3_), .S(n2504), .Z(n3202) );
  NAND2_X1 U3145 ( .A1(n3202), .A2(n3035), .ZN(n2492) );
  AOI22_X1 U3146 ( .A1(n4132), .A2(n3040), .B1(n3202), .B2(n4119), .ZN(n2494)
         );
  NAND2_X1 U3147 ( .A1(n3197), .A2(n3198), .ZN(n3189) );
  INV_X1 U31480 ( .A(n2493), .ZN(n2495) );
  NAND2_X1 U31490 ( .A1(n2495), .A2(n2494), .ZN(n3191) );
  NAND2_X1 U3150 ( .A1(n2465), .A2(REG0_REG_4__SCAN_IN), .ZN(n2501) );
  INV_X1 U3151 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2497) );
  XNOR2_X1 U3152 ( .A(n2497), .B(REG3_REG_3__SCAN_IN), .ZN(n3302) );
  NAND2_X1 U3153 ( .A1(n2496), .A2(n3302), .ZN(n2500) );
  NAND2_X1 U3154 ( .A1(n2950), .A2(REG2_REG_4__SCAN_IN), .ZN(n2499) );
  INV_X1 U3155 ( .A(REG1_REG_4__SCAN_IN), .ZN(n3125) );
  OR2_X1 U3156 ( .A1(n2482), .A2(n3125), .ZN(n2498) );
  NAND2_X1 U3157 ( .A1(n3200), .A2(n2714), .ZN(n2506) );
  NAND2_X1 U3158 ( .A1(n2502), .A2(IR_REG_31__SCAN_IN), .ZN(n2503) );
  XNOR2_X1 U3159 ( .A(n2503), .B(IR_REG_4__SCAN_IN), .ZN(n4680) );
  MUX2_X1 U3160 ( .A(n4680), .B(DATAI_4_), .S(n2943), .Z(n3295) );
  NAND2_X1 U3161 ( .A1(n3295), .A2(n3035), .ZN(n2505) );
  NAND2_X1 U3162 ( .A1(n2506), .A2(n2505), .ZN(n2507) );
  XNOR2_X1 U3163 ( .A(n2507), .B(n3038), .ZN(n2512) );
  AOI22_X1 U3164 ( .A1(n3200), .A2(n3040), .B1(n3295), .B2(n4119), .ZN(n2510)
         );
  XNOR2_X1 U3165 ( .A(n2512), .B(n2510), .ZN(n3190) );
  AND2_X1 U3166 ( .A1(n3191), .A2(n3190), .ZN(n2509) );
  NAND2_X1 U3167 ( .A1(n3189), .A2(n2509), .ZN(n3188) );
  INV_X1 U3168 ( .A(n2510), .ZN(n2511) );
  NAND2_X1 U3169 ( .A1(n2512), .A2(n2511), .ZN(n2513) );
  NAND2_X1 U3170 ( .A1(n3188), .A2(n2513), .ZN(n3253) );
  NAND2_X1 U3171 ( .A1(n2996), .A2(REG2_REG_5__SCAN_IN), .ZN(n2518) );
  AOI21_X1 U3172 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        REG3_REG_5__SCAN_IN), .ZN(n2514) );
  NOR2_X1 U3173 ( .A1(n2514), .A2(n2531), .ZN(n3267) );
  NAND2_X1 U3174 ( .A1(n2496), .A2(n3267), .ZN(n2517) );
  NAND2_X1 U3175 ( .A1(n2465), .A2(REG0_REG_5__SCAN_IN), .ZN(n2516) );
  INV_X1 U3176 ( .A(REG1_REG_5__SCAN_IN), .ZN(n3114) );
  OR2_X1 U3177 ( .A1(n3489), .A2(n3114), .ZN(n2515) );
  NAND2_X1 U3178 ( .A1(n4131), .A2(n2714), .ZN(n2525) );
  NAND2_X1 U3179 ( .A1(n2519), .A2(IR_REG_31__SCAN_IN), .ZN(n2520) );
  MUX2_X1 U3180 ( .A(IR_REG_31__SCAN_IN), .B(n2520), .S(IR_REG_5__SCAN_IN), 
        .Z(n2523) );
  AND2_X1 U3181 ( .A1(n2523), .A2(n2522), .ZN(n4679) );
  MUX2_X1 U3182 ( .A(n4679), .B(DATAI_5_), .S(n2233), .Z(n3273) );
  NAND2_X1 U3183 ( .A1(n3273), .A2(n3035), .ZN(n2524) );
  NAND2_X1 U3184 ( .A1(n2525), .A2(n2524), .ZN(n2526) );
  AOI22_X1 U3185 ( .A1(n4131), .A2(n3040), .B1(n3273), .B2(n4119), .ZN(n2528)
         );
  XNOR2_X1 U3186 ( .A(n2527), .B(n2528), .ZN(n3252) );
  INV_X1 U3187 ( .A(n2527), .ZN(n2529) );
  NOR2_X1 U3188 ( .A1(n2529), .A2(n2528), .ZN(n2530) );
  NAND2_X1 U3189 ( .A1(n2465), .A2(REG0_REG_6__SCAN_IN), .ZN(n2536) );
  NAND2_X1 U3190 ( .A1(n2531), .A2(REG3_REG_6__SCAN_IN), .ZN(n2548) );
  OAI21_X1 U3191 ( .B1(n2531), .B2(REG3_REG_6__SCAN_IN), .A(n2548), .ZN(n3340)
         );
  INV_X1 U3192 ( .A(n3340), .ZN(n3288) );
  NAND2_X1 U3193 ( .A1(n2949), .A2(n3288), .ZN(n2535) );
  NAND2_X1 U3194 ( .A1(n2996), .A2(REG2_REG_6__SCAN_IN), .ZN(n2534) );
  INV_X1 U3195 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2532) );
  OR2_X1 U3196 ( .A1(n3489), .A2(n2532), .ZN(n2533) );
  NAND4_X1 U3197 ( .A1(n2536), .A2(n2535), .A3(n2534), .A4(n2533), .ZN(n3503)
         );
  NAND2_X1 U3198 ( .A1(n3503), .A2(n2714), .ZN(n2539) );
  NAND2_X1 U3199 ( .A1(n2522), .A2(IR_REG_31__SCAN_IN), .ZN(n2537) );
  XNOR2_X1 U3200 ( .A(n2537), .B(IR_REG_6__SCAN_IN), .ZN(n4746) );
  MUX2_X1 U3201 ( .A(n4746), .B(DATAI_6_), .S(n2233), .Z(n3326) );
  NAND2_X1 U3202 ( .A1(n3326), .A2(n3035), .ZN(n2538) );
  NAND2_X1 U3203 ( .A1(n2539), .A2(n2538), .ZN(n2540) );
  XNOR2_X1 U3204 ( .A(n2540), .B(n3038), .ZN(n2543) );
  NAND2_X1 U3205 ( .A1(n3503), .A2(n3040), .ZN(n2542) );
  NAND2_X1 U3206 ( .A1(n3326), .A2(n2714), .ZN(n2541) );
  NAND2_X1 U3207 ( .A1(n2542), .A2(n2541), .ZN(n2544) );
  NAND2_X1 U3208 ( .A1(n2543), .A2(n2544), .ZN(n3282) );
  INV_X1 U3209 ( .A(n2543), .ZN(n2546) );
  INV_X1 U32100 ( .A(n2544), .ZN(n2545) );
  NAND2_X1 U32110 ( .A1(n2546), .A2(n2545), .ZN(n3281) );
  NAND2_X1 U32120 ( .A1(n2465), .A2(REG0_REG_7__SCAN_IN), .ZN(n2554) );
  INV_X1 U32130 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2547) );
  NOR2_X1 U32140 ( .A1(n2548), .A2(n2547), .ZN(n2566) );
  AND2_X1 U32150 ( .A1(n2548), .A2(n2547), .ZN(n2549) );
  NOR2_X1 U32160 ( .A1(n2566), .A2(n2549), .ZN(n3506) );
  NAND2_X1 U32170 ( .A1(n2949), .A2(n3506), .ZN(n2553) );
  NAND2_X1 U32180 ( .A1(n2996), .A2(REG2_REG_7__SCAN_IN), .ZN(n2552) );
  INV_X1 U32190 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2550) );
  OR2_X1 U32200 ( .A1(n3489), .A2(n2550), .ZN(n2551) );
  NAND4_X1 U32210 ( .A1(n2554), .A2(n2553), .A3(n2552), .A4(n2551), .ZN(n4130)
         );
  NAND2_X1 U32220 ( .A1(n4130), .A2(n2714), .ZN(n2558) );
  OAI21_X1 U32230 ( .B1(n2522), .B2(IR_REG_6__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2555) );
  NAND2_X1 U32240 ( .A1(n2555), .A2(n2590), .ZN(n2573) );
  OR2_X1 U32250 ( .A1(n2555), .A2(n2590), .ZN(n2556) );
  MUX2_X1 U32260 ( .A(n4754), .B(DATAI_7_), .S(n2233), .Z(n3312) );
  NAND2_X1 U32270 ( .A1(n3312), .A2(n3035), .ZN(n2557) );
  NAND2_X1 U32280 ( .A1(n2558), .A2(n2557), .ZN(n2559) );
  XNOR2_X1 U32290 ( .A(n2559), .B(n2846), .ZN(n2561) );
  AOI22_X1 U32300 ( .A1(n4130), .A2(n3040), .B1(n3312), .B2(n4119), .ZN(n2562)
         );
  XNOR2_X1 U32310 ( .A(n2561), .B(n2562), .ZN(n3498) );
  INV_X1 U32320 ( .A(n2561), .ZN(n2564) );
  INV_X1 U32330 ( .A(n2562), .ZN(n2563) );
  NAND2_X1 U32340 ( .A1(n2564), .A2(n2563), .ZN(n2565) );
  NAND2_X1 U32350 ( .A1(n2996), .A2(REG2_REG_8__SCAN_IN), .ZN(n2572) );
  NAND2_X1 U32360 ( .A1(n2566), .A2(REG3_REG_8__SCAN_IN), .ZN(n2583) );
  OR2_X1 U32370 ( .A1(n2566), .A2(REG3_REG_8__SCAN_IN), .ZN(n2567) );
  AND2_X1 U32380 ( .A1(n2583), .A2(n2567), .ZN(n3366) );
  NAND2_X1 U32390 ( .A1(n2949), .A2(n3366), .ZN(n2571) );
  NAND2_X1 U32400 ( .A1(n2465), .A2(REG0_REG_8__SCAN_IN), .ZN(n2570) );
  INV_X1 U32410 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2568) );
  OR2_X1 U32420 ( .A1(n3489), .A2(n2568), .ZN(n2569) );
  NAND4_X1 U32430 ( .A1(n2572), .A2(n2571), .A3(n2570), .A4(n2569), .ZN(n3502)
         );
  NAND2_X1 U32440 ( .A1(n3502), .A2(n2508), .ZN(n2576) );
  NAND2_X1 U32450 ( .A1(n2573), .A2(IR_REG_31__SCAN_IN), .ZN(n2574) );
  XNOR2_X1 U32460 ( .A(n2574), .B(IR_REG_8__SCAN_IN), .ZN(n3222) );
  MUX2_X1 U32470 ( .A(n3222), .B(DATAI_8_), .S(n2233), .Z(n2967) );
  NAND2_X1 U32480 ( .A1(n2967), .A2(n2714), .ZN(n2575) );
  NAND2_X1 U32490 ( .A1(n2576), .A2(n2575), .ZN(n3349) );
  NAND2_X1 U32500 ( .A1(n3502), .A2(n4119), .ZN(n2578) );
  NAND2_X1 U32510 ( .A1(n2967), .A2(n3035), .ZN(n2577) );
  NAND2_X1 U32520 ( .A1(n2578), .A2(n2577), .ZN(n2579) );
  XNOR2_X1 U32530 ( .A(n2579), .B(n3038), .ZN(n3348) );
  OAI21_X1 U32540 ( .B1(n3347), .B2(n3349), .A(n3348), .ZN(n2581) );
  NAND2_X1 U32550 ( .A1(n3347), .A2(n3349), .ZN(n2580) );
  NAND2_X1 U32560 ( .A1(n3487), .A2(REG0_REG_9__SCAN_IN), .ZN(n2589) );
  NAND2_X1 U32570 ( .A1(n2583), .A2(n2582), .ZN(n2584) );
  AND2_X1 U32580 ( .A1(n2602), .A2(n2584), .ZN(n3426) );
  NAND2_X1 U32590 ( .A1(n2949), .A2(n3426), .ZN(n2588) );
  NAND2_X1 U32600 ( .A1(n2996), .A2(REG2_REG_9__SCAN_IN), .ZN(n2587) );
  INV_X1 U32610 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2585) );
  OR2_X1 U32620 ( .A1(n3489), .A2(n2585), .ZN(n2586) );
  NAND4_X1 U32630 ( .A1(n2589), .A2(n2588), .A3(n2587), .A4(n2586), .ZN(n3432)
         );
  NAND2_X1 U32640 ( .A1(n3432), .A2(n4119), .ZN(n2600) );
  INV_X1 U32650 ( .A(IR_REG_6__SCAN_IN), .ZN(n2592) );
  INV_X1 U32660 ( .A(IR_REG_8__SCAN_IN), .ZN(n2591) );
  NAND3_X1 U32670 ( .A1(n2592), .A2(n2591), .A3(n2590), .ZN(n2593) );
  NOR2_X1 U32680 ( .A1(n2522), .A2(n2593), .ZN(n2596) );
  NOR2_X1 U32690 ( .A1(n2596), .A2(n2681), .ZN(n2594) );
  MUX2_X1 U32700 ( .A(n2681), .B(n2594), .S(IR_REG_9__SCAN_IN), .Z(n2598) );
  NAND2_X1 U32710 ( .A1(n2596), .A2(n2595), .ZN(n2626) );
  INV_X1 U32720 ( .A(n2626), .ZN(n2597) );
  MUX2_X1 U32730 ( .A(n4678), .B(DATAI_9_), .S(n2233), .Z(n3373) );
  NAND2_X1 U32740 ( .A1(n3373), .A2(n3035), .ZN(n2599) );
  NAND2_X1 U32750 ( .A1(n2600), .A2(n2599), .ZN(n2601) );
  XNOR2_X1 U32760 ( .A(n2601), .B(n2846), .ZN(n2614) );
  AOI22_X1 U32770 ( .A1(n3432), .A2(n3040), .B1(n3373), .B2(n4119), .ZN(n2613)
         );
  XNOR2_X1 U32780 ( .A(n2614), .B(n2613), .ZN(n3422) );
  NAND2_X1 U32790 ( .A1(n2996), .A2(REG2_REG_10__SCAN_IN), .ZN(n2608) );
  NAND2_X1 U32800 ( .A1(n2602), .A2(n3414), .ZN(n2603) );
  AND2_X1 U32810 ( .A1(n2620), .A2(n2603), .ZN(n3439) );
  NAND2_X1 U32820 ( .A1(n2949), .A2(n3439), .ZN(n2607) );
  NAND2_X1 U32830 ( .A1(n3487), .A2(REG0_REG_10__SCAN_IN), .ZN(n2606) );
  INV_X1 U32840 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2604) );
  OR2_X1 U32850 ( .A1(n3489), .A2(n2604), .ZN(n2605) );
  NAND4_X1 U32860 ( .A1(n2608), .A2(n2607), .A3(n2606), .A4(n2605), .ZN(n4862)
         );
  NAND2_X1 U32870 ( .A1(n4862), .A2(n2714), .ZN(n2611) );
  NAND2_X1 U32880 ( .A1(n2626), .A2(IR_REG_31__SCAN_IN), .ZN(n2609) );
  XNOR2_X1 U32890 ( .A(n2609), .B(IR_REG_10__SCAN_IN), .ZN(n4917) );
  MUX2_X1 U32900 ( .A(n4917), .B(DATAI_10_), .S(n2233), .Z(n3010) );
  NAND2_X1 U32910 ( .A1(n3010), .A2(n3035), .ZN(n2610) );
  NAND2_X1 U32920 ( .A1(n2611), .A2(n2610), .ZN(n2612) );
  XNOR2_X1 U32930 ( .A(n2612), .B(n3038), .ZN(n2616) );
  AOI22_X1 U32940 ( .A1(n4862), .A2(n3040), .B1(n3010), .B2(n4119), .ZN(n2617)
         );
  XNOR2_X1 U32950 ( .A(n2616), .B(n2617), .ZN(n3412) );
  NAND2_X1 U32960 ( .A1(n2614), .A2(n2613), .ZN(n3413) );
  AND2_X1 U32970 ( .A1(n3412), .A2(n3413), .ZN(n2615) );
  NAND2_X1 U32980 ( .A1(n3409), .A2(n2619), .ZN(n3446) );
  AND2_X1 U32990 ( .A1(n2620), .A2(n3695), .ZN(n2621) );
  NOR2_X1 U33000 ( .A1(n2640), .A2(n2621), .ZN(n4868) );
  NAND2_X1 U33010 ( .A1(n2949), .A2(n4868), .ZN(n2625) );
  NAND2_X1 U33020 ( .A1(n3487), .A2(REG0_REG_11__SCAN_IN), .ZN(n2624) );
  NAND2_X1 U33030 ( .A1(n2996), .A2(REG2_REG_11__SCAN_IN), .ZN(n2623) );
  INV_X1 U33040 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3395) );
  OR2_X1 U33050 ( .A1(n3489), .A2(n3395), .ZN(n2622) );
  NAND4_X1 U33060 ( .A1(n2625), .A2(n2624), .A3(n2623), .A4(n2622), .ZN(n4129)
         );
  NAND2_X1 U33070 ( .A1(n4129), .A2(n4119), .ZN(n2632) );
  OR2_X1 U33080 ( .A1(n2626), .A2(IR_REG_10__SCAN_IN), .ZN(n2627) );
  NAND2_X1 U33090 ( .A1(n2627), .A2(IR_REG_31__SCAN_IN), .ZN(n2629) );
  OR2_X1 U33100 ( .A1(n2629), .A2(n2628), .ZN(n2630) );
  NAND2_X1 U33110 ( .A1(n2629), .A2(n2628), .ZN(n2647) );
  MUX2_X1 U33120 ( .A(n4677), .B(DATAI_11_), .S(n2233), .Z(n4870) );
  NAND2_X1 U33130 ( .A1(n4870), .A2(n3035), .ZN(n2631) );
  NAND2_X1 U33140 ( .A1(n2632), .A2(n2631), .ZN(n2633) );
  XNOR2_X1 U33150 ( .A(n2633), .B(n2846), .ZN(n2635) );
  AOI22_X1 U33160 ( .A1(n4129), .A2(n3040), .B1(n4870), .B2(n4119), .ZN(n2636)
         );
  NAND2_X1 U33170 ( .A1(n2635), .A2(n2636), .ZN(n3444) );
  INV_X1 U33180 ( .A(n2635), .ZN(n2638) );
  INV_X1 U33190 ( .A(n2636), .ZN(n2637) );
  NAND2_X1 U33200 ( .A1(n2638), .A2(n2637), .ZN(n3445) );
  NAND2_X1 U33210 ( .A1(n3487), .A2(REG0_REG_12__SCAN_IN), .ZN(n2646) );
  OR2_X1 U33220 ( .A1(n2640), .A2(REG3_REG_12__SCAN_IN), .ZN(n2641) );
  NAND2_X1 U33230 ( .A1(n2640), .A2(REG3_REG_12__SCAN_IN), .ZN(n2654) );
  AND2_X1 U33240 ( .A1(n2641), .A2(n2654), .ZN(n3478) );
  NAND2_X1 U33250 ( .A1(n2949), .A2(n3478), .ZN(n2645) );
  NAND2_X1 U33260 ( .A1(n2996), .A2(REG2_REG_12__SCAN_IN), .ZN(n2644) );
  INV_X1 U33270 ( .A(REG1_REG_12__SCAN_IN), .ZN(n2642) );
  OR2_X1 U33280 ( .A1(n3489), .A2(n2642), .ZN(n2643) );
  NAND4_X1 U33290 ( .A1(n2646), .A2(n2645), .A3(n2644), .A4(n2643), .ZN(n4128)
         );
  NAND2_X1 U33300 ( .A1(n4128), .A2(n4119), .ZN(n2650) );
  NAND2_X1 U33310 ( .A1(n2647), .A2(IR_REG_31__SCAN_IN), .ZN(n2648) );
  XNOR2_X1 U33320 ( .A(n2648), .B(IR_REG_12__SCAN_IN), .ZN(n4190) );
  MUX2_X1 U33330 ( .A(n4190), .B(DATAI_12_), .S(n2233), .Z(n2971) );
  NAND2_X1 U33340 ( .A1(n2971), .A2(n3035), .ZN(n2649) );
  NAND2_X1 U33350 ( .A1(n2650), .A2(n2649), .ZN(n2651) );
  XNOR2_X1 U33360 ( .A(n2651), .B(n3038), .ZN(n3938) );
  NAND2_X1 U33370 ( .A1(n4128), .A2(n3040), .ZN(n2653) );
  NAND2_X1 U33380 ( .A1(n2971), .A2(n4119), .ZN(n2652) );
  NAND2_X1 U33390 ( .A1(n2653), .A2(n2652), .ZN(n3937) );
  AND2_X1 U33400 ( .A1(n3938), .A2(n3937), .ZN(n2667) );
  NAND2_X1 U33410 ( .A1(n2996), .A2(REG2_REG_13__SCAN_IN), .ZN(n2659) );
  NAND2_X1 U33420 ( .A1(n2654), .A2(n3944), .ZN(n2655) );
  AND2_X1 U33430 ( .A1(n2688), .A2(n2655), .ZN(n4527) );
  NAND2_X1 U33440 ( .A1(n2949), .A2(n4527), .ZN(n2658) );
  NAND2_X1 U33450 ( .A1(n3487), .A2(REG0_REG_13__SCAN_IN), .ZN(n2657) );
  INV_X1 U33460 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4613) );
  OR2_X1 U33470 ( .A1(n3489), .A2(n4613), .ZN(n2656) );
  NAND4_X1 U33480 ( .A1(n2659), .A2(n2658), .A3(n2657), .A4(n2656), .ZN(n4127)
         );
  NAND2_X1 U33490 ( .A1(n4127), .A2(n4119), .ZN(n2663) );
  OR2_X1 U33500 ( .A1(n2660), .A2(n2681), .ZN(n2661) );
  XNOR2_X1 U33510 ( .A(n2661), .B(IR_REG_13__SCAN_IN), .ZN(n4193) );
  MUX2_X1 U33520 ( .A(n4193), .B(DATAI_13_), .S(n2233), .Z(n4515) );
  NAND2_X1 U3353 ( .A1(n4515), .A2(n3035), .ZN(n2662) );
  NAND2_X1 U33540 ( .A1(n2663), .A2(n2662), .ZN(n2664) );
  XNOR2_X1 U3355 ( .A(n2664), .B(n3038), .ZN(n2669) );
  NAND2_X1 U3356 ( .A1(n4127), .A2(n3040), .ZN(n2666) );
  NAND2_X1 U3357 ( .A1(n4515), .A2(n4119), .ZN(n2665) );
  NAND2_X1 U3358 ( .A1(n2666), .A2(n2665), .ZN(n2670) );
  AND2_X1 U3359 ( .A1(n2669), .A2(n2670), .ZN(n2668) );
  INV_X1 U3360 ( .A(n2668), .ZN(n3936) );
  INV_X1 U3361 ( .A(n3937), .ZN(n3461) );
  INV_X1 U3362 ( .A(n3938), .ZN(n3940) );
  NAND3_X1 U3363 ( .A1(n3936), .A2(n3461), .A3(n3940), .ZN(n2673) );
  INV_X1 U3364 ( .A(n2669), .ZN(n2672) );
  INV_X1 U3365 ( .A(n2670), .ZN(n2671) );
  NAND2_X1 U3366 ( .A1(n2672), .A2(n2671), .ZN(n3935) );
  AND2_X1 U3367 ( .A1(n2673), .A2(n3935), .ZN(n2674) );
  NAND2_X1 U3368 ( .A1(n3487), .A2(REG0_REG_14__SCAN_IN), .ZN(n2679) );
  XNOR2_X1 U3369 ( .A(n2688), .B(REG3_REG_14__SCAN_IN), .ZN(n4501) );
  NAND2_X1 U3370 ( .A1(n2949), .A2(n4501), .ZN(n2678) );
  NAND2_X1 U3371 ( .A1(n2996), .A2(REG2_REG_14__SCAN_IN), .ZN(n2677) );
  INV_X1 U3372 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4803) );
  OR2_X1 U3373 ( .A1(n3489), .A2(n4803), .ZN(n2676) );
  NAND4_X1 U3374 ( .A1(n2679), .A2(n2678), .A3(n2677), .A4(n2676), .ZN(n4517)
         );
  NAND2_X1 U3375 ( .A1(n4517), .A2(n4119), .ZN(n2684) );
  OR2_X1 U3376 ( .A1(n2680), .A2(n2681), .ZN(n2682) );
  XNOR2_X1 U3377 ( .A(n2682), .B(IR_REG_14__SCAN_IN), .ZN(n4809) );
  MUX2_X1 U3378 ( .A(n4809), .B(DATAI_14_), .S(n2233), .Z(n4498) );
  NAND2_X1 U3379 ( .A1(n4498), .A2(n3035), .ZN(n2683) );
  NAND2_X1 U3380 ( .A1(n2684), .A2(n2683), .ZN(n2685) );
  INV_X1 U3381 ( .A(n4517), .ZN(n2919) );
  INV_X1 U3382 ( .A(n2508), .ZN(n2808) );
  INV_X1 U3383 ( .A(n4498), .ZN(n3513) );
  OAI22_X1 U3384 ( .A1(n2919), .A2(n2808), .B1(n3513), .B2(n2832), .ZN(n3511)
         );
  NAND2_X1 U3385 ( .A1(n2996), .A2(REG2_REG_15__SCAN_IN), .ZN(n2694) );
  INV_X1 U3386 ( .A(n2688), .ZN(n2686) );
  AOI21_X1 U3387 ( .B1(n2686), .B2(REG3_REG_14__SCAN_IN), .A(
        REG3_REG_15__SCAN_IN), .ZN(n2689) );
  NAND2_X1 U3388 ( .A1(REG3_REG_14__SCAN_IN), .A2(REG3_REG_15__SCAN_IN), .ZN(
        n2687) );
  OR2_X1 U3389 ( .A1(n2689), .A2(n2699), .ZN(n4475) );
  INV_X1 U3390 ( .A(n4475), .ZN(n2690) );
  NAND2_X1 U3391 ( .A1(n2949), .A2(n2690), .ZN(n2693) );
  NAND2_X1 U3392 ( .A1(n3487), .A2(REG0_REG_15__SCAN_IN), .ZN(n2692) );
  INV_X1 U3393 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4179) );
  OR2_X1 U3394 ( .A1(n3489), .A2(n4179), .ZN(n2691) );
  NAND4_X1 U3395 ( .A1(n2694), .A2(n2693), .A3(n2692), .A4(n2691), .ZN(n4494)
         );
  INV_X1 U3396 ( .A(n4494), .ZN(n4465) );
  INV_X1 U3397 ( .A(IR_REG_14__SCAN_IN), .ZN(n2695) );
  NAND2_X1 U3398 ( .A1(n2680), .A2(n2695), .ZN(n2696) );
  NAND2_X1 U3399 ( .A1(n2696), .A2(IR_REG_31__SCAN_IN), .ZN(n2706) );
  XNOR2_X1 U3400 ( .A(n2706), .B(IR_REG_15__SCAN_IN), .ZN(n4910) );
  INV_X1 U3401 ( .A(n4910), .ZN(n4196) );
  INV_X1 U3402 ( .A(DATAI_15_), .ZN(n2697) );
  MUX2_X1 U3403 ( .A(n4196), .B(n2697), .S(n2233), .Z(n4477) );
  OAI22_X1 U3404 ( .A1(n4465), .A2(n2832), .B1(n2843), .B2(n4477), .ZN(n2698)
         );
  XOR2_X1 U3405 ( .A(n3038), .B(n2698), .Z(n2715) );
  NOR2_X1 U3406 ( .A1(n2716), .A2(n2715), .ZN(n3896) );
  NAND2_X1 U3407 ( .A1(n2996), .A2(REG2_REG_16__SCAN_IN), .ZN(n2704) );
  NOR2_X1 U3408 ( .A1(n2699), .A2(REG3_REG_16__SCAN_IN), .ZN(n2700) );
  OR2_X1 U3409 ( .A1(n2725), .A2(n2700), .ZN(n4456) );
  INV_X1 U3410 ( .A(n4456), .ZN(n3901) );
  NAND2_X1 U3411 ( .A1(n2949), .A2(n3901), .ZN(n2703) );
  NAND2_X1 U3412 ( .A1(n3487), .A2(REG0_REG_16__SCAN_IN), .ZN(n2702) );
  INV_X1 U3413 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4827) );
  OR2_X1 U3414 ( .A1(n3489), .A2(n4827), .ZN(n2701) );
  NAND4_X1 U3415 ( .A1(n2704), .A2(n2703), .A3(n2702), .A4(n2701), .ZN(n4439)
         );
  NAND2_X1 U3416 ( .A1(n4439), .A2(n4119), .ZN(n2712) );
  INV_X1 U3417 ( .A(IR_REG_15__SCAN_IN), .ZN(n2705) );
  NAND2_X1 U3418 ( .A1(n2706), .A2(n2705), .ZN(n2707) );
  NAND2_X1 U3419 ( .A1(n2707), .A2(IR_REG_31__SCAN_IN), .ZN(n2709) );
  XNOR2_X1 U3420 ( .A(n2709), .B(n2708), .ZN(n4909) );
  INV_X1 U3421 ( .A(n4909), .ZN(n2710) );
  MUX2_X1 U3422 ( .A(n2710), .B(DATAI_16_), .S(n2233), .Z(n4462) );
  NAND2_X1 U3423 ( .A1(n4462), .A2(n3035), .ZN(n2711) );
  NAND2_X1 U3424 ( .A1(n2712), .A2(n2711), .ZN(n2713) );
  XNOR2_X1 U3425 ( .A(n2713), .B(n3038), .ZN(n2719) );
  INV_X1 U3426 ( .A(n4439), .ZN(n4478) );
  OAI22_X1 U3427 ( .A1(n4478), .A2(n2808), .B1(n4453), .B2(n2832), .ZN(n2720)
         );
  XNOR2_X1 U3428 ( .A(n2719), .B(n2720), .ZN(n3897) );
  NOR2_X1 U3429 ( .A1(n3896), .A2(n3897), .ZN(n2724) );
  NAND2_X1 U3430 ( .A1(n2716), .A2(n2715), .ZN(n3959) );
  NAND2_X1 U3431 ( .A1(n4474), .A2(n2714), .ZN(n2718) );
  NAND2_X1 U3432 ( .A1(n4494), .A2(n3040), .ZN(n2717) );
  NAND2_X1 U3433 ( .A1(n2718), .A2(n2717), .ZN(n3961) );
  NAND2_X1 U3434 ( .A1(n3959), .A2(n3961), .ZN(n2723) );
  INV_X1 U3435 ( .A(n2719), .ZN(n2722) );
  INV_X1 U3436 ( .A(n2720), .ZN(n2721) );
  NAND2_X1 U3437 ( .A1(n3487), .A2(REG0_REG_17__SCAN_IN), .ZN(n2730) );
  NAND2_X1 U3438 ( .A1(n2725), .A2(REG3_REG_17__SCAN_IN), .ZN(n2743) );
  OR2_X1 U3439 ( .A1(n2725), .A2(REG3_REG_17__SCAN_IN), .ZN(n2726) );
  AND2_X1 U3440 ( .A1(n2743), .A2(n2726), .ZN(n4445) );
  NAND2_X1 U3441 ( .A1(n2496), .A2(n4445), .ZN(n2729) );
  NAND2_X1 U3442 ( .A1(n2996), .A2(REG2_REG_17__SCAN_IN), .ZN(n2728) );
  INV_X1 U3443 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4597) );
  OR2_X1 U3444 ( .A1(n3489), .A2(n4597), .ZN(n2727) );
  NAND4_X1 U3445 ( .A1(n2730), .A2(n2729), .A3(n2728), .A4(n2727), .ZN(n4723)
         );
  NAND2_X1 U3446 ( .A1(n4723), .A2(n4119), .ZN(n2735) );
  NAND2_X1 U3447 ( .A1(n2731), .A2(IR_REG_31__SCAN_IN), .ZN(n2732) );
  MUX2_X1 U3448 ( .A(IR_REG_31__SCAN_IN), .B(n2732), .S(IR_REG_17__SCAN_IN), 
        .Z(n2733) );
  AND2_X1 U3449 ( .A1(n2733), .A2(n2240), .ZN(n4690) );
  MUX2_X1 U3450 ( .A(n4690), .B(DATAI_17_), .S(n2233), .Z(n4442) );
  NAND2_X1 U3451 ( .A1(n4442), .A2(n3035), .ZN(n2734) );
  NAND2_X1 U3452 ( .A1(n2735), .A2(n2734), .ZN(n2736) );
  XNOR2_X1 U3453 ( .A(n2736), .B(n2846), .ZN(n3906) );
  NAND2_X1 U3454 ( .A1(n4723), .A2(n3040), .ZN(n2738) );
  NAND2_X1 U3455 ( .A1(n4442), .A2(n4119), .ZN(n2737) );
  AND2_X1 U3456 ( .A1(n2738), .A2(n2737), .ZN(n2739) );
  NAND2_X1 U3457 ( .A1(n3906), .A2(n2739), .ZN(n2741) );
  INV_X1 U34580 ( .A(n3906), .ZN(n2740) );
  INV_X1 U34590 ( .A(n2739), .ZN(n3905) );
  NAND2_X1 U3460 ( .A1(n2743), .A2(n2742), .ZN(n2744) );
  NAND2_X1 U3461 ( .A1(n2753), .A2(n2744), .ZN(n4727) );
  INV_X1 U3462 ( .A(n4727), .ZN(n4427) );
  NAND2_X1 U3463 ( .A1(n2949), .A2(n4427), .ZN(n2748) );
  NAND2_X1 U3464 ( .A1(n3487), .A2(REG0_REG_18__SCAN_IN), .ZN(n2747) );
  NAND2_X1 U3465 ( .A1(n2996), .A2(REG2_REG_18__SCAN_IN), .ZN(n2746) );
  INV_X1 U3466 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4683) );
  OR2_X1 U34670 ( .A1(n3489), .A2(n4683), .ZN(n2745) );
  NAND4_X1 U3468 ( .A1(n2748), .A2(n2747), .A3(n2746), .A4(n2745), .ZN(n4402)
         );
  INV_X1 U34690 ( .A(n4402), .ZN(n4437) );
  NAND2_X1 U3470 ( .A1(n2240), .A2(IR_REG_31__SCAN_IN), .ZN(n2749) );
  XNOR2_X1 U34710 ( .A(n2749), .B(IR_REG_18__SCAN_IN), .ZN(n4847) );
  MUX2_X1 U3472 ( .A(n4847), .B(DATAI_18_), .S(n2233), .Z(n4713) );
  INV_X1 U34730 ( .A(n4713), .ZN(n2925) );
  OAI22_X1 U3474 ( .A1(n4437), .A2(n2832), .B1(n2925), .B2(n2843), .ZN(n2750)
         );
  XNOR2_X1 U34750 ( .A(n2750), .B(n3038), .ZN(n2752) );
  OAI22_X1 U3476 ( .A1(n4437), .A2(n2808), .B1(n2925), .B2(n2832), .ZN(n2751)
         );
  NAND2_X1 U34770 ( .A1(n2752), .A2(n2751), .ZN(n4716) );
  NOR2_X1 U3478 ( .A1(n2752), .A2(n2751), .ZN(n4715) );
  AND2_X1 U34790 ( .A1(n2753), .A2(n3872), .ZN(n2754) );
  NOR2_X1 U3480 ( .A1(n2764), .A2(n2754), .ZN(n4408) );
  NAND2_X1 U34810 ( .A1(n2949), .A2(n4408), .ZN(n2758) );
  NAND2_X1 U3482 ( .A1(n3487), .A2(REG0_REG_19__SCAN_IN), .ZN(n2757) );
  NAND2_X1 U34830 ( .A1(n2950), .A2(REG2_REG_19__SCAN_IN), .ZN(n2756) );
  INV_X1 U3484 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4589) );
  OR2_X1 U34850 ( .A1(n3489), .A2(n4589), .ZN(n2755) );
  NAND4_X1 U3486 ( .A1(n2758), .A2(n2757), .A3(n2756), .A4(n2755), .ZN(n4710)
         );
  INV_X1 U34870 ( .A(n4710), .ZN(n4380) );
  INV_X1 U3488 ( .A(DATAI_19_), .ZN(n3061) );
  MUX2_X1 U34890 ( .A(n4695), .B(n3061), .S(n2233), .Z(n4407) );
  OAI22_X1 U3490 ( .A1(n4380), .A2(n2832), .B1(n4407), .B2(n2843), .ZN(n2759)
         );
  XNOR2_X1 U34910 ( .A(n2759), .B(n3038), .ZN(n2762) );
  NAND2_X1 U3492 ( .A1(n4710), .A2(n3040), .ZN(n2760) );
  OAI21_X1 U34930 ( .B1(n2832), .B2(n4407), .A(n2760), .ZN(n2761) );
  XNOR2_X1 U3494 ( .A(n2762), .B(n2761), .ZN(n3871) );
  NAND2_X1 U34950 ( .A1(n2996), .A2(REG2_REG_20__SCAN_IN), .ZN(n2769) );
  NOR2_X1 U3496 ( .A1(n2764), .A2(REG3_REG_20__SCAN_IN), .ZN(n2765) );
  OR2_X1 U34970 ( .A1(n2776), .A2(n2765), .ZN(n4386) );
  INV_X1 U3498 ( .A(n4386), .ZN(n3931) );
  NAND2_X1 U34990 ( .A1(n2949), .A2(n3931), .ZN(n2768) );
  NAND2_X1 U3500 ( .A1(n3487), .A2(REG0_REG_20__SCAN_IN), .ZN(n2767) );
  INV_X1 U35010 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4585) );
  OR2_X1 U3502 ( .A1(n3489), .A2(n4585), .ZN(n2766) );
  NAND4_X1 U35030 ( .A1(n2769), .A2(n2768), .A3(n2767), .A4(n2766), .ZN(n4126)
         );
  NAND2_X1 U3504 ( .A1(n4126), .A2(n4119), .ZN(n2771) );
  OR2_X1 U35050 ( .A1(n4385), .A2(n2843), .ZN(n2770) );
  NAND2_X1 U35060 ( .A1(n2771), .A2(n2770), .ZN(n2772) );
  XNOR2_X1 U35070 ( .A(n2772), .B(n2846), .ZN(n2775) );
  NOR2_X1 U35080 ( .A1(n4385), .A2(n2832), .ZN(n2773) );
  AOI21_X1 U35090 ( .B1(n4126), .B2(n3040), .A(n2773), .ZN(n2774) );
  OR2_X1 U35100 ( .A1(n2775), .A2(n2774), .ZN(n3925) );
  NAND2_X1 U35110 ( .A1(n3924), .A2(n3925), .ZN(n3923) );
  NAND2_X1 U35120 ( .A1(n2775), .A2(n2774), .ZN(n3927) );
  NAND2_X1 U35130 ( .A1(n3923), .A2(n3927), .ZN(n3877) );
  NAND2_X1 U35140 ( .A1(n2996), .A2(REG2_REG_21__SCAN_IN), .ZN(n2781) );
  OR2_X1 U35150 ( .A1(n2776), .A2(REG3_REG_21__SCAN_IN), .ZN(n2777) );
  AND2_X1 U35160 ( .A1(n2790), .A2(n2777), .ZN(n4364) );
  NAND2_X1 U35170 ( .A1(n2949), .A2(n4364), .ZN(n2780) );
  NAND2_X1 U35180 ( .A1(n3487), .A2(REG0_REG_21__SCAN_IN), .ZN(n2779) );
  INV_X1 U35190 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4580) );
  OR2_X1 U35200 ( .A1(n3489), .A2(n4580), .ZN(n2778) );
  NAND4_X1 U35210 ( .A1(n2781), .A2(n2780), .A3(n2779), .A4(n2778), .ZN(n4378)
         );
  NAND2_X1 U35220 ( .A1(n4378), .A2(n4119), .ZN(n2783) );
  OR2_X1 U35230 ( .A1(n4362), .A2(n2843), .ZN(n2782) );
  NAND2_X1 U35240 ( .A1(n2783), .A2(n2782), .ZN(n2784) );
  XNOR2_X1 U35250 ( .A(n2784), .B(n3038), .ZN(n3879) );
  NAND2_X1 U35260 ( .A1(n4378), .A2(n2508), .ZN(n2786) );
  OR2_X1 U35270 ( .A1(n4362), .A2(n2832), .ZN(n2785) );
  NAND2_X1 U35280 ( .A1(n2786), .A2(n2785), .ZN(n3878) );
  NOR2_X1 U35290 ( .A1(n3879), .A2(n3878), .ZN(n2789) );
  INV_X1 U35300 ( .A(n3879), .ZN(n2788) );
  INV_X1 U35310 ( .A(n3878), .ZN(n2787) );
  NAND2_X1 U35320 ( .A1(n3487), .A2(REG0_REG_22__SCAN_IN), .ZN(n2796) );
  NAND2_X1 U35330 ( .A1(n2790), .A2(n3952), .ZN(n2791) );
  AND2_X1 U35340 ( .A1(n2802), .A2(n2791), .ZN(n4337) );
  NAND2_X1 U35350 ( .A1(n2949), .A2(n4337), .ZN(n2795) );
  NAND2_X1 U35360 ( .A1(n2996), .A2(REG2_REG_22__SCAN_IN), .ZN(n2794) );
  INV_X1 U35370 ( .A(REG1_REG_22__SCAN_IN), .ZN(n2792) );
  OR2_X1 U35380 ( .A1(n3489), .A2(n2792), .ZN(n2793) );
  NAND4_X1 U35390 ( .A1(n2796), .A2(n2795), .A3(n2794), .A4(n2793), .ZN(n4358)
         );
  OAI22_X1 U35400 ( .A1(n2932), .A2(n2832), .B1(n4345), .B2(n2843), .ZN(n2797)
         );
  XNOR2_X1 U35410 ( .A(n2797), .B(n3038), .ZN(n2799) );
  OAI22_X1 U35420 ( .A1(n2932), .A2(n2808), .B1(n4345), .B2(n2832), .ZN(n2798)
         );
  XNOR2_X1 U35430 ( .A(n2799), .B(n2798), .ZN(n3951) );
  NOR2_X2 U35440 ( .A1(n3950), .A2(n3951), .ZN(n3858) );
  NOR2_X1 U35450 ( .A1(n2799), .A2(n2798), .ZN(n3860) );
  NAND2_X1 U35460 ( .A1(n3487), .A2(REG0_REG_23__SCAN_IN), .ZN(n2801) );
  INV_X1 U35470 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4571) );
  OR2_X1 U35480 ( .A1(n3489), .A2(n4571), .ZN(n2800) );
  AND2_X1 U35490 ( .A1(n2801), .A2(n2800), .ZN(n2806) );
  NAND2_X1 U35500 ( .A1(n2802), .A2(n3863), .ZN(n2803) );
  AND2_X1 U35510 ( .A1(n2811), .A2(n2803), .ZN(n4327) );
  NAND2_X1 U35520 ( .A1(n4327), .A2(n2949), .ZN(n2805) );
  NAND2_X1 U35530 ( .A1(n2950), .A2(REG2_REG_23__SCAN_IN), .ZN(n2804) );
  OAI22_X1 U35540 ( .A1(n4348), .A2(n2832), .B1(n2843), .B2(n2934), .ZN(n2807)
         );
  XNOR2_X1 U35550 ( .A(n2807), .B(n3038), .ZN(n2810) );
  OAI22_X1 U35560 ( .A1(n4348), .A2(n2808), .B1(n2832), .B2(n2934), .ZN(n2809)
         );
  XNOR2_X1 U35570 ( .A(n2810), .B(n2809), .ZN(n3859) );
  AND2_X1 U35580 ( .A1(n2810), .A2(n2809), .ZN(n2823) );
  INV_X1 U35590 ( .A(n2823), .ZN(n2819) );
  AND2_X1 U35600 ( .A1(n2811), .A2(n3917), .ZN(n2812) );
  OR2_X1 U35610 ( .A1(n2812), .A2(n2837), .ZN(n4305) );
  INV_X1 U35620 ( .A(n3489), .ZN(n2813) );
  AOI22_X1 U35630 ( .A1(n2813), .A2(REG1_REG_24__SCAN_IN), .B1(n2996), .B2(
        REG2_REG_24__SCAN_IN), .ZN(n2815) );
  NAND2_X1 U35640 ( .A1(n3487), .A2(REG0_REG_24__SCAN_IN), .ZN(n2814) );
  NAND2_X1 U35650 ( .A1(n4321), .A2(n3040), .ZN(n2817) );
  OR2_X1 U35660 ( .A1(n4308), .A2(n2832), .ZN(n2816) );
  NAND2_X1 U35670 ( .A1(n2817), .A2(n2816), .ZN(n2822) );
  INV_X1 U35680 ( .A(n2822), .ZN(n2818) );
  INV_X1 U35690 ( .A(n4321), .ZN(n4283) );
  OAI22_X1 U35700 ( .A1(n4283), .A2(n2832), .B1(n4308), .B2(n2843), .ZN(n2821)
         );
  XOR2_X1 U35710 ( .A(n3038), .B(n2821), .Z(n3915) );
  INV_X1 U35720 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3891) );
  XNOR2_X1 U35730 ( .A(n2837), .B(n3891), .ZN(n4291) );
  NAND2_X1 U35740 ( .A1(n4291), .A2(n2949), .ZN(n2828) );
  INV_X1 U35750 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4563) );
  NAND2_X1 U35760 ( .A1(n2996), .A2(REG2_REG_25__SCAN_IN), .ZN(n2825) );
  NAND2_X1 U35770 ( .A1(n3487), .A2(REG0_REG_25__SCAN_IN), .ZN(n2824) );
  OAI211_X1 U35780 ( .C1(n3489), .C2(n4563), .A(n2825), .B(n2824), .ZN(n2826)
         );
  INV_X1 U35790 ( .A(n2826), .ZN(n2827) );
  NAND2_X1 U35800 ( .A1(n4302), .A2(n4119), .ZN(n2830) );
  OR2_X1 U35810 ( .A1(n4289), .A2(n2843), .ZN(n2829) );
  NAND2_X1 U3582 ( .A1(n2830), .A2(n2829), .ZN(n2831) );
  XNOR2_X1 U3583 ( .A(n2831), .B(n2846), .ZN(n2835) );
  NOR2_X1 U3584 ( .A1(n4289), .A2(n2832), .ZN(n2833) );
  AOI21_X1 U3585 ( .B1(n4302), .B2(n3040), .A(n2833), .ZN(n2834) );
  NAND2_X1 U3586 ( .A1(n2835), .A2(n2834), .ZN(n3888) );
  NOR2_X1 U3587 ( .A1(n2835), .A2(n2834), .ZN(n3889) );
  AND2_X1 U3588 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2836) );
  AOI21_X1 U3589 ( .B1(n2837), .B2(REG3_REG_25__SCAN_IN), .A(
        REG3_REG_26__SCAN_IN), .ZN(n2838) );
  INV_X1 U3590 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4559) );
  NAND2_X1 U3591 ( .A1(n2996), .A2(REG2_REG_26__SCAN_IN), .ZN(n2840) );
  NAND2_X1 U3592 ( .A1(n3487), .A2(REG0_REG_26__SCAN_IN), .ZN(n2839) );
  OAI211_X1 U3593 ( .C1(n3489), .C2(n4559), .A(n2840), .B(n2839), .ZN(n2841)
         );
  INV_X1 U3594 ( .A(n2841), .ZN(n2842) );
  OAI21_X2 U3595 ( .B1(n2885), .B2(n3001), .A(n2842), .ZN(n4285) );
  NAND2_X1 U3596 ( .A1(n4285), .A2(n4119), .ZN(n2845) );
  OR2_X1 U3597 ( .A1(n4264), .A2(n2843), .ZN(n2844) );
  NAND2_X1 U3598 ( .A1(n2845), .A2(n2844), .ZN(n2847) );
  XNOR2_X1 U3599 ( .A(n2847), .B(n2846), .ZN(n2850) );
  NOR2_X1 U3600 ( .A1(n4264), .A2(n2832), .ZN(n2848) );
  AOI21_X1 U3601 ( .B1(n4285), .B2(n2508), .A(n2848), .ZN(n2849) );
  AND2_X1 U3602 ( .A1(n2850), .A2(n2849), .ZN(n3019) );
  OR2_X1 U3603 ( .A1(n2850), .A2(n2849), .ZN(n3020) );
  NAND2_X1 U3604 ( .A1(n2360), .A2(n3020), .ZN(n2851) );
  XNOR2_X1 U3605 ( .A(n3021), .B(n2851), .ZN(n2898) );
  NAND2_X1 U3606 ( .A1(n2856), .A2(n2852), .ZN(n2853) );
  MUX2_X1 U3607 ( .A(n2852), .B(n2853), .S(B_REG_SCAN_IN), .Z(n2855) );
  INV_X1 U3608 ( .A(n2856), .ZN(n4674) );
  OAI22_X1 U3609 ( .A1(n3073), .A2(D_REG_1__SCAN_IN), .B1(n2854), .B2(n4674), 
        .ZN(n3145) );
  NOR4_X1 U3610 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_26__SCAN_IN), .ZN(n2865) );
  NOR4_X1 U3611 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_23__SCAN_IN), .ZN(n2864) );
  INV_X1 U3612 ( .A(D_REG_7__SCAN_IN), .ZN(n4899) );
  INV_X1 U3613 ( .A(D_REG_20__SCAN_IN), .ZN(n4896) );
  INV_X1 U3614 ( .A(D_REG_25__SCAN_IN), .ZN(n4891) );
  INV_X1 U3615 ( .A(D_REG_21__SCAN_IN), .ZN(n4895) );
  NAND4_X1 U3616 ( .A1(n4899), .A2(n4896), .A3(n4891), .A4(n4895), .ZN(n2862)
         );
  NOR4_X1 U3617 ( .A1(D_REG_8__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_11__SCAN_IN), .ZN(n2860) );
  NOR4_X1 U3618 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2859) );
  NOR4_X1 U3619 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2858) );
  NOR4_X1 U3620 ( .A1(D_REG_12__SCAN_IN), .A2(D_REG_13__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2857) );
  NAND4_X1 U3621 ( .A1(n2860), .A2(n2859), .A3(n2858), .A4(n2857), .ZN(n2861)
         );
  NOR4_X1 U3622 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(n2862), 
        .A4(n2861), .ZN(n2863) );
  AND3_X1 U3623 ( .A1(n2865), .A2(n2864), .A3(n2863), .ZN(n2866) );
  NOR2_X1 U3624 ( .A1(n3145), .A2(n3006), .ZN(n2867) );
  INV_X1 U3625 ( .A(n2852), .ZN(n3077) );
  INV_X1 U3626 ( .A(n3146), .ZN(n3009) );
  NAND2_X1 U3627 ( .A1(n2867), .A2(n3009), .ZN(n2887) );
  INV_X1 U3628 ( .A(n2887), .ZN(n2871) );
  NAND2_X1 U3629 ( .A1(n4111), .A2(n4695), .ZN(n2888) );
  AOI21_X1 U3630 ( .B1(n2872), .B2(n2888), .A(n3080), .ZN(n2873) );
  NAND2_X1 U3631 ( .A1(n2891), .A2(n2260), .ZN(n2877) );
  NAND2_X1 U3632 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2875) );
  NAND2_X1 U3633 ( .A1(n2874), .A2(n2875), .ZN(n2876) );
  NOR2_X2 U3634 ( .A1(n2877), .A2(n4673), .ZN(n4711) );
  OR2_X1 U3635 ( .A1(n2878), .A2(REG3_REG_27__SCAN_IN), .ZN(n2879) );
  NAND2_X1 U3636 ( .A1(n2878), .A2(REG3_REG_27__SCAN_IN), .ZN(n2947) );
  NAND2_X1 U3637 ( .A1(n4252), .A2(n2496), .ZN(n2884) );
  INV_X1 U3638 ( .A(REG1_REG_27__SCAN_IN), .ZN(n3587) );
  NAND2_X1 U3639 ( .A1(n2950), .A2(REG2_REG_27__SCAN_IN), .ZN(n2881) );
  NAND2_X1 U3640 ( .A1(n3487), .A2(REG0_REG_27__SCAN_IN), .ZN(n2880) );
  OAI211_X1 U3641 ( .C1(n3489), .C2(n3587), .A(n2881), .B(n2880), .ZN(n2882)
         );
  INV_X1 U3642 ( .A(n2882), .ZN(n2883) );
  AOI22_X1 U3643 ( .A1(n4724), .A2(n4302), .B1(n4711), .B2(n4266), .ZN(n2896)
         );
  INV_X1 U3644 ( .A(n2885), .ZN(n4273) );
  NOR2_X1 U3645 ( .A1(n4874), .A2(n4695), .ZN(n2886) );
  NAND2_X1 U3646 ( .A1(n4858), .A2(n2886), .ZN(n3007) );
  NAND2_X1 U3647 ( .A1(n2887), .A2(n3007), .ZN(n3135) );
  AND2_X1 U3648 ( .A1(n3080), .A2(n2888), .ZN(n3005) );
  INV_X1 U3649 ( .A(n3005), .ZN(n2889) );
  NAND4_X1 U3650 ( .A1(n3135), .A2(n3082), .A3(n3059), .A4(n2889), .ZN(n2890)
         );
  NAND2_X1 U3651 ( .A1(n2890), .A2(STATE_REG_SCAN_IN), .ZN(n4728) );
  NAND2_X1 U3652 ( .A1(n2891), .A2(n4543), .ZN(n2892) );
  INV_X1 U3653 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2893) );
  OAI22_X1 U3654 ( .A1(n3953), .A2(n4264), .B1(STATE_REG_SCAN_IN), .B2(n2893), 
        .ZN(n2894) );
  AOI21_X1 U3655 ( .B1(n4273), .B2(n3955), .A(n2894), .ZN(n2895) );
  OAI21_X1 U3656 ( .B1(n2898), .B2(n4719), .A(n2897), .ZN(U3237) );
  INV_X1 U3657 ( .A(REG1_REG_28__SCAN_IN), .ZN(n3835) );
  NAND2_X1 U3658 ( .A1(n4879), .A2(n3141), .ZN(n2959) );
  NAND2_X1 U3659 ( .A1(n2899), .A2(n3156), .ZN(n4044) );
  AND2_X1 U3660 ( .A1(n2900), .A2(n3136), .ZN(n3151) );
  CLKBUF_X1 U3661 ( .A(n2899), .Z(n4133) );
  NAND2_X1 U3662 ( .A1(n4133), .A2(n3141), .ZN(n2901) );
  NAND2_X1 U3663 ( .A1(n3153), .A2(n2901), .ZN(n3234) );
  INV_X1 U3664 ( .A(n3234), .ZN(n2902) );
  NAND2_X1 U3665 ( .A1(n3199), .A2(n3246), .ZN(n4051) );
  NAND2_X1 U3666 ( .A1(n2902), .A2(n3237), .ZN(n3233) );
  NAND2_X1 U3667 ( .A1(n3179), .A2(n3246), .ZN(n2903) );
  NAND2_X1 U3668 ( .A1(n3233), .A2(n2903), .ZN(n3176) );
  NOR2_X1 U3669 ( .A1(n4132), .A2(n3202), .ZN(n2904) );
  INV_X1 U3670 ( .A(n4132), .ZN(n3297) );
  INV_X1 U3671 ( .A(n3202), .ZN(n2961) );
  INV_X1 U3672 ( .A(n3200), .ZN(n3276) );
  NAND2_X1 U3673 ( .A1(n3276), .A2(n3295), .ZN(n4054) );
  NAND2_X1 U3674 ( .A1(n3200), .A2(n3291), .ZN(n4057) );
  NAND2_X1 U3675 ( .A1(n3293), .A2(n4023), .ZN(n2906) );
  NAND2_X1 U3676 ( .A1(n3200), .A2(n3295), .ZN(n2905) );
  NAND2_X1 U3677 ( .A1(n2906), .A2(n2905), .ZN(n3262) );
  AND2_X1 U3678 ( .A1(n4131), .A2(n3273), .ZN(n3321) );
  OR2_X1 U3679 ( .A1(n3503), .A2(n3326), .ZN(n2907) );
  INV_X1 U3680 ( .A(n4131), .ZN(n3328) );
  INV_X1 U3681 ( .A(n3273), .ZN(n3256) );
  NAND2_X1 U3682 ( .A1(n3328), .A2(n3256), .ZN(n3322) );
  AND2_X1 U3683 ( .A1(n2907), .A2(n3322), .ZN(n2908) );
  OAI21_X1 U3684 ( .B1(n3262), .B2(n3321), .A(n2908), .ZN(n2910) );
  NAND2_X1 U3685 ( .A1(n3503), .A2(n3326), .ZN(n2909) );
  NAND2_X1 U3686 ( .A1(n2910), .A2(n2909), .ZN(n3311) );
  INV_X1 U3687 ( .A(n4130), .ZN(n3285) );
  NAND2_X1 U3688 ( .A1(n3285), .A2(n3312), .ZN(n2965) );
  INV_X1 U3689 ( .A(n3312), .ZN(n3504) );
  NAND2_X1 U3690 ( .A1(n4130), .A2(n3504), .ZN(n4067) );
  NAND2_X1 U3691 ( .A1(n2965), .A2(n4067), .ZN(n4030) );
  NAND2_X1 U3692 ( .A1(n3311), .A2(n4030), .ZN(n2912) );
  NAND2_X1 U3693 ( .A1(n4130), .A2(n3312), .ZN(n2911) );
  AND2_X1 U3694 ( .A1(n3502), .A2(n2967), .ZN(n2913) );
  NOR2_X1 U3695 ( .A1(n3432), .A2(n3373), .ZN(n2914) );
  INV_X1 U3696 ( .A(n3432), .ZN(n3357) );
  INV_X1 U3697 ( .A(n3373), .ZN(n3423) );
  INV_X1 U3698 ( .A(n4862), .ZN(n2969) );
  INV_X1 U3699 ( .A(n4129), .ZN(n3463) );
  NAND2_X1 U3700 ( .A1(n3463), .A2(n4870), .ZN(n3470) );
  NAND2_X1 U3701 ( .A1(n4129), .A2(n4859), .ZN(n2970) );
  NOR2_X1 U3702 ( .A1(n4128), .A2(n2971), .ZN(n2917) );
  INV_X1 U3703 ( .A(n4128), .ZN(n4860) );
  OAI22_X2 U3704 ( .A1(n3474), .A2(n2917), .B1(n4860), .B2(n3476), .ZN(n4508)
         );
  NAND2_X1 U3705 ( .A1(n2919), .A2(n4498), .ZN(n3976) );
  NAND2_X1 U3706 ( .A1(n4517), .A2(n3513), .ZN(n3972) );
  NOR2_X1 U3707 ( .A1(n4465), .A2(n4477), .ZN(n2920) );
  INV_X1 U3708 ( .A(n4127), .ZN(n4497) );
  NOR2_X1 U3709 ( .A1(n4497), .A2(n4525), .ZN(n4469) );
  NOR3_X1 U3710 ( .A1(n4491), .A2(n2920), .A3(n4469), .ZN(n2922) );
  NAND2_X1 U3711 ( .A1(n2919), .A2(n3513), .ZN(n4471) );
  OAI22_X1 U3712 ( .A1(n2920), .A2(n4471), .B1(n4474), .B2(n4494), .ZN(n2921)
         );
  NAND2_X1 U3713 ( .A1(n4478), .A2(n4462), .ZN(n3974) );
  NAND2_X1 U3714 ( .A1(n4439), .A2(n4453), .ZN(n4088) );
  NAND2_X1 U3715 ( .A1(n3974), .A2(n4088), .ZN(n4451) );
  NAND2_X1 U3716 ( .A1(n4452), .A2(n4451), .ZN(n4450) );
  INV_X1 U3717 ( .A(n4723), .ZN(n4418) );
  INV_X1 U3718 ( .A(n4442), .ZN(n4436) );
  NAND2_X1 U3719 ( .A1(n4418), .A2(n4436), .ZN(n2924) );
  NAND2_X1 U3720 ( .A1(n4437), .A2(n4713), .ZN(n4395) );
  NAND2_X1 U3721 ( .A1(n4402), .A2(n2925), .ZN(n4396) );
  NAND2_X1 U3722 ( .A1(n4395), .A2(n4396), .ZN(n4422) );
  NAND2_X1 U3723 ( .A1(n4423), .A2(n4422), .ZN(n4421) );
  INV_X1 U3724 ( .A(n4407), .ZN(n2978) );
  NAND2_X1 U3725 ( .A1(n4710), .A2(n2978), .ZN(n2927) );
  INV_X1 U3726 ( .A(n4385), .ZN(n4377) );
  NAND2_X1 U3727 ( .A1(n4371), .A2(n2928), .ZN(n2929) );
  INV_X1 U3728 ( .A(n4126), .ZN(n4400) );
  NAND2_X1 U3729 ( .A1(n2929), .A2(n2377), .ZN(n4353) );
  INV_X1 U3730 ( .A(n4353), .ZN(n2931) );
  INV_X1 U3731 ( .A(n4378), .ZN(n2983) );
  NAND2_X1 U3732 ( .A1(n2932), .A2(n4336), .ZN(n4317) );
  NAND2_X1 U3733 ( .A1(n4358), .A2(n4345), .ZN(n2984) );
  NAND2_X1 U3734 ( .A1(n4317), .A2(n2984), .ZN(n4333) );
  NAND2_X1 U3735 ( .A1(n4348), .A2(n2934), .ZN(n2936) );
  INV_X1 U3736 ( .A(n4308), .ZN(n2937) );
  NAND2_X1 U3737 ( .A1(n4321), .A2(n2937), .ZN(n2938) );
  INV_X1 U3738 ( .A(n4302), .ZN(n4269) );
  NAND2_X1 U3739 ( .A1(n4269), .A2(n4289), .ZN(n2940) );
  NOR2_X1 U3740 ( .A1(n4269), .A2(n4289), .ZN(n2939) );
  NAND2_X1 U3741 ( .A1(n4285), .A2(n4270), .ZN(n2942) );
  NOR2_X1 U3742 ( .A1(n4285), .A2(n4270), .ZN(n2941) );
  INV_X1 U3743 ( .A(n4249), .ZN(n3027) );
  NAND2_X1 U3744 ( .A1(n4042), .A2(n3027), .ZN(n2945) );
  NOR2_X1 U3745 ( .A1(n4042), .A2(n3027), .ZN(n2944) );
  AOI21_X1 U3746 ( .B1(n4238), .B2(n2945), .A(n2944), .ZN(n4221) );
  INV_X1 U3747 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2946) );
  NAND2_X1 U3748 ( .A1(n2947), .A2(n2946), .ZN(n2948) );
  NAND2_X1 U3749 ( .A1(n4230), .A2(n2949), .ZN(n2955) );
  NAND2_X1 U3750 ( .A1(n2950), .A2(REG2_REG_28__SCAN_IN), .ZN(n2952) );
  NAND2_X1 U3751 ( .A1(n3487), .A2(REG0_REG_28__SCAN_IN), .ZN(n2951) );
  OAI211_X1 U3752 ( .C1(n3489), .C2(n3835), .A(n2952), .B(n2951), .ZN(n2953)
         );
  INV_X1 U3753 ( .A(n2953), .ZN(n2954) );
  NAND2_X1 U3754 ( .A1(n4243), .A2(n4217), .ZN(n4206) );
  NAND2_X1 U3755 ( .A1(n4207), .A2(n4206), .ZN(n4003) );
  XNOR2_X1 U3756 ( .A(n4221), .B(n4003), .ZN(n4229) );
  XNOR2_X1 U3757 ( .A(n3162), .B(n4675), .ZN(n2956) );
  NAND2_X1 U3758 ( .A1(n4111), .A2(n4685), .ZN(n4881) );
  INV_X1 U3759 ( .A(n2234), .ZN(n2958) );
  NAND2_X1 U3760 ( .A1(n2958), .A2(n3136), .ZN(n4043) );
  NAND2_X1 U3761 ( .A1(n3238), .A2(n4020), .ZN(n2960) );
  NAND2_X1 U3762 ( .A1(n2960), .A2(n4048), .ZN(n3177) );
  NAND2_X1 U3763 ( .A1(n3297), .A2(n3202), .ZN(n4053) );
  NAND2_X1 U3764 ( .A1(n4132), .A2(n2961), .ZN(n4050) );
  NAND2_X1 U3765 ( .A1(n3177), .A2(n4022), .ZN(n2962) );
  INV_X1 U3766 ( .A(n4054), .ZN(n2963) );
  AND2_X1 U3767 ( .A1(n4131), .A2(n3256), .ZN(n3263) );
  NAND2_X1 U3768 ( .A1(n3328), .A2(n3273), .ZN(n4071) );
  NAND2_X1 U3769 ( .A1(n3503), .A2(n2271), .ZN(n4068) );
  NAND2_X1 U3770 ( .A1(n3325), .A2(n4068), .ZN(n2964) );
  INV_X1 U3771 ( .A(n3503), .ZN(n3257) );
  NAND2_X1 U3772 ( .A1(n3257), .A2(n3326), .ZN(n4059) );
  INV_X1 U3773 ( .A(n2965), .ZN(n2966) );
  INV_X1 U3774 ( .A(n3502), .ZN(n3375) );
  NAND2_X1 U3775 ( .A1(n3375), .A2(n2967), .ZN(n4064) );
  NAND2_X1 U3776 ( .A1(n3502), .A2(n3363), .ZN(n4069) );
  NAND2_X1 U3777 ( .A1(n2968), .A2(n4069), .ZN(n3372) );
  AND2_X1 U3778 ( .A1(n3432), .A2(n3423), .ZN(n4077) );
  NAND2_X1 U3779 ( .A1(n3357), .A2(n3373), .ZN(n4063) );
  NAND2_X1 U3780 ( .A1(n4862), .A2(n3437), .ZN(n4079) );
  NAND2_X1 U3781 ( .A1(n2969), .A2(n3010), .ZN(n4076) );
  NAND2_X1 U3782 ( .A1(n4128), .A2(n3476), .ZN(n4510) );
  NAND2_X1 U3783 ( .A1(n4127), .A2(n4525), .ZN(n4005) );
  NAND2_X1 U3784 ( .A1(n4510), .A2(n4005), .ZN(n2972) );
  INV_X1 U3785 ( .A(n2970), .ZN(n3469) );
  NOR2_X1 U3786 ( .A1(n2972), .A2(n3469), .ZN(n4080) );
  NAND2_X1 U3787 ( .A1(n3468), .A2(n4080), .ZN(n2975) );
  NAND2_X1 U3788 ( .A1(n4860), .A2(n2971), .ZN(n4509) );
  NAND2_X1 U3789 ( .A1(n3470), .A2(n4509), .ZN(n2974) );
  INV_X1 U3790 ( .A(n2972), .ZN(n2973) );
  NOR2_X1 U3791 ( .A1(n4127), .A2(n4525), .ZN(n4006) );
  AOI21_X1 U3792 ( .B1(n2974), .B2(n2973), .A(n4006), .ZN(n4086) );
  NAND2_X1 U3793 ( .A1(n2975), .A2(n4086), .ZN(n4492) );
  NAND2_X1 U3794 ( .A1(n4465), .A2(n4474), .ZN(n3975) );
  NAND2_X1 U3795 ( .A1(n4494), .A2(n4477), .ZN(n3973) );
  NAND2_X1 U3796 ( .A1(n3975), .A2(n3973), .ZN(n4481) );
  NAND2_X1 U3797 ( .A1(n4479), .A2(n3973), .ZN(n4461) );
  INV_X1 U3798 ( .A(n4451), .ZN(n4460) );
  NAND2_X1 U3799 ( .A1(n4461), .A2(n4460), .ZN(n4459) );
  NAND2_X1 U3800 ( .A1(n4710), .A2(n4407), .ZN(n2976) );
  AND2_X1 U3801 ( .A1(n4396), .A2(n2976), .ZN(n3978) );
  NAND2_X1 U3802 ( .A1(n4436), .A2(n4723), .ZN(n4027) );
  NAND2_X1 U3803 ( .A1(n3978), .A2(n4027), .ZN(n4091) );
  NAND2_X1 U3804 ( .A1(n4418), .A2(n4442), .ZN(n4393) );
  NAND2_X1 U3805 ( .A1(n4395), .A2(n4393), .ZN(n2977) );
  NAND2_X1 U3806 ( .A1(n2977), .A2(n3978), .ZN(n2980) );
  NAND2_X1 U3807 ( .A1(n4380), .A2(n2978), .ZN(n2979) );
  NAND2_X1 U3808 ( .A1(n2980), .A2(n2979), .ZN(n4372) );
  NOR2_X1 U3809 ( .A1(n4126), .A2(n4385), .ZN(n2981) );
  OR2_X1 U3810 ( .A1(n4372), .A2(n2981), .ZN(n3981) );
  INV_X1 U3811 ( .A(n3981), .ZN(n4090) );
  NAND2_X1 U3812 ( .A1(n4126), .A2(n4385), .ZN(n4093) );
  NAND2_X1 U3813 ( .A1(n2983), .A2(n4357), .ZN(n4315) );
  AND2_X1 U3814 ( .A1(n4317), .A2(n4315), .ZN(n4097) );
  NAND2_X1 U3815 ( .A1(n4355), .A2(n4097), .ZN(n2987) );
  NAND2_X1 U3816 ( .A1(n4125), .A2(n2934), .ZN(n4013) );
  AND2_X1 U3817 ( .A1(n4013), .A2(n2984), .ZN(n4101) );
  AND2_X1 U3818 ( .A1(n4378), .A2(n4362), .ZN(n4314) );
  NAND2_X1 U3819 ( .A1(n4317), .A2(n4314), .ZN(n2985) );
  NAND2_X1 U3820 ( .A1(n4101), .A2(n2985), .ZN(n3983) );
  INV_X1 U3821 ( .A(n3983), .ZN(n2986) );
  NAND2_X1 U3822 ( .A1(n2987), .A2(n2986), .ZN(n4298) );
  OR2_X1 U3823 ( .A1(n4321), .A2(n4308), .ZN(n4004) );
  NAND2_X1 U3824 ( .A1(n4348), .A2(n4320), .ZN(n4297) );
  NAND2_X1 U3825 ( .A1(n4004), .A2(n4297), .ZN(n4099) );
  INV_X1 U3826 ( .A(n4099), .ZN(n2988) );
  NAND2_X1 U3827 ( .A1(n4298), .A2(n2988), .ZN(n4280) );
  OR2_X1 U3828 ( .A1(n4285), .A2(n4264), .ZN(n2989) );
  OR2_X1 U3829 ( .A1(n4302), .A2(n4289), .ZN(n4258) );
  AND2_X1 U3830 ( .A1(n2989), .A2(n4258), .ZN(n3986) );
  INV_X1 U3831 ( .A(n3986), .ZN(n4098) );
  NAND2_X1 U3832 ( .A1(n4302), .A2(n4289), .ZN(n4036) );
  NAND2_X1 U3833 ( .A1(n4321), .A2(n4308), .ZN(n4279) );
  AND2_X1 U3834 ( .A1(n4036), .A2(n4279), .ZN(n4260) );
  INV_X1 U3835 ( .A(n4260), .ZN(n2990) );
  NAND2_X1 U3836 ( .A1(n2990), .A2(n3986), .ZN(n2991) );
  NAND2_X1 U3837 ( .A1(n4285), .A2(n4264), .ZN(n3992) );
  NAND2_X1 U3838 ( .A1(n2991), .A2(n3992), .ZN(n4103) );
  INV_X1 U3839 ( .A(n4103), .ZN(n2992) );
  XNOR2_X1 U3840 ( .A(n4266), .B(n4249), .ZN(n4237) );
  INV_X1 U3841 ( .A(n4237), .ZN(n4239) );
  NAND2_X1 U3842 ( .A1(n4042), .A2(n4249), .ZN(n3985) );
  INV_X1 U3843 ( .A(n3985), .ZN(n3993) );
  XNOR2_X1 U3844 ( .A(n2237), .B(n4003), .ZN(n2995) );
  NAND2_X1 U3845 ( .A1(n4675), .A2(n4685), .ZN(n2994) );
  INV_X1 U3846 ( .A(n4111), .ZN(n4676) );
  NAND2_X1 U3847 ( .A1(n4676), .A2(n4046), .ZN(n4001) );
  NAND2_X1 U3848 ( .A1(n2995), .A2(n4876), .ZN(n3004) );
  INV_X1 U3849 ( .A(REG1_REG_29__SCAN_IN), .ZN(n3810) );
  NAND2_X1 U3850 ( .A1(n3487), .A2(REG0_REG_29__SCAN_IN), .ZN(n2998) );
  NAND2_X1 U3851 ( .A1(n2996), .A2(REG2_REG_29__SCAN_IN), .ZN(n2997) );
  OAI211_X1 U3852 ( .C1(n3489), .C2(n3810), .A(n2998), .B(n2997), .ZN(n2999)
         );
  INV_X1 U3853 ( .A(n2999), .ZN(n3000) );
  OAI21_X1 U3854 ( .B1(n4205), .B2(n3001), .A(n3000), .ZN(n3991) );
  NOR2_X1 U3855 ( .A1(n4217), .A2(n4858), .ZN(n3002) );
  AOI21_X1 U3856 ( .B1(n3991), .B2(n4516), .A(n3002), .ZN(n3003) );
  OAI211_X1 U3857 ( .C1(n4042), .C2(n4519), .A(n3004), .B(n3003), .ZN(n4234)
         );
  AOI21_X1 U3858 ( .B1(n4229), .B2(n4968), .A(n4234), .ZN(n3015) );
  AND2_X1 U3859 ( .A1(n3145), .A2(n3007), .ZN(n3008) );
  NAND2_X1 U3860 ( .A1(n3247), .A2(n3246), .ZN(n3183) );
  NAND2_X1 U3861 ( .A1(n3292), .A2(n3291), .ZN(n3266) );
  NAND2_X1 U3862 ( .A1(n4869), .A2(n3476), .ZN(n3475) );
  INV_X1 U3863 ( .A(n4289), .ZN(n3011) );
  OAI21_X1 U3864 ( .B1(n4248), .B2(n4217), .A(n4224), .ZN(n4232) );
  NAND2_X1 U3865 ( .A1(n3013), .A2(n3012), .ZN(U3546) );
  INV_X1 U3866 ( .A(REG0_REG_28__SCAN_IN), .ZN(n3016) );
  NAND2_X1 U3867 ( .A1(n3018), .A2(n3017), .ZN(U3514) );
  NAND2_X1 U3868 ( .A1(n4266), .A2(n4119), .ZN(n3023) );
  NAND2_X1 U3869 ( .A1(n4249), .A2(n3035), .ZN(n3022) );
  NAND2_X1 U3870 ( .A1(n3023), .A2(n3022), .ZN(n3024) );
  XNOR2_X1 U3871 ( .A(n3024), .B(n3038), .ZN(n3046) );
  AND2_X1 U3872 ( .A1(n4249), .A2(n2714), .ZN(n3025) );
  AOI21_X1 U3873 ( .B1(n4266), .B2(n3040), .A(n3025), .ZN(n3044) );
  XNOR2_X1 U3874 ( .A(n3046), .B(n3044), .ZN(n3033) );
  XNOR2_X1 U3875 ( .A(n3034), .B(n3033), .ZN(n3032) );
  AOI22_X1 U3876 ( .A1(n4724), .A2(n4285), .B1(n3963), .B2(n4243), .ZN(n3030)
         );
  INV_X1 U3877 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3026) );
  OAI22_X1 U3878 ( .A1(n3953), .A2(n3027), .B1(STATE_REG_SCAN_IN), .B2(n3026), 
        .ZN(n3028) );
  AOI21_X1 U3879 ( .B1(n4252), .B2(n3955), .A(n3028), .ZN(n3029) );
  AND2_X1 U3880 ( .A1(n3030), .A2(n3029), .ZN(n3031) );
  OAI21_X1 U3881 ( .B1(n3032), .B2(n4719), .A(n3031), .ZN(U3211) );
  NAND2_X1 U3882 ( .A1(n3034), .A2(n3033), .ZN(n3058) );
  NAND2_X1 U3883 ( .A1(n4243), .A2(n4119), .ZN(n3037) );
  INV_X1 U3884 ( .A(n4217), .ZN(n3049) );
  NAND2_X1 U3885 ( .A1(n3049), .A2(n3035), .ZN(n3036) );
  NAND2_X1 U3886 ( .A1(n3037), .A2(n3036), .ZN(n3039) );
  XNOR2_X1 U3887 ( .A(n3039), .B(n3038), .ZN(n3042) );
  AOI22_X1 U3888 ( .A1(n4243), .A2(n3040), .B1(n3049), .B2(n4119), .ZN(n3041)
         );
  XNOR2_X1 U3889 ( .A(n3042), .B(n3041), .ZN(n3048) );
  INV_X1 U3890 ( .A(n3048), .ZN(n3043) );
  NAND2_X1 U3891 ( .A1(n3043), .A2(n3968), .ZN(n3057) );
  INV_X1 U3892 ( .A(n3044), .ZN(n3045) );
  NAND2_X1 U3893 ( .A1(n3046), .A2(n3045), .ZN(n3047) );
  NAND2_X1 U3894 ( .A1(n3058), .A2(n2255), .ZN(n3056) );
  NOR3_X1 U3895 ( .A1(n3048), .A2(n4719), .A3(n3047), .ZN(n3054) );
  INV_X1 U3896 ( .A(n4230), .ZN(n3052) );
  AOI22_X1 U3897 ( .A1(n4724), .A2(n4266), .B1(n3963), .B2(n3991), .ZN(n3051)
         );
  AOI22_X1 U3898 ( .A1(n4712), .A2(n3049), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3050) );
  OAI211_X1 U3899 ( .C1(n4728), .C2(n3052), .A(n3051), .B(n3050), .ZN(n3053)
         );
  NOR2_X1 U3900 ( .A1(n3054), .A2(n3053), .ZN(n3055) );
  OAI211_X1 U3901 ( .C1(n3058), .C2(n3057), .A(n3056), .B(n3055), .ZN(U3217)
         );
  INV_X1 U3902 ( .A(DATAI_21_), .ZN(n3837) );
  NAND2_X1 U3903 ( .A1(n4046), .A2(STATE_REG_SCAN_IN), .ZN(n3060) );
  OAI21_X1 U3904 ( .B1(STATE_REG_SCAN_IN), .B2(n3837), .A(n3060), .ZN(U3331)
         );
  MUX2_X1 U3905 ( .A(n3061), .B(n4695), .S(STATE_REG_SCAN_IN), .Z(n3062) );
  INV_X1 U3906 ( .A(n3062), .ZN(U3333) );
  INV_X1 U3907 ( .A(DATAI_24_), .ZN(n3063) );
  MUX2_X1 U3908 ( .A(n3063), .B(n2852), .S(STATE_REG_SCAN_IN), .Z(n3064) );
  INV_X1 U3909 ( .A(n3064), .ZN(U3328) );
  INV_X1 U3910 ( .A(DATAI_29_), .ZN(n3067) );
  NAND2_X1 U3911 ( .A1(n3065), .A2(STATE_REG_SCAN_IN), .ZN(n3066) );
  OAI21_X1 U3912 ( .B1(STATE_REG_SCAN_IN), .B2(n3067), .A(n3066), .ZN(U3323)
         );
  INV_X1 U3913 ( .A(DATAI_27_), .ZN(n3069) );
  XNOR2_X1 U3914 ( .A(n2874), .B(IR_REG_27__SCAN_IN), .ZN(n4737) );
  NAND2_X1 U3915 ( .A1(n4737), .A2(STATE_REG_SCAN_IN), .ZN(n3068) );
  OAI21_X1 U3916 ( .B1(STATE_REG_SCAN_IN), .B2(n3069), .A(n3068), .ZN(U3325)
         );
  INV_X1 U3917 ( .A(DATAI_30_), .ZN(n3770) );
  INV_X1 U3918 ( .A(n3070), .ZN(n3071) );
  NAND2_X1 U3919 ( .A1(n3071), .A2(STATE_REG_SCAN_IN), .ZN(n3072) );
  OAI21_X1 U3920 ( .B1(STATE_REG_SCAN_IN), .B2(n3770), .A(n3072), .ZN(U3322)
         );
  INV_X1 U3921 ( .A(D_REG_1__SCAN_IN), .ZN(n3076) );
  NOR3_X1 U3922 ( .A1(n4674), .A2(n2854), .A3(n4904), .ZN(n3075) );
  AOI21_X1 U3923 ( .B1(n4903), .B2(n3076), .A(n3075), .ZN(U3459) );
  INV_X1 U3924 ( .A(D_REG_0__SCAN_IN), .ZN(n3079) );
  NOR3_X1 U3925 ( .A1(n2854), .A2(n3077), .A3(n4904), .ZN(n3078) );
  AOI21_X1 U3926 ( .B1(n4903), .B2(n3079), .A(n3078), .ZN(U3458) );
  NAND2_X1 U3927 ( .A1(n3080), .A2(n3082), .ZN(n3081) );
  INV_X1 U3928 ( .A(n3096), .ZN(n3084) );
  OR2_X1 U3929 ( .A1(n3082), .A2(U3149), .ZN(n4122) );
  NAND2_X1 U3930 ( .A1(n3083), .A2(n4122), .ZN(n3097) );
  NOR2_X1 U3931 ( .A1(n4825), .A2(U4043), .ZN(U3148) );
  INV_X1 U3932 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n3841) );
  NAND2_X1 U3933 ( .A1(n3200), .A2(U4043), .ZN(n3085) );
  OAI21_X1 U3934 ( .B1(n3841), .B2(U4043), .A(n3085), .ZN(U3554) );
  INV_X1 U3935 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n3790) );
  NAND2_X1 U3936 ( .A1(n3503), .A2(U4043), .ZN(n3086) );
  OAI21_X1 U3937 ( .B1(U4043), .B2(n3790), .A(n3086), .ZN(U3556) );
  INV_X1 U3938 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n3816) );
  NAND2_X1 U3939 ( .A1(n3502), .A2(U4043), .ZN(n3087) );
  OAI21_X1 U3940 ( .B1(U4043), .B2(n3816), .A(n3087), .ZN(U3558) );
  INV_X1 U3941 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n3606) );
  INV_X1 U3942 ( .A(REG1_REG_30__SCAN_IN), .ZN(n3090) );
  NAND2_X1 U3943 ( .A1(n2996), .A2(REG2_REG_30__SCAN_IN), .ZN(n3089) );
  NAND2_X1 U3944 ( .A1(n3487), .A2(REG0_REG_30__SCAN_IN), .ZN(n3088) );
  OAI211_X1 U3945 ( .C1(n3489), .C2(n3090), .A(n3089), .B(n3088), .ZN(n4212)
         );
  NAND2_X1 U3946 ( .A1(n4212), .A2(U4043), .ZN(n3091) );
  OAI21_X1 U3947 ( .B1(U4043), .B2(n3606), .A(n3091), .ZN(U3580) );
  INV_X1 U3948 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n3603) );
  NAND2_X1 U3949 ( .A1(n3199), .A2(U4043), .ZN(n3092) );
  OAI21_X1 U3950 ( .B1(U4043), .B2(n3603), .A(n3092), .ZN(U3552) );
  INV_X1 U3951 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n3793) );
  NAND2_X1 U3952 ( .A1(n3432), .A2(U4043), .ZN(n3093) );
  OAI21_X1 U3953 ( .B1(U4043), .B2(n3793), .A(n3093), .ZN(U3559) );
  INV_X1 U3954 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n3692) );
  NAND2_X1 U3955 ( .A1(n4710), .A2(U4043), .ZN(n3094) );
  OAI21_X1 U3956 ( .B1(U4043), .B2(n3692), .A(n3094), .ZN(U3569) );
  INV_X1 U3957 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n3783) );
  NAND2_X1 U3958 ( .A1(n4402), .A2(U4043), .ZN(n3095) );
  OAI21_X1 U3959 ( .B1(U4043), .B2(n3783), .A(n3095), .ZN(U3568) );
  INV_X1 U3960 ( .A(n4679), .ZN(n3217) );
  INV_X1 U3961 ( .A(REG3_REG_5__SCAN_IN), .ZN(n3098) );
  NOR2_X1 U3962 ( .A1(STATE_REG_SCAN_IN), .A2(n3098), .ZN(n3254) );
  INV_X1 U3963 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n3811) );
  INV_X1 U3964 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3099) );
  MUX2_X1 U3965 ( .A(REG2_REG_5__SCAN_IN), .B(n3099), .S(n4679), .Z(n3111) );
  INV_X1 U3966 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3100) );
  MUX2_X1 U3967 ( .A(REG2_REG_2__SCAN_IN), .B(n3100), .S(n4681), .Z(n4157) );
  INV_X1 U3968 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3101) );
  AND2_X1 U3969 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4150)
         );
  NAND2_X1 U3970 ( .A1(n4682), .A2(REG2_REG_1__SCAN_IN), .ZN(n3102) );
  INV_X1 U3971 ( .A(n4705), .ZN(n3120) );
  XNOR2_X1 U3972 ( .A(n3105), .B(n4680), .ZN(n4166) );
  INV_X1 U3973 ( .A(REG2_REG_4__SCAN_IN), .ZN(n3107) );
  INV_X1 U3974 ( .A(n3105), .ZN(n3106) );
  INV_X1 U3975 ( .A(n4680), .ZN(n3123) );
  NOR2_X1 U3976 ( .A1(n4149), .A2(n3108), .ZN(n3109) );
  NAND2_X1 U3977 ( .A1(n3208), .A2(n3111), .ZN(n3110) );
  OAI211_X1 U3978 ( .C1(n3111), .C2(n3208), .A(n4833), .B(n3110), .ZN(n3112)
         );
  OAI21_X1 U3979 ( .B1(n4853), .B2(n3811), .A(n3112), .ZN(n3113) );
  NOR2_X1 U3980 ( .A1(n3254), .A2(n3113), .ZN(n3129) );
  MUX2_X1 U3981 ( .A(REG1_REG_5__SCAN_IN), .B(n3114), .S(n4679), .Z(n3127) );
  AND2_X1 U3982 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n4140)
         );
  NAND2_X1 U3983 ( .A1(n4139), .A2(n4140), .ZN(n4138) );
  NAND2_X1 U3984 ( .A1(n4682), .A2(REG1_REG_1__SCAN_IN), .ZN(n3117) );
  NAND2_X1 U3985 ( .A1(n4138), .A2(n3117), .ZN(n4153) );
  NAND2_X1 U3986 ( .A1(n4153), .A2(n4154), .ZN(n4152) );
  OAI21_X1 U3987 ( .B1(n3121), .B2(n3120), .A(n4701), .ZN(n3122) );
  XNOR2_X1 U3988 ( .A(n3122), .B(n4680), .ZN(n4167) );
  INV_X1 U3989 ( .A(n3122), .ZN(n3124) );
  OAI211_X1 U3990 ( .C1(n3127), .C2(n3126), .A(n4835), .B(n3219), .ZN(n3128)
         );
  OAI211_X1 U3991 ( .C1(n4838), .C2(n3217), .A(n3129), .B(n3128), .ZN(U3245)
         );
  INV_X1 U3992 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n3834) );
  NAND2_X1 U3993 ( .A1(n3991), .A2(U4043), .ZN(n3130) );
  OAI21_X1 U3994 ( .B1(U4043), .B2(n3834), .A(n3130), .ZN(U3579) );
  XOR2_X1 U3995 ( .A(n3132), .B(n3131), .Z(n4147) );
  AOI22_X1 U3996 ( .A1(n4711), .A2(n4133), .B1(n4147), .B2(n3968), .ZN(n3138)
         );
  INV_X1 U3997 ( .A(n3133), .ZN(n3134) );
  NAND2_X1 U3998 ( .A1(n3135), .A2(n3134), .ZN(n3171) );
  AOI22_X1 U3999 ( .A1(n4712), .A2(n3136), .B1(REG3_REG_0__SCAN_IN), .B2(n3171), .ZN(n3137) );
  NAND2_X1 U4000 ( .A1(n3138), .A2(n3137), .ZN(U3229) );
  XNOR2_X1 U4001 ( .A(n3139), .B(n3140), .ZN(n3144) );
  AOI22_X1 U4002 ( .A1(n4724), .A2(n2234), .B1(n3963), .B2(n3199), .ZN(n3143)
         );
  AOI22_X1 U4003 ( .A1(n4712), .A2(n3141), .B1(REG3_REG_1__SCAN_IN), .B2(n3171), .ZN(n3142) );
  OAI211_X1 U4004 ( .C1(n3144), .C2(n4719), .A(n3143), .B(n3142), .ZN(U3219)
         );
  INV_X1 U4005 ( .A(n3145), .ZN(n3147) );
  NAND3_X1 U4006 ( .A1(n3148), .A2(n3147), .A3(n3146), .ZN(n3149) );
  AND2_X1 U4007 ( .A1(n4457), .A2(n4695), .ZN(n3315) );
  INV_X1 U4008 ( .A(n3247), .ZN(n3150) );
  OAI21_X1 U4009 ( .B1(n4875), .B2(n3156), .A(n3150), .ZN(n4930) );
  OR2_X1 U4010 ( .A1(n4024), .A2(n3151), .ZN(n3152) );
  NAND2_X1 U4011 ( .A1(n3153), .A2(n3152), .ZN(n4931) );
  NAND2_X1 U4012 ( .A1(n2234), .A2(n4863), .ZN(n3155) );
  NAND2_X1 U4013 ( .A1(n3199), .A2(n4516), .ZN(n3154) );
  OAI211_X1 U4014 ( .C1(n3156), .C2(n4858), .A(n3155), .B(n3154), .ZN(n3157)
         );
  INV_X1 U4015 ( .A(n3157), .ZN(n3160) );
  XNOR2_X1 U4016 ( .A(n4024), .B(n4043), .ZN(n3158) );
  NAND2_X1 U4017 ( .A1(n3158), .A2(n4876), .ZN(n3159) );
  OAI211_X1 U4018 ( .C1(n4931), .C2(n4523), .A(n3160), .B(n3159), .ZN(n4933)
         );
  MUX2_X1 U4019 ( .A(n4933), .B(REG2_REG_1__SCAN_IN), .S(n4888), .Z(n3161) );
  INV_X1 U4020 ( .A(n3161), .ZN(n3166) );
  INV_X1 U4021 ( .A(n4931), .ZN(n3164) );
  OR2_X1 U4022 ( .A1(n3162), .A2(n4695), .ZN(n3264) );
  INV_X1 U4023 ( .A(n3264), .ZN(n3163) );
  NAND2_X1 U4024 ( .A1(n4457), .A2(n3163), .ZN(n4535) );
  INV_X1 U4025 ( .A(n4535), .ZN(n4884) );
  AOI22_X1 U4026 ( .A1(n3164), .A2(n4884), .B1(REG3_REG_1__SCAN_IN), .B2(n4883), .ZN(n3165) );
  OAI211_X1 U4027 ( .C1(n4503), .C2(n4930), .A(n3166), .B(n3165), .ZN(U3289)
         );
  INV_X1 U4028 ( .A(n3169), .ZN(n3170) );
  AOI21_X1 U4029 ( .B1(n3167), .B2(n3168), .A(n3170), .ZN(n3175) );
  AOI22_X1 U4030 ( .A1(n4712), .A2(n3172), .B1(REG3_REG_2__SCAN_IN), .B2(n3171), .ZN(n3174) );
  AOI22_X1 U4031 ( .A1(n4724), .A2(n4133), .B1(n4711), .B2(n4132), .ZN(n3173)
         );
  OAI211_X1 U4032 ( .C1(n3175), .C2(n4719), .A(n3174), .B(n3173), .ZN(U3234)
         );
  XNOR2_X1 U4033 ( .A(n3176), .B(n4022), .ZN(n4942) );
  XNOR2_X1 U4034 ( .A(n3177), .B(n4022), .ZN(n3181) );
  AOI22_X1 U4035 ( .A1(n3200), .A2(n4516), .B1(n3202), .B2(n4543), .ZN(n3178)
         );
  OAI21_X1 U4036 ( .B1(n3179), .B2(n4519), .A(n3178), .ZN(n3180) );
  AOI21_X1 U4037 ( .B1(n3181), .B2(n4876), .A(n3180), .ZN(n3182) );
  OAI21_X1 U4038 ( .B1(n4942), .B2(n4523), .A(n3182), .ZN(n4943) );
  NAND2_X1 U4039 ( .A1(n4943), .A2(n4530), .ZN(n3187) );
  AOI21_X1 U4040 ( .B1(n3202), .B2(n3183), .A(n3292), .ZN(n4945) );
  INV_X1 U4041 ( .A(n4888), .ZN(n4530) );
  INV_X1 U4042 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3184) );
  OAI22_X1 U40430 ( .A1(n4530), .A2(n3184), .B1(n4528), .B2(
        REG3_REG_3__SCAN_IN), .ZN(n3185) );
  AOI21_X1 U4044 ( .B1(n4945), .B2(n4871), .A(n3185), .ZN(n3186) );
  OAI211_X1 U4045 ( .C1(n4942), .C2(n4535), .A(n3187), .B(n3186), .ZN(U3287)
         );
  NAND2_X1 U4046 ( .A1(n3188), .A2(n3968), .ZN(n3196) );
  AOI21_X1 U4047 ( .B1(n3189), .B2(n3191), .A(n3190), .ZN(n3195) );
  AOI22_X1 U4048 ( .A1(n4724), .A2(n4132), .B1(n4711), .B2(n4131), .ZN(n3194)
         );
  AND2_X1 U4049 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n4165) );
  NOR2_X1 U4050 ( .A1(n3953), .A2(n3291), .ZN(n3192) );
  AOI211_X1 U4051 ( .C1(n3302), .C2(n3955), .A(n4165), .B(n3192), .ZN(n3193)
         );
  OAI211_X1 U4052 ( .C1(n3196), .C2(n3195), .A(n3194), .B(n3193), .ZN(U3227)
         );
  OAI21_X1 U4053 ( .B1(n3198), .B2(n3197), .A(n3189), .ZN(n3206) );
  AOI22_X1 U4054 ( .A1(n4711), .A2(n3200), .B1(n4724), .B2(n3199), .ZN(n3204)
         );
  INV_X1 U4055 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3201) );
  NOR2_X1 U4056 ( .A1(STATE_REG_SCAN_IN), .A2(n3201), .ZN(n4700) );
  AOI21_X1 U4057 ( .B1(n4712), .B2(n3202), .A(n4700), .ZN(n3203) );
  OAI211_X1 U4058 ( .C1(REG3_REG_3__SCAN_IN), .C2(n4728), .A(n3204), .B(n3203), 
        .ZN(n3205) );
  AOI21_X1 U4059 ( .B1(n3206), .B2(n3968), .A(n3205), .ZN(n3207) );
  INV_X1 U4060 ( .A(n3207), .ZN(U3215) );
  INV_X1 U4061 ( .A(n4678), .ZN(n3232) );
  NAND2_X1 U4062 ( .A1(n4746), .A2(n3209), .ZN(n3210) );
  INV_X1 U4063 ( .A(n4746), .ZN(n4924) );
  NAND2_X1 U4064 ( .A1(n3210), .A2(n4749), .ZN(n4761) );
  INV_X1 U4065 ( .A(n4754), .ZN(n4922) );
  INV_X1 U4066 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3317) );
  AOI22_X1 U4067 ( .A1(REG2_REG_7__SCAN_IN), .A2(n4754), .B1(n4922), .B2(n3317), .ZN(n4762) );
  NAND2_X1 U4068 ( .A1(REG2_REG_7__SCAN_IN), .A2(n4754), .ZN(n3211) );
  INV_X1 U4069 ( .A(n3222), .ZN(n4920) );
  NAND2_X1 U4070 ( .A1(n3222), .A2(n3212), .ZN(n3213) );
  INV_X1 U4071 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3214) );
  MUX2_X1 U4072 ( .A(REG2_REG_9__SCAN_IN), .B(n3214), .S(n4678), .Z(n3215) );
  OAI211_X1 U4073 ( .C1(n3216), .C2(n3215), .A(n4833), .B(n3384), .ZN(n3231)
         );
  AND2_X1 U4074 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n3425) );
  NAND2_X1 U4075 ( .A1(REG1_REG_6__SCAN_IN), .A2(n4748), .ZN(n4747) );
  NAND2_X1 U4076 ( .A1(n4746), .A2(n3220), .ZN(n3221) );
  NOR2_X1 U4077 ( .A1(n4920), .A2(n3223), .ZN(n3224) );
  NOR2_X1 U4078 ( .A1(n3224), .A2(n4765), .ZN(n3228) );
  NAND2_X1 U4079 ( .A1(n4678), .A2(REG1_REG_9__SCAN_IN), .ZN(n3391) );
  OR2_X1 U4080 ( .A1(n4678), .A2(REG1_REG_9__SCAN_IN), .ZN(n3225) );
  NAND2_X1 U4081 ( .A1(n3391), .A2(n3225), .ZN(n3227) );
  INV_X1 U4082 ( .A(n3392), .ZN(n3226) );
  AOI211_X1 U4083 ( .C1(n3228), .C2(n3227), .A(n3226), .B(n4839), .ZN(n3229)
         );
  AOI211_X1 U4084 ( .C1(n4825), .C2(ADDR_REG_9__SCAN_IN), .A(n3425), .B(n3229), 
        .ZN(n3230) );
  OAI211_X1 U4085 ( .C1(n4838), .C2(n3232), .A(n3231), .B(n3230), .ZN(U3249)
         );
  NAND2_X1 U4086 ( .A1(n3234), .A2(n4020), .ZN(n3235) );
  NAND2_X1 U4087 ( .A1(n3236), .A2(n3235), .ZN(n4939) );
  INV_X1 U4088 ( .A(n4939), .ZN(n3251) );
  XNOR2_X1 U4089 ( .A(n3238), .B(n3237), .ZN(n3244) );
  INV_X1 U4090 ( .A(n4523), .ZN(n4877) );
  NAND2_X1 U4091 ( .A1(n4939), .A2(n4877), .ZN(n3243) );
  NAND2_X1 U4092 ( .A1(n4133), .A2(n4863), .ZN(n3240) );
  NAND2_X1 U4093 ( .A1(n4132), .A2(n4516), .ZN(n3239) );
  OAI211_X1 U4094 ( .C1(n3246), .C2(n4858), .A(n3240), .B(n3239), .ZN(n3241)
         );
  INV_X1 U4095 ( .A(n3241), .ZN(n3242) );
  OAI211_X1 U4096 ( .C1(n3244), .C2(n4865), .A(n3243), .B(n3242), .ZN(n4937)
         );
  MUX2_X1 U4097 ( .A(n4937), .B(REG2_REG_2__SCAN_IN), .S(n4888), .Z(n3245) );
  INV_X1 U4098 ( .A(n3245), .ZN(n3250) );
  INV_X1 U4099 ( .A(n3183), .ZN(n4935) );
  NOR2_X1 U4100 ( .A1(n3247), .A2(n3246), .ZN(n4936) );
  NOR3_X1 U4101 ( .A1(n4503), .A2(n4935), .A3(n4936), .ZN(n3248) );
  AOI21_X1 U4102 ( .B1(n4883), .B2(REG3_REG_2__SCAN_IN), .A(n3248), .ZN(n3249)
         );
  OAI211_X1 U4103 ( .C1(n3251), .C2(n4535), .A(n3250), .B(n3249), .ZN(U3288)
         );
  XNOR2_X1 U4104 ( .A(n3253), .B(n3252), .ZN(n3261) );
  INV_X1 U4105 ( .A(n3254), .ZN(n3255) );
  OAI21_X1 U4106 ( .B1(n3953), .B2(n3256), .A(n3255), .ZN(n3259) );
  OAI22_X1 U4107 ( .A1(n3276), .A2(n3514), .B1(n3515), .B2(n3257), .ZN(n3258)
         );
  AOI211_X1 U4108 ( .C1(n3267), .C2(n3955), .A(n3259), .B(n3258), .ZN(n3260)
         );
  OAI21_X1 U4109 ( .B1(n3261), .B2(n4719), .A(n3260), .ZN(U3224) );
  INV_X1 U4110 ( .A(n3263), .ZN(n4056) );
  XOR2_X1 U4111 ( .A(n3262), .B(n4021), .Z(n4953) );
  NAND2_X1 U4112 ( .A1(n4523), .A2(n3264), .ZN(n3265) );
  AOI21_X1 U4113 ( .B1(n3273), .B2(n3266), .A(n3332), .ZN(n4956) );
  INV_X1 U4114 ( .A(n3267), .ZN(n3268) );
  OAI22_X1 U4115 ( .A1(n4530), .A2(n3099), .B1(n3268), .B2(n4528), .ZN(n3269)
         );
  AOI21_X1 U4116 ( .B1(n4956), .B2(n4871), .A(n3269), .ZN(n3278) );
  INV_X1 U4117 ( .A(n4021), .ZN(n3270) );
  XNOR2_X1 U4118 ( .A(n3271), .B(n3270), .ZN(n3272) );
  NAND2_X1 U4119 ( .A1(n3272), .A2(n4876), .ZN(n3275) );
  AOI22_X1 U4120 ( .A1(n3503), .A2(n4516), .B1(n3273), .B2(n4543), .ZN(n3274)
         );
  OAI211_X1 U4121 ( .C1(n3276), .C2(n4519), .A(n3275), .B(n3274), .ZN(n4955)
         );
  NAND2_X1 U4122 ( .A1(n4955), .A2(n4530), .ZN(n3277) );
  OAI211_X1 U4123 ( .C1(n4953), .C2(n4506), .A(n3278), .B(n3277), .ZN(U3285)
         );
  NAND2_X1 U4124 ( .A1(n3282), .A2(n3281), .ZN(n3283) );
  XNOR2_X1 U4125 ( .A(n3280), .B(n3283), .ZN(n3290) );
  INV_X1 U4126 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3691) );
  NOR2_X1 U4127 ( .A1(STATE_REG_SCAN_IN), .A2(n3691), .ZN(n4745) );
  INV_X1 U4128 ( .A(n4745), .ZN(n3284) );
  OAI21_X1 U4129 ( .B1(n3953), .B2(n2271), .A(n3284), .ZN(n3287) );
  OAI22_X1 U4130 ( .A1(n3328), .A2(n3514), .B1(n3515), .B2(n3285), .ZN(n3286)
         );
  AOI211_X1 U4131 ( .C1(n3288), .C2(n3955), .A(n3287), .B(n3286), .ZN(n3289)
         );
  OAI21_X1 U4132 ( .B1(n3290), .B2(n4719), .A(n3289), .ZN(U3236) );
  OAI211_X1 U4133 ( .C1(n3292), .C2(n3291), .A(n3266), .B(n4971), .ZN(n4947)
         );
  NOR2_X1 U4134 ( .A1(n4947), .A2(n4685), .ZN(n3301) );
  XNOR2_X1 U4135 ( .A(n3293), .B(n4023), .ZN(n3303) );
  XOR2_X1 U4136 ( .A(n3294), .B(n4023), .Z(n3299) );
  AOI22_X1 U4137 ( .A1(n4131), .A2(n4516), .B1(n3295), .B2(n4543), .ZN(n3296)
         );
  OAI21_X1 U4138 ( .B1(n3297), .B2(n4519), .A(n3296), .ZN(n3298) );
  AOI21_X1 U4139 ( .B1(n3299), .B2(n4876), .A(n3298), .ZN(n3300) );
  OAI21_X1 U4140 ( .B1(n3303), .B2(n4523), .A(n3300), .ZN(n4948) );
  AOI211_X1 U4141 ( .C1(n4883), .C2(n3302), .A(n3301), .B(n4948), .ZN(n3305)
         );
  INV_X1 U4142 ( .A(n3303), .ZN(n4950) );
  AOI22_X1 U4143 ( .A1(n4950), .A2(n4884), .B1(REG2_REG_4__SCAN_IN), .B2(n4888), .ZN(n3304) );
  OAI21_X1 U4144 ( .B1(n3305), .B2(n4888), .A(n3304), .ZN(U3286) );
  INV_X1 U4145 ( .A(n4030), .ZN(n4060) );
  XNOR2_X1 U4146 ( .A(n3306), .B(n4060), .ZN(n3310) );
  NAND2_X1 U4147 ( .A1(n3503), .A2(n4863), .ZN(n3308) );
  NAND2_X1 U4148 ( .A1(n3502), .A2(n4516), .ZN(n3307) );
  OAI211_X1 U4149 ( .C1(n3504), .C2(n4858), .A(n3308), .B(n3307), .ZN(n3309)
         );
  AOI21_X1 U4150 ( .B1(n3310), .B2(n4876), .A(n3309), .ZN(n4961) );
  XNOR2_X1 U4151 ( .A(n3311), .B(n4060), .ZN(n4958) );
  NAND2_X1 U4152 ( .A1(n3331), .A2(n3312), .ZN(n3313) );
  NAND2_X1 U4153 ( .A1(n3313), .A2(n4971), .ZN(n3314) );
  OR2_X1 U4154 ( .A1(n3314), .A2(n3364), .ZN(n4959) );
  INV_X1 U4155 ( .A(n3315), .ZN(n4429) );
  NOR2_X1 U4156 ( .A1(n4959), .A2(n4429), .ZN(n3319) );
  INV_X1 U4157 ( .A(n3506), .ZN(n3316) );
  OAI22_X1 U4158 ( .A1(n4530), .A2(n3317), .B1(n3316), .B2(n4528), .ZN(n3318)
         );
  AOI211_X1 U4159 ( .C1(n4958), .C2(n4431), .A(n3319), .B(n3318), .ZN(n3320)
         );
  OAI21_X1 U4160 ( .B1(n4888), .B2(n4961), .A(n3320), .ZN(U3283) );
  NAND2_X1 U4161 ( .A1(n4059), .A2(n4068), .ZN(n4028) );
  OR2_X1 U4162 ( .A1(n3262), .A2(n3321), .ZN(n3323) );
  NAND2_X1 U4163 ( .A1(n3323), .A2(n3322), .ZN(n3324) );
  XOR2_X1 U4164 ( .A(n4028), .B(n3324), .Z(n3341) );
  XOR2_X1 U4165 ( .A(n4028), .B(n3325), .Z(n3330) );
  AOI22_X1 U4166 ( .A1(n4130), .A2(n4516), .B1(n3326), .B2(n4543), .ZN(n3327)
         );
  OAI21_X1 U4167 ( .B1(n3328), .B2(n4519), .A(n3327), .ZN(n3329) );
  AOI21_X1 U4168 ( .B1(n3330), .B2(n4876), .A(n3329), .ZN(n3346) );
  OAI21_X1 U4169 ( .B1(n3341), .B2(n4952), .A(n3346), .ZN(n3337) );
  OAI21_X1 U4170 ( .B1(n3332), .B2(n2271), .A(n3331), .ZN(n3339) );
  OAI22_X1 U4171 ( .A1(n3339), .A2(n4618), .B1(n4990), .B2(n2532), .ZN(n3333)
         );
  AOI21_X1 U4172 ( .B1(n3337), .B2(n4990), .A(n3333), .ZN(n3334) );
  INV_X1 U4173 ( .A(n3334), .ZN(U3524) );
  INV_X1 U4174 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3335) );
  OAI22_X1 U4175 ( .A1(n3339), .A2(n4671), .B1(n4978), .B2(n3335), .ZN(n3336)
         );
  AOI21_X1 U4176 ( .B1(n3337), .B2(n4978), .A(n3336), .ZN(n3338) );
  INV_X1 U4177 ( .A(n3338), .ZN(U3479) );
  INV_X1 U4178 ( .A(n3339), .ZN(n3344) );
  OAI22_X1 U4179 ( .A1(n4530), .A2(n3773), .B1(n3340), .B2(n4528), .ZN(n3343)
         );
  NOR2_X1 U4180 ( .A1(n3341), .A2(n4506), .ZN(n3342) );
  AOI211_X1 U4181 ( .C1(n3344), .C2(n4871), .A(n3343), .B(n3342), .ZN(n3345)
         );
  OAI21_X1 U4182 ( .B1(n4888), .B2(n3346), .A(n3345), .ZN(U3284) );
  XOR2_X1 U4183 ( .A(n3349), .B(n3348), .Z(n3350) );
  XNOR2_X1 U4184 ( .A(n3347), .B(n3350), .ZN(n3355) );
  AOI22_X1 U4185 ( .A1(n4724), .A2(n4130), .B1(n3963), .B2(n3432), .ZN(n3354)
         );
  INV_X1 U4186 ( .A(REG3_REG_8__SCAN_IN), .ZN(n3351) );
  NOR2_X1 U4187 ( .A1(STATE_REG_SCAN_IN), .A2(n3351), .ZN(n4768) );
  NOR2_X1 U4188 ( .A1(n3953), .A2(n3363), .ZN(n3352) );
  AOI211_X1 U4189 ( .C1(n3366), .C2(n3955), .A(n4768), .B(n3352), .ZN(n3353)
         );
  OAI211_X1 U4190 ( .C1(n3355), .C2(n4719), .A(n3354), .B(n3353), .ZN(U3218)
         );
  NAND2_X1 U4191 ( .A1(n4064), .A2(n4069), .ZN(n4029) );
  XOR2_X1 U4192 ( .A(n4029), .B(n3356), .Z(n3360) );
  OAI22_X1 U4193 ( .A1(n3357), .A2(n4878), .B1(n3363), .B2(n4858), .ZN(n3358)
         );
  AOI21_X1 U4194 ( .B1(n4863), .B2(n4130), .A(n3358), .ZN(n3359) );
  OAI21_X1 U4195 ( .B1(n3360), .B2(n4865), .A(n3359), .ZN(n3402) );
  INV_X1 U4196 ( .A(n3402), .ZN(n3370) );
  XOR2_X1 U4197 ( .A(n4029), .B(n3361), .Z(n3403) );
  OR2_X1 U4198 ( .A1(n3364), .A2(n3363), .ZN(n3365) );
  NAND2_X1 U4199 ( .A1(n3362), .A2(n3365), .ZN(n3408) );
  AOI22_X1 U4200 ( .A1(n4888), .A2(REG2_REG_8__SCAN_IN), .B1(n3366), .B2(n4883), .ZN(n3367) );
  OAI21_X1 U4201 ( .B1(n3408), .B2(n4503), .A(n3367), .ZN(n3368) );
  AOI21_X1 U4202 ( .B1(n3403), .B2(n4431), .A(n3368), .ZN(n3369) );
  OAI21_X1 U4203 ( .B1(n3370), .B2(n4888), .A(n3369), .ZN(U3282) );
  INV_X1 U4204 ( .A(n4077), .ZN(n3371) );
  NAND2_X1 U4205 ( .A1(n3371), .A2(n4063), .ZN(n4016) );
  XNOR2_X1 U4206 ( .A(n3372), .B(n4016), .ZN(n3377) );
  AOI22_X1 U4207 ( .A1(n4862), .A2(n4516), .B1(n3373), .B2(n4543), .ZN(n3374)
         );
  OAI21_X1 U4208 ( .B1(n3375), .B2(n4519), .A(n3374), .ZN(n3376) );
  AOI21_X1 U4209 ( .B1(n3377), .B2(n4876), .A(n3376), .ZN(n4963) );
  XNOR2_X1 U4210 ( .A(n3378), .B(n4016), .ZN(n4967) );
  INV_X1 U4211 ( .A(n3362), .ZN(n3379) );
  OAI21_X1 U4212 ( .B1(n3379), .B2(n3423), .A(n3436), .ZN(n4964) );
  NOR2_X1 U4213 ( .A1(n4964), .A2(n4503), .ZN(n3382) );
  INV_X1 U4214 ( .A(n3426), .ZN(n3380) );
  OAI22_X1 U4215 ( .A1(n4530), .A2(n3214), .B1(n3380), .B2(n4528), .ZN(n3381)
         );
  AOI211_X1 U4216 ( .C1(n4967), .C2(n4431), .A(n3382), .B(n3381), .ZN(n3383)
         );
  OAI21_X1 U4217 ( .B1(n4888), .B2(n4963), .A(n3383), .ZN(U3281) );
  INV_X1 U4218 ( .A(n4677), .ZN(n4187) );
  NAND2_X1 U4219 ( .A1(n4678), .A2(REG2_REG_9__SCAN_IN), .ZN(n3385) );
  NAND2_X1 U4220 ( .A1(n4917), .A2(n3386), .ZN(n3387) );
  XNOR2_X1 U4221 ( .A(n3386), .B(n3393), .ZN(n4778) );
  NAND2_X1 U4222 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4778), .ZN(n4777) );
  NAND2_X1 U4223 ( .A1(n3387), .A2(n4777), .ZN(n3390) );
  INV_X1 U4224 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3388) );
  MUX2_X1 U4225 ( .A(REG2_REG_11__SCAN_IN), .B(n3388), .S(n4677), .Z(n3389) );
  NAND2_X1 U4226 ( .A1(n3390), .A2(n3389), .ZN(n4189) );
  OAI211_X1 U4227 ( .C1(n3390), .C2(n3389), .A(n4189), .B(n4833), .ZN(n3401)
         );
  NOR2_X1 U4228 ( .A1(STATE_REG_SCAN_IN), .A2(n3695), .ZN(n3449) );
  NOR2_X1 U4229 ( .A1(n2245), .A2(n3393), .ZN(n3394) );
  MUX2_X1 U4230 ( .A(n3395), .B(REG1_REG_11__SCAN_IN), .S(n4677), .Z(n3397) );
  INV_X1 U4231 ( .A(n4174), .ZN(n3396) );
  AOI211_X1 U4232 ( .C1(n3398), .C2(n3397), .A(n3396), .B(n4839), .ZN(n3399)
         );
  AOI211_X1 U4233 ( .C1(n4825), .C2(ADDR_REG_11__SCAN_IN), .A(n3449), .B(n3399), .ZN(n3400) );
  OAI211_X1 U4234 ( .C1(n4838), .C2(n4187), .A(n3401), .B(n3400), .ZN(U3251)
         );
  AOI21_X1 U4235 ( .B1(n3403), .B2(n4968), .A(n3402), .ZN(n3405) );
  MUX2_X1 U4236 ( .A(n2568), .B(n3405), .S(n4990), .Z(n3404) );
  OAI21_X1 U4237 ( .B1(n3408), .B2(n4618), .A(n3404), .ZN(U3526) );
  INV_X1 U4238 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3406) );
  MUX2_X1 U4239 ( .A(n3406), .B(n3405), .S(n4978), .Z(n3407) );
  OAI21_X1 U4240 ( .B1(n3408), .B2(n4671), .A(n3407), .ZN(U3483) );
  NAND2_X1 U4241 ( .A1(n3409), .A2(n3968), .ZN(n3419) );
  AOI21_X1 U4242 ( .B1(n3411), .B2(n3413), .A(n3412), .ZN(n3418) );
  AOI22_X1 U4243 ( .A1(n4724), .A2(n3432), .B1(n3963), .B2(n4129), .ZN(n3417)
         );
  NOR2_X1 U4244 ( .A1(STATE_REG_SCAN_IN), .A2(n3414), .ZN(n4775) );
  NOR2_X1 U4245 ( .A1(n3953), .A2(n3437), .ZN(n3415) );
  AOI211_X1 U4246 ( .C1(n3439), .C2(n3955), .A(n4775), .B(n3415), .ZN(n3416)
         );
  OAI211_X1 U4247 ( .C1(n3419), .C2(n3418), .A(n3417), .B(n3416), .ZN(U3214)
         );
  INV_X1 U4248 ( .A(n3411), .ZN(n3420) );
  AOI21_X1 U4249 ( .B1(n3422), .B2(n3421), .A(n3420), .ZN(n3429) );
  AOI22_X1 U4250 ( .A1(n4724), .A2(n3502), .B1(n4711), .B2(n4862), .ZN(n3428)
         );
  NOR2_X1 U4251 ( .A1(n3953), .A2(n3423), .ZN(n3424) );
  AOI211_X1 U4252 ( .C1(n3426), .C2(n3955), .A(n3425), .B(n3424), .ZN(n3427)
         );
  OAI211_X1 U4253 ( .C1(n3429), .C2(n4719), .A(n3428), .B(n3427), .ZN(U3228)
         );
  NAND2_X1 U4254 ( .A1(n4076), .A2(n4079), .ZN(n4014) );
  XNOR2_X1 U4255 ( .A(n3430), .B(n4014), .ZN(n3434) );
  OAI22_X1 U4256 ( .A1(n3463), .A2(n4878), .B1(n3437), .B2(n4858), .ZN(n3431)
         );
  AOI21_X1 U4257 ( .B1(n4863), .B2(n3432), .A(n3431), .ZN(n3433) );
  OAI21_X1 U4258 ( .B1(n3434), .B2(n4865), .A(n3433), .ZN(n3453) );
  INV_X1 U4259 ( .A(n3453), .ZN(n3443) );
  XOR2_X1 U4260 ( .A(n4014), .B(n3435), .Z(n3454) );
  INV_X1 U4261 ( .A(n3436), .ZN(n3438) );
  OAI21_X1 U4262 ( .B1(n3438), .B2(n3437), .A(n2269), .ZN(n3459) );
  AOI22_X1 U4263 ( .A1(n4888), .A2(REG2_REG_10__SCAN_IN), .B1(n3439), .B2(
        n4883), .ZN(n3440) );
  OAI21_X1 U4264 ( .B1(n3459), .B2(n4503), .A(n3440), .ZN(n3441) );
  AOI21_X1 U4265 ( .B1(n3454), .B2(n4431), .A(n3441), .ZN(n3442) );
  OAI21_X1 U4266 ( .B1(n4888), .B2(n3443), .A(n3442), .ZN(U3280) );
  NAND2_X1 U4267 ( .A1(n3445), .A2(n3444), .ZN(n3447) );
  XOR2_X1 U4268 ( .A(n3447), .B(n3446), .Z(n3452) );
  AOI22_X1 U4269 ( .A1(n4724), .A2(n4862), .B1(n4711), .B2(n4128), .ZN(n3451)
         );
  NOR2_X1 U4270 ( .A1(n3953), .A2(n4859), .ZN(n3448) );
  AOI211_X1 U4271 ( .C1(n4868), .C2(n3955), .A(n3449), .B(n3448), .ZN(n3450)
         );
  OAI211_X1 U4272 ( .C1(n3452), .C2(n4719), .A(n3451), .B(n3450), .ZN(U3233)
         );
  INV_X1 U4273 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3455) );
  AOI21_X1 U4274 ( .B1(n3454), .B2(n4968), .A(n3453), .ZN(n3457) );
  MUX2_X1 U4275 ( .A(n3455), .B(n3457), .S(n4978), .Z(n3456) );
  OAI21_X1 U4276 ( .B1(n3459), .B2(n4671), .A(n3456), .ZN(U3487) );
  MUX2_X1 U4277 ( .A(n2604), .B(n3457), .S(n4990), .Z(n3458) );
  OAI21_X1 U4278 ( .B1(n3459), .B2(n4618), .A(n3458), .ZN(U3528) );
  XNOR2_X1 U4279 ( .A(n3938), .B(n3461), .ZN(n3462) );
  XNOR2_X1 U4280 ( .A(n3460), .B(n3462), .ZN(n3467) );
  NAND2_X1 U4281 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4783) );
  OAI21_X1 U4282 ( .B1(n3953), .B2(n3476), .A(n4783), .ZN(n3465) );
  OAI22_X1 U4283 ( .A1(n4497), .A2(n3515), .B1(n3514), .B2(n3463), .ZN(n3464)
         );
  AOI211_X1 U4284 ( .C1(n3478), .C2(n3955), .A(n3465), .B(n3464), .ZN(n3466)
         );
  OAI21_X1 U4285 ( .B1(n3467), .B2(n4719), .A(n3466), .ZN(U3221) );
  INV_X1 U4286 ( .A(n3468), .ZN(n4857) );
  AOI21_X1 U4287 ( .B1(n4857), .B2(n3470), .A(n3469), .ZN(n4512) );
  NAND2_X1 U4288 ( .A1(n4509), .A2(n4510), .ZN(n4015) );
  XNOR2_X1 U4289 ( .A(n4512), .B(n4015), .ZN(n3473) );
  OAI22_X1 U4290 ( .A1(n4497), .A2(n4878), .B1(n3476), .B2(n4858), .ZN(n3471)
         );
  AOI21_X1 U4291 ( .B1(n4863), .B2(n4129), .A(n3471), .ZN(n3472) );
  OAI21_X1 U4292 ( .B1(n3473), .B2(n4865), .A(n3472), .ZN(n4615) );
  INV_X1 U4293 ( .A(n4615), .ZN(n3482) );
  XNOR2_X1 U4294 ( .A(n3474), .B(n4015), .ZN(n4616) );
  OR2_X1 U4295 ( .A1(n4869), .A2(n3476), .ZN(n3477) );
  NAND2_X1 U4296 ( .A1(n3475), .A2(n3477), .ZN(n4672) );
  AOI22_X1 U4297 ( .A1(n4888), .A2(REG2_REG_12__SCAN_IN), .B1(n3478), .B2(
        n4883), .ZN(n3479) );
  OAI21_X1 U4298 ( .B1(n4672), .B2(n4503), .A(n3479), .ZN(n3480) );
  AOI21_X1 U4299 ( .B1(n4616), .B2(n4431), .A(n3480), .ZN(n3481) );
  OAI21_X1 U4300 ( .B1(n4888), .B2(n3482), .A(n3481), .ZN(U3278) );
  NAND3_X1 U4301 ( .A1(n2390), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3484) );
  INV_X1 U4302 ( .A(DATAI_31_), .ZN(n3483) );
  OAI22_X1 U4303 ( .A1(n3485), .A2(n3484), .B1(STATE_REG_SCAN_IN), .B2(n3483), 
        .ZN(U3321) );
  INV_X1 U4304 ( .A(REG0_REG_31__SCAN_IN), .ZN(n3497) );
  INV_X1 U4305 ( .A(n4008), .ZN(n3494) );
  NAND2_X1 U4306 ( .A1(n2233), .A2(DATAI_29_), .ZN(n3990) );
  INV_X1 U4307 ( .A(n4544), .ZN(n3971) );
  NAND2_X1 U4308 ( .A1(n4539), .A2(n3971), .ZN(n4540) );
  INV_X1 U4309 ( .A(n4671), .ZN(n3486) );
  NAND2_X1 U4310 ( .A1(n4730), .A2(n3486), .ZN(n3496) );
  NAND2_X1 U4311 ( .A1(n2996), .A2(REG2_REG_31__SCAN_IN), .ZN(n3492) );
  NAND2_X1 U4312 ( .A1(n3487), .A2(REG0_REG_31__SCAN_IN), .ZN(n3491) );
  INV_X1 U4313 ( .A(REG1_REG_31__SCAN_IN), .ZN(n3488) );
  OR2_X1 U4314 ( .A1(n3489), .A2(n3488), .ZN(n3490) );
  NAND2_X1 U4315 ( .A1(n4737), .A2(B_REG_SCAN_IN), .ZN(n3493) );
  AND2_X1 U4316 ( .A1(n4516), .A2(n3493), .ZN(n4211) );
  NAND2_X1 U4317 ( .A1(n4124), .A2(n4211), .ZN(n4546) );
  OAI21_X1 U4318 ( .B1(n3494), .B2(n4858), .A(n4546), .ZN(n4729) );
  NAND2_X1 U4319 ( .A1(n4978), .A2(n4729), .ZN(n3495) );
  OAI211_X1 U4320 ( .C1(n4978), .C2(n3497), .A(n3496), .B(n3495), .ZN(U3517)
         );
  AOI21_X1 U4321 ( .B1(n3499), .B2(n3498), .A(n4719), .ZN(n3501) );
  NAND2_X1 U4322 ( .A1(n3501), .A2(n3500), .ZN(n3509) );
  AOI22_X1 U4323 ( .A1(n4724), .A2(n3503), .B1(n4711), .B2(n3502), .ZN(n3508)
         );
  AND2_X1 U4324 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n4759) );
  NOR2_X1 U4325 ( .A1(n3953), .A2(n3504), .ZN(n3505) );
  AOI211_X1 U4326 ( .C1(n3506), .C2(n3955), .A(n4759), .B(n3505), .ZN(n3507)
         );
  NAND3_X1 U4327 ( .A1(n3509), .A2(n3508), .A3(n3507), .ZN(U3210) );
  XNOR2_X1 U4328 ( .A(n2236), .B(n3511), .ZN(n3512) );
  XNOR2_X1 U4329 ( .A(n3510), .B(n3512), .ZN(n3519) );
  NAND2_X1 U4330 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4810) );
  OAI21_X1 U4331 ( .B1(n3953), .B2(n3513), .A(n4810), .ZN(n3517) );
  OAI22_X1 U4332 ( .A1(n4465), .A2(n3515), .B1(n3514), .B2(n4497), .ZN(n3516)
         );
  AOI211_X1 U4333 ( .C1(n4501), .C2(n3955), .A(n3517), .B(n3516), .ZN(n3518)
         );
  OAI21_X1 U4334 ( .B1(n3519), .B2(n4719), .A(n3518), .ZN(U3212) );
  INV_X1 U4335 ( .A(D_REG_18__SCAN_IN), .ZN(n4897) );
  AOI22_X1 U4336 ( .A1(n4897), .A2(keyinput204), .B1(n4895), .B2(keyinput139), 
        .ZN(n3520) );
  OAI221_X1 U4337 ( .B1(n4897), .B2(keyinput204), .C1(n4895), .C2(keyinput139), 
        .A(n3520), .ZN(n3533) );
  INV_X1 U4338 ( .A(REG3_REG_1__SCAN_IN), .ZN(n4135) );
  AOI22_X1 U4339 ( .A1(n4135), .A2(keyinput153), .B1(n3917), .B2(keyinput141), 
        .ZN(n3521) );
  OAI221_X1 U4340 ( .B1(n4135), .B2(keyinput153), .C1(n3917), .C2(keyinput141), 
        .A(n3521), .ZN(n3532) );
  XNOR2_X1 U4341 ( .A(IR_REG_11__SCAN_IN), .B(keyinput220), .ZN(n3525) );
  XNOR2_X1 U4342 ( .A(IR_REG_19__SCAN_IN), .B(keyinput234), .ZN(n3524) );
  XNOR2_X1 U4343 ( .A(IR_REG_18__SCAN_IN), .B(keyinput130), .ZN(n3523) );
  XNOR2_X1 U4344 ( .A(IR_REG_27__SCAN_IN), .B(keyinput229), .ZN(n3522) );
  NAND4_X1 U4345 ( .A1(n3525), .A2(n3524), .A3(n3523), .A4(n3522), .ZN(n3531)
         );
  XNOR2_X1 U4346 ( .A(REG3_REG_17__SCAN_IN), .B(keyinput167), .ZN(n3529) );
  XNOR2_X1 U4347 ( .A(IR_REG_9__SCAN_IN), .B(keyinput218), .ZN(n3528) );
  XNOR2_X1 U4348 ( .A(IR_REG_5__SCAN_IN), .B(keyinput209), .ZN(n3527) );
  XNOR2_X1 U4349 ( .A(IR_REG_17__SCAN_IN), .B(keyinput237), .ZN(n3526) );
  NAND4_X1 U4350 ( .A1(n3529), .A2(n3528), .A3(n3527), .A4(n3526), .ZN(n3530)
         );
  OR4_X1 U4351 ( .A1(n3533), .A2(n3532), .A3(n3531), .A4(n3530), .ZN(n3575) );
  AOI22_X1 U4352 ( .A1(REG1_REG_15__SCAN_IN), .A2(keyinput140), .B1(
        REG1_REG_13__SCAN_IN), .B2(keyinput195), .ZN(n3534) );
  OAI221_X1 U4353 ( .B1(REG1_REG_15__SCAN_IN), .B2(keyinput140), .C1(
        REG1_REG_13__SCAN_IN), .C2(keyinput195), .A(n3534), .ZN(n3541) );
  AOI22_X1 U4354 ( .A1(REG1_REG_14__SCAN_IN), .A2(keyinput187), .B1(
        REG1_REG_16__SCAN_IN), .B2(keyinput180), .ZN(n3535) );
  OAI221_X1 U4355 ( .B1(REG1_REG_14__SCAN_IN), .B2(keyinput187), .C1(
        REG1_REG_16__SCAN_IN), .C2(keyinput180), .A(n3535), .ZN(n3540) );
  AOI22_X1 U4356 ( .A1(REG1_REG_18__SCAN_IN), .A2(keyinput230), .B1(
        REG1_REG_21__SCAN_IN), .B2(keyinput250), .ZN(n3536) );
  OAI221_X1 U4357 ( .B1(REG1_REG_18__SCAN_IN), .B2(keyinput230), .C1(
        REG1_REG_21__SCAN_IN), .C2(keyinput250), .A(n3536), .ZN(n3539) );
  AOI22_X1 U4358 ( .A1(REG1_REG_25__SCAN_IN), .A2(keyinput169), .B1(
        REG1_REG_29__SCAN_IN), .B2(keyinput223), .ZN(n3537) );
  OAI221_X1 U4359 ( .B1(REG1_REG_25__SCAN_IN), .B2(keyinput169), .C1(
        REG1_REG_29__SCAN_IN), .C2(keyinput223), .A(n3537), .ZN(n3538) );
  NOR4_X1 U4360 ( .A1(n3541), .A2(n3540), .A3(n3539), .A4(n3538), .ZN(n3569)
         );
  AOI22_X1 U4361 ( .A1(REG2_REG_4__SCAN_IN), .A2(keyinput163), .B1(
        REG2_REG_6__SCAN_IN), .B2(keyinput249), .ZN(n3542) );
  OAI221_X1 U4362 ( .B1(REG2_REG_4__SCAN_IN), .B2(keyinput163), .C1(
        REG2_REG_6__SCAN_IN), .C2(keyinput249), .A(n3542), .ZN(n3549) );
  AOI22_X1 U4363 ( .A1(REG2_REG_7__SCAN_IN), .A2(keyinput174), .B1(
        REG2_REG_8__SCAN_IN), .B2(keyinput217), .ZN(n3543) );
  OAI221_X1 U4364 ( .B1(REG2_REG_7__SCAN_IN), .B2(keyinput174), .C1(
        REG2_REG_8__SCAN_IN), .C2(keyinput217), .A(n3543), .ZN(n3548) );
  AOI22_X1 U4365 ( .A1(REG2_REG_15__SCAN_IN), .A2(keyinput194), .B1(
        REG2_REG_11__SCAN_IN), .B2(keyinput208), .ZN(n3544) );
  OAI221_X1 U4366 ( .B1(REG2_REG_15__SCAN_IN), .B2(keyinput194), .C1(
        REG2_REG_11__SCAN_IN), .C2(keyinput208), .A(n3544), .ZN(n3547) );
  AOI22_X1 U4367 ( .A1(REG2_REG_24__SCAN_IN), .A2(keyinput171), .B1(
        REG2_REG_18__SCAN_IN), .B2(keyinput142), .ZN(n3545) );
  OAI221_X1 U4368 ( .B1(REG2_REG_24__SCAN_IN), .B2(keyinput171), .C1(
        REG2_REG_18__SCAN_IN), .C2(keyinput142), .A(n3545), .ZN(n3546) );
  NOR4_X1 U4369 ( .A1(n3549), .A2(n3548), .A3(n3547), .A4(n3546), .ZN(n3568)
         );
  AOI22_X1 U4370 ( .A1(REG2_REG_22__SCAN_IN), .A2(keyinput241), .B1(
        REG2_REG_25__SCAN_IN), .B2(keyinput160), .ZN(n3550) );
  OAI221_X1 U4371 ( .B1(REG2_REG_22__SCAN_IN), .B2(keyinput241), .C1(
        REG2_REG_25__SCAN_IN), .C2(keyinput160), .A(n3550), .ZN(n3557) );
  AOI22_X1 U4372 ( .A1(ADDR_REG_15__SCAN_IN), .A2(keyinput137), .B1(
        REG2_REG_31__SCAN_IN), .B2(keyinput227), .ZN(n3551) );
  OAI221_X1 U4373 ( .B1(ADDR_REG_15__SCAN_IN), .B2(keyinput137), .C1(
        REG2_REG_31__SCAN_IN), .C2(keyinput227), .A(n3551), .ZN(n3556) );
  AOI22_X1 U4374 ( .A1(ADDR_REG_7__SCAN_IN), .A2(keyinput207), .B1(
        ADDR_REG_14__SCAN_IN), .B2(keyinput146), .ZN(n3552) );
  OAI221_X1 U4375 ( .B1(ADDR_REG_7__SCAN_IN), .B2(keyinput207), .C1(
        ADDR_REG_14__SCAN_IN), .C2(keyinput146), .A(n3552), .ZN(n3555) );
  AOI22_X1 U4376 ( .A1(ADDR_REG_4__SCAN_IN), .A2(keyinput135), .B1(
        ADDR_REG_8__SCAN_IN), .B2(keyinput155), .ZN(n3553) );
  OAI221_X1 U4377 ( .B1(ADDR_REG_4__SCAN_IN), .B2(keyinput135), .C1(
        ADDR_REG_8__SCAN_IN), .C2(keyinput155), .A(n3553), .ZN(n3554) );
  NOR4_X1 U4378 ( .A1(n3557), .A2(n3556), .A3(n3555), .A4(n3554), .ZN(n3567)
         );
  AOI22_X1 U4379 ( .A1(DATAO_REG_4__SCAN_IN), .A2(keyinput239), .B1(
        DATAO_REG_0__SCAN_IN), .B2(keyinput131), .ZN(n3558) );
  OAI221_X1 U4380 ( .B1(DATAO_REG_4__SCAN_IN), .B2(keyinput239), .C1(
        DATAO_REG_0__SCAN_IN), .C2(keyinput131), .A(n3558), .ZN(n3565) );
  AOI22_X1 U4381 ( .A1(DATAO_REG_6__SCAN_IN), .A2(keyinput201), .B1(
        DATAO_REG_8__SCAN_IN), .B2(keyinput184), .ZN(n3559) );
  OAI221_X1 U4382 ( .B1(DATAO_REG_6__SCAN_IN), .B2(keyinput201), .C1(
        DATAO_REG_8__SCAN_IN), .C2(keyinput184), .A(n3559), .ZN(n3564) );
  AOI22_X1 U4383 ( .A1(DATAO_REG_24__SCAN_IN), .A2(keyinput168), .B1(
        DATAO_REG_12__SCAN_IN), .B2(keyinput144), .ZN(n3560) );
  OAI221_X1 U4384 ( .B1(DATAO_REG_24__SCAN_IN), .B2(keyinput168), .C1(
        DATAO_REG_12__SCAN_IN), .C2(keyinput144), .A(n3560), .ZN(n3563) );
  AOI22_X1 U4385 ( .A1(DATAO_REG_28__SCAN_IN), .A2(keyinput232), .B1(
        D_REG_8__SCAN_IN), .B2(keyinput149), .ZN(n3561) );
  OAI221_X1 U4386 ( .B1(DATAO_REG_28__SCAN_IN), .B2(keyinput232), .C1(
        D_REG_8__SCAN_IN), .C2(keyinput149), .A(n3561), .ZN(n3562) );
  NOR4_X1 U4387 ( .A1(n3565), .A2(n3564), .A3(n3563), .A4(n3562), .ZN(n3566)
         );
  NAND4_X1 U4388 ( .A1(n3569), .A2(n3568), .A3(n3567), .A4(n3566), .ZN(n3574)
         );
  INV_X1 U4389 ( .A(D_REG_16__SCAN_IN), .ZN(n4898) );
  AOI22_X1 U4390 ( .A1(n4898), .A2(keyinput158), .B1(n4899), .B2(keyinput154), 
        .ZN(n3570) );
  OAI221_X1 U4391 ( .B1(n4898), .B2(keyinput158), .C1(n4899), .C2(keyinput154), 
        .A(n3570), .ZN(n3573) );
  INV_X1 U4392 ( .A(D_REG_4__SCAN_IN), .ZN(n4901) );
  AOI22_X1 U4393 ( .A1(n3079), .A2(keyinput162), .B1(keyinput143), .B2(n4901), 
        .ZN(n3571) );
  OAI221_X1 U4394 ( .B1(n3079), .B2(keyinput162), .C1(n4901), .C2(keyinput143), 
        .A(n3571), .ZN(n3572) );
  OR4_X1 U4395 ( .A1(n3575), .A2(n3574), .A3(n3573), .A4(n3572), .ZN(n3654) );
  INV_X1 U4396 ( .A(REG0_REG_27__SCAN_IN), .ZN(n3577) );
  INV_X1 U4397 ( .A(REG0_REG_29__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4398 ( .A1(n3577), .A2(keyinput147), .B1(n3809), .B2(keyinput133), 
        .ZN(n3576) );
  OAI221_X1 U4399 ( .B1(n3577), .B2(keyinput147), .C1(n3809), .C2(keyinput133), 
        .A(n3576), .ZN(n3584) );
  AOI22_X1 U4400 ( .A1(n2483), .A2(keyinput176), .B1(n3125), .B2(keyinput179), 
        .ZN(n3578) );
  OAI221_X1 U4401 ( .B1(n2483), .B2(keyinput176), .C1(n3125), .C2(keyinput179), 
        .A(n3578), .ZN(n3583) );
  AOI22_X1 U4402 ( .A1(n2604), .A2(keyinput231), .B1(n2642), .B2(keyinput189), 
        .ZN(n3579) );
  OAI221_X1 U4403 ( .B1(n2604), .B2(keyinput231), .C1(n2642), .C2(keyinput189), 
        .A(n3579), .ZN(n3582) );
  AOI22_X1 U4404 ( .A1(n4597), .A2(keyinput243), .B1(n4589), .B2(keyinput150), 
        .ZN(n3580) );
  OAI221_X1 U4405 ( .B1(n4597), .B2(keyinput243), .C1(n4589), .C2(keyinput150), 
        .A(n3580), .ZN(n3581) );
  NOR4_X1 U4406 ( .A1(n3584), .A2(n3583), .A3(n3582), .A4(n3581), .ZN(n3615)
         );
  AOI22_X1 U4407 ( .A1(n4585), .A2(keyinput224), .B1(n4571), .B2(keyinput211), 
        .ZN(n3585) );
  OAI221_X1 U4408 ( .B1(n4585), .B2(keyinput224), .C1(n4571), .C2(keyinput211), 
        .A(n3585), .ZN(n3593) );
  AOI22_X1 U4409 ( .A1(n3587), .A2(keyinput148), .B1(n3835), .B2(keyinput192), 
        .ZN(n3586) );
  OAI221_X1 U4410 ( .B1(n3587), .B2(keyinput148), .C1(n3835), .C2(keyinput192), 
        .A(n3586), .ZN(n3592) );
  AOI22_X1 U4411 ( .A1(n3100), .A2(keyinput197), .B1(n3099), .B2(keyinput152), 
        .ZN(n3588) );
  OAI221_X1 U4412 ( .B1(n3100), .B2(keyinput197), .C1(n3099), .C2(keyinput152), 
        .A(n3588), .ZN(n3591) );
  INV_X1 U4413 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4806) );
  AOI22_X1 U4414 ( .A1(n4806), .A2(keyinput214), .B1(n4688), .B2(keyinput129), 
        .ZN(n3589) );
  OAI221_X1 U4415 ( .B1(n4806), .B2(keyinput214), .C1(n4688), .C2(keyinput129), 
        .A(n3589), .ZN(n3590) );
  NOR4_X1 U4416 ( .A1(n3593), .A2(n3592), .A3(n3591), .A4(n3590), .ZN(n3614)
         );
  INV_X1 U4417 ( .A(ADDR_REG_17__SCAN_IN), .ZN(n3681) );
  INV_X1 U4418 ( .A(ADDR_REG_18__SCAN_IN), .ZN(n4854) );
  AOI22_X1 U4419 ( .A1(n3681), .A2(keyinput200), .B1(keyinput166), .B2(n4854), 
        .ZN(n3594) );
  OAI221_X1 U4420 ( .B1(n3681), .B2(keyinput200), .C1(n4854), .C2(keyinput166), 
        .A(n3594), .ZN(n3601) );
  INV_X1 U4421 ( .A(ADDR_REG_9__SCAN_IN), .ZN(n3678) );
  INV_X1 U4422 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n3682) );
  AOI22_X1 U4423 ( .A1(n3678), .A2(keyinput170), .B1(keyinput228), .B2(n3682), 
        .ZN(n3595) );
  OAI221_X1 U4424 ( .B1(n3678), .B2(keyinput170), .C1(n3682), .C2(keyinput228), 
        .A(n3595), .ZN(n3600) );
  INV_X1 U4425 ( .A(ADDR_REG_6__SCAN_IN), .ZN(n4743) );
  AOI22_X1 U4426 ( .A1(n4743), .A2(keyinput216), .B1(keyinput132), .B2(n3811), 
        .ZN(n3596) );
  OAI221_X1 U4427 ( .B1(n4743), .B2(keyinput216), .C1(n3811), .C2(keyinput132), 
        .A(n3596), .ZN(n3599) );
  INV_X1 U4428 ( .A(ADDR_REG_1__SCAN_IN), .ZN(n4136) );
  INV_X1 U4429 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n4742) );
  AOI22_X1 U4430 ( .A1(n4136), .A2(keyinput219), .B1(keyinput193), .B2(n4742), 
        .ZN(n3597) );
  OAI221_X1 U4431 ( .B1(n4136), .B2(keyinput219), .C1(n4742), .C2(keyinput193), 
        .A(n3597), .ZN(n3598) );
  NOR4_X1 U4432 ( .A1(n3601), .A2(n3600), .A3(n3599), .A4(n3598), .ZN(n3613)
         );
  AOI22_X1 U4433 ( .A1(n3603), .A2(keyinput172), .B1(keyinput165), .B2(n3793), 
        .ZN(n3602) );
  OAI221_X1 U4434 ( .B1(n3603), .B2(keyinput172), .C1(n3793), .C2(keyinput165), 
        .A(n3602), .ZN(n3611) );
  AOI22_X1 U4435 ( .A1(n3783), .A2(keyinput190), .B1(keyinput236), .B2(n3692), 
        .ZN(n3604) );
  OAI221_X1 U4436 ( .B1(n3783), .B2(keyinput190), .C1(n3692), .C2(keyinput236), 
        .A(n3604), .ZN(n3610) );
  AOI22_X1 U4437 ( .A1(n3834), .A2(keyinput185), .B1(keyinput245), .B2(n3606), 
        .ZN(n3605) );
  OAI221_X1 U4438 ( .B1(n3834), .B2(keyinput185), .C1(n3606), .C2(keyinput245), 
        .A(n3605), .ZN(n3609) );
  AOI22_X1 U4439 ( .A1(n3691), .A2(keyinput240), .B1(keyinput138), .B2(n3695), 
        .ZN(n3607) );
  OAI221_X1 U4440 ( .B1(n3691), .B2(keyinput240), .C1(n3695), .C2(keyinput138), 
        .A(n3607), .ZN(n3608) );
  NOR4_X1 U4441 ( .A1(n3611), .A2(n3610), .A3(n3609), .A4(n3608), .ZN(n3612)
         );
  NAND4_X1 U4442 ( .A1(n3615), .A2(n3614), .A3(n3613), .A4(n3612), .ZN(n3653)
         );
  AOI22_X1 U4443 ( .A1(DATAI_30_), .A2(keyinput196), .B1(DATAI_21_), .B2(
        keyinput235), .ZN(n3616) );
  OAI221_X1 U4444 ( .B1(DATAI_30_), .B2(keyinput196), .C1(DATAI_21_), .C2(
        keyinput235), .A(n3616), .ZN(n3623) );
  AOI22_X1 U4445 ( .A1(DATAI_10_), .A2(keyinput206), .B1(DATAI_16_), .B2(
        keyinput177), .ZN(n3617) );
  OAI221_X1 U4446 ( .B1(DATAI_10_), .B2(keyinput206), .C1(DATAI_16_), .C2(
        keyinput177), .A(n3617), .ZN(n3622) );
  AOI22_X1 U4447 ( .A1(DATAI_6_), .A2(keyinput251), .B1(REG3_REG_5__SCAN_IN), 
        .B2(keyinput238), .ZN(n3618) );
  OAI221_X1 U4448 ( .B1(DATAI_6_), .B2(keyinput251), .C1(REG3_REG_5__SCAN_IN), 
        .C2(keyinput238), .A(n3618), .ZN(n3621) );
  AOI22_X1 U4449 ( .A1(REG3_REG_20__SCAN_IN), .A2(keyinput255), .B1(
        IR_REG_1__SCAN_IN), .B2(keyinput183), .ZN(n3619) );
  OAI221_X1 U4450 ( .B1(REG3_REG_20__SCAN_IN), .B2(keyinput255), .C1(
        IR_REG_1__SCAN_IN), .C2(keyinput183), .A(n3619), .ZN(n3620) );
  NOR4_X1 U4451 ( .A1(n3623), .A2(n3622), .A3(n3621), .A4(n3620), .ZN(n3651)
         );
  AOI22_X1 U4452 ( .A1(IR_REG_4__SCAN_IN), .A2(keyinput198), .B1(
        IR_REG_3__SCAN_IN), .B2(keyinput136), .ZN(n3624) );
  OAI221_X1 U4453 ( .B1(IR_REG_4__SCAN_IN), .B2(keyinput198), .C1(
        IR_REG_3__SCAN_IN), .C2(keyinput136), .A(n3624), .ZN(n3631) );
  AOI22_X1 U4454 ( .A1(IR_REG_8__SCAN_IN), .A2(keyinput159), .B1(
        IR_REG_6__SCAN_IN), .B2(keyinput182), .ZN(n3625) );
  OAI221_X1 U4455 ( .B1(IR_REG_8__SCAN_IN), .B2(keyinput159), .C1(
        IR_REG_6__SCAN_IN), .C2(keyinput182), .A(n3625), .ZN(n3630) );
  AOI22_X1 U4456 ( .A1(IR_REG_25__SCAN_IN), .A2(keyinput203), .B1(
        IR_REG_24__SCAN_IN), .B2(keyinput248), .ZN(n3626) );
  OAI221_X1 U4457 ( .B1(IR_REG_25__SCAN_IN), .B2(keyinput203), .C1(
        IR_REG_24__SCAN_IN), .C2(keyinput248), .A(n3626), .ZN(n3629) );
  AOI22_X1 U4458 ( .A1(IR_REG_26__SCAN_IN), .A2(keyinput213), .B1(
        IR_REG_31__SCAN_IN), .B2(keyinput244), .ZN(n3627) );
  OAI221_X1 U4459 ( .B1(IR_REG_26__SCAN_IN), .B2(keyinput213), .C1(
        IR_REG_31__SCAN_IN), .C2(keyinput244), .A(n3627), .ZN(n3628) );
  NOR4_X1 U4460 ( .A1(n3631), .A2(n3630), .A3(n3629), .A4(n3628), .ZN(n3650)
         );
  AOI22_X1 U4461 ( .A1(D_REG_17__SCAN_IN), .A2(keyinput199), .B1(
        D_REG_6__SCAN_IN), .B2(keyinput181), .ZN(n3632) );
  OAI221_X1 U4462 ( .B1(D_REG_17__SCAN_IN), .B2(keyinput199), .C1(
        D_REG_6__SCAN_IN), .C2(keyinput181), .A(n3632), .ZN(n3639) );
  AOI22_X1 U4463 ( .A1(D_REG_24__SCAN_IN), .A2(keyinput188), .B1(
        D_REG_22__SCAN_IN), .B2(keyinput175), .ZN(n3633) );
  OAI221_X1 U4464 ( .B1(D_REG_24__SCAN_IN), .B2(keyinput188), .C1(
        D_REG_22__SCAN_IN), .C2(keyinput175), .A(n3633), .ZN(n3638) );
  AOI22_X1 U4465 ( .A1(D_REG_26__SCAN_IN), .A2(keyinput225), .B1(
        D_REG_28__SCAN_IN), .B2(keyinput221), .ZN(n3634) );
  OAI221_X1 U4466 ( .B1(D_REG_26__SCAN_IN), .B2(keyinput225), .C1(
        D_REG_28__SCAN_IN), .C2(keyinput221), .A(n3634), .ZN(n3637) );
  AOI22_X1 U4467 ( .A1(REG0_REG_15__SCAN_IN), .A2(keyinput151), .B1(
        REG0_REG_0__SCAN_IN), .B2(keyinput186), .ZN(n3635) );
  OAI221_X1 U4468 ( .B1(REG0_REG_15__SCAN_IN), .B2(keyinput151), .C1(
        REG0_REG_0__SCAN_IN), .C2(keyinput186), .A(n3635), .ZN(n3636) );
  NOR4_X1 U4469 ( .A1(n3639), .A2(n3638), .A3(n3637), .A4(n3636), .ZN(n3649)
         );
  AOI22_X1 U4470 ( .A1(REG0_REG_16__SCAN_IN), .A2(keyinput254), .B1(
        REG0_REG_19__SCAN_IN), .B2(keyinput226), .ZN(n3640) );
  OAI221_X1 U4471 ( .B1(REG0_REG_16__SCAN_IN), .B2(keyinput254), .C1(
        REG0_REG_19__SCAN_IN), .C2(keyinput226), .A(n3640), .ZN(n3647) );
  AOI22_X1 U4472 ( .A1(REG1_REG_0__SCAN_IN), .A2(keyinput164), .B1(
        REG0_REG_25__SCAN_IN), .B2(keyinput252), .ZN(n3641) );
  OAI221_X1 U4473 ( .B1(REG1_REG_0__SCAN_IN), .B2(keyinput164), .C1(
        REG0_REG_25__SCAN_IN), .C2(keyinput252), .A(n3641), .ZN(n3646) );
  AOI22_X1 U4474 ( .A1(REG0_REG_30__SCAN_IN), .A2(keyinput247), .B1(
        REG1_REG_2__SCAN_IN), .B2(keyinput161), .ZN(n3642) );
  OAI221_X1 U4475 ( .B1(REG0_REG_30__SCAN_IN), .B2(keyinput247), .C1(
        REG1_REG_2__SCAN_IN), .C2(keyinput161), .A(n3642), .ZN(n3645) );
  AOI22_X1 U4476 ( .A1(REG1_REG_5__SCAN_IN), .A2(keyinput242), .B1(
        REG1_REG_9__SCAN_IN), .B2(keyinput233), .ZN(n3643) );
  OAI221_X1 U4477 ( .B1(REG1_REG_5__SCAN_IN), .B2(keyinput242), .C1(
        REG1_REG_9__SCAN_IN), .C2(keyinput233), .A(n3643), .ZN(n3644) );
  NOR4_X1 U4478 ( .A1(n3647), .A2(n3646), .A3(n3645), .A4(n3644), .ZN(n3648)
         );
  NAND4_X1 U4479 ( .A1(n3651), .A2(n3650), .A3(n3649), .A4(n3648), .ZN(n3652)
         );
  NOR3_X1 U4480 ( .A1(n3654), .A2(n3653), .A3(n3652), .ZN(n3676) );
  INV_X1 U4481 ( .A(D_REG_23__SCAN_IN), .ZN(n4893) );
  AOI22_X1 U4482 ( .A1(n4896), .A2(keyinput145), .B1(keyinput156), .B2(n4893), 
        .ZN(n3655) );
  OAI221_X1 U4483 ( .B1(n4896), .B2(keyinput145), .C1(n4893), .C2(keyinput156), 
        .A(n3655), .ZN(n3662) );
  INV_X1 U4484 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4934) );
  AOI22_X1 U4485 ( .A1(n4891), .A2(keyinput173), .B1(keyinput128), .B2(n4934), 
        .ZN(n3656) );
  OAI221_X1 U4486 ( .B1(n4891), .B2(keyinput173), .C1(n4934), .C2(keyinput128), 
        .A(n3656), .ZN(n3661) );
  INV_X1 U4487 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4969) );
  INV_X1 U4488 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4951) );
  AOI22_X1 U4489 ( .A1(n4969), .A2(keyinput205), .B1(keyinput222), .B2(n4951), 
        .ZN(n3657) );
  OAI221_X1 U4490 ( .B1(n4969), .B2(keyinput205), .C1(n4951), .C2(keyinput222), 
        .A(n3657), .ZN(n3660) );
  INV_X1 U4491 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4977) );
  INV_X1 U4492 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4625) );
  AOI22_X1 U4493 ( .A1(n4977), .A2(keyinput253), .B1(n4625), .B2(keyinput178), 
        .ZN(n3658) );
  OAI221_X1 U4494 ( .B1(n4977), .B2(keyinput253), .C1(n4625), .C2(keyinput178), 
        .A(n3658), .ZN(n3659) );
  NOR4_X1 U4495 ( .A1(n3662), .A2(n3661), .A3(n3660), .A4(n3659), .ZN(n3675)
         );
  INV_X1 U4496 ( .A(DATAI_14_), .ZN(n4912) );
  AOI22_X1 U4497 ( .A1(IR_REG_30__SCAN_IN), .A2(keyinput191), .B1(n4912), .B2(
        keyinput215), .ZN(n3663) );
  OAI221_X1 U4498 ( .B1(IR_REG_30__SCAN_IN), .B2(keyinput191), .C1(n4912), 
        .C2(keyinput215), .A(n3663), .ZN(n3673) );
  INV_X1 U4499 ( .A(DATAI_13_), .ZN(n4913) );
  INV_X1 U4500 ( .A(DATAI_8_), .ZN(n4919) );
  AOI22_X1 U4501 ( .A1(n4913), .A2(keyinput157), .B1(n4919), .B2(keyinput202), 
        .ZN(n3664) );
  OAI221_X1 U4502 ( .B1(n4913), .B2(keyinput157), .C1(n4919), .C2(keyinput202), 
        .A(n3664), .ZN(n3672) );
  INV_X1 U4503 ( .A(DATAI_4_), .ZN(n3667) );
  INV_X1 U4504 ( .A(DATAI_5_), .ZN(n3666) );
  AOI22_X1 U4505 ( .A1(n3667), .A2(keyinput212), .B1(n3666), .B2(keyinput134), 
        .ZN(n3665) );
  OAI221_X1 U4506 ( .B1(n3667), .B2(keyinput212), .C1(n3666), .C2(keyinput134), 
        .A(n3665), .ZN(n3671) );
  INV_X1 U4507 ( .A(DATAI_3_), .ZN(n3669) );
  AOI22_X1 U4508 ( .A1(n3669), .A2(keyinput246), .B1(n3863), .B2(keyinput210), 
        .ZN(n3668) );
  OAI221_X1 U4509 ( .B1(n3669), .B2(keyinput246), .C1(n3863), .C2(keyinput210), 
        .A(n3668), .ZN(n3670) );
  NOR4_X1 U4510 ( .A1(n3673), .A2(n3672), .A3(n3671), .A4(n3670), .ZN(n3674)
         );
  NAND3_X1 U4511 ( .A1(n3676), .A2(n3675), .A3(n3674), .ZN(n3711) );
  INV_X1 U4512 ( .A(ADDR_REG_8__SCAN_IN), .ZN(n3679) );
  AOI22_X1 U4513 ( .A1(n3679), .A2(keyinput27), .B1(keyinput42), .B2(n3678), 
        .ZN(n3677) );
  OAI221_X1 U4514 ( .B1(n3679), .B2(keyinput27), .C1(n3678), .C2(keyinput42), 
        .A(n3677), .ZN(n3688) );
  AOI22_X1 U4515 ( .A1(n3682), .A2(keyinput100), .B1(n3681), .B2(keyinput72), 
        .ZN(n3680) );
  OAI221_X1 U4516 ( .B1(n3682), .B2(keyinput100), .C1(n3681), .C2(keyinput72), 
        .A(n3680), .ZN(n3687) );
  AOI22_X1 U4517 ( .A1(n3100), .A2(keyinput69), .B1(keyinput80), .B2(n3388), 
        .ZN(n3683) );
  OAI221_X1 U4518 ( .B1(n3100), .B2(keyinput69), .C1(n3388), .C2(keyinput80), 
        .A(n3683), .ZN(n3686) );
  AOI22_X1 U4519 ( .A1(n4597), .A2(keyinput115), .B1(keyinput86), .B2(n4806), 
        .ZN(n3684) );
  OAI221_X1 U4520 ( .B1(n4597), .B2(keyinput115), .C1(n4806), .C2(keyinput86), 
        .A(n3684), .ZN(n3685) );
  NOR4_X1 U4521 ( .A1(n3688), .A2(n3687), .A3(n3686), .A4(n3685), .ZN(n3710)
         );
  INV_X1 U4522 ( .A(DATAI_6_), .ZN(n4923) );
  AOI22_X1 U4523 ( .A1(n4580), .A2(keyinput122), .B1(keyinput123), .B2(n4923), 
        .ZN(n3689) );
  OAI221_X1 U4524 ( .B1(n4580), .B2(keyinput122), .C1(n4923), .C2(keyinput123), 
        .A(n3689), .ZN(n3699) );
  AOI22_X1 U4525 ( .A1(n3692), .A2(keyinput108), .B1(n3691), .B2(keyinput112), 
        .ZN(n3690) );
  OAI221_X1 U4526 ( .B1(n3692), .B2(keyinput108), .C1(n3691), .C2(keyinput112), 
        .A(n3690), .ZN(n3698) );
  INV_X1 U4527 ( .A(REG3_REG_17__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4528 ( .A1(n4899), .A2(keyinput26), .B1(keyinput39), .B2(n3909), 
        .ZN(n3693) );
  OAI221_X1 U4529 ( .B1(n4899), .B2(keyinput26), .C1(n3909), .C2(keyinput39), 
        .A(n3693), .ZN(n3697) );
  AOI22_X1 U4530 ( .A1(n3079), .A2(keyinput34), .B1(keyinput10), .B2(n3695), 
        .ZN(n3694) );
  OAI221_X1 U4531 ( .B1(n3079), .B2(keyinput34), .C1(n3695), .C2(keyinput10), 
        .A(n3694), .ZN(n3696) );
  NOR4_X1 U4532 ( .A1(n3699), .A2(n3698), .A3(n3697), .A4(n3696), .ZN(n3709)
         );
  AOI22_X1 U4533 ( .A1(DATAO_REG_0__SCAN_IN), .A2(keyinput3), .B1(
        REG2_REG_17__SCAN_IN), .B2(keyinput1), .ZN(n3700) );
  OAI221_X1 U4534 ( .B1(DATAO_REG_0__SCAN_IN), .B2(keyinput3), .C1(
        REG2_REG_17__SCAN_IN), .C2(keyinput1), .A(n3700), .ZN(n3707) );
  AOI22_X1 U4535 ( .A1(DATAO_REG_12__SCAN_IN), .A2(keyinput16), .B1(
        REG3_REG_20__SCAN_IN), .B2(keyinput127), .ZN(n3701) );
  OAI221_X1 U4536 ( .B1(DATAO_REG_12__SCAN_IN), .B2(keyinput16), .C1(
        REG3_REG_20__SCAN_IN), .C2(keyinput127), .A(n3701), .ZN(n3706) );
  AOI22_X1 U4537 ( .A1(REG0_REG_19__SCAN_IN), .A2(keyinput98), .B1(
        REG1_REG_25__SCAN_IN), .B2(keyinput41), .ZN(n3702) );
  OAI221_X1 U4538 ( .B1(REG0_REG_19__SCAN_IN), .B2(keyinput98), .C1(
        REG1_REG_25__SCAN_IN), .C2(keyinput41), .A(n3702), .ZN(n3705) );
  AOI22_X1 U4539 ( .A1(REG2_REG_24__SCAN_IN), .A2(keyinput43), .B1(
        REG2_REG_22__SCAN_IN), .B2(keyinput113), .ZN(n3703) );
  OAI221_X1 U4540 ( .B1(REG2_REG_24__SCAN_IN), .B2(keyinput43), .C1(
        REG2_REG_22__SCAN_IN), .C2(keyinput113), .A(n3703), .ZN(n3704) );
  NOR4_X1 U4541 ( .A1(n3707), .A2(n3706), .A3(n3705), .A4(n3704), .ZN(n3708)
         );
  NAND4_X1 U4542 ( .A1(n3711), .A2(n3710), .A3(n3709), .A4(n3708), .ZN(n3856)
         );
  OAI22_X1 U4543 ( .A1(IR_REG_31__SCAN_IN), .A2(keyinput116), .B1(DATAI_10_), 
        .B2(keyinput78), .ZN(n3712) );
  AOI221_X1 U4544 ( .B1(IR_REG_31__SCAN_IN), .B2(keyinput116), .C1(keyinput78), 
        .C2(DATAI_10_), .A(n3712), .ZN(n3719) );
  OAI22_X1 U4545 ( .A1(D_REG_8__SCAN_IN), .A2(keyinput21), .B1(
        IR_REG_30__SCAN_IN), .B2(keyinput63), .ZN(n3713) );
  AOI221_X1 U4546 ( .B1(D_REG_8__SCAN_IN), .B2(keyinput21), .C1(keyinput63), 
        .C2(IR_REG_30__SCAN_IN), .A(n3713), .ZN(n3718) );
  OAI22_X1 U4547 ( .A1(REG0_REG_27__SCAN_IN), .A2(keyinput19), .B1(keyinput20), 
        .B2(REG1_REG_27__SCAN_IN), .ZN(n3714) );
  AOI221_X1 U4548 ( .B1(REG0_REG_27__SCAN_IN), .B2(keyinput19), .C1(
        REG1_REG_27__SCAN_IN), .C2(keyinput20), .A(n3714), .ZN(n3717) );
  OAI22_X1 U4549 ( .A1(REG0_REG_0__SCAN_IN), .A2(keyinput58), .B1(
        DATAO_REG_24__SCAN_IN), .B2(keyinput40), .ZN(n3715) );
  AOI221_X1 U4550 ( .B1(REG0_REG_0__SCAN_IN), .B2(keyinput58), .C1(keyinput40), 
        .C2(DATAO_REG_24__SCAN_IN), .A(n3715), .ZN(n3716) );
  NAND4_X1 U4551 ( .A1(n3719), .A2(n3718), .A3(n3717), .A4(n3716), .ZN(n3767)
         );
  OAI22_X1 U4552 ( .A1(REG1_REG_13__SCAN_IN), .A2(keyinput67), .B1(keyinput12), 
        .B2(REG1_REG_15__SCAN_IN), .ZN(n3720) );
  AOI221_X1 U4553 ( .B1(REG1_REG_13__SCAN_IN), .B2(keyinput67), .C1(
        REG1_REG_15__SCAN_IN), .C2(keyinput12), .A(n3720), .ZN(n3727) );
  OAI22_X1 U4554 ( .A1(IR_REG_27__SCAN_IN), .A2(keyinput101), .B1(
        REG1_REG_16__SCAN_IN), .B2(keyinput52), .ZN(n3721) );
  AOI221_X1 U4555 ( .B1(IR_REG_27__SCAN_IN), .B2(keyinput101), .C1(keyinput52), 
        .C2(REG1_REG_16__SCAN_IN), .A(n3721), .ZN(n3726) );
  OAI22_X1 U4556 ( .A1(D_REG_17__SCAN_IN), .A2(keyinput71), .B1(keyinput114), 
        .B2(REG1_REG_5__SCAN_IN), .ZN(n3722) );
  AOI221_X1 U4557 ( .B1(D_REG_17__SCAN_IN), .B2(keyinput71), .C1(
        REG1_REG_5__SCAN_IN), .C2(keyinput114), .A(n3722), .ZN(n3725) );
  OAI22_X1 U4558 ( .A1(REG1_REG_9__SCAN_IN), .A2(keyinput105), .B1(
        REG1_REG_2__SCAN_IN), .B2(keyinput33), .ZN(n3723) );
  AOI221_X1 U4559 ( .B1(REG1_REG_9__SCAN_IN), .B2(keyinput105), .C1(keyinput33), .C2(REG1_REG_2__SCAN_IN), .A(n3723), .ZN(n3724) );
  NAND4_X1 U4560 ( .A1(n3727), .A2(n3726), .A3(n3725), .A4(n3724), .ZN(n3766)
         );
  AOI22_X1 U4561 ( .A1(DATAI_4_), .A2(keyinput84), .B1(D_REG_18__SCAN_IN), 
        .B2(keyinput76), .ZN(n3728) );
  OAI221_X1 U4562 ( .B1(DATAI_4_), .B2(keyinput84), .C1(D_REG_18__SCAN_IN), 
        .C2(keyinput76), .A(n3728), .ZN(n3735) );
  AOI22_X1 U4563 ( .A1(ADDR_REG_6__SCAN_IN), .A2(keyinput88), .B1(
        IR_REG_11__SCAN_IN), .B2(keyinput92), .ZN(n3729) );
  OAI221_X1 U4564 ( .B1(ADDR_REG_6__SCAN_IN), .B2(keyinput88), .C1(
        IR_REG_11__SCAN_IN), .C2(keyinput92), .A(n3729), .ZN(n3734) );
  AOI22_X1 U4565 ( .A1(REG0_REG_4__SCAN_IN), .A2(keyinput94), .B1(
        IR_REG_3__SCAN_IN), .B2(keyinput8), .ZN(n3730) );
  OAI221_X1 U4566 ( .B1(REG0_REG_4__SCAN_IN), .B2(keyinput94), .C1(
        IR_REG_3__SCAN_IN), .C2(keyinput8), .A(n3730), .ZN(n3733) );
  AOI22_X1 U4567 ( .A1(DATAO_REG_2__SCAN_IN), .A2(keyinput44), .B1(
        D_REG_23__SCAN_IN), .B2(keyinput28), .ZN(n3731) );
  OAI221_X1 U4568 ( .B1(DATAO_REG_2__SCAN_IN), .B2(keyinput44), .C1(
        D_REG_23__SCAN_IN), .C2(keyinput28), .A(n3731), .ZN(n3732) );
  NOR4_X1 U4569 ( .A1(n3735), .A2(n3734), .A3(n3733), .A4(n3732), .ZN(n3764)
         );
  AOI22_X1 U4570 ( .A1(REG0_REG_9__SCAN_IN), .A2(keyinput77), .B1(
        IR_REG_26__SCAN_IN), .B2(keyinput85), .ZN(n3736) );
  OAI221_X1 U4571 ( .B1(REG0_REG_9__SCAN_IN), .B2(keyinput77), .C1(
        IR_REG_26__SCAN_IN), .C2(keyinput85), .A(n3736), .ZN(n3743) );
  AOI22_X1 U4572 ( .A1(DATAO_REG_30__SCAN_IN), .A2(keyinput117), .B1(
        DATAO_REG_28__SCAN_IN), .B2(keyinput104), .ZN(n3737) );
  OAI221_X1 U4573 ( .B1(DATAO_REG_30__SCAN_IN), .B2(keyinput117), .C1(
        DATAO_REG_28__SCAN_IN), .C2(keyinput104), .A(n3737), .ZN(n3742) );
  AOI22_X1 U4574 ( .A1(REG1_REG_20__SCAN_IN), .A2(keyinput96), .B1(
        IR_REG_24__SCAN_IN), .B2(keyinput120), .ZN(n3738) );
  OAI221_X1 U4575 ( .B1(REG1_REG_20__SCAN_IN), .B2(keyinput96), .C1(
        IR_REG_24__SCAN_IN), .C2(keyinput120), .A(n3738), .ZN(n3741) );
  AOI22_X1 U4576 ( .A1(DATAI_13_), .A2(keyinput29), .B1(REG1_REG_12__SCAN_IN), 
        .B2(keyinput61), .ZN(n3739) );
  OAI221_X1 U4577 ( .B1(DATAI_13_), .B2(keyinput29), .C1(REG1_REG_12__SCAN_IN), 
        .C2(keyinput61), .A(n3739), .ZN(n3740) );
  NOR4_X1 U4578 ( .A1(n3743), .A2(n3742), .A3(n3741), .A4(n3740), .ZN(n3763)
         );
  INV_X1 U4579 ( .A(REG2_REG_25__SCAN_IN), .ZN(n3745) );
  AOI22_X1 U4580 ( .A1(REG0_REG_1__SCAN_IN), .A2(keyinput0), .B1(n3745), .B2(
        keyinput32), .ZN(n3744) );
  OAI221_X1 U4581 ( .B1(REG0_REG_1__SCAN_IN), .B2(keyinput0), .C1(n3745), .C2(
        keyinput32), .A(n3744), .ZN(n3752) );
  AOI22_X1 U4582 ( .A1(IR_REG_25__SCAN_IN), .A2(keyinput75), .B1(
        IR_REG_8__SCAN_IN), .B2(keyinput31), .ZN(n3746) );
  OAI221_X1 U4583 ( .B1(IR_REG_25__SCAN_IN), .B2(keyinput75), .C1(
        IR_REG_8__SCAN_IN), .C2(keyinput31), .A(n3746), .ZN(n3751) );
  INV_X1 U4584 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4687) );
  AOI22_X1 U4585 ( .A1(n4687), .A2(keyinput14), .B1(n2483), .B2(keyinput48), 
        .ZN(n3747) );
  OAI221_X1 U4586 ( .B1(n4687), .B2(keyinput14), .C1(n2483), .C2(keyinput48), 
        .A(n3747), .ZN(n3750) );
  AOI22_X1 U4587 ( .A1(n4589), .A2(keyinput22), .B1(keyinput102), .B2(n4683), 
        .ZN(n3748) );
  OAI221_X1 U4588 ( .B1(n4589), .B2(keyinput22), .C1(n4683), .C2(keyinput102), 
        .A(n3748), .ZN(n3749) );
  NOR4_X1 U4589 ( .A1(n3752), .A2(n3751), .A3(n3750), .A4(n3749), .ZN(n3762)
         );
  AOI22_X1 U4590 ( .A1(ADDR_REG_18__SCAN_IN), .A2(keyinput38), .B1(DATAI_5_), 
        .B2(keyinput6), .ZN(n3753) );
  OAI221_X1 U4591 ( .B1(ADDR_REG_18__SCAN_IN), .B2(keyinput38), .C1(DATAI_5_), 
        .C2(keyinput6), .A(n3753), .ZN(n3760) );
  AOI22_X1 U4592 ( .A1(DATAI_3_), .A2(keyinput118), .B1(D_REG_16__SCAN_IN), 
        .B2(keyinput30), .ZN(n3754) );
  OAI221_X1 U4593 ( .B1(DATAI_3_), .B2(keyinput118), .C1(D_REG_16__SCAN_IN), 
        .C2(keyinput30), .A(n3754), .ZN(n3759) );
  AOI22_X1 U4594 ( .A1(D_REG_4__SCAN_IN), .A2(keyinput15), .B1(
        D_REG_21__SCAN_IN), .B2(keyinput11), .ZN(n3755) );
  OAI221_X1 U4595 ( .B1(D_REG_4__SCAN_IN), .B2(keyinput15), .C1(
        D_REG_21__SCAN_IN), .C2(keyinput11), .A(n3755), .ZN(n3758) );
  AOI22_X1 U4596 ( .A1(IR_REG_6__SCAN_IN), .A2(keyinput54), .B1(
        IR_REG_18__SCAN_IN), .B2(keyinput2), .ZN(n3756) );
  OAI221_X1 U4597 ( .B1(IR_REG_6__SCAN_IN), .B2(keyinput54), .C1(
        IR_REG_18__SCAN_IN), .C2(keyinput2), .A(n3756), .ZN(n3757) );
  NOR4_X1 U4598 ( .A1(n3760), .A2(n3759), .A3(n3758), .A4(n3757), .ZN(n3761)
         );
  NAND4_X1 U4599 ( .A1(n3764), .A2(n3763), .A3(n3762), .A4(n3761), .ZN(n3765)
         );
  NOR3_X1 U4600 ( .A1(n3767), .A2(n3766), .A3(n3765), .ZN(n3854) );
  INV_X1 U4601 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4732) );
  AOI22_X1 U4602 ( .A1(n3917), .A2(keyinput13), .B1(keyinput99), .B2(n4732), 
        .ZN(n3768) );
  OAI221_X1 U4603 ( .B1(n3917), .B2(keyinput13), .C1(n4732), .C2(keyinput99), 
        .A(n3768), .ZN(n3777) );
  AOI22_X1 U4604 ( .A1(n3770), .A2(keyinput68), .B1(n4979), .B2(keyinput36), 
        .ZN(n3769) );
  OAI221_X1 U4605 ( .B1(n3770), .B2(keyinput68), .C1(n4979), .C2(keyinput36), 
        .A(n3769), .ZN(n3776) );
  INV_X1 U4606 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n4163) );
  AOI22_X1 U4607 ( .A1(n4163), .A2(keyinput7), .B1(n3125), .B2(keyinput51), 
        .ZN(n3771) );
  OAI221_X1 U4608 ( .B1(n4163), .B2(keyinput7), .C1(n3125), .C2(keyinput51), 
        .A(n3771), .ZN(n3775) );
  INV_X1 U4609 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4610 ( .A1(n3107), .A2(keyinput35), .B1(n3773), .B2(keyinput121), 
        .ZN(n3772) );
  OAI221_X1 U4611 ( .B1(n3107), .B2(keyinput35), .C1(n3773), .C2(keyinput121), 
        .A(n3772), .ZN(n3774) );
  NOR4_X1 U4612 ( .A1(n3777), .A2(n3776), .A3(n3775), .A4(n3774), .ZN(n3853)
         );
  INV_X1 U4613 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3779) );
  INV_X1 U4614 ( .A(ADDR_REG_14__SCAN_IN), .ZN(n4812) );
  AOI22_X1 U4615 ( .A1(n3779), .A2(keyinput23), .B1(keyinput18), .B2(n4812), 
        .ZN(n3778) );
  OAI221_X1 U4616 ( .B1(n3779), .B2(keyinput23), .C1(n4812), .C2(keyinput18), 
        .A(n3778), .ZN(n3788) );
  AOI22_X1 U4617 ( .A1(n4919), .A2(keyinput74), .B1(n3781), .B2(keyinput70), 
        .ZN(n3780) );
  OAI221_X1 U4618 ( .B1(n4919), .B2(keyinput74), .C1(n3781), .C2(keyinput70), 
        .A(n3780), .ZN(n3787) );
  AOI22_X1 U4619 ( .A1(n3783), .A2(keyinput62), .B1(n4912), .B2(keyinput87), 
        .ZN(n3782) );
  OAI221_X1 U4620 ( .B1(n3783), .B2(keyinput62), .C1(n4912), .C2(keyinput87), 
        .A(n3782), .ZN(n3786) );
  AOI22_X1 U4621 ( .A1(n3863), .A2(keyinput82), .B1(keyinput83), .B2(n4571), 
        .ZN(n3784) );
  OAI221_X1 U4622 ( .B1(n3863), .B2(keyinput82), .C1(n4571), .C2(keyinput83), 
        .A(n3784), .ZN(n3785) );
  NOR4_X1 U4623 ( .A1(n3788), .A2(n3787), .A3(n3786), .A4(n3785), .ZN(n3852)
         );
  INV_X1 U4624 ( .A(D_REG_28__SCAN_IN), .ZN(n4889) );
  AOI22_X1 U4625 ( .A1(n4889), .A2(keyinput93), .B1(keyinput73), .B2(n3790), 
        .ZN(n3789) );
  OAI221_X1 U4626 ( .B1(n4889), .B2(keyinput93), .C1(n3790), .C2(keyinput73), 
        .A(n3789), .ZN(n3798) );
  INV_X1 U4627 ( .A(DATAI_16_), .ZN(n4908) );
  AOI22_X1 U4628 ( .A1(n4742), .A2(keyinput65), .B1(n4908), .B2(keyinput49), 
        .ZN(n3791) );
  OAI221_X1 U4629 ( .B1(n4742), .B2(keyinput65), .C1(n4908), .C2(keyinput49), 
        .A(n3791), .ZN(n3797) );
  INV_X1 U4630 ( .A(D_REG_6__SCAN_IN), .ZN(n4900) );
  AOI22_X1 U4631 ( .A1(n4900), .A2(keyinput53), .B1(keyinput37), .B2(n3793), 
        .ZN(n3792) );
  OAI221_X1 U4632 ( .B1(n4900), .B2(keyinput53), .C1(n3793), .C2(keyinput37), 
        .A(n3792), .ZN(n3796) );
  AOI22_X1 U4633 ( .A1(n4891), .A2(keyinput45), .B1(n4896), .B2(keyinput17), 
        .ZN(n3794) );
  OAI221_X1 U4634 ( .B1(n4891), .B2(keyinput45), .C1(n4896), .C2(keyinput17), 
        .A(n3794), .ZN(n3795) );
  NOR4_X1 U4635 ( .A1(n3798), .A2(n3797), .A3(n3796), .A4(n3795), .ZN(n3850)
         );
  AOI22_X1 U4636 ( .A1(ADDR_REG_7__SCAN_IN), .A2(keyinput79), .B1(
        REG2_REG_8__SCAN_IN), .B2(keyinput89), .ZN(n3799) );
  OAI221_X1 U4637 ( .B1(ADDR_REG_7__SCAN_IN), .B2(keyinput79), .C1(
        REG2_REG_8__SCAN_IN), .C2(keyinput89), .A(n3799), .ZN(n3806) );
  AOI22_X1 U4638 ( .A1(REG3_REG_1__SCAN_IN), .A2(keyinput25), .B1(
        REG0_REG_16__SCAN_IN), .B2(keyinput126), .ZN(n3800) );
  OAI221_X1 U4639 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput25), .C1(
        REG0_REG_16__SCAN_IN), .C2(keyinput126), .A(n3800), .ZN(n3805) );
  AOI22_X1 U4640 ( .A1(REG2_REG_5__SCAN_IN), .A2(keyinput24), .B1(
        REG2_REG_7__SCAN_IN), .B2(keyinput46), .ZN(n3801) );
  OAI221_X1 U4641 ( .B1(REG2_REG_5__SCAN_IN), .B2(keyinput24), .C1(
        REG2_REG_7__SCAN_IN), .C2(keyinput46), .A(n3801), .ZN(n3804) );
  AOI22_X1 U4642 ( .A1(ADDR_REG_15__SCAN_IN), .A2(keyinput9), .B1(
        REG2_REG_15__SCAN_IN), .B2(keyinput66), .ZN(n3802) );
  OAI221_X1 U4643 ( .B1(ADDR_REG_15__SCAN_IN), .B2(keyinput9), .C1(
        REG2_REG_15__SCAN_IN), .C2(keyinput66), .A(n3802), .ZN(n3803) );
  NOR4_X1 U4644 ( .A1(n3806), .A2(n3805), .A3(n3804), .A4(n3803), .ZN(n3849)
         );
  INV_X1 U4645 ( .A(D_REG_22__SCAN_IN), .ZN(n4894) );
  AOI22_X1 U4646 ( .A1(n4894), .A2(keyinput47), .B1(keyinput59), .B2(n4803), 
        .ZN(n3807) );
  OAI221_X1 U4647 ( .B1(n4894), .B2(keyinput47), .C1(n4803), .C2(keyinput59), 
        .A(n3807), .ZN(n3814) );
  AOI22_X1 U4648 ( .A1(n3810), .A2(keyinput95), .B1(keyinput5), .B2(n3809), 
        .ZN(n3808) );
  OAI221_X1 U4649 ( .B1(n3810), .B2(keyinput95), .C1(n3809), .C2(keyinput5), 
        .A(n3808), .ZN(n3813) );
  XNOR2_X1 U4650 ( .A(n3811), .B(keyinput4), .ZN(n3812) );
  NOR3_X1 U4651 ( .A1(n3814), .A2(n3813), .A3(n3812), .ZN(n3832) );
  INV_X1 U4652 ( .A(D_REG_24__SCAN_IN), .ZN(n4892) );
  AOI22_X1 U4653 ( .A1(n4892), .A2(keyinput60), .B1(keyinput56), .B2(n3816), 
        .ZN(n3815) );
  OAI221_X1 U4654 ( .B1(n4892), .B2(keyinput60), .C1(n3816), .C2(keyinput56), 
        .A(n3815), .ZN(n3822) );
  INV_X1 U4655 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4629) );
  AOI22_X1 U4656 ( .A1(n4629), .A2(keyinput124), .B1(n4625), .B2(keyinput50), 
        .ZN(n3817) );
  OAI221_X1 U4657 ( .B1(n4629), .B2(keyinput124), .C1(n4625), .C2(keyinput50), 
        .A(n3817), .ZN(n3821) );
  XNOR2_X1 U4658 ( .A(IR_REG_17__SCAN_IN), .B(keyinput109), .ZN(n3819) );
  XNOR2_X1 U4659 ( .A(keyinput110), .B(REG3_REG_5__SCAN_IN), .ZN(n3818) );
  NAND2_X1 U4660 ( .A1(n3819), .A2(n3818), .ZN(n3820) );
  NOR3_X1 U4661 ( .A1(n3822), .A2(n3821), .A3(n3820), .ZN(n3831) );
  INV_X1 U4662 ( .A(D_REG_26__SCAN_IN), .ZN(n4890) );
  AOI22_X1 U4663 ( .A1(n4977), .A2(keyinput125), .B1(n4890), .B2(keyinput97), 
        .ZN(n3823) );
  OAI221_X1 U4664 ( .B1(n4977), .B2(keyinput125), .C1(n4890), .C2(keyinput97), 
        .A(n3823), .ZN(n3829) );
  XNOR2_X1 U4665 ( .A(IR_REG_19__SCAN_IN), .B(keyinput106), .ZN(n3827) );
  XNOR2_X1 U4666 ( .A(IR_REG_9__SCAN_IN), .B(keyinput90), .ZN(n3826) );
  XNOR2_X1 U4667 ( .A(IR_REG_5__SCAN_IN), .B(keyinput81), .ZN(n3825) );
  XNOR2_X1 U4668 ( .A(IR_REG_1__SCAN_IN), .B(keyinput55), .ZN(n3824) );
  NAND4_X1 U4669 ( .A1(n3827), .A2(n3826), .A3(n3825), .A4(n3824), .ZN(n3828)
         );
  NOR2_X1 U4670 ( .A1(n3829), .A2(n3828), .ZN(n3830) );
  NAND3_X1 U4671 ( .A1(n3832), .A2(n3831), .A3(n3830), .ZN(n3847) );
  AOI22_X1 U4672 ( .A1(n3835), .A2(keyinput64), .B1(keyinput57), .B2(n3834), 
        .ZN(n3833) );
  OAI221_X1 U4673 ( .B1(n3835), .B2(keyinput64), .C1(n3834), .C2(keyinput57), 
        .A(n3833), .ZN(n3839) );
  INV_X1 U4674 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4619) );
  AOI22_X1 U4675 ( .A1(n3837), .A2(keyinput107), .B1(keyinput119), .B2(n4619), 
        .ZN(n3836) );
  OAI221_X1 U4676 ( .B1(n3837), .B2(keyinput107), .C1(n4619), .C2(keyinput119), 
        .A(n3836), .ZN(n3838) );
  NOR2_X1 U4677 ( .A1(n3839), .A2(n3838), .ZN(n3845) );
  AOI22_X1 U4678 ( .A1(n4136), .A2(keyinput91), .B1(n2604), .B2(keyinput103), 
        .ZN(n3840) );
  OAI221_X1 U4679 ( .B1(n4136), .B2(keyinput91), .C1(n2604), .C2(keyinput103), 
        .A(n3840), .ZN(n3843) );
  XNOR2_X1 U4680 ( .A(n3841), .B(keyinput111), .ZN(n3842) );
  NOR2_X1 U4681 ( .A1(n3843), .A2(n3842), .ZN(n3844) );
  NAND2_X1 U4682 ( .A1(n3845), .A2(n3844), .ZN(n3846) );
  NOR2_X1 U4683 ( .A1(n3847), .A2(n3846), .ZN(n3848) );
  AND3_X1 U4684 ( .A1(n3850), .A2(n3849), .A3(n3848), .ZN(n3851) );
  NAND4_X1 U4685 ( .A1(n3854), .A2(n3853), .A3(n3852), .A4(n3851), .ZN(n3855)
         );
  NOR2_X1 U4686 ( .A1(n3856), .A2(n3855), .ZN(n3869) );
  OAI21_X1 U4687 ( .B1(n3949), .B2(n3860), .A(n3859), .ZN(n3861) );
  NAND3_X1 U4688 ( .A1(n3862), .A2(n3968), .A3(n3861), .ZN(n3867) );
  AOI22_X1 U4689 ( .A1(n4724), .A2(n4358), .B1(n3963), .B2(n4321), .ZN(n3866)
         );
  OAI22_X1 U4690 ( .A1(n3953), .A2(n2934), .B1(STATE_REG_SCAN_IN), .B2(n3863), 
        .ZN(n3864) );
  AOI21_X1 U4691 ( .B1(n4327), .B2(n3955), .A(n3864), .ZN(n3865) );
  NAND3_X1 U4692 ( .A1(n3867), .A2(n3866), .A3(n3865), .ZN(n3868) );
  XOR2_X1 U4693 ( .A(n3869), .B(n3868), .Z(U3213) );
  XOR2_X1 U4694 ( .A(n3871), .B(n3870), .Z(n3876) );
  AOI22_X1 U4695 ( .A1(n4724), .A2(n4402), .B1(n3963), .B2(n4126), .ZN(n3875)
         );
  NOR2_X1 U4696 ( .A1(n3872), .A2(STATE_REG_SCAN_IN), .ZN(n4693) );
  NOR2_X1 U4697 ( .A1(n3953), .A2(n4407), .ZN(n3873) );
  AOI211_X1 U4698 ( .C1(n4408), .C2(n3955), .A(n4693), .B(n3873), .ZN(n3874)
         );
  OAI211_X1 U4699 ( .C1(n3876), .C2(n4719), .A(n3875), .B(n3874), .ZN(U3216)
         );
  XNOR2_X1 U4700 ( .A(n3879), .B(n3878), .ZN(n3880) );
  XNOR2_X1 U4701 ( .A(n3881), .B(n3880), .ZN(n3886) );
  AOI22_X1 U4702 ( .A1(n4724), .A2(n4126), .B1(n3963), .B2(n4358), .ZN(n3885)
         );
  INV_X1 U4703 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3882) );
  OAI22_X1 U4704 ( .A1(n3953), .A2(n4362), .B1(STATE_REG_SCAN_IN), .B2(n3882), 
        .ZN(n3883) );
  AOI21_X1 U4705 ( .B1(n4364), .B2(n3955), .A(n3883), .ZN(n3884) );
  OAI211_X1 U4706 ( .C1(n3886), .C2(n4719), .A(n3885), .B(n3884), .ZN(U3220)
         );
  NOR2_X1 U4707 ( .A1(n3889), .A2(n2361), .ZN(n3890) );
  XNOR2_X1 U4708 ( .A(n3887), .B(n3890), .ZN(n3895) );
  AOI22_X1 U4709 ( .A1(n4724), .A2(n4321), .B1(n3963), .B2(n4285), .ZN(n3894)
         );
  OAI22_X1 U4710 ( .A1(n3953), .A2(n4289), .B1(STATE_REG_SCAN_IN), .B2(n3891), 
        .ZN(n3892) );
  AOI21_X1 U4711 ( .B1(n4291), .B2(n3955), .A(n3892), .ZN(n3893) );
  OAI211_X1 U4712 ( .C1(n3895), .C2(n4719), .A(n3894), .B(n3893), .ZN(U3222)
         );
  OAI21_X1 U4713 ( .B1(n3896), .B2(n3961), .A(n3959), .ZN(n3898) );
  XNOR2_X1 U4714 ( .A(n3898), .B(n3897), .ZN(n3904) );
  AOI22_X1 U4715 ( .A1(n4711), .A2(n4723), .B1(n4724), .B2(n4494), .ZN(n3903)
         );
  INV_X1 U4716 ( .A(REG3_REG_16__SCAN_IN), .ZN(n3899) );
  NOR2_X1 U4717 ( .A1(STATE_REG_SCAN_IN), .A2(n3899), .ZN(n4824) );
  NOR2_X1 U4718 ( .A1(n3953), .A2(n4453), .ZN(n3900) );
  AOI211_X1 U4719 ( .C1(n3901), .C2(n3955), .A(n4824), .B(n3900), .ZN(n3902)
         );
  OAI211_X1 U4720 ( .C1(n3904), .C2(n4719), .A(n3903), .B(n3902), .ZN(U3223)
         );
  XNOR2_X1 U4721 ( .A(n3906), .B(n3905), .ZN(n3907) );
  XNOR2_X1 U4722 ( .A(n3908), .B(n3907), .ZN(n3913) );
  AOI22_X1 U4723 ( .A1(n4724), .A2(n4439), .B1(n3963), .B2(n4402), .ZN(n3912)
         );
  NOR2_X1 U4724 ( .A1(STATE_REG_SCAN_IN), .A2(n3909), .ZN(n4185) );
  NOR2_X1 U4725 ( .A1(n3953), .A2(n4436), .ZN(n3910) );
  AOI211_X1 U4726 ( .C1(n4445), .C2(n3955), .A(n4185), .B(n3910), .ZN(n3911)
         );
  OAI211_X1 U4727 ( .C1(n3913), .C2(n4719), .A(n3912), .B(n3911), .ZN(U3225)
         );
  NAND2_X1 U4728 ( .A1(n2250), .A2(n3914), .ZN(n3916) );
  XNOR2_X1 U4729 ( .A(n3916), .B(n3915), .ZN(n3922) );
  AOI22_X1 U4730 ( .A1(n4724), .A2(n4125), .B1(n4711), .B2(n4302), .ZN(n3921)
         );
  INV_X1 U4731 ( .A(n4305), .ZN(n3919) );
  OAI22_X1 U4732 ( .A1(n3953), .A2(n4308), .B1(STATE_REG_SCAN_IN), .B2(n3917), 
        .ZN(n3918) );
  AOI21_X1 U4733 ( .B1(n3919), .B2(n3955), .A(n3918), .ZN(n3920) );
  OAI211_X1 U4734 ( .C1(n3922), .C2(n4719), .A(n3921), .B(n3920), .ZN(U3226)
         );
  INV_X1 U4735 ( .A(n3923), .ZN(n3928) );
  AOI21_X1 U4736 ( .B1(n3927), .B2(n3925), .A(n3924), .ZN(n3926) );
  AOI21_X1 U4737 ( .B1(n3928), .B2(n3927), .A(n3926), .ZN(n3934) );
  AOI22_X1 U4738 ( .A1(n4724), .A2(n4710), .B1(n3963), .B2(n4378), .ZN(n3933)
         );
  INV_X1 U4739 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3929) );
  OAI22_X1 U4740 ( .A1(n3953), .A2(n4385), .B1(STATE_REG_SCAN_IN), .B2(n3929), 
        .ZN(n3930) );
  AOI21_X1 U4741 ( .B1(n3931), .B2(n3955), .A(n3930), .ZN(n3932) );
  OAI211_X1 U4742 ( .C1(n3934), .C2(n4719), .A(n3933), .B(n3932), .ZN(U3230)
         );
  NAND2_X1 U4743 ( .A1(n3936), .A2(n3935), .ZN(n3943) );
  INV_X1 U4744 ( .A(n3460), .ZN(n3941) );
  OAI21_X1 U4745 ( .B1(n3460), .B2(n3938), .A(n3937), .ZN(n3939) );
  OAI21_X1 U4746 ( .B1(n3941), .B2(n3940), .A(n3939), .ZN(n3942) );
  XOR2_X1 U4747 ( .A(n3943), .B(n3942), .Z(n3948) );
  AOI22_X1 U4748 ( .A1(n4711), .A2(n4517), .B1(n4724), .B2(n4128), .ZN(n3947)
         );
  NOR2_X1 U4749 ( .A1(STATE_REG_SCAN_IN), .A2(n3944), .ZN(n4793) );
  NOR2_X1 U4750 ( .A1(n3953), .A2(n4525), .ZN(n3945) );
  AOI211_X1 U4751 ( .C1(n4527), .C2(n3955), .A(n4793), .B(n3945), .ZN(n3946)
         );
  OAI211_X1 U4752 ( .C1(n3948), .C2(n4719), .A(n3947), .B(n3946), .ZN(U3231)
         );
  AOI21_X1 U4753 ( .B1(n3951), .B2(n3950), .A(n3949), .ZN(n3958) );
  AOI22_X1 U4754 ( .A1(n4711), .A2(n4125), .B1(n4724), .B2(n4378), .ZN(n3957)
         );
  OAI22_X1 U4755 ( .A1(n3953), .A2(n4345), .B1(STATE_REG_SCAN_IN), .B2(n3952), 
        .ZN(n3954) );
  AOI21_X1 U4756 ( .B1(n4337), .B2(n3955), .A(n3954), .ZN(n3956) );
  OAI211_X1 U4757 ( .C1(n3958), .C2(n4719), .A(n3957), .B(n3956), .ZN(U3232)
         );
  INV_X1 U4758 ( .A(n3896), .ZN(n3960) );
  NAND2_X1 U4759 ( .A1(n3960), .A2(n3959), .ZN(n3962) );
  XNOR2_X1 U4760 ( .A(n3962), .B(n3961), .ZN(n3969) );
  AOI22_X1 U4761 ( .A1(n4724), .A2(n4517), .B1(n3963), .B2(n4439), .ZN(n3966)
         );
  NAND2_X1 U4762 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4821) );
  INV_X1 U4763 ( .A(n4821), .ZN(n3964) );
  AOI21_X1 U4764 ( .B1(n4712), .B2(n4474), .A(n3964), .ZN(n3965) );
  OAI211_X1 U4765 ( .C1(n4728), .C2(n4475), .A(n3966), .B(n3965), .ZN(n3967)
         );
  AOI21_X1 U4766 ( .B1(n3969), .B2(n3968), .A(n3967), .ZN(n3970) );
  INV_X1 U4767 ( .A(n3970), .ZN(U3238) );
  NAND2_X1 U4768 ( .A1(n4212), .A2(n3971), .ZN(n4010) );
  NAND2_X1 U4769 ( .A1(n4124), .A2(n4010), .ZN(n4002) );
  NAND2_X1 U4770 ( .A1(n3973), .A2(n3972), .ZN(n4066) );
  AND2_X1 U4771 ( .A1(n4066), .A2(n3975), .ZN(n4085) );
  INV_X1 U4772 ( .A(n4085), .ZN(n3977) );
  INV_X1 U4773 ( .A(n3974), .ZN(n4087) );
  AOI21_X1 U4774 ( .B1(n3976), .B2(n3975), .A(n4085), .ZN(n4082) );
  AOI211_X1 U4775 ( .C1(n4492), .C2(n3977), .A(n4087), .B(n4082), .ZN(n3980)
         );
  INV_X1 U4776 ( .A(n4027), .ZN(n4394) );
  INV_X1 U4777 ( .A(n3978), .ZN(n3979) );
  NOR4_X1 U4778 ( .A1(n3980), .A2(n2278), .A3(n4394), .A4(n3979), .ZN(n3982)
         );
  OAI21_X1 U4779 ( .B1(n3982), .B2(n3981), .A(n4093), .ZN(n3984) );
  AOI21_X1 U4780 ( .B1(n4097), .B2(n3984), .A(n3983), .ZN(n3988) );
  OR2_X1 U4781 ( .A1(n3991), .A2(n3990), .ZN(n4035) );
  NAND4_X1 U4782 ( .A1(n3986), .A2(n4035), .A3(n4207), .A4(n3985), .ZN(n3987)
         );
  AOI221_X1 U4783 ( .B1(n3988), .B2(n4260), .C1(n4099), .C2(n4260), .A(n3987), 
        .ZN(n3998) );
  INV_X1 U4784 ( .A(n4212), .ZN(n3989) );
  NOR2_X1 U4785 ( .A1(n4009), .A2(n4008), .ZN(n4107) );
  AOI21_X1 U4786 ( .B1(n4544), .B2(n3989), .A(n4107), .ZN(n4037) );
  NAND2_X1 U4787 ( .A1(n3991), .A2(n3990), .ZN(n4034) );
  NAND4_X1 U4788 ( .A1(n4237), .A2(n4034), .A3(n4206), .A4(n3992), .ZN(n3997)
         );
  NAND2_X1 U4789 ( .A1(n4034), .A2(n4206), .ZN(n4102) );
  INV_X1 U4790 ( .A(n4207), .ZN(n3994) );
  NOR2_X1 U4791 ( .A1(n3994), .A2(n3993), .ZN(n3995) );
  OAI211_X1 U4792 ( .C1(n4102), .C2(n3995), .A(n4035), .B(n4037), .ZN(n4108)
         );
  INV_X1 U4793 ( .A(n4108), .ZN(n3996) );
  AOI22_X1 U4794 ( .A1(n3998), .A2(n4037), .B1(n3997), .B2(n3996), .ZN(n3999)
         );
  AOI21_X1 U4795 ( .B1(n4009), .B2(n4544), .A(n3999), .ZN(n4000) );
  AOI211_X1 U4796 ( .C1(n4008), .C2(n4002), .A(n4001), .B(n4000), .ZN(n4115)
         );
  INV_X1 U4797 ( .A(n4003), .ZN(n4220) );
  XNOR2_X1 U4798 ( .A(n4126), .B(n4385), .ZN(n4376) );
  XNOR2_X1 U4799 ( .A(n4710), .B(n4407), .ZN(n4399) );
  NOR2_X1 U4800 ( .A1(n4376), .A2(n4399), .ZN(n4019) );
  NAND2_X1 U4801 ( .A1(n4004), .A2(n4279), .ZN(n4299) );
  INV_X1 U4802 ( .A(n4005), .ZN(n4007) );
  NAND2_X1 U4803 ( .A1(n4009), .A2(n4008), .ZN(n4011) );
  AND2_X1 U4804 ( .A1(n4011), .A2(n4010), .ZN(n4106) );
  INV_X1 U4805 ( .A(n4106), .ZN(n4012) );
  NOR4_X1 U4806 ( .A1(n4299), .A2(n4513), .A3(n4046), .A4(n4012), .ZN(n4018)
         );
  NAND2_X1 U4807 ( .A1(n4013), .A2(n4297), .ZN(n4318) );
  NOR4_X1 U4808 ( .A1(n4318), .A2(n4016), .A3(n4015), .A4(n4014), .ZN(n4017)
         );
  NAND4_X1 U4809 ( .A1(n4220), .A2(n4019), .A3(n4018), .A4(n4017), .ZN(n4041)
         );
  INV_X1 U4810 ( .A(n4422), .ZN(n4415) );
  NAND4_X1 U4811 ( .A1(n4415), .A2(n4021), .A3(n4856), .A4(n4020), .ZN(n4026)
         );
  NAND2_X1 U4812 ( .A1(n4491), .A2(n4022), .ZN(n4025) );
  NOR4_X1 U4813 ( .A1(n4026), .A2(n4025), .A3(n4024), .A4(n4023), .ZN(n4033)
         );
  INV_X1 U4814 ( .A(n4314), .ZN(n4094) );
  NAND2_X1 U4815 ( .A1(n4094), .A2(n4315), .ZN(n4354) );
  NAND2_X1 U4816 ( .A1(n4393), .A2(n4027), .ZN(n4435) );
  NOR4_X1 U4817 ( .A1(n4354), .A2(n4435), .A3(n4029), .A4(n4028), .ZN(n4032)
         );
  NOR4_X1 U4818 ( .A1(n4333), .A2(n4451), .A3(n4481), .A4(n4030), .ZN(n4031)
         );
  NAND4_X1 U4819 ( .A1(n4033), .A2(n4237), .A3(n4032), .A4(n4031), .ZN(n4040)
         );
  NAND2_X1 U4820 ( .A1(n4258), .A2(n4036), .ZN(n4282) );
  INV_X1 U4821 ( .A(n4282), .ZN(n4038) );
  NAND2_X1 U4822 ( .A1(n4875), .A2(n2234), .ZN(n4045) );
  NAND4_X1 U4823 ( .A1(n4222), .A2(n4038), .A3(n4037), .A4(n4882), .ZN(n4039)
         );
  XNOR2_X1 U4824 ( .A(n4285), .B(n4264), .ZN(n4261) );
  NOR4_X1 U4825 ( .A1(n4041), .A2(n4040), .A3(n4039), .A4(n4261), .ZN(n4113)
         );
  NOR2_X1 U4826 ( .A1(n4042), .A2(n4249), .ZN(n4105) );
  INV_X1 U4827 ( .A(n4043), .ZN(n4047) );
  OAI211_X1 U4828 ( .C1(n4047), .C2(n4046), .A(n4045), .B(n4044), .ZN(n4049)
         );
  NAND3_X1 U4829 ( .A1(n4049), .A2(n4048), .A3(n2959), .ZN(n4052) );
  NAND3_X1 U4830 ( .A1(n4052), .A2(n4051), .A3(n4050), .ZN(n4055) );
  NAND3_X1 U4831 ( .A1(n4055), .A2(n4054), .A3(n4053), .ZN(n4058) );
  NAND4_X1 U4832 ( .A1(n4058), .A2(n4057), .A3(n4056), .A4(n4068), .ZN(n4061)
         );
  NAND3_X1 U4833 ( .A1(n4061), .A2(n4060), .A3(n4059), .ZN(n4062) );
  NAND3_X1 U4834 ( .A1(n4062), .A2(n4067), .A3(n4069), .ZN(n4065) );
  NAND3_X1 U4835 ( .A1(n4065), .A2(n4064), .A3(n4063), .ZN(n4075) );
  INV_X1 U4836 ( .A(n4066), .ZN(n4074) );
  INV_X1 U4837 ( .A(n4067), .ZN(n4072) );
  NAND2_X1 U4838 ( .A1(n4069), .A2(n4068), .ZN(n4070) );
  NOR4_X1 U4839 ( .A1(n4085), .A2(n4072), .A3(n4071), .A4(n4070), .ZN(n4073)
         );
  AOI21_X1 U4840 ( .B1(n4075), .B2(n4074), .A(n4073), .ZN(n4078) );
  OAI22_X1 U4841 ( .A1(n4078), .A2(n4077), .B1(n4085), .B2(n4076), .ZN(n4081)
         );
  NAND3_X1 U4842 ( .A1(n4081), .A2(n4080), .A3(n4079), .ZN(n4084) );
  INV_X1 U4843 ( .A(n4082), .ZN(n4083) );
  OAI211_X1 U4844 ( .C1(n4086), .C2(n4085), .A(n4084), .B(n4083), .ZN(n4089)
         );
  AOI21_X1 U4845 ( .B1(n4089), .B2(n4088), .A(n4087), .ZN(n4092) );
  OAI21_X1 U4846 ( .B1(n4092), .B2(n4091), .A(n4090), .ZN(n4095) );
  NAND3_X1 U4847 ( .A1(n4095), .A2(n4094), .A3(n4093), .ZN(n4096) );
  NAND2_X1 U4848 ( .A1(n4097), .A2(n4096), .ZN(n4100) );
  AOI211_X1 U4849 ( .C1(n4101), .C2(n4100), .A(n4099), .B(n4098), .ZN(n4104)
         );
  NOR4_X1 U4850 ( .A1(n4105), .A2(n4104), .A3(n4103), .A4(n4102), .ZN(n4109)
         );
  OAI22_X1 U4851 ( .A1(n4109), .A2(n4108), .B1(n4107), .B2(n4106), .ZN(n4110)
         );
  INV_X1 U4852 ( .A(n4110), .ZN(n4112) );
  MUX2_X1 U4853 ( .A(n4113), .B(n4112), .S(n4111), .Z(n4114) );
  NOR2_X1 U4854 ( .A1(n4115), .A2(n4114), .ZN(n4116) );
  XNOR2_X1 U4855 ( .A(n4116), .B(n4695), .ZN(n4123) );
  NOR2_X1 U4856 ( .A1(n4904), .A2(n4117), .ZN(n4118) );
  NAND4_X1 U4857 ( .A1(n4119), .A2(n4737), .A3(n4118), .A4(n4673), .ZN(n4120)
         );
  OAI211_X1 U4858 ( .C1(n4675), .C2(n4122), .A(n4120), .B(B_REG_SCAN_IN), .ZN(
        n4121) );
  OAI21_X1 U4859 ( .B1(n4123), .B2(n4122), .A(n4121), .ZN(U3239) );
  MUX2_X1 U4860 ( .A(n4124), .B(DATAO_REG_31__SCAN_IN), .S(n4134), .Z(U3581)
         );
  MUX2_X1 U4861 ( .A(n4243), .B(DATAO_REG_28__SCAN_IN), .S(n4134), .Z(U3578)
         );
  MUX2_X1 U4862 ( .A(n4266), .B(DATAO_REG_27__SCAN_IN), .S(n4134), .Z(U3577)
         );
  MUX2_X1 U4863 ( .A(n4285), .B(DATAO_REG_26__SCAN_IN), .S(n4134), .Z(U3576)
         );
  MUX2_X1 U4864 ( .A(n4302), .B(DATAO_REG_25__SCAN_IN), .S(n4134), .Z(U3575)
         );
  MUX2_X1 U4865 ( .A(n4321), .B(DATAO_REG_24__SCAN_IN), .S(n4134), .Z(U3574)
         );
  MUX2_X1 U4866 ( .A(n4125), .B(DATAO_REG_23__SCAN_IN), .S(n4134), .Z(U3573)
         );
  MUX2_X1 U4867 ( .A(n4358), .B(DATAO_REG_22__SCAN_IN), .S(n4134), .Z(U3572)
         );
  MUX2_X1 U4868 ( .A(n4378), .B(DATAO_REG_21__SCAN_IN), .S(n4134), .Z(U3571)
         );
  MUX2_X1 U4869 ( .A(n4126), .B(DATAO_REG_20__SCAN_IN), .S(n4134), .Z(U3570)
         );
  MUX2_X1 U4870 ( .A(n4723), .B(DATAO_REG_17__SCAN_IN), .S(n4134), .Z(U3567)
         );
  MUX2_X1 U4871 ( .A(n4439), .B(DATAO_REG_16__SCAN_IN), .S(n4134), .Z(U3566)
         );
  MUX2_X1 U4872 ( .A(n4494), .B(DATAO_REG_15__SCAN_IN), .S(n4134), .Z(U3565)
         );
  MUX2_X1 U4873 ( .A(n4517), .B(DATAO_REG_14__SCAN_IN), .S(n4134), .Z(U3564)
         );
  MUX2_X1 U4874 ( .A(n4127), .B(DATAO_REG_13__SCAN_IN), .S(n4134), .Z(U3563)
         );
  MUX2_X1 U4875 ( .A(n4128), .B(DATAO_REG_12__SCAN_IN), .S(n4134), .Z(U3562)
         );
  MUX2_X1 U4876 ( .A(n4129), .B(DATAO_REG_11__SCAN_IN), .S(n4134), .Z(U3561)
         );
  MUX2_X1 U4877 ( .A(n4862), .B(DATAO_REG_10__SCAN_IN), .S(n4134), .Z(U3560)
         );
  MUX2_X1 U4878 ( .A(n4130), .B(DATAO_REG_7__SCAN_IN), .S(n4134), .Z(U3557) );
  MUX2_X1 U4879 ( .A(n4131), .B(DATAO_REG_5__SCAN_IN), .S(n4134), .Z(U3555) );
  MUX2_X1 U4880 ( .A(n4132), .B(DATAO_REG_3__SCAN_IN), .S(n4134), .Z(U3553) );
  MUX2_X1 U4881 ( .A(n4133), .B(DATAO_REG_1__SCAN_IN), .S(n4134), .Z(U3551) );
  MUX2_X1 U4882 ( .A(n2234), .B(DATAO_REG_0__SCAN_IN), .S(n4134), .Z(U3550) );
  OAI22_X1 U4883 ( .A1(n4853), .A2(n4136), .B1(STATE_REG_SCAN_IN), .B2(n4135), 
        .ZN(n4137) );
  AOI21_X1 U4884 ( .B1(n4682), .B2(n4848), .A(n4137), .ZN(n4145) );
  OAI211_X1 U4885 ( .C1(n4140), .C2(n4139), .A(n4835), .B(n4138), .ZN(n4144)
         );
  OAI211_X1 U4886 ( .C1(n4150), .C2(n4142), .A(n4833), .B(n4141), .ZN(n4143)
         );
  NAND3_X1 U4887 ( .A1(n4145), .A2(n4144), .A3(n4143), .ZN(U3241) );
  INV_X1 U4888 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4886) );
  NAND2_X1 U4889 ( .A1(n4737), .A2(n4886), .ZN(n4146) );
  AND2_X1 U4890 ( .A1(n4673), .A2(n4146), .ZN(n4736) );
  NAND2_X1 U4891 ( .A1(n4147), .A2(n4149), .ZN(n4148) );
  OAI211_X1 U4892 ( .C1(n4150), .C2(n4149), .A(n4148), .B(n4673), .ZN(n4151)
         );
  OAI211_X1 U4893 ( .C1(IR_REG_0__SCAN_IN), .C2(n4736), .A(n4151), .B(U4043), 
        .ZN(n4172) );
  AOI22_X1 U4894 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4825), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4162) );
  OAI211_X1 U4895 ( .C1(n4154), .C2(n4153), .A(n4835), .B(n4152), .ZN(n4160)
         );
  OAI211_X1 U4896 ( .C1(n4157), .C2(n4156), .A(n4833), .B(n4155), .ZN(n4159)
         );
  NAND2_X1 U4897 ( .A1(n4848), .A2(n4681), .ZN(n4158) );
  AND3_X1 U4898 ( .A1(n4160), .A2(n4159), .A3(n4158), .ZN(n4161) );
  NAND3_X1 U4899 ( .A1(n4172), .A2(n4162), .A3(n4161), .ZN(U3242) );
  NOR2_X1 U4900 ( .A1(n4853), .A2(n4163), .ZN(n4164) );
  AOI211_X1 U4901 ( .C1(n4848), .C2(n4680), .A(n4165), .B(n4164), .ZN(n4171)
         );
  XNOR2_X1 U4902 ( .A(n4166), .B(REG2_REG_4__SCAN_IN), .ZN(n4169) );
  XNOR2_X1 U4903 ( .A(n4167), .B(REG1_REG_4__SCAN_IN), .ZN(n4168) );
  AOI22_X1 U4904 ( .A1(n4833), .A2(n4169), .B1(n4835), .B2(n4168), .ZN(n4170)
         );
  NAND3_X1 U4905 ( .A1(n4172), .A2(n4171), .A3(n4170), .ZN(U3244) );
  XOR2_X1 U4906 ( .A(REG1_REG_17__SCAN_IN), .B(n4690), .Z(n4183) );
  NAND2_X1 U4907 ( .A1(n4677), .A2(REG1_REG_11__SCAN_IN), .ZN(n4173) );
  INV_X1 U4908 ( .A(n4190), .ZN(n4916) );
  NOR2_X1 U4909 ( .A1(n4175), .A2(n4916), .ZN(n4176) );
  INV_X1 U4910 ( .A(n4193), .ZN(n4914) );
  AOI22_X1 U4911 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4914), .B1(n4193), .B2(
        n4613), .ZN(n4791) );
  NOR2_X1 U4912 ( .A1(n4177), .A2(n2313), .ZN(n4178) );
  XNOR2_X1 U4913 ( .A(n2313), .B(n4177), .ZN(n4802) );
  NOR2_X1 U4914 ( .A1(n4803), .A2(n4802), .ZN(n4801) );
  NOR2_X1 U4915 ( .A1(n4178), .A2(n4801), .ZN(n4815) );
  AOI22_X1 U4916 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4196), .B1(n4910), .B2(
        n4179), .ZN(n4814) );
  NOR2_X1 U4917 ( .A1(n4815), .A2(n4814), .ZN(n4813) );
  NAND2_X1 U4918 ( .A1(n4180), .A2(n4909), .ZN(n4181) );
  NAND2_X1 U4919 ( .A1(n4182), .A2(n4183), .ZN(n4684) );
  OAI21_X1 U4920 ( .B1(n4183), .B2(n4182), .A(n4684), .ZN(n4184) );
  AOI22_X1 U4921 ( .A1(n4690), .A2(n4848), .B1(n4835), .B2(n4184), .ZN(n4204)
         );
  AOI21_X1 U4922 ( .B1(n4825), .B2(ADDR_REG_17__SCAN_IN), .A(n4185), .ZN(n4203) );
  NOR2_X1 U4923 ( .A1(n4690), .A2(REG2_REG_17__SCAN_IN), .ZN(n4186) );
  AOI21_X1 U4924 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4690), .A(n4186), .ZN(n4200) );
  INV_X1 U4925 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4795) );
  NOR2_X1 U4926 ( .A1(n4795), .A2(n4914), .ZN(n4794) );
  NAND2_X1 U4927 ( .A1(n4190), .A2(n4191), .ZN(n4192) );
  NOR2_X1 U4928 ( .A1(n2313), .A2(n4194), .ZN(n4195) );
  NOR2_X1 U4929 ( .A1(n4806), .A2(n4805), .ZN(n4804) );
  NOR2_X1 U4930 ( .A1(n4195), .A2(n4804), .ZN(n4818) );
  INV_X1 U4931 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4476) );
  AOI22_X1 U4932 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4196), .B1(n4910), .B2(
        n4476), .ZN(n4817) );
  NOR2_X1 U4933 ( .A1(n4818), .A2(n4817), .ZN(n4816) );
  NAND2_X1 U4934 ( .A1(n4197), .A2(n4909), .ZN(n4198) );
  INV_X1 U4935 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4830) );
  NAND2_X1 U4936 ( .A1(n4689), .A2(n4200), .ZN(n4199) );
  OAI21_X1 U4937 ( .B1(n4200), .B2(n4689), .A(n4199), .ZN(n4201) );
  NAND2_X1 U4938 ( .A1(n4833), .A2(n4201), .ZN(n4202) );
  NAND3_X1 U4939 ( .A1(n4204), .A2(n4203), .A3(n4202), .ZN(U3257) );
  INV_X1 U4940 ( .A(n4205), .ZN(n4216) );
  INV_X1 U4941 ( .A(n4206), .ZN(n4208) );
  INV_X1 U4942 ( .A(n4222), .ZN(n4209) );
  XNOR2_X1 U4943 ( .A(n4210), .B(n4209), .ZN(n4215) );
  AOI22_X1 U4944 ( .A1(n4212), .A2(n4211), .B1(n4225), .B2(n4543), .ZN(n4214)
         );
  NAND2_X1 U4945 ( .A1(n4243), .A2(n4863), .ZN(n4213) );
  OAI211_X1 U4946 ( .C1(n4215), .C2(n4865), .A(n4214), .B(n4213), .ZN(n4549)
         );
  AOI21_X1 U4947 ( .B1(n4216), .B2(n4883), .A(n4549), .ZN(n4228) );
  INV_X1 U4948 ( .A(n4243), .ZN(n4218) );
  XNOR2_X1 U4949 ( .A(n4223), .B(n4222), .ZN(n4548) );
  NAND2_X1 U4950 ( .A1(n4548), .A2(n4431), .ZN(n4227) );
  AOI21_X1 U4951 ( .B1(n4225), .B2(n4224), .A(n4539), .ZN(n4550) );
  AOI22_X1 U4952 ( .A1(n4550), .A2(n4871), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4888), .ZN(n4226) );
  OAI211_X1 U4953 ( .C1(n4888), .C2(n4228), .A(n4227), .B(n4226), .ZN(U3354)
         );
  INV_X1 U4954 ( .A(n4229), .ZN(n4236) );
  AOI22_X1 U4955 ( .A1(n4230), .A2(n4883), .B1(n4888), .B2(
        REG2_REG_28__SCAN_IN), .ZN(n4231) );
  OAI21_X1 U4956 ( .B1(n4232), .B2(n4503), .A(n4231), .ZN(n4233) );
  AOI21_X1 U4957 ( .B1(n4234), .B2(n4530), .A(n4233), .ZN(n4235) );
  OAI21_X1 U4958 ( .B1(n4236), .B2(n4506), .A(n4235), .ZN(U3262) );
  XNOR2_X1 U4959 ( .A(n4238), .B(n4237), .ZN(n4553) );
  AND2_X1 U4960 ( .A1(n4240), .A2(n4239), .ZN(n4242) );
  OR2_X1 U4961 ( .A1(n4242), .A2(n4241), .ZN(n4247) );
  NAND2_X1 U4962 ( .A1(n4243), .A2(n4516), .ZN(n4245) );
  AOI22_X1 U4963 ( .A1(n4285), .A2(n4863), .B1(n4249), .B2(n4543), .ZN(n4244)
         );
  NAND2_X1 U4964 ( .A1(n4245), .A2(n4244), .ZN(n4246) );
  AOI21_X1 U4965 ( .B1(n4247), .B2(n4876), .A(n4246), .ZN(n4554) );
  NOR2_X1 U4966 ( .A1(n4554), .A2(n4888), .ZN(n4255) );
  INV_X1 U4967 ( .A(n4248), .ZN(n4251) );
  NAND2_X1 U4968 ( .A1(n4272), .A2(n4249), .ZN(n4250) );
  NAND2_X1 U4969 ( .A1(n4251), .A2(n4250), .ZN(n4556) );
  AOI22_X1 U4970 ( .A1(n4888), .A2(REG2_REG_27__SCAN_IN), .B1(n4252), .B2(
        n4883), .ZN(n4253) );
  OAI21_X1 U4971 ( .B1(n4556), .B2(n4503), .A(n4253), .ZN(n4254) );
  AOI211_X1 U4972 ( .C1(n4553), .C2(n4431), .A(n4255), .B(n4254), .ZN(n4256)
         );
  INV_X1 U4973 ( .A(n4256), .ZN(U3263) );
  XNOR2_X1 U4974 ( .A(n4257), .B(n4261), .ZN(n4558) );
  INV_X1 U4975 ( .A(n4558), .ZN(n4277) );
  INV_X1 U4976 ( .A(n4258), .ZN(n4259) );
  AOI21_X1 U4977 ( .B1(n4280), .B2(n4260), .A(n4259), .ZN(n4262) );
  XNOR2_X1 U4978 ( .A(n4262), .B(n4261), .ZN(n4263) );
  NAND2_X1 U4979 ( .A1(n4263), .A2(n4876), .ZN(n4268) );
  NOR2_X1 U4980 ( .A1(n4264), .A2(n4858), .ZN(n4265) );
  AOI21_X1 U4981 ( .B1(n4266), .B2(n4516), .A(n4265), .ZN(n4267) );
  OAI211_X1 U4982 ( .C1(n4269), .C2(n4519), .A(n4268), .B(n4267), .ZN(n4557)
         );
  NAND2_X1 U4983 ( .A1(n4288), .A2(n4270), .ZN(n4271) );
  NAND2_X1 U4984 ( .A1(n4272), .A2(n4271), .ZN(n4627) );
  AOI22_X1 U4985 ( .A1(n4888), .A2(REG2_REG_26__SCAN_IN), .B1(n4273), .B2(
        n4883), .ZN(n4274) );
  OAI21_X1 U4986 ( .B1(n4627), .B2(n4503), .A(n4274), .ZN(n4275) );
  AOI21_X1 U4987 ( .B1(n4557), .B2(n4530), .A(n4275), .ZN(n4276) );
  OAI21_X1 U4988 ( .B1(n4277), .B2(n4506), .A(n4276), .ZN(U3264) );
  XOR2_X1 U4989 ( .A(n4282), .B(n4278), .Z(n4562) );
  INV_X1 U4990 ( .A(n4562), .ZN(n4295) );
  NAND2_X1 U4991 ( .A1(n4280), .A2(n4279), .ZN(n4281) );
  XOR2_X1 U4992 ( .A(n4282), .B(n4281), .Z(n4287) );
  OAI22_X1 U4993 ( .A1(n4283), .A2(n4519), .B1(n4289), .B2(n4858), .ZN(n4284)
         );
  AOI21_X1 U4994 ( .B1(n4516), .B2(n4285), .A(n4284), .ZN(n4286) );
  OAI21_X1 U4995 ( .B1(n4287), .B2(n4865), .A(n4286), .ZN(n4561) );
  INV_X1 U4996 ( .A(n4307), .ZN(n4290) );
  OAI21_X1 U4997 ( .B1(n4290), .B2(n4289), .A(n4288), .ZN(n4631) );
  AOI22_X1 U4998 ( .A1(n4888), .A2(REG2_REG_25__SCAN_IN), .B1(n4291), .B2(
        n4883), .ZN(n4292) );
  OAI21_X1 U4999 ( .B1(n4631), .B2(n4503), .A(n4292), .ZN(n4293) );
  AOI21_X1 U5000 ( .B1(n4561), .B2(n4530), .A(n4293), .ZN(n4294) );
  OAI21_X1 U5001 ( .B1(n4295), .B2(n4506), .A(n4294), .ZN(U3265) );
  XNOR2_X1 U5002 ( .A(n4296), .B(n4299), .ZN(n4566) );
  INV_X1 U5003 ( .A(n4566), .ZN(n4312) );
  NAND2_X1 U5004 ( .A1(n4298), .A2(n4297), .ZN(n4300) );
  XNOR2_X1 U5005 ( .A(n4300), .B(n4299), .ZN(n4304) );
  OAI22_X1 U5006 ( .A1(n4348), .A2(n4519), .B1(n4308), .B2(n4858), .ZN(n4301)
         );
  AOI21_X1 U5007 ( .B1(n4516), .B2(n4302), .A(n4301), .ZN(n4303) );
  OAI21_X1 U5008 ( .B1(n4304), .B2(n4865), .A(n4303), .ZN(n4565) );
  INV_X1 U5009 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4306) );
  OAI22_X1 U5010 ( .A1(n4530), .A2(n4306), .B1(n4305), .B2(n4528), .ZN(n4310)
         );
  OAI21_X1 U5011 ( .B1(n4326), .B2(n4308), .A(n4307), .ZN(n4635) );
  NOR2_X1 U5012 ( .A1(n4635), .A2(n4503), .ZN(n4309) );
  AOI211_X1 U5013 ( .C1(n4565), .C2(n4457), .A(n4310), .B(n4309), .ZN(n4311)
         );
  OAI21_X1 U5014 ( .B1(n4312), .B2(n4506), .A(n4311), .ZN(U3266) );
  XOR2_X1 U5015 ( .A(n4318), .B(n4313), .Z(n4570) );
  INV_X1 U5016 ( .A(n4570), .ZN(n4331) );
  OR2_X1 U5017 ( .A1(n4355), .A2(n4314), .ZN(n4316) );
  NAND2_X1 U5018 ( .A1(n4316), .A2(n4315), .ZN(n4343) );
  INV_X1 U5019 ( .A(n4333), .ZN(n4344) );
  NAND2_X1 U5020 ( .A1(n4343), .A2(n4344), .ZN(n4342) );
  NAND2_X1 U5021 ( .A1(n4342), .A2(n4317), .ZN(n4319) );
  XNOR2_X1 U5022 ( .A(n4319), .B(n4318), .ZN(n4324) );
  AOI22_X1 U5023 ( .A1(n4321), .A2(n4516), .B1(n4543), .B2(n4320), .ZN(n4323)
         );
  NAND2_X1 U5024 ( .A1(n4358), .A2(n4863), .ZN(n4322) );
  OAI211_X1 U5025 ( .C1(n4324), .C2(n4865), .A(n4323), .B(n4322), .ZN(n4569)
         );
  NOR2_X1 U5026 ( .A1(n4335), .A2(n2934), .ZN(n4325) );
  OR2_X1 U5027 ( .A1(n4326), .A2(n4325), .ZN(n4639) );
  AOI22_X1 U5028 ( .A1(n4888), .A2(REG2_REG_23__SCAN_IN), .B1(n4327), .B2(
        n4883), .ZN(n4328) );
  OAI21_X1 U5029 ( .B1(n4639), .B2(n4503), .A(n4328), .ZN(n4329) );
  AOI21_X1 U5030 ( .B1(n4569), .B2(n4457), .A(n4329), .ZN(n4330) );
  OAI21_X1 U5031 ( .B1(n4331), .B2(n4506), .A(n4330), .ZN(U3267) );
  OAI21_X1 U5032 ( .B1(n4334), .B2(n4333), .A(n4332), .ZN(n4577) );
  INV_X1 U5033 ( .A(n4335), .ZN(n4574) );
  NAND2_X1 U5034 ( .A1(n4361), .A2(n4336), .ZN(n4573) );
  AND2_X1 U5035 ( .A1(n4573), .A2(n4871), .ZN(n4341) );
  INV_X1 U5036 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4339) );
  INV_X1 U5037 ( .A(n4337), .ZN(n4338) );
  OAI22_X1 U5038 ( .A1(n4530), .A2(n4339), .B1(n4338), .B2(n4528), .ZN(n4340)
         );
  AOI21_X1 U5039 ( .B1(n4574), .B2(n4341), .A(n4340), .ZN(n4352) );
  OAI21_X1 U5040 ( .B1(n4344), .B2(n4343), .A(n4342), .ZN(n4350) );
  OR2_X1 U5041 ( .A1(n4345), .A2(n4858), .ZN(n4347) );
  NAND2_X1 U5042 ( .A1(n4378), .A2(n4863), .ZN(n4346) );
  OAI211_X1 U5043 ( .C1(n4348), .C2(n4878), .A(n4347), .B(n4346), .ZN(n4349)
         );
  AOI21_X1 U5044 ( .B1(n4350), .B2(n4876), .A(n4349), .ZN(n4576) );
  OR2_X1 U5045 ( .A1(n4576), .A2(n4888), .ZN(n4351) );
  OAI211_X1 U5046 ( .C1(n4577), .C2(n4506), .A(n4352), .B(n4351), .ZN(U3268)
         );
  XOR2_X1 U5047 ( .A(n4354), .B(n4353), .Z(n4579) );
  INV_X1 U5048 ( .A(n4579), .ZN(n4370) );
  XNOR2_X1 U5049 ( .A(n4355), .B(n4354), .ZN(n4356) );
  NAND2_X1 U5050 ( .A1(n4356), .A2(n4876), .ZN(n4360) );
  AOI22_X1 U5051 ( .A1(n4358), .A2(n4516), .B1(n4543), .B2(n4357), .ZN(n4359)
         );
  OAI211_X1 U5052 ( .C1(n4400), .C2(n4519), .A(n4360), .B(n4359), .ZN(n4578)
         );
  INV_X1 U5053 ( .A(n4384), .ZN(n4363) );
  OAI21_X1 U5054 ( .B1(n4363), .B2(n4362), .A(n4361), .ZN(n4644) );
  NOR2_X1 U5055 ( .A1(n4644), .A2(n4503), .ZN(n4368) );
  INV_X1 U5056 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4366) );
  INV_X1 U5057 ( .A(n4364), .ZN(n4365) );
  OAI22_X1 U5058 ( .A1(n4530), .A2(n4366), .B1(n4365), .B2(n4528), .ZN(n4367)
         );
  AOI211_X1 U5059 ( .C1(n4578), .C2(n4457), .A(n4368), .B(n4367), .ZN(n4369)
         );
  OAI21_X1 U5060 ( .B1(n4370), .B2(n4506), .A(n4369), .ZN(U3269) );
  XNOR2_X1 U5061 ( .A(n4371), .B(n4376), .ZN(n4582) );
  INV_X1 U5062 ( .A(n4372), .ZN(n4373) );
  NAND2_X1 U5063 ( .A1(n4374), .A2(n4373), .ZN(n4375) );
  XOR2_X1 U5064 ( .A(n4376), .B(n4375), .Z(n4382) );
  AOI22_X1 U5065 ( .A1(n4378), .A2(n4516), .B1(n4543), .B2(n4377), .ZN(n4379)
         );
  OAI21_X1 U5066 ( .B1(n4380), .B2(n4519), .A(n4379), .ZN(n4381) );
  AOI21_X1 U5067 ( .B1(n4382), .B2(n4876), .A(n4381), .ZN(n4383) );
  OAI21_X1 U5068 ( .B1(n4582), .B2(n4523), .A(n4383), .ZN(n4583) );
  NAND2_X1 U5069 ( .A1(n4583), .A2(n4530), .ZN(n4391) );
  OAI21_X1 U5070 ( .B1(n4405), .B2(n4385), .A(n4384), .ZN(n4648) );
  INV_X1 U5071 ( .A(n4648), .ZN(n4389) );
  INV_X1 U5072 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4387) );
  OAI22_X1 U5073 ( .A1(n4457), .A2(n4387), .B1(n4386), .B2(n4528), .ZN(n4388)
         );
  AOI21_X1 U5074 ( .B1(n4389), .B2(n4871), .A(n4388), .ZN(n4390) );
  OAI211_X1 U5075 ( .C1(n4582), .C2(n4535), .A(n4391), .B(n4390), .ZN(U3270)
         );
  XNOR2_X1 U5076 ( .A(n4392), .B(n4399), .ZN(n4588) );
  INV_X1 U5077 ( .A(n4588), .ZN(n4414) );
  OAI21_X1 U5078 ( .B1(n4434), .B2(n4394), .A(n4393), .ZN(n4416) );
  INV_X1 U5079 ( .A(n4395), .ZN(n4397) );
  OAI21_X1 U5080 ( .B1(n4416), .B2(n4397), .A(n4396), .ZN(n4398) );
  XOR2_X1 U5081 ( .A(n4399), .B(n4398), .Z(n4404) );
  OAI22_X1 U5082 ( .A1(n4400), .A2(n4878), .B1(n4858), .B2(n4407), .ZN(n4401)
         );
  AOI21_X1 U5083 ( .B1(n4863), .B2(n4402), .A(n4401), .ZN(n4403) );
  OAI21_X1 U5084 ( .B1(n4404), .B2(n4865), .A(n4403), .ZN(n4587) );
  INV_X1 U5085 ( .A(n4405), .ZN(n4406) );
  OAI21_X1 U5086 ( .B1(n4425), .B2(n4407), .A(n4406), .ZN(n4652) );
  NOR2_X1 U5087 ( .A1(n4652), .A2(n4503), .ZN(n4412) );
  INV_X1 U5088 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4410) );
  INV_X1 U5089 ( .A(n4408), .ZN(n4409) );
  OAI22_X1 U5090 ( .A1(n4457), .A2(n4410), .B1(n4409), .B2(n4528), .ZN(n4411)
         );
  AOI211_X1 U5091 ( .C1(n4587), .C2(n4457), .A(n4412), .B(n4411), .ZN(n4413)
         );
  OAI21_X1 U5092 ( .B1(n4414), .B2(n4506), .A(n4413), .ZN(U3271) );
  XNOR2_X1 U5093 ( .A(n4416), .B(n4415), .ZN(n4420) );
  AOI22_X1 U5094 ( .A1(n4710), .A2(n4516), .B1(n4713), .B2(n4543), .ZN(n4417)
         );
  OAI21_X1 U5095 ( .B1(n4418), .B2(n4519), .A(n4417), .ZN(n4419) );
  AOI21_X1 U5096 ( .B1(n4420), .B2(n4876), .A(n4419), .ZN(n4593) );
  OAI21_X1 U5097 ( .B1(n4423), .B2(n4422), .A(n4421), .ZN(n4591) );
  NAND2_X1 U5098 ( .A1(n4444), .A2(n4713), .ZN(n4424) );
  NAND2_X1 U5099 ( .A1(n4424), .A2(n4971), .ZN(n4426) );
  OR2_X1 U5100 ( .A1(n4426), .A2(n4425), .ZN(n4592) );
  AOI22_X1 U5101 ( .A1(n4888), .A2(REG2_REG_18__SCAN_IN), .B1(n4427), .B2(
        n4883), .ZN(n4428) );
  OAI21_X1 U5102 ( .B1(n4592), .B2(n4429), .A(n4428), .ZN(n4430) );
  AOI21_X1 U5103 ( .B1(n4591), .B2(n4431), .A(n4430), .ZN(n4432) );
  OAI21_X1 U5104 ( .B1(n4888), .B2(n4593), .A(n4432), .ZN(U3272) );
  XOR2_X1 U5105 ( .A(n4435), .B(n4433), .Z(n4596) );
  INV_X1 U5106 ( .A(n4596), .ZN(n4449) );
  XOR2_X1 U5107 ( .A(n4435), .B(n4434), .Z(n4441) );
  OAI22_X1 U5108 ( .A1(n4437), .A2(n4878), .B1(n4436), .B2(n4858), .ZN(n4438)
         );
  AOI21_X1 U5109 ( .B1(n4863), .B2(n4439), .A(n4438), .ZN(n4440) );
  OAI21_X1 U5110 ( .B1(n4441), .B2(n4865), .A(n4440), .ZN(n4595) );
  NAND2_X1 U5111 ( .A1(n4454), .A2(n4442), .ZN(n4443) );
  NAND2_X1 U5112 ( .A1(n4444), .A2(n4443), .ZN(n4657) );
  AOI22_X1 U5113 ( .A1(n4888), .A2(REG2_REG_17__SCAN_IN), .B1(n4445), .B2(
        n4883), .ZN(n4446) );
  OAI21_X1 U5114 ( .B1(n4657), .B2(n4503), .A(n4446), .ZN(n4447) );
  AOI21_X1 U5115 ( .B1(n4595), .B2(n4457), .A(n4447), .ZN(n4448) );
  OAI21_X1 U5116 ( .B1(n4449), .B2(n4506), .A(n4448), .ZN(U3273) );
  OAI21_X1 U5117 ( .B1(n4452), .B2(n4451), .A(n4450), .ZN(n4602) );
  OR2_X1 U5118 ( .A1(n4473), .A2(n4453), .ZN(n4455) );
  AND2_X1 U5119 ( .A1(n4455), .A2(n4454), .ZN(n4600) );
  OAI22_X1 U5120 ( .A1(n4457), .A2(n4830), .B1(n4456), .B2(n4528), .ZN(n4458)
         );
  AOI21_X1 U5121 ( .B1(n4600), .B2(n4871), .A(n4458), .ZN(n4467) );
  OAI211_X1 U5122 ( .C1(n4461), .C2(n4460), .A(n4459), .B(n4876), .ZN(n4464)
         );
  AOI22_X1 U5123 ( .A1(n4723), .A2(n4516), .B1(n4462), .B2(n4543), .ZN(n4463)
         );
  OAI211_X1 U5124 ( .C1(n4465), .C2(n4519), .A(n4464), .B(n4463), .ZN(n4599)
         );
  NAND2_X1 U5125 ( .A1(n4599), .A2(n4530), .ZN(n4466) );
  OAI211_X1 U5126 ( .C1(n4602), .C2(n4506), .A(n4467), .B(n4466), .ZN(U3274)
         );
  INV_X1 U5127 ( .A(n4468), .ZN(n4470) );
  NOR2_X1 U5128 ( .A1(n4470), .A2(n4469), .ZN(n4490) );
  INV_X1 U5129 ( .A(n4491), .ZN(n4489) );
  NAND2_X1 U5130 ( .A1(n4490), .A2(n4489), .ZN(n4488) );
  NAND2_X1 U5131 ( .A1(n4488), .A2(n4471), .ZN(n4472) );
  XOR2_X1 U5132 ( .A(n4481), .B(n4472), .Z(n4606) );
  AOI21_X1 U5133 ( .B1(n4474), .B2(n4500), .A(n4473), .ZN(n4603) );
  OAI22_X1 U5134 ( .A1(n4530), .A2(n4476), .B1(n4475), .B2(n4528), .ZN(n4486)
         );
  OAI22_X1 U5135 ( .A1(n4478), .A2(n4878), .B1(n4858), .B2(n4477), .ZN(n4484)
         );
  INV_X1 U5136 ( .A(n4479), .ZN(n4480) );
  AOI211_X1 U5137 ( .C1(n4482), .C2(n4481), .A(n4865), .B(n4480), .ZN(n4483)
         );
  AOI211_X1 U5138 ( .C1(n4863), .C2(n4517), .A(n4484), .B(n4483), .ZN(n4605)
         );
  NOR2_X1 U5139 ( .A1(n4605), .A2(n4888), .ZN(n4485) );
  AOI211_X1 U5140 ( .C1(n4603), .C2(n4871), .A(n4486), .B(n4485), .ZN(n4487)
         );
  OAI21_X1 U5141 ( .B1(n4606), .B2(n4506), .A(n4487), .ZN(U3275) );
  OAI21_X1 U5142 ( .B1(n4490), .B2(n4489), .A(n4488), .ZN(n4608) );
  INV_X1 U5143 ( .A(n4608), .ZN(n4507) );
  XNOR2_X1 U5144 ( .A(n4492), .B(n4491), .ZN(n4493) );
  NAND2_X1 U5145 ( .A1(n4493), .A2(n4876), .ZN(n4496) );
  AOI22_X1 U5146 ( .A1(n4494), .A2(n4516), .B1(n4498), .B2(n4543), .ZN(n4495)
         );
  OAI211_X1 U5147 ( .C1(n4497), .C2(n4519), .A(n4496), .B(n4495), .ZN(n4607)
         );
  NAND2_X1 U5148 ( .A1(n4524), .A2(n4498), .ZN(n4499) );
  NAND2_X1 U5149 ( .A1(n4500), .A2(n4499), .ZN(n4663) );
  AOI22_X1 U5150 ( .A1(n4888), .A2(REG2_REG_14__SCAN_IN), .B1(n4501), .B2(
        n4883), .ZN(n4502) );
  OAI21_X1 U5151 ( .B1(n4663), .B2(n4503), .A(n4502), .ZN(n4504) );
  AOI21_X1 U5152 ( .B1(n4607), .B2(n4530), .A(n4504), .ZN(n4505) );
  OAI21_X1 U5153 ( .B1(n4507), .B2(n4506), .A(n4505), .ZN(U3276) );
  XNOR2_X1 U5154 ( .A(n4508), .B(n4513), .ZN(n4610) );
  INV_X1 U5155 ( .A(n4509), .ZN(n4511) );
  OAI21_X1 U5156 ( .B1(n4512), .B2(n4511), .A(n4510), .ZN(n4514) );
  XNOR2_X1 U5157 ( .A(n4514), .B(n4513), .ZN(n4521) );
  AOI22_X1 U5158 ( .A1(n4517), .A2(n4516), .B1(n4515), .B2(n4543), .ZN(n4518)
         );
  OAI21_X1 U5159 ( .B1(n4860), .B2(n4519), .A(n4518), .ZN(n4520) );
  AOI21_X1 U5160 ( .B1(n4521), .B2(n4876), .A(n4520), .ZN(n4522) );
  OAI21_X1 U5161 ( .B1(n4610), .B2(n4523), .A(n4522), .ZN(n4611) );
  NAND2_X1 U5162 ( .A1(n4611), .A2(n4530), .ZN(n4534) );
  INV_X1 U5163 ( .A(n3475), .ZN(n4526) );
  OAI21_X1 U5164 ( .B1(n4526), .B2(n4525), .A(n4524), .ZN(n4667) );
  INV_X1 U5165 ( .A(n4667), .ZN(n4532) );
  INV_X1 U5166 ( .A(n4527), .ZN(n4529) );
  OAI22_X1 U5167 ( .A1(n4530), .A2(n4795), .B1(n4529), .B2(n4528), .ZN(n4531)
         );
  AOI21_X1 U5168 ( .B1(n4532), .B2(n4871), .A(n4531), .ZN(n4533) );
  OAI211_X1 U5169 ( .C1(n4610), .C2(n4535), .A(n4534), .B(n4533), .ZN(U3277)
         );
  INV_X1 U5170 ( .A(n4618), .ZN(n4536) );
  NAND2_X1 U5171 ( .A1(n4730), .A2(n4536), .ZN(n4538) );
  NAND2_X1 U5172 ( .A1(n4990), .A2(n4729), .ZN(n4537) );
  OAI211_X1 U5173 ( .C1(n4990), .C2(n3488), .A(n4538), .B(n4537), .ZN(U3549)
         );
  INV_X1 U5174 ( .A(n4539), .ZN(n4542) );
  INV_X1 U5175 ( .A(n4540), .ZN(n4541) );
  AOI21_X1 U5176 ( .B1(n4544), .B2(n4542), .A(n4541), .ZN(n4733) );
  INV_X1 U5177 ( .A(n4733), .ZN(n4621) );
  NAND2_X1 U5178 ( .A1(n4544), .A2(n4543), .ZN(n4545) );
  AND2_X1 U5179 ( .A1(n4546), .A2(n4545), .ZN(n4735) );
  MUX2_X1 U5180 ( .A(n3090), .B(n4735), .S(n4990), .Z(n4547) );
  OAI21_X1 U5181 ( .B1(n4621), .B2(n4618), .A(n4547), .ZN(U3548) );
  NAND2_X1 U5182 ( .A1(n4548), .A2(n4968), .ZN(n4552) );
  AOI21_X1 U5183 ( .B1(n4971), .B2(n4550), .A(n4549), .ZN(n4551) );
  NAND2_X1 U5184 ( .A1(n4552), .A2(n4551), .ZN(n4622) );
  MUX2_X1 U5185 ( .A(REG1_REG_29__SCAN_IN), .B(n4622), .S(n4990), .Z(U3547) );
  NAND2_X1 U5186 ( .A1(n4553), .A2(n4968), .ZN(n4555) );
  OAI211_X1 U5187 ( .C1(n4965), .C2(n4556), .A(n4555), .B(n4554), .ZN(n4623)
         );
  MUX2_X1 U5188 ( .A(REG1_REG_27__SCAN_IN), .B(n4623), .S(n4990), .Z(U3545) );
  AOI21_X1 U5189 ( .B1(n4558), .B2(n4968), .A(n4557), .ZN(n4624) );
  MUX2_X1 U5190 ( .A(n4559), .B(n4624), .S(n4990), .Z(n4560) );
  OAI21_X1 U5191 ( .B1(n4618), .B2(n4627), .A(n4560), .ZN(U3544) );
  AOI21_X1 U5192 ( .B1(n4562), .B2(n4968), .A(n4561), .ZN(n4628) );
  MUX2_X1 U5193 ( .A(n4563), .B(n4628), .S(n4990), .Z(n4564) );
  OAI21_X1 U5194 ( .B1(n4618), .B2(n4631), .A(n4564), .ZN(U3543) );
  INV_X1 U5195 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4567) );
  AOI21_X1 U5196 ( .B1(n4566), .B2(n4968), .A(n4565), .ZN(n4632) );
  MUX2_X1 U5197 ( .A(n4567), .B(n4632), .S(n4990), .Z(n4568) );
  OAI21_X1 U5198 ( .B1(n4618), .B2(n4635), .A(n4568), .ZN(U3542) );
  AOI21_X1 U5199 ( .B1(n4570), .B2(n4968), .A(n4569), .ZN(n4636) );
  MUX2_X1 U5200 ( .A(n4571), .B(n4636), .S(n4990), .Z(n4572) );
  OAI21_X1 U5201 ( .B1(n4618), .B2(n4639), .A(n4572), .ZN(U3541) );
  NAND3_X1 U5202 ( .A1(n4574), .A2(n4573), .A3(n4971), .ZN(n4575) );
  OAI211_X1 U5203 ( .C1(n4577), .C2(n4952), .A(n4576), .B(n4575), .ZN(n4640)
         );
  MUX2_X1 U5204 ( .A(REG1_REG_22__SCAN_IN), .B(n4640), .S(n4990), .Z(U3540) );
  AOI21_X1 U5205 ( .B1(n4579), .B2(n4968), .A(n4578), .ZN(n4641) );
  MUX2_X1 U5206 ( .A(n4580), .B(n4641), .S(n4990), .Z(n4581) );
  OAI21_X1 U5207 ( .B1(n4618), .B2(n4644), .A(n4581), .ZN(U3539) );
  INV_X1 U5208 ( .A(n4941), .ZN(n4972) );
  INV_X1 U5209 ( .A(n4582), .ZN(n4584) );
  AOI21_X1 U5210 ( .B1(n4972), .B2(n4584), .A(n4583), .ZN(n4645) );
  MUX2_X1 U5211 ( .A(n4585), .B(n4645), .S(n4990), .Z(n4586) );
  OAI21_X1 U5212 ( .B1(n4618), .B2(n4648), .A(n4586), .ZN(U3538) );
  AOI21_X1 U5213 ( .B1(n4588), .B2(n4968), .A(n4587), .ZN(n4649) );
  MUX2_X1 U5214 ( .A(n4589), .B(n4649), .S(n4990), .Z(n4590) );
  OAI21_X1 U5215 ( .B1(n4618), .B2(n4652), .A(n4590), .ZN(U3537) );
  INV_X1 U5216 ( .A(n4591), .ZN(n4594) );
  OAI211_X1 U5217 ( .C1(n4594), .C2(n4952), .A(n4593), .B(n4592), .ZN(n4653)
         );
  MUX2_X1 U5218 ( .A(REG1_REG_18__SCAN_IN), .B(n4653), .S(n4990), .Z(U3536) );
  AOI21_X1 U5219 ( .B1(n4596), .B2(n4968), .A(n4595), .ZN(n4654) );
  MUX2_X1 U5220 ( .A(n4597), .B(n4654), .S(n4990), .Z(n4598) );
  OAI21_X1 U5221 ( .B1(n4618), .B2(n4657), .A(n4598), .ZN(U3535) );
  AOI21_X1 U5222 ( .B1(n4971), .B2(n4600), .A(n4599), .ZN(n4601) );
  OAI21_X1 U5223 ( .B1(n4602), .B2(n4952), .A(n4601), .ZN(n4658) );
  MUX2_X1 U5224 ( .A(REG1_REG_16__SCAN_IN), .B(n4658), .S(n4990), .Z(U3534) );
  NAND2_X1 U5225 ( .A1(n4603), .A2(n4971), .ZN(n4604) );
  OAI211_X1 U5226 ( .C1(n4606), .C2(n4952), .A(n4605), .B(n4604), .ZN(n4659)
         );
  MUX2_X1 U5227 ( .A(REG1_REG_15__SCAN_IN), .B(n4659), .S(n4990), .Z(U3533) );
  AOI21_X1 U5228 ( .B1(n4608), .B2(n4968), .A(n4607), .ZN(n4660) );
  MUX2_X1 U5229 ( .A(n4803), .B(n4660), .S(n4990), .Z(n4609) );
  OAI21_X1 U5230 ( .B1(n4618), .B2(n4663), .A(n4609), .ZN(U3532) );
  INV_X1 U5231 ( .A(n4610), .ZN(n4612) );
  AOI21_X1 U5232 ( .B1(n4972), .B2(n4612), .A(n4611), .ZN(n4664) );
  MUX2_X1 U5233 ( .A(n4613), .B(n4664), .S(n4990), .Z(n4614) );
  OAI21_X1 U5234 ( .B1(n4618), .B2(n4667), .A(n4614), .ZN(U3531) );
  AOI21_X1 U5235 ( .B1(n4616), .B2(n4968), .A(n4615), .ZN(n4668) );
  MUX2_X1 U5236 ( .A(n2642), .B(n4668), .S(n4990), .Z(n4617) );
  OAI21_X1 U5237 ( .B1(n4672), .B2(n4618), .A(n4617), .ZN(U3530) );
  MUX2_X1 U5238 ( .A(n4619), .B(n4735), .S(n4978), .Z(n4620) );
  OAI21_X1 U5239 ( .B1(n4621), .B2(n4671), .A(n4620), .ZN(U3516) );
  MUX2_X1 U5240 ( .A(REG0_REG_29__SCAN_IN), .B(n4622), .S(n4978), .Z(U3515) );
  MUX2_X1 U5241 ( .A(REG0_REG_27__SCAN_IN), .B(n4623), .S(n4978), .Z(U3513) );
  MUX2_X1 U5242 ( .A(n4625), .B(n4624), .S(n4978), .Z(n4626) );
  OAI21_X1 U5243 ( .B1(n4627), .B2(n4671), .A(n4626), .ZN(U3512) );
  MUX2_X1 U5244 ( .A(n4629), .B(n4628), .S(n4978), .Z(n4630) );
  OAI21_X1 U5245 ( .B1(n4631), .B2(n4671), .A(n4630), .ZN(U3511) );
  INV_X1 U5246 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4633) );
  MUX2_X1 U5247 ( .A(n4633), .B(n4632), .S(n4978), .Z(n4634) );
  OAI21_X1 U5248 ( .B1(n4635), .B2(n4671), .A(n4634), .ZN(U3510) );
  INV_X1 U5249 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4637) );
  MUX2_X1 U5250 ( .A(n4637), .B(n4636), .S(n4978), .Z(n4638) );
  OAI21_X1 U5251 ( .B1(n4639), .B2(n4671), .A(n4638), .ZN(U3509) );
  MUX2_X1 U5252 ( .A(REG0_REG_22__SCAN_IN), .B(n4640), .S(n4978), .Z(U3508) );
  INV_X1 U5253 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4642) );
  MUX2_X1 U5254 ( .A(n4642), .B(n4641), .S(n4978), .Z(n4643) );
  OAI21_X1 U5255 ( .B1(n4644), .B2(n4671), .A(n4643), .ZN(U3507) );
  INV_X1 U5256 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4646) );
  MUX2_X1 U5257 ( .A(n4646), .B(n4645), .S(n4978), .Z(n4647) );
  OAI21_X1 U5258 ( .B1(n4648), .B2(n4671), .A(n4647), .ZN(U3506) );
  INV_X1 U5259 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4650) );
  MUX2_X1 U5260 ( .A(n4650), .B(n4649), .S(n4978), .Z(n4651) );
  OAI21_X1 U5261 ( .B1(n4652), .B2(n4671), .A(n4651), .ZN(U3505) );
  MUX2_X1 U5262 ( .A(REG0_REG_18__SCAN_IN), .B(n4653), .S(n4978), .Z(U3503) );
  INV_X1 U5263 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4655) );
  MUX2_X1 U5264 ( .A(n4655), .B(n4654), .S(n4978), .Z(n4656) );
  OAI21_X1 U5265 ( .B1(n4657), .B2(n4671), .A(n4656), .ZN(U3501) );
  MUX2_X1 U5266 ( .A(REG0_REG_16__SCAN_IN), .B(n4658), .S(n4978), .Z(U3499) );
  MUX2_X1 U5267 ( .A(REG0_REG_15__SCAN_IN), .B(n4659), .S(n4978), .Z(U3497) );
  INV_X1 U5268 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4661) );
  MUX2_X1 U5269 ( .A(n4661), .B(n4660), .S(n4978), .Z(n4662) );
  OAI21_X1 U5270 ( .B1(n4663), .B2(n4671), .A(n4662), .ZN(U3495) );
  INV_X1 U5271 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4665) );
  MUX2_X1 U5272 ( .A(n4665), .B(n4664), .S(n4978), .Z(n4666) );
  OAI21_X1 U5273 ( .B1(n4667), .B2(n4671), .A(n4666), .ZN(U3493) );
  INV_X1 U5274 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4669) );
  MUX2_X1 U5275 ( .A(n4669), .B(n4668), .S(n4978), .Z(n4670) );
  OAI21_X1 U5276 ( .B1(n4672), .B2(n4671), .A(n4670), .ZN(U3491) );
  MUX2_X1 U5277 ( .A(DATAI_28_), .B(n4673), .S(STATE_REG_SCAN_IN), .Z(U3324)
         );
  MUX2_X1 U5278 ( .A(n2854), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5279 ( .A(n4674), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U5280 ( .A(DATAI_22_), .B(n4675), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U5281 ( .A(DATAI_20_), .B(n4676), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5282 ( .A(n4690), .B(DATAI_17_), .S(U3149), .Z(U3335) );
  MUX2_X1 U5283 ( .A(n4677), .B(DATAI_11_), .S(U3149), .Z(U3341) );
  MUX2_X1 U5284 ( .A(DATAI_9_), .B(n4678), .S(STATE_REG_SCAN_IN), .Z(U3343) );
  MUX2_X1 U5285 ( .A(n4679), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5286 ( .A(DATAI_4_), .B(n4680), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5287 ( .A(n4705), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5288 ( .A(n4681), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5289 ( .A(n4682), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  INV_X1 U5290 ( .A(n4847), .ZN(n4907) );
  AOI22_X1 U5291 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4907), .B1(n4847), .B2(
        n4683), .ZN(n4840) );
  XNOR2_X1 U5292 ( .A(n4685), .B(REG1_REG_19__SCAN_IN), .ZN(n4686) );
  AOI22_X1 U5293 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4907), .B1(n4847), .B2(
        n4687), .ZN(n4846) );
  INV_X1 U5294 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4688) );
  AOI21_X1 U5295 ( .B1(n4847), .B2(REG2_REG_18__SCAN_IN), .A(n4844), .ZN(n4692) );
  MUX2_X1 U5296 ( .A(n4410), .B(REG2_REG_19__SCAN_IN), .S(n4695), .Z(n4691) );
  XNOR2_X1 U5297 ( .A(n4692), .B(n4691), .ZN(n4697) );
  AOI21_X1 U5298 ( .B1(n4825), .B2(ADDR_REG_19__SCAN_IN), .A(n4693), .ZN(n4694) );
  OAI21_X1 U5299 ( .B1(n4838), .B2(n4695), .A(n4694), .ZN(n4696) );
  AOI21_X1 U5300 ( .B1(n4697), .B2(n4833), .A(n4696), .ZN(n4698) );
  OAI21_X1 U5301 ( .B1(n4699), .B2(n4839), .A(n4698), .ZN(U3259) );
  AOI21_X1 U5302 ( .B1(n4825), .B2(ADDR_REG_3__SCAN_IN), .A(n4700), .ZN(n4709)
         );
  OAI211_X1 U5303 ( .C1(REG1_REG_3__SCAN_IN), .C2(n4702), .A(n4835), .B(n4701), 
        .ZN(n4708) );
  OAI211_X1 U5304 ( .C1(REG2_REG_3__SCAN_IN), .C2(n4704), .A(n4833), .B(n4703), 
        .ZN(n4707) );
  NAND2_X1 U5305 ( .A1(n4848), .A2(n4705), .ZN(n4706) );
  NAND4_X1 U5306 ( .A1(n4709), .A2(n4708), .A3(n4707), .A4(n4706), .ZN(U3243)
         );
  AOI22_X1 U5307 ( .A1(n4713), .A2(n4712), .B1(n4711), .B2(n4710), .ZN(n4726)
         );
  NAND2_X1 U5308 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4851) );
  INV_X1 U5309 ( .A(n4851), .ZN(n4722) );
  INV_X1 U5310 ( .A(n4715), .ZN(n4717) );
  NAND2_X1 U5311 ( .A1(n4717), .A2(n4716), .ZN(n4718) );
  XNOR2_X1 U5312 ( .A(n4714), .B(n4718), .ZN(n4720) );
  NOR2_X1 U5313 ( .A1(n4720), .A2(n4719), .ZN(n4721) );
  AOI211_X1 U5314 ( .C1(n4724), .C2(n4723), .A(n4722), .B(n4721), .ZN(n4725)
         );
  OAI211_X1 U5315 ( .C1(n4728), .C2(n4727), .A(n4726), .B(n4725), .ZN(U3235)
         );
  AOI22_X1 U5316 ( .A1(n4730), .A2(n4871), .B1(n4530), .B2(n4729), .ZN(n4731)
         );
  OAI21_X1 U5317 ( .B1(n4530), .B2(n4732), .A(n4731), .ZN(U3260) );
  AOI22_X1 U5318 ( .A1(n4733), .A2(n4871), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4888), .ZN(n4734) );
  OAI21_X1 U5319 ( .B1(n4888), .B2(n4735), .A(n4734), .ZN(U3261) );
  OAI21_X1 U5320 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4737), .A(n4736), .ZN(n4738)
         );
  XOR2_X1 U5321 ( .A(n2444), .B(n4738), .Z(n4740) );
  AOI22_X1 U5322 ( .A1(n4740), .A2(n4739), .B1(REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4741) );
  OAI21_X1 U5323 ( .B1(n4742), .B2(n4853), .A(n4741), .ZN(U3240) );
  NOR2_X1 U5324 ( .A1(n4743), .A2(n4853), .ZN(n4744) );
  AOI211_X1 U5325 ( .C1(n4848), .C2(n4746), .A(n4745), .B(n4744), .ZN(n4753)
         );
  OAI211_X1 U5326 ( .C1(REG1_REG_6__SCAN_IN), .C2(n4748), .A(n4835), .B(n4747), 
        .ZN(n4752) );
  OAI211_X1 U5327 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4750), .A(n4833), .B(n4749), 
        .ZN(n4751) );
  NAND3_X1 U5328 ( .A1(n4753), .A2(n4752), .A3(n4751), .ZN(U3246) );
  AOI22_X1 U5329 ( .A1(REG1_REG_7__SCAN_IN), .A2(n4754), .B1(n4922), .B2(n2550), .ZN(n4757) );
  OAI21_X1 U5330 ( .B1(n4757), .B2(n4756), .A(n4835), .ZN(n4755) );
  AOI21_X1 U5331 ( .B1(n4757), .B2(n4756), .A(n4755), .ZN(n4758) );
  AOI211_X1 U5332 ( .C1(n4825), .C2(ADDR_REG_7__SCAN_IN), .A(n4759), .B(n4758), 
        .ZN(n4764) );
  OAI211_X1 U5333 ( .C1(n4762), .C2(n4761), .A(n4833), .B(n4760), .ZN(n4763)
         );
  OAI211_X1 U5334 ( .C1(n4838), .C2(n4922), .A(n4764), .B(n4763), .ZN(U3247)
         );
  AOI211_X1 U5335 ( .C1(n2568), .C2(n4766), .A(n4765), .B(n4839), .ZN(n4767)
         );
  AOI211_X1 U5336 ( .C1(n4825), .C2(ADDR_REG_8__SCAN_IN), .A(n4768), .B(n4767), 
        .ZN(n4772) );
  OAI211_X1 U5337 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4770), .A(n4833), .B(n4769), 
        .ZN(n4771) );
  OAI211_X1 U5338 ( .C1(n4838), .C2(n4920), .A(n4772), .B(n4771), .ZN(U3248)
         );
  AOI211_X1 U5339 ( .C1(n2604), .C2(n4774), .A(n4773), .B(n4839), .ZN(n4776)
         );
  AOI211_X1 U5340 ( .C1(n4825), .C2(ADDR_REG_10__SCAN_IN), .A(n4776), .B(n4775), .ZN(n4780) );
  OAI211_X1 U5341 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4778), .A(n4833), .B(n4777), .ZN(n4779) );
  OAI211_X1 U5342 ( .C1(n4838), .C2(n3393), .A(n4780), .B(n4779), .ZN(U3250)
         );
  AOI211_X1 U5343 ( .C1(n2642), .C2(n4782), .A(n4781), .B(n4839), .ZN(n4785)
         );
  INV_X1 U5344 ( .A(n4783), .ZN(n4784) );
  AOI211_X1 U5345 ( .C1(n4825), .C2(ADDR_REG_12__SCAN_IN), .A(n4785), .B(n4784), .ZN(n4789) );
  OAI211_X1 U5346 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4787), .A(n4833), .B(n4786), .ZN(n4788) );
  OAI211_X1 U5347 ( .C1(n4838), .C2(n4916), .A(n4789), .B(n4788), .ZN(U3252)
         );
  AOI211_X1 U5348 ( .C1(n2256), .C2(n4791), .A(n4790), .B(n4839), .ZN(n4792)
         );
  AOI211_X1 U5349 ( .C1(ADDR_REG_13__SCAN_IN), .C2(n4825), .A(n4793), .B(n4792), .ZN(n4800) );
  AOI21_X1 U5350 ( .B1(n4795), .B2(n4914), .A(n4794), .ZN(n4798) );
  INV_X1 U5351 ( .A(n4833), .ZN(n4843) );
  AOI21_X1 U5352 ( .B1(n4798), .B2(n4797), .A(n4843), .ZN(n4796) );
  OAI21_X1 U5353 ( .B1(n4798), .B2(n4797), .A(n4796), .ZN(n4799) );
  OAI211_X1 U5354 ( .C1(n4838), .C2(n4914), .A(n4800), .B(n4799), .ZN(U3253)
         );
  AOI211_X1 U5355 ( .C1(n4803), .C2(n4802), .A(n4801), .B(n4839), .ZN(n4808)
         );
  AOI211_X1 U5356 ( .C1(n4806), .C2(n4805), .A(n4804), .B(n4843), .ZN(n4807)
         );
  AOI211_X1 U5357 ( .C1(n4848), .C2(n4809), .A(n4808), .B(n4807), .ZN(n4811)
         );
  OAI211_X1 U5358 ( .C1(n4812), .C2(n4853), .A(n4811), .B(n4810), .ZN(U3254)
         );
  INV_X1 U5359 ( .A(ADDR_REG_15__SCAN_IN), .ZN(n4823) );
  AOI211_X1 U5360 ( .C1(n4815), .C2(n4814), .A(n4813), .B(n4839), .ZN(n4820)
         );
  AOI211_X1 U5361 ( .C1(n4818), .C2(n4817), .A(n4816), .B(n4843), .ZN(n4819)
         );
  AOI211_X1 U5362 ( .C1(n4848), .C2(n4910), .A(n4820), .B(n4819), .ZN(n4822)
         );
  OAI211_X1 U5363 ( .C1(n4823), .C2(n4853), .A(n4822), .B(n4821), .ZN(U3255)
         );
  AOI21_X1 U5364 ( .B1(n4825), .B2(ADDR_REG_16__SCAN_IN), .A(n4824), .ZN(n4837) );
  OAI21_X1 U5365 ( .B1(n4828), .B2(n4827), .A(n4826), .ZN(n4834) );
  OAI21_X1 U5366 ( .B1(n4831), .B2(n4830), .A(n4829), .ZN(n4832) );
  AOI22_X1 U5367 ( .A1(n4835), .A2(n4834), .B1(n4833), .B2(n4832), .ZN(n4836)
         );
  OAI211_X1 U5368 ( .C1(n4909), .C2(n4838), .A(n4837), .B(n4836), .ZN(U3256)
         );
  AOI21_X1 U5369 ( .B1(n4841), .B2(n4840), .A(n4839), .ZN(n4850) );
  INV_X1 U5370 ( .A(n4842), .ZN(n4849) );
  OAI211_X1 U5371 ( .C1(n4854), .C2(n4853), .A(n4852), .B(n4851), .ZN(U3258)
         );
  XNOR2_X1 U5372 ( .A(n4855), .B(n4856), .ZN(n4973) );
  XNOR2_X1 U5373 ( .A(n4857), .B(n4856), .ZN(n4866) );
  OAI22_X1 U5374 ( .A1(n4860), .A2(n4878), .B1(n4859), .B2(n4858), .ZN(n4861)
         );
  AOI21_X1 U5375 ( .B1(n4863), .B2(n4862), .A(n4861), .ZN(n4864) );
  OAI21_X1 U5376 ( .B1(n4866), .B2(n4865), .A(n4864), .ZN(n4867) );
  AOI21_X1 U5377 ( .B1(n4973), .B2(n4877), .A(n4867), .ZN(n4975) );
  AOI22_X1 U5378 ( .A1(n4868), .A2(n4883), .B1(REG2_REG_11__SCAN_IN), .B2(
        n4888), .ZN(n4873) );
  AOI21_X1 U5379 ( .B1(n4870), .B2(n2269), .A(n4869), .ZN(n4970) );
  AOI22_X1 U5380 ( .A1(n4973), .A2(n4884), .B1(n4871), .B2(n4970), .ZN(n4872)
         );
  OAI211_X1 U5381 ( .C1(n4888), .C2(n4975), .A(n4873), .B(n4872), .ZN(U3279)
         );
  NOR2_X1 U5382 ( .A1(n4875), .A2(n4874), .ZN(n4927) );
  NOR2_X1 U5383 ( .A1(n4877), .A2(n4876), .ZN(n4880) );
  OAI22_X1 U5384 ( .A1(n4882), .A2(n4880), .B1(n4879), .B2(n4878), .ZN(n4926)
         );
  AOI21_X1 U5385 ( .B1(n4927), .B2(n4881), .A(n4926), .ZN(n4887) );
  INV_X1 U5386 ( .A(n4882), .ZN(n4928) );
  AOI22_X1 U5387 ( .A1(n4884), .A2(n4928), .B1(REG3_REG_0__SCAN_IN), .B2(n4883), .ZN(n4885) );
  OAI221_X1 U5388 ( .B1(n4888), .B2(n4887), .C1(n4530), .C2(n4886), .A(n4885), 
        .ZN(U3290) );
  AND2_X1 U5389 ( .A1(D_REG_31__SCAN_IN), .A2(n4903), .ZN(U3291) );
  AND2_X1 U5390 ( .A1(D_REG_30__SCAN_IN), .A2(n4903), .ZN(U3292) );
  AND2_X1 U5391 ( .A1(D_REG_29__SCAN_IN), .A2(n4903), .ZN(U3293) );
  NOR2_X1 U5392 ( .A1(n4902), .A2(n4889), .ZN(U3294) );
  AND2_X1 U5393 ( .A1(D_REG_27__SCAN_IN), .A2(n4903), .ZN(U3295) );
  NOR2_X1 U5394 ( .A1(n4902), .A2(n4890), .ZN(U3296) );
  NOR2_X1 U5395 ( .A1(n4902), .A2(n4891), .ZN(U3297) );
  NOR2_X1 U5396 ( .A1(n4902), .A2(n4892), .ZN(U3298) );
  NOR2_X1 U5397 ( .A1(n4902), .A2(n4893), .ZN(U3299) );
  NOR2_X1 U5398 ( .A1(n4902), .A2(n4894), .ZN(U3300) );
  NOR2_X1 U5399 ( .A1(n4902), .A2(n4895), .ZN(U3301) );
  NOR2_X1 U5400 ( .A1(n4902), .A2(n4896), .ZN(U3302) );
  AND2_X1 U5401 ( .A1(D_REG_19__SCAN_IN), .A2(n4903), .ZN(U3303) );
  NOR2_X1 U5402 ( .A1(n4902), .A2(n4897), .ZN(U3304) );
  AND2_X1 U5403 ( .A1(n4903), .A2(D_REG_17__SCAN_IN), .ZN(U3305) );
  NOR2_X1 U5404 ( .A1(n4902), .A2(n4898), .ZN(U3306) );
  AND2_X1 U5405 ( .A1(D_REG_15__SCAN_IN), .A2(n4903), .ZN(U3307) );
  AND2_X1 U5406 ( .A1(D_REG_14__SCAN_IN), .A2(n4903), .ZN(U3308) );
  AND2_X1 U5407 ( .A1(D_REG_13__SCAN_IN), .A2(n4903), .ZN(U3309) );
  AND2_X1 U5408 ( .A1(D_REG_12__SCAN_IN), .A2(n4903), .ZN(U3310) );
  AND2_X1 U5409 ( .A1(D_REG_11__SCAN_IN), .A2(n4903), .ZN(U3311) );
  AND2_X1 U5410 ( .A1(D_REG_10__SCAN_IN), .A2(n4903), .ZN(U3312) );
  AND2_X1 U5411 ( .A1(D_REG_9__SCAN_IN), .A2(n4903), .ZN(U3313) );
  AND2_X1 U5412 ( .A1(n4903), .A2(D_REG_8__SCAN_IN), .ZN(U3314) );
  NOR2_X1 U5413 ( .A1(n4902), .A2(n4899), .ZN(U3315) );
  NOR2_X1 U5414 ( .A1(n4902), .A2(n4900), .ZN(U3316) );
  AND2_X1 U5415 ( .A1(D_REG_5__SCAN_IN), .A2(n4903), .ZN(U3317) );
  NOR2_X1 U5416 ( .A1(n4902), .A2(n4901), .ZN(U3318) );
  AND2_X1 U5417 ( .A1(D_REG_3__SCAN_IN), .A2(n4903), .ZN(U3319) );
  AND2_X1 U5418 ( .A1(D_REG_2__SCAN_IN), .A2(n4903), .ZN(U3320) );
  OAI21_X1 U5419 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4904), .ZN(
        n4905) );
  INV_X1 U5420 ( .A(n4905), .ZN(U3329) );
  INV_X1 U5421 ( .A(DATAI_18_), .ZN(n4906) );
  AOI22_X1 U5422 ( .A1(STATE_REG_SCAN_IN), .A2(n4907), .B1(n4906), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5423 ( .A1(STATE_REG_SCAN_IN), .A2(n4909), .B1(n4908), .B2(U3149), 
        .ZN(U3336) );
  OAI22_X1 U5424 ( .A1(U3149), .A2(n4910), .B1(DATAI_15_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4911) );
  INV_X1 U5425 ( .A(n4911), .ZN(U3337) );
  AOI22_X1 U5426 ( .A1(STATE_REG_SCAN_IN), .A2(n2313), .B1(n4912), .B2(U3149), 
        .ZN(U3338) );
  AOI22_X1 U5427 ( .A1(STATE_REG_SCAN_IN), .A2(n4914), .B1(n4913), .B2(U3149), 
        .ZN(U3339) );
  INV_X1 U5428 ( .A(DATAI_12_), .ZN(n4915) );
  AOI22_X1 U5429 ( .A1(STATE_REG_SCAN_IN), .A2(n4916), .B1(n4915), .B2(U3149), 
        .ZN(U3340) );
  OAI22_X1 U5430 ( .A1(U3149), .A2(n4917), .B1(DATAI_10_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4918) );
  INV_X1 U5431 ( .A(n4918), .ZN(U3342) );
  AOI22_X1 U5432 ( .A1(STATE_REG_SCAN_IN), .A2(n4920), .B1(n4919), .B2(U3149), 
        .ZN(U3344) );
  INV_X1 U5433 ( .A(DATAI_7_), .ZN(n4921) );
  AOI22_X1 U5434 ( .A1(STATE_REG_SCAN_IN), .A2(n4922), .B1(n4921), .B2(U3149), 
        .ZN(U3345) );
  AOI22_X1 U5435 ( .A1(STATE_REG_SCAN_IN), .A2(n4924), .B1(n4923), .B2(U3149), 
        .ZN(U3346) );
  OAI22_X1 U5436 ( .A1(U3149), .A2(IR_REG_0__SCAN_IN), .B1(DATAI_0_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4925) );
  INV_X1 U5437 ( .A(n4925), .ZN(U3352) );
  AOI211_X1 U5438 ( .C1(n4972), .C2(n4928), .A(n4927), .B(n4926), .ZN(n4980)
         );
  INV_X1 U5439 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4929) );
  AOI22_X1 U5440 ( .A1(n4978), .A2(n4980), .B1(n4929), .B2(n4976), .ZN(U3467)
         );
  OAI22_X1 U5441 ( .A1(n4931), .A2(n4941), .B1(n4965), .B2(n4930), .ZN(n4932)
         );
  NOR2_X1 U5442 ( .A1(n4933), .A2(n4932), .ZN(n4981) );
  AOI22_X1 U5443 ( .A1(n4978), .A2(n4981), .B1(n4934), .B2(n4976), .ZN(U3469)
         );
  NOR3_X1 U5444 ( .A1(n4936), .A2(n4935), .A3(n4965), .ZN(n4938) );
  AOI211_X1 U5445 ( .C1(n4972), .C2(n4939), .A(n4938), .B(n4937), .ZN(n4982)
         );
  INV_X1 U5446 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4940) );
  AOI22_X1 U5447 ( .A1(n4978), .A2(n4982), .B1(n4940), .B2(n4976), .ZN(U3471)
         );
  NOR2_X1 U5448 ( .A1(n4942), .A2(n4941), .ZN(n4944) );
  AOI211_X1 U5449 ( .C1(n4971), .C2(n4945), .A(n4944), .B(n4943), .ZN(n4983)
         );
  INV_X1 U5450 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4946) );
  AOI22_X1 U5451 ( .A1(n4978), .A2(n4983), .B1(n4946), .B2(n4976), .ZN(U3473)
         );
  INV_X1 U5452 ( .A(n4947), .ZN(n4949) );
  AOI211_X1 U5453 ( .C1(n4950), .C2(n4972), .A(n4949), .B(n4948), .ZN(n4984)
         );
  AOI22_X1 U5454 ( .A1(n4978), .A2(n4984), .B1(n4951), .B2(n4976), .ZN(U3475)
         );
  NOR2_X1 U5455 ( .A1(n4953), .A2(n4952), .ZN(n4954) );
  AOI211_X1 U5456 ( .C1(n4971), .C2(n4956), .A(n4955), .B(n4954), .ZN(n4985)
         );
  INV_X1 U5457 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4957) );
  AOI22_X1 U5458 ( .A1(n4978), .A2(n4985), .B1(n4957), .B2(n4976), .ZN(U3477)
         );
  NAND2_X1 U5459 ( .A1(n4958), .A2(n4968), .ZN(n4960) );
  AND3_X1 U5460 ( .A1(n4961), .A2(n4960), .A3(n4959), .ZN(n4986) );
  INV_X1 U5461 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4962) );
  AOI22_X1 U5462 ( .A1(n4978), .A2(n4986), .B1(n4962), .B2(n4976), .ZN(U3481)
         );
  OAI21_X1 U5463 ( .B1(n4965), .B2(n4964), .A(n4963), .ZN(n4966) );
  AOI21_X1 U5464 ( .B1(n4968), .B2(n4967), .A(n4966), .ZN(n4987) );
  AOI22_X1 U5465 ( .A1(n4978), .A2(n4987), .B1(n4969), .B2(n4976), .ZN(U3485)
         );
  AOI22_X1 U5466 ( .A1(n4973), .A2(n4972), .B1(n4971), .B2(n4970), .ZN(n4974)
         );
  AND2_X1 U5467 ( .A1(n4975), .A2(n4974), .ZN(n4989) );
  AOI22_X1 U5468 ( .A1(n4978), .A2(n4989), .B1(n4977), .B2(n4976), .ZN(U3489)
         );
  AOI22_X1 U5469 ( .A1(n4990), .A2(n4980), .B1(n4979), .B2(n4988), .ZN(U3518)
         );
  AOI22_X1 U5470 ( .A1(n4990), .A2(n4981), .B1(n3116), .B2(n4988), .ZN(U3519)
         );
  AOI22_X1 U5471 ( .A1(n4990), .A2(n4982), .B1(n3119), .B2(n4988), .ZN(U3520)
         );
  AOI22_X1 U5472 ( .A1(n4990), .A2(n4983), .B1(n2483), .B2(n4988), .ZN(U3521)
         );
  AOI22_X1 U5473 ( .A1(n4990), .A2(n4984), .B1(n3125), .B2(n4988), .ZN(U3522)
         );
  AOI22_X1 U5474 ( .A1(n4990), .A2(n4985), .B1(n3114), .B2(n4988), .ZN(U3523)
         );
  AOI22_X1 U5475 ( .A1(n4990), .A2(n4986), .B1(n2550), .B2(n4988), .ZN(U3525)
         );
  AOI22_X1 U5476 ( .A1(n4990), .A2(n4987), .B1(n2585), .B2(n4988), .ZN(U3527)
         );
  AOI22_X1 U5477 ( .A1(n4990), .A2(n4989), .B1(n3395), .B2(n4988), .ZN(U3529)
         );
  NOR2_X1 U2490 ( .A1(n2470), .A2(n2469), .ZN(n2472) );
  AND2_X1 U2952 ( .A1(n2413), .A2(n2296), .ZN(n2392) );
  CLKBUF_X1 U2482 ( .A(n2504), .Z(n2943) );
  CLKBUF_X1 U2485 ( .A(n2465), .Z(n3487) );
  CLKBUF_X1 U3039 ( .A(n3858), .Z(n3949) );
endmodule

