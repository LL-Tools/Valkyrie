

module b21_C_gen_AntiSAT_k_256_7 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2, 
        keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7, 
        keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12, 
        keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17, 
        keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22, 
        keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27, 
        keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32, 
        keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37, 
        keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42, 
        keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47, 
        keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52, 
        keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57, 
        keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62, 
        keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67, 
        keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72, 
        keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77, 
        keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82, 
        keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87, 
        keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92, 
        keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97, 
        keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515;

  INV_X4 U4982 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  OAI21_X1 U4983 ( .B1(n5687), .B2(n4947), .A(n5712), .ZN(n4943) );
  AND3_X1 U4984 ( .A1(n6006), .A2(n6005), .A3(n6004), .ZN(n9839) );
  CLKBUF_X2 U4985 ( .A(n5148), .Z(n5772) );
  INV_X4 U4986 ( .A(n5148), .ZN(n5137) );
  NAND2_X1 U4987 ( .A1(n4940), .A2(n4939), .ZN(n7839) );
  INV_X1 U4988 ( .A(n5199), .ZN(n7823) );
  INV_X1 U4989 ( .A(n5915), .ZN(n8754) );
  NAND2_X1 U4990 ( .A1(n9617), .A2(n7832), .ZN(n6018) );
  NAND2_X1 U4991 ( .A1(n5921), .A2(n4578), .ZN(n6680) );
  AOI22_X1 U4992 ( .A1(n4536), .A2(P1_IR_REG_0__SCAN_IN), .B1(n4579), .B2(
        n5860), .ZN(n4578) );
  INV_X2 U4993 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5860) );
  INV_X1 U4994 ( .A(n7984), .ZN(n7976) );
  INV_X1 U4995 ( .A(n6556), .ZN(n5568) );
  NAND2_X1 U4996 ( .A1(n6556), .A2(n7832), .ZN(n5196) );
  INV_X1 U4997 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5807) );
  INV_X2 U4998 ( .A(n6345), .ZN(n7773) );
  INV_X1 U4999 ( .A(n7304), .ZN(n7776) );
  INV_X2 U5000 ( .A(n7839), .ZN(n5771) );
  INV_X1 U5001 ( .A(n5579), .ZN(n5822) );
  NAND2_X2 U5002 ( .A1(n8243), .A2(n5818), .ZN(n6556) );
  NAND2_X2 U5003 ( .A1(n6450), .A2(n9613), .ZN(n9617) );
  BUF_X1 U5004 ( .A(n5991), .Z(n4478) );
  NAND2_X1 U5005 ( .A1(n8899), .A2(n8896), .ZN(n9771) );
  AND3_X1 U5006 ( .A1(n5942), .A2(n5941), .A3(n5940), .ZN(n9819) );
  OR2_X1 U5007 ( .A1(n5861), .A2(n5860), .ZN(n5862) );
  INV_X1 U5008 ( .A(n5576), .ZN(n7827) );
  NAND2_X1 U5009 ( .A1(n5325), .A2(n5324), .ZN(n10014) );
  NAND2_X1 U5010 ( .A1(n4497), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5778) );
  INV_X2 U5011 ( .A(n6492), .ZN(n7832) );
  AND2_X1 U5012 ( .A1(n6461), .A2(n6460), .ZN(n9356) );
  OAI21_X1 U5013 ( .B1(n9243), .B2(n9244), .A(n9088), .ZN(n9228) );
  INV_X2 U5014 ( .A(n6018), .ZN(n6048) );
  NAND2_X1 U5015 ( .A1(n9497), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5859) );
  NAND2_X1 U5016 ( .A1(n4795), .A2(n4793), .ZN(n9506) );
  XNOR2_X1 U5017 ( .A(n5894), .B(n5893), .ZN(n6450) );
  OAI21_X2 U5018 ( .B1(n5117), .B2(n8020), .A(n6946), .ZN(n5148) );
  AND3_X2 U5019 ( .A1(n4720), .A2(n4719), .A3(n4607), .ZN(n5878) );
  XNOR2_X2 U5020 ( .A(n5859), .B(n9498), .ZN(n5865) );
  AOI21_X2 U5021 ( .B1(n8203), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8202), .ZN(
        n8206) );
  NAND2_X1 U5022 ( .A1(n9726), .A2(n7314), .ZN(n7360) );
  AOI21_X2 U5023 ( .B1(n9104), .B2(n9103), .A(n9102), .ZN(n9311) );
  AOI21_X2 U5024 ( .B1(n5219), .B2(n5218), .A(n5217), .ZN(n5244) );
  AOI211_X2 U5025 ( .C1(n9012), .C2(n9011), .A(n9013), .B(n9010), .ZN(n9015)
         );
  OAI22_X2 U5026 ( .A1(n8106), .A2(n8107), .B1(n5606), .B2(n5605), .ZN(n8072)
         );
  OAI21_X2 U5027 ( .B1(n8126), .B2(n4957), .A(n4954), .ZN(n8106) );
  NOR2_X2 U5028 ( .A1(n7186), .A2(n10014), .ZN(n7185) );
  NAND2_X1 U5029 ( .A1(n5737), .A2(n5736), .ZN(n8037) );
  MUX2_X1 U5030 ( .A(n9460), .B(n9459), .S(n9888), .Z(n9461) );
  AND2_X1 U5031 ( .A1(n9140), .A2(n9139), .ZN(n9349) );
  AND2_X1 U5032 ( .A1(n4999), .A2(n6367), .ZN(n8637) );
  OR2_X1 U5033 ( .A1(n7990), .A2(n8022), .ZN(n8026) );
  AND2_X1 U5034 ( .A1(n4712), .A2(n4612), .ZN(n8622) );
  XNOR2_X1 U5035 ( .A(n4841), .B(n4563), .ZN(n9503) );
  NAND2_X1 U5036 ( .A1(n7772), .A2(n7771), .ZN(n9352) );
  OR2_X1 U5037 ( .A1(n9162), .A2(n9172), .ZN(n9096) );
  NAND2_X1 U5038 ( .A1(n5514), .A2(n5513), .ZN(n8090) );
  NAND2_X1 U5039 ( .A1(n6384), .A2(n6383), .ZN(n9364) );
  NAND2_X1 U5040 ( .A1(n5636), .A2(n5635), .ZN(n8546) );
  NAND2_X1 U5041 ( .A1(n6308), .A2(n6307), .ZN(n9400) );
  NAND2_X1 U5042 ( .A1(n5043), .A2(n5041), .ZN(n7755) );
  OAI21_X1 U5043 ( .B1(n7507), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7506), .ZN(
        n7738) );
  AND2_X1 U5044 ( .A1(n6408), .A2(n6407), .ZN(n9172) );
  NAND2_X1 U5045 ( .A1(n6823), .A2(n5241), .ZN(n6833) );
  OR2_X1 U5046 ( .A1(n7333), .A2(n8961), .ZN(n9731) );
  AOI21_X1 U5047 ( .B1(n4937), .B2(n4935), .A(n4510), .ZN(n4934) );
  NAND2_X1 U5048 ( .A1(n4886), .A2(n4885), .ZN(n7059) );
  XNOR2_X1 U5049 ( .A(n4698), .B(n4553), .ZN(n6535) );
  NAND2_X1 U5050 ( .A1(n9035), .A2(n9831), .ZN(n8896) );
  OR2_X1 U5051 ( .A1(n5317), .A2(n5316), .ZN(n5347) );
  NAND2_X1 U5052 ( .A1(n5292), .A2(n5291), .ZN(n5317) );
  AND3_X1 U5053 ( .A1(n5978), .A2(n5977), .A3(n5976), .ZN(n9831) );
  AND2_X1 U5054 ( .A1(n5225), .A2(n5224), .ZN(n9989) );
  NAND2_X1 U5055 ( .A1(n4634), .A2(n5198), .ZN(n9922) );
  INV_X1 U5056 ( .A(n9825), .ZN(n7251) );
  AND3_X1 U5057 ( .A1(n5964), .A2(n5963), .A3(n5962), .ZN(n9825) );
  NAND4_X2 U5058 ( .A1(n5999), .A2(n5998), .A3(n5997), .A4(n5996), .ZN(n9844)
         );
  INV_X1 U5059 ( .A(n4478), .ZN(n8750) );
  NOR2_X1 U5060 ( .A1(n7716), .A2(n9963), .ZN(n9945) );
  INV_X1 U5061 ( .A(n5993), .ZN(n6537) );
  CLKBUF_X1 U5062 ( .A(n5929), .Z(n7784) );
  BUF_X2 U5063 ( .A(n5196), .Z(n5221) );
  AND4_X1 U5064 ( .A1(n5102), .A2(n5101), .A3(n5100), .A4(n5099), .ZN(n7804)
         );
  CLKBUF_X3 U5065 ( .A(n8754), .Z(n4479) );
  NAND2_X2 U5066 ( .A1(n9617), .A2(n4876), .ZN(n8855) );
  NAND2_X1 U5067 ( .A1(n6443), .A2(n7135), .ZN(n6345) );
  NAND2_X1 U5068 ( .A1(n5184), .A2(n5183), .ZN(n5189) );
  AND2_X1 U5069 ( .A1(n8030), .A2(n8356), .ZN(n8020) );
  NAND2_X1 U5070 ( .A1(n5827), .A2(n7840), .ZN(n7984) );
  AOI21_X1 U5071 ( .B1(n6600), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6599), .ZN(
        n6602) );
  OR2_X1 U5072 ( .A1(n9013), .A2(n4721), .ZN(n7135) );
  XNOR2_X1 U5073 ( .A(n5900), .B(n5899), .ZN(n9013) );
  INV_X1 U5074 ( .A(n5864), .ZN(n5869) );
  BUF_X1 U5075 ( .A(n6450), .Z(n4480) );
  NAND2_X1 U5076 ( .A1(n4630), .A2(n4745), .ZN(n8243) );
  NAND2_X1 U5077 ( .A1(n5006), .A2(n8610), .ZN(n5199) );
  OR2_X2 U5078 ( .A1(n8606), .A2(n8610), .ZN(n5726) );
  AND2_X1 U5079 ( .A1(n9525), .A2(n4786), .ZN(n9523) );
  NAND2_X1 U5080 ( .A1(n4835), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5891) );
  NAND2_X1 U5081 ( .A1(n5892), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U5082 ( .A1(n5889), .A2(n5133), .ZN(n5161) );
  OR2_X1 U5083 ( .A1(n9511), .A2(n6570), .ZN(n9525) );
  NAND2_X1 U5084 ( .A1(n5121), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4629) );
  INV_X2 U5085 ( .A(n9502), .ZN(n8036) );
  INV_X1 U5086 ( .A(n6492), .ZN(n4877) );
  AND2_X1 U5087 ( .A1(n5078), .A2(n5880), .ZN(n5077) );
  OR2_X1 U5088 ( .A1(n5854), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n5855) );
  AND4_X1 U5089 ( .A1(n5844), .A2(n5843), .A3(n5842), .A4(n5841), .ZN(n5847)
         );
  AND2_X1 U5090 ( .A1(n5849), .A2(n5848), .ZN(n5907) );
  NOR2_X2 U5091 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5920) );
  INV_X1 U5092 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5112) );
  INV_X1 U5093 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5103) );
  NOR2_X1 U5094 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5087) );
  NOR2_X1 U5095 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5088) );
  INV_X1 U5096 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5475) );
  INV_X1 U5097 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5442) );
  INV_X1 U5098 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5445) );
  NOR2_X1 U5099 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5842) );
  INV_X1 U5100 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5902) );
  NOR2_X1 U5101 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5843) );
  INV_X1 U5102 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5899) );
  NOR2_X1 U5103 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5849) );
  NOR2_X1 U5104 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5852) );
  NOR2_X2 U5105 ( .A1(n8485), .A2(n8568), .ZN(n8471) );
  NOR2_X2 U5106 ( .A1(n4882), .A2(n7658), .ZN(n7653) );
  OAI22_X2 U5107 ( .A1(n7755), .A2(n7609), .B1(n7762), .B2(n9568), .ZN(n7671)
         );
  NOR2_X2 U5108 ( .A1(n8354), .A2(n8523), .ZN(n8339) );
  NOR2_X2 U5109 ( .A1(n8382), .A2(n8533), .ZN(n4888) );
  OAI222_X1 U5110 ( .A1(n7729), .A2(n7705), .B1(P2_U3152), .B2(n5818), .C1(
        n8612), .C2(n8035), .ZN(P2_U3330) );
  NAND2_X1 U5111 ( .A1(n4862), .A2(n4861), .ZN(n7725) );
  AOI21_X1 U5112 ( .B1(n4864), .B2(n4866), .A(n4562), .ZN(n4861) );
  NAND2_X1 U5113 ( .A1(n5758), .A2(n4864), .ZN(n4862) );
  NOR2_X1 U5114 ( .A1(n7841), .A2(n4685), .ZN(n4684) );
  AND2_X1 U5115 ( .A1(n9437), .A2(n9442), .ZN(n9102) );
  NAND2_X1 U5116 ( .A1(n5294), .A2(n5293), .ZN(n5343) );
  NAND2_X1 U5117 ( .A1(n8857), .A2(n8856), .ZN(n9126) );
  NAND2_X1 U5118 ( .A1(n4738), .A2(n7934), .ZN(n7941) );
  OAI21_X1 U5119 ( .B1(n4742), .B2(n4739), .A(n7933), .ZN(n4738) );
  NOR2_X1 U5120 ( .A1(n6877), .A2(n4938), .ZN(n4937) );
  INV_X1 U5121 ( .A(n5265), .ZN(n4938) );
  AND2_X1 U5122 ( .A1(n8503), .A2(n4682), .ZN(n4681) );
  NAND2_X1 U5123 ( .A1(n4683), .A2(n7977), .ZN(n4682) );
  OR2_X1 U5124 ( .A1(n8511), .A2(n8257), .ZN(n7819) );
  OR2_X1 U5125 ( .A1(n8533), .A2(n8149), .ZN(n7961) );
  INV_X1 U5126 ( .A(n8272), .ZN(n4913) );
  OR2_X1 U5127 ( .A1(n8571), .A2(n8130), .ZN(n7848) );
  NOR2_X1 U5128 ( .A1(n7534), .A2(n7424), .ZN(n4881) );
  AND2_X1 U5129 ( .A1(n4621), .A2(n4618), .ZN(n4617) );
  NAND2_X1 U5130 ( .A1(n4586), .A2(n4589), .ZN(n4584) );
  AND2_X1 U5131 ( .A1(n9150), .A2(n4810), .ZN(n4809) );
  NAND2_X1 U5132 ( .A1(n9192), .A2(n9204), .ZN(n8948) );
  INV_X1 U5133 ( .A(n5069), .ZN(n5068) );
  OAI21_X1 U5134 ( .B1(n5070), .B2(n9244), .A(n9109), .ZN(n5069) );
  OR2_X1 U5135 ( .A1(n9239), .A2(n9254), .ZN(n9109) );
  INV_X1 U5136 ( .A(n4871), .ZN(n4870) );
  OAI21_X1 U5137 ( .B1(n4874), .B2(n4550), .A(n5713), .ZN(n4871) );
  NAND2_X1 U5138 ( .A1(n5672), .A2(n5671), .ZN(n5674) );
  OAI21_X1 U5139 ( .B1(n5591), .B2(n5590), .A(n5589), .ZN(n5608) );
  NAND2_X1 U5140 ( .A1(n4858), .A2(n5466), .ZN(n4857) );
  INV_X1 U5141 ( .A(n5491), .ZN(n4858) );
  XNOR2_X1 U5142 ( .A(n5465), .B(n10223), .ZN(n5464) );
  NAND2_X1 U5143 ( .A1(n5343), .A2(n5296), .ZN(n5316) );
  AND2_X2 U5144 ( .A1(n8606), .A2(n8610), .ZN(n5576) );
  AND2_X1 U5145 ( .A1(n4953), .A2(n4503), .ZN(n4951) );
  OR2_X1 U5146 ( .A1(n5403), .A2(n10394), .ZN(n5429) );
  AOI21_X1 U5147 ( .B1(n4684), .B2(n4683), .A(n4564), .ZN(n4679) );
  NAND2_X1 U5148 ( .A1(n8606), .A2(n5098), .ZN(n5579) );
  NAND2_X1 U5149 ( .A1(n7821), .A2(n7820), .ZN(n8288) );
  NAND2_X1 U5150 ( .A1(n4891), .A2(n4890), .ZN(n8330) );
  AOI21_X1 U5151 ( .B1(n4486), .B2(n4895), .A(n4525), .ZN(n4890) );
  OR2_X1 U5152 ( .A1(n8554), .A2(n8151), .ZN(n7948) );
  OR2_X1 U5153 ( .A1(n7658), .A2(n8093), .ZN(n7927) );
  AND2_X1 U5154 ( .A1(n4628), .A2(n4917), .ZN(n7426) );
  NAND2_X1 U5155 ( .A1(n7269), .A2(n4916), .ZN(n4628) );
  NAND2_X1 U5156 ( .A1(n4924), .A2(n4484), .ZN(n4917) );
  AND2_X1 U5157 ( .A1(n4926), .A2(n4918), .ZN(n4916) );
  OR2_X1 U5158 ( .A1(n5356), .A2(n6957), .ZN(n5376) );
  OR2_X1 U5159 ( .A1(n7269), .A2(n7105), .ZN(n4922) );
  INV_X1 U5160 ( .A(n7992), .ZN(n8284) );
  NAND2_X1 U5161 ( .A1(n8649), .A2(n8644), .ZN(n8658) );
  AOI21_X1 U5162 ( .B1(n4705), .B2(n4597), .A(n4596), .ZN(n4595) );
  INV_X1 U5163 ( .A(n7521), .ZN(n4596) );
  INV_X1 U5164 ( .A(n4599), .ZN(n4597) );
  INV_X1 U5165 ( .A(n4705), .ZN(n4598) );
  INV_X2 U5166 ( .A(n6537), .ZN(n8751) );
  NOR2_X1 U5167 ( .A1(n7028), .A2(n7027), .ZN(n7227) );
  OR2_X1 U5168 ( .A1(n7229), .A2(n7611), .ZN(n4572) );
  OR2_X1 U5169 ( .A1(n9159), .A2(n9352), .ZN(n9143) );
  OR2_X1 U5170 ( .A1(n9192), .A2(n9204), .ZN(n9167) );
  NOR2_X1 U5171 ( .A1(n9406), .A2(n9106), .ZN(n9107) );
  AND2_X1 U5172 ( .A1(n9406), .A2(n9106), .ZN(n5062) );
  INV_X1 U5173 ( .A(n9415), .ZN(n9265) );
  NAND2_X1 U5174 ( .A1(n7672), .A2(n9441), .ZN(n5052) );
  NOR2_X1 U5175 ( .A1(n7672), .A2(n9441), .ZN(n5051) );
  INV_X1 U5176 ( .A(n8855), .ZN(n6276) );
  AND2_X1 U5177 ( .A1(n5077), .A2(n5893), .ZN(n4668) );
  NOR2_X1 U5178 ( .A1(n5855), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4607) );
  OR2_X1 U5179 ( .A1(n6514), .A2(n5818), .ZN(n8426) );
  OAI21_X1 U5180 ( .B1(n8238), .B2(n9907), .A(n4791), .ZN(n4790) );
  AOI21_X1 U5181 ( .B1(n8239), .B2(n9904), .A(n9527), .ZN(n4791) );
  INV_X1 U5182 ( .A(n9617), .ZN(n6485) );
  AOI21_X1 U5183 ( .B1(n5074), .B2(n9150), .A(n4538), .ZN(n5073) );
  INV_X1 U5184 ( .A(n7881), .ZN(n4735) );
  NOR2_X1 U5185 ( .A1(n4731), .A2(n7111), .ZN(n4730) );
  INV_X1 U5186 ( .A(n7927), .ZN(n4741) );
  OAI211_X1 U5187 ( .C1(n7913), .C2(n7976), .A(n4749), .B(n8008), .ZN(n7926)
         );
  INV_X1 U5188 ( .A(n4750), .ZN(n4749) );
  NAND2_X1 U5189 ( .A1(n4659), .A2(n4658), .ZN(n4657) );
  AOI21_X1 U5190 ( .B1(n8783), .B2(n8864), .A(n8807), .ZN(n4658) );
  NAND2_X1 U5191 ( .A1(n4661), .A2(n4660), .ZN(n4659) );
  AOI21_X1 U5192 ( .B1(n7935), .B2(n7944), .A(n4727), .ZN(n4726) );
  NAND2_X1 U5193 ( .A1(n7948), .A2(n7942), .ZN(n4727) );
  NAND2_X1 U5194 ( .A1(n7939), .A2(n4517), .ZN(n4753) );
  AOI21_X1 U5195 ( .B1(n8388), .B2(n8273), .A(n7984), .ZN(n4754) );
  NAND2_X1 U5196 ( .A1(n4640), .A2(n4641), .ZN(n8825) );
  AOI21_X1 U5197 ( .B1(n8923), .B2(n4643), .A(n4642), .ZN(n4641) );
  MUX2_X1 U5198 ( .A(n8832), .B(n8831), .S(n8864), .Z(n8833) );
  AOI21_X1 U5199 ( .B1(n8827), .B2(n8865), .A(n8835), .ZN(n4665) );
  OAI22_X1 U5200 ( .A1(n8845), .A2(n9364), .B1(n8864), .B2(n8948), .ZN(n4663)
         );
  INV_X1 U5201 ( .A(n7849), .ZN(n7860) );
  INV_X1 U5202 ( .A(n6156), .ZN(n4993) );
  INV_X1 U5203 ( .A(n7603), .ZN(n5047) );
  NAND2_X1 U5204 ( .A1(n5391), .A2(n10363), .ZN(n5417) );
  NOR2_X1 U5205 ( .A1(n5345), .A2(n4553), .ZN(n4850) );
  NAND2_X1 U5206 ( .A1(n5349), .A2(n5348), .ZN(n5367) );
  OAI21_X1 U5207 ( .B1(n7832), .B2(n5192), .A(n5191), .ZN(n5211) );
  NAND2_X1 U5208 ( .A1(n4877), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5191) );
  NAND2_X1 U5209 ( .A1(n7446), .A2(n5416), .ZN(n4972) );
  AND2_X1 U5210 ( .A1(n7819), .A2(n7818), .ZN(n7993) );
  NOR2_X1 U5211 ( .A1(n7914), .A2(n7416), .ZN(n4692) );
  INV_X1 U5212 ( .A(n8004), .ZN(n7105) );
  NOR2_X1 U5213 ( .A1(n4481), .A2(n6945), .ZN(n4615) );
  NAND2_X1 U5214 ( .A1(n9922), .A2(n4755), .ZN(n7849) );
  OR2_X1 U5215 ( .A1(n5726), .A2(n10365), .ZN(n5153) );
  NAND2_X1 U5216 ( .A1(n7426), .A2(n7425), .ZN(n7427) );
  NOR2_X1 U5217 ( .A1(n7860), .A2(n5014), .ZN(n5021) );
  INV_X1 U5218 ( .A(n5021), .ZN(n5017) );
  NOR2_X1 U5219 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5083) );
  AND2_X1 U5220 ( .A1(n4980), .A2(n6036), .ZN(n4979) );
  INV_X1 U5221 ( .A(n7194), .ZN(n6036) );
  NAND2_X1 U5222 ( .A1(n6031), .A2(n4507), .ZN(n4980) );
  NAND2_X1 U5223 ( .A1(n6841), .A2(n5989), .ZN(n7092) );
  OR2_X1 U5224 ( .A1(n6348), .A2(n6347), .ZN(n4604) );
  INV_X1 U5225 ( .A(n7436), .ZN(n4709) );
  AND2_X1 U5226 ( .A1(n6104), .A2(n6079), .ZN(n4994) );
  AND2_X1 U5227 ( .A1(n9012), .A2(n4670), .ZN(n4669) );
  INV_X1 U5228 ( .A(n4671), .ZN(n4670) );
  OAI22_X1 U5229 ( .A1(n9341), .A2(n8865), .B1(n9347), .B2(n8864), .ZN(n4671)
         );
  NAND2_X1 U5230 ( .A1(n9341), .A2(n9347), .ZN(n4672) );
  INV_X1 U5231 ( .A(n5865), .ZN(n5870) );
  OR2_X1 U5232 ( .A1(n5929), .A2(n5863), .ZN(n5868) );
  NAND2_X1 U5233 ( .A1(n4807), .A2(n8873), .ZN(n4806) );
  NAND2_X1 U5234 ( .A1(n9137), .A2(n4808), .ZN(n4807) );
  INV_X1 U5235 ( .A(n9096), .ZN(n4808) );
  NOR2_X1 U5236 ( .A1(n4806), .A2(n4805), .ZN(n4804) );
  INV_X1 U5237 ( .A(n9095), .ZN(n4805) );
  NAND2_X1 U5238 ( .A1(n9162), .A2(n9172), .ZN(n8875) );
  AND2_X1 U5239 ( .A1(n9364), .A2(n9153), .ZN(n9094) );
  AND2_X1 U5240 ( .A1(n8948), .A2(n9182), .ZN(n9093) );
  OR2_X1 U5241 ( .A1(n9364), .A2(n9186), .ZN(n9119) );
  NOR2_X1 U5242 ( .A1(n9400), .A2(n9239), .ZN(n4767) );
  NOR2_X1 U5243 ( .A1(n9303), .A2(n9307), .ZN(n9281) );
  OR2_X1 U5244 ( .A1(n9307), .A2(n9424), .ZN(n8953) );
  OR2_X1 U5245 ( .A1(n9437), .A2(n9423), .ZN(n9075) );
  AND2_X1 U5246 ( .A1(n9592), .A2(n7607), .ZN(n7608) );
  NOR2_X1 U5247 ( .A1(n7608), .A2(n7472), .ZN(n5044) );
  AND2_X1 U5248 ( .A1(n5048), .A2(n5047), .ZN(n9561) );
  NAND2_X1 U5249 ( .A1(n7605), .A2(n7604), .ZN(n5048) );
  NOR2_X1 U5250 ( .A1(n7469), .A2(n4760), .ZN(n4759) );
  NAND2_X1 U5251 ( .A1(n7527), .A2(n4761), .ZN(n4760) );
  INV_X1 U5252 ( .A(n9744), .ZN(n4762) );
  NAND2_X1 U5253 ( .A1(n8997), .A2(n4816), .ZN(n4815) );
  NAND2_X1 U5254 ( .A1(n7316), .A2(n8896), .ZN(n4816) );
  OR2_X1 U5255 ( .A1(n9843), .A2(n9861), .ZN(n9730) );
  NAND2_X1 U5256 ( .A1(n8760), .A2(n7397), .ZN(n8962) );
  XNOR2_X1 U5257 ( .A(n9794), .B(n9813), .ZN(n7124) );
  NAND2_X1 U5258 ( .A1(n4800), .A2(n9799), .ZN(n4801) );
  INV_X1 U5259 ( .A(n8886), .ZN(n4800) );
  NOR2_X1 U5260 ( .A1(n9364), .A2(n9190), .ZN(n9173) );
  OAI21_X1 U5261 ( .B1(n7725), .B2(n7724), .A(n7723), .ZN(n7831) );
  AOI21_X1 U5262 ( .B1(n4855), .B2(n4857), .A(n4852), .ZN(n4851) );
  INV_X1 U5263 ( .A(n4856), .ZN(n4855) );
  OAI21_X1 U5264 ( .B1(n4859), .B2(n4857), .A(n5490), .ZN(n4856) );
  NOR2_X1 U5265 ( .A1(n5467), .A2(n4860), .ZN(n4859) );
  INV_X1 U5266 ( .A(n5464), .ZN(n5467) );
  INV_X1 U5267 ( .A(n5440), .ZN(n4860) );
  NAND2_X1 U5268 ( .A1(n5490), .A2(n5472), .ZN(n5491) );
  NAND2_X1 U5269 ( .A1(n5439), .A2(n5080), .ZN(n5441) );
  OAI21_X1 U5270 ( .B1(n5419), .B2(n5418), .A(n5417), .ZN(n5439) );
  AOI21_X1 U5271 ( .B1(n4850), .B2(n4848), .A(n4847), .ZN(n4846) );
  INV_X1 U5272 ( .A(n5367), .ZN(n4847) );
  INV_X1 U5273 ( .A(n5346), .ZN(n4848) );
  INV_X1 U5274 ( .A(n4850), .ZN(n4849) );
  AND2_X1 U5275 ( .A1(n5343), .A2(n5342), .ZN(n5346) );
  XNOR2_X1 U5276 ( .A(n5290), .B(SI_7_), .ZN(n5287) );
  AOI21_X1 U5277 ( .B1(n5267), .B2(n4839), .A(n4529), .ZN(n4838) );
  XNOR2_X1 U5278 ( .A(n5211), .B(SI_4_), .ZN(n5213) );
  OR2_X1 U5279 ( .A1(n5549), .A2(n5548), .ZN(n5574) );
  NAND2_X1 U5280 ( .A1(n5572), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5597) );
  INV_X1 U5281 ( .A(n5574), .ZN(n5572) );
  NAND2_X1 U5282 ( .A1(n8126), .A2(n8125), .ZN(n4960) );
  INV_X1 U5283 ( .A(n4937), .ZN(n4936) );
  INV_X1 U5284 ( .A(n6834), .ZN(n4935) );
  NAND2_X1 U5285 ( .A1(n5327), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5356) );
  INV_X1 U5286 ( .A(n5329), .ZN(n5327) );
  INV_X1 U5287 ( .A(n4958), .ZN(n4957) );
  AOI21_X1 U5288 ( .B1(n4958), .B2(n4956), .A(n4955), .ZN(n4954) );
  INV_X1 U5289 ( .A(n5588), .ZN(n4955) );
  NAND2_X1 U5290 ( .A1(n4966), .A2(n5341), .ZN(n4965) );
  INV_X1 U5291 ( .A(n8053), .ZN(n4966) );
  INV_X1 U5292 ( .A(n4965), .ZN(n4961) );
  NOR2_X1 U5293 ( .A1(n7623), .A2(n4969), .ZN(n4968) );
  INV_X1 U5294 ( .A(n5518), .ZN(n4969) );
  INV_X1 U5295 ( .A(n8078), .ZN(n4947) );
  INV_X1 U5296 ( .A(n8099), .ZN(n4948) );
  OR2_X1 U5297 ( .A1(n8321), .A2(n8511), .ZN(n8304) );
  XNOR2_X1 U5298 ( .A(n8281), .B(n8280), .ZN(n8313) );
  OR2_X1 U5299 ( .A1(n8529), .A2(n8370), .ZN(n7842) );
  XNOR2_X1 U5300 ( .A(n8523), .B(n8278), .ZN(n8333) );
  NAND2_X1 U5301 ( .A1(n4894), .A2(n8276), .ZN(n4893) );
  INV_X1 U5302 ( .A(n8276), .ZN(n4895) );
  AND2_X1 U5303 ( .A1(n7842), .A2(n7843), .ZN(n8348) );
  NOR2_X1 U5304 ( .A1(n4637), .A2(n4636), .ZN(n8275) );
  INV_X1 U5305 ( .A(n8274), .ZN(n4636) );
  INV_X1 U5306 ( .A(n8389), .ZN(n4637) );
  AOI21_X1 U5307 ( .B1(n4912), .B2(n4911), .A(n4915), .ZN(n4910) );
  NOR2_X1 U5308 ( .A1(n8546), .A2(n8410), .ZN(n4915) );
  INV_X1 U5309 ( .A(n8270), .ZN(n4911) );
  NAND2_X1 U5310 ( .A1(n4909), .A2(n4912), .ZN(n4908) );
  AND2_X1 U5311 ( .A1(n5620), .A2(n5619), .ZN(n8429) );
  NAND2_X1 U5312 ( .A1(n5009), .A2(n4697), .ZN(n8431) );
  AND2_X1 U5313 ( .A1(n5007), .A2(n7817), .ZN(n4697) );
  NAND2_X1 U5314 ( .A1(n8471), .A2(n8454), .ZN(n8450) );
  OR2_X1 U5315 ( .A1(n8568), .A2(n8152), .ZN(n8445) );
  NAND2_X1 U5316 ( .A1(n4906), .A2(n4905), .ZN(n8463) );
  AOI21_X1 U5317 ( .B1(n4485), .B2(n8262), .A(n4526), .ZN(n4905) );
  NAND2_X1 U5318 ( .A1(n7561), .A2(n4689), .ZN(n4688) );
  NOR2_X1 U5319 ( .A1(n5005), .A2(n4690), .ZN(n4689) );
  NAND2_X1 U5320 ( .A1(n8262), .A2(n7927), .ZN(n5005) );
  NAND2_X1 U5321 ( .A1(n5004), .A2(n7927), .ZN(n5003) );
  NAND2_X1 U5322 ( .A1(n7378), .A2(n4491), .ZN(n4882) );
  NAND2_X1 U5323 ( .A1(n7561), .A2(n7915), .ZN(n7563) );
  AND2_X1 U5324 ( .A1(n7915), .A2(n7917), .ZN(n8009) );
  INV_X1 U5325 ( .A(n9552), .ZN(n4625) );
  AND4_X1 U5326 ( .A1(n5457), .A2(n5456), .A3(n5455), .A4(n5454), .ZN(n7642)
         );
  AND2_X1 U5327 ( .A1(n7377), .A2(n10029), .ZN(n7378) );
  AND4_X1 U5328 ( .A1(n5434), .A2(n5433), .A3(n5432), .A4(n5431), .ZN(n7554)
         );
  AND2_X1 U5329 ( .A1(n5024), .A2(n7908), .ZN(n5025) );
  NAND2_X1 U5330 ( .A1(n7273), .A2(n4700), .ZN(n5024) );
  AND2_X1 U5331 ( .A1(n8004), .A2(n7894), .ZN(n4700) );
  AND4_X1 U5332 ( .A1(n5382), .A2(n5381), .A3(n5380), .A4(n5379), .ZN(n7392)
         );
  NAND2_X1 U5333 ( .A1(n8005), .A2(n4925), .ZN(n4924) );
  NAND2_X1 U5334 ( .A1(n7105), .A2(n4927), .ZN(n4925) );
  INV_X1 U5335 ( .A(n4924), .ZN(n4923) );
  AND4_X1 U5336 ( .A1(n5409), .A2(n5408), .A3(n5407), .A4(n5406), .ZN(n7449)
         );
  NOR2_X1 U5337 ( .A1(n5027), .A2(n5026), .ZN(n7272) );
  INV_X1 U5338 ( .A(n7894), .ZN(n5026) );
  INV_X1 U5339 ( .A(n7271), .ZN(n5027) );
  AND2_X1 U5340 ( .A1(n7185), .A2(n10022), .ZN(n7377) );
  NAND2_X1 U5341 ( .A1(n7174), .A2(n7115), .ZN(n7269) );
  NAND2_X1 U5342 ( .A1(n7106), .A2(n7105), .ZN(n7271) );
  AOI21_X1 U5343 ( .B1(n4900), .B2(n4899), .A(n4898), .ZN(n7175) );
  AND2_X1 U5344 ( .A1(n7111), .A2(n7063), .ZN(n4899) );
  NAND2_X1 U5345 ( .A1(n4901), .A2(n4500), .ZN(n4898) );
  INV_X1 U5346 ( .A(n7061), .ZN(n4900) );
  NAND2_X1 U5347 ( .A1(n7065), .A2(n5000), .ZN(n7102) );
  NOR2_X1 U5348 ( .A1(n7111), .A2(n5001), .ZN(n5000) );
  INV_X1 U5349 ( .A(n7886), .ZN(n5001) );
  NAND2_X1 U5350 ( .A1(n4884), .A2(n4883), .ZN(n7186) );
  INV_X1 U5351 ( .A(n7059), .ZN(n4884) );
  OR2_X1 U5352 ( .A1(n7882), .A2(n6917), .ZN(n7065) );
  INV_X1 U5353 ( .A(n7004), .ZN(n4620) );
  NAND2_X1 U5354 ( .A1(n4622), .A2(n7013), .ZN(n4621) );
  NAND2_X1 U5355 ( .A1(n7849), .A2(n7876), .ZN(n9920) );
  NAND2_X1 U5356 ( .A1(n4531), .A2(n9945), .ZN(n9923) );
  NAND2_X1 U5357 ( .A1(n9936), .A2(n9935), .ZN(n9934) );
  OR2_X1 U5358 ( .A1(n7720), .A2(n6779), .ZN(n6934) );
  NAND2_X1 U5359 ( .A1(n5504), .A2(n5503), .ZN(n8578) );
  NAND2_X1 U5360 ( .A1(n4903), .A2(n7063), .ZN(n7110) );
  NAND2_X1 U5361 ( .A1(n7061), .A2(n7882), .ZN(n4903) );
  INV_X1 U5362 ( .A(n6852), .ZN(n4589) );
  AND2_X1 U5363 ( .A1(n5985), .A2(n4587), .ZN(n4586) );
  NAND2_X1 U5364 ( .A1(n6852), .A2(n4588), .ZN(n4587) );
  INV_X1 U5365 ( .A(n5951), .ZN(n4588) );
  INV_X1 U5366 ( .A(n9831), .ZN(n7321) );
  NAND2_X1 U5367 ( .A1(n7210), .A2(n6076), .ZN(n6080) );
  AND2_X1 U5368 ( .A1(n5913), .A2(n4613), .ZN(n6582) );
  NAND2_X1 U5369 ( .A1(n4611), .A2(n4983), .ZN(n4724) );
  NAND2_X1 U5370 ( .A1(n8622), .A2(n8623), .ZN(n4611) );
  OAI21_X1 U5371 ( .B1(n4981), .B2(n4535), .A(n4492), .ZN(n8685) );
  NAND2_X1 U5372 ( .A1(n4703), .A2(n6768), .ZN(n8695) );
  AND2_X1 U5373 ( .A1(n5951), .A2(n5950), .ZN(n8696) );
  NAND2_X1 U5374 ( .A1(n5949), .A2(n5948), .ZN(n5950) );
  OAI21_X1 U5375 ( .B1(n8658), .B2(n4711), .A(n4534), .ZN(n8703) );
  OR2_X1 U5376 ( .A1(n8659), .A2(n4711), .ZN(n4710) );
  INV_X1 U5377 ( .A(n6258), .ZN(n4711) );
  NAND2_X1 U5378 ( .A1(n8657), .A2(n4520), .ZN(n4712) );
  INV_X1 U5379 ( .A(n6394), .ZN(n7779) );
  NOR2_X1 U5380 ( .A1(n4716), .A2(n4512), .ZN(n8714) );
  INV_X1 U5381 ( .A(n4997), .ZN(n4716) );
  NAND2_X1 U5382 ( .A1(n4998), .A2(n4996), .ZN(n4995) );
  NAND2_X2 U5383 ( .A1(n5870), .A2(n5869), .ZN(n5991) );
  INV_X1 U5384 ( .A(n6709), .ZN(n4571) );
  INV_X1 U5385 ( .A(n6758), .ZN(n4574) );
  AND2_X1 U5386 ( .A1(n7024), .A2(n7023), .ZN(n7028) );
  AND2_X1 U5387 ( .A1(n4572), .A2(n4541), .ZN(n7730) );
  OR2_X1 U5388 ( .A1(n9039), .A2(n9038), .ZN(n4568) );
  NAND2_X1 U5389 ( .A1(n9125), .A2(n4774), .ZN(n9071) );
  NOR2_X1 U5390 ( .A1(n9143), .A2(n9126), .ZN(n9125) );
  INV_X1 U5391 ( .A(n9186), .ZN(n9153) );
  INV_X1 U5392 ( .A(n9094), .ZN(n4810) );
  NAND2_X1 U5393 ( .A1(n6369), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6386) );
  INV_X1 U5394 ( .A(n6371), .ZN(n6369) );
  NAND2_X1 U5395 ( .A1(n9200), .A2(n9093), .ZN(n9168) );
  OR2_X1 U5396 ( .A1(n9192), .A2(n9372), .ZN(n9116) );
  NAND2_X1 U5397 ( .A1(n9214), .A2(n4823), .ZN(n9200) );
  NOR2_X1 U5398 ( .A1(n9092), .A2(n8828), .ZN(n4823) );
  NAND2_X1 U5399 ( .A1(n5067), .A2(n5066), .ZN(n9219) );
  AOI21_X1 U5400 ( .B1(n5068), .B2(n5070), .A(n4521), .ZN(n5066) );
  AND2_X1 U5401 ( .A1(n8949), .A2(n9089), .ZN(n9229) );
  AOI21_X1 U5402 ( .B1(n5058), .B2(n5055), .A(n4539), .ZN(n5054) );
  NAND2_X1 U5403 ( .A1(n5058), .A2(n5057), .ZN(n5056) );
  OR2_X1 U5404 ( .A1(n5061), .A2(n4487), .ZN(n5055) );
  NAND2_X1 U5405 ( .A1(n9083), .A2(n4827), .ZN(n9275) );
  NOR2_X1 U5406 ( .A1(n9279), .A2(n4828), .ZN(n4827) );
  INV_X1 U5407 ( .A(n9082), .ZN(n4828) );
  OR2_X1 U5408 ( .A1(n9314), .A2(n9079), .ZN(n9083) );
  OAI21_X1 U5409 ( .B1(n9312), .B2(n9105), .A(n5060), .ZN(n9297) );
  NOR2_X1 U5410 ( .A1(n8974), .A2(n4822), .ZN(n4821) );
  INV_X1 U5411 ( .A(n8911), .ZN(n4822) );
  NAND2_X1 U5412 ( .A1(n7765), .A2(n7599), .ZN(n7673) );
  NOR2_X1 U5413 ( .A1(n9574), .A2(n9586), .ZN(n7756) );
  NAND2_X1 U5414 ( .A1(n7341), .A2(n8961), .ZN(n5065) );
  NAND2_X1 U5415 ( .A1(n7404), .A2(n9861), .ZN(n9743) );
  OR2_X1 U5416 ( .A1(n9844), .A2(n9839), .ZN(n8760) );
  NAND2_X1 U5417 ( .A1(n9839), .A2(n4756), .ZN(n9751) );
  INV_X1 U5418 ( .A(n9784), .ZN(n4756) );
  NAND2_X1 U5419 ( .A1(n9770), .A2(n9771), .ZN(n5072) );
  INV_X1 U5420 ( .A(n8962), .ZN(n9766) );
  NAND2_X1 U5421 ( .A1(n6181), .A2(n6180), .ZN(n7672) );
  INV_X1 U5422 ( .A(n9857), .ZN(n9735) );
  NAND2_X1 U5423 ( .A1(n6124), .A2(n6123), .ZN(n9601) );
  OR3_X1 U5424 ( .A1(n7544), .A2(n7635), .A3(n7620), .ZN(n6443) );
  XNOR2_X1 U5425 ( .A(n7831), .B(n7830), .ZN(n7829) );
  NAND2_X1 U5426 ( .A1(n5741), .A2(n5740), .ZN(n5758) );
  NAND2_X1 U5427 ( .A1(n4869), .A2(n4867), .ZN(n5741) );
  AOI21_X1 U5428 ( .B1(n4870), .B2(n4550), .A(n4868), .ZN(n4867) );
  INV_X1 U5429 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5876) );
  XNOR2_X1 U5430 ( .A(n5739), .B(n5738), .ZN(n7631) );
  OAI21_X1 U5431 ( .B1(n5674), .B2(n4550), .A(n4870), .ZN(n5739) );
  INV_X1 U5432 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5882) );
  NAND2_X1 U5433 ( .A1(n5874), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5883) );
  NOR2_X1 U5434 ( .A1(n5855), .A2(n4609), .ZN(n4608) );
  NAND2_X1 U5435 ( .A1(n6437), .A2(n5880), .ZN(n4609) );
  XNOR2_X1 U5436 ( .A(n5715), .B(n5714), .ZN(n7617) );
  INV_X1 U5437 ( .A(n5855), .ZN(n4610) );
  OR2_X1 U5438 ( .A1(n6068), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n6069) );
  XNOR2_X1 U5439 ( .A(n5322), .B(n5321), .ZN(n6529) );
  NAND2_X1 U5440 ( .A1(n4840), .A2(n5246), .ZN(n5268) );
  NAND2_X1 U5441 ( .A1(n5244), .A2(n5243), .ZN(n4840) );
  NAND2_X1 U5442 ( .A1(n5181), .A2(n5180), .ZN(n5184) );
  NAND2_X1 U5443 ( .A1(n5611), .A2(n5610), .ZN(n8549) );
  AND3_X1 U5444 ( .A1(n5488), .A2(n5487), .A3(n5486), .ZN(n8093) );
  AND3_X1 U5445 ( .A1(n5533), .A2(n5532), .A3(n5531), .ZN(n8130) );
  NAND2_X1 U5446 ( .A1(n5677), .A2(n5676), .ZN(n8533) );
  NOR2_X1 U5447 ( .A1(n6810), .A2(n4950), .ZN(n4949) );
  INV_X1 U5448 ( .A(n5171), .ZN(n4950) );
  NAND2_X1 U5449 ( .A1(n5596), .A2(n5595), .ZN(n8554) );
  AND4_X1 U5450 ( .A1(n5284), .A2(n5283), .A3(n5282), .A4(n5281), .ZN(n7062)
         );
  NAND2_X1 U5451 ( .A1(n4737), .A2(n8027), .ZN(n4701) );
  NAND2_X1 U5452 ( .A1(n8026), .A2(n8025), .ZN(n8027) );
  OR3_X1 U5453 ( .A1(n8026), .A2(n8020), .A3(n4940), .ZN(n4737) );
  XNOR2_X1 U5454 ( .A(n7837), .B(n8340), .ZN(n4702) );
  AOI21_X1 U5455 ( .B1(n4679), .B2(n4680), .A(n4675), .ZN(n4674) );
  AND4_X1 U5456 ( .A1(n5362), .A2(n5361), .A3(n5360), .A4(n5359), .ZN(n8158)
         );
  OR3_X1 U5457 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n5178) );
  NOR2_X1 U5458 ( .A1(n6613), .A2(n4502), .ZN(n6617) );
  NOR2_X1 U5459 ( .A1(n6617), .A2(n6616), .ZN(n6629) );
  AND2_X1 U5460 ( .A1(n5116), .A2(n5115), .ZN(n8356) );
  NAND2_X1 U5461 ( .A1(n4789), .A2(n8241), .ZN(n4788) );
  OR2_X1 U5462 ( .A1(n8242), .A2(n5128), .ZN(n4789) );
  AOI21_X1 U5463 ( .B1(n9503), .B2(n5220), .A(n7834), .ZN(n8246) );
  INV_X1 U5464 ( .A(n9922), .ZN(n9981) );
  INV_X1 U5466 ( .A(n8506), .ZN(n8507) );
  XNOR2_X1 U5467 ( .A(n8285), .B(n8284), .ZN(n8509) );
  NOR2_X1 U5468 ( .A1(n5123), .A2(n5122), .ZN(n4630) );
  NAND2_X1 U5469 ( .A1(n5789), .A2(n4746), .ZN(n4745) );
  XNOR2_X1 U5470 ( .A(n5112), .B(n5111), .ZN(n7249) );
  INV_X1 U5471 ( .A(n8356), .ZN(n8340) );
  NAND2_X1 U5472 ( .A1(n6278), .A2(n6277), .ZN(n9283) );
  AND2_X1 U5473 ( .A1(n7782), .A2(n8732), .ZN(n4714) );
  NOR2_X1 U5474 ( .A1(n8714), .A2(n4715), .ZN(n7800) );
  OR2_X1 U5475 ( .A1(n6415), .A2(n6416), .ZN(n4715) );
  NAND2_X1 U5476 ( .A1(n4592), .A2(n4591), .ZN(n7579) );
  AOI21_X1 U5477 ( .B1(n4595), .B2(n4598), .A(n4509), .ZN(n4591) );
  INV_X1 U5478 ( .A(n9215), .ZN(n9113) );
  AND2_X1 U5479 ( .A1(n6318), .A2(n6317), .ZN(n9266) );
  AND2_X1 U5480 ( .A1(n4833), .A2(n4832), .ZN(n9340) );
  NAND2_X1 U5481 ( .A1(n9099), .A2(n9100), .ZN(n4832) );
  NAND2_X1 U5482 ( .A1(n9101), .A2(n9427), .ZN(n4833) );
  NAND2_X1 U5483 ( .A1(n9149), .A2(n9096), .ZN(n9134) );
  NAND2_X1 U5484 ( .A1(n9154), .A2(n5074), .ZN(n9140) );
  NAND2_X1 U5485 ( .A1(n9154), .A2(n9122), .ZN(n9138) );
  INV_X1 U5486 ( .A(n9804), .ZN(n9319) );
  NAND2_X1 U5487 ( .A1(n7770), .A2(n6048), .ZN(n7772) );
  AOI21_X2 U5488 ( .B1(n9503), .B2(n6048), .A(n4560), .ZN(n9454) );
  INV_X1 U5489 ( .A(n9352), .ZN(n9462) );
  INV_X1 U5490 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9498) );
  AND2_X1 U5491 ( .A1(n4668), .A2(n5858), .ZN(n4667) );
  NOR2_X1 U5492 ( .A1(n4514), .A2(n4732), .ZN(n4731) );
  INV_X1 U5493 ( .A(n7888), .ZN(n4732) );
  AND2_X1 U5494 ( .A1(n4736), .A2(n7888), .ZN(n4733) );
  AOI21_X1 U5495 ( .B1(n7907), .B2(n7909), .A(n4751), .ZN(n4750) );
  NAND2_X1 U5496 ( .A1(n7910), .A2(n7976), .ZN(n4751) );
  NAND2_X1 U5497 ( .A1(n4662), .A2(n8782), .ZN(n4661) );
  NAND2_X1 U5498 ( .A1(n8781), .A2(n8780), .ZN(n4662) );
  NOR2_X1 U5499 ( .A1(n8903), .A2(n8864), .ZN(n4660) );
  OAI21_X1 U5500 ( .B1(n7928), .B2(n7984), .A(n4513), .ZN(n4739) );
  NAND2_X1 U5501 ( .A1(n4741), .A2(n7984), .ZN(n4740) );
  AOI211_X1 U5502 ( .C1(n7918), .C2(n7984), .A(n4743), .B(n5004), .ZN(n4742)
         );
  NOR2_X1 U5503 ( .A1(n4744), .A2(n7984), .ZN(n4743) );
  INV_X1 U5504 ( .A(n7917), .ZN(n4744) );
  NAND2_X1 U5505 ( .A1(n4657), .A2(n8806), .ZN(n8809) );
  AND2_X1 U5506 ( .A1(n8923), .A2(n9086), .ZN(n4639) );
  INV_X1 U5507 ( .A(n9089), .ZN(n4642) );
  INV_X1 U5508 ( .A(n9088), .ZN(n4643) );
  NAND2_X1 U5509 ( .A1(n8818), .A2(n4646), .ZN(n4644) );
  AND2_X1 U5510 ( .A1(n8922), .A2(n8865), .ZN(n4646) );
  NOR2_X1 U5511 ( .A1(n4648), .A2(n8865), .ZN(n4647) );
  NAND2_X1 U5512 ( .A1(n8951), .A2(n9084), .ZN(n4648) );
  OAI211_X1 U5513 ( .C1(n7957), .C2(n7976), .A(n4753), .B(n7959), .ZN(n4752)
         );
  NAND2_X1 U5514 ( .A1(n4666), .A2(n4665), .ZN(n4664) );
  NAND2_X1 U5515 ( .A1(n8826), .A2(n8864), .ZN(n4666) );
  INV_X1 U5516 ( .A(n4865), .ZN(n4864) );
  OAI21_X1 U5517 ( .B1(n5757), .B2(n4866), .A(n7706), .ZN(n4865) );
  INV_X1 U5518 ( .A(n5759), .ZN(n4866) );
  INV_X1 U5519 ( .A(n5519), .ZN(n4852) );
  NOR2_X1 U5520 ( .A1(n5266), .A2(n5242), .ZN(n4837) );
  INV_X1 U5521 ( .A(n5246), .ZN(n4839) );
  INV_X1 U5522 ( .A(n8125), .ZN(n4956) );
  AOI21_X1 U5523 ( .B1(n4934), .B2(n4936), .A(n4931), .ZN(n4930) );
  NAND2_X1 U5524 ( .A1(n4941), .A2(n7839), .ZN(n5138) );
  OR2_X1 U5525 ( .A1(n8496), .A2(n8245), .ZN(n7983) );
  AND2_X1 U5526 ( .A1(n4486), .A2(n8274), .ZN(n4638) );
  AND2_X1 U5527 ( .A1(n7955), .A2(n5038), .ZN(n5034) );
  NOR2_X1 U5528 ( .A1(n8419), .A2(n5039), .ZN(n5038) );
  INV_X1 U5529 ( .A(n7948), .ZN(n5039) );
  AND2_X1 U5530 ( .A1(n7816), .A2(n5011), .ZN(n5010) );
  NAND2_X1 U5531 ( .A1(n8465), .A2(n5012), .ZN(n5011) );
  INV_X1 U5532 ( .A(n7848), .ZN(n5012) );
  NOR2_X1 U5533 ( .A1(n5002), .A2(n4527), .ZN(n4687) );
  NOR2_X1 U5534 ( .A1(n4928), .A2(n4920), .ZN(n4918) );
  NAND2_X1 U5535 ( .A1(n7111), .A2(n4902), .ZN(n4901) );
  NOR2_X1 U5536 ( .A1(n7882), .A2(n4904), .ZN(n4902) );
  INV_X1 U5537 ( .A(n7063), .ZN(n4904) );
  NAND2_X1 U5538 ( .A1(n6983), .A2(n6695), .ZN(n7855) );
  AND2_X1 U5539 ( .A1(n7977), .A2(n7978), .ZN(n7992) );
  NAND2_X1 U5540 ( .A1(n4888), .A2(n4887), .ZN(n8354) );
  OR2_X1 U5541 ( .A1(n8456), .A2(n8455), .ZN(n8458) );
  NAND2_X1 U5542 ( .A1(n4889), .A2(n6940), .ZN(n9921) );
  NAND2_X1 U5543 ( .A1(n6994), .A2(n7996), .ZN(n4889) );
  NAND2_X1 U5544 ( .A1(n7852), .A2(n7870), .ZN(n9942) );
  AND2_X1 U5545 ( .A1(n5082), .A2(n5103), .ZN(n4974) );
  INV_X1 U5546 ( .A(n8623), .ZN(n4984) );
  NOR2_X1 U5547 ( .A1(n4498), .A2(n4983), .ZN(n4982) );
  NAND2_X1 U5548 ( .A1(n8630), .A2(n4990), .ZN(n4989) );
  INV_X1 U5549 ( .A(n8675), .ZN(n4990) );
  AND2_X1 U5550 ( .A1(n4987), .A2(n4549), .ZN(n4986) );
  NAND2_X1 U5551 ( .A1(n8630), .A2(n4988), .ZN(n4987) );
  NAND2_X1 U5552 ( .A1(n4979), .A2(n6030), .ZN(n4976) );
  INV_X1 U5553 ( .A(n8716), .ZN(n4996) );
  AOI21_X1 U5554 ( .B1(n4482), .B2(n7580), .A(n4494), .ZN(n4991) );
  AND2_X1 U5555 ( .A1(n9068), .A2(n8859), .ZN(n8985) );
  INV_X1 U5556 ( .A(n9013), .ZN(n8947) );
  AND2_X1 U5557 ( .A1(n9267), .A2(n4764), .ZN(n9189) );
  NOR2_X1 U5558 ( .A1(n9210), .A2(n4765), .ZN(n4764) );
  INV_X1 U5559 ( .A(n4766), .ZN(n4765) );
  INV_X1 U5560 ( .A(n4499), .ZN(n5070) );
  AND2_X1 U5561 ( .A1(n9476), .A2(n4767), .ZN(n4766) );
  OR2_X1 U5562 ( .A1(n9400), .A2(n9266), .ZN(n8950) );
  INV_X1 U5563 ( .A(n9105), .ZN(n5057) );
  INV_X1 U5564 ( .A(n5059), .ZN(n5058) );
  OAI21_X1 U5565 ( .B1(n4487), .B2(n9296), .A(n4522), .ZN(n5059) );
  AND2_X1 U5566 ( .A1(n4770), .A2(n4769), .ZN(n4768) );
  AND2_X1 U5567 ( .A1(n4772), .A2(n4771), .ZN(n4770) );
  NOR2_X1 U5568 ( .A1(n9443), .A2(n7672), .ZN(n4772) );
  NAND2_X1 U5569 ( .A1(n4817), .A2(n8899), .ZN(n7399) );
  INV_X1 U5570 ( .A(n9772), .ZN(n4817) );
  NAND2_X1 U5571 ( .A1(n9189), .A2(n9471), .ZN(n9190) );
  INV_X1 U5572 ( .A(n9617), .ZN(n4797) );
  NAND2_X1 U5573 ( .A1(n6492), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4796) );
  NOR2_X1 U5574 ( .A1(n5856), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4834) );
  INV_X1 U5575 ( .A(n5738), .ZN(n4868) );
  INV_X1 U5576 ( .A(n5690), .ZN(n4872) );
  NOR2_X1 U5577 ( .A1(n5691), .A2(n4875), .ZN(n4874) );
  INV_X1 U5578 ( .A(n5673), .ZN(n4875) );
  AOI21_X1 U5579 ( .B1(n4488), .B2(n4849), .A(n4528), .ZN(n4843) );
  NAND2_X1 U5580 ( .A1(n5417), .A2(n5393), .ZN(n5418) );
  NOR2_X1 U5581 ( .A1(n5216), .A2(n5215), .ZN(n5217) );
  NAND2_X1 U5582 ( .A1(n5189), .A2(n5188), .ZN(n5219) );
  NAND2_X1 U5583 ( .A1(n4972), .A2(n4971), .ZN(n4970) );
  INV_X1 U5584 ( .A(n5438), .ZN(n4971) );
  INV_X1 U5585 ( .A(n5638), .ZN(n5637) );
  OR2_X1 U5586 ( .A1(n5658), .A2(n8047), .ZN(n5678) );
  NAND2_X1 U5587 ( .A1(n8114), .A2(n5649), .ZN(n5668) );
  AND2_X1 U5588 ( .A1(n4959), .A2(n5557), .ZN(n4958) );
  INV_X1 U5589 ( .A(n8063), .ZN(n4959) );
  OR2_X1 U5590 ( .A1(n5597), .A2(n10318), .ZN(n5613) );
  NAND2_X1 U5591 ( .A1(n5612), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5638) );
  INV_X1 U5592 ( .A(n5613), .ZN(n5612) );
  INV_X1 U5593 ( .A(n5529), .ZN(n5528) );
  OR2_X1 U5594 ( .A1(n5429), .A2(n5428), .ZN(n5451) );
  NAND2_X1 U5595 ( .A1(n4973), .A2(n5415), .ZN(n7386) );
  INV_X1 U5596 ( .A(n7389), .ZN(n4973) );
  NAND2_X1 U5597 ( .A1(n5479), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5505) );
  AND2_X1 U5598 ( .A1(n7983), .A2(n7981), .ZN(n8017) );
  INV_X1 U5599 ( .A(n4684), .ZN(n4680) );
  AND2_X1 U5600 ( .A1(n4681), .A2(n4685), .ZN(n4675) );
  NAND2_X1 U5601 ( .A1(n4678), .A2(n4677), .ZN(n4676) );
  INV_X1 U5602 ( .A(n4681), .ZN(n4677) );
  INV_X1 U5603 ( .A(n4679), .ZN(n4678) );
  AND3_X1 U5604 ( .A1(n5509), .A2(n5508), .A3(n5507), .ZN(n7650) );
  AND4_X1 U5605 ( .A1(n5334), .A2(n5333), .A3(n5332), .A4(n5331), .ZN(n7114)
         );
  NOR2_X1 U5606 ( .A1(n9509), .A2(n4792), .ZN(n9511) );
  NAND2_X1 U5607 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n4792) );
  OR2_X1 U5608 ( .A1(n9523), .A2(n4506), .ZN(n4785) );
  AND2_X1 U5609 ( .A1(n6952), .A2(n6951), .ZN(n6955) );
  NAND2_X1 U5610 ( .A1(n8188), .A2(n8189), .ZN(n8191) );
  NOR2_X1 U5611 ( .A1(n8191), .A2(n8190), .ZN(n8202) );
  XNOR2_X1 U5612 ( .A(n8226), .B(n8232), .ZN(n8214) );
  NAND2_X1 U5613 ( .A1(n5109), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5113) );
  INV_X1 U5614 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5128) );
  NOR2_X1 U5615 ( .A1(n8213), .A2(n4775), .ZN(n8226) );
  NOR2_X1 U5616 ( .A1(n4777), .A2(n4776), .ZN(n4775) );
  INV_X1 U5617 ( .A(n8218), .ZN(n4777) );
  NAND2_X1 U5618 ( .A1(n8214), .A2(n8473), .ZN(n8228) );
  NOR2_X2 U5619 ( .A1(n8250), .A2(n8287), .ZN(n8249) );
  AND2_X1 U5620 ( .A1(n5770), .A2(n5769), .ZN(n8257) );
  NAND2_X1 U5621 ( .A1(n8299), .A2(n7819), .ZN(n8254) );
  OR2_X1 U5622 ( .A1(n5763), .A2(n5762), .ZN(n5821) );
  INV_X1 U5623 ( .A(n7993), .ZN(n8302) );
  NAND2_X1 U5624 ( .A1(n8312), .A2(n7969), .ZN(n8294) );
  INV_X1 U5625 ( .A(n8313), .ZN(n8319) );
  NAND2_X1 U5626 ( .A1(n8332), .A2(n5029), .ZN(n8312) );
  AND2_X1 U5627 ( .A1(n8313), .A2(n7965), .ZN(n5029) );
  NAND2_X1 U5628 ( .A1(n5722), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5763) );
  INV_X1 U5629 ( .A(n5724), .ZN(n5722) );
  NAND2_X1 U5630 ( .A1(n8346), .A2(n5030), .ZN(n8332) );
  AND2_X1 U5631 ( .A1(n8333), .A2(n7842), .ZN(n5030) );
  NAND2_X1 U5632 ( .A1(n8372), .A2(n7961), .ZN(n8347) );
  NAND2_X1 U5633 ( .A1(n8347), .A2(n8348), .ZN(n8346) );
  AND2_X1 U5634 ( .A1(n5708), .A2(n5707), .ZN(n8370) );
  OR2_X1 U5635 ( .A1(n8368), .A2(n8367), .ZN(n8372) );
  NAND2_X1 U5636 ( .A1(n4908), .A2(n4508), .ZN(n8389) );
  NAND2_X1 U5637 ( .A1(n5033), .A2(n5031), .ZN(n8379) );
  NAND2_X1 U5638 ( .A1(n5032), .A2(n7955), .ZN(n5031) );
  NAND2_X1 U5639 ( .A1(n8431), .A2(n5034), .ZN(n5033) );
  INV_X1 U5640 ( .A(n5035), .ZN(n5032) );
  NOR2_X1 U5641 ( .A1(n8394), .A2(n5036), .ZN(n5035) );
  INV_X1 U5642 ( .A(n7950), .ZN(n5036) );
  NAND2_X1 U5643 ( .A1(n8431), .A2(n5038), .ZN(n5037) );
  AND2_X1 U5644 ( .A1(n5582), .A2(n5581), .ZN(n8427) );
  AOI21_X1 U5645 ( .B1(n5010), .B2(n5013), .A(n5008), .ZN(n5007) );
  INV_X1 U5646 ( .A(n7944), .ZN(n5008) );
  INV_X1 U5647 ( .A(n8465), .ZN(n5013) );
  NAND2_X1 U5648 ( .A1(n7814), .A2(n7848), .ZN(n8464) );
  OAI21_X1 U5649 ( .B1(n7428), .B2(n4627), .A(n4623), .ZN(n7657) );
  AOI21_X1 U5650 ( .B1(n4626), .B2(n8008), .A(n4524), .ZN(n4623) );
  NAND2_X1 U5651 ( .A1(n7378), .A2(n4881), .ZN(n7568) );
  NAND2_X1 U5652 ( .A1(n4530), .A2(n7530), .ZN(n4693) );
  NAND2_X1 U5653 ( .A1(n7378), .A2(n10035), .ZN(n7420) );
  NAND2_X1 U5654 ( .A1(n5374), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U5655 ( .A1(n7894), .A2(n7899), .ZN(n8004) );
  INV_X1 U5656 ( .A(n7113), .ZN(n8003) );
  AND4_X1 U5657 ( .A1(n5310), .A2(n5309), .A3(n5308), .A4(n5307), .ZN(n7177)
         );
  NAND2_X1 U5658 ( .A1(n5277), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5304) );
  INV_X1 U5659 ( .A(n5279), .ZN(n5277) );
  INV_X1 U5660 ( .A(n6978), .ZN(n4886) );
  NAND2_X1 U5661 ( .A1(n4616), .A2(n4614), .ZN(n7061) );
  AOI21_X1 U5662 ( .B1(n4621), .B2(n4615), .A(n4523), .ZN(n4614) );
  NAND2_X1 U5663 ( .A1(n5227), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U5664 ( .A1(n5251), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5279) );
  INV_X1 U5665 ( .A(n5252), .ZN(n5251) );
  NAND2_X1 U5666 ( .A1(n5019), .A2(n5017), .ZN(n5016) );
  NOR2_X1 U5667 ( .A1(n5020), .A2(n6943), .ZN(n5019) );
  INV_X1 U5668 ( .A(n4635), .ZN(n4634) );
  OAI21_X1 U5669 ( .B1(n5221), .B2(n5192), .A(n5197), .ZN(n4635) );
  NAND2_X1 U5670 ( .A1(n9945), .A2(n9967), .ZN(n9947) );
  OR2_X1 U5671 ( .A1(n6924), .A2(n6923), .ZN(n6927) );
  OAI211_X1 U5672 ( .C1(n6556), .C2(n6488), .A(n5165), .B(n5164), .ZN(n6914)
         );
  INV_X1 U5673 ( .A(n9942), .ZN(n9935) );
  AND2_X1 U5674 ( .A1(n7855), .A2(n7853), .ZN(n9936) );
  AND4_X1 U5675 ( .A1(n5156), .A2(n5155), .A3(n5154), .A4(n5153), .ZN(n6937)
         );
  OR2_X1 U5676 ( .A1(n5254), .A2(n5152), .ZN(n5154) );
  NAND2_X1 U5677 ( .A1(n5761), .A2(n5760), .ZN(n8511) );
  OAI211_X1 U5678 ( .C1(n6995), .C2(n5017), .A(n5015), .B(n7876), .ZN(n7005)
         );
  NAND2_X1 U5679 ( .A1(n7996), .A2(n5021), .ZN(n5015) );
  INV_X1 U5680 ( .A(n10034), .ZN(n10002) );
  AND2_X1 U5681 ( .A1(n5791), .A2(n5792), .ZN(n9955) );
  AND2_X1 U5682 ( .A1(n5119), .A2(n5079), .ZN(n5093) );
  NAND2_X1 U5683 ( .A1(n5497), .A2(n5093), .ZN(n5121) );
  NOR2_X1 U5684 ( .A1(n5120), .A2(n5399), .ZN(n4746) );
  INV_X1 U5685 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5120) );
  INV_X1 U5686 ( .A(n5121), .ZN(n5123) );
  NAND2_X1 U5687 ( .A1(n4748), .A2(n4747), .ZN(n5789) );
  INV_X1 U5688 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4747) );
  INV_X1 U5689 ( .A(n5787), .ZN(n4748) );
  NAND2_X1 U5690 ( .A1(n5119), .A2(n5497), .ZN(n5787) );
  OR2_X1 U5691 ( .A1(n5300), .A2(n5299), .ZN(n5323) );
  INV_X1 U5692 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6038) );
  NAND2_X1 U5693 ( .A1(n4704), .A2(n4979), .ZN(n7038) );
  AND2_X1 U5694 ( .A1(n6031), .A2(n5989), .ZN(n4590) );
  NOR2_X1 U5695 ( .A1(n6182), .A2(n7219), .ZN(n6201) );
  NAND2_X1 U5696 ( .A1(n4992), .A2(n4991), .ZN(n7688) );
  NOR2_X1 U5697 ( .A1(n6039), .A2(n6038), .ZN(n6060) );
  OR2_X1 U5698 ( .A1(n6367), .A2(n8636), .ZN(n4998) );
  AOI21_X1 U5699 ( .B1(n4604), .B2(n4605), .A(n4540), .ZN(n4603) );
  OR2_X1 U5700 ( .A1(n8645), .A2(n8646), .ZN(n8649) );
  INV_X1 U5701 ( .A(n8615), .ZN(n4605) );
  OR2_X1 U5702 ( .A1(n8667), .A2(n8666), .ZN(n4999) );
  NAND2_X1 U5703 ( .A1(n6582), .A2(n6581), .ZN(n6580) );
  NAND2_X1 U5704 ( .A1(n6309), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6328) );
  INV_X1 U5705 ( .A(n6311), .ZN(n6309) );
  AOI21_X1 U5706 ( .B1(n4724), .B2(n4723), .A(n4722), .ZN(n8684) );
  INV_X1 U5707 ( .A(n4989), .ZN(n4723) );
  NAND2_X1 U5708 ( .A1(n4986), .A2(n6336), .ZN(n4722) );
  NOR2_X1 U5709 ( .A1(n6126), .A2(n6125), .ZN(n6143) );
  NOR2_X1 U5710 ( .A1(n4706), .A2(n4600), .ZN(n4599) );
  INV_X1 U5711 ( .A(n6076), .ZN(n4600) );
  NAND2_X1 U5712 ( .A1(n6105), .A2(n4709), .ZN(n4706) );
  NAND2_X1 U5713 ( .A1(n4707), .A2(n4709), .ZN(n4705) );
  OAI21_X1 U5714 ( .B1(n4994), .B2(n4708), .A(n7435), .ZN(n4707) );
  OR2_X1 U5715 ( .A1(n6266), .A2(n6265), .ZN(n6280) );
  NAND2_X1 U5716 ( .A1(n6243), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6266) );
  INV_X1 U5717 ( .A(n6245), .ZN(n6243) );
  AND3_X1 U5718 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6012) );
  NAND2_X1 U5719 ( .A1(n6012), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6039) );
  OAI21_X1 U5720 ( .B1(n4992), .B2(n4582), .A(n4580), .ZN(n8728) );
  INV_X1 U5721 ( .A(n4581), .ZN(n4580) );
  OAI21_X1 U5722 ( .B1(n4991), .B2(n4582), .A(n6211), .ZN(n4581) );
  INV_X1 U5723 ( .A(n6215), .ZN(n4582) );
  OAI21_X1 U5724 ( .B1(n8863), .B2(n4672), .A(n4669), .ZN(n8868) );
  NOR2_X1 U5725 ( .A1(n9010), .A2(n4655), .ZN(n4654) );
  OR2_X1 U5726 ( .A1(n8872), .A2(n8946), .ZN(n4655) );
  AND2_X1 U5727 ( .A1(n9454), .A2(n9066), .ZN(n9010) );
  OR2_X1 U5728 ( .A1(n5991), .A2(n5954), .ZN(n5956) );
  NAND2_X1 U5729 ( .A1(n5952), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5932) );
  OAI211_X1 U5730 ( .C1(n8754), .C2(n5895), .A(n5873), .B(n5872), .ZN(n7123)
         );
  INV_X1 U5731 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5845) );
  OR2_X1 U5732 ( .A1(n5938), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n6002) );
  INV_X1 U5733 ( .A(n6711), .ZN(n4570) );
  OR2_X1 U5734 ( .A1(n6759), .A2(n6758), .ZN(n4577) );
  AND2_X1 U5735 ( .A1(n9699), .A2(n6904), .ZN(n6907) );
  NOR2_X1 U5736 ( .A1(n7227), .A2(n4561), .ZN(n7514) );
  XNOR2_X1 U5737 ( .A(n9126), .B(n9028), .ZN(n9123) );
  OR2_X1 U5738 ( .A1(n4544), .A2(n4806), .ZN(n4803) );
  NAND2_X1 U5739 ( .A1(n9167), .A2(n8948), .ZN(n9181) );
  OR2_X1 U5740 ( .A1(n6340), .A2(n6339), .ZN(n6353) );
  OR2_X1 U5741 ( .A1(n6328), .A2(n8689), .ZN(n6340) );
  NAND2_X1 U5742 ( .A1(n9090), .A2(n4490), .ZN(n9214) );
  NAND2_X1 U5743 ( .A1(n9267), .A2(n4767), .ZN(n9235) );
  NAND2_X1 U5744 ( .A1(n9267), .A2(n9256), .ZN(n9246) );
  AND2_X1 U5745 ( .A1(n9282), .A2(n9272), .ZN(n9267) );
  NAND2_X1 U5746 ( .A1(n9087), .A2(n9086), .ZN(n9243) );
  NOR2_X1 U5747 ( .A1(n9085), .A2(n4826), .ZN(n4825) );
  NAND2_X1 U5748 ( .A1(n6279), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6293) );
  INV_X1 U5749 ( .A(n6280), .ZN(n6279) );
  AND2_X1 U5750 ( .A1(n9281), .A2(n9486), .ZN(n9282) );
  AND2_X1 U5751 ( .A1(n9292), .A2(n9291), .ZN(n9313) );
  NAND2_X1 U5752 ( .A1(n6201), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6222) );
  NAND2_X1 U5753 ( .A1(n6221), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6245) );
  INV_X1 U5754 ( .A(n6222), .ZN(n6221) );
  NAND2_X1 U5755 ( .A1(n7756), .A2(n4770), .ZN(n9316) );
  INV_X1 U5756 ( .A(n4819), .ZN(n4818) );
  OAI21_X1 U5757 ( .B1(n7599), .B2(n4820), .A(n8917), .ZN(n4819) );
  INV_X1 U5758 ( .A(n4821), .ZN(n4820) );
  NAND2_X1 U5759 ( .A1(n5049), .A2(n4501), .ZN(n9104) );
  OR2_X1 U5760 ( .A1(n9443), .A2(n9031), .ZN(n5050) );
  NAND2_X1 U5761 ( .A1(n7756), .A2(n4772), .ZN(n7697) );
  AND2_X1 U5762 ( .A1(n7756), .A2(n8788), .ZN(n7676) );
  NAND2_X1 U5763 ( .A1(n4762), .A2(n4489), .ZN(n9574) );
  NAND2_X1 U5764 ( .A1(n5046), .A2(n5042), .ZN(n5041) );
  INV_X1 U5765 ( .A(n7608), .ZN(n5042) );
  AND2_X1 U5766 ( .A1(n5048), .A2(n5045), .ZN(n9563) );
  NAND2_X1 U5767 ( .A1(n4762), .A2(n4759), .ZN(n9573) );
  OR2_X1 U5768 ( .A1(n7469), .A2(n9879), .ZN(n4758) );
  NOR2_X1 U5769 ( .A1(n9744), .A2(n9879), .ZN(n7365) );
  OR2_X1 U5770 ( .A1(n9743), .A2(n7322), .ZN(n9744) );
  NOR2_X1 U5771 ( .A1(n9729), .A2(n5064), .ZN(n5063) );
  INV_X1 U5772 ( .A(n7312), .ZN(n5064) );
  NAND2_X1 U5773 ( .A1(n4813), .A2(n4814), .ZN(n4812) );
  INV_X1 U5774 ( .A(n8896), .ZN(n4814) );
  NOR2_X1 U5775 ( .A1(n9751), .A2(n7412), .ZN(n7404) );
  NAND2_X1 U5776 ( .A1(n7399), .A2(n8896), .ZN(n9756) );
  NAND2_X1 U5777 ( .A1(n4757), .A2(n9831), .ZN(n9784) );
  NOR2_X1 U5778 ( .A1(n8698), .A2(n7164), .ZN(n7256) );
  NAND2_X1 U5779 ( .A1(n7158), .A2(n4801), .ZN(n4798) );
  INV_X1 U5780 ( .A(n7154), .ZN(n8956) );
  NAND2_X1 U5781 ( .A1(n7159), .A2(n7158), .ZN(n8894) );
  CLKBUF_X1 U5782 ( .A(n5904), .Z(n5905) );
  INV_X1 U5783 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5848) );
  CLKBUF_X1 U5784 ( .A(n7124), .Z(n8959) );
  NAND2_X1 U5785 ( .A1(n9813), .A2(n4773), .ZN(n7164) );
  INV_X1 U5786 ( .A(n4801), .ZN(n8955) );
  OR2_X1 U5787 ( .A1(n8959), .A2(n4801), .ZN(n7159) );
  INV_X1 U5788 ( .A(n8959), .ZN(n7139) );
  NAND2_X1 U5789 ( .A1(n7631), .A2(n6048), .ZN(n6384) );
  AND4_X1 U5790 ( .A1(n6228), .A2(n6227), .A3(n6226), .A4(n6225), .ZN(n9423)
         );
  NAND2_X1 U5791 ( .A1(n6162), .A2(n6161), .ZN(n9586) );
  AND2_X1 U5792 ( .A1(n4480), .A2(n7138), .ZN(n9857) );
  INV_X1 U5793 ( .A(SI_30_), .ZN(n4842) );
  XNOR2_X1 U5794 ( .A(n7829), .B(SI_30_), .ZN(n8746) );
  XNOR2_X1 U5795 ( .A(n7725), .B(n7710), .ZN(n8853) );
  NOR2_X1 U5796 ( .A1(n5856), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n5078) );
  XNOR2_X1 U5797 ( .A(n7707), .B(n7706), .ZN(n7770) );
  NAND2_X1 U5798 ( .A1(n4863), .A2(n5759), .ZN(n7707) );
  NAND2_X1 U5799 ( .A1(n5758), .A2(n5757), .ZN(n4863) );
  NAND2_X1 U5800 ( .A1(n5674), .A2(n5673), .ZN(n5692) );
  OAI21_X1 U5801 ( .B1(n5652), .B2(n5651), .A(n5650), .ZN(n5672) );
  AND2_X1 U5802 ( .A1(n5673), .A2(n5655), .ZN(n5671) );
  NAND2_X1 U5803 ( .A1(n4878), .A2(n5609), .ZN(n5626) );
  OAI21_X1 U5804 ( .B1(n5441), .B2(n4857), .A(n4855), .ZN(n5520) );
  NAND2_X1 U5805 ( .A1(n4854), .A2(n5466), .ZN(n5492) );
  NAND2_X1 U5806 ( .A1(n5441), .A2(n4859), .ZN(n4854) );
  NAND2_X1 U5807 ( .A1(n5441), .A2(n5440), .ZN(n5468) );
  NAND2_X1 U5808 ( .A1(n4845), .A2(n4846), .ZN(n5390) );
  OR2_X1 U5809 ( .A1(n5347), .A2(n4849), .ZN(n4845) );
  NAND2_X1 U5810 ( .A1(n4699), .A2(n5344), .ZN(n4698) );
  NAND2_X1 U5811 ( .A1(n5347), .A2(n5346), .ZN(n4699) );
  OR2_X1 U5812 ( .A1(n6046), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n6068) );
  XNOR2_X1 U5813 ( .A(n5182), .B(n10398), .ZN(n5180) );
  NAND2_X1 U5814 ( .A1(n4877), .A2(n5132), .ZN(n5889) );
  NAND2_X1 U5815 ( .A1(n6832), .A2(n5265), .ZN(n6878) );
  NAND2_X1 U5816 ( .A1(n5746), .A2(n5745), .ZN(n8281) );
  XNOR2_X1 U5817 ( .A(n5668), .B(n5666), .ZN(n8046) );
  NAND2_X1 U5818 ( .A1(n5341), .A2(n7081), .ZN(n8052) );
  NAND2_X1 U5819 ( .A1(n5571), .A2(n5570), .ZN(n8559) );
  INV_X1 U5820 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10250) );
  NAND2_X1 U5821 ( .A1(n4933), .A2(n4934), .ZN(n6474) );
  OR2_X1 U5822 ( .A1(n6833), .A2(n4936), .ZN(n4933) );
  AND4_X1 U5823 ( .A1(n5146), .A2(n5145), .A3(n5144), .A4(n5143), .ZN(n7720)
         );
  OR2_X1 U5824 ( .A1(n5254), .A2(n5141), .ZN(n5145) );
  NAND2_X1 U5825 ( .A1(n5687), .A2(n4946), .ZN(n8079) );
  NAND2_X1 U5826 ( .A1(n8100), .A2(n8099), .ZN(n4946) );
  NAND2_X1 U5827 ( .A1(n8090), .A2(n5518), .ZN(n7624) );
  NAND2_X1 U5828 ( .A1(n5527), .A2(n5526), .ZN(n8571) );
  CLKBUF_X1 U5829 ( .A(n7080), .Z(n7084) );
  AND2_X1 U5830 ( .A1(n7386), .A2(n5416), .ZN(n7447) );
  OAI22_X1 U5831 ( .A1(n5340), .A2(n4965), .B1(n5365), .B2(n5366), .ZN(n4963)
         );
  NAND2_X1 U5832 ( .A1(n5539), .A2(n5538), .ZN(n8126) );
  NAND2_X1 U5833 ( .A1(n6833), .A2(n6834), .ZN(n6832) );
  INV_X1 U5834 ( .A(n7717), .ZN(n8131) );
  NAND2_X1 U5835 ( .A1(n4944), .A2(n4942), .ZN(n8136) );
  INV_X1 U5836 ( .A(n4943), .ZN(n4942) );
  NOR2_X1 U5837 ( .A1(n4947), .A2(n4948), .ZN(n4945) );
  INV_X1 U5838 ( .A(n6937), .ZN(n8165) );
  AND2_X1 U5839 ( .A1(n4785), .A2(n4784), .ZN(n6599) );
  INV_X1 U5840 ( .A(n6575), .ZN(n4784) );
  INV_X1 U5841 ( .A(n4785), .ZN(n6576) );
  NOR2_X1 U5842 ( .A1(n6602), .A2(n6601), .ZN(n6613) );
  NOR2_X1 U5843 ( .A1(n6629), .A2(n4552), .ZN(n6633) );
  AOI21_X1 U5844 ( .B1(n6665), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6664), .ZN(
        n6668) );
  AOI21_X1 U5845 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n6866), .A(n6865), .ZN(
        n6870) );
  NOR2_X1 U5846 ( .A1(n6870), .A2(n6869), .ZN(n6961) );
  NOR2_X1 U5847 ( .A1(n6965), .A2(n6964), .ZN(n7044) );
  NOR2_X1 U5848 ( .A1(n6961), .A2(n4780), .ZN(n6965) );
  AND2_X1 U5849 ( .A1(n6962), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4780) );
  NOR2_X1 U5850 ( .A1(n7044), .A2(n4778), .ZN(n7046) );
  NOR2_X1 U5851 ( .A1(n4779), .A2(n7117), .ZN(n4778) );
  INV_X1 U5852 ( .A(n7050), .ZN(n4779) );
  NOR2_X1 U5853 ( .A1(n7243), .A2(n7244), .ZN(n7282) );
  NOR2_X1 U5854 ( .A1(n7282), .A2(n4782), .ZN(n7286) );
  AND2_X1 U5855 ( .A1(n7283), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4782) );
  NAND2_X1 U5856 ( .A1(n7286), .A2(n7285), .ZN(n7454) );
  NAND2_X1 U5857 ( .A1(n7454), .A2(n4781), .ZN(n7455) );
  OR2_X1 U5858 ( .A1(n7458), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4781) );
  XNOR2_X1 U5859 ( .A(n8186), .B(n4783), .ZN(n8169) );
  NAND2_X1 U5860 ( .A1(n8169), .A2(n7571), .ZN(n8188) );
  AND2_X1 U5861 ( .A1(n6574), .A2(n5818), .ZN(n9527) );
  NOR2_X1 U5862 ( .A1(n8206), .A2(n8205), .ZN(n8213) );
  NAND2_X1 U5863 ( .A1(n5721), .A2(n5720), .ZN(n8523) );
  OAI21_X1 U5864 ( .B1(n8275), .B2(n4895), .A(n4486), .ZN(n8351) );
  NAND2_X1 U5865 ( .A1(n4892), .A2(n8276), .ZN(n8353) );
  NAND2_X1 U5866 ( .A1(n8275), .A2(n8367), .ZN(n4892) );
  NAND2_X1 U5867 ( .A1(n8420), .A2(n8270), .ZN(n4914) );
  INV_X1 U5868 ( .A(n8433), .ZN(n8414) );
  NAND2_X1 U5869 ( .A1(n8431), .A2(n7948), .ZN(n8408) );
  NAND2_X1 U5870 ( .A1(n5547), .A2(n5546), .ZN(n8568) );
  AND2_X1 U5871 ( .A1(n4907), .A2(n8261), .ZN(n8483) );
  NAND2_X1 U5872 ( .A1(n4907), .A2(n4485), .ZN(n8482) );
  OR2_X1 U5873 ( .A1(n8263), .A2(n8262), .ZN(n4907) );
  NOR2_X1 U5874 ( .A1(n4686), .A2(n5002), .ZN(n8479) );
  INV_X1 U5875 ( .A(n4688), .ZN(n4686) );
  NAND2_X1 U5876 ( .A1(n7649), .A2(n7927), .ZN(n7812) );
  INV_X1 U5877 ( .A(n4882), .ZN(n7569) );
  NAND2_X1 U5878 ( .A1(n9552), .A2(n4626), .ZN(n7560) );
  NOR2_X1 U5879 ( .A1(n4625), .A2(n4624), .ZN(n7536) );
  INV_X1 U5880 ( .A(n7535), .ZN(n4624) );
  NAND2_X1 U5881 ( .A1(n5426), .A2(n5425), .ZN(n7534) );
  NAND2_X1 U5882 ( .A1(n7428), .A2(n7528), .ZN(n9552) );
  NAND2_X1 U5883 ( .A1(n4695), .A2(n7910), .ZN(n7529) );
  NAND2_X1 U5884 ( .A1(n5025), .A2(n4696), .ZN(n7417) );
  OAI21_X1 U5885 ( .B1(n7269), .B2(n4924), .A(n4919), .ZN(n7375) );
  AOI21_X1 U5886 ( .B1(n4923), .B2(n4928), .A(n4920), .ZN(n4919) );
  NAND2_X1 U5887 ( .A1(n4922), .A2(n4927), .ZN(n7270) );
  NAND2_X1 U5888 ( .A1(n7269), .A2(n4927), .ZN(n4921) );
  NAND2_X1 U5889 ( .A1(n7271), .A2(n5028), .ZN(n7370) );
  NAND2_X1 U5890 ( .A1(n7065), .A2(n7886), .ZN(n7066) );
  NAND2_X1 U5891 ( .A1(n4619), .A2(n4621), .ZN(n6970) );
  NAND2_X1 U5892 ( .A1(n4620), .A2(n4481), .ZN(n4619) );
  NAND2_X1 U5893 ( .A1(n5022), .A2(n7859), .ZN(n9914) );
  NAND2_X1 U5894 ( .A1(n6995), .A2(n7858), .ZN(n5022) );
  OAI22_X1 U5895 ( .A1(n5196), .A2(n6491), .B1(n6490), .B2(n6556), .ZN(n4897)
         );
  OR2_X1 U5896 ( .A1(n5194), .A2(n6498), .ZN(n5136) );
  AND2_X1 U5897 ( .A1(n9927), .A2(n6947), .ZN(n9944) );
  OR2_X1 U5898 ( .A1(n9956), .A2(n6925), .ZN(n9924) );
  INV_X1 U5899 ( .A(n9944), .ZN(n8478) );
  AND2_X1 U5900 ( .A1(n5830), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9962) );
  NAND4_X1 U5901 ( .A1(n5093), .A2(n5497), .A3(n5040), .A4(n5118), .ZN(n8602)
         );
  INV_X1 U5902 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5040) );
  XNOR2_X1 U5903 ( .A(n5094), .B(n8600), .ZN(n8606) );
  NAND2_X1 U5904 ( .A1(n8602), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5094) );
  NOR2_X1 U5905 ( .A1(n5157), .A2(n4794), .ZN(n4793) );
  NAND2_X1 U5906 ( .A1(n4537), .A2(P2_IR_REG_1__SCAN_IN), .ZN(n4795) );
  NOR2_X1 U5907 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4794) );
  NAND2_X1 U5908 ( .A1(n7832), .A2(P2_U3152), .ZN(n7729) );
  AND2_X1 U5909 ( .A1(n6050), .A2(n6049), .ZN(n9861) );
  NAND2_X1 U5910 ( .A1(n7345), .A2(n6105), .ZN(n7439) );
  NAND2_X1 U5911 ( .A1(n8694), .A2(n5951), .ZN(n4975) );
  NAND2_X1 U5912 ( .A1(n8703), .A2(n8706), .ZN(n4612) );
  NAND2_X1 U5913 ( .A1(n4985), .A2(n8674), .ZN(n8629) );
  OR2_X1 U5914 ( .A1(n8677), .A2(n8675), .ZN(n4985) );
  INV_X1 U5915 ( .A(n9032), .ZN(n9568) );
  NAND2_X1 U5916 ( .A1(n7617), .A2(n6048), .ZN(n4566) );
  OR2_X1 U5917 ( .A1(n6018), .A2(n6504), .ZN(n6006) );
  NAND2_X1 U5918 ( .A1(n8614), .A2(n4601), .ZN(n8667) );
  NAND2_X1 U5919 ( .A1(n4606), .A2(n4605), .ZN(n4601) );
  NAND2_X1 U5920 ( .A1(n4583), .A2(n4586), .ZN(n6841) );
  NAND2_X1 U5921 ( .A1(n4975), .A2(n6852), .ZN(n6851) );
  INV_X1 U5922 ( .A(n4724), .ZN(n8677) );
  NAND2_X1 U5923 ( .A1(n7577), .A2(n6156), .ZN(n7589) );
  NAND2_X1 U5924 ( .A1(n4593), .A2(n4595), .ZN(n7520) );
  OR2_X1 U5925 ( .A1(n7210), .A2(n4598), .ZN(n4593) );
  NAND2_X1 U5926 ( .A1(n4594), .A2(n4705), .ZN(n7522) );
  NAND2_X1 U5927 ( .A1(n7210), .A2(n4599), .ZN(n4594) );
  INV_X1 U5928 ( .A(n4712), .ZN(n8705) );
  AND3_X1 U5929 ( .A1(n6024), .A2(n6023), .A3(n6022), .ZN(n9847) );
  AND2_X1 U5930 ( .A1(n6377), .A2(n6376), .ZN(n9204) );
  INV_X1 U5931 ( .A(n9027), .ZN(n4651) );
  INV_X1 U5932 ( .A(n9204), .ZN(n9372) );
  NAND2_X1 U5933 ( .A1(n6360), .A2(n6359), .ZN(n9215) );
  AND4_X1 U5934 ( .A1(n6149), .A2(n6148), .A3(n6147), .A4(n6146), .ZN(n9597)
         );
  INV_X1 U5935 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6544) );
  AND4_X1 U5936 ( .A1(n6115), .A2(n6114), .A3(n6113), .A4(n6112), .ZN(n9598)
         );
  INV_X1 U5937 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6546) );
  AND4_X1 U5938 ( .A1(n6066), .A2(n6065), .A3(n6064), .A4(n6063), .ZN(n7348)
         );
  CLKBUF_X1 U5939 ( .A(n7123), .Z(n8886) );
  NAND2_X1 U5940 ( .A1(n6652), .A2(n6651), .ZN(n6708) );
  NAND2_X1 U5941 ( .A1(n6708), .A2(n6709), .ZN(n9646) );
  OAI22_X1 U5942 ( .A1(n6759), .A2(n4573), .B1(n4575), .B2(n6899), .ZN(n9669)
         );
  AND2_X1 U5943 ( .A1(n6900), .A2(n4496), .ZN(n4575) );
  NAND2_X1 U5944 ( .A1(n4576), .A2(n4574), .ZN(n4573) );
  XNOR2_X1 U5945 ( .A(n7514), .B(n7513), .ZN(n7229) );
  INV_X1 U5946 ( .A(n4572), .ZN(n7515) );
  NOR2_X1 U5947 ( .A1(n7731), .A2(n7732), .ZN(n9039) );
  INV_X1 U5948 ( .A(n4568), .ZN(n9037) );
  NOR2_X1 U5949 ( .A1(n9052), .A2(n9051), .ZN(n9050) );
  AND2_X1 U5950 ( .A1(n4568), .A2(n4567), .ZN(n9052) );
  NAND2_X1 U5951 ( .A1(n7742), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4567) );
  XNOR2_X1 U5952 ( .A(n9071), .B(n9454), .ZN(n9062) );
  OAI21_X1 U5953 ( .B1(n9153), .B2(n9757), .A(n9152), .ZN(n9358) );
  NAND2_X1 U5954 ( .A1(n7726), .A2(n6048), .ZN(n6403) );
  AND2_X1 U5955 ( .A1(n6455), .A2(n6387), .ZN(n9174) );
  NAND2_X1 U5956 ( .A1(n9394), .A2(n4499), .ZN(n9230) );
  NAND2_X1 U5957 ( .A1(n6327), .A2(n6326), .ZN(n9239) );
  NAND2_X1 U5958 ( .A1(n9245), .A2(n9244), .ZN(n9394) );
  NAND2_X1 U5959 ( .A1(n9275), .A2(n9084), .ZN(n9263) );
  AOI21_X1 U5960 ( .B1(n9297), .B2(n9296), .A(n4487), .ZN(n9280) );
  NAND2_X1 U5961 ( .A1(n9083), .A2(n9082), .ZN(n9277) );
  NAND2_X1 U5962 ( .A1(n6264), .A2(n6263), .ZN(n9307) );
  NAND2_X1 U5963 ( .A1(n7673), .A2(n4821), .ZN(n7701) );
  NAND2_X1 U5964 ( .A1(n7673), .A2(n8911), .ZN(n7674) );
  OR2_X1 U5965 ( .A1(n9807), .A2(n9755), .ZN(n9781) );
  NAND2_X1 U5966 ( .A1(n5072), .A2(n7309), .ZN(n9765) );
  INV_X1 U5967 ( .A(n9813), .ZN(n8888) );
  INV_X1 U5968 ( .A(n9781), .ZN(n9572) );
  AND2_X1 U5969 ( .A1(n9332), .A2(n9335), .ZN(n9451) );
  NOR2_X1 U5970 ( .A1(n9343), .A2(n4830), .ZN(n4829) );
  INV_X1 U5971 ( .A(n9342), .ZN(n4831) );
  AOI21_X1 U5972 ( .B1(n9349), .B2(n9867), .A(n9348), .ZN(n9459) );
  INV_X1 U5973 ( .A(n9192), .ZN(n9471) );
  AOI211_X1 U5974 ( .C1(n9382), .C2(n9867), .A(n9381), .B(n9380), .ZN(n9473)
         );
  INV_X1 U5975 ( .A(n9283), .ZN(n9486) );
  AND2_X1 U5976 ( .A1(n6443), .A2(n6439), .ZN(n9810) );
  OAI21_X1 U5977 ( .B1(n7829), .B2(n4842), .A(n4532), .ZN(n4841) );
  XNOR2_X1 U5978 ( .A(n5758), .B(n5757), .ZN(n7726) );
  XNOR2_X1 U5979 ( .A(n5877), .B(n5876), .ZN(n7635) );
  XNOR2_X1 U5980 ( .A(n5672), .B(n5671), .ZN(n7486) );
  INV_X1 U5981 ( .A(n8871), .ZN(n9761) );
  INV_X1 U5982 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10192) );
  XNOR2_X1 U5983 ( .A(n6083), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9672) );
  INV_X1 U5984 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6528) );
  XNOR2_X1 U5985 ( .A(n5189), .B(n5188), .ZN(n6496) );
  NOR2_X1 U5986 ( .A1(n10093), .A2(n10494), .ZN(n10119) );
  NAND2_X1 U5987 ( .A1(n4952), .A2(n4503), .ZN(n6817) );
  AOI21_X1 U5988 ( .B1(n4702), .B2(n8028), .A(n4701), .ZN(n8034) );
  OAI21_X1 U5989 ( .B1(n8240), .B2(n8356), .A(n4787), .ZN(P2_U3264) );
  AOI21_X1 U5990 ( .B1(n4790), .B2(n8356), .A(n4788), .ZN(n4787) );
  NAND2_X1 U5991 ( .A1(n10062), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n4929) );
  AOI21_X1 U5992 ( .B1(n4483), .B2(n10043), .A(n4495), .ZN(n4632) );
  NOR2_X1 U5993 ( .A1(n10042), .A2(n9995), .ZN(n4633) );
  NAND2_X1 U5994 ( .A1(n7800), .A2(n4714), .ZN(n7798) );
  OR2_X1 U5995 ( .A1(n9026), .A2(n9025), .ZN(n4649) );
  INV_X1 U5996 ( .A(n6067), .ZN(n6000) );
  OR2_X1 U5997 ( .A1(n7013), .A2(n9918), .ZN(n4481) );
  OAI21_X1 U5998 ( .B1(n8011), .B2(n5003), .A(n7929), .ZN(n5002) );
  NAND2_X1 U5999 ( .A1(n5320), .A2(SI_9_), .ZN(n5344) );
  NOR2_X1 U6000 ( .A1(n6176), .A2(n4993), .ZN(n4482) );
  NAND2_X1 U6001 ( .A1(n8508), .A2(n8507), .ZN(n4483) );
  AND2_X1 U6002 ( .A1(n4926), .A2(n7373), .ZN(n4484) );
  AND2_X1 U6003 ( .A1(n7927), .A2(n7923), .ZN(n7562) );
  INV_X1 U6004 ( .A(n7562), .ZN(n5004) );
  AND2_X1 U6005 ( .A1(n4527), .A2(n8261), .ZN(n4485) );
  AND2_X1 U6006 ( .A1(n8352), .A2(n4893), .ZN(n4486) );
  AND2_X1 U6007 ( .A1(n9307), .A2(n9324), .ZN(n4487) );
  NAND2_X1 U6008 ( .A1(n6292), .A2(n6291), .ZN(n9406) );
  INV_X1 U6009 ( .A(n9799), .ZN(n4773) );
  INV_X1 U6010 ( .A(n9084), .ZN(n4826) );
  AND2_X1 U6011 ( .A1(n4846), .A2(n5388), .ZN(n4488) );
  INV_X1 U6012 ( .A(n7978), .ZN(n4683) );
  NAND2_X1 U6013 ( .A1(n5657), .A2(n5656), .ZN(n8538) );
  NAND2_X1 U6014 ( .A1(n9096), .A2(n8875), .ZN(n9155) );
  AND2_X1 U6015 ( .A1(n4759), .A2(n4763), .ZN(n4489) );
  AND2_X1 U6016 ( .A1(n4824), .A2(n9089), .ZN(n4490) );
  INV_X1 U6017 ( .A(n5266), .ZN(n5267) );
  XNOR2_X1 U6018 ( .A(n5269), .B(SI_6_), .ZN(n5266) );
  AND2_X1 U6019 ( .A1(n4880), .A2(n4881), .ZN(n4491) );
  INV_X1 U6020 ( .A(n7373), .ZN(n4920) );
  NOR2_X1 U6021 ( .A1(n4546), .A2(n4982), .ZN(n4492) );
  NAND2_X1 U6022 ( .A1(n5037), .A2(n5035), .ZN(n4493) );
  AND2_X1 U6023 ( .A1(n6175), .A2(n7586), .ZN(n4494) );
  NAND2_X1 U6024 ( .A1(n5065), .A2(n7312), .ZN(n9725) );
  NAND2_X1 U6025 ( .A1(n4960), .A2(n5557), .ZN(n8062) );
  NAND2_X1 U6026 ( .A1(n7249), .A2(n8340), .ZN(n8029) );
  INV_X1 U6027 ( .A(n8029), .ZN(n4939) );
  NAND2_X1 U6028 ( .A1(n6080), .A2(n6079), .ZN(n7344) );
  AND2_X1 U6029 ( .A1(n10042), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n4495) );
  INV_X2 U6030 ( .A(n5194), .ZN(n5220) );
  NAND2_X1 U6031 ( .A1(n4566), .A2(n6368), .ZN(n9192) );
  OR2_X1 U6032 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6760), .ZN(n4496) );
  INV_X1 U6033 ( .A(n8164), .ZN(n4755) );
  OR2_X1 U6034 ( .A1(n8546), .A2(n8150), .ZN(n7955) );
  AND2_X1 U6035 ( .A1(n5865), .A2(n5864), .ZN(n5915) );
  OR2_X1 U6036 ( .A1(n5105), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n4497) );
  OR2_X1 U6037 ( .A1(n4989), .A2(n6336), .ZN(n4498) );
  INV_X1 U6038 ( .A(n4928), .ZN(n4927) );
  NOR2_X1 U6039 ( .A1(n10022), .A2(n8158), .ZN(n4928) );
  OR2_X1 U6040 ( .A1(n9256), .A2(n9266), .ZN(n4499) );
  NAND2_X1 U6041 ( .A1(n7112), .A2(n8161), .ZN(n4500) );
  OR2_X1 U6042 ( .A1(n8744), .A2(n8652), .ZN(n4501) );
  INV_X1 U6043 ( .A(n5929), .ZN(n5952) );
  NAND2_X1 U6044 ( .A1(n5478), .A2(n5477), .ZN(n7658) );
  OAI21_X1 U6045 ( .B1(n6496), .B2(n5194), .A(n4896), .ZN(n6999) );
  INV_X1 U6046 ( .A(n6999), .ZN(n4879) );
  INV_X1 U6047 ( .A(n8367), .ZN(n4894) );
  INV_X1 U6048 ( .A(n4627), .ZN(n4626) );
  NAND2_X1 U6049 ( .A1(n7921), .A2(n7535), .ZN(n4627) );
  AND2_X1 U6050 ( .A1(n6614), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4502) );
  OR2_X1 U6051 ( .A1(n5187), .A2(n5186), .ZN(n4503) );
  INV_X1 U6052 ( .A(n7859), .ZN(n5014) );
  OR3_X1 U6053 ( .A1(n9010), .A2(n9024), .A3(n8745), .ZN(n4504) );
  NOR2_X1 U6054 ( .A1(n9647), .A2(n4571), .ZN(n4505) );
  AND2_X1 U6055 ( .A1(n9526), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4506) );
  AND2_X1 U6056 ( .A1(n7090), .A2(n7094), .ZN(n4507) );
  XNOR2_X1 U6057 ( .A(n5096), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5098) );
  OR2_X1 U6058 ( .A1(n9221), .A2(n9207), .ZN(n9091) );
  AND2_X1 U6059 ( .A1(n4910), .A2(n8390), .ZN(n4508) );
  OR2_X1 U6060 ( .A1(n7424), .A2(n7449), .ZN(n7910) );
  INV_X1 U6061 ( .A(n7910), .ZN(n4694) );
  NAND2_X1 U6062 ( .A1(n8749), .A2(n8748), .ZN(n9070) );
  INV_X1 U6063 ( .A(n9070), .ZN(n4774) );
  AND2_X1 U6064 ( .A1(n6138), .A2(n6137), .ZN(n4509) );
  OR2_X1 U6065 ( .A1(n7567), .A2(n7642), .ZN(n7915) );
  INV_X1 U6066 ( .A(n7915), .ZN(n4690) );
  AND2_X1 U6067 ( .A1(n5286), .A2(n5285), .ZN(n4510) );
  INV_X1 U6068 ( .A(n6275), .ZN(n4713) );
  AND2_X1 U6069 ( .A1(n4908), .A2(n4910), .ZN(n4511) );
  INV_X1 U6070 ( .A(n9443), .ZN(n8744) );
  NAND2_X1 U6071 ( .A1(n6200), .A2(n6199), .ZN(n9443) );
  OR2_X1 U6072 ( .A1(n8715), .A2(n4995), .ZN(n4512) );
  AND2_X1 U6073 ( .A1(n8262), .A2(n4740), .ZN(n4513) );
  NAND2_X1 U6074 ( .A1(n5402), .A2(n5401), .ZN(n7424) );
  AND2_X1 U6075 ( .A1(n6916), .A2(n7885), .ZN(n4514) );
  AND2_X1 U6076 ( .A1(n9214), .A2(n9091), .ZN(n4515) );
  INV_X1 U6077 ( .A(n6899), .ZN(n4576) );
  NAND2_X1 U6078 ( .A1(n5920), .A2(n5845), .ZN(n5938) );
  XNOR2_X1 U6079 ( .A(n5389), .B(n5368), .ZN(n5388) );
  OR2_X1 U6080 ( .A1(n4797), .A2(n4796), .ZN(n4516) );
  NOR2_X1 U6081 ( .A1(n8396), .A2(n4913), .ZN(n4912) );
  AND2_X1 U6082 ( .A1(n4894), .A2(n4754), .ZN(n4517) );
  NAND2_X1 U6083 ( .A1(n7637), .A2(n5510), .ZN(n4518) );
  AND2_X1 U6084 ( .A1(n9090), .A2(n9089), .ZN(n4519) );
  AND2_X1 U6085 ( .A1(n4713), .A2(n6258), .ZN(n4520) );
  INV_X1 U6086 ( .A(n4888), .ZN(n8363) );
  INV_X1 U6087 ( .A(n5242), .ZN(n5243) );
  XNOR2_X1 U6088 ( .A(n5245), .B(SI_5_), .ZN(n5242) );
  INV_X1 U6089 ( .A(n9210), .ZN(n9375) );
  NAND2_X1 U6090 ( .A1(n6350), .A2(n6349), .ZN(n9210) );
  AND2_X1 U6091 ( .A1(n9239), .A2(n9254), .ZN(n4521) );
  OR2_X1 U6092 ( .A1(n9283), .A2(n9415), .ZN(n4522) );
  OR2_X1 U6093 ( .A1(n9352), .A2(n9356), .ZN(n8873) );
  NOR2_X2 U6094 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5157) );
  NOR2_X1 U6095 ( .A1(n7884), .A2(n8163), .ZN(n4523) );
  INV_X1 U6096 ( .A(n9729), .ZN(n7313) );
  AND2_X1 U6097 ( .A1(n8778), .A2(n8774), .ZN(n9729) );
  NOR2_X1 U6098 ( .A1(n7567), .A2(n8154), .ZN(n4524) );
  NOR2_X1 U6099 ( .A1(n8529), .A2(n8277), .ZN(n4525) );
  NOR2_X1 U6100 ( .A1(n8571), .A2(n8466), .ZN(n4526) );
  NAND2_X1 U6101 ( .A1(n6242), .A2(n6241), .ZN(n9317) );
  INV_X1 U6102 ( .A(n9317), .ZN(n4769) );
  NAND2_X1 U6103 ( .A1(n7848), .A2(n7846), .ZN(n4527) );
  AND2_X1 U6104 ( .A1(n5389), .A2(SI_11_), .ZN(n4528) );
  AND2_X1 U6105 ( .A1(n5269), .A2(SI_6_), .ZN(n4529) );
  INV_X1 U6106 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5399) );
  INV_X1 U6107 ( .A(n6945), .ZN(n4618) );
  AND2_X1 U6108 ( .A1(n8873), .A2(n8876), .ZN(n9137) );
  INV_X1 U6109 ( .A(n9137), .ZN(n5076) );
  INV_X1 U6110 ( .A(n9839), .ZN(n9750) );
  OR2_X1 U6111 ( .A1(n7528), .A2(n4694), .ZN(n4530) );
  AND2_X1 U6112 ( .A1(n9967), .A2(n4879), .ZN(n4531) );
  NAND2_X1 U6113 ( .A1(n7831), .A2(n7830), .ZN(n4532) );
  AND2_X1 U6114 ( .A1(n5037), .A2(n7950), .ZN(n4533) );
  AND2_X1 U6115 ( .A1(n4710), .A2(n6275), .ZN(n4534) );
  INV_X1 U6116 ( .A(n6105), .ZN(n4708) );
  OR2_X1 U6117 ( .A1(n4498), .A2(n4984), .ZN(n4535) );
  AND2_X1 U6118 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4536) );
  AND2_X1 U6119 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4537) );
  NOR2_X1 U6120 ( .A1(n9462), .A2(n9356), .ZN(n4538) );
  NOR2_X1 U6121 ( .A1(n9265), .A2(n9486), .ZN(n4539) );
  OR2_X1 U6122 ( .A1(n8636), .A2(n8666), .ZN(n4540) );
  INV_X1 U6123 ( .A(n5046), .ZN(n5045) );
  NAND2_X1 U6124 ( .A1(n9560), .A2(n5047), .ZN(n5046) );
  NOR2_X1 U6125 ( .A1(n5085), .A2(n5084), .ZN(n5119) );
  OR2_X1 U6126 ( .A1(n8288), .A2(n8296), .ZN(n7977) );
  INV_X1 U6127 ( .A(n7977), .ZN(n4685) );
  INV_X1 U6128 ( .A(n8503), .ZN(n8250) );
  AOI21_X1 U6129 ( .B1(n8746), .B2(n5220), .A(n7822), .ZN(n8503) );
  OR2_X1 U6130 ( .A1(n7514), .A2(n7513), .ZN(n4541) );
  AND2_X1 U6131 ( .A1(n7123), .A2(n5912), .ZN(n4542) );
  AND2_X1 U6132 ( .A1(n6651), .A2(n4570), .ZN(n4543) );
  AND2_X1 U6133 ( .A1(n4809), .A2(n9137), .ZN(n4544) );
  INV_X1 U6134 ( .A(n5061), .ZN(n5060) );
  NOR2_X1 U6135 ( .A1(n4769), .A2(n9302), .ZN(n5061) );
  AND2_X1 U6136 ( .A1(n8346), .A2(n7842), .ZN(n4545) );
  INV_X1 U6137 ( .A(n9476), .ZN(n9221) );
  AND2_X1 U6138 ( .A1(n6338), .A2(n6337), .ZN(n9476) );
  NOR2_X1 U6139 ( .A1(n4986), .A2(n6336), .ZN(n4546) );
  INV_X1 U6140 ( .A(n7035), .ZN(n4978) );
  AND2_X1 U6141 ( .A1(n8332), .A2(n7965), .ZN(n4547) );
  OR2_X1 U6142 ( .A1(n7388), .A2(n5438), .ZN(n4548) );
  NAND2_X1 U6143 ( .A1(n6325), .A2(n6324), .ZN(n4549) );
  INV_X1 U6144 ( .A(n5023), .ZN(n5028) );
  NAND2_X1 U6145 ( .A1(n7273), .A2(n7894), .ZN(n5023) );
  INV_X1 U6146 ( .A(n5075), .ZN(n5074) );
  NAND2_X1 U6147 ( .A1(n5076), .A2(n9122), .ZN(n5075) );
  OR2_X1 U6148 ( .A1(n7106), .A2(n5023), .ZN(n4696) );
  OR2_X1 U6149 ( .A1(n5714), .A2(n4872), .ZN(n4550) );
  NAND2_X1 U6150 ( .A1(n8464), .A2(n8465), .ZN(n8444) );
  AND2_X1 U6151 ( .A1(n9267), .A2(n4766), .ZN(n4551) );
  AND2_X1 U6152 ( .A1(n6630), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4552) );
  INV_X1 U6153 ( .A(n8674), .ZN(n4988) );
  INV_X1 U6154 ( .A(n9441), .ZN(n9583) );
  NAND2_X1 U6155 ( .A1(n5367), .A2(n5351), .ZN(n4553) );
  NAND2_X1 U6156 ( .A1(n5698), .A2(n5697), .ZN(n8529) );
  INV_X1 U6157 ( .A(n8529), .ZN(n4887) );
  NAND2_X1 U6158 ( .A1(n5009), .A2(n5007), .ZN(n8424) );
  NAND2_X1 U6159 ( .A1(n7563), .A2(n7562), .ZN(n7649) );
  NAND2_X1 U6160 ( .A1(n9091), .A2(n9002), .ZN(n9220) );
  INV_X1 U6161 ( .A(n9220), .ZN(n4824) );
  AND2_X1 U6162 ( .A1(n4960), .A2(n4958), .ZN(n4554) );
  NAND2_X1 U6163 ( .A1(n6289), .A2(n6290), .ZN(n4983) );
  OR2_X1 U6164 ( .A1(n7579), .A2(n7580), .ZN(n7577) );
  INV_X1 U6165 ( .A(n9162), .ZN(n9466) );
  NAND2_X1 U6166 ( .A1(n6403), .A2(n6402), .ZN(n9162) );
  NAND3_X1 U6167 ( .A1(n4720), .A2(n4719), .A3(n4610), .ZN(n4555) );
  NAND2_X1 U6168 ( .A1(n5497), .A2(n5082), .ZN(n4556) );
  AND2_X1 U6169 ( .A1(n5627), .A2(n5609), .ZN(n4557) );
  NAND2_X1 U6170 ( .A1(n6220), .A2(n6219), .ZN(n9437) );
  INV_X1 U6171 ( .A(n9437), .ZN(n4771) );
  NAND2_X1 U6172 ( .A1(n5449), .A2(n5448), .ZN(n7567) );
  INV_X1 U6173 ( .A(n7567), .ZN(n4880) );
  AND2_X1 U6174 ( .A1(n7434), .A2(n8871), .ZN(n8864) );
  OR2_X1 U6175 ( .A1(n4758), .A2(n9744), .ZN(n4558) );
  AND2_X1 U6176 ( .A1(n4577), .A2(n4496), .ZN(n4559) );
  NOR2_X1 U6177 ( .A1(n8855), .A2(n10261), .ZN(n4560) );
  AND2_X1 U6178 ( .A1(n7228), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4561) );
  NAND2_X1 U6179 ( .A1(n4967), .A2(n5340), .ZN(n7081) );
  NAND2_X1 U6180 ( .A1(n6080), .A2(n4994), .ZN(n7345) );
  AND2_X1 U6181 ( .A1(n7910), .A2(n7909), .ZN(n8007) );
  INV_X1 U6182 ( .A(n8007), .ZN(n4926) );
  INV_X1 U6183 ( .A(n7876), .ZN(n5020) );
  NAND2_X1 U6184 ( .A1(n9981), .A2(n8164), .ZN(n7876) );
  AND2_X1 U6185 ( .A1(n7709), .A2(n10392), .ZN(n4562) );
  INV_X1 U6186 ( .A(n7996), .ZN(n7858) );
  NAND2_X1 U6187 ( .A1(n7875), .A2(n7859), .ZN(n7996) );
  INV_X1 U6188 ( .A(n7234), .ZN(n4721) );
  INV_X1 U6189 ( .A(n8187), .ZN(n4783) );
  NAND2_X1 U6190 ( .A1(n5303), .A2(n5302), .ZN(n7112) );
  INV_X1 U6191 ( .A(n7112), .ZN(n4883) );
  INV_X1 U6192 ( .A(n10001), .ZN(n4885) );
  INV_X1 U6193 ( .A(n9879), .ZN(n4761) );
  NAND2_X1 U6194 ( .A1(n6142), .A2(n6141), .ZN(n9592) );
  INV_X1 U6195 ( .A(n9592), .ZN(n4763) );
  XOR2_X1 U6196 ( .A(n7833), .B(n10204), .Z(n4563) );
  INV_X1 U6197 ( .A(n9783), .ZN(n4757) );
  OR2_X1 U6198 ( .A1(n5928), .A2(n5927), .ZN(n6767) );
  NOR2_X1 U6199 ( .A1(n7835), .A2(n7828), .ZN(n4564) );
  AND2_X1 U6200 ( .A1(n4505), .A2(n6708), .ZN(n4565) );
  INV_X1 U6201 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4717) );
  NAND2_X1 U6202 ( .A1(n5827), .A2(n7828), .ZN(n7991) );
  INV_X1 U6203 ( .A(n7991), .ZN(n4940) );
  INV_X1 U6204 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5880) );
  INV_X1 U6205 ( .A(n9522), .ZN(n4786) );
  INV_X1 U6206 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n4776) );
  INV_X2 U6207 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  OAI21_X1 U6208 ( .B1(n7389), .B2(n4548), .A(n4970), .ZN(n7550) );
  NAND2_X1 U6209 ( .A1(n5631), .A2(n5630), .ZN(n5652) );
  OAI21_X1 U6210 ( .B1(n5544), .B2(n5543), .A(n5542), .ZN(n5560) );
  OAI21_X1 U6211 ( .B1(n4656), .B2(n4504), .A(n4653), .ZN(n4652) );
  NAND3_X1 U6212 ( .A1(n8863), .A2(n9028), .A3(n8864), .ZN(n8867) );
  NAND2_X1 U6213 ( .A1(n4652), .A2(n4651), .ZN(n4650) );
  NAND2_X1 U6214 ( .A1(n5522), .A2(n5521), .ZN(n5544) );
  AOI21_X1 U6215 ( .B1(n4656), .B2(n4654), .A(n9022), .ZN(n4653) );
  AOI211_X1 U6216 ( .C1(n9019), .C2(n9018), .A(n9017), .B(n9016), .ZN(n9020)
         );
  NAND2_X1 U6217 ( .A1(n4952), .A2(n4951), .ZN(n6814) );
  NAND2_X1 U6218 ( .A1(n4964), .A2(n4962), .ZN(n7205) );
  OR2_X2 U6219 ( .A1(n5138), .A2(n5139), .ZN(n5140) );
  NAND2_X1 U6220 ( .A1(n7549), .A2(n5463), .ZN(n7638) );
  XNOR2_X1 U6221 ( .A(n5161), .B(n5134), .ZN(n5160) );
  NAND2_X1 U6222 ( .A1(n7695), .A2(n5050), .ZN(n5049) );
  INV_X1 U6223 ( .A(n7671), .ZN(n5053) );
  NAND2_X1 U6224 ( .A1(n9344), .A2(n4831), .ZN(n4830) );
  INV_X1 U6225 ( .A(n4963), .ZN(n4962) );
  NAND2_X1 U6226 ( .A1(n9340), .A2(n4829), .ZN(n9458) );
  NAND2_X1 U6227 ( .A1(n8339), .A2(n8516), .ZN(n8321) );
  NOR2_X2 U6228 ( .A1(n8546), .A2(n8412), .ZN(n8400) );
  NOR2_X1 U6229 ( .A1(n9923), .A2(n9922), .ZN(n7009) );
  NAND2_X1 U6230 ( .A1(n5124), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n5125) );
  NAND2_X1 U6231 ( .A1(n5608), .A2(n5607), .ZN(n4878) );
  NAND2_X1 U6232 ( .A1(n4836), .A2(n4838), .ZN(n5289) );
  NAND2_X1 U6233 ( .A1(n4844), .A2(n4843), .ZN(n5419) );
  NAND2_X1 U6234 ( .A1(n5563), .A2(n5562), .ZN(n5591) );
  NAND2_X1 U6235 ( .A1(n4873), .A2(n5690), .ZN(n5715) );
  NAND2_X1 U6236 ( .A1(n4853), .A2(n4851), .ZN(n5522) );
  NAND2_X1 U6237 ( .A1(n4650), .A2(n4649), .ZN(P1_U3240) );
  NAND2_X1 U6238 ( .A1(n4663), .A2(n9153), .ZN(n8840) );
  NAND2_X1 U6239 ( .A1(n4664), .A2(n8834), .ZN(n8845) );
  NOR2_X1 U6240 ( .A1(n8869), .A2(n8870), .ZN(n4656) );
  NAND2_X1 U6241 ( .A1(n6652), .A2(n4543), .ZN(n4569) );
  OAI21_X1 U6242 ( .B1(n4505), .B2(n6711), .A(n4569), .ZN(n6713) );
  INV_X1 U6243 ( .A(n4577), .ZN(n6757) );
  NOR2_X1 U6244 ( .A1(n9669), .A2(n9668), .ZN(n9667) );
  MUX2_X1 U6245 ( .A(n6647), .B(P1_REG2_REG_1__SCAN_IN), .S(n6680), .Z(n6682)
         );
  INV_X1 U6246 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4579) );
  NAND2_X1 U6247 ( .A1(n8728), .A2(n8730), .ZN(n6217) );
  OR2_X1 U6248 ( .A1(n8694), .A2(n4589), .ZN(n4583) );
  NAND2_X1 U6249 ( .A1(n8694), .A2(n4586), .ZN(n4585) );
  NAND3_X1 U6250 ( .A1(n4585), .A2(n4590), .A3(n4584), .ZN(n4704) );
  NAND2_X1 U6251 ( .A1(n7210), .A2(n4595), .ZN(n4592) );
  OR2_X1 U6252 ( .A1(n8684), .A2(n4604), .ZN(n4606) );
  NAND3_X1 U6253 ( .A1(n8614), .A2(n4602), .A3(n4603), .ZN(n4997) );
  NAND2_X1 U6254 ( .A1(n8684), .A2(n4605), .ZN(n4602) );
  NAND2_X1 U6255 ( .A1(n4720), .A2(n4719), .ZN(n5884) );
  NAND3_X1 U6256 ( .A1(n4720), .A2(n4719), .A3(n4608), .ZN(n5874) );
  NAND2_X1 U6257 ( .A1(n4542), .A2(n7773), .ZN(n4613) );
  AND2_X2 U6258 ( .A1(n7773), .A2(n5912), .ZN(n6394) );
  NAND2_X1 U6259 ( .A1(n7004), .A2(n4617), .ZN(n4616) );
  INV_X1 U6260 ( .A(n7997), .ZN(n4622) );
  XNOR2_X2 U6261 ( .A(n4629), .B(n5118), .ZN(n5818) );
  NAND2_X1 U6262 ( .A1(n8509), .A2(n4633), .ZN(n4631) );
  NAND2_X1 U6263 ( .A1(n4631), .A2(n4632), .ZN(P2_U3517) );
  AOI21_X1 U6264 ( .B1(n8509), .B2(n10041), .A(n4483), .ZN(n8585) );
  NAND2_X1 U6265 ( .A1(n8389), .A2(n4638), .ZN(n4891) );
  INV_X1 U6266 ( .A(n8275), .ZN(n8362) );
  NAND3_X1 U6267 ( .A1(n4645), .A2(n4644), .A3(n4639), .ZN(n4640) );
  NAND2_X1 U6268 ( .A1(n8820), .A2(n4647), .ZN(n4645) );
  AND2_X1 U6269 ( .A1(n4645), .A2(n4644), .ZN(n8823) );
  NAND2_X1 U6270 ( .A1(n6067), .A2(n9794), .ZN(n5925) );
  NAND4_X2 U6271 ( .A1(n5916), .A2(n5917), .A3(n5918), .A4(n5919), .ZN(n9794)
         );
  AND2_X1 U6272 ( .A1(n5878), .A2(n4668), .ZN(n5861) );
  NAND2_X1 U6273 ( .A1(n5878), .A2(n4667), .ZN(n9497) );
  NAND2_X1 U6274 ( .A1(n5878), .A2(n5077), .ZN(n5892) );
  NAND2_X1 U6275 ( .A1(n4673), .A2(n4674), .ZN(n7836) );
  NAND2_X1 U6276 ( .A1(n8254), .A2(n4676), .ZN(n4673) );
  NAND2_X1 U6277 ( .A1(n4688), .A2(n4687), .ZN(n7814) );
  NAND2_X1 U6278 ( .A1(n4691), .A2(n4693), .ZN(n7531) );
  NAND3_X1 U6279 ( .A1(n5025), .A2(n4692), .A3(n4696), .ZN(n4691) );
  NAND3_X1 U6280 ( .A1(n4696), .A2(n5025), .A3(n7909), .ZN(n4695) );
  MUX2_X1 U6281 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n6492), .Z(n5182) );
  NAND2_X1 U6282 ( .A1(n6767), .A2(n6769), .ZN(n4703) );
  INV_X1 U6283 ( .A(n7038), .ZN(n6057) );
  NAND2_X1 U6284 ( .A1(n8658), .A2(n8659), .ZN(n8657) );
  NAND2_X1 U6285 ( .A1(n4718), .A2(n4717), .ZN(n5886) );
  INV_X1 U6286 ( .A(n5884), .ZN(n4718) );
  NOR2_X2 U6287 ( .A1(n5853), .A2(n5906), .ZN(n4719) );
  INV_X2 U6288 ( .A(n5904), .ZN(n4720) );
  OAI21_X1 U6289 ( .B1(n4726), .B2(n4725), .A(n7947), .ZN(n7936) );
  NAND2_X1 U6290 ( .A1(n7950), .A2(n7945), .ZN(n4725) );
  OR2_X1 U6291 ( .A1(n7873), .A2(n4735), .ZN(n4729) );
  NAND2_X1 U6292 ( .A1(n4728), .A2(n4730), .ZN(n7892) );
  NAND3_X1 U6293 ( .A1(n4729), .A2(n4734), .A3(n4733), .ZN(n4728) );
  NAND2_X1 U6294 ( .A1(n7880), .A2(n7976), .ZN(n4736) );
  OR2_X1 U6295 ( .A1(n7872), .A2(n4735), .ZN(n4734) );
  AOI21_X1 U6296 ( .B1(n4752), .B2(n7963), .A(n7962), .ZN(n7967) );
  NAND2_X1 U6297 ( .A1(n7756), .A2(n4768), .ZN(n9303) );
  AND3_X2 U6298 ( .A1(n5923), .A2(n5922), .A3(n4516), .ZN(n9813) );
  MUX2_X1 U6299 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6569), .S(n9506), .Z(n9509)
         );
  NAND2_X1 U6300 ( .A1(n8959), .A2(n7158), .ZN(n4799) );
  NAND3_X1 U6301 ( .A1(n4799), .A2(n8956), .A3(n4798), .ZN(n7259) );
  NAND2_X1 U6302 ( .A1(n9168), .A2(n4804), .ZN(n4802) );
  NAND2_X1 U6303 ( .A1(n9168), .A2(n9095), .ZN(n4811) );
  NAND2_X1 U6304 ( .A1(n4802), .A2(n4803), .ZN(n9098) );
  NAND2_X1 U6305 ( .A1(n4811), .A2(n4809), .ZN(n9149) );
  AND2_X1 U6306 ( .A1(n4811), .A2(n4810), .ZN(n9151) );
  INV_X1 U6307 ( .A(n4815), .ZN(n4813) );
  OAI211_X1 U6308 ( .C1(n9772), .C2(n4815), .A(n4812), .B(n8900), .ZN(n7333)
         );
  OAI21_X1 U6309 ( .B1(n7765), .B2(n4820), .A(n4818), .ZN(n9076) );
  NAND2_X1 U6310 ( .A1(n9275), .A2(n4825), .ZN(n9087) );
  NAND2_X1 U6311 ( .A1(n5878), .A2(n4834), .ZN(n4835) );
  NAND2_X1 U6312 ( .A1(n5244), .A2(n4837), .ZN(n4836) );
  NAND2_X1 U6313 ( .A1(n5347), .A2(n4488), .ZN(n4844) );
  NAND2_X1 U6314 ( .A1(n5441), .A2(n4855), .ZN(n4853) );
  NAND2_X1 U6315 ( .A1(n5674), .A2(n4870), .ZN(n4869) );
  NAND2_X1 U6316 ( .A1(n5674), .A2(n4874), .ZN(n4873) );
  CLKBUF_X1 U6317 ( .A(n6492), .Z(n4876) );
  MUX2_X1 U6318 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n6492), .Z(n5190) );
  MUX2_X1 U6319 ( .A(n10192), .B(n5318), .S(n6492), .Z(n5319) );
  MUX2_X1 U6320 ( .A(n10463), .B(n6544), .S(n6492), .Z(n5349) );
  MUX2_X1 U6321 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n4876), .Z(n5389) );
  MUX2_X1 U6322 ( .A(n6777), .B(n6775), .S(n4876), .Z(n5420) );
  MUX2_X1 U6323 ( .A(n10454), .B(n6875), .S(n4876), .Z(n5470) );
  MUX2_X1 U6324 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n4876), .Z(n5541) );
  MUX2_X1 U6325 ( .A(n10389), .B(n7150), .S(n4876), .Z(n5565) );
  MUX2_X1 U6326 ( .A(n7303), .B(n7331), .S(n4876), .Z(n5628) );
  MUX2_X1 U6327 ( .A(n10465), .B(n7485), .S(n4876), .Z(n5653) );
  MUX2_X1 U6328 ( .A(n10437), .B(n7619), .S(n4876), .Z(n5694) );
  MUX2_X1 U6329 ( .A(n10272), .B(n7728), .S(n4876), .Z(n5742) );
  MUX2_X1 U6330 ( .A(n8854), .B(n8609), .S(n4876), .Z(n7721) );
  NAND2_X1 U6331 ( .A1(n4878), .A2(n4557), .ZN(n5631) );
  AND3_X2 U6332 ( .A1(n5092), .A2(n5091), .A3(n5223), .ZN(n5497) );
  AND2_X2 U6333 ( .A1(n5090), .A2(n5157), .ZN(n5223) );
  AND4_X2 U6334 ( .A1(n5089), .A2(n5087), .A3(n5298), .A4(n5088), .ZN(n5091)
         );
  AND2_X2 U6335 ( .A1(n5498), .A2(n5086), .ZN(n5092) );
  NOR2_X2 U6336 ( .A1(n8450), .A2(n8554), .ZN(n8433) );
  INV_X1 U6337 ( .A(n4897), .ZN(n4896) );
  NAND2_X1 U6338 ( .A1(n6556), .A2(n6492), .ZN(n5194) );
  NAND2_X1 U6339 ( .A1(n8263), .A2(n4485), .ZN(n4906) );
  INV_X1 U6340 ( .A(n8420), .ZN(n4909) );
  NAND2_X1 U6341 ( .A1(n4914), .A2(n8272), .ZN(n8395) );
  NAND2_X1 U6342 ( .A1(n4921), .A2(n4923), .ZN(n7374) );
  OAI21_X1 U6343 ( .B1(n8585), .B2(n10062), .A(n4929), .ZN(P2_U3549) );
  NAND2_X1 U6344 ( .A1(n6833), .A2(n4934), .ZN(n4932) );
  INV_X1 U6345 ( .A(n6473), .ZN(n4931) );
  NAND2_X1 U6346 ( .A1(n4932), .A2(n4930), .ZN(n5315) );
  INV_X1 U6347 ( .A(n7804), .ZN(n4941) );
  NAND2_X1 U6348 ( .A1(n8100), .A2(n4945), .ZN(n4944) );
  INV_X1 U6349 ( .A(n6816), .ZN(n4953) );
  NAND2_X1 U6350 ( .A1(n7805), .A2(n4949), .ZN(n4952) );
  NAND2_X1 U6351 ( .A1(n6814), .A2(n5210), .ZN(n6824) );
  NAND2_X1 U6352 ( .A1(n7805), .A2(n5171), .ZN(n6809) );
  NAND2_X1 U6353 ( .A1(n7080), .A2(n4961), .ZN(n4964) );
  INV_X1 U6354 ( .A(n7084), .ZN(n4967) );
  NAND2_X1 U6355 ( .A1(n8090), .A2(n4968), .ZN(n5539) );
  INV_X1 U6356 ( .A(n5109), .ZN(n5108) );
  NAND4_X1 U6357 ( .A1(n5092), .A2(n5091), .A3(n4974), .A4(n5223), .ZN(n5109)
         );
  OAI21_X1 U6358 ( .B1(n6852), .B2(n4975), .A(n6851), .ZN(n6857) );
  NAND3_X1 U6359 ( .A1(n4977), .A2(n4976), .A3(n7035), .ZN(n6056) );
  NAND2_X1 U6360 ( .A1(n7092), .A2(n4979), .ZN(n4977) );
  INV_X1 U6361 ( .A(n8622), .ZN(n4981) );
  NAND2_X1 U6362 ( .A1(n7579), .A2(n4482), .ZN(n4992) );
  NAND2_X1 U6363 ( .A1(n4997), .A2(n4998), .ZN(n8717) );
  INV_X1 U6364 ( .A(n4999), .ZN(n8665) );
  INV_X1 U6365 ( .A(n8606), .ZN(n5006) );
  NAND2_X1 U6366 ( .A1(n7814), .A2(n5010), .ZN(n5009) );
  NAND3_X1 U6367 ( .A1(n5018), .A2(n5016), .A3(n7863), .ZN(n6971) );
  NAND3_X1 U6368 ( .A1(n7858), .A2(n5019), .A3(n6995), .ZN(n5018) );
  NAND3_X1 U6369 ( .A1(n5093), .A2(n5497), .A3(n5118), .ZN(n5095) );
  NAND2_X1 U6370 ( .A1(n7255), .A2(n7306), .ZN(n7308) );
  NAND2_X1 U6371 ( .A1(n7254), .A2(n7253), .ZN(n7255) );
  XNOR2_X2 U6372 ( .A(n5891), .B(n5857), .ZN(n9613) );
  NAND2_X1 U6373 ( .A1(n7605), .A2(n5044), .ZN(n5043) );
  AOI21_X2 U6374 ( .B1(n5053), .B2(n5052), .A(n5051), .ZN(n7695) );
  OAI21_X1 U6375 ( .B1(n9311), .B2(n5056), .A(n5054), .ZN(n9261) );
  NOR2_X1 U6376 ( .A1(n9261), .A2(n5062), .ZN(n9108) );
  NAND2_X1 U6377 ( .A1(n5065), .A2(n5063), .ZN(n9726) );
  NAND2_X1 U6378 ( .A1(n9245), .A2(n5068), .ZN(n5067) );
  NAND2_X1 U6379 ( .A1(n5071), .A2(n5072), .ZN(n9763) );
  AND2_X1 U6380 ( .A1(n8962), .A2(n7309), .ZN(n5071) );
  OAI21_X1 U6381 ( .B1(n9156), .B2(n5075), .A(n5073), .ZN(n9124) );
  NAND2_X1 U6382 ( .A1(n9156), .A2(n9155), .ZN(n9154) );
  XNOR2_X2 U6383 ( .A(n5686), .B(n5684), .ZN(n8100) );
  CLKBUF_X1 U6384 ( .A(n8106), .Z(n8108) );
  INV_X1 U6385 ( .A(n5930), .ZN(n5993) );
  OR2_X1 U6386 ( .A1(n5930), .A2(n5866), .ZN(n5867) );
  NAND2_X1 U6387 ( .A1(n5489), .A2(n4518), .ZN(n5514) );
  OR2_X1 U6388 ( .A1(n8754), .A2(n9892), .ZN(n5935) );
  NAND2_X1 U6389 ( .A1(n5138), .A2(n5139), .ZN(n5149) );
  NAND2_X1 U6390 ( .A1(n7839), .A2(n7838), .ZN(n8028) );
  NAND2_X2 U6391 ( .A1(n5670), .A2(n5669), .ZN(n5686) );
  INV_X1 U6392 ( .A(n5938), .ZN(n5846) );
  OR2_X1 U6393 ( .A1(n9813), .A2(n6345), .ZN(n5924) );
  CLKBUF_X1 U6394 ( .A(n9311), .Z(n9312) );
  INV_X1 U6395 ( .A(n5576), .ZN(n5254) );
  INV_X1 U6396 ( .A(n6914), .ZN(n9967) );
  INV_X1 U6397 ( .A(n7929), .ZN(n7813) );
  NOR2_X1 U6398 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n5079) );
  INV_X1 U6399 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5192) );
  AND2_X1 U6400 ( .A1(n5440), .A2(n5422), .ZN(n5080) );
  INV_X1 U6401 ( .A(n7528), .ZN(n8008) );
  OR2_X1 U6402 ( .A1(n6581), .A2(n7776), .ZN(n5081) );
  INV_X1 U6403 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5841) );
  INV_X1 U6404 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5851) );
  INV_X1 U6405 ( .A(n5701), .ZN(n5699) );
  INV_X1 U6406 ( .A(n5451), .ZN(n5450) );
  INV_X1 U6407 ( .A(n7083), .ZN(n5340) );
  INV_X1 U6408 ( .A(n5481), .ZN(n5479) );
  NAND2_X1 U6409 ( .A1(n5699), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5724) );
  INV_X1 U6410 ( .A(n5376), .ZN(n5374) );
  INV_X1 U6411 ( .A(n5229), .ZN(n5227) );
  INV_X1 U6412 ( .A(n6030), .ZN(n6031) );
  INV_X1 U6413 ( .A(n7347), .ZN(n6104) );
  INV_X1 U6414 ( .A(n6353), .ZN(n6351) );
  INV_X1 U6415 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6087) );
  INV_X1 U6416 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6259) );
  INV_X1 U6417 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6157) );
  INV_X1 U6418 ( .A(n5287), .ZN(n5288) );
  INV_X1 U6419 ( .A(n5213), .ZN(n5216) );
  NAND2_X1 U6420 ( .A1(n5450), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5481) );
  NOR2_X1 U6421 ( .A1(n8297), .A2(n8129), .ZN(n5819) );
  NAND2_X1 U6422 ( .A1(n5149), .A2(n5140), .ZN(n7711) );
  NAND2_X1 U6423 ( .A1(n5528), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5549) );
  INV_X1 U6424 ( .A(n7388), .ZN(n5415) );
  NAND2_X1 U6425 ( .A1(n5637), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5658) );
  OR2_X1 U6426 ( .A1(n5678), .A2(n10253), .ZN(n5701) );
  NAND2_X1 U6427 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5229) );
  AND2_X1 U6428 ( .A1(n5764), .A2(n5821), .ZN(n8306) );
  INV_X1 U6429 ( .A(n7882), .ZN(n6916) );
  OR2_X1 U6430 ( .A1(n6109), .A2(n7441), .ZN(n6126) );
  NAND2_X1 U6431 ( .A1(n6351), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6371) );
  OR2_X1 U6432 ( .A1(n6293), .A2(n8678), .ZN(n6311) );
  OR2_X1 U6433 ( .A1(n6164), .A2(n6163), .ZN(n6182) );
  INV_X1 U6434 ( .A(n9155), .ZN(n9150) );
  INV_X1 U6435 ( .A(n9560), .ZN(n7606) );
  OR2_X1 U6436 ( .A1(n6088), .A2(n6087), .ZN(n6109) );
  INV_X1 U6437 ( .A(n9847), .ZN(n7412) );
  NAND2_X1 U6438 ( .A1(n5470), .A2(n5469), .ZN(n5490) );
  OR2_X1 U6439 ( .A1(n5304), .A2(n10250), .ZN(n5329) );
  OR2_X1 U6440 ( .A1(n5505), .A2(n10436), .ZN(n5529) );
  INV_X1 U6441 ( .A(n8511), .ZN(n8309) );
  INV_X1 U6442 ( .A(n8438), .ZN(n7817) );
  AND2_X1 U6443 ( .A1(n7906), .A2(n7908), .ZN(n7273) );
  INV_X1 U6444 ( .A(n8009), .ZN(n7921) );
  OR2_X1 U6445 ( .A1(n6514), .A2(n5820), .ZN(n8428) );
  NOR2_X1 U6446 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5122) );
  INV_X1 U6447 ( .A(n5497), .ZN(n5524) );
  OR2_X1 U6448 ( .A1(n6386), .A2(n6385), .ZN(n6455) );
  OR2_X1 U6449 ( .A1(n5929), .A2(n7144), .ZN(n5916) );
  INV_X1 U6450 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7441) );
  INV_X1 U6451 ( .A(n9400), .ZN(n9256) );
  INV_X1 U6452 ( .A(n9406), .ZN(n9272) );
  INV_X1 U6453 ( .A(n9031), .ZN(n8652) );
  AOI21_X1 U6454 ( .B1(n7360), .B2(n7359), .A(n7358), .ZN(n7361) );
  OR2_X1 U6455 ( .A1(n9797), .A2(n6442), .ZN(n9869) );
  INV_X1 U6456 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6437) );
  AND2_X1 U6457 ( .A1(n5609), .A2(n5594), .ZN(n5607) );
  AND2_X1 U6458 ( .A1(n5521), .A2(n5496), .ZN(n5519) );
  INV_X1 U6459 ( .A(n8123), .ZN(n8143) );
  AND2_X1 U6460 ( .A1(n5645), .A2(n5644), .ZN(n8150) );
  AND2_X1 U6461 ( .A1(n6558), .A2(n6557), .ZN(n9904) );
  AND2_X1 U6462 ( .A1(n8445), .A2(n7940), .ZN(n8465) );
  OR2_X1 U6463 ( .A1(n8020), .A2(n6697), .ZN(n9938) );
  INV_X1 U6464 ( .A(n9951), .ZN(n8490) );
  OR2_X1 U6465 ( .A1(n7991), .A2(n4939), .ZN(n10034) );
  AND2_X1 U6466 ( .A1(n5827), .A2(n5828), .ZN(n10020) );
  OR3_X1 U6467 ( .A1(n6922), .A2(n6691), .A3(n6923), .ZN(n6705) );
  AND2_X1 U6468 ( .A1(n6401), .A2(n6400), .ZN(n6416) );
  INV_X1 U6469 ( .A(n8735), .ZN(n8725) );
  INV_X1 U6470 ( .A(n8712), .ZN(n8732) );
  AND4_X1 U6471 ( .A1(n6271), .A2(n6270), .A3(n6269), .A4(n6268), .ZN(n9424)
         );
  AND2_X1 U6472 ( .A1(n8906), .A2(n8909), .ZN(n8971) );
  INV_X1 U6473 ( .A(n9331), .ZN(n9767) );
  INV_X1 U6474 ( .A(n9819), .ZN(n8698) );
  AND2_X1 U6475 ( .A1(n9810), .A2(n6466), .ZN(n9804) );
  AND2_X1 U6476 ( .A1(n8864), .A2(n7234), .ZN(n9875) );
  OR3_X1 U6477 ( .A1(n6421), .A2(n6420), .A3(n7635), .ZN(n7130) );
  XNOR2_X1 U6478 ( .A(n5190), .B(n5185), .ZN(n5188) );
  OR2_X1 U6479 ( .A1(n8141), .A2(n8426), .ZN(n8129) );
  OR3_X1 U6480 ( .A1(n5817), .A2(n10002), .A3(n6552), .ZN(n8145) );
  INV_X1 U6481 ( .A(n8370), .ZN(n8277) );
  AND2_X1 U6482 ( .A1(n8350), .A2(n8349), .ZN(n8531) );
  OR2_X1 U6483 ( .A1(n6927), .A2(n7839), .ZN(n9948) );
  OR2_X1 U6484 ( .A1(n6705), .A2(n6921), .ZN(n10062) );
  OR2_X1 U6485 ( .A1(n6705), .A2(n6692), .ZN(n10042) );
  OR2_X1 U6486 ( .A1(n9956), .A2(n9955), .ZN(n9959) );
  OR2_X1 U6487 ( .A1(n6465), .A2(n6440), .ZN(n8712) );
  INV_X1 U6488 ( .A(n8710), .ZN(n8743) );
  NAND2_X1 U6489 ( .A1(n6393), .A2(n6392), .ZN(n9186) );
  OR3_X1 U6490 ( .A1(n6285), .A2(n6284), .A3(n6283), .ZN(n9415) );
  AND2_X1 U6491 ( .A1(n7134), .A2(n9319), .ZN(n9779) );
  OR2_X1 U6492 ( .A1(n9807), .A2(n7305), .ZN(n9331) );
  INV_X1 U6493 ( .A(n9222), .ZN(n9807) );
  INV_X1 U6494 ( .A(n9351), .ZN(n9434) );
  INV_X1 U6495 ( .A(n7672), .ZN(n8788) );
  INV_X1 U6496 ( .A(n9888), .ZN(n9887) );
  INV_X1 U6497 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10463) );
  NOR2_X1 U6498 ( .A1(n10119), .A2(n10118), .ZN(n10117) );
  INV_X1 U6499 ( .A(n9036), .ZN(P1_U4006) );
  INV_X1 U6500 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5082) );
  NAND4_X1 U6501 ( .A1(n5083), .A2(n5103), .A3(n5807), .A4(n5082), .ZN(n5085)
         );
  INV_X1 U6502 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5110) );
  INV_X1 U6503 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5106) );
  INV_X1 U6504 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5781) );
  NAND4_X1 U6505 ( .A1(n5110), .A2(n5106), .A3(n5112), .A4(n5781), .ZN(n5084)
         );
  AND3_X2 U6506 ( .A1(n5445), .A2(n5442), .A3(n5475), .ZN(n5498) );
  NOR2_X1 U6507 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5086) );
  NOR2_X2 U6508 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5298) );
  NOR2_X1 U6509 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5089) );
  NOR2_X1 U6510 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5090) );
  INV_X1 U6511 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5118) );
  INV_X1 U6512 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8600) );
  NAND2_X1 U6513 ( .A1(n5095), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5096) );
  INV_X1 U6514 ( .A(n5098), .ZN(n8610) );
  INV_X1 U6515 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5097) );
  OR2_X1 U6516 ( .A1(n5254), .A2(n5097), .ZN(n5102) );
  INV_X1 U6517 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6569) );
  OR2_X1 U6518 ( .A1(n5199), .A2(n6569), .ZN(n5101) );
  INV_X1 U6519 ( .A(n5579), .ZN(n5150) );
  NAND2_X1 U6520 ( .A1(n5150), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5100) );
  INV_X1 U6521 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10448) );
  OR2_X1 U6522 ( .A1(n5726), .A2(n10448), .ZN(n5099) );
  NOR2_X1 U6523 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5104) );
  NAND2_X1 U6524 ( .A1(n5108), .A2(n5104), .ZN(n5105) );
  INV_X1 U6525 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5782) );
  XNOR2_X2 U6526 ( .A(n5778), .B(n5782), .ZN(n5827) );
  NAND2_X1 U6527 ( .A1(n5105), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5107) );
  XNOR2_X1 U6528 ( .A(n5107), .B(n5106), .ZN(n7828) );
  NAND2_X1 U6529 ( .A1(n5113), .A2(n5110), .ZN(n5115) );
  NAND2_X1 U6530 ( .A1(n5115), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5111) );
  INV_X1 U6531 ( .A(n5113), .ZN(n5114) );
  NAND2_X1 U6532 ( .A1(n5114), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n5116) );
  NAND2_X1 U6533 ( .A1(n7991), .A2(n7828), .ZN(n5117) );
  INV_X1 U6534 ( .A(n5827), .ZN(n8030) );
  INV_X1 U6535 ( .A(n7828), .ZN(n8023) );
  NAND2_X1 U6536 ( .A1(n8023), .A2(n7249), .ZN(n6946) );
  INV_X2 U6537 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5124) );
  NAND2_X2 U6538 ( .A1(n5125), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5131) );
  INV_X1 U6539 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5127) );
  INV_X1 U6540 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5126) );
  NAND2_X1 U6541 ( .A1(n5127), .A2(n5126), .ZN(n5129) );
  NAND2_X2 U6542 ( .A1(n5129), .A2(n5128), .ZN(n5130) );
  NAND2_X4 U6543 ( .A1(n5131), .A2(n5130), .ZN(n6492) );
  AND2_X1 U6544 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5132) );
  NAND3_X1 U6545 ( .A1(n6492), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n5133) );
  INV_X1 U6546 ( .A(SI_1_), .ZN(n5134) );
  MUX2_X1 U6547 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4877), .Z(n5159) );
  XNOR2_X1 U6548 ( .A(n5160), .B(n5159), .ZN(n6498) );
  INV_X1 U6549 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6487) );
  OR2_X1 U6550 ( .A1(n5196), .A2(n6487), .ZN(n5135) );
  OAI211_X2 U6551 ( .C1(n6556), .C2(n9506), .A(n5136), .B(n5135), .ZN(n7716)
         );
  XNOR2_X1 U6552 ( .A(n5137), .B(n7716), .ZN(n5139) );
  NAND2_X1 U6553 ( .A1(n5150), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5146) );
  INV_X1 U6554 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5141) );
  INV_X1 U6555 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5142) );
  OR2_X1 U6556 ( .A1(n5199), .A2(n5142), .ZN(n5144) );
  INV_X1 U6557 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6984) );
  OR2_X1 U6558 ( .A1(n5726), .A2(n6984), .ZN(n5143) );
  NAND2_X1 U6559 ( .A1(n6492), .A2(SI_0_), .ZN(n5147) );
  XNOR2_X1 U6560 ( .A(n5147), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8613) );
  MUX2_X1 U6561 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8613), .S(n6556), .Z(n9963) );
  INV_X1 U6562 ( .A(n9963), .ZN(n6779) );
  OAI22_X1 U6563 ( .A1(n6934), .A2(n5771), .B1(n9963), .B2(n5772), .ZN(n7712)
         );
  OR2_X1 U6564 ( .A1(n7711), .A2(n7712), .ZN(n7714) );
  NAND2_X1 U6565 ( .A1(n7714), .A2(n5149), .ZN(n7806) );
  NAND2_X1 U6566 ( .A1(n5150), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5156) );
  INV_X1 U6567 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5151) );
  OR2_X1 U6568 ( .A1(n5199), .A2(n5151), .ZN(n5155) );
  INV_X1 U6569 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5152) );
  INV_X1 U6570 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10365) );
  NOR2_X1 U6571 ( .A1(n6937), .A2(n5771), .ZN(n5166) );
  OR2_X1 U6572 ( .A1(n5157), .A2(n5399), .ZN(n5158) );
  XNOR2_X1 U6573 ( .A(n5158), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9526) );
  INV_X1 U6574 ( .A(n9526), .ZN(n6488) );
  NAND2_X1 U6575 ( .A1(n5160), .A2(n5159), .ZN(n5163) );
  NAND2_X1 U6576 ( .A1(n5161), .A2(SI_1_), .ZN(n5162) );
  NAND2_X1 U6577 ( .A1(n5163), .A2(n5162), .ZN(n5181) );
  INV_X1 U6578 ( .A(SI_2_), .ZN(n10398) );
  XNOR2_X1 U6579 ( .A(n5181), .B(n5180), .ZN(n6493) );
  OR2_X1 U6580 ( .A1(n5194), .A2(n6493), .ZN(n5165) );
  INV_X1 U6581 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6489) );
  OR2_X1 U6582 ( .A1(n5196), .A2(n6489), .ZN(n5164) );
  XNOR2_X1 U6583 ( .A(n5772), .B(n6914), .ZN(n5167) );
  NAND2_X1 U6584 ( .A1(n5166), .A2(n5167), .ZN(n5170) );
  INV_X1 U6585 ( .A(n5166), .ZN(n5169) );
  INV_X1 U6586 ( .A(n5167), .ZN(n5168) );
  NAND2_X1 U6587 ( .A1(n5169), .A2(n5168), .ZN(n5171) );
  AND2_X1 U6588 ( .A1(n5170), .A2(n5171), .ZN(n7807) );
  NAND2_X1 U6589 ( .A1(n7806), .A2(n7807), .ZN(n7805) );
  NAND2_X1 U6590 ( .A1(n5822), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5177) );
  INV_X1 U6591 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5172) );
  OR2_X1 U6592 ( .A1(n5199), .A2(n5172), .ZN(n5176) );
  INV_X1 U6593 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5173) );
  OR2_X1 U6594 ( .A1(n7827), .A2(n5173), .ZN(n5175) );
  OR2_X1 U6595 ( .A1(n5726), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5174) );
  AND4_X1 U6596 ( .A1(n5177), .A2(n5176), .A3(n5175), .A4(n5174), .ZN(n7803)
         );
  OR2_X1 U6597 ( .A1(n7803), .A2(n5771), .ZN(n5186) );
  NAND2_X1 U6598 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5178), .ZN(n5179) );
  XNOR2_X1 U6599 ( .A(n5179), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6600) );
  INV_X1 U6600 ( .A(n6600), .ZN(n6490) );
  NAND2_X1 U6601 ( .A1(n5182), .A2(SI_2_), .ZN(n5183) );
  INV_X1 U6602 ( .A(SI_3_), .ZN(n5185) );
  INV_X1 U6603 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6491) );
  XNOR2_X1 U6604 ( .A(n5137), .B(n6999), .ZN(n5187) );
  XNOR2_X1 U6605 ( .A(n5186), .B(n5187), .ZN(n6810) );
  NAND2_X1 U6606 ( .A1(n5190), .A2(SI_3_), .ZN(n5212) );
  NAND2_X1 U6607 ( .A1(n5219), .A2(n5212), .ZN(n5193) );
  XNOR2_X1 U6608 ( .A(n5193), .B(n5213), .ZN(n5974) );
  NAND2_X1 U6609 ( .A1(n5974), .A2(n5220), .ZN(n5198) );
  OR2_X1 U6610 ( .A1(n5223), .A2(n5399), .ZN(n5195) );
  XNOR2_X1 U6611 ( .A(n5195), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6614) );
  NAND2_X1 U6612 ( .A1(n5568), .A2(n6614), .ZN(n5197) );
  XNOR2_X1 U6613 ( .A(n9981), .B(n5772), .ZN(n5205) );
  NAND2_X1 U6614 ( .A1(n7823), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5204) );
  INV_X1 U6615 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6588) );
  OR2_X1 U6616 ( .A1(n5579), .A2(n6588), .ZN(n5203) );
  OAI21_X1 U6617 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n5229), .ZN(n9925) );
  OR2_X1 U6618 ( .A1(n5726), .A2(n9925), .ZN(n5202) );
  INV_X1 U6619 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5200) );
  OR2_X1 U6620 ( .A1(n7827), .A2(n5200), .ZN(n5201) );
  NAND4_X1 U6621 ( .A1(n5204), .A2(n5203), .A3(n5202), .A4(n5201), .ZN(n8164)
         );
  NAND2_X1 U6622 ( .A1(n8164), .A2(n7839), .ZN(n5206) );
  NAND2_X1 U6623 ( .A1(n5205), .A2(n5206), .ZN(n5210) );
  INV_X1 U6624 ( .A(n5205), .ZN(n5208) );
  INV_X1 U6625 ( .A(n5206), .ZN(n5207) );
  NAND2_X1 U6626 ( .A1(n5208), .A2(n5207), .ZN(n5209) );
  NAND2_X1 U6627 ( .A1(n5210), .A2(n5209), .ZN(n6816) );
  NAND2_X1 U6628 ( .A1(n5211), .A2(SI_4_), .ZN(n5214) );
  AND2_X1 U6629 ( .A1(n5212), .A2(n5214), .ZN(n5218) );
  INV_X1 U6630 ( .A(n5214), .ZN(n5215) );
  MUX2_X1 U6631 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n7832), .Z(n5245) );
  XNOR2_X1 U6632 ( .A(n5244), .B(n5242), .ZN(n6001) );
  NAND2_X1 U6633 ( .A1(n6001), .A2(n5220), .ZN(n5225) );
  INV_X2 U6634 ( .A(n5221), .ZN(n5569) );
  INV_X1 U6635 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5222) );
  NAND2_X1 U6636 ( .A1(n5223), .A2(n5222), .ZN(n5300) );
  NAND2_X1 U6637 ( .A1(n5300), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5247) );
  XNOR2_X1 U6638 ( .A(n5247), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6630) );
  AOI22_X1 U6639 ( .A1(n5569), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n5568), .B2(
        n6630), .ZN(n5224) );
  XNOR2_X1 U6640 ( .A(n9989), .B(n5772), .ZN(n5236) );
  NAND2_X1 U6641 ( .A1(n7823), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5235) );
  INV_X1 U6642 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5226) );
  OR2_X1 U6643 ( .A1(n5579), .A2(n5226), .ZN(n5234) );
  INV_X1 U6644 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5228) );
  NAND2_X1 U6645 ( .A1(n5229), .A2(n5228), .ZN(n5230) );
  NAND2_X1 U6646 ( .A1(n5252), .A2(n5230), .ZN(n7010) );
  OR2_X1 U6647 ( .A1(n5726), .A2(n7010), .ZN(n5233) );
  INV_X1 U6648 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5231) );
  OR2_X1 U6649 ( .A1(n7827), .A2(n5231), .ZN(n5232) );
  NAND4_X1 U6650 ( .A1(n5235), .A2(n5234), .A3(n5233), .A4(n5232), .ZN(n9918)
         );
  NAND2_X1 U6651 ( .A1(n9918), .A2(n7839), .ZN(n5237) );
  NAND2_X1 U6652 ( .A1(n5236), .A2(n5237), .ZN(n5241) );
  INV_X1 U6653 ( .A(n5236), .ZN(n5239) );
  INV_X1 U6654 ( .A(n5237), .ZN(n5238) );
  NAND2_X1 U6655 ( .A1(n5239), .A2(n5238), .ZN(n5240) );
  AND2_X1 U6656 ( .A1(n5241), .A2(n5240), .ZN(n6825) );
  NAND2_X1 U6657 ( .A1(n6824), .A2(n6825), .ZN(n6823) );
  NAND2_X1 U6658 ( .A1(n5245), .A2(SI_5_), .ZN(n5246) );
  MUX2_X1 U6659 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7832), .Z(n5269) );
  XNOR2_X1 U6660 ( .A(n5268), .B(n5266), .ZN(n6506) );
  NAND2_X1 U6661 ( .A1(n6506), .A2(n5220), .ZN(n5250) );
  INV_X1 U6662 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5297) );
  NAND2_X1 U6663 ( .A1(n5247), .A2(n5297), .ZN(n5248) );
  NAND2_X1 U6664 ( .A1(n5248), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5271) );
  XNOR2_X1 U6665 ( .A(n5271), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6665) );
  AOI22_X1 U6666 ( .A1(n5569), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n5568), .B2(
        n6665), .ZN(n5249) );
  NAND2_X1 U6667 ( .A1(n5250), .A2(n5249), .ZN(n7884) );
  XNOR2_X1 U6668 ( .A(n7884), .B(n5137), .ZN(n5260) );
  NAND2_X1 U6669 ( .A1(n5822), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5259) );
  INV_X1 U6670 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6979) );
  OR2_X1 U6671 ( .A1(n5199), .A2(n6979), .ZN(n5258) );
  INV_X1 U6672 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10275) );
  NAND2_X1 U6673 ( .A1(n5252), .A2(n10275), .ZN(n5253) );
  NAND2_X1 U6674 ( .A1(n5279), .A2(n5253), .ZN(n6975) );
  OR2_X1 U6675 ( .A1(n5726), .A2(n6975), .ZN(n5257) );
  INV_X1 U6676 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5255) );
  OR2_X1 U6677 ( .A1(n7827), .A2(n5255), .ZN(n5256) );
  NAND4_X1 U6678 ( .A1(n5259), .A2(n5258), .A3(n5257), .A4(n5256), .ZN(n8163)
         );
  NAND2_X1 U6679 ( .A1(n8163), .A2(n7839), .ZN(n5261) );
  NAND2_X1 U6680 ( .A1(n5260), .A2(n5261), .ZN(n5265) );
  INV_X1 U6681 ( .A(n5260), .ZN(n5263) );
  INV_X1 U6682 ( .A(n5261), .ZN(n5262) );
  NAND2_X1 U6683 ( .A1(n5263), .A2(n5262), .ZN(n5264) );
  AND2_X1 U6684 ( .A1(n5265), .A2(n5264), .ZN(n6834) );
  MUX2_X1 U6685 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7832), .Z(n5290) );
  XNOR2_X1 U6686 ( .A(n5289), .B(n5287), .ZN(n6510) );
  NAND2_X1 U6687 ( .A1(n6510), .A2(n5220), .ZN(n5275) );
  INV_X1 U6688 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5270) );
  NAND2_X1 U6689 ( .A1(n5271), .A2(n5270), .ZN(n5272) );
  NAND2_X1 U6690 ( .A1(n5272), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5273) );
  XNOR2_X1 U6691 ( .A(n5273), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6795) );
  AOI22_X1 U6692 ( .A1(n5569), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5568), .B2(
        n6795), .ZN(n5274) );
  NAND2_X1 U6693 ( .A1(n5275), .A2(n5274), .ZN(n10001) );
  XNOR2_X1 U6694 ( .A(n10001), .B(n5772), .ZN(n5286) );
  NAND2_X1 U6695 ( .A1(n5822), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5284) );
  INV_X1 U6696 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5276) );
  OR2_X1 U6697 ( .A1(n7827), .A2(n5276), .ZN(n5283) );
  INV_X1 U6698 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U6699 ( .A1(n5279), .A2(n5278), .ZN(n5280) );
  NAND2_X1 U6700 ( .A1(n5304), .A2(n5280), .ZN(n6928) );
  OR2_X1 U6701 ( .A1(n5726), .A2(n6928), .ZN(n5282) );
  INV_X1 U6702 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6929) );
  OR2_X1 U6703 ( .A1(n5199), .A2(n6929), .ZN(n5281) );
  NOR2_X1 U6704 ( .A1(n7062), .A2(n5771), .ZN(n5285) );
  XNOR2_X1 U6705 ( .A(n5286), .B(n5285), .ZN(n6877) );
  NAND2_X1 U6706 ( .A1(n5289), .A2(n5288), .ZN(n5292) );
  NAND2_X1 U6707 ( .A1(n5290), .A2(SI_7_), .ZN(n5291) );
  MUX2_X1 U6708 ( .A(n6546), .B(n6528), .S(n7832), .Z(n5294) );
  INV_X1 U6709 ( .A(SI_8_), .ZN(n5293) );
  INV_X1 U6710 ( .A(n5294), .ZN(n5295) );
  NAND2_X1 U6711 ( .A1(n5295), .A2(SI_8_), .ZN(n5296) );
  XNOR2_X1 U6712 ( .A(n5317), .B(n5316), .ZN(n6518) );
  NAND2_X1 U6713 ( .A1(n6518), .A2(n5220), .ZN(n5303) );
  NAND2_X1 U6714 ( .A1(n5298), .A2(n5297), .ZN(n5299) );
  NAND2_X1 U6715 ( .A1(n5323), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5301) );
  XNOR2_X1 U6716 ( .A(n5301), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6866) );
  AOI22_X1 U6717 ( .A1(n5569), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5568), .B2(
        n6866), .ZN(n5302) );
  XNOR2_X1 U6718 ( .A(n7112), .B(n5137), .ZN(n5311) );
  NAND2_X1 U6719 ( .A1(n5822), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5310) );
  INV_X1 U6720 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7073) );
  OR2_X1 U6721 ( .A1(n5199), .A2(n7073), .ZN(n5309) );
  NAND2_X1 U6722 ( .A1(n5304), .A2(n10250), .ZN(n5305) );
  NAND2_X1 U6723 ( .A1(n5329), .A2(n5305), .ZN(n7072) );
  OR2_X1 U6724 ( .A1(n5726), .A2(n7072), .ZN(n5308) );
  INV_X1 U6725 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5306) );
  OR2_X1 U6726 ( .A1(n7827), .A2(n5306), .ZN(n5307) );
  NOR2_X1 U6727 ( .A1(n7177), .A2(n5771), .ZN(n5312) );
  XNOR2_X1 U6728 ( .A(n5311), .B(n5312), .ZN(n6473) );
  INV_X1 U6729 ( .A(n5311), .ZN(n5313) );
  NAND2_X1 U6730 ( .A1(n5313), .A2(n5312), .ZN(n5314) );
  NAND2_X1 U6731 ( .A1(n5315), .A2(n5314), .ZN(n7080) );
  NAND2_X1 U6732 ( .A1(n5347), .A2(n5343), .ZN(n5322) );
  INV_X1 U6733 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5318) );
  INV_X1 U6734 ( .A(SI_9_), .ZN(n10395) );
  NAND2_X1 U6735 ( .A1(n5319), .A2(n10395), .ZN(n5342) );
  INV_X1 U6736 ( .A(n5319), .ZN(n5320) );
  AND2_X1 U6737 ( .A1(n5342), .A2(n5344), .ZN(n5321) );
  NAND2_X1 U6738 ( .A1(n6529), .A2(n5220), .ZN(n5325) );
  NOR2_X1 U6739 ( .A1(n5323), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5398) );
  OR2_X1 U6740 ( .A1(n5398), .A2(n5399), .ZN(n5352) );
  XNOR2_X1 U6741 ( .A(n5352), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6962) );
  AOI22_X1 U6742 ( .A1(n5569), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5568), .B2(
        n6962), .ZN(n5324) );
  XNOR2_X1 U6743 ( .A(n10014), .B(n5137), .ZN(n5335) );
  NAND2_X1 U6744 ( .A1(n5822), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5334) );
  INV_X1 U6745 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5326) );
  OR2_X1 U6746 ( .A1(n7827), .A2(n5326), .ZN(n5333) );
  INV_X1 U6747 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5328) );
  NAND2_X1 U6748 ( .A1(n5329), .A2(n5328), .ZN(n5330) );
  NAND2_X1 U6749 ( .A1(n5356), .A2(n5330), .ZN(n7182) );
  OR2_X1 U6750 ( .A1(n5726), .A2(n7182), .ZN(n5332) );
  INV_X1 U6751 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7183) );
  OR2_X1 U6752 ( .A1(n5199), .A2(n7183), .ZN(n5331) );
  OR2_X1 U6753 ( .A1(n7114), .A2(n5771), .ZN(n5336) );
  NAND2_X1 U6754 ( .A1(n5335), .A2(n5336), .ZN(n5341) );
  INV_X1 U6755 ( .A(n5335), .ZN(n5338) );
  INV_X1 U6756 ( .A(n5336), .ZN(n5337) );
  NAND2_X1 U6757 ( .A1(n5338), .A2(n5337), .ZN(n5339) );
  NAND2_X1 U6758 ( .A1(n5341), .A2(n5339), .ZN(n7083) );
  INV_X1 U6759 ( .A(n5344), .ZN(n5345) );
  INV_X1 U6760 ( .A(SI_10_), .ZN(n5348) );
  INV_X1 U6761 ( .A(n5349), .ZN(n5350) );
  NAND2_X1 U6762 ( .A1(n5350), .A2(SI_10_), .ZN(n5351) );
  NAND2_X1 U6763 ( .A1(n6535), .A2(n5220), .ZN(n5355) );
  INV_X1 U6764 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5395) );
  NAND2_X1 U6765 ( .A1(n5352), .A2(n5395), .ZN(n5353) );
  NAND2_X1 U6766 ( .A1(n5353), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5369) );
  XNOR2_X1 U6767 ( .A(n5369), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7050) );
  AOI22_X1 U6768 ( .A1(n5569), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5568), .B2(
        n7050), .ZN(n5354) );
  NAND2_X1 U6769 ( .A1(n5355), .A2(n5354), .ZN(n7119) );
  XNOR2_X1 U6770 ( .A(n7119), .B(n5772), .ZN(n5363) );
  NAND2_X1 U6771 ( .A1(n5822), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5362) );
  INV_X1 U6772 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7117) );
  OR2_X1 U6773 ( .A1(n5199), .A2(n7117), .ZN(n5361) );
  INV_X1 U6774 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6957) );
  NAND2_X1 U6775 ( .A1(n5356), .A2(n6957), .ZN(n5357) );
  NAND2_X1 U6776 ( .A1(n5376), .A2(n5357), .ZN(n8057) );
  OR2_X1 U6777 ( .A1(n5726), .A2(n8057), .ZN(n5360) );
  INV_X1 U6778 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5358) );
  OR2_X1 U6779 ( .A1(n7827), .A2(n5358), .ZN(n5359) );
  NOR2_X1 U6780 ( .A1(n8158), .A2(n5771), .ZN(n5364) );
  XNOR2_X1 U6781 ( .A(n5363), .B(n5364), .ZN(n8053) );
  INV_X1 U6782 ( .A(n5363), .ZN(n5366) );
  INV_X1 U6783 ( .A(n5364), .ZN(n5365) );
  INV_X1 U6784 ( .A(SI_11_), .ZN(n5368) );
  XNOR2_X1 U6785 ( .A(n5390), .B(n5388), .ZN(n6548) );
  NAND2_X1 U6786 ( .A1(n6548), .A2(n5220), .ZN(n5373) );
  INV_X1 U6787 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5396) );
  NAND2_X1 U6788 ( .A1(n5369), .A2(n5396), .ZN(n5370) );
  NAND2_X1 U6789 ( .A1(n5370), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5371) );
  XNOR2_X1 U6790 ( .A(n5371), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7242) );
  AOI22_X1 U6791 ( .A1(n5569), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5568), .B2(
        n7242), .ZN(n5372) );
  NAND2_X1 U6792 ( .A1(n5373), .A2(n5372), .ZN(n7372) );
  XNOR2_X1 U6793 ( .A(n7372), .B(n5137), .ZN(n5383) );
  NAND2_X1 U6794 ( .A1(n5822), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5382) );
  INV_X1 U6795 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7277) );
  OR2_X1 U6796 ( .A1(n5199), .A2(n7277), .ZN(n5381) );
  INV_X1 U6797 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5375) );
  NAND2_X1 U6798 ( .A1(n5376), .A2(n5375), .ZN(n5377) );
  NAND2_X1 U6799 ( .A1(n5403), .A2(n5377), .ZN(n7276) );
  OR2_X1 U6800 ( .A1(n5726), .A2(n7276), .ZN(n5380) );
  INV_X1 U6801 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5378) );
  OR2_X1 U6802 ( .A1(n7827), .A2(n5378), .ZN(n5379) );
  NOR2_X1 U6803 ( .A1(n7392), .A2(n5771), .ZN(n5384) );
  XNOR2_X1 U6804 ( .A(n5383), .B(n5384), .ZN(n7204) );
  NAND2_X1 U6805 ( .A1(n7205), .A2(n7204), .ZN(n5387) );
  INV_X1 U6806 ( .A(n5383), .ZN(n5385) );
  NAND2_X1 U6807 ( .A1(n5385), .A2(n5384), .ZN(n5386) );
  NAND2_X1 U6808 ( .A1(n5387), .A2(n5386), .ZN(n7389) );
  INV_X1 U6809 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6673) );
  INV_X1 U6810 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6675) );
  MUX2_X1 U6811 ( .A(n6673), .B(n6675), .S(n7832), .Z(n5391) );
  INV_X1 U6812 ( .A(SI_12_), .ZN(n10363) );
  INV_X1 U6813 ( .A(n5391), .ZN(n5392) );
  NAND2_X1 U6814 ( .A1(n5392), .A2(SI_12_), .ZN(n5393) );
  XNOR2_X1 U6815 ( .A(n5419), .B(n5418), .ZN(n6672) );
  NAND2_X1 U6816 ( .A1(n6672), .A2(n5220), .ZN(n5402) );
  INV_X1 U6817 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5394) );
  AND3_X1 U6818 ( .A1(n5396), .A2(n5395), .A3(n5394), .ZN(n5397) );
  AND2_X1 U6819 ( .A1(n5398), .A2(n5397), .ZN(n5424) );
  OR2_X1 U6820 ( .A1(n5424), .A2(n5399), .ZN(n5400) );
  XNOR2_X1 U6821 ( .A(n5400), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7283) );
  AOI22_X1 U6822 ( .A1(n5569), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5568), .B2(
        n7283), .ZN(n5401) );
  XNOR2_X1 U6823 ( .A(n7424), .B(n5137), .ZN(n5410) );
  NAND2_X1 U6824 ( .A1(n7823), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5409) );
  INV_X1 U6825 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7289) );
  OR2_X1 U6826 ( .A1(n5579), .A2(n7289), .ZN(n5408) );
  INV_X1 U6827 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10394) );
  NAND2_X1 U6828 ( .A1(n5403), .A2(n10394), .ZN(n5404) );
  NAND2_X1 U6829 ( .A1(n5429), .A2(n5404), .ZN(n7391) );
  OR2_X1 U6830 ( .A1(n5726), .A2(n7391), .ZN(n5407) );
  INV_X1 U6831 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n5405) );
  OR2_X1 U6832 ( .A1(n7827), .A2(n5405), .ZN(n5406) );
  OR2_X1 U6833 ( .A1(n7449), .A2(n5771), .ZN(n5411) );
  NAND2_X1 U6834 ( .A1(n5410), .A2(n5411), .ZN(n5416) );
  INV_X1 U6835 ( .A(n5410), .ZN(n5413) );
  INV_X1 U6836 ( .A(n5411), .ZN(n5412) );
  NAND2_X1 U6837 ( .A1(n5413), .A2(n5412), .ZN(n5414) );
  NAND2_X1 U6838 ( .A1(n5416), .A2(n5414), .ZN(n7388) );
  INV_X1 U6839 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6775) );
  INV_X1 U6840 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6777) );
  INV_X1 U6841 ( .A(SI_13_), .ZN(n10379) );
  NAND2_X1 U6842 ( .A1(n5420), .A2(n10379), .ZN(n5440) );
  INV_X1 U6843 ( .A(n5420), .ZN(n5421) );
  NAND2_X1 U6844 ( .A1(n5421), .A2(SI_13_), .ZN(n5422) );
  XNOR2_X1 U6845 ( .A(n5439), .B(n5080), .ZN(n6774) );
  NAND2_X1 U6846 ( .A1(n6774), .A2(n5220), .ZN(n5426) );
  INV_X1 U6847 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5423) );
  NAND2_X1 U6848 ( .A1(n5424), .A2(n5423), .ZN(n5500) );
  NAND2_X1 U6849 ( .A1(n5500), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5443) );
  XNOR2_X1 U6850 ( .A(n5443), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7458) );
  AOI22_X1 U6851 ( .A1(n5569), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5568), .B2(
        n7458), .ZN(n5425) );
  XNOR2_X1 U6852 ( .A(n7534), .B(n5137), .ZN(n5435) );
  NAND2_X1 U6853 ( .A1(n5576), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5434) );
  INV_X1 U6854 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5427) );
  OR2_X1 U6855 ( .A1(n5579), .A2(n5427), .ZN(n5433) );
  INV_X1 U6856 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5428) );
  NAND2_X1 U6857 ( .A1(n5429), .A2(n5428), .ZN(n5430) );
  NAND2_X1 U6858 ( .A1(n5451), .A2(n5430), .ZN(n7448) );
  OR2_X1 U6859 ( .A1(n5726), .A2(n7448), .ZN(n5432) );
  INV_X1 U6860 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7419) );
  OR2_X1 U6861 ( .A1(n5199), .A2(n7419), .ZN(n5431) );
  NOR2_X1 U6862 ( .A1(n7554), .A2(n5771), .ZN(n5436) );
  XNOR2_X1 U6863 ( .A(n5435), .B(n5436), .ZN(n7446) );
  INV_X1 U6864 ( .A(n5435), .ZN(n5437) );
  AND2_X1 U6865 ( .A1(n5437), .A2(n5436), .ZN(n5438) );
  MUX2_X1 U6866 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n7832), .Z(n5465) );
  INV_X1 U6867 ( .A(SI_14_), .ZN(n10223) );
  XNOR2_X1 U6868 ( .A(n5468), .B(n5464), .ZN(n6801) );
  NAND2_X1 U6869 ( .A1(n6801), .A2(n5220), .ZN(n5449) );
  NAND2_X1 U6870 ( .A1(n5443), .A2(n5442), .ZN(n5444) );
  NAND2_X1 U6871 ( .A1(n5444), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5446) );
  NAND2_X1 U6872 ( .A1(n5446), .A2(n5445), .ZN(n5473) );
  OR2_X1 U6873 ( .A1(n5446), .A2(n5445), .ZN(n5447) );
  AND2_X1 U6874 ( .A1(n5473), .A2(n5447), .ZN(n8174) );
  AOI22_X1 U6875 ( .A1(n5569), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8174), .B2(
        n5568), .ZN(n5448) );
  XNOR2_X1 U6876 ( .A(n7567), .B(n5137), .ZN(n5458) );
  NAND2_X1 U6877 ( .A1(n5576), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5457) );
  INV_X1 U6878 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10442) );
  NAND2_X1 U6879 ( .A1(n5451), .A2(n10442), .ZN(n5452) );
  NAND2_X1 U6880 ( .A1(n5481), .A2(n5452), .ZN(n7553) );
  OR2_X1 U6881 ( .A1(n7553), .A2(n5726), .ZN(n5456) );
  INV_X1 U6882 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n5453) );
  OR2_X1 U6883 ( .A1(n5579), .A2(n5453), .ZN(n5455) );
  INV_X1 U6884 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7537) );
  OR2_X1 U6885 ( .A1(n5199), .A2(n7537), .ZN(n5454) );
  INV_X1 U6886 ( .A(n7642), .ZN(n8154) );
  NAND2_X1 U6887 ( .A1(n8154), .A2(n7839), .ZN(n5459) );
  NAND2_X1 U6888 ( .A1(n5458), .A2(n5459), .ZN(n5463) );
  INV_X1 U6889 ( .A(n5458), .ZN(n5461) );
  INV_X1 U6890 ( .A(n5459), .ZN(n5460) );
  NAND2_X1 U6891 ( .A1(n5461), .A2(n5460), .ZN(n5462) );
  AND2_X1 U6892 ( .A1(n5463), .A2(n5462), .ZN(n7551) );
  NAND2_X1 U6893 ( .A1(n7550), .A2(n7551), .ZN(n7549) );
  INV_X1 U6894 ( .A(n7638), .ZN(n5489) );
  NAND2_X1 U6895 ( .A1(n5465), .A2(SI_14_), .ZN(n5466) );
  INV_X1 U6896 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6875) );
  INV_X1 U6897 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10454) );
  INV_X1 U6898 ( .A(SI_15_), .ZN(n5469) );
  INV_X1 U6899 ( .A(n5470), .ZN(n5471) );
  NAND2_X1 U6900 ( .A1(n5471), .A2(SI_15_), .ZN(n5472) );
  XNOR2_X1 U6901 ( .A(n5492), .B(n5491), .ZN(n6874) );
  NAND2_X1 U6902 ( .A1(n6874), .A2(n5220), .ZN(n5478) );
  NAND2_X1 U6903 ( .A1(n5473), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5474) );
  XNOR2_X1 U6904 ( .A(n5475), .B(n5474), .ZN(n8187) );
  OAI22_X1 U6905 ( .A1(n8187), .A2(n6556), .B1(n5221), .B2(n6875), .ZN(n5476)
         );
  INV_X1 U6906 ( .A(n5476), .ZN(n5477) );
  XNOR2_X1 U6907 ( .A(n7658), .B(n5137), .ZN(n7637) );
  INV_X1 U6908 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5480) );
  NAND2_X1 U6909 ( .A1(n5481), .A2(n5480), .ZN(n5482) );
  NAND2_X1 U6910 ( .A1(n5505), .A2(n5482), .ZN(n7641) );
  OR2_X1 U6911 ( .A1(n7641), .A2(n5726), .ZN(n5488) );
  INV_X1 U6912 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n5483) );
  OR2_X1 U6913 ( .A1(n5579), .A2(n5483), .ZN(n5485) );
  INV_X1 U6914 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7571) );
  OR2_X1 U6915 ( .A1(n5199), .A2(n7571), .ZN(n5484) );
  AND2_X1 U6916 ( .A1(n5485), .A2(n5484), .ZN(n5487) );
  NAND2_X1 U6917 ( .A1(n5576), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5486) );
  OR2_X1 U6918 ( .A1(n8093), .A2(n5771), .ZN(n5510) );
  INV_X1 U6919 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5493) );
  INV_X1 U6920 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10194) );
  MUX2_X1 U6921 ( .A(n5493), .B(n10194), .S(n7832), .Z(n5494) );
  INV_X1 U6922 ( .A(SI_16_), .ZN(n10455) );
  NAND2_X1 U6923 ( .A1(n5494), .A2(n10455), .ZN(n5521) );
  INV_X1 U6924 ( .A(n5494), .ZN(n5495) );
  NAND2_X1 U6925 ( .A1(n5495), .A2(SI_16_), .ZN(n5496) );
  XNOR2_X1 U6926 ( .A(n5520), .B(n5519), .ZN(n6849) );
  NAND2_X1 U6927 ( .A1(n6849), .A2(n5220), .ZN(n5504) );
  INV_X1 U6928 ( .A(n5498), .ZN(n5499) );
  OAI21_X1 U6929 ( .B1(n5500), .B2(n5499), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5501) );
  MUX2_X1 U6930 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5501), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5502) );
  AND2_X1 U6931 ( .A1(n5524), .A2(n5502), .ZN(n8203) );
  AOI22_X1 U6932 ( .A1(n5569), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5568), .B2(
        n8203), .ZN(n5503) );
  XNOR2_X1 U6933 ( .A(n8578), .B(n5137), .ZN(n5517) );
  INV_X1 U6934 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10436) );
  NAND2_X1 U6935 ( .A1(n5505), .A2(n10436), .ZN(n5506) );
  AND2_X1 U6936 ( .A1(n5529), .A2(n5506), .ZN(n8095) );
  INV_X1 U6937 ( .A(n5726), .ZN(n5826) );
  NAND2_X1 U6938 ( .A1(n8095), .A2(n5826), .ZN(n5509) );
  AOI22_X1 U6939 ( .A1(n5822), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n7823), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n5508) );
  NAND2_X1 U6940 ( .A1(n5576), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5507) );
  NOR2_X1 U6941 ( .A1(n7650), .A2(n5771), .ZN(n5515) );
  XNOR2_X1 U6942 ( .A(n5517), .B(n5515), .ZN(n8087) );
  INV_X1 U6943 ( .A(n7637), .ZN(n5511) );
  INV_X1 U6944 ( .A(n5510), .ZN(n7640) );
  NAND2_X1 U6945 ( .A1(n5511), .A2(n7640), .ZN(n5512) );
  AND2_X1 U6946 ( .A1(n8087), .A2(n5512), .ZN(n5513) );
  INV_X1 U6947 ( .A(n5515), .ZN(n5516) );
  NAND2_X1 U6948 ( .A1(n5517), .A2(n5516), .ZN(n5518) );
  INV_X1 U6949 ( .A(SI_17_), .ZN(n5523) );
  XNOR2_X1 U6950 ( .A(n5541), .B(n5523), .ZN(n5540) );
  XNOR2_X1 U6951 ( .A(n5544), .B(n5540), .ZN(n6886) );
  NAND2_X1 U6952 ( .A1(n6886), .A2(n5220), .ZN(n5527) );
  NAND2_X1 U6953 ( .A1(n5524), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5525) );
  XNOR2_X1 U6954 ( .A(n5525), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8218) );
  AOI22_X1 U6955 ( .A1(n5569), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5568), .B2(
        n8218), .ZN(n5526) );
  XNOR2_X1 U6956 ( .A(n8571), .B(n5137), .ZN(n5534) );
  INV_X1 U6957 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10407) );
  NAND2_X1 U6958 ( .A1(n5529), .A2(n10407), .ZN(n5530) );
  NAND2_X1 U6959 ( .A1(n5549), .A2(n5530), .ZN(n8488) );
  OR2_X1 U6960 ( .A1(n8488), .A2(n5726), .ZN(n5533) );
  AOI22_X1 U6961 ( .A1(n5822), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n7823), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U6962 ( .A1(n5576), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5531) );
  INV_X1 U6963 ( .A(n8130), .ZN(n8466) );
  NAND2_X1 U6964 ( .A1(n8466), .A2(n7839), .ZN(n5535) );
  XNOR2_X1 U6965 ( .A(n5534), .B(n5535), .ZN(n7623) );
  INV_X1 U6966 ( .A(n5534), .ZN(n5537) );
  INV_X1 U6967 ( .A(n5535), .ZN(n5536) );
  NAND2_X1 U6968 ( .A1(n5537), .A2(n5536), .ZN(n5538) );
  INV_X1 U6969 ( .A(n5540), .ZN(n5543) );
  NAND2_X1 U6970 ( .A1(n5541), .A2(SI_17_), .ZN(n5542) );
  MUX2_X1 U6971 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7832), .Z(n5561) );
  XNOR2_X1 U6972 ( .A(n5561), .B(SI_18_), .ZN(n5558) );
  XNOR2_X1 U6973 ( .A(n5560), .B(n5558), .ZN(n7077) );
  NAND2_X1 U6974 ( .A1(n7077), .A2(n5220), .ZN(n5547) );
  NAND2_X1 U6975 ( .A1(n4556), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5545) );
  XNOR2_X1 U6976 ( .A(n5545), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8232) );
  AOI22_X1 U6977 ( .A1(n5569), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5568), .B2(
        n8232), .ZN(n5546) );
  XNOR2_X1 U6978 ( .A(n8568), .B(n5137), .ZN(n5554) );
  INV_X1 U6979 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U6980 ( .A1(n5549), .A2(n5548), .ZN(n5550) );
  AND2_X1 U6981 ( .A1(n5574), .A2(n5550), .ZN(n8127) );
  INV_X1 U6982 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8473) );
  NAND2_X1 U6983 ( .A1(n5822), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U6984 ( .A1(n5576), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5551) );
  OAI211_X1 U6985 ( .C1(n5199), .C2(n8473), .A(n5552), .B(n5551), .ZN(n5553)
         );
  AOI21_X1 U6986 ( .B1(n8127), .B2(n5826), .A(n5553), .ZN(n8152) );
  NOR2_X1 U6987 ( .A1(n8152), .A2(n5771), .ZN(n5555) );
  XNOR2_X1 U6988 ( .A(n5554), .B(n5555), .ZN(n8125) );
  INV_X1 U6989 ( .A(n5554), .ZN(n5556) );
  NAND2_X1 U6990 ( .A1(n5556), .A2(n5555), .ZN(n5557) );
  INV_X1 U6991 ( .A(n5558), .ZN(n5559) );
  NAND2_X1 U6992 ( .A1(n5560), .A2(n5559), .ZN(n5563) );
  NAND2_X1 U6993 ( .A1(n5561), .A2(SI_18_), .ZN(n5562) );
  INV_X1 U6994 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7150) );
  INV_X1 U6995 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10389) );
  INV_X1 U6996 ( .A(SI_19_), .ZN(n5564) );
  NAND2_X1 U6997 ( .A1(n5565), .A2(n5564), .ZN(n5589) );
  INV_X1 U6998 ( .A(n5565), .ZN(n5566) );
  NAND2_X1 U6999 ( .A1(n5566), .A2(SI_19_), .ZN(n5567) );
  NAND2_X1 U7000 ( .A1(n5589), .A2(n5567), .ZN(n5590) );
  XNOR2_X1 U7001 ( .A(n5591), .B(n5590), .ZN(n7148) );
  NAND2_X1 U7002 ( .A1(n7148), .A2(n5220), .ZN(n5571) );
  AOI22_X1 U7003 ( .A1(n5569), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5568), .B2(
        n8356), .ZN(n5570) );
  XNOR2_X1 U7004 ( .A(n8559), .B(n5137), .ZN(n5583) );
  INV_X1 U7005 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U7006 ( .A1(n5574), .A2(n5573), .ZN(n5575) );
  NAND2_X1 U7007 ( .A1(n5597), .A2(n5575), .ZN(n8451) );
  OR2_X1 U7008 ( .A1(n8451), .A2(n5726), .ZN(n5582) );
  INV_X1 U7009 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8235) );
  NAND2_X1 U7010 ( .A1(n7823), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U7011 ( .A1(n5576), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5577) );
  OAI211_X1 U7012 ( .C1(n5579), .C2(n8235), .A(n5578), .B(n5577), .ZN(n5580)
         );
  INV_X1 U7013 ( .A(n5580), .ZN(n5581) );
  INV_X1 U7014 ( .A(n8427), .ZN(n8467) );
  NAND2_X1 U7015 ( .A1(n8467), .A2(n7839), .ZN(n5584) );
  NAND2_X1 U7016 ( .A1(n5583), .A2(n5584), .ZN(n5588) );
  INV_X1 U7017 ( .A(n5583), .ZN(n5586) );
  INV_X1 U7018 ( .A(n5584), .ZN(n5585) );
  NAND2_X1 U7019 ( .A1(n5586), .A2(n5585), .ZN(n5587) );
  NAND2_X1 U7020 ( .A1(n5588), .A2(n5587), .ZN(n8063) );
  INV_X1 U7021 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7250) );
  INV_X1 U7022 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10451) );
  MUX2_X1 U7023 ( .A(n7250), .B(n10451), .S(n7832), .Z(n5592) );
  INV_X1 U7024 ( .A(SI_20_), .ZN(n10404) );
  NAND2_X1 U7025 ( .A1(n5592), .A2(n10404), .ZN(n5609) );
  INV_X1 U7026 ( .A(n5592), .ZN(n5593) );
  NAND2_X1 U7027 ( .A1(n5593), .A2(SI_20_), .ZN(n5594) );
  XNOR2_X1 U7028 ( .A(n5608), .B(n5607), .ZN(n7233) );
  NAND2_X1 U7029 ( .A1(n7233), .A2(n5220), .ZN(n5596) );
  OR2_X1 U7030 ( .A1(n5221), .A2(n7250), .ZN(n5595) );
  XNOR2_X1 U7031 ( .A(n8554), .B(n5772), .ZN(n5603) );
  INV_X1 U7032 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10318) );
  NAND2_X1 U7033 ( .A1(n5597), .A2(n10318), .ZN(n5598) );
  AND2_X1 U7034 ( .A1(n5613), .A2(n5598), .ZN(n8434) );
  INV_X1 U7035 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n5601) );
  NAND2_X1 U7036 ( .A1(n7823), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U7037 ( .A1(n5822), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5599) );
  OAI211_X1 U7038 ( .C1(n5601), .C2(n7827), .A(n5600), .B(n5599), .ZN(n5602)
         );
  AOI21_X1 U7039 ( .B1(n8434), .B2(n5826), .A(n5602), .ZN(n8151) );
  NOR2_X1 U7040 ( .A1(n8151), .A2(n5771), .ZN(n5604) );
  XNOR2_X1 U7041 ( .A(n5603), .B(n5604), .ZN(n8107) );
  INV_X1 U7042 ( .A(n5603), .ZN(n5606) );
  INV_X1 U7043 ( .A(n5604), .ZN(n5605) );
  INV_X1 U7044 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7331) );
  INV_X1 U7045 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7303) );
  XNOR2_X1 U7046 ( .A(n5628), .B(SI_21_), .ZN(n5627) );
  XNOR2_X1 U7047 ( .A(n5626), .B(n5627), .ZN(n7302) );
  NAND2_X1 U7048 ( .A1(n7302), .A2(n5220), .ZN(n5611) );
  OR2_X1 U7049 ( .A1(n5221), .A2(n7331), .ZN(n5610) );
  XNOR2_X1 U7050 ( .A(n8549), .B(n5137), .ZN(n5621) );
  INV_X1 U7051 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8073) );
  NAND2_X1 U7052 ( .A1(n5613), .A2(n8073), .ZN(n5614) );
  NAND2_X1 U7053 ( .A1(n5638), .A2(n5614), .ZN(n8415) );
  OR2_X1 U7054 ( .A1(n8415), .A2(n5726), .ZN(n5620) );
  INV_X1 U7055 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U7056 ( .A1(n5822), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5616) );
  NAND2_X1 U7057 ( .A1(n7823), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5615) );
  OAI211_X1 U7058 ( .C1(n7827), .C2(n5617), .A(n5616), .B(n5615), .ZN(n5618)
         );
  INV_X1 U7059 ( .A(n5618), .ZN(n5619) );
  NOR2_X1 U7060 ( .A1(n8429), .A2(n5771), .ZN(n5622) );
  XNOR2_X1 U7061 ( .A(n5621), .B(n5622), .ZN(n8071) );
  NAND2_X1 U7062 ( .A1(n8072), .A2(n8071), .ZN(n5625) );
  INV_X1 U7063 ( .A(n5621), .ZN(n5623) );
  NAND2_X1 U7064 ( .A1(n5623), .A2(n5622), .ZN(n5624) );
  NAND2_X1 U7065 ( .A1(n5625), .A2(n5624), .ZN(n5648) );
  INV_X1 U7066 ( .A(n5628), .ZN(n5629) );
  NAND2_X1 U7067 ( .A1(n5629), .A2(SI_21_), .ZN(n5630) );
  INV_X1 U7068 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7802) );
  INV_X1 U7069 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10434) );
  MUX2_X1 U7070 ( .A(n7802), .B(n10434), .S(n7832), .Z(n5632) );
  INV_X1 U7071 ( .A(SI_22_), .ZN(n10423) );
  NAND2_X1 U7072 ( .A1(n5632), .A2(n10423), .ZN(n5650) );
  INV_X1 U7073 ( .A(n5632), .ZN(n5633) );
  NAND2_X1 U7074 ( .A1(n5633), .A2(SI_22_), .ZN(n5634) );
  NAND2_X1 U7075 ( .A1(n5650), .A2(n5634), .ZN(n5651) );
  XNOR2_X1 U7076 ( .A(n5652), .B(n5651), .ZN(n7433) );
  NAND2_X1 U7077 ( .A1(n7433), .A2(n5220), .ZN(n5636) );
  OR2_X1 U7078 ( .A1(n5221), .A2(n7802), .ZN(n5635) );
  XNOR2_X1 U7079 ( .A(n8546), .B(n5137), .ZN(n5646) );
  XNOR2_X1 U7080 ( .A(n5648), .B(n5646), .ZN(n8116) );
  INV_X1 U7081 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10424) );
  NAND2_X1 U7082 ( .A1(n5638), .A2(n10424), .ZN(n5639) );
  NAND2_X1 U7083 ( .A1(n5658), .A2(n5639), .ZN(n8402) );
  OR2_X1 U7084 ( .A1(n8402), .A2(n5726), .ZN(n5645) );
  INV_X1 U7085 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n5642) );
  NAND2_X1 U7086 ( .A1(n5822), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U7087 ( .A1(n7823), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5640) );
  OAI211_X1 U7088 ( .C1(n7827), .C2(n5642), .A(n5641), .B(n5640), .ZN(n5643)
         );
  INV_X1 U7089 ( .A(n5643), .ZN(n5644) );
  OR2_X1 U7090 ( .A1(n8150), .A2(n5771), .ZN(n8115) );
  NAND2_X1 U7091 ( .A1(n8116), .A2(n8115), .ZN(n8114) );
  INV_X1 U7092 ( .A(n5646), .ZN(n5647) );
  OR2_X1 U7093 ( .A1(n5648), .A2(n5647), .ZN(n5649) );
  INV_X1 U7094 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7485) );
  INV_X1 U7095 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n10465) );
  INV_X1 U7096 ( .A(SI_23_), .ZN(n10390) );
  NAND2_X1 U7097 ( .A1(n5653), .A2(n10390), .ZN(n5673) );
  INV_X1 U7098 ( .A(n5653), .ZN(n5654) );
  NAND2_X1 U7099 ( .A1(n5654), .A2(SI_23_), .ZN(n5655) );
  NAND2_X1 U7100 ( .A1(n7486), .A2(n5220), .ZN(n5657) );
  OR2_X1 U7101 ( .A1(n5221), .A2(n7485), .ZN(n5656) );
  XNOR2_X1 U7102 ( .A(n8538), .B(n5772), .ZN(n5666) );
  INV_X1 U7103 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8047) );
  NAND2_X1 U7104 ( .A1(n5658), .A2(n8047), .ZN(n5659) );
  NAND2_X1 U7105 ( .A1(n5678), .A2(n5659), .ZN(n8385) );
  OR2_X1 U7106 ( .A1(n8385), .A2(n5726), .ZN(n5665) );
  INV_X1 U7107 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n5662) );
  NAND2_X1 U7108 ( .A1(n5150), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U7109 ( .A1(n7823), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5660) );
  OAI211_X1 U7110 ( .C1(n5662), .C2(n7827), .A(n5661), .B(n5660), .ZN(n5663)
         );
  INV_X1 U7111 ( .A(n5663), .ZN(n5664) );
  NAND2_X1 U7112 ( .A1(n5665), .A2(n5664), .ZN(n8273) );
  AND2_X1 U7113 ( .A1(n8273), .A2(n7839), .ZN(n8045) );
  NAND2_X1 U7114 ( .A1(n8046), .A2(n8045), .ZN(n5670) );
  INV_X1 U7115 ( .A(n5666), .ZN(n5667) );
  OR2_X1 U7116 ( .A1(n5668), .A2(n5667), .ZN(n5669) );
  MUX2_X1 U7117 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n7832), .Z(n5689) );
  INV_X1 U7118 ( .A(SI_24_), .ZN(n5675) );
  XNOR2_X1 U7119 ( .A(n5689), .B(n5675), .ZN(n5688) );
  XNOR2_X1 U7120 ( .A(n5692), .B(n5688), .ZN(n7543) );
  NAND2_X1 U7121 ( .A1(n7543), .A2(n5220), .ZN(n5677) );
  INV_X1 U7122 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7546) );
  OR2_X1 U7123 ( .A1(n5221), .A2(n7546), .ZN(n5676) );
  XNOR2_X1 U7124 ( .A(n8533), .B(n5137), .ZN(n5684) );
  INV_X1 U7125 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10253) );
  NAND2_X1 U7126 ( .A1(n5678), .A2(n10253), .ZN(n5679) );
  AND2_X1 U7127 ( .A1(n5701), .A2(n5679), .ZN(n8364) );
  INV_X1 U7128 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n5682) );
  NAND2_X1 U7129 ( .A1(n5822), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5681) );
  NAND2_X1 U7130 ( .A1(n7823), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5680) );
  OAI211_X1 U7131 ( .C1(n7827), .C2(n5682), .A(n5681), .B(n5680), .ZN(n5683)
         );
  AOI21_X1 U7132 ( .B1(n8364), .B2(n5826), .A(n5683), .ZN(n8149) );
  NOR2_X1 U7133 ( .A1(n8149), .A2(n5771), .ZN(n8099) );
  INV_X1 U7134 ( .A(n5684), .ZN(n5685) );
  NAND2_X1 U7135 ( .A1(n5686), .A2(n5685), .ZN(n5687) );
  INV_X1 U7136 ( .A(n5688), .ZN(n5691) );
  NAND2_X1 U7137 ( .A1(n5689), .A2(SI_24_), .ZN(n5690) );
  INV_X1 U7138 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7619) );
  INV_X1 U7139 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10437) );
  INV_X1 U7140 ( .A(SI_25_), .ZN(n5693) );
  NAND2_X1 U7141 ( .A1(n5694), .A2(n5693), .ZN(n5713) );
  INV_X1 U7142 ( .A(n5694), .ZN(n5695) );
  NAND2_X1 U7143 ( .A1(n5695), .A2(SI_25_), .ZN(n5696) );
  NAND2_X1 U7144 ( .A1(n5713), .A2(n5696), .ZN(n5714) );
  NAND2_X1 U7145 ( .A1(n7617), .A2(n5220), .ZN(n5698) );
  OR2_X1 U7146 ( .A1(n5221), .A2(n7619), .ZN(n5697) );
  XNOR2_X1 U7147 ( .A(n8529), .B(n5772), .ZN(n5711) );
  INV_X1 U7148 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U7149 ( .A1(n5701), .A2(n5700), .ZN(n5702) );
  NAND2_X1 U7150 ( .A1(n5724), .A2(n5702), .ZN(n8081) );
  OR2_X1 U7151 ( .A1(n8081), .A2(n5726), .ZN(n5708) );
  INV_X1 U7152 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n5705) );
  NAND2_X1 U7153 ( .A1(n5822), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5704) );
  NAND2_X1 U7154 ( .A1(n7823), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5703) );
  OAI211_X1 U7155 ( .C1(n5705), .C2(n7827), .A(n5704), .B(n5703), .ZN(n5706)
         );
  INV_X1 U7156 ( .A(n5706), .ZN(n5707) );
  NAND2_X1 U7157 ( .A1(n8277), .A2(n7839), .ZN(n5709) );
  XNOR2_X1 U7158 ( .A(n5711), .B(n5709), .ZN(n8078) );
  INV_X1 U7159 ( .A(n5709), .ZN(n5710) );
  NAND2_X1 U7160 ( .A1(n5711), .A2(n5710), .ZN(n5712) );
  INV_X1 U7161 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7632) );
  INV_X1 U7162 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10449) );
  MUX2_X1 U7163 ( .A(n7632), .B(n10449), .S(n7832), .Z(n5717) );
  INV_X1 U7164 ( .A(SI_26_), .ZN(n5716) );
  NAND2_X1 U7165 ( .A1(n5717), .A2(n5716), .ZN(n5740) );
  INV_X1 U7166 ( .A(n5717), .ZN(n5718) );
  NAND2_X1 U7167 ( .A1(n5718), .A2(SI_26_), .ZN(n5719) );
  AND2_X1 U7168 ( .A1(n5740), .A2(n5719), .ZN(n5738) );
  NAND2_X1 U7169 ( .A1(n7631), .A2(n5220), .ZN(n5721) );
  OR2_X1 U7170 ( .A1(n5221), .A2(n7632), .ZN(n5720) );
  XNOR2_X1 U7171 ( .A(n8523), .B(n5772), .ZN(n5735) );
  INV_X1 U7172 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n5723) );
  NAND2_X1 U7173 ( .A1(n5724), .A2(n5723), .ZN(n5725) );
  NAND2_X1 U7174 ( .A1(n5763), .A2(n5725), .ZN(n8342) );
  OR2_X1 U7175 ( .A1(n8342), .A2(n5726), .ZN(n5732) );
  INV_X1 U7176 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n5729) );
  NAND2_X1 U7177 ( .A1(n5822), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5728) );
  NAND2_X1 U7178 ( .A1(n7823), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5727) );
  OAI211_X1 U7179 ( .C1(n5729), .C2(n7827), .A(n5728), .B(n5727), .ZN(n5730)
         );
  INV_X1 U7180 ( .A(n5730), .ZN(n5731) );
  NAND2_X1 U7181 ( .A1(n5732), .A2(n5731), .ZN(n8278) );
  NAND2_X1 U7182 ( .A1(n8278), .A2(n7839), .ZN(n5733) );
  XNOR2_X1 U7183 ( .A(n5735), .B(n5733), .ZN(n8137) );
  NAND2_X1 U7184 ( .A1(n8136), .A2(n8137), .ZN(n5737) );
  INV_X1 U7185 ( .A(n5733), .ZN(n5734) );
  NAND2_X1 U7186 ( .A1(n5735), .A2(n5734), .ZN(n5736) );
  INV_X1 U7187 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7728) );
  INV_X1 U7188 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10272) );
  INV_X1 U7189 ( .A(SI_27_), .ZN(n10428) );
  NAND2_X1 U7190 ( .A1(n5742), .A2(n10428), .ZN(n5759) );
  INV_X1 U7191 ( .A(n5742), .ZN(n5743) );
  NAND2_X1 U7192 ( .A1(n5743), .A2(SI_27_), .ZN(n5744) );
  AND2_X1 U7193 ( .A1(n5759), .A2(n5744), .ZN(n5757) );
  NAND2_X1 U7194 ( .A1(n7726), .A2(n5220), .ZN(n5746) );
  OR2_X1 U7195 ( .A1(n5221), .A2(n7728), .ZN(n5745) );
  XNOR2_X1 U7196 ( .A(n8281), .B(n5772), .ZN(n5755) );
  XNOR2_X1 U7197 ( .A(n5763), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8322) );
  NAND2_X1 U7198 ( .A1(n8322), .A2(n5826), .ZN(n5752) );
  INV_X1 U7199 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n5749) );
  NAND2_X1 U7200 ( .A1(n5822), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5748) );
  NAND2_X1 U7201 ( .A1(n7823), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5747) );
  OAI211_X1 U7202 ( .C1(n5749), .C2(n7827), .A(n5748), .B(n5747), .ZN(n5750)
         );
  INV_X1 U7203 ( .A(n5750), .ZN(n5751) );
  NAND2_X1 U7204 ( .A1(n5752), .A2(n5751), .ZN(n8280) );
  NAND2_X1 U7205 ( .A1(n8280), .A2(n7839), .ZN(n5753) );
  XNOR2_X1 U7206 ( .A(n5755), .B(n5753), .ZN(n8038) );
  INV_X1 U7207 ( .A(n5753), .ZN(n5754) );
  AND2_X1 U7208 ( .A1(n5755), .A2(n5754), .ZN(n5756) );
  AOI21_X1 U7209 ( .B1(n8037), .B2(n8038), .A(n5756), .ZN(n5816) );
  MUX2_X1 U7210 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7832), .Z(n7708) );
  INV_X1 U7211 ( .A(SI_28_), .ZN(n10392) );
  XNOR2_X1 U7212 ( .A(n7708), .B(n10392), .ZN(n7706) );
  NAND2_X1 U7213 ( .A1(n7770), .A2(n5220), .ZN(n5761) );
  INV_X1 U7214 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7705) );
  OR2_X1 U7215 ( .A1(n5221), .A2(n7705), .ZN(n5760) );
  NOR2_X1 U7216 ( .A1(n8309), .A2(n10002), .ZN(n5776) );
  INV_X1 U7217 ( .A(n5776), .ZN(n5774) );
  INV_X1 U7218 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8039) );
  INV_X1 U7219 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5834) );
  OAI21_X1 U7220 ( .B1(n5763), .B2(n8039), .A(n5834), .ZN(n5764) );
  NAND2_X1 U7221 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n5762) );
  NAND2_X1 U7222 ( .A1(n8306), .A2(n5826), .ZN(n5770) );
  INV_X1 U7223 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5767) );
  NAND2_X1 U7224 ( .A1(n7823), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5766) );
  NAND2_X1 U7225 ( .A1(n5822), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5765) );
  OAI211_X1 U7226 ( .C1(n5767), .C2(n7827), .A(n5766), .B(n5765), .ZN(n5768)
         );
  INV_X1 U7227 ( .A(n5768), .ZN(n5769) );
  NOR2_X1 U7228 ( .A1(n8257), .A2(n5771), .ZN(n5773) );
  XNOR2_X1 U7229 ( .A(n5773), .B(n5772), .ZN(n5775) );
  MUX2_X1 U7230 ( .A(n5774), .B(n8511), .S(n5775), .Z(n5815) );
  MUX2_X1 U7231 ( .A(n8309), .B(n5776), .S(n5775), .Z(n5777) );
  NAND2_X1 U7232 ( .A1(n5816), .A2(n5777), .ZN(n5814) );
  NAND2_X1 U7233 ( .A1(n5778), .A2(n5782), .ZN(n5779) );
  NAND2_X1 U7234 ( .A1(n5779), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5808) );
  NAND2_X1 U7235 ( .A1(n5808), .A2(n5807), .ZN(n5810) );
  NAND2_X1 U7236 ( .A1(n5810), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5780) );
  XNOR2_X1 U7237 ( .A(n5780), .B(P2_IR_REG_24__SCAN_IN), .ZN(n7545) );
  INV_X1 U7238 ( .A(P2_B_REG_SCAN_IN), .ZN(n10262) );
  XNOR2_X1 U7239 ( .A(n7545), .B(n10262), .ZN(n5786) );
  NAND3_X1 U7240 ( .A1(n5782), .A2(n5807), .A3(n5781), .ZN(n5783) );
  OAI21_X1 U7241 ( .B1(n4497), .B2(n5783), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5784) );
  MUX2_X1 U7242 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5784), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5785) );
  NAND2_X1 U7243 ( .A1(n5785), .A2(n5787), .ZN(n7618) );
  NAND2_X1 U7244 ( .A1(n5786), .A2(n7618), .ZN(n5791) );
  NAND2_X1 U7245 ( .A1(n5787), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5788) );
  MUX2_X1 U7246 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5788), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5790) );
  NAND2_X1 U7247 ( .A1(n5790), .A2(n5789), .ZN(n7633) );
  INV_X1 U7248 ( .A(n7633), .ZN(n5792) );
  INV_X1 U7249 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9957) );
  NAND2_X1 U7250 ( .A1(n9955), .A2(n9957), .ZN(n5794) );
  NOR2_X1 U7251 ( .A1(n7545), .A2(n5792), .ZN(n9958) );
  INV_X1 U7252 ( .A(n9958), .ZN(n5793) );
  NAND2_X1 U7253 ( .A1(n5794), .A2(n5793), .ZN(n6921) );
  INV_X1 U7254 ( .A(n6921), .ZN(n6692) );
  INV_X1 U7255 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9960) );
  AND2_X1 U7256 ( .A1(n7618), .A2(n7633), .ZN(n9961) );
  AOI21_X1 U7257 ( .B1(n9955), .B2(n9960), .A(n9961), .ZN(n6922) );
  NOR2_X1 U7258 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n5798) );
  NOR4_X1 U7259 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n5797) );
  NOR4_X1 U7260 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5796) );
  NOR4_X1 U7261 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5795) );
  AND4_X1 U7262 ( .A1(n5798), .A2(n5797), .A3(n5796), .A4(n5795), .ZN(n5804)
         );
  NOR4_X1 U7263 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5802) );
  NOR4_X1 U7264 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5801) );
  NOR4_X1 U7265 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5800) );
  NOR4_X1 U7266 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5799) );
  AND4_X1 U7267 ( .A1(n5802), .A2(n5801), .A3(n5800), .A4(n5799), .ZN(n5803)
         );
  NAND2_X1 U7268 ( .A1(n5804), .A2(n5803), .ZN(n5805) );
  NAND2_X1 U7269 ( .A1(n9955), .A2(n5805), .ZN(n6690) );
  NAND3_X1 U7270 ( .A1(n6692), .A2(n6922), .A3(n6690), .ZN(n5829) );
  NOR2_X1 U7271 ( .A1(n7618), .A2(n7633), .ZN(n5806) );
  NAND2_X1 U7272 ( .A1(n7545), .A2(n5806), .ZN(n6554) );
  OR2_X1 U7273 ( .A1(n5808), .A2(n5807), .ZN(n5809) );
  NAND2_X1 U7274 ( .A1(n5810), .A2(n5809), .ZN(n5830) );
  NAND2_X1 U7275 ( .A1(n6554), .A2(n9962), .ZN(n9956) );
  OR2_X1 U7276 ( .A1(n5829), .A2(n9956), .ZN(n5817) );
  INV_X1 U7277 ( .A(n7249), .ZN(n8022) );
  OR2_X1 U7278 ( .A1(n9956), .A2(n8022), .ZN(n5811) );
  NAND2_X1 U7279 ( .A1(n5817), .A2(n5811), .ZN(n5812) );
  NAND2_X1 U7280 ( .A1(n5812), .A2(n10002), .ZN(n8123) );
  NAND2_X1 U7281 ( .A1(n8030), .A2(n8023), .ZN(n6514) );
  INV_X1 U7282 ( .A(n6514), .ZN(n6552) );
  OAI21_X1 U7283 ( .B1(n8309), .B2(n8123), .A(n8145), .ZN(n5813) );
  OAI211_X1 U7284 ( .C1(n5816), .C2(n5815), .A(n5814), .B(n5813), .ZN(n5840)
         );
  INV_X1 U7285 ( .A(n8280), .ZN(n8297) );
  OR2_X1 U7286 ( .A1(n5817), .A2(n8029), .ZN(n8141) );
  INV_X1 U7287 ( .A(n5818), .ZN(n5820) );
  NOR2_X1 U7288 ( .A1(n8141), .A2(n8428), .ZN(n7717) );
  INV_X1 U7289 ( .A(n5821), .ZN(n8289) );
  INV_X1 U7290 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8586) );
  NAND2_X1 U7291 ( .A1(n5822), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5824) );
  NAND2_X1 U7292 ( .A1(n7823), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5823) );
  OAI211_X1 U7293 ( .C1(n7827), .C2(n8586), .A(n5824), .B(n5823), .ZN(n5825)
         );
  AOI21_X1 U7294 ( .B1(n8289), .B2(n5826), .A(n5825), .ZN(n8296) );
  INV_X1 U7295 ( .A(n8296), .ZN(n8148) );
  INV_X1 U7296 ( .A(n8306), .ZN(n5835) );
  AND2_X1 U7297 ( .A1(n7249), .A2(n8356), .ZN(n5828) );
  AND2_X1 U7298 ( .A1(n10020), .A2(n7828), .ZN(n6691) );
  INV_X1 U7299 ( .A(n6691), .ZN(n6925) );
  NAND2_X1 U7300 ( .A1(n5829), .A2(n6925), .ZN(n5833) );
  NOR2_X1 U7301 ( .A1(n6514), .A2(n4939), .ZN(n6688) );
  INV_X1 U7302 ( .A(n5830), .ZN(n6515) );
  NOR2_X1 U7303 ( .A1(n6688), .A2(n6515), .ZN(n5831) );
  AND2_X1 U7304 ( .A1(n6554), .A2(n5831), .ZN(n5832) );
  NAND2_X1 U7305 ( .A1(n5833), .A2(n5832), .ZN(n6778) );
  NAND2_X1 U7306 ( .A1(n6778), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8128) );
  OAI22_X1 U7307 ( .A1(n5835), .A2(n8128), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5834), .ZN(n5836) );
  AOI21_X1 U7308 ( .B1(n7717), .B2(n8148), .A(n5836), .ZN(n5837) );
  INV_X1 U7309 ( .A(n5837), .ZN(n5838) );
  NOR2_X1 U7310 ( .A1(n5819), .A2(n5838), .ZN(n5839) );
  NAND2_X1 U7311 ( .A1(n5840), .A2(n5839), .ZN(P2_U3222) );
  NOR2_X1 U7312 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5844) );
  NAND2_X1 U7313 ( .A1(n5847), .A2(n5846), .ZN(n5904) );
  NOR2_X1 U7314 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5850) );
  NAND2_X1 U7315 ( .A1(n5907), .A2(n5850), .ZN(n5853) );
  NAND4_X1 U7316 ( .A1(n5852), .A2(n6259), .A3(n5851), .A4(n6157), .ZN(n5906)
         );
  NAND2_X1 U7317 ( .A1(n5902), .A2(n5899), .ZN(n5854) );
  NAND2_X1 U7318 ( .A1(n5876), .A2(n5882), .ZN(n5856) );
  INV_X1 U7319 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5857) );
  INV_X1 U7320 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5893) );
  INV_X1 U7321 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5858) );
  XNOR2_X2 U7322 ( .A(n5862), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5864) );
  INV_X1 U7323 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5895) );
  NAND2_X2 U7324 ( .A1(n5870), .A2(n5864), .ZN(n5929) );
  INV_X1 U7325 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5863) );
  NAND2_X1 U7326 ( .A1(n5865), .A2(n5869), .ZN(n5930) );
  INV_X1 U7327 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5866) );
  AND2_X1 U7328 ( .A1(n5868), .A2(n5867), .ZN(n5873) );
  INV_X1 U7329 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5871) );
  OR2_X1 U7330 ( .A1(n5991), .A2(n5871), .ZN(n5872) );
  NAND2_X1 U7331 ( .A1(n5883), .A2(n5882), .ZN(n5875) );
  NAND2_X1 U7332 ( .A1(n5875), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5877) );
  INV_X1 U7333 ( .A(n5878), .ZN(n5879) );
  NAND2_X1 U7334 ( .A1(n5879), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5881) );
  XNOR2_X1 U7335 ( .A(n5881), .B(n5880), .ZN(n7544) );
  XNOR2_X1 U7336 ( .A(n5883), .B(n5882), .ZN(n7620) );
  NAND2_X1 U7337 ( .A1(n5886), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U7338 ( .A1(n5884), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5885) );
  MUX2_X1 U7339 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5885), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n5887) );
  NAND2_X1 U7340 ( .A1(n5887), .A2(n5886), .ZN(n7234) );
  INV_X1 U7341 ( .A(n7135), .ZN(n6449) );
  AND2_X2 U7342 ( .A1(n6443), .A2(n6449), .ZN(n6067) );
  NAND2_X1 U7343 ( .A1(n7123), .A2(n6067), .ZN(n5898) );
  INV_X1 U7344 ( .A(SI_0_), .ZN(n10439) );
  INV_X1 U7345 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5888) );
  OAI21_X1 U7346 ( .B1(n4876), .B2(n10439), .A(n5888), .ZN(n5890) );
  AND2_X1 U7347 ( .A1(n5890), .A2(n5889), .ZN(n9505) );
  MUX2_X1 U7348 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9505), .S(n9617), .Z(n9799) );
  NOR2_X1 U7349 ( .A1(n6443), .A2(n5895), .ZN(n5896) );
  AOI21_X1 U7350 ( .B1(n9799), .B2(n7773), .A(n5896), .ZN(n5897) );
  NAND2_X1 U7351 ( .A1(n5898), .A2(n5897), .ZN(n6581) );
  NAND2_X1 U7352 ( .A1(n5900), .A2(n5899), .ZN(n5901) );
  NAND2_X1 U7353 ( .A1(n5901), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5903) );
  XNOR2_X1 U7354 ( .A(n5903), .B(n5902), .ZN(n7434) );
  INV_X1 U7355 ( .A(n7434), .ZN(n9024) );
  INV_X1 U7356 ( .A(n5906), .ZN(n5908) );
  INV_X1 U7357 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6139) );
  NAND3_X1 U7358 ( .A1(n5908), .A2(n5907), .A3(n6139), .ZN(n5909) );
  OAI21_X1 U7359 ( .B1(n5905), .B2(n5909), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5910) );
  XNOR2_X1 U7360 ( .A(n5910), .B(P1_IR_REG_19__SCAN_IN), .ZN(n8871) );
  NAND2_X1 U7361 ( .A1(n9024), .A2(n9761), .ZN(n5911) );
  NAND2_X2 U7362 ( .A1(n5911), .A2(n7135), .ZN(n7304) );
  AND2_X1 U7363 ( .A1(n7234), .A2(n9761), .ZN(n6442) );
  NAND2_X1 U7364 ( .A1(n7434), .A2(n6442), .ZN(n5912) );
  INV_X1 U7365 ( .A(n6443), .ZN(n6471) );
  AOI22_X1 U7366 ( .A1(n9799), .A2(n6067), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n6471), .ZN(n5913) );
  NAND2_X1 U7367 ( .A1(n5081), .A2(n6580), .ZN(n5928) );
  INV_X1 U7368 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6647) );
  OR2_X1 U7369 ( .A1(n5991), .A2(n6647), .ZN(n5919) );
  INV_X1 U7370 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5914) );
  OR2_X1 U7371 ( .A1(n5930), .A2(n5914), .ZN(n5918) );
  NAND2_X1 U7372 ( .A1(n5915), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5917) );
  INV_X1 U7373 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7144) );
  INV_X1 U7374 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6499) );
  OR2_X1 U7375 ( .A1(n6018), .A2(n6498), .ZN(n5923) );
  INV_X1 U7376 ( .A(n5920), .ZN(n5921) );
  OR2_X1 U7377 ( .A1(n9617), .A2(n6680), .ZN(n5922) );
  NAND2_X1 U7378 ( .A1(n5925), .A2(n5924), .ZN(n5926) );
  XNOR2_X1 U7379 ( .A(n5926), .B(n7776), .ZN(n5927) );
  AOI22_X1 U7380 ( .A1(n9794), .A2(n6394), .B1(n8888), .B2(n6067), .ZN(n6769)
         );
  NAND2_X1 U7381 ( .A1(n5928), .A2(n5927), .ZN(n6768) );
  INV_X1 U7382 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9892) );
  NAND2_X1 U7383 ( .A1(n5993), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5931) );
  AND2_X1 U7384 ( .A1(n5932), .A2(n5931), .ZN(n5934) );
  INV_X1 U7385 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7168) );
  OR2_X1 U7386 ( .A1(n5991), .A2(n7168), .ZN(n5933) );
  NAND3_X2 U7387 ( .A1(n5935), .A2(n5934), .A3(n5933), .ZN(n7151) );
  NAND2_X1 U7388 ( .A1(n7151), .A2(n6067), .ZN(n5944) );
  OR2_X1 U7389 ( .A1(n6018), .A2(n6493), .ZN(n5942) );
  INV_X1 U7390 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6494) );
  OR2_X1 U7391 ( .A1(n8855), .A2(n6494), .ZN(n5941) );
  NOR2_X1 U7392 ( .A1(n5920), .A2(n5860), .ZN(n5936) );
  MUX2_X1 U7393 ( .A(n5860), .B(n5936), .S(P1_IR_REG_2__SCAN_IN), .Z(n5937) );
  INV_X1 U7394 ( .A(n5937), .ZN(n5939) );
  AND2_X1 U7395 ( .A1(n5939), .A2(n5938), .ZN(n6646) );
  INV_X1 U7396 ( .A(n6646), .ZN(n9630) );
  OR2_X1 U7397 ( .A1(n9617), .A2(n9630), .ZN(n5940) );
  OR2_X1 U7398 ( .A1(n9819), .A2(n6345), .ZN(n5943) );
  NAND2_X1 U7399 ( .A1(n5944), .A2(n5943), .ZN(n5945) );
  XNOR2_X1 U7400 ( .A(n5945), .B(n7776), .ZN(n5946) );
  AOI22_X1 U7401 ( .A1(n7151), .A2(n6394), .B1(n8698), .B2(n6067), .ZN(n5947)
         );
  NAND2_X1 U7402 ( .A1(n5946), .A2(n5947), .ZN(n5951) );
  INV_X1 U7403 ( .A(n5946), .ZN(n5949) );
  INV_X1 U7404 ( .A(n5947), .ZN(n5948) );
  NAND2_X1 U7405 ( .A1(n8695), .A2(n8696), .ZN(n8694) );
  OR2_X1 U7406 ( .A1(n5929), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5960) );
  INV_X1 U7407 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5953) );
  NOR2_X1 U7408 ( .A1(n4479), .A2(n5953), .ZN(n5958) );
  INV_X1 U7409 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U7410 ( .A1(n5993), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5955) );
  NAND2_X1 U7411 ( .A1(n5956), .A2(n5955), .ZN(n5957) );
  NOR2_X1 U7412 ( .A1(n5958), .A2(n5957), .ZN(n5959) );
  NAND2_X2 U7413 ( .A1(n5960), .A2(n5959), .ZN(n9773) );
  NAND2_X1 U7414 ( .A1(n9773), .A2(n6067), .ZN(n5966) );
  OR2_X1 U7415 ( .A1(n6018), .A2(n6496), .ZN(n5964) );
  INV_X1 U7416 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6497) );
  OR2_X1 U7417 ( .A1(n8855), .A2(n6497), .ZN(n5963) );
  NAND2_X1 U7418 ( .A1(n5938), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5961) );
  XNOR2_X1 U7419 ( .A(n5961), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6718) );
  INV_X1 U7420 ( .A(n6718), .ZN(n6495) );
  OR2_X1 U7421 ( .A1(n9617), .A2(n6495), .ZN(n5962) );
  OR2_X1 U7422 ( .A1(n9825), .A2(n6345), .ZN(n5965) );
  NAND2_X1 U7423 ( .A1(n5966), .A2(n5965), .ZN(n5967) );
  XNOR2_X1 U7424 ( .A(n5967), .B(n7304), .ZN(n5982) );
  AOI22_X1 U7425 ( .A1(n9773), .A2(n6394), .B1(n7251), .B2(n6067), .ZN(n5983)
         );
  XNOR2_X1 U7426 ( .A(n5982), .B(n5983), .ZN(n6852) );
  NAND2_X1 U7427 ( .A1(n5993), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5973) );
  INV_X1 U7428 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5968) );
  OR2_X1 U7429 ( .A1(n5991), .A2(n5968), .ZN(n5972) );
  XNOR2_X1 U7430 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n9777) );
  OR2_X1 U7431 ( .A1(n5929), .A2(n9777), .ZN(n5971) );
  INV_X1 U7432 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5969) );
  OR2_X1 U7433 ( .A1(n4479), .A2(n5969), .ZN(n5970) );
  NAND4_X2 U7434 ( .A1(n5973), .A2(n5972), .A3(n5971), .A4(n5970), .ZN(n9035)
         );
  NAND2_X1 U7435 ( .A1(n9035), .A2(n6067), .ZN(n5980) );
  INV_X1 U7436 ( .A(n5974), .ZN(n6501) );
  OR2_X1 U7437 ( .A1(n6018), .A2(n6501), .ZN(n5978) );
  INV_X1 U7438 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6502) );
  OR2_X1 U7439 ( .A1(n8855), .A2(n6502), .ZN(n5977) );
  NAND2_X1 U7440 ( .A1(n6002), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5975) );
  XNOR2_X1 U7441 ( .A(n5975), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9645) );
  INV_X1 U7442 ( .A(n9645), .ZN(n6710) );
  OR2_X1 U7443 ( .A1(n9617), .A2(n6710), .ZN(n5976) );
  OR2_X1 U7444 ( .A1(n9831), .A2(n6345), .ZN(n5979) );
  NAND2_X1 U7445 ( .A1(n5980), .A2(n5979), .ZN(n5981) );
  XNOR2_X1 U7446 ( .A(n5981), .B(n7304), .ZN(n5986) );
  AOI22_X1 U7447 ( .A1(n9035), .A2(n6394), .B1(n7321), .B2(n6067), .ZN(n5987)
         );
  XNOR2_X1 U7448 ( .A(n5986), .B(n5987), .ZN(n6842) );
  INV_X1 U7449 ( .A(n5982), .ZN(n5984) );
  NAND2_X1 U7450 ( .A1(n5984), .A2(n5983), .ZN(n6843) );
  AND2_X1 U7451 ( .A1(n6842), .A2(n6843), .ZN(n5985) );
  INV_X1 U7452 ( .A(n5986), .ZN(n5988) );
  OR2_X1 U7453 ( .A1(n5988), .A2(n5987), .ZN(n5989) );
  AOI21_X1 U7454 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5990) );
  NOR2_X1 U7455 ( .A1(n5990), .A2(n6012), .ZN(n9753) );
  NAND2_X1 U7456 ( .A1(n5952), .A2(n9753), .ZN(n5999) );
  INV_X1 U7457 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5992) );
  OR2_X1 U7458 ( .A1(n4478), .A2(n5992), .ZN(n5998) );
  INV_X1 U7459 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5994) );
  OR2_X1 U7460 ( .A1(n6537), .A2(n5994), .ZN(n5997) );
  INV_X1 U7461 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5995) );
  OR2_X1 U7462 ( .A1(n4479), .A2(n5995), .ZN(n5996) );
  NAND2_X1 U7463 ( .A1(n9844), .A2(n6067), .ZN(n6008) );
  INV_X1 U7464 ( .A(n6001), .ZN(n6504) );
  INV_X1 U7465 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6505) );
  OR2_X1 U7466 ( .A1(n8855), .A2(n6505), .ZN(n6005) );
  NOR2_X1 U7467 ( .A1(n6002), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6020) );
  OR2_X1 U7468 ( .A1(n6020), .A2(n5860), .ZN(n6003) );
  XNOR2_X1 U7469 ( .A(n6003), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6741) );
  INV_X1 U7470 ( .A(n6741), .ZN(n6727) );
  OR2_X1 U7471 ( .A1(n9617), .A2(n6727), .ZN(n6004) );
  OR2_X1 U7472 ( .A1(n9839), .A2(n6345), .ZN(n6007) );
  NAND2_X1 U7473 ( .A1(n6008), .A2(n6007), .ZN(n6009) );
  XNOR2_X1 U7474 ( .A(n6009), .B(n7776), .ZN(n7090) );
  NAND2_X1 U7475 ( .A1(n9844), .A2(n6394), .ZN(n6011) );
  OR2_X1 U7476 ( .A1(n9839), .A2(n6000), .ZN(n6010) );
  AND2_X1 U7477 ( .A1(n6011), .A2(n6010), .ZN(n7094) );
  NAND2_X1 U7478 ( .A1(n8751), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6017) );
  INV_X1 U7479 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6744) );
  OR2_X1 U7480 ( .A1(n4478), .A2(n6744), .ZN(n6016) );
  OAI21_X1 U7481 ( .B1(n6012), .B2(P1_REG3_REG_6__SCAN_IN), .A(n6039), .ZN(
        n7407) );
  OR2_X1 U7482 ( .A1(n5929), .A2(n7407), .ZN(n6015) );
  INV_X1 U7483 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6013) );
  OR2_X1 U7484 ( .A1(n4479), .A2(n6013), .ZN(n6014) );
  NAND4_X1 U7485 ( .A1(n6017), .A2(n6016), .A3(n6015), .A4(n6014), .ZN(n9855)
         );
  NAND2_X1 U7486 ( .A1(n9855), .A2(n6067), .ZN(n6026) );
  NAND2_X1 U7487 ( .A1(n6048), .A2(n6506), .ZN(n6024) );
  INV_X1 U7488 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U7489 ( .A1(n6020), .A2(n6019), .ZN(n6046) );
  NAND2_X1 U7490 ( .A1(n6046), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6021) );
  XNOR2_X1 U7491 ( .A(n6021), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9654) );
  INV_X1 U7492 ( .A(n9654), .ZN(n6508) );
  OR2_X1 U7493 ( .A1(n9617), .A2(n6508), .ZN(n6023) );
  INV_X1 U7494 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10397) );
  OR2_X1 U7495 ( .A1(n8855), .A2(n10397), .ZN(n6022) );
  OR2_X1 U7496 ( .A1(n9847), .A2(n6345), .ZN(n6025) );
  NAND2_X1 U7497 ( .A1(n6026), .A2(n6025), .ZN(n6027) );
  XNOR2_X1 U7498 ( .A(n6027), .B(n7304), .ZN(n6032) );
  NAND2_X1 U7499 ( .A1(n9855), .A2(n6394), .ZN(n6029) );
  OR2_X1 U7500 ( .A1(n9847), .A2(n6000), .ZN(n6028) );
  NAND2_X1 U7501 ( .A1(n6029), .A2(n6028), .ZN(n6033) );
  NAND2_X1 U7502 ( .A1(n6032), .A2(n6033), .ZN(n7193) );
  OAI21_X1 U7503 ( .B1(n7090), .B2(n7094), .A(n7193), .ZN(n6030) );
  INV_X1 U7504 ( .A(n6032), .ZN(n6035) );
  INV_X1 U7505 ( .A(n6033), .ZN(n6034) );
  AND2_X1 U7506 ( .A1(n6035), .A2(n6034), .ZN(n7194) );
  NAND2_X1 U7507 ( .A1(n8750), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6045) );
  INV_X1 U7508 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n6037) );
  OR2_X1 U7509 ( .A1(n6537), .A2(n6037), .ZN(n6044) );
  AND2_X1 U7510 ( .A1(n6039), .A2(n6038), .ZN(n6040) );
  OR2_X1 U7511 ( .A1(n6040), .A2(n6060), .ZN(n7334) );
  OR2_X1 U7512 ( .A1(n7784), .A2(n7334), .ZN(n6043) );
  INV_X1 U7513 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6041) );
  OR2_X1 U7514 ( .A1(n4479), .A2(n6041), .ZN(n6042) );
  NAND4_X1 U7515 ( .A1(n6045), .A2(n6044), .A3(n6043), .A4(n6042), .ZN(n9843)
         );
  NAND2_X1 U7516 ( .A1(n9843), .A2(n6394), .ZN(n6052) );
  NAND2_X1 U7517 ( .A1(n6068), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6047) );
  XNOR2_X1 U7518 ( .A(n6047), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6760) );
  AOI22_X1 U7519 ( .A1(n6276), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6485), .B2(
        n6760), .ZN(n6050) );
  NAND2_X1 U7520 ( .A1(n6510), .A2(n6048), .ZN(n6049) );
  OR2_X1 U7521 ( .A1(n9861), .A2(n6000), .ZN(n6051) );
  AND2_X1 U7522 ( .A1(n6052), .A2(n6051), .ZN(n7035) );
  NAND2_X1 U7523 ( .A1(n9843), .A2(n6067), .ZN(n6054) );
  OR2_X1 U7524 ( .A1(n9861), .A2(n6345), .ZN(n6053) );
  NAND2_X1 U7525 ( .A1(n6054), .A2(n6053), .ZN(n6055) );
  XNOR2_X1 U7526 ( .A(n6055), .B(n7304), .ZN(n7036) );
  NAND2_X1 U7527 ( .A1(n6056), .A2(n7036), .ZN(n6059) );
  NAND2_X1 U7528 ( .A1(n6057), .A2(n4978), .ZN(n6058) );
  NAND2_X1 U7529 ( .A1(n6059), .A2(n6058), .ZN(n7210) );
  NAND2_X1 U7530 ( .A1(n8751), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6066) );
  INV_X1 U7531 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6746) );
  OR2_X1 U7532 ( .A1(n4478), .A2(n6746), .ZN(n6065) );
  NAND2_X1 U7533 ( .A1(n6060), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6088) );
  OR2_X1 U7534 ( .A1(n6060), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7535 ( .A1(n6088), .A2(n6061), .ZN(n9739) );
  OR2_X1 U7536 ( .A1(n5929), .A2(n9739), .ZN(n6064) );
  INV_X1 U7537 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6062) );
  OR2_X1 U7538 ( .A1(n4479), .A2(n6062), .ZN(n6063) );
  NAND2_X1 U7539 ( .A1(n6518), .A2(n6048), .ZN(n6071) );
  NAND2_X1 U7540 ( .A1(n6069), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6081) );
  XNOR2_X1 U7541 ( .A(n6081), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6892) );
  AOI22_X1 U7542 ( .A1(n6276), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6485), .B2(
        n6892), .ZN(n6070) );
  NAND2_X1 U7543 ( .A1(n6071), .A2(n6070), .ZN(n7322) );
  NAND2_X1 U7544 ( .A1(n7322), .A2(n7773), .ZN(n6072) );
  OAI21_X1 U7545 ( .B1(n7348), .B2(n6000), .A(n6072), .ZN(n6073) );
  XNOR2_X1 U7546 ( .A(n6073), .B(n7776), .ZN(n7212) );
  OR2_X1 U7547 ( .A1(n7348), .A2(n7779), .ZN(n6075) );
  NAND2_X1 U7548 ( .A1(n7322), .A2(n6067), .ZN(n6074) );
  AND2_X1 U7549 ( .A1(n6075), .A2(n6074), .ZN(n7211) );
  NAND2_X1 U7550 ( .A1(n7212), .A2(n7211), .ZN(n6076) );
  INV_X1 U7551 ( .A(n7212), .ZN(n6078) );
  INV_X1 U7552 ( .A(n7211), .ZN(n6077) );
  NAND2_X1 U7553 ( .A1(n6078), .A2(n6077), .ZN(n6079) );
  NAND2_X1 U7554 ( .A1(n6529), .A2(n6048), .ZN(n6085) );
  NAND2_X1 U7555 ( .A1(n6081), .A2(n10452), .ZN(n6082) );
  NAND2_X1 U7556 ( .A1(n6082), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6083) );
  AOI22_X1 U7557 ( .A1(n6276), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6485), .B2(
        n9672), .ZN(n6084) );
  NAND2_X2 U7558 ( .A1(n6085), .A2(n6084), .ZN(n9879) );
  NAND2_X1 U7559 ( .A1(n9879), .A2(n7773), .ZN(n6096) );
  NAND2_X1 U7560 ( .A1(n8750), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6094) );
  INV_X1 U7561 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n6086) );
  OR2_X1 U7562 ( .A1(n6537), .A2(n6086), .ZN(n6093) );
  NAND2_X1 U7563 ( .A1(n6088), .A2(n6087), .ZN(n6089) );
  NAND2_X1 U7564 ( .A1(n6109), .A2(n6089), .ZN(n7349) );
  OR2_X1 U7565 ( .A1(n7784), .A2(n7349), .ZN(n6092) );
  INV_X1 U7566 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6090) );
  OR2_X1 U7567 ( .A1(n4479), .A2(n6090), .ZN(n6091) );
  NAND4_X1 U7568 ( .A1(n6094), .A2(n6093), .A3(n6092), .A4(n6091), .ZN(n9034)
         );
  NAND2_X1 U7569 ( .A1(n9034), .A2(n6067), .ZN(n6095) );
  NAND2_X1 U7570 ( .A1(n6096), .A2(n6095), .ZN(n6097) );
  XNOR2_X1 U7571 ( .A(n6097), .B(n7776), .ZN(n6099) );
  AND2_X1 U7572 ( .A1(n9034), .A2(n6394), .ZN(n6098) );
  AOI21_X1 U7573 ( .B1(n9879), .B2(n6067), .A(n6098), .ZN(n6100) );
  NAND2_X1 U7574 ( .A1(n6099), .A2(n6100), .ZN(n6105) );
  INV_X1 U7575 ( .A(n6099), .ZN(n6102) );
  INV_X1 U7576 ( .A(n6100), .ZN(n6101) );
  NAND2_X1 U7577 ( .A1(n6102), .A2(n6101), .ZN(n6103) );
  NAND2_X1 U7578 ( .A1(n6105), .A2(n6103), .ZN(n7347) );
  NAND2_X1 U7579 ( .A1(n6535), .A2(n6048), .ZN(n6108) );
  NAND2_X1 U7580 ( .A1(n5905), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6106) );
  XNOR2_X1 U7581 ( .A(n6106), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9689) );
  AOI22_X1 U7582 ( .A1(n6276), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6485), .B2(
        n9689), .ZN(n6107) );
  NAND2_X1 U7583 ( .A1(n6108), .A2(n6107), .ZN(n7469) );
  NAND2_X1 U7584 ( .A1(n7469), .A2(n7773), .ZN(n6117) );
  NAND2_X1 U7585 ( .A1(n8751), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6115) );
  INV_X1 U7586 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7362) );
  OR2_X1 U7587 ( .A1(n4478), .A2(n7362), .ZN(n6114) );
  NAND2_X1 U7588 ( .A1(n6109), .A2(n7441), .ZN(n6110) );
  NAND2_X1 U7589 ( .A1(n6126), .A2(n6110), .ZN(n7442) );
  OR2_X1 U7590 ( .A1(n5929), .A2(n7442), .ZN(n6113) );
  INV_X1 U7591 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6111) );
  OR2_X1 U7592 ( .A1(n4479), .A2(n6111), .ZN(n6112) );
  OR2_X1 U7593 ( .A1(n9598), .A2(n6000), .ZN(n6116) );
  NAND2_X1 U7594 ( .A1(n6117), .A2(n6116), .ZN(n6118) );
  XNOR2_X1 U7595 ( .A(n6118), .B(n7776), .ZN(n6121) );
  NOR2_X1 U7596 ( .A1(n9598), .A2(n7779), .ZN(n6119) );
  AOI21_X1 U7597 ( .B1(n7469), .B2(n6067), .A(n6119), .ZN(n6120) );
  OR2_X1 U7598 ( .A1(n6121), .A2(n6120), .ZN(n7435) );
  AND2_X1 U7599 ( .A1(n6121), .A2(n6120), .ZN(n7436) );
  NAND2_X1 U7600 ( .A1(n6548), .A2(n6048), .ZN(n6124) );
  NOR2_X1 U7601 ( .A1(n5905), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6140) );
  OR2_X1 U7602 ( .A1(n6140), .A2(n5860), .ZN(n6122) );
  XNOR2_X1 U7603 ( .A(n6122), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9694) );
  AOI22_X1 U7604 ( .A1(n6276), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6485), .B2(
        n9694), .ZN(n6123) );
  NAND2_X1 U7605 ( .A1(n9601), .A2(n7773), .ZN(n6133) );
  NAND2_X1 U7606 ( .A1(n8751), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6131) );
  INV_X1 U7607 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7474) );
  OR2_X1 U7608 ( .A1(n4478), .A2(n7474), .ZN(n6130) );
  INV_X1 U7609 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6125) );
  AND2_X1 U7610 ( .A1(n6126), .A2(n6125), .ZN(n6127) );
  OR2_X1 U7611 ( .A1(n6127), .A2(n6143), .ZN(n7523) );
  OR2_X1 U7612 ( .A1(n7784), .A2(n7523), .ZN(n6129) );
  INV_X1 U7613 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6894) );
  OR2_X1 U7614 ( .A1(n4479), .A2(n6894), .ZN(n6128) );
  NAND4_X1 U7615 ( .A1(n6131), .A2(n6130), .A3(n6129), .A4(n6128), .ZN(n9033)
         );
  NAND2_X1 U7616 ( .A1(n9033), .A2(n6067), .ZN(n6132) );
  NAND2_X1 U7617 ( .A1(n6133), .A2(n6132), .ZN(n6134) );
  XNOR2_X1 U7618 ( .A(n6134), .B(n7304), .ZN(n6138) );
  AND2_X1 U7619 ( .A1(n9033), .A2(n6394), .ZN(n6135) );
  AOI21_X1 U7620 ( .B1(n9601), .B2(n6067), .A(n6135), .ZN(n6136) );
  XNOR2_X1 U7621 ( .A(n6138), .B(n6136), .ZN(n7521) );
  INV_X1 U7622 ( .A(n6136), .ZN(n6137) );
  NAND2_X1 U7623 ( .A1(n6672), .A2(n6048), .ZN(n6142) );
  AND2_X1 U7624 ( .A1(n6140), .A2(n6139), .ZN(n6178) );
  OR2_X1 U7625 ( .A1(n6178), .A2(n5860), .ZN(n6158) );
  XNOR2_X1 U7626 ( .A(n6158), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7018) );
  AOI22_X1 U7627 ( .A1(n6276), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6485), .B2(
        n7018), .ZN(n6141) );
  NAND2_X1 U7628 ( .A1(n9592), .A2(n7773), .ZN(n6151) );
  NAND2_X1 U7629 ( .A1(n8751), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7630 ( .A1(n6143), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6164) );
  OR2_X1 U7631 ( .A1(n6143), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U7632 ( .A1(n6164), .A2(n6144), .ZN(n9570) );
  OR2_X1 U7633 ( .A1(n5929), .A2(n9570), .ZN(n6148) );
  INV_X1 U7634 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6145) );
  OR2_X1 U7635 ( .A1(n4478), .A2(n6145), .ZN(n6147) );
  INV_X1 U7636 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6889) );
  OR2_X1 U7637 ( .A1(n4479), .A2(n6889), .ZN(n6146) );
  OR2_X1 U7638 ( .A1(n9597), .A2(n6000), .ZN(n6150) );
  NAND2_X1 U7639 ( .A1(n6151), .A2(n6150), .ZN(n6152) );
  XNOR2_X1 U7640 ( .A(n6152), .B(n7776), .ZN(n6155) );
  NOR2_X1 U7641 ( .A1(n9597), .A2(n7779), .ZN(n6153) );
  AOI21_X1 U7642 ( .B1(n9592), .B2(n6067), .A(n6153), .ZN(n6154) );
  XNOR2_X1 U7643 ( .A(n6155), .B(n6154), .ZN(n7580) );
  NAND2_X1 U7644 ( .A1(n6155), .A2(n6154), .ZN(n6156) );
  NAND2_X1 U7645 ( .A1(n6774), .A2(n6048), .ZN(n6162) );
  NAND2_X1 U7646 ( .A1(n6158), .A2(n6157), .ZN(n6159) );
  NAND2_X1 U7647 ( .A1(n6159), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6160) );
  XNOR2_X1 U7648 ( .A(n6160), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7228) );
  AOI22_X1 U7649 ( .A1(n6276), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6485), .B2(
        n7228), .ZN(n6161) );
  NAND2_X1 U7650 ( .A1(n9586), .A2(n7773), .ZN(n6171) );
  NAND2_X1 U7651 ( .A1(n8751), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6169) );
  INV_X1 U7652 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7758) );
  OR2_X1 U7653 ( .A1(n4478), .A2(n7758), .ZN(n6168) );
  INV_X1 U7654 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U7655 ( .A1(n6164), .A2(n6163), .ZN(n6165) );
  NAND2_X1 U7656 ( .A1(n6182), .A2(n6165), .ZN(n7757) );
  OR2_X1 U7657 ( .A1(n7784), .A2(n7757), .ZN(n6167) );
  INV_X1 U7658 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7019) );
  OR2_X1 U7659 ( .A1(n4479), .A2(n7019), .ZN(n6166) );
  NAND4_X1 U7660 ( .A1(n6169), .A2(n6168), .A3(n6167), .A4(n6166), .ZN(n9032)
         );
  NAND2_X1 U7661 ( .A1(n9032), .A2(n6067), .ZN(n6170) );
  NAND2_X1 U7662 ( .A1(n6171), .A2(n6170), .ZN(n6172) );
  XNOR2_X1 U7663 ( .A(n6172), .B(n7776), .ZN(n7587) );
  AND2_X1 U7664 ( .A1(n9032), .A2(n6394), .ZN(n6173) );
  AOI21_X1 U7665 ( .B1(n9586), .B2(n6067), .A(n6173), .ZN(n6174) );
  AND2_X1 U7666 ( .A1(n7587), .A2(n6174), .ZN(n6176) );
  INV_X1 U7667 ( .A(n7587), .ZN(n6175) );
  INV_X1 U7668 ( .A(n6174), .ZN(n7586) );
  NAND2_X1 U7669 ( .A1(n6801), .A2(n6048), .ZN(n6181) );
  NOR2_X1 U7670 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n6177) );
  NAND2_X1 U7671 ( .A1(n6178), .A2(n6177), .ZN(n6195) );
  NAND2_X1 U7672 ( .A1(n6195), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6179) );
  XNOR2_X1 U7673 ( .A(n6179), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7507) );
  AOI22_X1 U7674 ( .A1(n6276), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6485), .B2(
        n7507), .ZN(n6180) );
  NAND2_X1 U7675 ( .A1(n7672), .A2(n7773), .ZN(n6189) );
  NAND2_X1 U7676 ( .A1(n8751), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6187) );
  INV_X1 U7677 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7611) );
  OR2_X1 U7678 ( .A1(n4478), .A2(n7611), .ZN(n6186) );
  INV_X1 U7679 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7219) );
  AND2_X1 U7680 ( .A1(n6182), .A2(n7219), .ZN(n6183) );
  OR2_X1 U7681 ( .A1(n6183), .A2(n6201), .ZN(n7690) );
  OR2_X1 U7682 ( .A1(n5929), .A2(n7690), .ZN(n6185) );
  INV_X1 U7683 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7221) );
  OR2_X1 U7684 ( .A1(n4479), .A2(n7221), .ZN(n6184) );
  NAND4_X1 U7685 ( .A1(n6187), .A2(n6186), .A3(n6185), .A4(n6184), .ZN(n9441)
         );
  NAND2_X1 U7686 ( .A1(n9441), .A2(n6067), .ZN(n6188) );
  NAND2_X1 U7687 ( .A1(n6189), .A2(n6188), .ZN(n6190) );
  XNOR2_X1 U7688 ( .A(n6190), .B(n7304), .ZN(n7686) );
  INV_X1 U7689 ( .A(n7686), .ZN(n6194) );
  NAND2_X1 U7690 ( .A1(n7672), .A2(n6067), .ZN(n6192) );
  NAND2_X1 U7691 ( .A1(n9441), .A2(n6394), .ZN(n6191) );
  NAND2_X1 U7692 ( .A1(n6192), .A2(n6191), .ZN(n7685) );
  INV_X1 U7693 ( .A(n7685), .ZN(n6193) );
  NAND2_X1 U7694 ( .A1(n6194), .A2(n6193), .ZN(n6215) );
  NAND2_X1 U7695 ( .A1(n6874), .A2(n6048), .ZN(n6200) );
  OR2_X1 U7696 ( .A1(n6195), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n6218) );
  NAND2_X1 U7697 ( .A1(n6218), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6197) );
  INV_X1 U7698 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6196) );
  XNOR2_X1 U7699 ( .A(n6197), .B(n6196), .ZN(n7739) );
  INV_X1 U7700 ( .A(n7739), .ZN(n6198) );
  AOI22_X1 U7701 ( .A1(n6276), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6485), .B2(
        n6198), .ZN(n6199) );
  NAND2_X1 U7702 ( .A1(n9443), .A2(n7773), .ZN(n6207) );
  NAND2_X1 U7703 ( .A1(n8751), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6205) );
  INV_X1 U7704 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7677) );
  OR2_X1 U7705 ( .A1(n4478), .A2(n7677), .ZN(n6204) );
  INV_X1 U7706 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7509) );
  OR2_X1 U7707 ( .A1(n4479), .A2(n7509), .ZN(n6203) );
  OAI21_X1 U7708 ( .B1(n6201), .B2(P1_REG3_REG_15__SCAN_IN), .A(n6222), .ZN(
        n8737) );
  OR2_X1 U7709 ( .A1(n7784), .A2(n8737), .ZN(n6202) );
  NAND4_X1 U7710 ( .A1(n6205), .A2(n6204), .A3(n6203), .A4(n6202), .ZN(n9031)
         );
  NAND2_X1 U7711 ( .A1(n9031), .A2(n6067), .ZN(n6206) );
  NAND2_X1 U7712 ( .A1(n6207), .A2(n6206), .ZN(n6208) );
  XNOR2_X1 U7713 ( .A(n6208), .B(n7304), .ZN(n6214) );
  INV_X1 U7714 ( .A(n6214), .ZN(n6210) );
  AND2_X1 U7715 ( .A1(n7686), .A2(n7685), .ZN(n6216) );
  INV_X1 U7716 ( .A(n6216), .ZN(n6209) );
  AND2_X1 U7717 ( .A1(n6210), .A2(n6209), .ZN(n6211) );
  NAND2_X1 U7718 ( .A1(n9443), .A2(n6067), .ZN(n6213) );
  NAND2_X1 U7719 ( .A1(n9031), .A2(n6394), .ZN(n6212) );
  NAND2_X1 U7720 ( .A1(n6213), .A2(n6212), .ZN(n8730) );
  OAI211_X1 U7721 ( .C1(n7688), .C2(n6216), .A(n6215), .B(n6214), .ZN(n8729)
         );
  NAND2_X1 U7722 ( .A1(n6217), .A2(n8729), .ZN(n8645) );
  NAND2_X1 U7723 ( .A1(n6849), .A2(n6048), .ZN(n6220) );
  OAI21_X1 U7724 ( .B1(n6218), .B2(P1_IR_REG_15__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6239) );
  XNOR2_X1 U7725 ( .A(n6239), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7742) );
  AOI22_X1 U7726 ( .A1(n6276), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6485), .B2(
        n7742), .ZN(n6219) );
  NAND2_X1 U7727 ( .A1(n9437), .A2(n7773), .ZN(n6230) );
  NAND2_X1 U7728 ( .A1(n8751), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6228) );
  INV_X1 U7729 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7698) );
  OR2_X1 U7730 ( .A1(n4478), .A2(n7698), .ZN(n6227) );
  INV_X1 U7731 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8651) );
  NAND2_X1 U7732 ( .A1(n6222), .A2(n8651), .ZN(n6223) );
  NAND2_X1 U7733 ( .A1(n6245), .A2(n6223), .ZN(n8653) );
  OR2_X1 U7734 ( .A1(n7784), .A2(n8653), .ZN(n6226) );
  INV_X1 U7735 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n6224) );
  OR2_X1 U7736 ( .A1(n4479), .A2(n6224), .ZN(n6225) );
  OR2_X1 U7737 ( .A1(n9423), .A2(n6000), .ZN(n6229) );
  NAND2_X1 U7738 ( .A1(n6230), .A2(n6229), .ZN(n6231) );
  XNOR2_X1 U7739 ( .A(n6231), .B(n7304), .ZN(n6234) );
  NAND2_X1 U7740 ( .A1(n9437), .A2(n6067), .ZN(n6233) );
  OR2_X1 U7741 ( .A1(n9423), .A2(n7779), .ZN(n6232) );
  NAND2_X1 U7742 ( .A1(n6233), .A2(n6232), .ZN(n6235) );
  AND2_X1 U7743 ( .A1(n6234), .A2(n6235), .ZN(n8646) );
  INV_X1 U7744 ( .A(n6234), .ZN(n6237) );
  INV_X1 U7745 ( .A(n6235), .ZN(n6236) );
  NAND2_X1 U7746 ( .A1(n6237), .A2(n6236), .ZN(n8644) );
  NAND2_X1 U7747 ( .A1(n6886), .A2(n6048), .ZN(n6242) );
  INV_X1 U7748 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6238) );
  NAND2_X1 U7749 ( .A1(n6239), .A2(n6238), .ZN(n6240) );
  NAND2_X1 U7750 ( .A1(n6240), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6260) );
  XNOR2_X1 U7751 ( .A(n6260), .B(P1_IR_REG_17__SCAN_IN), .ZN(n7743) );
  AOI22_X1 U7752 ( .A1(n6276), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6485), .B2(
        n7743), .ZN(n6241) );
  NAND2_X1 U7753 ( .A1(n9317), .A2(n7773), .ZN(n6252) );
  NAND2_X1 U7754 ( .A1(n8751), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6250) );
  INV_X1 U7755 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9321) );
  OR2_X1 U7756 ( .A1(n4478), .A2(n9321), .ZN(n6249) );
  INV_X1 U7757 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6244) );
  NAND2_X1 U7758 ( .A1(n6245), .A2(n6244), .ZN(n6246) );
  NAND2_X1 U7759 ( .A1(n6266), .A2(n6246), .ZN(n9320) );
  OR2_X1 U7760 ( .A1(n7784), .A2(n9320), .ZN(n6248) );
  INV_X1 U7761 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9432) );
  OR2_X1 U7762 ( .A1(n4479), .A2(n9432), .ZN(n6247) );
  NAND4_X1 U7763 ( .A1(n6250), .A2(n6249), .A3(n6248), .A4(n6247), .ZN(n9414)
         );
  NAND2_X1 U7764 ( .A1(n9414), .A2(n6067), .ZN(n6251) );
  NAND2_X1 U7765 ( .A1(n6252), .A2(n6251), .ZN(n6253) );
  XNOR2_X1 U7766 ( .A(n6253), .B(n7304), .ZN(n6255) );
  AND2_X1 U7767 ( .A1(n9414), .A2(n6394), .ZN(n6254) );
  AOI21_X1 U7768 ( .B1(n9317), .B2(n6067), .A(n6254), .ZN(n6256) );
  XNOR2_X1 U7769 ( .A(n6255), .B(n6256), .ZN(n8659) );
  INV_X1 U7770 ( .A(n6255), .ZN(n6257) );
  NAND2_X1 U7771 ( .A1(n6257), .A2(n6256), .ZN(n6258) );
  NAND2_X1 U7772 ( .A1(n7077), .A2(n6048), .ZN(n6264) );
  NAND2_X1 U7773 ( .A1(n6260), .A2(n6259), .ZN(n6261) );
  NAND2_X1 U7774 ( .A1(n6261), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6262) );
  XNOR2_X1 U7775 ( .A(n6262), .B(P1_IR_REG_18__SCAN_IN), .ZN(n7744) );
  AOI22_X1 U7776 ( .A1(n6276), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6485), .B2(
        n7744), .ZN(n6263) );
  NAND2_X1 U7777 ( .A1(n9307), .A2(n7773), .ZN(n6273) );
  NAND2_X1 U7778 ( .A1(n8751), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6271) );
  INV_X1 U7779 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9299) );
  OR2_X1 U7780 ( .A1(n4478), .A2(n9299), .ZN(n6270) );
  INV_X1 U7781 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6265) );
  NAND2_X1 U7782 ( .A1(n6266), .A2(n6265), .ZN(n6267) );
  NAND2_X1 U7783 ( .A1(n6280), .A2(n6267), .ZN(n9298) );
  OR2_X1 U7784 ( .A1(n9298), .A2(n7784), .ZN(n6269) );
  INV_X1 U7785 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9421) );
  OR2_X1 U7786 ( .A1(n4479), .A2(n9421), .ZN(n6268) );
  INV_X1 U7787 ( .A(n9424), .ZN(n9324) );
  NAND2_X1 U7788 ( .A1(n9324), .A2(n6067), .ZN(n6272) );
  NAND2_X1 U7789 ( .A1(n6273), .A2(n6272), .ZN(n6274) );
  XNOR2_X1 U7790 ( .A(n6274), .B(n7776), .ZN(n6275) );
  INV_X1 U7791 ( .A(n9307), .ZN(n9490) );
  OAI22_X1 U7792 ( .A1(n9490), .A2(n6000), .B1(n9424), .B2(n7779), .ZN(n8706)
         );
  NAND2_X1 U7793 ( .A1(n7148), .A2(n6048), .ZN(n6278) );
  AOI22_X1 U7794 ( .A1(n6276), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n8871), .B2(
        n6485), .ZN(n6277) );
  INV_X1 U7795 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8624) );
  NAND2_X1 U7796 ( .A1(n6280), .A2(n8624), .ZN(n6281) );
  NAND2_X1 U7797 ( .A1(n6293), .A2(n6281), .ZN(n9284) );
  NOR2_X1 U7798 ( .A1(n9284), .A2(n7784), .ZN(n6285) );
  INV_X1 U7799 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9412) );
  NOR2_X1 U7800 ( .A1(n4479), .A2(n9412), .ZN(n6284) );
  INV_X1 U7801 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9285) );
  NAND2_X1 U7802 ( .A1(n8751), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6282) );
  OAI21_X1 U7803 ( .B1(n9285), .B2(n4478), .A(n6282), .ZN(n6283) );
  OAI22_X1 U7804 ( .A1(n9486), .A2(n6000), .B1(n9265), .B2(n7779), .ZN(n6287)
         );
  OAI22_X1 U7805 ( .A1(n9486), .A2(n6345), .B1(n9265), .B2(n6000), .ZN(n6286)
         );
  XNOR2_X1 U7806 ( .A(n6286), .B(n7304), .ZN(n6288) );
  XOR2_X1 U7807 ( .A(n6287), .B(n6288), .Z(n8623) );
  INV_X1 U7808 ( .A(n6287), .ZN(n6290) );
  INV_X1 U7809 ( .A(n6288), .ZN(n6289) );
  NAND2_X1 U7810 ( .A1(n7233), .A2(n6048), .ZN(n6292) );
  OR2_X1 U7811 ( .A1(n8855), .A2(n10451), .ZN(n6291) );
  NAND2_X1 U7812 ( .A1(n9406), .A2(n7773), .ZN(n6302) );
  INV_X1 U7813 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8678) );
  NAND2_X1 U7814 ( .A1(n6293), .A2(n8678), .ZN(n6294) );
  AND2_X1 U7815 ( .A1(n6311), .A2(n6294), .ZN(n9269) );
  NAND2_X1 U7816 ( .A1(n9269), .A2(n5952), .ZN(n6300) );
  INV_X1 U7817 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n6297) );
  NAND2_X1 U7818 ( .A1(n8751), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U7819 ( .A1(n8750), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6295) );
  OAI211_X1 U7820 ( .C1(n6297), .C2(n4479), .A(n6296), .B(n6295), .ZN(n6298)
         );
  INV_X1 U7821 ( .A(n6298), .ZN(n6299) );
  NAND2_X1 U7822 ( .A1(n6300), .A2(n6299), .ZN(n9106) );
  NAND2_X1 U7823 ( .A1(n9106), .A2(n6067), .ZN(n6301) );
  NAND2_X1 U7824 ( .A1(n6302), .A2(n6301), .ZN(n6303) );
  XNOR2_X1 U7825 ( .A(n6303), .B(n7776), .ZN(n6306) );
  AND2_X1 U7826 ( .A1(n9106), .A2(n6394), .ZN(n6304) );
  AOI21_X1 U7827 ( .B1(n9406), .B2(n6067), .A(n6304), .ZN(n6305) );
  NOR2_X1 U7828 ( .A1(n6306), .A2(n6305), .ZN(n8675) );
  NAND2_X1 U7829 ( .A1(n6306), .A2(n6305), .ZN(n8674) );
  NAND2_X1 U7830 ( .A1(n7302), .A2(n6048), .ZN(n6308) );
  OR2_X1 U7831 ( .A1(n8855), .A2(n7303), .ZN(n6307) );
  INV_X1 U7832 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6310) );
  NAND2_X1 U7833 ( .A1(n6311), .A2(n6310), .ZN(n6312) );
  NAND2_X1 U7834 ( .A1(n6328), .A2(n6312), .ZN(n9250) );
  OR2_X1 U7835 ( .A1(n9250), .A2(n7784), .ZN(n6318) );
  INV_X1 U7836 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n6315) );
  NAND2_X1 U7837 ( .A1(n8751), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6314) );
  NAND2_X1 U7838 ( .A1(n8750), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6313) );
  OAI211_X1 U7839 ( .C1(n6315), .C2(n4479), .A(n6314), .B(n6313), .ZN(n6316)
         );
  INV_X1 U7840 ( .A(n6316), .ZN(n6317) );
  OAI22_X1 U7841 ( .A1(n9256), .A2(n6000), .B1(n9266), .B2(n7779), .ZN(n6323)
         );
  NAND2_X1 U7842 ( .A1(n9400), .A2(n7773), .ZN(n6320) );
  INV_X1 U7843 ( .A(n9266), .ZN(n9385) );
  NAND2_X1 U7844 ( .A1(n9385), .A2(n6067), .ZN(n6319) );
  NAND2_X1 U7845 ( .A1(n6320), .A2(n6319), .ZN(n6321) );
  XNOR2_X1 U7846 ( .A(n6321), .B(n7304), .ZN(n6322) );
  XOR2_X1 U7847 ( .A(n6323), .B(n6322), .Z(n8630) );
  INV_X1 U7848 ( .A(n6322), .ZN(n6325) );
  INV_X1 U7849 ( .A(n6323), .ZN(n6324) );
  NAND2_X1 U7850 ( .A1(n7433), .A2(n6048), .ZN(n6327) );
  OR2_X1 U7851 ( .A1(n8855), .A2(n10434), .ZN(n6326) );
  INV_X1 U7852 ( .A(n9239), .ZN(n9480) );
  INV_X1 U7853 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8689) );
  NAND2_X1 U7854 ( .A1(n6328), .A2(n8689), .ZN(n6329) );
  NAND2_X1 U7855 ( .A1(n6340), .A2(n6329), .ZN(n9231) );
  OR2_X1 U7856 ( .A1(n9231), .A2(n7784), .ZN(n6334) );
  INV_X1 U7857 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9392) );
  NAND2_X1 U7858 ( .A1(n8750), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6331) );
  NAND2_X1 U7859 ( .A1(n8751), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6330) );
  OAI211_X1 U7860 ( .C1(n9392), .C2(n4479), .A(n6331), .B(n6330), .ZN(n6332)
         );
  INV_X1 U7861 ( .A(n6332), .ZN(n6333) );
  NAND2_X1 U7862 ( .A1(n6334), .A2(n6333), .ZN(n9254) );
  INV_X1 U7863 ( .A(n9254), .ZN(n9397) );
  OAI22_X1 U7864 ( .A1(n9480), .A2(n6000), .B1(n9397), .B2(n7779), .ZN(n6336)
         );
  AOI22_X1 U7865 ( .A1(n9239), .A2(n7773), .B1(n6067), .B2(n9254), .ZN(n6335)
         );
  XNOR2_X1 U7866 ( .A(n6335), .B(n7304), .ZN(n8686) );
  NOR2_X1 U7867 ( .A1(n8685), .A2(n8686), .ZN(n6348) );
  NAND2_X1 U7868 ( .A1(n7486), .A2(n6048), .ZN(n6338) );
  OR2_X1 U7869 ( .A1(n8855), .A2(n10465), .ZN(n6337) );
  INV_X1 U7870 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6339) );
  NAND2_X1 U7871 ( .A1(n6340), .A2(n6339), .ZN(n6341) );
  AND2_X1 U7872 ( .A1(n6353), .A2(n6341), .ZN(n9218) );
  INV_X1 U7873 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9383) );
  NAND2_X1 U7874 ( .A1(n8750), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6343) );
  NAND2_X1 U7875 ( .A1(n8751), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6342) );
  OAI211_X1 U7876 ( .C1(n4479), .C2(n9383), .A(n6343), .B(n6342), .ZN(n6344)
         );
  AOI21_X1 U7877 ( .B1(n9218), .B2(n5952), .A(n6344), .ZN(n9207) );
  OAI22_X1 U7878 ( .A1(n9476), .A2(n6345), .B1(n9207), .B2(n6000), .ZN(n6346)
         );
  XNOR2_X1 U7879 ( .A(n6346), .B(n7304), .ZN(n6347) );
  INV_X1 U7880 ( .A(n9207), .ZN(n9386) );
  AOI22_X1 U7881 ( .A1(n9221), .A2(n6067), .B1(n6394), .B2(n9386), .ZN(n8615)
         );
  OAI21_X1 U7882 ( .B1(n6348), .B2(n8684), .A(n6347), .ZN(n8614) );
  NAND2_X1 U7883 ( .A1(n7543), .A2(n6048), .ZN(n6350) );
  INV_X1 U7884 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10368) );
  OR2_X1 U7885 ( .A1(n8855), .A2(n10368), .ZN(n6349) );
  NAND2_X1 U7886 ( .A1(n9210), .A2(n7773), .ZN(n6362) );
  INV_X1 U7887 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6352) );
  NAND2_X1 U7888 ( .A1(n6353), .A2(n6352), .ZN(n6354) );
  NAND2_X1 U7889 ( .A1(n6371), .A2(n6354), .ZN(n8668) );
  OR2_X1 U7890 ( .A1(n8668), .A2(n7784), .ZN(n6360) );
  INV_X1 U7891 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6357) );
  NAND2_X1 U7892 ( .A1(n8750), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U7893 ( .A1(n8751), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6355) );
  OAI211_X1 U7894 ( .C1(n4479), .C2(n6357), .A(n6356), .B(n6355), .ZN(n6358)
         );
  INV_X1 U7895 ( .A(n6358), .ZN(n6359) );
  NAND2_X1 U7896 ( .A1(n9215), .A2(n6067), .ZN(n6361) );
  NAND2_X1 U7897 ( .A1(n6362), .A2(n6361), .ZN(n6363) );
  XNOR2_X1 U7898 ( .A(n6363), .B(n7776), .ZN(n6366) );
  AND2_X1 U7899 ( .A1(n9215), .A2(n6394), .ZN(n6364) );
  AOI21_X1 U7900 ( .B1(n9210), .B2(n6067), .A(n6364), .ZN(n6365) );
  NAND2_X1 U7901 ( .A1(n6366), .A2(n6365), .ZN(n6367) );
  OAI21_X1 U7902 ( .B1(n6366), .B2(n6365), .A(n6367), .ZN(n8666) );
  OR2_X1 U7903 ( .A1(n8855), .A2(n10437), .ZN(n6368) );
  NAND2_X1 U7904 ( .A1(n9192), .A2(n7773), .ZN(n6379) );
  INV_X1 U7905 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6370) );
  NAND2_X1 U7906 ( .A1(n6371), .A2(n6370), .ZN(n6372) );
  NAND2_X1 U7907 ( .A1(n6386), .A2(n6372), .ZN(n8638) );
  OR2_X1 U7908 ( .A1(n8638), .A2(n7784), .ZN(n6377) );
  INV_X1 U7909 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9370) );
  NAND2_X1 U7910 ( .A1(n8751), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6374) );
  NAND2_X1 U7911 ( .A1(n8750), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6373) );
  OAI211_X1 U7912 ( .C1(n9370), .C2(n4479), .A(n6374), .B(n6373), .ZN(n6375)
         );
  INV_X1 U7913 ( .A(n6375), .ZN(n6376) );
  NAND2_X1 U7914 ( .A1(n9372), .A2(n6067), .ZN(n6378) );
  NAND2_X1 U7915 ( .A1(n6379), .A2(n6378), .ZN(n6380) );
  XNOR2_X1 U7916 ( .A(n6380), .B(n7304), .ZN(n6382) );
  OAI22_X1 U7917 ( .A1(n9471), .A2(n6000), .B1(n9204), .B2(n7779), .ZN(n6381)
         );
  XNOR2_X1 U7918 ( .A(n6382), .B(n6381), .ZN(n8636) );
  NOR2_X1 U7919 ( .A1(n6382), .A2(n6381), .ZN(n8716) );
  OR2_X1 U7920 ( .A1(n8855), .A2(n10449), .ZN(n6383) );
  INV_X1 U7921 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6385) );
  NAND2_X1 U7922 ( .A1(n6386), .A2(n6385), .ZN(n6387) );
  NAND2_X1 U7923 ( .A1(n9174), .A2(n5952), .ZN(n6393) );
  INV_X1 U7924 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n6390) );
  NAND2_X1 U7925 ( .A1(n8750), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6389) );
  NAND2_X1 U7926 ( .A1(n8751), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6388) );
  OAI211_X1 U7927 ( .C1(n6390), .C2(n4479), .A(n6389), .B(n6388), .ZN(n6391)
         );
  INV_X1 U7928 ( .A(n6391), .ZN(n6392) );
  AND2_X1 U7929 ( .A1(n9186), .A2(n6394), .ZN(n6395) );
  AOI21_X1 U7930 ( .B1(n9364), .B2(n6067), .A(n6395), .ZN(n6399) );
  NAND2_X1 U7931 ( .A1(n9364), .A2(n7773), .ZN(n6397) );
  NAND2_X1 U7932 ( .A1(n9186), .A2(n6067), .ZN(n6396) );
  NAND2_X1 U7933 ( .A1(n6397), .A2(n6396), .ZN(n6398) );
  XNOR2_X1 U7934 ( .A(n6398), .B(n7304), .ZN(n6401) );
  XOR2_X1 U7935 ( .A(n6399), .B(n6401), .Z(n8715) );
  INV_X1 U7936 ( .A(n6399), .ZN(n6400) );
  OR2_X1 U7937 ( .A1(n8855), .A2(n10272), .ZN(n6402) );
  NAND2_X1 U7938 ( .A1(n9162), .A2(n7773), .ZN(n6410) );
  XNOR2_X1 U7939 ( .A(n6455), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9157) );
  NAND2_X1 U7940 ( .A1(n9157), .A2(n5952), .ZN(n6408) );
  INV_X1 U7941 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9360) );
  NAND2_X1 U7942 ( .A1(n8750), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6405) );
  NAND2_X1 U7943 ( .A1(n8751), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6404) );
  OAI211_X1 U7944 ( .C1(n4479), .C2(n9360), .A(n6405), .B(n6404), .ZN(n6406)
         );
  INV_X1 U7945 ( .A(n6406), .ZN(n6407) );
  INV_X1 U7946 ( .A(n9172), .ZN(n9030) );
  NAND2_X1 U7947 ( .A1(n9030), .A2(n6067), .ZN(n6409) );
  NAND2_X1 U7948 ( .A1(n6410), .A2(n6409), .ZN(n6411) );
  XNOR2_X1 U7949 ( .A(n6411), .B(n7776), .ZN(n6414) );
  NOR2_X1 U7950 ( .A1(n9172), .A2(n7779), .ZN(n6412) );
  AOI21_X1 U7951 ( .B1(n9162), .B2(n6067), .A(n6412), .ZN(n6413) );
  NAND2_X1 U7952 ( .A1(n6414), .A2(n6413), .ZN(n7793) );
  OAI21_X1 U7953 ( .B1(n6414), .B2(n6413), .A(n7793), .ZN(n6415) );
  OAI21_X1 U7954 ( .B1(n8714), .B2(n6416), .A(n6415), .ZN(n6417) );
  INV_X1 U7955 ( .A(n6417), .ZN(n6441) );
  INV_X1 U7956 ( .A(n7544), .ZN(n6419) );
  INV_X1 U7957 ( .A(P1_B_REG_SCAN_IN), .ZN(n6418) );
  AND2_X1 U7958 ( .A1(n6419), .A2(n6418), .ZN(n6421) );
  AND3_X1 U7959 ( .A1(n7620), .A2(P1_B_REG_SCAN_IN), .A3(n7544), .ZN(n6420) );
  INV_X1 U7960 ( .A(n7635), .ZN(n6423) );
  INV_X1 U7961 ( .A(n7620), .ZN(n6422) );
  OAI22_X1 U7962 ( .A1(n7130), .A2(P1_D_REG_1__SCAN_IN), .B1(n6423), .B2(n6422), .ZN(n7492) );
  INV_X1 U7963 ( .A(n7492), .ZN(n6436) );
  INV_X1 U7964 ( .A(n7130), .ZN(n7128) );
  NOR4_X1 U7965 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6427) );
  NOR4_X1 U7966 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6426) );
  NOR4_X1 U7967 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6425) );
  NOR4_X1 U7968 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6424) );
  NAND4_X1 U7969 ( .A1(n6427), .A2(n6426), .A3(n6425), .A4(n6424), .ZN(n6433)
         );
  NOR2_X1 U7970 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .ZN(
        n6431) );
  NOR4_X1 U7971 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6430) );
  NOR4_X1 U7972 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6429) );
  NOR4_X1 U7973 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6428) );
  NAND4_X1 U7974 ( .A1(n6431), .A2(n6430), .A3(n6429), .A4(n6428), .ZN(n6432)
         );
  NOR2_X1 U7975 ( .A1(n6433), .A2(n6432), .ZN(n7126) );
  NAND2_X1 U7976 ( .A1(n7126), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6434) );
  NAND2_X1 U7977 ( .A1(n7128), .A2(n6434), .ZN(n6435) );
  NAND2_X1 U7978 ( .A1(n7635), .A2(n7544), .ZN(n7129) );
  AND2_X1 U7979 ( .A1(n6435), .A2(n7129), .ZN(n7493) );
  NAND2_X1 U7980 ( .A1(n6436), .A2(n7493), .ZN(n6447) );
  NAND2_X1 U7981 ( .A1(n4555), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6438) );
  XNOR2_X1 U7982 ( .A(n6438), .B(n6437), .ZN(n7487) );
  AND2_X1 U7983 ( .A1(n7487), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6439) );
  INV_X1 U7984 ( .A(n9810), .ZN(n9023) );
  OR2_X1 U7985 ( .A1(n6447), .A2(n9023), .ZN(n6465) );
  NAND2_X1 U7986 ( .A1(n7434), .A2(n9013), .ZN(n9797) );
  NAND2_X1 U7987 ( .A1(n9024), .A2(n8947), .ZN(n8872) );
  NAND2_X1 U7988 ( .A1(n9869), .A2(n8872), .ZN(n6440) );
  OAI21_X1 U7989 ( .B1(n7800), .B2(n6441), .A(n8732), .ZN(n6470) );
  NAND2_X1 U7990 ( .A1(n6447), .A2(n9869), .ZN(n6584) );
  OR2_X1 U7991 ( .A1(n8872), .A2(n6442), .ZN(n7489) );
  AND3_X1 U7992 ( .A1(n6443), .A2(n7487), .A3(n7489), .ZN(n6444) );
  AOI21_X1 U7993 ( .B1(n6584), .B2(n6444), .A(P1_U3084), .ZN(n6448) );
  OR2_X1 U7994 ( .A1(n9797), .A2(n7234), .ZN(n9755) );
  INV_X1 U7995 ( .A(n9755), .ZN(n6445) );
  AND2_X1 U7996 ( .A1(n9810), .A2(n6445), .ZN(n6446) );
  AND2_X1 U7997 ( .A1(n6447), .A2(n6446), .ZN(n6583) );
  OR2_X1 U7998 ( .A1(n6448), .A2(n6583), .ZN(n8721) );
  NAND3_X1 U7999 ( .A1(n6449), .A2(n9024), .A3(n9761), .ZN(n9791) );
  NOR2_X1 U8000 ( .A1(n6465), .A2(n9791), .ZN(n6462) );
  INV_X1 U8001 ( .A(n4480), .ZN(n7137) );
  NAND2_X1 U8002 ( .A1(n6462), .A2(n7137), .ZN(n8723) );
  INV_X1 U8003 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6454) );
  OAI22_X1 U8004 ( .A1(n9153), .A2(n8723), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6454), .ZN(n6464) );
  INV_X1 U8005 ( .A(n6455), .ZN(n6452) );
  AND2_X1 U8006 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6451) );
  NAND2_X1 U8007 ( .A1(n6452), .A2(n6451), .ZN(n9127) );
  INV_X1 U8008 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6453) );
  OAI21_X1 U8009 ( .B1(n6455), .B2(n6454), .A(n6453), .ZN(n6456) );
  NAND2_X1 U8010 ( .A1(n9127), .A2(n6456), .ZN(n7783) );
  OR2_X1 U8011 ( .A1(n7783), .A2(n7784), .ZN(n6461) );
  INV_X1 U8012 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9350) );
  NAND2_X1 U8013 ( .A1(n8750), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6458) );
  NAND2_X1 U8014 ( .A1(n8751), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6457) );
  OAI211_X1 U8015 ( .C1(n9350), .C2(n4479), .A(n6458), .B(n6457), .ZN(n6459)
         );
  INV_X1 U8016 ( .A(n6459), .ZN(n6460) );
  NAND2_X1 U8017 ( .A1(n6462), .A2(n4480), .ZN(n8735) );
  NOR2_X1 U8018 ( .A1(n9356), .A2(n8735), .ZN(n6463) );
  AOI211_X1 U8019 ( .C1(n9157), .C2(n8721), .A(n6464), .B(n6463), .ZN(n6469)
         );
  OR2_X1 U8020 ( .A1(n6465), .A2(n9755), .ZN(n6467) );
  NAND2_X1 U8021 ( .A1(n9875), .A2(n9013), .ZN(n7490) );
  INV_X1 U8022 ( .A(n7490), .ZN(n6466) );
  NAND2_X1 U8023 ( .A1(n6467), .A2(n9319), .ZN(n8710) );
  NAND2_X1 U8024 ( .A1(n9162), .A2(n8710), .ZN(n6468) );
  NAND3_X1 U8025 ( .A1(n6470), .A2(n6469), .A3(n6468), .ZN(P1_U3212) );
  NAND2_X1 U8026 ( .A1(n6471), .A2(n7487), .ZN(n6637) );
  OR2_X2 U8027 ( .A1(n6637), .A2(P1_U3084), .ZN(n9036) );
  INV_X1 U8028 ( .A(n9962), .ZN(n6472) );
  OR2_X2 U8029 ( .A1(n6554), .A2(n6472), .ZN(n8166) );
  INV_X1 U8030 ( .A(n8166), .ZN(P2_U3966) );
  XNOR2_X1 U8031 ( .A(n6473), .B(n6474), .ZN(n6475) );
  NOR2_X1 U8032 ( .A1(n6475), .A2(n8145), .ZN(n6482) );
  NOR2_X1 U8033 ( .A1(n8123), .A2(n4883), .ZN(n6481) );
  NOR2_X1 U8034 ( .A1(n8128), .A2(n7072), .ZN(n6480) );
  OR2_X1 U8035 ( .A1(n7114), .A2(n8428), .ZN(n6477) );
  OR2_X1 U8036 ( .A1(n7062), .A2(n8426), .ZN(n6476) );
  NAND2_X1 U8037 ( .A1(n6477), .A2(n6476), .ZN(n7069) );
  INV_X1 U8038 ( .A(n7069), .ZN(n6478) );
  OAI22_X1 U8039 ( .A1(n8141), .A2(n6478), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10250), .ZN(n6479) );
  OR4_X1 U8040 ( .A1(n6482), .A2(n6481), .A3(n6480), .A4(n6479), .ZN(P2_U3223)
         );
  INV_X1 U8041 ( .A(n7487), .ZN(n6483) );
  OR2_X1 U8042 ( .A1(n6483), .A2(n8872), .ZN(n6484) );
  NAND2_X1 U8043 ( .A1(n6637), .A2(n6484), .ZN(n9618) );
  OR2_X1 U8044 ( .A1(n9618), .A2(n6485), .ZN(n6486) );
  NAND2_X1 U8045 ( .A1(n6486), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  AND2_X1 U8046 ( .A1(n6492), .A2(P2_U3152), .ZN(n8604) );
  INV_X2 U8047 ( .A(n8604), .ZN(n8612) );
  OAI222_X1 U8048 ( .A1(n7729), .A2(n6487), .B1(n8612), .B2(n6498), .C1(
        P2_U3152), .C2(n9506), .ZN(P2_U3357) );
  OAI222_X1 U8049 ( .A1(n7729), .A2(n6489), .B1(n8612), .B2(n6493), .C1(
        P2_U3152), .C2(n6488), .ZN(P2_U3356) );
  OAI222_X1 U8050 ( .A1(n7729), .A2(n6491), .B1(n8612), .B2(n6496), .C1(
        P2_U3152), .C2(n6490), .ZN(P2_U3355) );
  NAND2_X1 U8051 ( .A1(n6492), .A2(P1_U3084), .ZN(n7622) );
  CLKBUF_X1 U8052 ( .A(n7622), .Z(n9499) );
  NOR2_X1 U8053 ( .A1(n6492), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9502) );
  OAI222_X1 U8054 ( .A1(n9499), .A2(n6494), .B1(n8036), .B2(n6493), .C1(
        P1_U3084), .C2(n9630), .ZN(P1_U3351) );
  OAI222_X1 U8055 ( .A1(n9499), .A2(n6497), .B1(n8036), .B2(n6496), .C1(
        P1_U3084), .C2(n6495), .ZN(P1_U3350) );
  OAI222_X1 U8056 ( .A1(n7622), .A2(n6499), .B1(n8036), .B2(n6498), .C1(
        P1_U3084), .C2(n6680), .ZN(P1_U3352) );
  INV_X1 U8057 ( .A(n6614), .ZN(n6500) );
  OAI222_X1 U8058 ( .A1(n7729), .A2(n5192), .B1(n8612), .B2(n6501), .C1(
        P2_U3152), .C2(n6500), .ZN(P2_U3354) );
  OAI222_X1 U8059 ( .A1(n9499), .A2(n6502), .B1(n8036), .B2(n6501), .C1(
        P1_U3084), .C2(n6710), .ZN(P1_U3349) );
  INV_X1 U8060 ( .A(n7729), .ZN(n6887) );
  AOI22_X1 U8061 ( .A1(n6630), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n6887), .ZN(n6503) );
  OAI21_X1 U8062 ( .B1(n6504), .B2(n8612), .A(n6503), .ZN(P2_U3353) );
  OAI222_X1 U8063 ( .A1(n9499), .A2(n6505), .B1(n8036), .B2(n6504), .C1(
        P1_U3084), .C2(n6727), .ZN(P1_U3348) );
  INV_X1 U8064 ( .A(n6506), .ZN(n6509) );
  AOI22_X1 U8065 ( .A1(n6665), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n6887), .ZN(n6507) );
  OAI21_X1 U8066 ( .B1(n6509), .B2(n8612), .A(n6507), .ZN(P2_U3352) );
  OAI222_X1 U8067 ( .A1(n9499), .A2(n10397), .B1(n8036), .B2(n6509), .C1(
        P1_U3084), .C2(n6508), .ZN(P1_U3347) );
  INV_X1 U8068 ( .A(n6510), .ZN(n6513) );
  AOI22_X1 U8069 ( .A1(n6795), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n6887), .ZN(n6511) );
  OAI21_X1 U8070 ( .B1(n6513), .B2(n8612), .A(n6511), .ZN(P2_U3351) );
  INV_X1 U8071 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10380) );
  INV_X1 U8072 ( .A(n6760), .ZN(n6512) );
  OAI222_X1 U8073 ( .A1(n9499), .A2(n10380), .B1(n8036), .B2(n6513), .C1(
        P1_U3084), .C2(n6512), .ZN(P1_U3346) );
  OAI21_X1 U8074 ( .B1(n9956), .B2(n6514), .A(n6556), .ZN(n6517) );
  NAND2_X1 U8075 ( .A1(n6515), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8033) );
  NAND2_X1 U8076 ( .A1(n9956), .A2(n8033), .ZN(n6516) );
  NAND2_X1 U8077 ( .A1(n6517), .A2(n6516), .ZN(n8242) );
  INV_X1 U8078 ( .A(n8242), .ZN(n9909) );
  NOR2_X1 U8079 ( .A1(n9909), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8080 ( .A(n6518), .ZN(n6527) );
  AOI22_X1 U8081 ( .A1(n6866), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n6887), .ZN(n6519) );
  OAI21_X1 U8082 ( .B1(n6527), .B2(n8612), .A(n6519), .ZN(P2_U3350) );
  INV_X1 U8083 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10261) );
  INV_X1 U8084 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6522) );
  NAND2_X1 U8085 ( .A1(n7823), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6521) );
  NAND2_X1 U8086 ( .A1(n5150), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6520) );
  OAI211_X1 U8087 ( .C1(n7827), .C2(n6522), .A(n6521), .B(n6520), .ZN(n7835)
         );
  NAND2_X1 U8088 ( .A1(P2_U3966), .A2(n7835), .ZN(n6523) );
  OAI21_X1 U8089 ( .B1(P2_U3966), .B2(n10261), .A(n6523), .ZN(P2_U3583) );
  INV_X1 U8090 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6526) );
  NAND2_X1 U8091 ( .A1(n9810), .A2(n7130), .ZN(n9808) );
  INV_X1 U8092 ( .A(n9808), .ZN(n6524) );
  OAI21_X1 U8093 ( .B1(n6524), .B2(P1_D_REG_0__SCAN_IN), .A(n7129), .ZN(n6525)
         );
  OAI21_X1 U8094 ( .B1(n6526), .B2(n9810), .A(n6525), .ZN(P1_U3440) );
  INV_X1 U8095 ( .A(n6892), .ZN(n6898) );
  OAI222_X1 U8096 ( .A1(n9499), .A2(n6528), .B1(n8036), .B2(n6527), .C1(
        P1_U3084), .C2(n6898), .ZN(P1_U3345) );
  INV_X1 U8097 ( .A(n6529), .ZN(n6534) );
  AOI22_X1 U8098 ( .A1(n6962), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n6887), .ZN(n6530) );
  OAI21_X1 U8099 ( .B1(n6534), .B2(n8612), .A(n6530), .ZN(P2_U3349) );
  INV_X1 U8100 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6532) );
  NAND2_X1 U8101 ( .A1(n8886), .A2(P1_U4006), .ZN(n6531) );
  OAI21_X1 U8102 ( .B1(P1_U4006), .B2(n6532), .A(n6531), .ZN(P1_U3555) );
  INV_X1 U8103 ( .A(n9672), .ZN(n6533) );
  OAI222_X1 U8104 ( .A1(n9499), .A2(n10192), .B1(n8036), .B2(n6534), .C1(n6533), .C2(P1_U3084), .ZN(P1_U3344) );
  INV_X1 U8105 ( .A(n6535), .ZN(n6542) );
  AOI22_X1 U8106 ( .A1(n7050), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n6887), .ZN(n6536) );
  OAI21_X1 U8107 ( .B1(n6542), .B2(n8612), .A(n6536), .ZN(P2_U3348) );
  INV_X1 U8108 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6541) );
  INV_X1 U8109 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9063) );
  NAND2_X1 U8110 ( .A1(n5915), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6539) );
  INV_X1 U8111 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9452) );
  OR2_X1 U8112 ( .A1(n6537), .A2(n9452), .ZN(n6538) );
  OAI211_X1 U8113 ( .C1(n4478), .C2(n9063), .A(n6539), .B(n6538), .ZN(n9066)
         );
  NAND2_X1 U8114 ( .A1(n9066), .A2(P1_U4006), .ZN(n6540) );
  OAI21_X1 U8115 ( .B1(P1_U4006), .B2(n6541), .A(n6540), .ZN(P1_U3586) );
  INV_X1 U8116 ( .A(n9689), .ZN(n6890) );
  OAI222_X1 U8117 ( .A1(n9499), .A2(n10463), .B1(n8036), .B2(n6542), .C1(n6890), .C2(P1_U3084), .ZN(P1_U3343) );
  MUX2_X1 U8118 ( .A(n6673), .B(n9597), .S(P1_U4006), .Z(n6543) );
  INV_X1 U8119 ( .A(n6543), .ZN(P1_U3567) );
  MUX2_X1 U8120 ( .A(n6544), .B(n9598), .S(P1_U4006), .Z(n6545) );
  INV_X1 U8121 ( .A(n6545), .ZN(P1_U3565) );
  MUX2_X1 U8122 ( .A(n6546), .B(n7348), .S(P1_U4006), .Z(n6547) );
  INV_X1 U8123 ( .A(n6547), .ZN(P1_U3563) );
  INV_X1 U8124 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6549) );
  INV_X1 U8125 ( .A(n6548), .ZN(n6550) );
  INV_X1 U8126 ( .A(n9694), .ZN(n6903) );
  OAI222_X1 U8127 ( .A1(n9499), .A2(n6549), .B1(n8036), .B2(n6550), .C1(n6903), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  INV_X1 U8128 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6551) );
  INV_X1 U8129 ( .A(n7242), .ZN(n7058) );
  OAI222_X1 U8130 ( .A1(n7729), .A2(n6551), .B1(n8612), .B2(n6550), .C1(n7058), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  OR2_X1 U8131 ( .A1(n9956), .A2(n6552), .ZN(n6553) );
  OAI211_X1 U8132 ( .C1(P2_U3152), .C2(n6554), .A(n6553), .B(n8033), .ZN(n6558) );
  NAND2_X1 U8133 ( .A1(n6558), .A2(n6556), .ZN(n6555) );
  NAND2_X1 U8134 ( .A1(n6555), .A2(n8166), .ZN(n6574) );
  INV_X1 U8135 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6568) );
  AND2_X1 U8136 ( .A1(n6556), .A2(n8243), .ZN(n6557) );
  INV_X1 U8137 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9912) );
  INV_X1 U8138 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10044) );
  INV_X1 U8139 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6559) );
  MUX2_X1 U8140 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6559), .S(n9506), .Z(n9514)
         );
  NOR3_X1 U8141 ( .A1(n9912), .A2(n10044), .A3(n9514), .ZN(n9512) );
  NOR2_X1 U8142 ( .A1(n9506), .A2(n6559), .ZN(n6560) );
  NOR2_X1 U8143 ( .A1(n9512), .A2(n6560), .ZN(n9530) );
  NAND2_X1 U8144 ( .A1(n9526), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6561) );
  OAI21_X1 U8145 ( .B1(n9526), .B2(P2_REG1_REG_2__SCAN_IN), .A(n6561), .ZN(
        n9529) );
  NOR2_X1 U8146 ( .A1(n9530), .A2(n9529), .ZN(n9528) );
  AOI21_X1 U8147 ( .B1(n9526), .B2(P2_REG1_REG_2__SCAN_IN), .A(n9528), .ZN(
        n6564) );
  OR2_X1 U8148 ( .A1(n6600), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6562) );
  NAND2_X1 U8149 ( .A1(n6600), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6591) );
  NAND2_X1 U8150 ( .A1(n6562), .A2(n6591), .ZN(n6563) );
  NOR2_X1 U8151 ( .A1(n6564), .A2(n6563), .ZN(n6589) );
  AOI21_X1 U8152 ( .B1(n6564), .B2(n6563), .A(n6589), .ZN(n6565) );
  NAND2_X1 U8153 ( .A1(n9904), .A2(n6565), .ZN(n6567) );
  INV_X1 U8154 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6808) );
  NOR2_X1 U8155 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6808), .ZN(n6807) );
  INV_X1 U8156 ( .A(n6807), .ZN(n6566) );
  OAI211_X1 U8157 ( .C1(n6568), .C2(n8242), .A(n6567), .B(n6566), .ZN(n6578)
         );
  NOR2_X1 U8158 ( .A1(n9506), .A2(n6569), .ZN(n6570) );
  NAND2_X1 U8159 ( .A1(n9526), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6571) );
  OAI21_X1 U8160 ( .B1(n9526), .B2(P2_REG2_REG_2__SCAN_IN), .A(n6571), .ZN(
        n9522) );
  NAND2_X1 U8161 ( .A1(n6600), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6572) );
  OAI21_X1 U8162 ( .B1(n6600), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6572), .ZN(
        n6575) );
  NOR2_X1 U8163 ( .A1(n5818), .A2(n8243), .ZN(n6573) );
  NAND2_X1 U8164 ( .A1(n6574), .A2(n6573), .ZN(n9907) );
  AOI211_X1 U8165 ( .C1(n6576), .C2(n6575), .A(n6599), .B(n9907), .ZN(n6577)
         );
  AOI211_X1 U8166 ( .C1(n9527), .C2(n6600), .A(n6578), .B(n6577), .ZN(n6579)
         );
  INV_X1 U8167 ( .A(n6579), .ZN(P2_U3248) );
  INV_X1 U8168 ( .A(n9794), .ZN(n8889) );
  OAI21_X1 U8169 ( .B1(n6582), .B2(n6581), .A(n6580), .ZN(n9635) );
  NAND2_X1 U8170 ( .A1(n9635), .A2(n8732), .ZN(n6587) );
  INV_X1 U8171 ( .A(n6583), .ZN(n6585) );
  NAND4_X1 U8172 ( .A1(n6585), .A2(n9810), .A3(n7489), .A4(n6584), .ZN(n8699)
         );
  AOI22_X1 U8173 ( .A1(n8699), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n8710), .B2(
        n9799), .ZN(n6586) );
  OAI211_X1 U8174 ( .C1(n8889), .C2(n8735), .A(n6587), .B(n6586), .ZN(P1_U3230) );
  INV_X1 U8175 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6598) );
  XNOR2_X1 U8176 ( .A(n6614), .B(n6588), .ZN(n6592) );
  INV_X1 U8177 ( .A(n6589), .ZN(n6590) );
  NAND2_X1 U8178 ( .A1(n6591), .A2(n6590), .ZN(n6593) );
  NAND2_X1 U8179 ( .A1(n6592), .A2(n6593), .ZN(n6608) );
  INV_X1 U8180 ( .A(n6592), .ZN(n6595) );
  INV_X1 U8181 ( .A(n6593), .ZN(n6594) );
  NAND2_X1 U8182 ( .A1(n6595), .A2(n6594), .ZN(n6596) );
  NAND3_X1 U8183 ( .A1(n9904), .A2(n6608), .A3(n6596), .ZN(n6597) );
  NAND2_X1 U8184 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n6818) );
  OAI211_X1 U8185 ( .C1(n6598), .C2(n8242), .A(n6597), .B(n6818), .ZN(n6604)
         );
  XNOR2_X1 U8186 ( .A(n6614), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n6601) );
  AOI211_X1 U8187 ( .C1(n6602), .C2(n6601), .A(n6613), .B(n9907), .ZN(n6603)
         );
  AOI211_X1 U8188 ( .C1(n9527), .C2(n6614), .A(n6604), .B(n6603), .ZN(n6605)
         );
  INV_X1 U8189 ( .A(n6605), .ZN(P2_U3249) );
  INV_X1 U8190 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6612) );
  OR2_X1 U8191 ( .A1(n6630), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6606) );
  NAND2_X1 U8192 ( .A1(n6630), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6621) );
  AND2_X1 U8193 ( .A1(n6606), .A2(n6621), .ZN(n6610) );
  NAND2_X1 U8194 ( .A1(n6614), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6607) );
  NAND2_X1 U8195 ( .A1(n6608), .A2(n6607), .ZN(n6609) );
  NAND2_X1 U8196 ( .A1(n6609), .A2(n6610), .ZN(n6622) );
  OAI211_X1 U8197 ( .C1(n6610), .C2(n6609), .A(n9904), .B(n6622), .ZN(n6611)
         );
  NAND2_X1 U8198 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3152), .ZN(n6826) );
  OAI211_X1 U8199 ( .C1(n6612), .C2(n8242), .A(n6611), .B(n6826), .ZN(n6619)
         );
  NAND2_X1 U8200 ( .A1(n6630), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6615) );
  OAI21_X1 U8201 ( .B1(n6630), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6615), .ZN(
        n6616) );
  AOI211_X1 U8202 ( .C1(n6617), .C2(n6616), .A(n6629), .B(n9907), .ZN(n6618)
         );
  AOI211_X1 U8203 ( .C1(n9527), .C2(n6630), .A(n6619), .B(n6618), .ZN(n6620)
         );
  INV_X1 U8204 ( .A(n6620), .ZN(P2_U3250) );
  INV_X1 U8205 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10510) );
  AND2_X1 U8206 ( .A1(n6622), .A2(n6621), .ZN(n6626) );
  OR2_X1 U8207 ( .A1(n6665), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6624) );
  NAND2_X1 U8208 ( .A1(n6665), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6623) );
  NAND2_X1 U8209 ( .A1(n6624), .A2(n6623), .ZN(n6625) );
  NOR2_X1 U8210 ( .A1(n6626), .A2(n6625), .ZN(n6658) );
  AOI21_X1 U8211 ( .B1(n6626), .B2(n6625), .A(n6658), .ZN(n6627) );
  NAND2_X1 U8212 ( .A1(n9904), .A2(n6627), .ZN(n6628) );
  NAND2_X1 U8213 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n6835) );
  OAI211_X1 U8214 ( .C1(n10510), .C2(n8242), .A(n6628), .B(n6835), .ZN(n6635)
         );
  NAND2_X1 U8215 ( .A1(n6665), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6631) );
  OAI21_X1 U8216 ( .B1(n6665), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6631), .ZN(
        n6632) );
  NOR2_X1 U8217 ( .A1(n6633), .A2(n6632), .ZN(n6664) );
  AOI211_X1 U8218 ( .C1(n6633), .C2(n6632), .A(n6664), .B(n9907), .ZN(n6634)
         );
  AOI211_X1 U8219 ( .C1(n9527), .C2(n6665), .A(n6635), .B(n6634), .ZN(n6636)
         );
  INV_X1 U8220 ( .A(n6636), .ZN(P2_U3251) );
  INV_X1 U8221 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6655) );
  INV_X1 U8222 ( .A(n6637), .ZN(n6638) );
  NOR2_X2 U8223 ( .A1(P1_U3083), .A2(n6638), .ZN(n9690) );
  INV_X1 U8224 ( .A(n9690), .ZN(n9724) );
  OR2_X1 U8225 ( .A1(n9613), .A2(P1_U3084), .ZN(n7647) );
  NOR2_X1 U8226 ( .A1(n9618), .A2(n7647), .ZN(n7747) );
  NAND2_X1 U8227 ( .A1(n7747), .A2(n4480), .ZN(n9715) );
  INV_X1 U8228 ( .A(n9715), .ZN(n9695) );
  AND2_X1 U8229 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6853) );
  INV_X1 U8230 ( .A(n6680), .ZN(n6640) );
  INV_X1 U8231 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9890) );
  MUX2_X1 U8232 ( .A(n9890), .B(P1_REG1_REG_1__SCAN_IN), .S(n6680), .Z(n6678)
         );
  NAND3_X1 U8233 ( .A1(n6678), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_REG1_REG_0__SCAN_IN), .ZN(n6676) );
  INV_X1 U8234 ( .A(n6676), .ZN(n6639) );
  AOI21_X1 U8235 ( .B1(n6640), .B2(P1_REG1_REG_1__SCAN_IN), .A(n6639), .ZN(
        n9626) );
  XNOR2_X1 U8236 ( .A(n6646), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9625) );
  NOR2_X1 U8237 ( .A1(n9626), .A2(n9625), .ZN(n9624) );
  AOI21_X1 U8238 ( .B1(P1_REG1_REG_2__SCAN_IN), .B2(n6646), .A(n9624), .ZN(
        n6644) );
  NAND2_X1 U8239 ( .A1(n6718), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6641) );
  OAI21_X1 U8240 ( .B1(n6718), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6641), .ZN(
        n6643) );
  NOR2_X1 U8241 ( .A1(n6644), .A2(n6643), .ZN(n6717) );
  INV_X1 U8242 ( .A(n9613), .ZN(n9064) );
  OR2_X1 U8243 ( .A1(n4480), .A2(n9064), .ZN(n9634) );
  INV_X1 U8244 ( .A(n9634), .ZN(n9638) );
  NAND2_X1 U8245 ( .A1(n9638), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6642) );
  OR2_X1 U8246 ( .A1(n6642), .A2(n9618), .ZN(n9623) );
  AOI211_X1 U8247 ( .C1(n6644), .C2(n6643), .A(n6717), .B(n9623), .ZN(n6645)
         );
  AOI211_X1 U8248 ( .C1(n9695), .C2(n6718), .A(n6853), .B(n6645), .ZN(n6654)
         );
  NAND2_X1 U8249 ( .A1(n6646), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6648) );
  AOI22_X1 U8250 ( .A1(n6646), .A2(P1_REG2_REG_2__SCAN_IN), .B1(n7168), .B2(
        n9630), .ZN(n9629) );
  NAND3_X1 U8251 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .A3(n6682), .ZN(n6681) );
  OAI21_X1 U8252 ( .B1(n6647), .B2(n6680), .A(n6681), .ZN(n9628) );
  NAND2_X1 U8253 ( .A1(n9629), .A2(n9628), .ZN(n9627) );
  NAND2_X1 U8254 ( .A1(n6648), .A2(n9627), .ZN(n6652) );
  MUX2_X1 U8255 ( .A(n5954), .B(P1_REG2_REG_3__SCAN_IN), .S(n6718), .Z(n6649)
         );
  INV_X1 U8256 ( .A(n6649), .ZN(n6651) );
  INV_X1 U8257 ( .A(n7747), .ZN(n6650) );
  NOR2_X1 U8258 ( .A1(n6650), .A2(n4480), .ZN(n9711) );
  OAI211_X1 U8259 ( .C1(n6652), .C2(n6651), .A(n9711), .B(n6708), .ZN(n6653)
         );
  OAI211_X1 U8260 ( .C1(n6655), .C2(n9724), .A(n6654), .B(n6653), .ZN(P1_U3244) );
  INV_X1 U8261 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10497) );
  OR2_X1 U8262 ( .A1(n6795), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6657) );
  NAND2_X1 U8263 ( .A1(n6795), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6656) );
  NAND2_X1 U8264 ( .A1(n6657), .A2(n6656), .ZN(n6660) );
  AOI21_X1 U8265 ( .B1(n6665), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6658), .ZN(
        n6659) );
  NOR2_X1 U8266 ( .A1(n6659), .A2(n6660), .ZN(n6786) );
  AOI21_X1 U8267 ( .B1(n6660), .B2(n6659), .A(n6786), .ZN(n6661) );
  NAND2_X1 U8268 ( .A1(n9904), .A2(n6661), .ZN(n6663) );
  NOR2_X1 U8269 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5278), .ZN(n6880) );
  INV_X1 U8270 ( .A(n6880), .ZN(n6662) );
  OAI211_X1 U8271 ( .C1(n10497), .C2(n8242), .A(n6663), .B(n6662), .ZN(n6670)
         );
  NAND2_X1 U8272 ( .A1(n6795), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6666) );
  OAI21_X1 U8273 ( .B1(n6795), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6666), .ZN(
        n6667) );
  NOR2_X1 U8274 ( .A1(n6668), .A2(n6667), .ZN(n6794) );
  AOI211_X1 U8275 ( .C1(n6668), .C2(n6667), .A(n6794), .B(n9907), .ZN(n6669)
         );
  AOI211_X1 U8276 ( .C1(n9527), .C2(n6795), .A(n6670), .B(n6669), .ZN(n6671)
         );
  INV_X1 U8277 ( .A(n6671), .ZN(P2_U3252) );
  INV_X1 U8278 ( .A(n6672), .ZN(n6674) );
  INV_X1 U8279 ( .A(n7283), .ZN(n7290) );
  OAI222_X1 U8280 ( .A1(n7729), .A2(n6673), .B1(n8612), .B2(n6674), .C1(
        P2_U3152), .C2(n7290), .ZN(P2_U3346) );
  INV_X1 U8281 ( .A(n7018), .ZN(n6910) );
  OAI222_X1 U8282 ( .A1(n7622), .A2(n6675), .B1(n8036), .B2(n6674), .C1(
        P1_U3084), .C2(n6910), .ZN(P1_U3341) );
  AND2_X1 U8283 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6677) );
  INV_X1 U8284 ( .A(n9623), .ZN(n9720) );
  OAI211_X1 U8285 ( .C1(n6678), .C2(n6677), .A(n9720), .B(n6676), .ZN(n6679)
         );
  OAI21_X1 U8286 ( .B1(n9715), .B2(n6680), .A(n6679), .ZN(n6686) );
  AND2_X1 U8287 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6683) );
  OAI211_X1 U8288 ( .C1(n6683), .C2(n6682), .A(n9711), .B(n6681), .ZN(n6684)
         );
  OAI21_X1 U8289 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n7144), .A(n6684), .ZN(n6685) );
  AOI211_X1 U8290 ( .C1(n9690), .C2(P1_ADDR_REG_1__SCAN_IN), .A(n6686), .B(
        n6685), .ZN(n6687) );
  INV_X1 U8291 ( .A(n6687), .ZN(P1_U3242) );
  NOR2_X1 U8292 ( .A1(n9956), .A2(n6688), .ZN(n6689) );
  NAND2_X1 U8293 ( .A1(n6690), .A2(n6689), .ZN(n6923) );
  INV_X2 U8294 ( .A(n10042), .ZN(n10043) );
  NAND2_X1 U8295 ( .A1(n7804), .A2(n7716), .ZN(n6695) );
  INV_X1 U8296 ( .A(n7716), .ZN(n6933) );
  NAND2_X1 U8297 ( .A1(n4941), .A2(n6933), .ZN(n7853) );
  AND2_X1 U8298 ( .A1(n6695), .A2(n7853), .ZN(n7994) );
  XOR2_X1 U8299 ( .A(n6934), .B(n7994), .Z(n6988) );
  INV_X1 U8300 ( .A(n6988), .ZN(n6703) );
  XNOR2_X1 U8301 ( .A(n6946), .B(n5827), .ZN(n6693) );
  OR2_X1 U8302 ( .A1(n6693), .A2(n8356), .ZN(n7064) );
  INV_X1 U8303 ( .A(n10020), .ZN(n6694) );
  NAND2_X1 U8304 ( .A1(n7064), .A2(n6694), .ZN(n10041) );
  INV_X1 U8305 ( .A(n10041), .ZN(n9995) );
  NAND2_X1 U8306 ( .A1(n7720), .A2(n9963), .ZN(n6983) );
  INV_X1 U8307 ( .A(n7853), .ZN(n6696) );
  OR2_X1 U8308 ( .A1(n7855), .A2(n6696), .ZN(n6698) );
  NAND2_X1 U8309 ( .A1(n8022), .A2(n8023), .ZN(n7838) );
  INV_X1 U8310 ( .A(n7838), .ZN(n6697) );
  OAI211_X1 U8311 ( .C1(n7994), .C2(n6983), .A(n6698), .B(n9938), .ZN(n6701)
         );
  OAI22_X1 U8312 ( .A1(n7720), .A2(n8426), .B1(n6937), .B2(n8428), .ZN(n6699)
         );
  INV_X1 U8313 ( .A(n6699), .ZN(n6700) );
  AND2_X1 U8314 ( .A1(n6701), .A2(n6700), .ZN(n6993) );
  XNOR2_X1 U8315 ( .A(n6779), .B(n7716), .ZN(n6990) );
  OR2_X1 U8316 ( .A1(n7991), .A2(n8022), .ZN(n10036) );
  INV_X1 U8317 ( .A(n10036), .ZN(n10003) );
  AOI22_X1 U8318 ( .A1(n6990), .A2(n10003), .B1(n10002), .B2(n7716), .ZN(n6702) );
  OAI211_X1 U8319 ( .C1(n6703), .C2(n9995), .A(n6993), .B(n6702), .ZN(n6706)
         );
  NAND2_X1 U8320 ( .A1(n6706), .A2(n10043), .ZN(n6704) );
  OAI21_X1 U8321 ( .B1(n10043), .B2(n5097), .A(n6704), .ZN(P2_U3454) );
  INV_X2 U8322 ( .A(n10062), .ZN(n10064) );
  NAND2_X1 U8323 ( .A1(n6706), .A2(n10064), .ZN(n6707) );
  OAI21_X1 U8324 ( .B1(n10064), .B2(n6559), .A(n6707), .ZN(P2_U3521) );
  INV_X1 U8325 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6715) );
  NOR2_X1 U8326 ( .A1(n9645), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6711) );
  NAND2_X1 U8327 ( .A1(n6718), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6709) );
  AOI22_X1 U8328 ( .A1(n9645), .A2(n5968), .B1(P1_REG2_REG_4__SCAN_IN), .B2(
        n6710), .ZN(n9647) );
  AOI22_X1 U8329 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6727), .B1(n6741), .B2(
        n5992), .ZN(n6712) );
  NOR2_X1 U8330 ( .A1(n6713), .A2(n6712), .ZN(n6742) );
  AOI21_X1 U8331 ( .B1(n6713), .B2(n6712), .A(n6742), .ZN(n6714) );
  INV_X1 U8332 ( .A(n9711), .ZN(n9682) );
  OAI22_X1 U8333 ( .A1(n9724), .A2(n6715), .B1(n6714), .B2(n9682), .ZN(n6729)
         );
  NAND2_X1 U8334 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7096) );
  NOR2_X1 U8335 ( .A1(n9645), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6716) );
  AOI21_X1 U8336 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9645), .A(n6716), .ZN(
        n9643) );
  AOI21_X1 U8337 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n6718), .A(n6717), .ZN(
        n9642) );
  NAND2_X1 U8338 ( .A1(n9643), .A2(n9642), .ZN(n9641) );
  OR2_X1 U8339 ( .A1(n9645), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6719) );
  NAND2_X1 U8340 ( .A1(n9641), .A2(n6719), .ZN(n6722) );
  OR2_X1 U8341 ( .A1(n6741), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6721) );
  NAND2_X1 U8342 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6741), .ZN(n6720) );
  NAND2_X1 U8343 ( .A1(n6721), .A2(n6720), .ZN(n6723) );
  NAND2_X1 U8344 ( .A1(n6722), .A2(n6723), .ZN(n6725) );
  NOR2_X1 U8345 ( .A1(n6723), .A2(n6722), .ZN(n6732) );
  INV_X1 U8346 ( .A(n6732), .ZN(n6724) );
  NAND3_X1 U8347 ( .A1(n9720), .A2(n6725), .A3(n6724), .ZN(n6726) );
  OAI211_X1 U8348 ( .C1(n9715), .C2(n6727), .A(n7096), .B(n6726), .ZN(n6728)
         );
  OR2_X1 U8349 ( .A1(n6729), .A2(n6728), .ZN(P1_U3246) );
  NAND2_X1 U8350 ( .A1(n6892), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6730) );
  OAI21_X1 U8351 ( .B1(n6892), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6730), .ZN(
        n6736) );
  OR2_X1 U8352 ( .A1(n6760), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6734) );
  NOR2_X1 U8353 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6760), .ZN(n6731) );
  AOI21_X1 U8354 ( .B1(n6760), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6731), .ZN(
        n6755) );
  AOI21_X1 U8355 ( .B1(n6741), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6732), .ZN(
        n9657) );
  NOR2_X1 U8356 ( .A1(n9654), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6733) );
  AOI21_X1 U8357 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n9654), .A(n6733), .ZN(
        n9658) );
  NAND2_X1 U8358 ( .A1(n9657), .A2(n9658), .ZN(n9656) );
  OAI21_X1 U8359 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n9654), .A(n9656), .ZN(
        n6756) );
  NAND2_X1 U8360 ( .A1(n6755), .A2(n6756), .ZN(n6754) );
  NAND2_X1 U8361 ( .A1(n6734), .A2(n6754), .ZN(n6735) );
  NOR2_X1 U8362 ( .A1(n6736), .A2(n6735), .ZN(n6891) );
  AOI21_X1 U8363 ( .B1(n6736), .B2(n6735), .A(n6891), .ZN(n6738) );
  INV_X1 U8364 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6737) );
  NOR2_X1 U8365 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6737), .ZN(n7216) );
  AOI21_X1 U8366 ( .B1(n9720), .B2(n6738), .A(n7216), .ZN(n6739) );
  OAI21_X1 U8367 ( .B1(n9715), .B2(n6898), .A(n6739), .ZN(n6752) );
  INV_X1 U8368 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6740) );
  MUX2_X1 U8369 ( .A(n6740), .B(P1_REG2_REG_7__SCAN_IN), .S(n6760), .Z(n6758)
         );
  NAND2_X1 U8370 ( .A1(n9654), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6745) );
  NOR2_X1 U8371 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6741), .ZN(n6743) );
  NOR2_X1 U8372 ( .A1(n6743), .A2(n6742), .ZN(n9662) );
  MUX2_X1 U8373 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6744), .S(n9654), .Z(n9661)
         );
  NAND2_X1 U8374 ( .A1(n9662), .A2(n9661), .ZN(n9660) );
  NAND2_X1 U8375 ( .A1(n6745), .A2(n9660), .ZN(n6759) );
  NOR2_X1 U8376 ( .A1(n6898), .A2(n6746), .ZN(n6899) );
  XNOR2_X1 U8377 ( .A(n4559), .B(n6746), .ZN(n6748) );
  NOR2_X1 U8378 ( .A1(n4559), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6747) );
  MUX2_X1 U8379 ( .A(n6748), .B(n6747), .S(n6892), .Z(n6749) );
  AOI21_X1 U8380 ( .B1(n4559), .B2(n6899), .A(n6749), .ZN(n6750) );
  NOR2_X1 U8381 ( .A1(n6750), .A2(n9682), .ZN(n6751) );
  AOI211_X1 U8382 ( .C1(n9690), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n6752), .B(
        n6751), .ZN(n6753) );
  INV_X1 U8383 ( .A(n6753), .ZN(P1_U3249) );
  OAI21_X1 U8384 ( .B1(n6756), .B2(n6755), .A(n6754), .ZN(n6765) );
  AOI21_X1 U8385 ( .B1(n6759), .B2(n6758), .A(n6757), .ZN(n6763) );
  AND2_X1 U8386 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7041) );
  AOI21_X1 U8387 ( .B1(n9695), .B2(n6760), .A(n7041), .ZN(n6762) );
  NAND2_X1 U8388 ( .A1(n9690), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n6761) );
  OAI211_X1 U8389 ( .C1(n6763), .C2(n9682), .A(n6762), .B(n6761), .ZN(n6764)
         );
  AOI21_X1 U8390 ( .B1(n9720), .B2(n6765), .A(n6764), .ZN(n6766) );
  INV_X1 U8391 ( .A(n6766), .ZN(P1_U3248) );
  NAND2_X1 U8392 ( .A1(n6767), .A2(n6768), .ZN(n6770) );
  XNOR2_X1 U8393 ( .A(n6770), .B(n6769), .ZN(n6773) );
  AOI22_X1 U8394 ( .A1(n8699), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n8710), .B2(
        n8888), .ZN(n6772) );
  INV_X1 U8395 ( .A(n8723), .ZN(n8740) );
  AOI22_X1 U8396 ( .A1(n8740), .A2(n8886), .B1(n8725), .B2(n7151), .ZN(n6771)
         );
  OAI211_X1 U8397 ( .C1(n6773), .C2(n8712), .A(n6772), .B(n6771), .ZN(P1_U3220) );
  INV_X1 U8398 ( .A(n6774), .ZN(n6776) );
  INV_X1 U8399 ( .A(n7458), .ZN(n7288) );
  OAI222_X1 U8400 ( .A1(n7729), .A2(n6775), .B1(n8612), .B2(n6776), .C1(n7288), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8401 ( .A(n7228), .ZN(n7031) );
  OAI222_X1 U8402 ( .A1(n7622), .A2(n6777), .B1(n8036), .B2(n6776), .C1(n7031), 
        .C2(P1_U3084), .ZN(P1_U3340) );
  OR2_X1 U8403 ( .A1(n6778), .A2(P2_U3152), .ZN(n7809) );
  INV_X1 U8404 ( .A(n7809), .ZN(n6785) );
  AOI22_X1 U8405 ( .A1(n7717), .A2(n4941), .B1(n8143), .B2(n9963), .ZN(n6784)
         );
  INV_X1 U8406 ( .A(n6983), .ZN(n6782) );
  INV_X1 U8407 ( .A(n7720), .ZN(n8167) );
  NAND2_X1 U8408 ( .A1(n8167), .A2(n6779), .ZN(n7867) );
  INV_X1 U8409 ( .A(n7867), .ZN(n6780) );
  MUX2_X1 U8410 ( .A(n9963), .B(n6780), .S(n7839), .Z(n6781) );
  INV_X1 U8411 ( .A(n8145), .ZN(n8117) );
  OAI21_X1 U8412 ( .B1(n6782), .B2(n6781), .A(n8117), .ZN(n6783) );
  OAI211_X1 U8413 ( .C1(n6785), .C2(n6984), .A(n6784), .B(n6783), .ZN(P2_U3234) );
  INV_X1 U8414 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10508) );
  AOI21_X1 U8415 ( .B1(n6795), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6786), .ZN(
        n6790) );
  INV_X1 U8416 ( .A(n6790), .ZN(n6788) );
  XNOR2_X1 U8417 ( .A(n6866), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n6789) );
  INV_X1 U8418 ( .A(n6789), .ZN(n6787) );
  NAND2_X1 U8419 ( .A1(n6788), .A2(n6787), .ZN(n6860) );
  NAND2_X1 U8420 ( .A1(n6790), .A2(n6789), .ZN(n6791) );
  NAND3_X1 U8421 ( .A1(n9904), .A2(n6860), .A3(n6791), .ZN(n6793) );
  NAND2_X1 U8422 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n6792) );
  OAI211_X1 U8423 ( .C1(n10508), .C2(n8242), .A(n6793), .B(n6792), .ZN(n6799)
         );
  AOI21_X1 U8424 ( .B1(n6795), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6794), .ZN(
        n6797) );
  XNOR2_X1 U8425 ( .A(n6866), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n6796) );
  NOR2_X1 U8426 ( .A1(n6797), .A2(n6796), .ZN(n6865) );
  AOI211_X1 U8427 ( .C1(n6797), .C2(n6796), .A(n6865), .B(n9907), .ZN(n6798)
         );
  AOI211_X1 U8428 ( .C1(n9527), .C2(n6866), .A(n6799), .B(n6798), .ZN(n6800)
         );
  INV_X1 U8429 ( .A(n6800), .ZN(P2_U3253) );
  INV_X1 U8430 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6802) );
  INV_X1 U8431 ( .A(n6801), .ZN(n6803) );
  INV_X1 U8432 ( .A(n8174), .ZN(n7464) );
  OAI222_X1 U8433 ( .A1(n7729), .A2(n6802), .B1(n8612), .B2(n6803), .C1(n7464), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8434 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10252) );
  INV_X1 U8435 ( .A(n7507), .ZN(n7513) );
  OAI222_X1 U8436 ( .A1(n7622), .A2(n10252), .B1(n8036), .B2(n6803), .C1(n7513), .C2(P1_U3084), .ZN(P1_U3339) );
  INV_X1 U8437 ( .A(n8128), .ZN(n8138) );
  OR2_X1 U8438 ( .A1(n6937), .A2(n8426), .ZN(n6805) );
  INV_X1 U8439 ( .A(n8428), .ZN(n9917) );
  NAND2_X1 U8440 ( .A1(n8164), .A2(n9917), .ZN(n6804) );
  AND2_X1 U8441 ( .A1(n6805), .A2(n6804), .ZN(n6997) );
  NOR2_X1 U8442 ( .A1(n8141), .A2(n6997), .ZN(n6806) );
  AOI211_X1 U8443 ( .C1(n8138), .C2(n6808), .A(n6807), .B(n6806), .ZN(n6813)
         );
  XOR2_X1 U8444 ( .A(n6810), .B(n6809), .Z(n6811) );
  NAND2_X1 U8445 ( .A1(n6811), .A2(n8117), .ZN(n6812) );
  OAI211_X1 U8446 ( .C1(n4879), .C2(n8123), .A(n6813), .B(n6812), .ZN(P2_U3220) );
  INV_X1 U8447 ( .A(n6814), .ZN(n6815) );
  AOI21_X1 U8448 ( .B1(n6817), .B2(n6816), .A(n6815), .ZN(n6822) );
  INV_X1 U8449 ( .A(n8129), .ZN(n6881) );
  INV_X1 U8450 ( .A(n7803), .ZN(n9916) );
  OAI21_X1 U8451 ( .B1(n8128), .B2(n9925), .A(n6818), .ZN(n6820) );
  INV_X1 U8452 ( .A(n9918), .ZN(n6944) );
  OAI22_X1 U8453 ( .A1(n8131), .A2(n6944), .B1(n9981), .B2(n8123), .ZN(n6819)
         );
  AOI211_X1 U8454 ( .C1(n6881), .C2(n9916), .A(n6820), .B(n6819), .ZN(n6821)
         );
  OAI21_X1 U8455 ( .B1(n6822), .B2(n8145), .A(n6821), .ZN(P2_U3232) );
  OAI21_X1 U8456 ( .B1(n6825), .B2(n6824), .A(n6823), .ZN(n6830) );
  NAND2_X1 U8457 ( .A1(n6881), .A2(n8164), .ZN(n6827) );
  OAI211_X1 U8458 ( .C1(n8128), .C2(n7010), .A(n6827), .B(n6826), .ZN(n6829)
         );
  INV_X1 U8459 ( .A(n8163), .ZN(n7883) );
  OAI22_X1 U8460 ( .A1(n8131), .A2(n7883), .B1(n9989), .B2(n8123), .ZN(n6828)
         );
  AOI211_X1 U8461 ( .C1(n8117), .C2(n6830), .A(n6829), .B(n6828), .ZN(n6831)
         );
  INV_X1 U8462 ( .A(n6831), .ZN(P2_U3229) );
  OAI21_X1 U8463 ( .B1(n6834), .B2(n6833), .A(n6832), .ZN(n6839) );
  INV_X1 U8464 ( .A(n7884), .ZN(n9992) );
  OAI22_X1 U8465 ( .A1(n8131), .A2(n7062), .B1(n9992), .B2(n8123), .ZN(n6838)
         );
  NAND2_X1 U8466 ( .A1(n6881), .A2(n9918), .ZN(n6836) );
  OAI211_X1 U8467 ( .C1(n8128), .C2(n6975), .A(n6836), .B(n6835), .ZN(n6837)
         );
  AOI211_X1 U8468 ( .C1(n6839), .C2(n8117), .A(n6838), .B(n6837), .ZN(n6840)
         );
  INV_X1 U8469 ( .A(n6840), .ZN(P2_U3241) );
  NAND2_X1 U8470 ( .A1(n6841), .A2(n8732), .ZN(n6848) );
  AOI21_X1 U8471 ( .B1(n6851), .B2(n6843), .A(n6842), .ZN(n6847) );
  AOI22_X1 U8472 ( .A1(n8740), .A2(n9773), .B1(n8725), .B2(n9844), .ZN(n6846)
         );
  AND2_X1 U8473 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9650) );
  INV_X1 U8474 ( .A(n8721), .ZN(n8736) );
  NOR2_X1 U8475 ( .A1(n8736), .A2(n9777), .ZN(n6844) );
  AOI211_X1 U8476 ( .C1(n7321), .C2(n8710), .A(n9650), .B(n6844), .ZN(n6845)
         );
  OAI211_X1 U8477 ( .C1(n6848), .C2(n6847), .A(n6846), .B(n6845), .ZN(P1_U3228) );
  INV_X1 U8478 ( .A(n6849), .ZN(n6885) );
  AOI22_X1 U8479 ( .A1(n8203), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n6887), .ZN(n6850) );
  OAI21_X1 U8480 ( .B1(n6885), .B2(n8612), .A(n6850), .ZN(P2_U3342) );
  AOI22_X1 U8481 ( .A1(n8740), .A2(n7151), .B1(n8725), .B2(n9035), .ZN(n6855)
         );
  AOI21_X1 U8482 ( .B1(n8710), .B2(n7251), .A(n6853), .ZN(n6854) );
  OAI211_X1 U8483 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n8736), .A(n6855), .B(
        n6854), .ZN(n6856) );
  AOI21_X1 U8484 ( .B1(n6857), .B2(n8732), .A(n6856), .ZN(n6858) );
  INV_X1 U8485 ( .A(n6858), .ZN(P1_U3216) );
  INV_X1 U8486 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n6864) );
  INV_X1 U8487 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10058) );
  MUX2_X1 U8488 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10058), .S(n6962), .Z(n6862)
         );
  NAND2_X1 U8489 ( .A1(n6866), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6859) );
  NAND2_X1 U8490 ( .A1(n6860), .A2(n6859), .ZN(n6861) );
  NAND2_X1 U8491 ( .A1(n6861), .A2(n6862), .ZN(n6952) );
  OAI211_X1 U8492 ( .C1(n6862), .C2(n6861), .A(n9904), .B(n6952), .ZN(n6863)
         );
  NAND2_X1 U8493 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7085) );
  OAI211_X1 U8494 ( .C1(n6864), .C2(n8242), .A(n6863), .B(n7085), .ZN(n6872)
         );
  OR2_X1 U8495 ( .A1(n6962), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6868) );
  NAND2_X1 U8496 ( .A1(n6962), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6867) );
  NAND2_X1 U8497 ( .A1(n6868), .A2(n6867), .ZN(n6869) );
  AOI211_X1 U8498 ( .C1(n6870), .C2(n6869), .A(n6961), .B(n9907), .ZN(n6871)
         );
  AOI211_X1 U8499 ( .C1(n9527), .C2(n6962), .A(n6872), .B(n6871), .ZN(n6873)
         );
  INV_X1 U8500 ( .A(n6873), .ZN(P2_U3254) );
  INV_X1 U8501 ( .A(n6874), .ZN(n6876) );
  OAI222_X1 U8502 ( .A1(n7729), .A2(n6875), .B1(n8612), .B2(n6876), .C1(
        P2_U3152), .C2(n8187), .ZN(P2_U3343) );
  OAI222_X1 U8503 ( .A1(n7622), .A2(n10454), .B1(n8036), .B2(n6876), .C1(
        P1_U3084), .C2(n7739), .ZN(P1_U3338) );
  XNOR2_X1 U8504 ( .A(n6878), .B(n6877), .ZN(n6884) );
  INV_X1 U8505 ( .A(n7177), .ZN(n8161) );
  AOI22_X1 U8506 ( .A1(n7717), .A2(n8161), .B1(n8143), .B2(n10001), .ZN(n6883)
         );
  NOR2_X1 U8507 ( .A1(n8128), .A2(n6928), .ZN(n6879) );
  AOI211_X1 U8508 ( .C1(n6881), .C2(n8163), .A(n6880), .B(n6879), .ZN(n6882)
         );
  OAI211_X1 U8509 ( .C1(n6884), .C2(n8145), .A(n6883), .B(n6882), .ZN(P2_U3215) );
  INV_X1 U8510 ( .A(n7742), .ZN(n9046) );
  OAI222_X1 U8511 ( .A1(n7622), .A2(n10194), .B1(n8036), .B2(n6885), .C1(n9046), .C2(P1_U3084), .ZN(P1_U3337) );
  INV_X1 U8512 ( .A(n6886), .ZN(n6950) );
  AOI22_X1 U8513 ( .A1(n8218), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n6887), .ZN(n6888) );
  OAI21_X1 U8514 ( .B1(n6950), .B2(n8612), .A(n6888), .ZN(P2_U3341) );
  MUX2_X1 U8515 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6889), .S(n7018), .Z(n6896)
         );
  AOI22_X1 U8516 ( .A1(n9689), .A2(P1_REG1_REG_10__SCAN_IN), .B1(n6111), .B2(
        n6890), .ZN(n9681) );
  AOI21_X1 U8517 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n6892), .A(n6891), .ZN(
        n9674) );
  NOR2_X1 U8518 ( .A1(n9672), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6893) );
  AOI21_X1 U8519 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9672), .A(n6893), .ZN(
        n9675) );
  NAND2_X1 U8520 ( .A1(n9674), .A2(n9675), .ZN(n9673) );
  OAI21_X1 U8521 ( .B1(n9672), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9673), .ZN(
        n9680) );
  NAND2_X1 U8522 ( .A1(n9681), .A2(n9680), .ZN(n9679) );
  OAI21_X1 U8523 ( .B1(n9689), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9679), .ZN(
        n9698) );
  MUX2_X1 U8524 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n6894), .S(n9694), .Z(n9697)
         );
  NAND2_X1 U8525 ( .A1(n9698), .A2(n9697), .ZN(n9696) );
  OAI21_X1 U8526 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9694), .A(n9696), .ZN(
        n6895) );
  NAND2_X1 U8527 ( .A1(n6895), .A2(n6896), .ZN(n7017) );
  OAI21_X1 U8528 ( .B1(n6896), .B2(n6895), .A(n7017), .ZN(n6897) );
  NAND2_X1 U8529 ( .A1(n6897), .A2(n9720), .ZN(n6913) );
  MUX2_X1 U8530 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n7474), .S(n9694), .Z(n9700)
         );
  NAND2_X1 U8531 ( .A1(n6898), .A2(n6746), .ZN(n6900) );
  NAND2_X1 U8532 ( .A1(n9672), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6901) );
  OAI21_X1 U8533 ( .B1(n9672), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6901), .ZN(
        n9668) );
  AOI21_X1 U8534 ( .B1(n9672), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9667), .ZN(
        n9685) );
  NAND2_X1 U8535 ( .A1(n9689), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6902) );
  OAI21_X1 U8536 ( .B1(n9689), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6902), .ZN(
        n9684) );
  NOR2_X1 U8537 ( .A1(n9685), .A2(n9684), .ZN(n9683) );
  AOI21_X1 U8538 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9689), .A(n9683), .ZN(
        n9701) );
  NAND2_X1 U8539 ( .A1(n9700), .A2(n9701), .ZN(n9699) );
  NAND2_X1 U8540 ( .A1(n6903), .A2(n7474), .ZN(n6904) );
  NAND2_X1 U8541 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7018), .ZN(n7023) );
  OAI21_X1 U8542 ( .B1(n7018), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7023), .ZN(
        n6905) );
  INV_X1 U8543 ( .A(n6905), .ZN(n6906) );
  NAND2_X1 U8544 ( .A1(n6907), .A2(n6906), .ZN(n7024) );
  OAI211_X1 U8545 ( .C1(n6907), .C2(n6906), .A(n9711), .B(n7024), .ZN(n6909)
         );
  NAND2_X1 U8546 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n6908) );
  OAI211_X1 U8547 ( .C1(n9715), .C2(n6910), .A(n6909), .B(n6908), .ZN(n6911)
         );
  AOI21_X1 U8548 ( .B1(n9690), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n6911), .ZN(
        n6912) );
  NAND2_X1 U8549 ( .A1(n6913), .A2(n6912), .ZN(P1_U3253) );
  NAND2_X1 U8550 ( .A1(n8165), .A2(n9967), .ZN(n7852) );
  NAND2_X1 U8551 ( .A1(n6937), .A2(n6914), .ZN(n7870) );
  NAND2_X1 U8552 ( .A1(n9934), .A2(n7870), .ZN(n6995) );
  NAND2_X1 U8553 ( .A1(n7803), .A2(n6999), .ZN(n7859) );
  NAND2_X1 U8554 ( .A1(n9916), .A2(n4879), .ZN(n7875) );
  AND2_X1 U8555 ( .A1(n9989), .A2(n9918), .ZN(n6943) );
  INV_X1 U8556 ( .A(n9989), .ZN(n7013) );
  NAND2_X1 U8557 ( .A1(n6944), .A2(n7013), .ZN(n7863) );
  XNOR2_X1 U8558 ( .A(n7884), .B(n8163), .ZN(n7999) );
  NAND2_X1 U8559 ( .A1(n6971), .A2(n7999), .ZN(n6915) );
  NAND2_X1 U8560 ( .A1(n7884), .A2(n7883), .ZN(n7861) );
  NAND2_X1 U8561 ( .A1(n6915), .A2(n7861), .ZN(n6917) );
  OR2_X1 U8562 ( .A1(n10001), .A2(n7062), .ZN(n7886) );
  NAND2_X1 U8563 ( .A1(n10001), .A2(n7062), .ZN(n7887) );
  NAND2_X1 U8564 ( .A1(n7886), .A2(n7887), .ZN(n7882) );
  NAND2_X1 U8565 ( .A1(n6917), .A2(n7882), .ZN(n6918) );
  NAND3_X1 U8566 ( .A1(n7065), .A2(n9938), .A3(n6918), .ZN(n6920) );
  INV_X1 U8567 ( .A(n8426), .ZN(n9915) );
  AOI22_X1 U8568 ( .A1(n8161), .A2(n9917), .B1(n9915), .B2(n8163), .ZN(n6919)
         );
  AND2_X1 U8569 ( .A1(n6920), .A2(n6919), .ZN(n10007) );
  NAND2_X1 U8570 ( .A1(n6922), .A2(n6921), .ZN(n6924) );
  NAND2_X1 U8571 ( .A1(n6927), .A2(n9924), .ZN(n8406) );
  INV_X2 U8572 ( .A(n8406), .ZN(n9941) );
  AND2_X1 U8573 ( .A1(n7009), .A2(n9989), .ZN(n7007) );
  NAND2_X1 U8574 ( .A1(n7007), .A2(n9992), .ZN(n6978) );
  NAND2_X1 U8575 ( .A1(n6978), .A2(n10001), .ZN(n6926) );
  AND2_X1 U8576 ( .A1(n7059), .A2(n6926), .ZN(n10004) );
  INV_X1 U8577 ( .A(n9948), .ZN(n8442) );
  OAI22_X1 U8578 ( .A1(n9927), .A2(n6929), .B1(n6928), .B2(n9924), .ZN(n6932)
         );
  NOR2_X1 U8579 ( .A1(n7991), .A2(n7249), .ZN(n6930) );
  NAND2_X1 U8580 ( .A1(n9927), .A2(n6930), .ZN(n9951) );
  NOR2_X1 U8581 ( .A1(n9951), .A2(n4885), .ZN(n6931) );
  AOI211_X1 U8582 ( .C1(n10004), .C2(n8442), .A(n6932), .B(n6931), .ZN(n6949)
         );
  OAI21_X1 U8583 ( .B1(n6934), .B2(n6933), .A(n7804), .ZN(n6936) );
  NAND2_X1 U8584 ( .A1(n6934), .A2(n6933), .ZN(n6935) );
  NAND2_X1 U8585 ( .A1(n6936), .A2(n6935), .ZN(n9943) );
  NAND2_X1 U8586 ( .A1(n9943), .A2(n9942), .ZN(n6939) );
  NAND2_X1 U8587 ( .A1(n6937), .A2(n9967), .ZN(n6938) );
  NAND2_X1 U8588 ( .A1(n6939), .A2(n6938), .ZN(n6994) );
  NAND2_X1 U8589 ( .A1(n7803), .A2(n4879), .ZN(n6940) );
  NAND2_X1 U8590 ( .A1(n9921), .A2(n9920), .ZN(n6942) );
  NAND2_X1 U8591 ( .A1(n4755), .A2(n9981), .ZN(n6941) );
  NAND2_X1 U8592 ( .A1(n6942), .A2(n6941), .ZN(n7004) );
  INV_X1 U8593 ( .A(n6943), .ZN(n7877) );
  NAND2_X1 U8594 ( .A1(n7863), .A2(n7877), .ZN(n7997) );
  AND2_X1 U8595 ( .A1(n7884), .A2(n8163), .ZN(n6945) );
  XNOR2_X1 U8596 ( .A(n7061), .B(n7882), .ZN(n10000) );
  OR2_X1 U8597 ( .A1(n6946), .A2(n8340), .ZN(n7173) );
  NAND2_X1 U8598 ( .A1(n7064), .A2(n7173), .ZN(n6947) );
  NAND2_X1 U8599 ( .A1(n10000), .A2(n9944), .ZN(n6948) );
  OAI211_X1 U8600 ( .C1(n10007), .C2(n9941), .A(n6949), .B(n6948), .ZN(
        P2_U3289) );
  INV_X1 U8601 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10377) );
  INV_X1 U8602 ( .A(n7743), .ZN(n9058) );
  OAI222_X1 U8603 ( .A1(n7622), .A2(n10377), .B1(n8036), .B2(n6950), .C1(n9058), .C2(P1_U3084), .ZN(P1_U3336) );
  INV_X1 U8604 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n6960) );
  NAND2_X1 U8605 ( .A1(n6962), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6951) );
  INV_X1 U8606 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6953) );
  MUX2_X1 U8607 ( .A(n6953), .B(P2_REG1_REG_10__SCAN_IN), .S(n7050), .Z(n6954)
         );
  NOR2_X1 U8608 ( .A1(n6955), .A2(n6954), .ZN(n7049) );
  AOI21_X1 U8609 ( .B1(n6955), .B2(n6954), .A(n7049), .ZN(n6956) );
  NAND2_X1 U8610 ( .A1(n9904), .A2(n6956), .ZN(n6959) );
  NOR2_X1 U8611 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6957), .ZN(n8055) );
  INV_X1 U8612 ( .A(n8055), .ZN(n6958) );
  OAI211_X1 U8613 ( .C1(n6960), .C2(n8242), .A(n6959), .B(n6958), .ZN(n6967)
         );
  NAND2_X1 U8614 ( .A1(n7050), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6963) );
  OAI21_X1 U8615 ( .B1(n7050), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6963), .ZN(
        n6964) );
  AOI211_X1 U8616 ( .C1(n6965), .C2(n6964), .A(n7044), .B(n9907), .ZN(n6966)
         );
  AOI211_X1 U8617 ( .C1(n9527), .C2(n7050), .A(n6967), .B(n6966), .ZN(n6968)
         );
  INV_X1 U8618 ( .A(n6968), .ZN(P2_U3255) );
  INV_X1 U8619 ( .A(n7999), .ZN(n6969) );
  XNOR2_X1 U8620 ( .A(n6970), .B(n6969), .ZN(n9996) );
  XNOR2_X1 U8621 ( .A(n6971), .B(n7999), .ZN(n6974) );
  NAND2_X1 U8622 ( .A1(n9918), .A2(n9915), .ZN(n6972) );
  OAI21_X1 U8623 ( .B1(n7062), .B2(n8428), .A(n6972), .ZN(n6973) );
  AOI21_X1 U8624 ( .B1(n6974), .B2(n9938), .A(n6973), .ZN(n9999) );
  OAI21_X1 U8625 ( .B1(n6975), .B2(n9924), .A(n9999), .ZN(n6976) );
  NAND2_X1 U8626 ( .A1(n6976), .A2(n9927), .ZN(n6982) );
  OR2_X1 U8627 ( .A1(n7007), .A2(n9992), .ZN(n6977) );
  NAND2_X1 U8628 ( .A1(n6978), .A2(n6977), .ZN(n9993) );
  OAI22_X1 U8629 ( .A1(n9948), .A2(n9993), .B1(n9927), .B2(n6979), .ZN(n6980)
         );
  AOI21_X1 U8630 ( .B1(n8490), .B2(n7884), .A(n6980), .ZN(n6981) );
  OAI211_X1 U8631 ( .C1(n9996), .C2(n8478), .A(n6982), .B(n6981), .ZN(P2_U3290) );
  AND2_X1 U8632 ( .A1(n6983), .A2(n7867), .ZN(n7995) );
  INV_X1 U8633 ( .A(n7995), .ZN(n9964) );
  AOI22_X1 U8634 ( .A1(n9964), .A2(n9938), .B1(n9917), .B2(n4941), .ZN(n9966)
         );
  OAI22_X1 U8635 ( .A1(n9941), .A2(n9966), .B1(n6984), .B2(n9924), .ZN(n6985)
         );
  AOI21_X1 U8636 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n9941), .A(n6985), .ZN(
        n6987) );
  OAI21_X1 U8637 ( .B1(n8490), .B2(n8442), .A(n9963), .ZN(n6986) );
  OAI211_X1 U8638 ( .C1(n7995), .C2(n8478), .A(n6987), .B(n6986), .ZN(P2_U3296) );
  AOI22_X1 U8639 ( .A1(n8490), .A2(n7716), .B1(n9944), .B2(n6988), .ZN(n6992)
         );
  OAI22_X1 U8640 ( .A1(n6569), .A2(n9927), .B1(n10448), .B2(n9924), .ZN(n6989)
         );
  AOI21_X1 U8641 ( .B1(n8442), .B2(n6990), .A(n6989), .ZN(n6991) );
  OAI211_X1 U8642 ( .C1(n9941), .C2(n6993), .A(n6992), .B(n6991), .ZN(P2_U3295) );
  XNOR2_X1 U8643 ( .A(n6994), .B(n7858), .ZN(n9976) );
  XNOR2_X1 U8644 ( .A(n6995), .B(n7858), .ZN(n6996) );
  NAND2_X1 U8645 ( .A1(n6996), .A2(n9938), .ZN(n6998) );
  NAND2_X1 U8646 ( .A1(n6998), .A2(n6997), .ZN(n9975) );
  AOI22_X1 U8647 ( .A1(n8490), .A2(n6999), .B1(n9975), .B2(n9927), .ZN(n7003)
         );
  NAND2_X1 U8648 ( .A1(n9947), .A2(n6999), .ZN(n7000) );
  NAND2_X1 U8649 ( .A1(n9923), .A2(n7000), .ZN(n9973) );
  OAI22_X1 U8650 ( .A1(n9948), .A2(n9973), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9924), .ZN(n7001) );
  AOI21_X1 U8651 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n9941), .A(n7001), .ZN(
        n7002) );
  OAI211_X1 U8652 ( .C1(n9976), .C2(n8478), .A(n7003), .B(n7002), .ZN(P2_U3293) );
  XNOR2_X1 U8653 ( .A(n7004), .B(n7997), .ZN(n9991) );
  INV_X1 U8654 ( .A(n9991), .ZN(n7016) );
  XNOR2_X1 U8655 ( .A(n7005), .B(n7997), .ZN(n7006) );
  AOI222_X1 U8656 ( .A1(n9938), .A2(n7006), .B1(n8163), .B2(n9917), .C1(n8164), 
        .C2(n9915), .ZN(n9988) );
  INV_X1 U8657 ( .A(n9988), .ZN(n7012) );
  INV_X1 U8658 ( .A(n7007), .ZN(n7008) );
  OAI211_X1 U8659 ( .C1(n9989), .C2(n7009), .A(n7008), .B(n10003), .ZN(n9987)
         );
  OAI22_X1 U8660 ( .A1(n9987), .A2(n8356), .B1(n9924), .B2(n7010), .ZN(n7011)
         );
  OAI21_X1 U8661 ( .B1(n7012), .B2(n7011), .A(n8406), .ZN(n7015) );
  AOI22_X1 U8662 ( .A1(n8490), .A2(n7013), .B1(n9941), .B2(
        P2_REG2_REG_5__SCAN_IN), .ZN(n7014) );
  OAI211_X1 U8663 ( .C1(n7016), .C2(n8478), .A(n7015), .B(n7014), .ZN(P2_U3291) );
  OAI21_X1 U8664 ( .B1(n7018), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7017), .ZN(
        n7021) );
  MUX2_X1 U8665 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7019), .S(n7228), .Z(n7020)
         );
  NAND2_X1 U8666 ( .A1(n7020), .A2(n7021), .ZN(n7220) );
  OAI21_X1 U8667 ( .B1(n7021), .B2(n7020), .A(n7220), .ZN(n7022) );
  NAND2_X1 U8668 ( .A1(n7022), .A2(n9720), .ZN(n7034) );
  OR2_X1 U8669 ( .A1(n7228), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7026) );
  NAND2_X1 U8670 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7228), .ZN(n7025) );
  NAND2_X1 U8671 ( .A1(n7026), .A2(n7025), .ZN(n7027) );
  AOI21_X1 U8672 ( .B1(n7028), .B2(n7027), .A(n7227), .ZN(n7029) );
  NAND2_X1 U8673 ( .A1(n9711), .A2(n7029), .ZN(n7030) );
  NAND2_X1 U8674 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7591) );
  OAI211_X1 U8675 ( .C1(n9715), .C2(n7031), .A(n7030), .B(n7591), .ZN(n7032)
         );
  AOI21_X1 U8676 ( .B1(n9690), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n7032), .ZN(
        n7033) );
  NAND2_X1 U8677 ( .A1(n7034), .A2(n7033), .ZN(P1_U3254) );
  XNOR2_X1 U8678 ( .A(n7036), .B(n7035), .ZN(n7037) );
  XNOR2_X1 U8679 ( .A(n7038), .B(n7037), .ZN(n7039) );
  NAND2_X1 U8680 ( .A1(n7039), .A2(n8732), .ZN(n7043) );
  OAI22_X1 U8681 ( .A1(n8736), .A2(n7334), .B1(n8735), .B2(n7348), .ZN(n7040)
         );
  AOI211_X1 U8682 ( .C1(n8740), .C2(n9855), .A(n7041), .B(n7040), .ZN(n7042)
         );
  OAI211_X1 U8683 ( .C1(n9861), .C2(n8743), .A(n7043), .B(n7042), .ZN(P1_U3211) );
  INV_X1 U8684 ( .A(n9527), .ZN(n9906) );
  AOI22_X1 U8685 ( .A1(n7242), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7277), .B2(
        n7058), .ZN(n7045) );
  NAND2_X1 U8686 ( .A1(n7046), .A2(n7045), .ZN(n7241) );
  OAI21_X1 U8687 ( .B1(n7046), .B2(n7045), .A(n7241), .ZN(n7047) );
  INV_X1 U8688 ( .A(n9907), .ZN(n9903) );
  NAND2_X1 U8689 ( .A1(n7047), .A2(n9903), .ZN(n7057) );
  INV_X1 U8690 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7048) );
  NOR2_X1 U8691 ( .A1(n8242), .A2(n7048), .ZN(n7055) );
  AOI21_X1 U8692 ( .B1(n7050), .B2(P2_REG1_REG_10__SCAN_IN), .A(n7049), .ZN(
        n7053) );
  INV_X1 U8693 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7051) );
  MUX2_X1 U8694 ( .A(n7051), .B(P2_REG1_REG_11__SCAN_IN), .S(n7242), .Z(n7052)
         );
  NOR2_X1 U8695 ( .A1(n7053), .A2(n7052), .ZN(n7235) );
  INV_X1 U8696 ( .A(n9904), .ZN(n8199) );
  AOI211_X1 U8697 ( .C1(n7053), .C2(n7052), .A(n7235), .B(n8199), .ZN(n7054)
         );
  AOI211_X1 U8698 ( .C1(P2_REG3_REG_11__SCAN_IN), .C2(P2_U3152), .A(n7055), 
        .B(n7054), .ZN(n7056) );
  OAI211_X1 U8699 ( .C1(n9906), .C2(n7058), .A(n7057), .B(n7056), .ZN(P2_U3256) );
  NAND2_X1 U8700 ( .A1(n7059), .A2(n7112), .ZN(n7060) );
  NAND2_X1 U8701 ( .A1(n7186), .A2(n7060), .ZN(n10008) );
  INV_X1 U8702 ( .A(n7062), .ZN(n8162) );
  OR2_X1 U8703 ( .A1(n10001), .A2(n8162), .ZN(n7063) );
  OR2_X1 U8704 ( .A1(n7112), .A2(n7177), .ZN(n7889) );
  NAND2_X1 U8705 ( .A1(n7112), .A2(n7177), .ZN(n7890) );
  NAND2_X1 U8706 ( .A1(n7889), .A2(n7890), .ZN(n7111) );
  XNOR2_X1 U8707 ( .A(n7110), .B(n7111), .ZN(n10012) );
  INV_X1 U8708 ( .A(n10012), .ZN(n7070) );
  INV_X1 U8709 ( .A(n7064), .ZN(n9978) );
  NAND2_X1 U8710 ( .A1(n7066), .A2(n7111), .ZN(n7067) );
  INV_X1 U8711 ( .A(n9938), .ZN(n8425) );
  AOI21_X1 U8712 ( .B1(n7102), .B2(n7067), .A(n8425), .ZN(n7068) );
  AOI211_X1 U8713 ( .C1(n9978), .C2(n10012), .A(n7069), .B(n7068), .ZN(n10009)
         );
  OAI21_X1 U8714 ( .B1(n7070), .B2(n7173), .A(n10009), .ZN(n7071) );
  NAND2_X1 U8715 ( .A1(n7071), .A2(n8406), .ZN(n7076) );
  OAI22_X1 U8716 ( .A1(n9927), .A2(n7073), .B1(n7072), .B2(n9924), .ZN(n7074)
         );
  AOI21_X1 U8717 ( .B1(n8490), .B2(n7112), .A(n7074), .ZN(n7075) );
  OAI211_X1 U8718 ( .C1(n9948), .C2(n10008), .A(n7076), .B(n7075), .ZN(
        P2_U3288) );
  INV_X1 U8719 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10238) );
  INV_X1 U8720 ( .A(n7077), .ZN(n7078) );
  INV_X1 U8721 ( .A(n7744), .ZN(n9714) );
  OAI222_X1 U8722 ( .A1(n7622), .A2(n10238), .B1(n8036), .B2(n7078), .C1(
        P1_U3084), .C2(n9714), .ZN(P1_U3335) );
  INV_X1 U8723 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7079) );
  INV_X1 U8724 ( .A(n8232), .ZN(n8225) );
  OAI222_X1 U8725 ( .A1(n7729), .A2(n7079), .B1(n8612), .B2(n7078), .C1(
        P2_U3152), .C2(n8225), .ZN(P2_U3340) );
  INV_X1 U8726 ( .A(n7081), .ZN(n7082) );
  AOI21_X1 U8727 ( .B1(n7084), .B2(n7083), .A(n7082), .ZN(n7089) );
  OAI21_X1 U8728 ( .B1(n8128), .B2(n7182), .A(n7085), .ZN(n7087) );
  OAI22_X1 U8729 ( .A1(n8131), .A2(n8158), .B1(n7177), .B2(n8129), .ZN(n7086)
         );
  AOI211_X1 U8730 ( .C1(n8143), .C2(n10014), .A(n7087), .B(n7086), .ZN(n7088)
         );
  OAI21_X1 U8731 ( .B1(n7089), .B2(n8145), .A(n7088), .ZN(P2_U3233) );
  INV_X1 U8732 ( .A(n7090), .ZN(n7091) );
  NOR2_X1 U8733 ( .A1(n7092), .A2(n7091), .ZN(n7190) );
  AOI21_X1 U8734 ( .B1(n7092), .B2(n7091), .A(n7190), .ZN(n7093) );
  NAND2_X1 U8735 ( .A1(n7093), .A2(n7094), .ZN(n7192) );
  OAI21_X1 U8736 ( .B1(n7094), .B2(n7093), .A(n7192), .ZN(n7095) );
  NAND2_X1 U8737 ( .A1(n7095), .A2(n8732), .ZN(n7101) );
  INV_X1 U8738 ( .A(n7096), .ZN(n7099) );
  INV_X1 U8739 ( .A(n9753), .ZN(n7097) );
  INV_X1 U8740 ( .A(n9035), .ZN(n9758) );
  OAI22_X1 U8741 ( .A1(n8736), .A2(n7097), .B1(n8723), .B2(n9758), .ZN(n7098)
         );
  AOI211_X1 U8742 ( .C1(n8725), .C2(n9855), .A(n7099), .B(n7098), .ZN(n7100)
         );
  OAI211_X1 U8743 ( .C1(n9839), .C2(n8743), .A(n7101), .B(n7100), .ZN(P1_U3225) );
  NAND2_X1 U8744 ( .A1(n7102), .A2(n7890), .ZN(n7176) );
  OR2_X1 U8745 ( .A1(n10014), .A2(n7114), .ZN(n7893) );
  NAND2_X1 U8746 ( .A1(n10014), .A2(n7114), .ZN(n7897) );
  AND2_X1 U8747 ( .A1(n7893), .A2(n7897), .ZN(n7113) );
  NAND2_X1 U8748 ( .A1(n7176), .A2(n7113), .ZN(n7103) );
  NAND2_X1 U8749 ( .A1(n7103), .A2(n7897), .ZN(n7104) );
  OR2_X1 U8750 ( .A1(n7119), .A2(n8158), .ZN(n7894) );
  NAND2_X1 U8751 ( .A1(n7119), .A2(n8158), .ZN(n7899) );
  AOI21_X1 U8752 ( .B1(n7104), .B2(n8004), .A(n8425), .ZN(n7109) );
  INV_X1 U8753 ( .A(n7104), .ZN(n7106) );
  OR2_X1 U8754 ( .A1(n7392), .A2(n8428), .ZN(n7108) );
  OR2_X1 U8755 ( .A1(n7114), .A2(n8426), .ZN(n7107) );
  NAND2_X1 U8756 ( .A1(n7108), .A2(n7107), .ZN(n8056) );
  AOI21_X1 U8757 ( .B1(n7109), .B2(n7271), .A(n8056), .ZN(n10027) );
  INV_X1 U8758 ( .A(n7111), .ZN(n8001) );
  NAND2_X1 U8759 ( .A1(n7175), .A2(n8003), .ZN(n7174) );
  INV_X1 U8760 ( .A(n7114), .ZN(n8160) );
  OR2_X1 U8761 ( .A1(n10014), .A2(n8160), .ZN(n7115) );
  XNOR2_X1 U8762 ( .A(n7269), .B(n8004), .ZN(n10021) );
  INV_X1 U8763 ( .A(n7119), .ZN(n10022) );
  NOR2_X1 U8764 ( .A1(n7185), .A2(n10022), .ZN(n7116) );
  OR2_X1 U8765 ( .A1(n7377), .A2(n7116), .ZN(n10023) );
  OAI22_X1 U8766 ( .A1(n9927), .A2(n7117), .B1(n8057), .B2(n9924), .ZN(n7118)
         );
  AOI21_X1 U8767 ( .B1(n8490), .B2(n7119), .A(n7118), .ZN(n7120) );
  OAI21_X1 U8768 ( .B1(n10023), .B2(n9948), .A(n7120), .ZN(n7121) );
  AOI21_X1 U8769 ( .B1(n10021), .B2(n9944), .A(n7121), .ZN(n7122) );
  OAI21_X1 U8770 ( .B1(n10027), .B2(n9941), .A(n7122), .ZN(P2_U3286) );
  AND2_X1 U8771 ( .A1(n7123), .A2(n9799), .ZN(n7125) );
  NAND2_X1 U8772 ( .A1(n7125), .A2(n7124), .ZN(n7153) );
  OAI21_X1 U8773 ( .B1(n8959), .B2(n7125), .A(n7153), .ZN(n9811) );
  INV_X1 U8774 ( .A(n7126), .ZN(n7127) );
  NAND2_X1 U8775 ( .A1(n7128), .A2(n7127), .ZN(n7132) );
  OAI21_X1 U8776 ( .B1(n7130), .B2(P1_D_REG_0__SCAN_IN), .A(n7129), .ZN(n7131)
         );
  AND2_X1 U8777 ( .A1(n7132), .A2(n7131), .ZN(n7500) );
  INV_X1 U8778 ( .A(n7500), .ZN(n7133) );
  OR2_X1 U8779 ( .A1(n9023), .A2(n7492), .ZN(n9809) );
  NOR2_X1 U8780 ( .A1(n7133), .A2(n9809), .ZN(n7166) );
  NAND2_X1 U8781 ( .A1(n7166), .A2(n7489), .ZN(n7134) );
  OR2_X1 U8782 ( .A1(n7135), .A2(n9761), .ZN(n7136) );
  NOR2_X1 U8783 ( .A1(n9779), .A2(n7136), .ZN(n9788) );
  INV_X1 U8784 ( .A(n9788), .ZN(n9577) );
  NAND3_X1 U8785 ( .A1(n7304), .A2(n9791), .A3(n9761), .ZN(n9849) );
  INV_X1 U8786 ( .A(n8872), .ZN(n7138) );
  NAND2_X1 U8787 ( .A1(n7137), .A2(n7138), .ZN(n9757) );
  INV_X1 U8788 ( .A(n9757), .ZN(n9856) );
  AOI22_X1 U8789 ( .A1(n9856), .A2(n8886), .B1(n7151), .B2(n9857), .ZN(n7143)
         );
  OAI21_X1 U8790 ( .B1(n7139), .B2(n8955), .A(n7159), .ZN(n7141) );
  NAND2_X1 U8791 ( .A1(n9024), .A2(n8871), .ZN(n7140) );
  NAND2_X1 U8792 ( .A1(n8947), .A2(n4721), .ZN(n8745) );
  NAND2_X1 U8793 ( .A1(n7140), .A2(n8745), .ZN(n9427) );
  NAND2_X1 U8794 ( .A1(n7141), .A2(n9427), .ZN(n7142) );
  OAI211_X1 U8795 ( .C1(n9811), .C2(n9849), .A(n7143), .B(n7142), .ZN(n9814)
         );
  OR2_X1 U8796 ( .A1(n9797), .A2(n4721), .ZN(n9749) );
  INV_X1 U8797 ( .A(n9749), .ZN(n9785) );
  OAI211_X1 U8798 ( .C1(n4773), .C2(n9813), .A(n9785), .B(n7164), .ZN(n9812)
         );
  OAI22_X1 U8799 ( .A1(n9812), .A2(n8871), .B1(n9319), .B2(n7144), .ZN(n7145)
         );
  INV_X1 U8800 ( .A(n9779), .ZN(n9222) );
  OAI21_X1 U8801 ( .B1(n9814), .B2(n7145), .A(n9222), .ZN(n7147) );
  AOI22_X1 U8802 ( .A1(n9572), .A2(n8888), .B1(n9779), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7146) );
  OAI211_X1 U8803 ( .C1(n9811), .C2(n9577), .A(n7147), .B(n7146), .ZN(P1_U3290) );
  INV_X1 U8804 ( .A(n7148), .ZN(n7149) );
  OAI222_X1 U8805 ( .A1(n7622), .A2(n10389), .B1(n8036), .B2(n7149), .C1(
        P1_U3084), .C2(n9761), .ZN(P1_U3334) );
  OAI222_X1 U8806 ( .A1(n7729), .A2(n7150), .B1(n8612), .B2(n7149), .C1(n8340), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OR2_X1 U8807 ( .A1(n7151), .A2(n9819), .ZN(n8890) );
  NAND2_X1 U8808 ( .A1(n7151), .A2(n9819), .ZN(n8892) );
  NAND2_X1 U8809 ( .A1(n8890), .A2(n8892), .ZN(n7154) );
  NAND2_X1 U8810 ( .A1(n9794), .A2(n8888), .ZN(n7152) );
  NAND2_X1 U8811 ( .A1(n7153), .A2(n7152), .ZN(n7157) );
  INV_X1 U8812 ( .A(n7157), .ZN(n7155) );
  NAND2_X1 U8813 ( .A1(n7155), .A2(n7154), .ZN(n7254) );
  INV_X1 U8814 ( .A(n7254), .ZN(n7156) );
  AOI21_X1 U8815 ( .B1(n8956), .B2(n7157), .A(n7156), .ZN(n9817) );
  AOI22_X1 U8816 ( .A1(n9856), .A2(n9794), .B1(n9773), .B2(n9857), .ZN(n7162)
         );
  OR2_X1 U8817 ( .A1(n9794), .A2(n9813), .ZN(n7158) );
  OAI21_X1 U8818 ( .B1(n8956), .B2(n8894), .A(n7259), .ZN(n7160) );
  NAND2_X1 U8819 ( .A1(n7160), .A2(n9427), .ZN(n7161) );
  OAI211_X1 U8820 ( .C1(n9817), .C2(n9849), .A(n7162), .B(n7161), .ZN(n9820)
         );
  NAND2_X1 U8821 ( .A1(n9820), .A2(n9222), .ZN(n7172) );
  NAND2_X1 U8822 ( .A1(n8698), .A2(n7164), .ZN(n7163) );
  NAND2_X1 U8823 ( .A1(n7163), .A2(n9785), .ZN(n7165) );
  OR2_X1 U8824 ( .A1(n7165), .A2(n7256), .ZN(n9818) );
  AND2_X1 U8825 ( .A1(n7166), .A2(n9761), .ZN(n9787) );
  INV_X1 U8826 ( .A(n9787), .ZN(n9576) );
  NOR2_X1 U8827 ( .A1(n9818), .A2(n9576), .ZN(n7170) );
  INV_X1 U8828 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7167) );
  OAI22_X1 U8829 ( .A1(n9222), .A2(n7168), .B1(n7167), .B2(n9319), .ZN(n7169)
         );
  AOI211_X1 U8830 ( .C1(n9572), .C2(n8698), .A(n7170), .B(n7169), .ZN(n7171)
         );
  OAI211_X1 U8831 ( .C1(n9817), .C2(n9577), .A(n7172), .B(n7171), .ZN(P1_U3289) );
  INV_X1 U8832 ( .A(n7173), .ZN(n7181) );
  OAI21_X1 U8833 ( .B1(n7175), .B2(n8003), .A(n7174), .ZN(n10019) );
  XNOR2_X1 U8834 ( .A(n7176), .B(n8003), .ZN(n7180) );
  OAI22_X1 U8835 ( .A1(n7177), .A2(n8426), .B1(n8158), .B2(n8428), .ZN(n7178)
         );
  AOI21_X1 U8836 ( .B1(n10019), .B2(n9978), .A(n7178), .ZN(n7179) );
  OAI21_X1 U8837 ( .B1(n8425), .B2(n7180), .A(n7179), .ZN(n10017) );
  AOI21_X1 U8838 ( .B1(n7181), .B2(n10019), .A(n10017), .ZN(n7189) );
  OAI22_X1 U8839 ( .A1(n9927), .A2(n7183), .B1(n7182), .B2(n9924), .ZN(n7184)
         );
  AOI21_X1 U8840 ( .B1(n8490), .B2(n10014), .A(n7184), .ZN(n7188) );
  AOI21_X1 U8841 ( .B1(n10014), .B2(n7186), .A(n7185), .ZN(n10013) );
  NAND2_X1 U8842 ( .A1(n10013), .A2(n8442), .ZN(n7187) );
  OAI211_X1 U8843 ( .C1(n7189), .C2(n9941), .A(n7188), .B(n7187), .ZN(P2_U3287) );
  INV_X1 U8844 ( .A(n7190), .ZN(n7191) );
  NAND2_X1 U8845 ( .A1(n7192), .A2(n7191), .ZN(n7197) );
  INV_X1 U8846 ( .A(n7193), .ZN(n7195) );
  NOR2_X1 U8847 ( .A1(n7195), .A2(n7194), .ZN(n7196) );
  XNOR2_X1 U8848 ( .A(n7197), .B(n7196), .ZN(n7198) );
  NAND2_X1 U8849 ( .A1(n7198), .A2(n8732), .ZN(n7203) );
  INV_X1 U8850 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7199) );
  NOR2_X1 U8851 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7199), .ZN(n9655) );
  INV_X1 U8852 ( .A(n9844), .ZN(n7200) );
  OAI22_X1 U8853 ( .A1(n8736), .A2(n7407), .B1(n8723), .B2(n7200), .ZN(n7201)
         );
  AOI211_X1 U8854 ( .C1(n8725), .C2(n9843), .A(n9655), .B(n7201), .ZN(n7202)
         );
  OAI211_X1 U8855 ( .C1(n9847), .C2(n8743), .A(n7203), .B(n7202), .ZN(P1_U3237) );
  XNOR2_X1 U8856 ( .A(n7205), .B(n7204), .ZN(n7209) );
  OAI22_X1 U8857 ( .A1(n8128), .A2(n7276), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5375), .ZN(n7207) );
  OAI22_X1 U8858 ( .A1(n8131), .A2(n7449), .B1(n8158), .B2(n8129), .ZN(n7206)
         );
  AOI211_X1 U8859 ( .C1(n8143), .C2(n7372), .A(n7207), .B(n7206), .ZN(n7208)
         );
  OAI21_X1 U8860 ( .B1(n7209), .B2(n8145), .A(n7208), .ZN(P2_U3238) );
  INV_X1 U8861 ( .A(n7322), .ZN(n9870) );
  XNOR2_X1 U8862 ( .A(n7212), .B(n7211), .ZN(n7213) );
  XNOR2_X1 U8863 ( .A(n7210), .B(n7213), .ZN(n7214) );
  NAND2_X1 U8864 ( .A1(n7214), .A2(n8732), .ZN(n7218) );
  INV_X1 U8865 ( .A(n9034), .ZN(n9736) );
  OAI22_X1 U8866 ( .A1(n8736), .A2(n9739), .B1(n8735), .B2(n9736), .ZN(n7215)
         );
  AOI211_X1 U8867 ( .C1(n8740), .C2(n9843), .A(n7216), .B(n7215), .ZN(n7217)
         );
  OAI211_X1 U8868 ( .C1(n9870), .C2(n8743), .A(n7218), .B(n7217), .ZN(P1_U3219) );
  NOR2_X1 U8869 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7219), .ZN(n7692) );
  INV_X1 U8870 ( .A(n7692), .ZN(n7226) );
  OAI21_X1 U8871 ( .B1(n7228), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7220), .ZN(
        n7223) );
  MUX2_X1 U8872 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n7221), .S(n7507), .Z(n7222)
         );
  NAND2_X1 U8873 ( .A1(n7222), .A2(n7223), .ZN(n7506) );
  OAI21_X1 U8874 ( .B1(n7223), .B2(n7222), .A(n7506), .ZN(n7224) );
  NAND2_X1 U8875 ( .A1(n9720), .A2(n7224), .ZN(n7225) );
  OAI211_X1 U8876 ( .C1(n9715), .C2(n7513), .A(n7226), .B(n7225), .ZN(n7231)
         );
  AOI211_X1 U8877 ( .C1(n7229), .C2(n7611), .A(n7515), .B(n9682), .ZN(n7230)
         );
  AOI211_X1 U8878 ( .C1(P1_ADDR_REG_14__SCAN_IN), .C2(n9690), .A(n7231), .B(
        n7230), .ZN(n7232) );
  INV_X1 U8879 ( .A(n7232), .ZN(P1_U3255) );
  INV_X1 U8880 ( .A(n7233), .ZN(n7248) );
  OAI222_X1 U8881 ( .A1(n7622), .A2(n10451), .B1(n8036), .B2(n7248), .C1(n7234), .C2(P1_U3084), .ZN(P1_U3333) );
  INV_X1 U8882 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7240) );
  AOI21_X1 U8883 ( .B1(n7242), .B2(P2_REG1_REG_11__SCAN_IN), .A(n7235), .ZN(
        n7237) );
  MUX2_X1 U8884 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7289), .S(n7283), .Z(n7236)
         );
  NAND2_X1 U8885 ( .A1(n7237), .A2(n7236), .ZN(n7292) );
  OAI21_X1 U8886 ( .B1(n7237), .B2(n7236), .A(n7292), .ZN(n7238) );
  NAND2_X1 U8887 ( .A1(n9904), .A2(n7238), .ZN(n7239) );
  NAND2_X1 U8888 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7390) );
  OAI211_X1 U8889 ( .C1(n7240), .C2(n8242), .A(n7239), .B(n7390), .ZN(n7246)
         );
  XNOR2_X1 U8890 ( .A(n7283), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n7244) );
  OAI21_X1 U8891 ( .B1(n7242), .B2(P2_REG2_REG_11__SCAN_IN), .A(n7241), .ZN(
        n7243) );
  AOI211_X1 U8892 ( .C1(n7244), .C2(n7243), .A(n9907), .B(n7282), .ZN(n7245)
         );
  AOI211_X1 U8893 ( .C1(n9527), .C2(n7283), .A(n7246), .B(n7245), .ZN(n7247)
         );
  INV_X1 U8894 ( .A(n7247), .ZN(P2_U3257) );
  OAI222_X1 U8895 ( .A1(n7729), .A2(n7250), .B1(P2_U3152), .B2(n7249), .C1(
        n8612), .C2(n7248), .ZN(P2_U3338) );
  INV_X1 U8896 ( .A(n9773), .ZN(n7252) );
  NAND2_X1 U8897 ( .A1(n7252), .A2(n7251), .ZN(n8989) );
  NAND2_X1 U8898 ( .A1(n9773), .A2(n9825), .ZN(n8895) );
  NAND2_X1 U8899 ( .A1(n8989), .A2(n8895), .ZN(n7306) );
  OR2_X1 U8900 ( .A1(n7151), .A2(n8698), .ZN(n7253) );
  XNOR2_X1 U8901 ( .A(n7306), .B(n7255), .ZN(n9828) );
  NAND2_X1 U8902 ( .A1(n7256), .A2(n9825), .ZN(n9783) );
  OAI211_X1 U8903 ( .C1(n7256), .C2(n9825), .A(n9783), .B(n9785), .ZN(n9824)
         );
  INV_X1 U8904 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7257) );
  AOI22_X1 U8905 ( .A1(n9572), .A2(n7251), .B1(n9804), .B2(n7257), .ZN(n7258)
         );
  OAI21_X1 U8906 ( .B1(n9576), .B2(n9824), .A(n7258), .ZN(n7267) );
  INV_X1 U8907 ( .A(n7306), .ZN(n8957) );
  NAND2_X1 U8908 ( .A1(n7259), .A2(n8890), .ZN(n8993) );
  NAND2_X1 U8909 ( .A1(n8993), .A2(n8957), .ZN(n7315) );
  OAI21_X1 U8910 ( .B1(n8957), .B2(n8993), .A(n7315), .ZN(n7263) );
  NAND2_X1 U8911 ( .A1(n7151), .A2(n9856), .ZN(n7261) );
  NAND2_X1 U8912 ( .A1(n9035), .A2(n9857), .ZN(n7260) );
  NAND2_X1 U8913 ( .A1(n7261), .A2(n7260), .ZN(n7262) );
  AOI21_X1 U8914 ( .B1(n7263), .B2(n9427), .A(n7262), .ZN(n7265) );
  INV_X1 U8915 ( .A(n9849), .ZN(n9886) );
  NAND2_X1 U8916 ( .A1(n9828), .A2(n9886), .ZN(n7264) );
  NAND2_X1 U8917 ( .A1(n7265), .A2(n7264), .ZN(n9826) );
  MUX2_X1 U8918 ( .A(n9826), .B(P1_REG2_REG_3__SCAN_IN), .S(n9807), .Z(n7266)
         );
  AOI211_X1 U8919 ( .C1(n9788), .C2(n9828), .A(n7267), .B(n7266), .ZN(n7268)
         );
  INV_X1 U8920 ( .A(n7268), .ZN(P1_U3288) );
  OR2_X1 U8921 ( .A1(n7372), .A2(n7392), .ZN(n7906) );
  NAND2_X1 U8922 ( .A1(n7372), .A2(n7392), .ZN(n7908) );
  INV_X1 U8923 ( .A(n7273), .ZN(n8005) );
  OAI21_X1 U8924 ( .B1(n7270), .B2(n8005), .A(n7374), .ZN(n10028) );
  OAI21_X1 U8925 ( .B1(n7273), .B2(n7272), .A(n7370), .ZN(n7274) );
  INV_X1 U8926 ( .A(n7274), .ZN(n7275) );
  OAI222_X1 U8927 ( .A1(n8428), .A2(n7449), .B1(n8426), .B2(n8158), .C1(n8425), 
        .C2(n7275), .ZN(n10031) );
  NAND2_X1 U8928 ( .A1(n10031), .A2(n8406), .ZN(n7281) );
  OAI22_X1 U8929 ( .A1(n9927), .A2(n7277), .B1(n7276), .B2(n9924), .ZN(n7279)
         );
  INV_X1 U8930 ( .A(n7372), .ZN(n10029) );
  XNOR2_X1 U8931 ( .A(n7377), .B(n10029), .ZN(n10030) );
  NOR2_X1 U8932 ( .A1(n10030), .A2(n9948), .ZN(n7278) );
  AOI211_X1 U8933 ( .C1(n8490), .C2(n7372), .A(n7279), .B(n7278), .ZN(n7280)
         );
  OAI211_X1 U8934 ( .C1(n8478), .C2(n10028), .A(n7281), .B(n7280), .ZN(
        P2_U3285) );
  NOR2_X1 U8935 ( .A1(n7458), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7284) );
  AOI21_X1 U8936 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n7458), .A(n7284), .ZN(
        n7285) );
  OAI21_X1 U8937 ( .B1(n7286), .B2(n7285), .A(n7454), .ZN(n7287) );
  NAND2_X1 U8938 ( .A1(n7287), .A2(n9903), .ZN(n7301) );
  INV_X1 U8939 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7298) );
  AOI22_X1 U8940 ( .A1(n7458), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n5427), .B2(
        n7288), .ZN(n7294) );
  NAND2_X1 U8941 ( .A1(n7290), .A2(n7289), .ZN(n7291) );
  NAND2_X1 U8942 ( .A1(n7292), .A2(n7291), .ZN(n7293) );
  NAND2_X1 U8943 ( .A1(n7294), .A2(n7293), .ZN(n7457) );
  OAI21_X1 U8944 ( .B1(n7294), .B2(n7293), .A(n7457), .ZN(n7295) );
  NAND2_X1 U8945 ( .A1(n9904), .A2(n7295), .ZN(n7297) );
  NAND2_X1 U8946 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7296) );
  OAI211_X1 U8947 ( .C1(n8242), .C2(n7298), .A(n7297), .B(n7296), .ZN(n7299)
         );
  AOI21_X1 U8948 ( .B1(n7458), .B2(n9527), .A(n7299), .ZN(n7300) );
  NAND2_X1 U8949 ( .A1(n7301), .A2(n7300), .ZN(P2_U3258) );
  INV_X1 U8950 ( .A(n7302), .ZN(n7330) );
  OAI222_X1 U8951 ( .A1(n7622), .A2(n7303), .B1(n8036), .B2(n7330), .C1(n9013), 
        .C2(P1_U3084), .ZN(P1_U3332) );
  NAND2_X1 U8952 ( .A1(n7304), .A2(n9791), .ZN(n7305) );
  OR2_X1 U8953 ( .A1(n9773), .A2(n7251), .ZN(n7307) );
  NAND2_X1 U8954 ( .A1(n7308), .A2(n7307), .ZN(n9770) );
  OR2_X1 U8955 ( .A1(n9035), .A2(n9831), .ZN(n8899) );
  OR2_X1 U8956 ( .A1(n9035), .A2(n7321), .ZN(n7309) );
  NAND2_X1 U8957 ( .A1(n9844), .A2(n9839), .ZN(n7397) );
  NAND2_X1 U8958 ( .A1(n9844), .A2(n9750), .ZN(n7310) );
  AND2_X1 U8959 ( .A1(n9763), .A2(n7310), .ZN(n7403) );
  OR2_X1 U8960 ( .A1(n9855), .A2(n9847), .ZN(n8772) );
  NAND2_X1 U8961 ( .A1(n9855), .A2(n9847), .ZN(n8764) );
  NAND2_X1 U8962 ( .A1(n8772), .A2(n8764), .ZN(n8757) );
  NAND2_X1 U8963 ( .A1(n7403), .A2(n8757), .ZN(n7402) );
  OR2_X1 U8964 ( .A1(n9855), .A2(n7412), .ZN(n7311) );
  NAND2_X1 U8965 ( .A1(n7402), .A2(n7311), .ZN(n7341) );
  NAND2_X1 U8966 ( .A1(n9843), .A2(n9861), .ZN(n8901) );
  NAND2_X1 U8967 ( .A1(n9730), .A2(n8901), .ZN(n8961) );
  INV_X1 U8968 ( .A(n9861), .ZN(n7340) );
  OR2_X1 U8969 ( .A1(n7340), .A2(n9843), .ZN(n7312) );
  NAND2_X1 U8970 ( .A1(n7348), .A2(n7322), .ZN(n8778) );
  INV_X1 U8971 ( .A(n7348), .ZN(n9858) );
  NAND2_X1 U8972 ( .A1(n9870), .A2(n9858), .ZN(n8774) );
  NAND2_X1 U8973 ( .A1(n7322), .A2(n9858), .ZN(n7314) );
  OR2_X1 U8974 ( .A1(n9879), .A2(n9736), .ZN(n8780) );
  NAND2_X1 U8975 ( .A1(n9879), .A2(n9736), .ZN(n8777) );
  NAND2_X1 U8976 ( .A1(n8780), .A2(n8777), .ZN(n8966) );
  XNOR2_X1 U8977 ( .A(n7360), .B(n8966), .ZN(n9882) );
  INV_X1 U8978 ( .A(n9427), .ZN(n9862) );
  NAND2_X1 U8979 ( .A1(n7315), .A2(n8989), .ZN(n9772) );
  INV_X1 U8980 ( .A(n8899), .ZN(n7316) );
  AND2_X1 U8981 ( .A1(n8772), .A2(n8760), .ZN(n8997) );
  NAND2_X1 U8982 ( .A1(n8764), .A2(n7397), .ZN(n7317) );
  NAND2_X1 U8983 ( .A1(n7317), .A2(n8772), .ZN(n8900) );
  INV_X1 U8984 ( .A(n9730), .ZN(n8775) );
  NOR2_X1 U8985 ( .A1(n7313), .A2(n8775), .ZN(n7318) );
  NAND2_X1 U8986 ( .A1(n9731), .A2(n7318), .ZN(n9728) );
  NAND2_X1 U8987 ( .A1(n9728), .A2(n8774), .ZN(n7319) );
  XOR2_X1 U8988 ( .A(n8966), .B(n7319), .Z(n7320) );
  OAI222_X1 U8989 ( .A1(n9735), .A2(n9598), .B1(n9757), .B2(n7348), .C1(n9862), 
        .C2(n7320), .ZN(n9877) );
  NAND2_X1 U8990 ( .A1(n9877), .A2(n9222), .ZN(n7329) );
  NAND2_X1 U8991 ( .A1(n9744), .A2(n9879), .ZN(n7323) );
  NAND2_X1 U8992 ( .A1(n7323), .A2(n9785), .ZN(n7324) );
  NOR2_X1 U8993 ( .A1(n7365), .A2(n7324), .ZN(n9878) );
  NOR2_X1 U8994 ( .A1(n9781), .A2(n4761), .ZN(n7327) );
  INV_X1 U8995 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7325) );
  OAI22_X1 U8996 ( .A1(n9222), .A2(n7325), .B1(n7349), .B2(n9319), .ZN(n7326)
         );
  AOI211_X1 U8997 ( .C1(n9878), .C2(n9787), .A(n7327), .B(n7326), .ZN(n7328)
         );
  OAI211_X1 U8998 ( .C1(n9331), .C2(n9882), .A(n7329), .B(n7328), .ZN(P1_U3282) );
  OAI222_X1 U8999 ( .A1(n7729), .A2(n7331), .B1(P2_U3152), .B2(n7828), .C1(
        n8612), .C2(n7330), .ZN(P2_U3337) );
  INV_X1 U9000 ( .A(n9731), .ZN(n7332) );
  AOI21_X1 U9001 ( .B1(n8961), .B2(n7333), .A(n7332), .ZN(n9863) );
  NOR2_X1 U9002 ( .A1(n9779), .A2(n9862), .ZN(n9329) );
  INV_X1 U9003 ( .A(n9329), .ZN(n9310) );
  OR2_X1 U9004 ( .A1(n9807), .A2(n9735), .ZN(n9203) );
  OR2_X1 U9005 ( .A1(n9807), .A2(n9757), .ZN(n9318) );
  INV_X1 U9006 ( .A(n9318), .ZN(n7409) );
  NAND2_X1 U9007 ( .A1(n7409), .A2(n9855), .ZN(n7337) );
  INV_X1 U9008 ( .A(n7334), .ZN(n7335) );
  AOI22_X1 U9009 ( .A1(n9779), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7335), .B2(
        n9804), .ZN(n7336) );
  OAI211_X1 U9010 ( .C1(n7348), .C2(n9203), .A(n7337), .B(n7336), .ZN(n7339)
         );
  OAI211_X1 U9011 ( .C1(n7404), .C2(n9861), .A(n9743), .B(n9785), .ZN(n9860)
         );
  NOR2_X1 U9012 ( .A1(n9860), .A2(n9576), .ZN(n7338) );
  AOI211_X1 U9013 ( .C1(n9572), .C2(n7340), .A(n7339), .B(n7338), .ZN(n7343)
         );
  XNOR2_X1 U9014 ( .A(n7341), .B(n8961), .ZN(n9866) );
  NAND2_X1 U9015 ( .A1(n9866), .A2(n9767), .ZN(n7342) );
  OAI211_X1 U9016 ( .C1(n9863), .C2(n9310), .A(n7343), .B(n7342), .ZN(P1_U3284) );
  INV_X1 U9017 ( .A(n7345), .ZN(n7346) );
  AOI21_X1 U9018 ( .B1(n7347), .B2(n7344), .A(n7346), .ZN(n7353) );
  INV_X1 U9019 ( .A(n9598), .ZN(n7468) );
  AND2_X1 U9020 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9671) );
  OAI22_X1 U9021 ( .A1(n8736), .A2(n7349), .B1(n8723), .B2(n7348), .ZN(n7350)
         );
  AOI211_X1 U9022 ( .C1(n8725), .C2(n7468), .A(n9671), .B(n7350), .ZN(n7352)
         );
  NAND2_X1 U9023 ( .A1(n9879), .A2(n8710), .ZN(n7351) );
  OAI211_X1 U9024 ( .C1(n7353), .C2(n8712), .A(n7352), .B(n7351), .ZN(P1_U3229) );
  AND2_X1 U9025 ( .A1(n8780), .A2(n8774), .ZN(n8767) );
  NAND2_X1 U9026 ( .A1(n9728), .A2(n8767), .ZN(n7355) );
  NAND2_X1 U9027 ( .A1(n7355), .A2(n8777), .ZN(n7354) );
  OR2_X1 U9028 ( .A1(n7469), .A2(n9598), .ZN(n8769) );
  NAND2_X1 U9029 ( .A1(n7469), .A2(n9598), .ZN(n8782) );
  NAND2_X1 U9030 ( .A1(n8769), .A2(n8782), .ZN(n8967) );
  AOI21_X1 U9031 ( .B1(n7354), .B2(n8967), .A(n9862), .ZN(n7357) );
  AND2_X1 U9032 ( .A1(n8782), .A2(n8777), .ZN(n8905) );
  NAND2_X1 U9033 ( .A1(n7355), .A2(n8905), .ZN(n7478) );
  INV_X1 U9034 ( .A(n8769), .ZN(n8903) );
  OR2_X1 U9035 ( .A1(n7478), .A2(n8903), .ZN(n7356) );
  NAND2_X1 U9036 ( .A1(n7357), .A2(n7356), .ZN(n7496) );
  OR2_X1 U9037 ( .A1(n9879), .A2(n9034), .ZN(n7359) );
  AND2_X1 U9038 ( .A1(n9879), .A2(n9034), .ZN(n7358) );
  NAND2_X1 U9039 ( .A1(n7361), .A2(n8967), .ZN(n7471) );
  OAI21_X1 U9040 ( .B1(n7361), .B2(n8967), .A(n7471), .ZN(n7498) );
  NAND2_X1 U9041 ( .A1(n7498), .A2(n9767), .ZN(n7369) );
  INV_X1 U9042 ( .A(n9033), .ZN(n9569) );
  OAI22_X1 U9043 ( .A1(n9222), .A2(n7362), .B1(n7442), .B2(n9319), .ZN(n7363)
         );
  AOI21_X1 U9044 ( .B1(n7409), .B2(n9034), .A(n7363), .ZN(n7364) );
  OAI21_X1 U9045 ( .B1(n9569), .B2(n9203), .A(n7364), .ZN(n7367) );
  INV_X1 U9046 ( .A(n7469), .ZN(n7505) );
  OAI211_X1 U9047 ( .C1(n7505), .C2(n7365), .A(n4558), .B(n9785), .ZN(n7494)
         );
  NOR2_X1 U9048 ( .A1(n7494), .A2(n9576), .ZN(n7366) );
  AOI211_X1 U9049 ( .C1(n9572), .C2(n7469), .A(n7367), .B(n7366), .ZN(n7368)
         );
  OAI211_X1 U9050 ( .C1(n9807), .C2(n7496), .A(n7369), .B(n7368), .ZN(P1_U3281) );
  AND2_X1 U9051 ( .A1(n7424), .A2(n7449), .ZN(n7416) );
  INV_X1 U9052 ( .A(n7416), .ZN(n7909) );
  XOR2_X1 U9053 ( .A(n7417), .B(n8007), .Z(n7371) );
  OAI222_X1 U9054 ( .A1(n8428), .A2(n7554), .B1(n8426), .B2(n7392), .C1(n7371), 
        .C2(n8425), .ZN(n10038) );
  INV_X1 U9055 ( .A(n10038), .ZN(n7385) );
  INV_X1 U9056 ( .A(n7392), .ZN(n8157) );
  NAND2_X1 U9057 ( .A1(n7372), .A2(n8157), .ZN(n7373) );
  INV_X1 U9058 ( .A(n7375), .ZN(n7376) );
  OAI21_X1 U9059 ( .B1(n7376), .B2(n4926), .A(n7426), .ZN(n10040) );
  INV_X1 U9060 ( .A(n7424), .ZN(n10035) );
  OR2_X1 U9061 ( .A1(n7378), .A2(n10035), .ZN(n7379) );
  NAND2_X1 U9062 ( .A1(n7420), .A2(n7379), .ZN(n10037) );
  INV_X1 U9063 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7380) );
  OAI22_X1 U9064 ( .A1(n9927), .A2(n7380), .B1(n7391), .B2(n9924), .ZN(n7381)
         );
  AOI21_X1 U9065 ( .B1(n7424), .B2(n8490), .A(n7381), .ZN(n7382) );
  OAI21_X1 U9066 ( .B1(n10037), .B2(n9948), .A(n7382), .ZN(n7383) );
  AOI21_X1 U9067 ( .B1(n10040), .B2(n9944), .A(n7383), .ZN(n7384) );
  OAI21_X1 U9068 ( .B1(n7385), .B2(n9941), .A(n7384), .ZN(P2_U3284) );
  INV_X1 U9069 ( .A(n7386), .ZN(n7387) );
  AOI21_X1 U9070 ( .B1(n7389), .B2(n7388), .A(n7387), .ZN(n7396) );
  OAI21_X1 U9071 ( .B1(n8128), .B2(n7391), .A(n7390), .ZN(n7394) );
  OAI22_X1 U9072 ( .A1(n8131), .A2(n7554), .B1(n7392), .B2(n8129), .ZN(n7393)
         );
  AOI211_X1 U9073 ( .C1(n8143), .C2(n7424), .A(n7394), .B(n7393), .ZN(n7395)
         );
  OAI21_X1 U9074 ( .B1(n7396), .B2(n8145), .A(n7395), .ZN(P2_U3226) );
  NAND2_X1 U9075 ( .A1(n8896), .A2(n7397), .ZN(n8996) );
  INV_X1 U9076 ( .A(n8996), .ZN(n7398) );
  NAND2_X1 U9077 ( .A1(n7399), .A2(n7398), .ZN(n8763) );
  NAND2_X1 U9078 ( .A1(n8763), .A2(n8760), .ZN(n7400) );
  INV_X1 U9079 ( .A(n8757), .ZN(n8963) );
  XNOR2_X1 U9080 ( .A(n7400), .B(n8963), .ZN(n7401) );
  NAND2_X1 U9081 ( .A1(n7401), .A2(n9427), .ZN(n9848) );
  OAI21_X1 U9082 ( .B1(n7403), .B2(n8757), .A(n7402), .ZN(n9853) );
  INV_X1 U9083 ( .A(n7404), .ZN(n7406) );
  AOI21_X1 U9084 ( .B1(n9751), .B2(n7412), .A(n9749), .ZN(n7405) );
  NAND2_X1 U9085 ( .A1(n7406), .A2(n7405), .ZN(n9846) );
  INV_X1 U9086 ( .A(n9843), .ZN(n9734) );
  OAI22_X1 U9087 ( .A1(n9222), .A2(n6744), .B1(n7407), .B2(n9319), .ZN(n7408)
         );
  AOI21_X1 U9088 ( .B1(n7409), .B2(n9844), .A(n7408), .ZN(n7410) );
  OAI21_X1 U9089 ( .B1(n9734), .B2(n9203), .A(n7410), .ZN(n7411) );
  AOI21_X1 U9090 ( .B1(n9572), .B2(n7412), .A(n7411), .ZN(n7413) );
  OAI21_X1 U9091 ( .B1(n9576), .B2(n9846), .A(n7413), .ZN(n7414) );
  AOI21_X1 U9092 ( .B1(n9853), .B2(n9767), .A(n7414), .ZN(n7415) );
  OAI21_X1 U9093 ( .B1(n9807), .B2(n9848), .A(n7415), .ZN(P1_U3285) );
  OR2_X1 U9094 ( .A1(n7534), .A2(n7554), .ZN(n7919) );
  NAND2_X1 U9095 ( .A1(n7534), .A2(n7554), .ZN(n7530) );
  NAND2_X1 U9096 ( .A1(n7919), .A2(n7530), .ZN(n7528) );
  XNOR2_X1 U9097 ( .A(n7529), .B(n8008), .ZN(n7418) );
  OAI222_X1 U9098 ( .A1(n8428), .A2(n7642), .B1(n8426), .B2(n7449), .C1(n8425), 
        .C2(n7418), .ZN(n9550) );
  INV_X1 U9099 ( .A(n9550), .ZN(n7432) );
  OAI22_X1 U9100 ( .A1(n9927), .A2(n7419), .B1(n7448), .B2(n9924), .ZN(n7423)
         );
  INV_X1 U9101 ( .A(n7420), .ZN(n7421) );
  INV_X1 U9102 ( .A(n7534), .ZN(n9548) );
  OAI21_X1 U9103 ( .B1(n7421), .B2(n9548), .A(n7568), .ZN(n9549) );
  NOR2_X1 U9104 ( .A1(n9549), .A2(n9948), .ZN(n7422) );
  AOI211_X1 U9105 ( .C1(n8490), .C2(n7534), .A(n7423), .B(n7422), .ZN(n7431)
         );
  INV_X1 U9106 ( .A(n7449), .ZN(n8156) );
  OR2_X1 U9107 ( .A1(n7424), .A2(n8156), .ZN(n7425) );
  AND2_X1 U9108 ( .A1(n7427), .A2(n8008), .ZN(n9547) );
  INV_X1 U9109 ( .A(n9547), .ZN(n7429) );
  INV_X1 U9110 ( .A(n7427), .ZN(n7428) );
  NAND3_X1 U9111 ( .A1(n7429), .A2(n9944), .A3(n9552), .ZN(n7430) );
  OAI211_X1 U9112 ( .C1(n7432), .C2(n9941), .A(n7431), .B(n7430), .ZN(P2_U3283) );
  INV_X1 U9113 ( .A(n7433), .ZN(n7801) );
  OAI222_X1 U9114 ( .A1(n7622), .A2(n10434), .B1(n8036), .B2(n7801), .C1(
        P1_U3084), .C2(n7434), .ZN(P1_U3331) );
  INV_X1 U9115 ( .A(n7435), .ZN(n7437) );
  NOR2_X1 U9116 ( .A1(n7437), .A2(n7436), .ZN(n7438) );
  XNOR2_X1 U9117 ( .A(n7439), .B(n7438), .ZN(n7440) );
  NAND2_X1 U9118 ( .A1(n7440), .A2(n8732), .ZN(n7445) );
  NOR2_X1 U9119 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7441), .ZN(n9687) );
  OAI22_X1 U9120 ( .A1(n8736), .A2(n7442), .B1(n8723), .B2(n9736), .ZN(n7443)
         );
  AOI211_X1 U9121 ( .C1(n8725), .C2(n9033), .A(n9687), .B(n7443), .ZN(n7444)
         );
  OAI211_X1 U9122 ( .C1(n7505), .C2(n8743), .A(n7445), .B(n7444), .ZN(P1_U3215) );
  XNOR2_X1 U9123 ( .A(n7447), .B(n7446), .ZN(n7453) );
  OAI22_X1 U9124 ( .A1(n8128), .A2(n7448), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5428), .ZN(n7451) );
  OAI22_X1 U9125 ( .A1(n8131), .A2(n7642), .B1(n7449), .B2(n8129), .ZN(n7450)
         );
  AOI211_X1 U9126 ( .C1(n8143), .C2(n7534), .A(n7451), .B(n7450), .ZN(n7452)
         );
  OAI21_X1 U9127 ( .B1(n7453), .B2(n8145), .A(n7452), .ZN(P2_U3236) );
  AOI22_X1 U9128 ( .A1(n8174), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7537), .B2(
        n7464), .ZN(n7456) );
  NAND2_X1 U9129 ( .A1(n7456), .A2(n7455), .ZN(n8168) );
  OAI21_X1 U9130 ( .B1(n7456), .B2(n7455), .A(n8168), .ZN(n7466) );
  AOI22_X1 U9131 ( .A1(n8174), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n5453), .B2(
        n7464), .ZN(n7460) );
  OAI21_X1 U9132 ( .B1(n7458), .B2(P2_REG1_REG_13__SCAN_IN), .A(n7457), .ZN(
        n7459) );
  NAND2_X1 U9133 ( .A1(n7460), .A2(n7459), .ZN(n8173) );
  OAI21_X1 U9134 ( .B1(n7460), .B2(n7459), .A(n8173), .ZN(n7461) );
  NAND2_X1 U9135 ( .A1(n7461), .A2(n9904), .ZN(n7463) );
  NOR2_X1 U9136 ( .A1(n10442), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7556) );
  AOI21_X1 U9137 ( .B1(n9909), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n7556), .ZN(
        n7462) );
  OAI211_X1 U9138 ( .C1(n9906), .C2(n7464), .A(n7463), .B(n7462), .ZN(n7465)
         );
  AOI21_X1 U9139 ( .B1(n9903), .B2(n7466), .A(n7465), .ZN(n7467) );
  INV_X1 U9140 ( .A(n7467), .ZN(P2_U3259) );
  OR2_X1 U9141 ( .A1(n7469), .A2(n7468), .ZN(n7470) );
  NAND2_X1 U9142 ( .A1(n7471), .A2(n7470), .ZN(n7605) );
  NOR2_X1 U9143 ( .A1(n9601), .A2(n9033), .ZN(n7603) );
  NAND2_X1 U9144 ( .A1(n9601), .A2(n9033), .ZN(n7604) );
  INV_X1 U9145 ( .A(n7604), .ZN(n7472) );
  OR2_X1 U9146 ( .A1(n7603), .A2(n7472), .ZN(n8969) );
  XOR2_X1 U9147 ( .A(n7605), .B(n8969), .Z(n9606) );
  INV_X1 U9148 ( .A(n9606), .ZN(n9604) );
  INV_X1 U9149 ( .A(n9601), .ZN(n7527) );
  INV_X1 U9150 ( .A(n9573), .ZN(n7473) );
  AOI211_X1 U9151 ( .C1(n9601), .C2(n4558), .A(n9749), .B(n7473), .ZN(n9599)
         );
  INV_X1 U9152 ( .A(n9203), .ZN(n9325) );
  INV_X1 U9153 ( .A(n9597), .ZN(n7607) );
  NOR2_X1 U9154 ( .A1(n9318), .A2(n9598), .ZN(n7476) );
  OAI22_X1 U9155 ( .A1(n9222), .A2(n7474), .B1(n7523), .B2(n9319), .ZN(n7475)
         );
  AOI211_X1 U9156 ( .C1(n9325), .C2(n7607), .A(n7476), .B(n7475), .ZN(n7477)
         );
  OAI21_X1 U9157 ( .B1(n7527), .B2(n9781), .A(n7477), .ZN(n7482) );
  NAND2_X1 U9158 ( .A1(n7478), .A2(n8769), .ZN(n7596) );
  INV_X1 U9159 ( .A(n8969), .ZN(n7479) );
  XNOR2_X1 U9160 ( .A(n7596), .B(n7479), .ZN(n7480) );
  NAND2_X1 U9161 ( .A1(n7480), .A2(n9427), .ZN(n9602) );
  NOR2_X1 U9162 ( .A1(n9602), .A2(n9779), .ZN(n7481) );
  AOI211_X1 U9163 ( .C1(n9599), .C2(n9787), .A(n7482), .B(n7481), .ZN(n7483)
         );
  OAI21_X1 U9164 ( .B1(n9604), .B2(n9331), .A(n7483), .ZN(P1_U3280) );
  NAND2_X1 U9165 ( .A1(n7486), .A2(n8604), .ZN(n7484) );
  OAI211_X1 U9166 ( .C1(n7485), .C2(n7729), .A(n7484), .B(n8033), .ZN(P2_U3335) );
  NAND2_X1 U9167 ( .A1(n7486), .A2(n9502), .ZN(n7488) );
  OR2_X1 U9168 ( .A1(n7487), .A2(P1_U3084), .ZN(n9027) );
  OAI211_X1 U9169 ( .C1(n10465), .C2(n9499), .A(n7488), .B(n9027), .ZN(
        P1_U3330) );
  AND2_X1 U9170 ( .A1(n7490), .A2(n7489), .ZN(n7491) );
  AND3_X1 U9171 ( .A1(n7492), .A2(n9810), .A3(n7491), .ZN(n7501) );
  AND2_X2 U9172 ( .A1(n7501), .A2(n7493), .ZN(n9902) );
  INV_X1 U9173 ( .A(n9869), .ZN(n9880) );
  AND2_X1 U9174 ( .A1(n9902), .A2(n9880), .ZN(n9351) );
  INV_X1 U9175 ( .A(n9875), .ZN(n9883) );
  NAND2_X1 U9176 ( .A1(n9849), .A2(n9883), .ZN(n9867) );
  AOI22_X1 U9177 ( .A1(n9856), .A2(n9034), .B1(n9033), .B2(n9857), .ZN(n7495)
         );
  NAND3_X1 U9178 ( .A1(n7496), .A2(n7495), .A3(n7494), .ZN(n7497) );
  AOI21_X1 U9179 ( .B1(n7498), .B2(n9867), .A(n7497), .ZN(n7502) );
  MUX2_X1 U9180 ( .A(n6111), .B(n7502), .S(n9902), .Z(n7499) );
  OAI21_X1 U9181 ( .B1(n7505), .B2(n9434), .A(n7499), .ZN(P1_U3533) );
  AND2_X2 U9182 ( .A1(n7501), .A2(n7500), .ZN(n9888) );
  NAND2_X1 U9183 ( .A1(n9888), .A2(n9880), .ZN(n9494) );
  INV_X1 U9184 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7503) );
  MUX2_X1 U9185 ( .A(n7503), .B(n7502), .S(n9888), .Z(n7504) );
  OAI21_X1 U9186 ( .B1(n7505), .B2(n9494), .A(n7504), .ZN(P1_U3484) );
  NAND2_X1 U9187 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8734) );
  XNOR2_X1 U9188 ( .A(n7739), .B(n7738), .ZN(n7508) );
  INV_X1 U9189 ( .A(n7508), .ZN(n7511) );
  NOR2_X1 U9190 ( .A1(n7509), .A2(n7508), .ZN(n7740) );
  INV_X1 U9191 ( .A(n7740), .ZN(n7510) );
  OAI211_X1 U9192 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n7511), .A(n9720), .B(
        n7510), .ZN(n7512) );
  OAI211_X1 U9193 ( .C1(n9715), .C2(n7739), .A(n8734), .B(n7512), .ZN(n7518)
         );
  XNOR2_X1 U9194 ( .A(n7730), .B(n7739), .ZN(n7516) );
  NOR2_X1 U9195 ( .A1(n7677), .A2(n7516), .ZN(n7731) );
  AOI211_X1 U9196 ( .C1(n7516), .C2(n7677), .A(n7731), .B(n9682), .ZN(n7517)
         );
  AOI211_X1 U9197 ( .C1(n9690), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n7518), .B(
        n7517), .ZN(n7519) );
  INV_X1 U9198 ( .A(n7519), .ZN(P1_U3256) );
  OAI211_X1 U9199 ( .C1(n7522), .C2(n7521), .A(n7520), .B(n8732), .ZN(n7526)
         );
  AND2_X1 U9200 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9693) );
  OAI22_X1 U9201 ( .A1(n8736), .A2(n7523), .B1(n8723), .B2(n9598), .ZN(n7524)
         );
  AOI211_X1 U9202 ( .C1(n8725), .C2(n7607), .A(n9693), .B(n7524), .ZN(n7525)
         );
  OAI211_X1 U9203 ( .C1(n7527), .C2(n8743), .A(n7526), .B(n7525), .ZN(P1_U3234) );
  NAND2_X1 U9204 ( .A1(n7567), .A2(n7642), .ZN(n7917) );
  INV_X1 U9205 ( .A(n7530), .ZN(n7914) );
  NAND2_X1 U9206 ( .A1(n7531), .A2(n8009), .ZN(n7561) );
  OAI211_X1 U9207 ( .C1(n8009), .C2(n7531), .A(n7561), .B(n9938), .ZN(n7533)
         );
  INV_X1 U9208 ( .A(n8093), .ZN(n8153) );
  INV_X1 U9209 ( .A(n7554), .ZN(n8155) );
  AOI22_X1 U9210 ( .A1(n8153), .A2(n9917), .B1(n8155), .B2(n9915), .ZN(n7532)
         );
  NAND2_X1 U9211 ( .A1(n7533), .A2(n7532), .ZN(n9544) );
  INV_X1 U9212 ( .A(n9544), .ZN(n7542) );
  NAND2_X1 U9213 ( .A1(n7534), .A2(n8155), .ZN(n7535) );
  OAI21_X1 U9214 ( .B1(n7536), .B2(n7921), .A(n7560), .ZN(n9546) );
  XNOR2_X1 U9215 ( .A(n7568), .B(n7567), .ZN(n9543) );
  OAI22_X1 U9216 ( .A1(n9927), .A2(n7537), .B1(n7553), .B2(n9924), .ZN(n7538)
         );
  AOI21_X1 U9217 ( .B1(n7567), .B2(n8490), .A(n7538), .ZN(n7539) );
  OAI21_X1 U9218 ( .B1(n9543), .B2(n9948), .A(n7539), .ZN(n7540) );
  AOI21_X1 U9219 ( .B1(n9546), .B2(n9944), .A(n7540), .ZN(n7541) );
  OAI21_X1 U9220 ( .B1(n7542), .B2(n9941), .A(n7541), .ZN(P2_U3282) );
  INV_X1 U9221 ( .A(n7543), .ZN(n7547) );
  OAI222_X1 U9222 ( .A1(P1_U3084), .A2(n7544), .B1(n8036), .B2(n7547), .C1(
        n10368), .C2(n7622), .ZN(P1_U3329) );
  INV_X1 U9223 ( .A(n7545), .ZN(n7548) );
  OAI222_X1 U9224 ( .A1(P2_U3152), .A2(n7548), .B1(n8612), .B2(n7547), .C1(
        n7546), .C2(n7729), .ZN(P2_U3334) );
  OAI21_X1 U9225 ( .B1(n7551), .B2(n7550), .A(n7549), .ZN(n7552) );
  NAND2_X1 U9226 ( .A1(n7552), .A2(n8117), .ZN(n7559) );
  INV_X1 U9227 ( .A(n7553), .ZN(n7557) );
  OAI22_X1 U9228 ( .A1(n8131), .A2(n8093), .B1(n7554), .B2(n8129), .ZN(n7555)
         );
  AOI211_X1 U9229 ( .C1(n8138), .C2(n7557), .A(n7556), .B(n7555), .ZN(n7558)
         );
  OAI211_X1 U9230 ( .C1(n4880), .C2(n8123), .A(n7559), .B(n7558), .ZN(P2_U3217) );
  NAND2_X1 U9231 ( .A1(n7658), .A2(n8093), .ZN(n7923) );
  XNOR2_X1 U9232 ( .A(n7657), .B(n5004), .ZN(n9542) );
  INV_X1 U9233 ( .A(n9542), .ZN(n7576) );
  NAND3_X1 U9234 ( .A1(n7561), .A2(n5004), .A3(n7915), .ZN(n7564) );
  NAND3_X1 U9235 ( .A1(n7649), .A2(n9938), .A3(n7564), .ZN(n7566) );
  INV_X1 U9236 ( .A(n7650), .ZN(n8260) );
  AOI22_X1 U9237 ( .A1(n8260), .A2(n9917), .B1(n9915), .B2(n8154), .ZN(n7565)
         );
  NAND2_X1 U9238 ( .A1(n7566), .A2(n7565), .ZN(n9540) );
  INV_X1 U9239 ( .A(n7658), .ZN(n9538) );
  NOR2_X1 U9240 ( .A1(n7569), .A2(n9538), .ZN(n7570) );
  OR2_X1 U9241 ( .A1(n7653), .A2(n7570), .ZN(n9539) );
  OAI22_X1 U9242 ( .A1(n9927), .A2(n7571), .B1(n7641), .B2(n9924), .ZN(n7572)
         );
  AOI21_X1 U9243 ( .B1(n7658), .B2(n8490), .A(n7572), .ZN(n7573) );
  OAI21_X1 U9244 ( .B1(n9539), .B2(n9948), .A(n7573), .ZN(n7574) );
  AOI21_X1 U9245 ( .B1(n9540), .B2(n9927), .A(n7574), .ZN(n7575) );
  OAI21_X1 U9246 ( .B1(n7576), .B2(n8478), .A(n7575), .ZN(P2_U3281) );
  INV_X1 U9247 ( .A(n7577), .ZN(n7578) );
  AOI21_X1 U9248 ( .B1(n7580), .B2(n7579), .A(n7578), .ZN(n7585) );
  INV_X1 U9249 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7581) );
  OAI22_X1 U9250 ( .A1(n8735), .A2(n9568), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7581), .ZN(n7583) );
  OAI22_X1 U9251 ( .A1(n8736), .A2(n9570), .B1(n8723), .B2(n9569), .ZN(n7582)
         );
  AOI211_X1 U9252 ( .C1(n9592), .C2(n8710), .A(n7583), .B(n7582), .ZN(n7584)
         );
  OAI21_X1 U9253 ( .B1(n7585), .B2(n8712), .A(n7584), .ZN(P1_U3222) );
  INV_X1 U9254 ( .A(n9586), .ZN(n7762) );
  XNOR2_X1 U9255 ( .A(n7587), .B(n7586), .ZN(n7588) );
  XNOR2_X1 U9256 ( .A(n7589), .B(n7588), .ZN(n7590) );
  NAND2_X1 U9257 ( .A1(n7590), .A2(n8732), .ZN(n7595) );
  INV_X1 U9258 ( .A(n7591), .ZN(n7593) );
  OAI22_X1 U9259 ( .A1(n8736), .A2(n7757), .B1(n8723), .B2(n9597), .ZN(n7592)
         );
  AOI211_X1 U9260 ( .C1(n8725), .C2(n9441), .A(n7593), .B(n7592), .ZN(n7594)
         );
  OAI211_X1 U9261 ( .C1(n7762), .C2(n8743), .A(n7595), .B(n7594), .ZN(P1_U3232) );
  NAND2_X1 U9262 ( .A1(n9601), .A2(n9569), .ZN(n8795) );
  NAND2_X1 U9263 ( .A1(n7596), .A2(n8795), .ZN(n9565) );
  OR2_X1 U9264 ( .A1(n9592), .A2(n9597), .ZN(n8798) );
  OR2_X1 U9265 ( .A1(n9601), .A2(n9569), .ZN(n9564) );
  AND2_X1 U9266 ( .A1(n8798), .A2(n9564), .ZN(n8908) );
  NAND2_X1 U9267 ( .A1(n9565), .A2(n8908), .ZN(n7597) );
  NAND2_X1 U9268 ( .A1(n9592), .A2(n9597), .ZN(n8796) );
  NAND2_X1 U9269 ( .A1(n7597), .A2(n8796), .ZN(n7763) );
  OR2_X1 U9270 ( .A1(n9586), .A2(n9568), .ZN(n8906) );
  NAND2_X1 U9271 ( .A1(n9586), .A2(n9568), .ZN(n8909) );
  NAND2_X1 U9272 ( .A1(n7763), .A2(n8971), .ZN(n7765) );
  OR2_X1 U9273 ( .A1(n7672), .A2(n9583), .ZN(n8911) );
  NAND2_X1 U9274 ( .A1(n7672), .A2(n9583), .ZN(n8916) );
  NAND2_X1 U9275 ( .A1(n8911), .A2(n8916), .ZN(n8973) );
  INV_X1 U9276 ( .A(n8909), .ZN(n7598) );
  NOR2_X1 U9277 ( .A1(n8973), .A2(n7598), .ZN(n7599) );
  NAND2_X1 U9278 ( .A1(n7673), .A2(n9427), .ZN(n7602) );
  INV_X1 U9279 ( .A(n8973), .ZN(n8784) );
  AOI21_X1 U9280 ( .B1(n7765), .B2(n8909), .A(n8784), .ZN(n7601) );
  AOI22_X1 U9281 ( .A1(n9856), .A2(n9032), .B1(n9031), .B2(n9857), .ZN(n7600)
         );
  OAI21_X1 U9282 ( .B1(n7602), .B2(n7601), .A(n7600), .ZN(n7664) );
  INV_X1 U9283 ( .A(n7664), .ZN(n7616) );
  NAND2_X1 U9284 ( .A1(n8798), .A2(n8796), .ZN(n9560) );
  NOR2_X1 U9285 ( .A1(n9586), .A2(n9032), .ZN(n7609) );
  XNOR2_X1 U9286 ( .A(n7671), .B(n8784), .ZN(n7666) );
  NAND2_X1 U9287 ( .A1(n7666), .A2(n9767), .ZN(n7615) );
  INV_X1 U9288 ( .A(n7756), .ZN(n7610) );
  AOI211_X1 U9289 ( .C1(n7672), .C2(n7610), .A(n9749), .B(n7676), .ZN(n7665)
         );
  NOR2_X1 U9290 ( .A1(n8788), .A2(n9781), .ZN(n7613) );
  OAI22_X1 U9291 ( .A1(n9222), .A2(n7611), .B1(n7690), .B2(n9319), .ZN(n7612)
         );
  AOI211_X1 U9292 ( .C1(n7665), .C2(n9787), .A(n7613), .B(n7612), .ZN(n7614)
         );
  OAI211_X1 U9293 ( .C1(n9807), .C2(n7616), .A(n7615), .B(n7614), .ZN(P1_U3277) );
  INV_X1 U9294 ( .A(n7617), .ZN(n7621) );
  OAI222_X1 U9295 ( .A1(n7729), .A2(n7619), .B1(n8612), .B2(n7621), .C1(
        P2_U3152), .C2(n7618), .ZN(P2_U3333) );
  OAI222_X1 U9296 ( .A1(n7622), .A2(n10437), .B1(n8036), .B2(n7621), .C1(
        P1_U3084), .C2(n7620), .ZN(P1_U3328) );
  XNOR2_X1 U9297 ( .A(n7624), .B(n7623), .ZN(n7630) );
  INV_X1 U9298 ( .A(n8141), .ZN(n8066) );
  OR2_X1 U9299 ( .A1(n8152), .A2(n8428), .ZN(n7626) );
  OR2_X1 U9300 ( .A1(n7650), .A2(n8426), .ZN(n7625) );
  NAND2_X1 U9301 ( .A1(n7626), .A2(n7625), .ZN(n8480) );
  AOI22_X1 U9302 ( .A1(n8066), .A2(n8480), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3152), .ZN(n7627) );
  OAI21_X1 U9303 ( .B1(n8488), .B2(n8128), .A(n7627), .ZN(n7628) );
  AOI21_X1 U9304 ( .B1(n8571), .B2(n8143), .A(n7628), .ZN(n7629) );
  OAI21_X1 U9305 ( .B1(n7630), .B2(n8145), .A(n7629), .ZN(P2_U3230) );
  INV_X1 U9306 ( .A(n7631), .ZN(n7634) );
  OAI222_X1 U9307 ( .A1(P2_U3152), .A2(n7633), .B1(n8612), .B2(n7634), .C1(
        n7632), .C2(n7729), .ZN(P2_U3332) );
  OAI222_X1 U9308 ( .A1(P1_U3084), .A2(n7635), .B1(n8036), .B2(n7634), .C1(
        n10449), .C2(n9499), .ZN(P1_U3327) );
  NAND2_X1 U9309 ( .A1(n7638), .A2(n7637), .ZN(n8086) );
  OAI21_X1 U9310 ( .B1(n7638), .B2(n7637), .A(n8086), .ZN(n7639) );
  NOR2_X1 U9311 ( .A1(n7639), .A2(n7640), .ZN(n8089) );
  AOI21_X1 U9312 ( .B1(n7640), .B2(n7639), .A(n8089), .ZN(n7646) );
  NAND2_X1 U9313 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n8170) );
  OAI21_X1 U9314 ( .B1(n8128), .B2(n7641), .A(n8170), .ZN(n7644) );
  OAI22_X1 U9315 ( .A1(n8131), .A2(n7650), .B1(n7642), .B2(n8129), .ZN(n7643)
         );
  AOI211_X1 U9316 ( .C1(n7658), .C2(n8143), .A(n7644), .B(n7643), .ZN(n7645)
         );
  OAI21_X1 U9317 ( .B1(n7646), .B2(n8145), .A(n7645), .ZN(P2_U3243) );
  NAND2_X1 U9318 ( .A1(n7726), .A2(n9502), .ZN(n7648) );
  OAI211_X1 U9319 ( .C1(n9499), .C2(n10272), .A(n7648), .B(n7647), .ZN(
        P1_U3326) );
  OR2_X1 U9320 ( .A1(n8578), .A2(n7650), .ZN(n7930) );
  NAND2_X1 U9321 ( .A1(n8578), .A2(n7650), .ZN(n7929) );
  NAND2_X1 U9322 ( .A1(n7930), .A2(n7929), .ZN(n8011) );
  XNOR2_X1 U9323 ( .A(n7812), .B(n8011), .ZN(n7652) );
  OAI22_X1 U9324 ( .A1(n8130), .A2(n8428), .B1(n8093), .B2(n8426), .ZN(n7651)
         );
  AOI21_X1 U9325 ( .B1(n7652), .B2(n9938), .A(n7651), .ZN(n8581) );
  INV_X1 U9326 ( .A(n8578), .ZN(n8098) );
  NAND2_X1 U9327 ( .A1(n8098), .A2(n7653), .ZN(n8484) );
  INV_X1 U9328 ( .A(n7653), .ZN(n7654) );
  NAND2_X1 U9329 ( .A1(n7654), .A2(n8578), .ZN(n7655) );
  AND2_X1 U9330 ( .A1(n8484), .A2(n7655), .ZN(n8579) );
  INV_X1 U9331 ( .A(n9924), .ZN(n9940) );
  AOI22_X1 U9332 ( .A1(n9941), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8095), .B2(
        n9940), .ZN(n7656) );
  OAI21_X1 U9333 ( .B1(n8098), .B2(n9951), .A(n7656), .ZN(n7662) );
  NAND2_X1 U9334 ( .A1(n7657), .A2(n5004), .ZN(n7660) );
  OR2_X1 U9335 ( .A1(n7658), .A2(n8153), .ZN(n7659) );
  NAND2_X1 U9336 ( .A1(n7660), .A2(n7659), .ZN(n8263) );
  INV_X1 U9337 ( .A(n8011), .ZN(n8262) );
  XNOR2_X1 U9338 ( .A(n8263), .B(n8262), .ZN(n8582) );
  NOR2_X1 U9339 ( .A1(n8582), .A2(n8478), .ZN(n7661) );
  AOI211_X1 U9340 ( .C1(n8579), .C2(n8442), .A(n7662), .B(n7661), .ZN(n7663)
         );
  OAI21_X1 U9341 ( .B1(n9941), .B2(n8581), .A(n7663), .ZN(P2_U3280) );
  AOI211_X1 U9342 ( .C1(n7666), .C2(n9867), .A(n7665), .B(n7664), .ZN(n7668)
         );
  MUX2_X1 U9343 ( .A(n7221), .B(n7668), .S(n9902), .Z(n7667) );
  OAI21_X1 U9344 ( .B1(n8788), .B2(n9434), .A(n7667), .ZN(P1_U3537) );
  INV_X1 U9345 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n7669) );
  MUX2_X1 U9346 ( .A(n7669), .B(n7668), .S(n9888), .Z(n7670) );
  OAI21_X1 U9347 ( .B1(n8788), .B2(n9494), .A(n7670), .ZN(P1_U3496) );
  OR2_X1 U9348 ( .A1(n9443), .A2(n8652), .ZN(n8919) );
  NAND2_X1 U9349 ( .A1(n9443), .A2(n8652), .ZN(n8917) );
  NAND2_X1 U9350 ( .A1(n8919), .A2(n8917), .ZN(n8974) );
  INV_X1 U9351 ( .A(n8974), .ZN(n8808) );
  XNOR2_X1 U9352 ( .A(n7695), .B(n8808), .ZN(n9449) );
  INV_X1 U9353 ( .A(n9449), .ZN(n7684) );
  NAND2_X1 U9354 ( .A1(n7674), .A2(n8974), .ZN(n7675) );
  AOI21_X1 U9355 ( .B1(n7701), .B2(n7675), .A(n9862), .ZN(n9448) );
  OAI211_X1 U9356 ( .C1(n7676), .C2(n8744), .A(n9785), .B(n7697), .ZN(n9446)
         );
  INV_X1 U9357 ( .A(n9423), .ZN(n9442) );
  NOR2_X1 U9358 ( .A1(n9318), .A2(n9583), .ZN(n7679) );
  OAI22_X1 U9359 ( .A1(n9222), .A2(n7677), .B1(n8737), .B2(n9319), .ZN(n7678)
         );
  AOI211_X1 U9360 ( .C1(n9325), .C2(n9442), .A(n7679), .B(n7678), .ZN(n7681)
         );
  NAND2_X1 U9361 ( .A1(n9443), .A2(n9572), .ZN(n7680) );
  OAI211_X1 U9362 ( .C1(n9446), .C2(n9576), .A(n7681), .B(n7680), .ZN(n7682)
         );
  AOI21_X1 U9363 ( .B1(n9448), .B2(n9222), .A(n7682), .ZN(n7683) );
  OAI21_X1 U9364 ( .B1(n7684), .B2(n9331), .A(n7683), .ZN(P1_U3276) );
  XNOR2_X1 U9365 ( .A(n7686), .B(n7685), .ZN(n7687) );
  XNOR2_X1 U9366 ( .A(n7688), .B(n7687), .ZN(n7689) );
  NAND2_X1 U9367 ( .A1(n7689), .A2(n8732), .ZN(n7694) );
  OAI22_X1 U9368 ( .A1(n8736), .A2(n7690), .B1(n8735), .B2(n8652), .ZN(n7691)
         );
  AOI211_X1 U9369 ( .C1(n8740), .C2(n9032), .A(n7692), .B(n7691), .ZN(n7693)
         );
  OAI211_X1 U9370 ( .C1(n8788), .C2(n8743), .A(n7694), .B(n7693), .ZN(P1_U3213) );
  NAND2_X1 U9371 ( .A1(n9437), .A2(n9423), .ZN(n9077) );
  NAND2_X1 U9372 ( .A1(n9075), .A2(n9077), .ZN(n9103) );
  XNOR2_X1 U9373 ( .A(n9104), .B(n9103), .ZN(n9440) );
  INV_X1 U9374 ( .A(n9316), .ZN(n7696) );
  AOI211_X1 U9375 ( .C1(n9437), .C2(n7697), .A(n9749), .B(n7696), .ZN(n9436)
         );
  NOR2_X1 U9376 ( .A1(n4771), .A2(n9781), .ZN(n7700) );
  OAI22_X1 U9377 ( .A1(n9222), .A2(n7698), .B1(n8653), .B2(n9319), .ZN(n7699)
         );
  AOI211_X1 U9378 ( .C1(n9436), .C2(n9787), .A(n7700), .B(n7699), .ZN(n7704)
         );
  INV_X1 U9379 ( .A(n9414), .ZN(n9302) );
  XNOR2_X1 U9380 ( .A(n9076), .B(n9103), .ZN(n7702) );
  OAI222_X1 U9381 ( .A1(n9757), .A2(n8652), .B1(n9735), .B2(n9302), .C1(n7702), 
        .C2(n9862), .ZN(n9435) );
  NAND2_X1 U9382 ( .A1(n9435), .A2(n9222), .ZN(n7703) );
  OAI211_X1 U9383 ( .C1(n9440), .C2(n9331), .A(n7704), .B(n7703), .ZN(P1_U3275) );
  INV_X1 U9384 ( .A(n7770), .ZN(n8035) );
  INV_X1 U9385 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8854) );
  INV_X1 U9386 ( .A(n7708), .ZN(n7709) );
  INV_X1 U9387 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8609) );
  XNOR2_X1 U9388 ( .A(n7721), .B(SI_29_), .ZN(n7710) );
  INV_X1 U9389 ( .A(n8853), .ZN(n8611) );
  OAI222_X1 U9390 ( .A1(n9499), .A2(n8854), .B1(P1_U3084), .B2(n5869), .C1(
        n8036), .C2(n8611), .ZN(P1_U3324) );
  NAND2_X1 U9391 ( .A1(n7712), .A2(n7711), .ZN(n7713) );
  AOI21_X1 U9392 ( .B1(n7714), .B2(n7713), .A(n8145), .ZN(n7715) );
  AOI21_X1 U9393 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7809), .A(n7715), .ZN(
        n7719) );
  AOI22_X1 U9394 ( .A1(n7717), .A2(n8165), .B1(n8143), .B2(n7716), .ZN(n7718)
         );
  OAI211_X1 U9395 ( .C1(n7720), .C2(n8129), .A(n7719), .B(n7718), .ZN(P2_U3224) );
  INV_X1 U9396 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8747) );
  INV_X1 U9397 ( .A(n7721), .ZN(n7722) );
  NOR2_X1 U9398 ( .A1(n7722), .A2(SI_29_), .ZN(n7724) );
  NAND2_X1 U9399 ( .A1(n7722), .A2(SI_29_), .ZN(n7723) );
  MUX2_X1 U9400 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n7832), .Z(n7830) );
  INV_X1 U9401 ( .A(n8746), .ZN(n8607) );
  OAI222_X1 U9402 ( .A1(n9499), .A2(n8747), .B1(n8036), .B2(n8607), .C1(n5865), 
        .C2(P1_U3084), .ZN(P1_U3323) );
  INV_X1 U9403 ( .A(n7726), .ZN(n7727) );
  OAI222_X1 U9404 ( .A1(n7729), .A2(n7728), .B1(n8612), .B2(n7727), .C1(n8243), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  NOR2_X1 U9405 ( .A1(n7730), .A2(n7739), .ZN(n7732) );
  NAND2_X1 U9406 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n7742), .ZN(n7733) );
  OAI21_X1 U9407 ( .B1(n7742), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7733), .ZN(
        n9038) );
  NAND2_X1 U9408 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n7743), .ZN(n7734) );
  OAI21_X1 U9409 ( .B1(n7743), .B2(P1_REG2_REG_17__SCAN_IN), .A(n7734), .ZN(
        n9051) );
  AOI21_X1 U9410 ( .B1(n7743), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9050), .ZN(
        n9708) );
  OR2_X1 U9411 ( .A1(n7744), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7736) );
  NAND2_X1 U9412 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n7744), .ZN(n7735) );
  NAND2_X1 U9413 ( .A1(n7736), .A2(n7735), .ZN(n9709) );
  NOR2_X1 U9414 ( .A1(n9708), .A2(n9709), .ZN(n9707) );
  AOI21_X1 U9415 ( .B1(n7744), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9707), .ZN(
        n7737) );
  XNOR2_X1 U9416 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n7737), .ZN(n7750) );
  INV_X1 U9417 ( .A(n7750), .ZN(n7748) );
  AOI22_X1 U9418 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n7744), .B1(n9714), .B2(
        n9421), .ZN(n9718) );
  NOR2_X1 U9419 ( .A1(n7739), .A2(n7738), .ZN(n7741) );
  NOR2_X1 U9420 ( .A1(n7741), .A2(n7740), .ZN(n9042) );
  XNOR2_X1 U9421 ( .A(n7742), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9041) );
  NOR2_X1 U9422 ( .A1(n9042), .A2(n9041), .ZN(n9040) );
  AOI21_X1 U9423 ( .B1(n7742), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9040), .ZN(
        n9055) );
  XNOR2_X1 U9424 ( .A(n7743), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9054) );
  NOR2_X1 U9425 ( .A1(n9055), .A2(n9054), .ZN(n9053) );
  AOI21_X1 U9426 ( .B1(n7743), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9053), .ZN(
        n9719) );
  NAND2_X1 U9427 ( .A1(n9718), .A2(n9719), .ZN(n9717) );
  OAI21_X1 U9428 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n7744), .A(n9717), .ZN(
        n7745) );
  XNOR2_X1 U9429 ( .A(n7745), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n7749) );
  OAI21_X1 U9430 ( .B1(n7749), .B2(n9623), .A(n9715), .ZN(n7746) );
  AOI21_X1 U9431 ( .B1(n7748), .B2(n7747), .A(n7746), .ZN(n7752) );
  AOI22_X1 U9432 ( .A1(n7750), .A2(n9711), .B1(n9720), .B2(n7749), .ZN(n7751)
         );
  MUX2_X1 U9433 ( .A(n7752), .B(n7751), .S(n9761), .Z(n7754) );
  NAND2_X1 U9434 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3084), .ZN(n7753) );
  OAI211_X1 U9435 ( .C1(n5127), .C2(n9724), .A(n7754), .B(n7753), .ZN(P1_U3260) );
  XNOR2_X1 U9436 ( .A(n7755), .B(n8971), .ZN(n9589) );
  AOI211_X1 U9437 ( .C1(n9586), .C2(n9574), .A(n9749), .B(n7756), .ZN(n9584)
         );
  NOR2_X1 U9438 ( .A1(n9318), .A2(n9597), .ZN(n7760) );
  OAI22_X1 U9439 ( .A1(n9222), .A2(n7758), .B1(n7757), .B2(n9319), .ZN(n7759)
         );
  AOI211_X1 U9440 ( .C1(n9325), .C2(n9441), .A(n7760), .B(n7759), .ZN(n7761)
         );
  OAI21_X1 U9441 ( .B1(n7762), .B2(n9781), .A(n7761), .ZN(n7768) );
  OR2_X1 U9442 ( .A1(n7763), .A2(n8971), .ZN(n7764) );
  NAND2_X1 U9443 ( .A1(n7765), .A2(n7764), .ZN(n7766) );
  NAND2_X1 U9444 ( .A1(n7766), .A2(n9427), .ZN(n9587) );
  NOR2_X1 U9445 ( .A1(n9587), .A2(n9779), .ZN(n7767) );
  AOI211_X1 U9446 ( .C1(n9584), .C2(n9787), .A(n7768), .B(n7767), .ZN(n7769)
         );
  OAI21_X1 U9447 ( .B1(n9589), .B2(n9331), .A(n7769), .ZN(P1_U3278) );
  INV_X1 U9448 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10426) );
  OR2_X1 U9449 ( .A1(n8855), .A2(n10426), .ZN(n7771) );
  NAND2_X1 U9450 ( .A1(n9352), .A2(n7773), .ZN(n7775) );
  INV_X1 U9451 ( .A(n9356), .ZN(n9029) );
  NAND2_X1 U9452 ( .A1(n9029), .A2(n6067), .ZN(n7774) );
  NAND2_X1 U9453 ( .A1(n7775), .A2(n7774), .ZN(n7777) );
  XNOR2_X1 U9454 ( .A(n7777), .B(n7776), .ZN(n7781) );
  NAND2_X1 U9455 ( .A1(n9352), .A2(n6067), .ZN(n7778) );
  OAI21_X1 U9456 ( .B1(n9356), .B2(n7779), .A(n7778), .ZN(n7780) );
  XNOR2_X1 U9457 ( .A(n7781), .B(n7780), .ZN(n7782) );
  INV_X1 U9458 ( .A(n7782), .ZN(n7794) );
  NAND3_X1 U9459 ( .A1(n7794), .A2(n8732), .A3(n7793), .ZN(n7799) );
  INV_X1 U9460 ( .A(n7783), .ZN(n9141) );
  AOI22_X1 U9461 ( .A1(n9141), .A2(n8721), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n7792) );
  OR2_X1 U9462 ( .A1(n9127), .A2(n7784), .ZN(n7790) );
  INV_X1 U9463 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7787) );
  NAND2_X1 U9464 ( .A1(n8750), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n7786) );
  NAND2_X1 U9465 ( .A1(n8751), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7785) );
  OAI211_X1 U9466 ( .C1(n4479), .C2(n7787), .A(n7786), .B(n7785), .ZN(n7788)
         );
  INV_X1 U9467 ( .A(n7788), .ZN(n7789) );
  NAND2_X1 U9468 ( .A1(n7790), .A2(n7789), .ZN(n9028) );
  NAND2_X1 U9469 ( .A1(n9028), .A2(n8725), .ZN(n7791) );
  OAI211_X1 U9470 ( .C1(n9172), .C2(n8723), .A(n7792), .B(n7791), .ZN(n7796)
         );
  NOR3_X1 U9471 ( .A1(n7794), .A2(n8712), .A3(n7793), .ZN(n7795) );
  AOI211_X1 U9472 ( .C1(n9352), .C2(n8710), .A(n7796), .B(n7795), .ZN(n7797)
         );
  OAI211_X1 U9473 ( .C1(n7800), .C2(n7799), .A(n7798), .B(n7797), .ZN(P1_U3218) );
  OAI222_X1 U9474 ( .A1(n7729), .A2(n7802), .B1(n8612), .B2(n7801), .C1(n5827), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  OAI22_X1 U9475 ( .A1(n7804), .A2(n8426), .B1(n7803), .B2(n8428), .ZN(n9937)
         );
  OAI21_X1 U9476 ( .B1(n7807), .B2(n7806), .A(n7805), .ZN(n7808) );
  AOI22_X1 U9477 ( .A1(n8066), .A2(n9937), .B1(n8117), .B2(n7808), .ZN(n7811)
         );
  NAND2_X1 U9478 ( .A1(n7809), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7810) );
  OAI211_X1 U9479 ( .C1(n9967), .C2(n8123), .A(n7811), .B(n7810), .ZN(P2_U3239) );
  NAND2_X1 U9480 ( .A1(n8571), .A2(n8130), .ZN(n7846) );
  NAND2_X1 U9481 ( .A1(n8568), .A2(n8152), .ZN(n7940) );
  OR2_X1 U9482 ( .A1(n8559), .A2(n8427), .ZN(n7942) );
  NAND2_X1 U9483 ( .A1(n8559), .A2(n8427), .ZN(n7944) );
  NAND2_X1 U9484 ( .A1(n7942), .A2(n7944), .ZN(n8446) );
  INV_X1 U9485 ( .A(n8445), .ZN(n7815) );
  NOR2_X1 U9486 ( .A1(n8446), .A2(n7815), .ZN(n7816) );
  NAND2_X1 U9487 ( .A1(n8554), .A2(n8151), .ZN(n7945) );
  NAND2_X1 U9488 ( .A1(n7948), .A2(n7945), .ZN(n8438) );
  XNOR2_X1 U9489 ( .A(n8549), .B(n8429), .ZN(n8419) );
  NAND2_X1 U9490 ( .A1(n8549), .A2(n8429), .ZN(n7950) );
  NAND2_X1 U9491 ( .A1(n8546), .A2(n8150), .ZN(n7952) );
  NAND2_X1 U9492 ( .A1(n7955), .A2(n7952), .ZN(n8394) );
  XNOR2_X1 U9493 ( .A(n8538), .B(n8273), .ZN(n8378) );
  NAND2_X1 U9494 ( .A1(n8379), .A2(n8378), .ZN(n8377) );
  INV_X1 U9495 ( .A(n8273), .ZN(n8369) );
  NAND2_X1 U9496 ( .A1(n8538), .A2(n8369), .ZN(n7958) );
  NAND2_X1 U9497 ( .A1(n8377), .A2(n7958), .ZN(n8368) );
  NAND2_X1 U9498 ( .A1(n8533), .A2(n8149), .ZN(n7959) );
  NAND2_X1 U9499 ( .A1(n7961), .A2(n7959), .ZN(n8367) );
  NAND2_X1 U9500 ( .A1(n8529), .A2(n8370), .ZN(n7843) );
  INV_X1 U9501 ( .A(n8278), .ZN(n8317) );
  NAND2_X1 U9502 ( .A1(n8523), .A2(n8317), .ZN(n7965) );
  OR2_X1 U9503 ( .A1(n8281), .A2(n8297), .ZN(n7969) );
  NAND2_X1 U9504 ( .A1(n8511), .A2(n8257), .ZN(n7818) );
  NAND2_X1 U9505 ( .A1(n8294), .A2(n7993), .ZN(n8299) );
  NAND2_X1 U9506 ( .A1(n8853), .A2(n5220), .ZN(n7821) );
  OR2_X1 U9507 ( .A1(n5221), .A2(n8609), .ZN(n7820) );
  NAND2_X1 U9508 ( .A1(n8288), .A2(n8296), .ZN(n7978) );
  INV_X1 U9509 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8608) );
  NOR2_X1 U9510 ( .A1(n5221), .A2(n8608), .ZN(n7822) );
  INV_X1 U9511 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n7826) );
  NAND2_X1 U9512 ( .A1(n5822), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n7825) );
  NAND2_X1 U9513 ( .A1(n7823), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7824) );
  OAI211_X1 U9514 ( .C1(n7827), .C2(n7826), .A(n7825), .B(n7824), .ZN(n8147)
         );
  AND2_X1 U9515 ( .A1(n8503), .A2(n8147), .ZN(n7841) );
  MUX2_X1 U9516 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7832), .Z(n7833) );
  INV_X1 U9517 ( .A(SI_31_), .ZN(n10204) );
  NOR2_X1 U9518 ( .A1(n5221), .A2(n6541), .ZN(n7834) );
  INV_X1 U9519 ( .A(n8246), .ZN(n8496) );
  INV_X1 U9520 ( .A(n7835), .ZN(n8245) );
  INV_X1 U9521 ( .A(n8147), .ZN(n8256) );
  NAND2_X1 U9522 ( .A1(n8250), .A2(n8256), .ZN(n7981) );
  NOR2_X1 U9523 ( .A1(n8246), .A2(n7835), .ZN(n7986) );
  AOI21_X1 U9524 ( .B1(n7836), .B2(n8017), .A(n7986), .ZN(n7837) );
  NOR2_X1 U9525 ( .A1(n7986), .A2(n7841), .ZN(n8018) );
  AND2_X1 U9526 ( .A1(n8023), .A2(n8356), .ZN(n7840) );
  MUX2_X1 U9527 ( .A(n8017), .B(n8018), .S(n7984), .Z(n7989) );
  INV_X1 U9528 ( .A(n7841), .ZN(n7982) );
  OR2_X1 U9529 ( .A1(n8523), .A2(n8317), .ZN(n7964) );
  NAND2_X1 U9530 ( .A1(n7964), .A2(n7842), .ZN(n7845) );
  NAND2_X1 U9531 ( .A1(n8333), .A2(n7843), .ZN(n7844) );
  MUX2_X1 U9532 ( .A(n7845), .B(n7844), .S(n7984), .Z(n7968) );
  AND2_X1 U9533 ( .A1(n7940), .A2(n7846), .ZN(n7847) );
  MUX2_X1 U9534 ( .A(n7848), .B(n7847), .S(n7976), .Z(n7934) );
  AND2_X1 U9535 ( .A1(n7877), .A2(n7876), .ZN(n7851) );
  AND2_X1 U9536 ( .A1(n7863), .A2(n7849), .ZN(n7850) );
  MUX2_X1 U9537 ( .A(n7851), .B(n7850), .S(n7976), .Z(n7874) );
  AND2_X1 U9538 ( .A1(n7867), .A2(n8023), .ZN(n7854) );
  AND2_X1 U9539 ( .A1(n7853), .A2(n7852), .ZN(n7866) );
  OAI21_X1 U9540 ( .B1(n7855), .B2(n7854), .A(n7866), .ZN(n7856) );
  NAND3_X1 U9541 ( .A1(n7856), .A2(n7870), .A3(n7984), .ZN(n7857) );
  NAND3_X1 U9542 ( .A1(n7874), .A2(n7858), .A3(n7857), .ZN(n7865) );
  OAI21_X1 U9543 ( .B1(n7860), .B2(n5014), .A(n7874), .ZN(n7862) );
  NAND4_X1 U9544 ( .A1(n7865), .A2(n7863), .A3(n7862), .A4(n7861), .ZN(n7864)
         );
  NAND2_X1 U9545 ( .A1(n7864), .A2(n7984), .ZN(n7873) );
  INV_X1 U9546 ( .A(n7865), .ZN(n7871) );
  INV_X1 U9547 ( .A(n6695), .ZN(n7868) );
  OAI21_X1 U9548 ( .B1(n7868), .B2(n7867), .A(n7866), .ZN(n7869) );
  NAND3_X1 U9549 ( .A1(n7871), .A2(n7870), .A3(n7869), .ZN(n7872) );
  OR2_X1 U9550 ( .A1(n7884), .A2(n7883), .ZN(n7881) );
  INV_X1 U9551 ( .A(n7874), .ZN(n7879) );
  AND2_X1 U9552 ( .A1(n7876), .A2(n7875), .ZN(n7878) );
  OAI211_X1 U9553 ( .C1(n7879), .C2(n7878), .A(n7877), .B(n7881), .ZN(n7880)
         );
  NAND3_X1 U9554 ( .A1(n7884), .A2(n7883), .A3(n7976), .ZN(n7885) );
  MUX2_X1 U9555 ( .A(n7887), .B(n7886), .S(n7976), .Z(n7888) );
  MUX2_X1 U9556 ( .A(n7890), .B(n7889), .S(n7976), .Z(n7891) );
  NAND2_X1 U9557 ( .A1(n7892), .A2(n7891), .ZN(n7898) );
  AOI21_X1 U9558 ( .B1(n7899), .B2(n7897), .A(n7976), .ZN(n7895) );
  NAND2_X1 U9559 ( .A1(n7894), .A2(n7893), .ZN(n7900) );
  OR2_X1 U9560 ( .A1(n7895), .A2(n7900), .ZN(n7896) );
  AOI21_X1 U9561 ( .B1(n7898), .B2(n7897), .A(n7896), .ZN(n7905) );
  NAND2_X1 U9562 ( .A1(n7908), .A2(n7899), .ZN(n7903) );
  NAND2_X1 U9563 ( .A1(n7900), .A2(n7899), .ZN(n7901) );
  NAND2_X1 U9564 ( .A1(n7906), .A2(n7901), .ZN(n7902) );
  MUX2_X1 U9565 ( .A(n7903), .B(n7902), .S(n7984), .Z(n7904) );
  OR2_X1 U9566 ( .A1(n7905), .A2(n7904), .ZN(n7912) );
  NAND2_X1 U9567 ( .A1(n7912), .A2(n7906), .ZN(n7907) );
  AND2_X1 U9568 ( .A1(n7909), .A2(n7908), .ZN(n7911) );
  AOI21_X1 U9569 ( .B1(n7912), .B2(n7911), .A(n4694), .ZN(n7913) );
  NOR2_X1 U9570 ( .A1(n7921), .A2(n7914), .ZN(n7916) );
  AOI21_X1 U9571 ( .B1(n7926), .B2(n7916), .A(n4690), .ZN(n7918) );
  INV_X1 U9572 ( .A(n7919), .ZN(n7920) );
  OR2_X1 U9573 ( .A1(n7921), .A2(n7920), .ZN(n7922) );
  NOR2_X1 U9574 ( .A1(n5004), .A2(n7922), .ZN(n7925) );
  INV_X1 U9575 ( .A(n7923), .ZN(n7924) );
  AOI21_X1 U9576 ( .B1(n7926), .B2(n7925), .A(n7924), .ZN(n7928) );
  INV_X1 U9577 ( .A(n7930), .ZN(n7931) );
  MUX2_X1 U9578 ( .A(n7813), .B(n7931), .S(n7976), .Z(n7932) );
  NOR2_X1 U9579 ( .A1(n4527), .A2(n7932), .ZN(n7933) );
  NAND2_X1 U9580 ( .A1(n7941), .A2(n8445), .ZN(n7935) );
  OR2_X1 U9581 ( .A1(n8549), .A2(n8429), .ZN(n7947) );
  NAND2_X1 U9582 ( .A1(n7936), .A2(n7952), .ZN(n7937) );
  NAND2_X1 U9583 ( .A1(n7937), .A2(n7955), .ZN(n7938) );
  NAND2_X1 U9584 ( .A1(n8378), .A2(n7938), .ZN(n7939) );
  INV_X1 U9585 ( .A(n8378), .ZN(n8390) );
  NAND2_X1 U9586 ( .A1(n7941), .A2(n7940), .ZN(n7943) );
  NAND3_X1 U9587 ( .A1(n7943), .A2(n7942), .A3(n8445), .ZN(n7946) );
  NAND3_X1 U9588 ( .A1(n7946), .A2(n7945), .A3(n7944), .ZN(n7949) );
  NAND3_X1 U9589 ( .A1(n7949), .A2(n7948), .A3(n7947), .ZN(n7951) );
  NAND2_X1 U9590 ( .A1(n7951), .A2(n7950), .ZN(n7954) );
  INV_X1 U9591 ( .A(n7952), .ZN(n7953) );
  AOI21_X1 U9592 ( .B1(n7955), .B2(n7954), .A(n7953), .ZN(n7956) );
  NOR2_X1 U9593 ( .A1(n8390), .A2(n7956), .ZN(n7957) );
  NAND2_X1 U9594 ( .A1(n7959), .A2(n7958), .ZN(n7960) );
  NAND2_X1 U9595 ( .A1(n7960), .A2(n7984), .ZN(n7963) );
  OAI21_X1 U9596 ( .B1(n7976), .B2(n7961), .A(n8348), .ZN(n7962) );
  MUX2_X1 U9597 ( .A(n7965), .B(n7964), .S(n7984), .Z(n7966) );
  OAI211_X1 U9598 ( .C1(n7968), .C2(n7967), .A(n8313), .B(n7966), .ZN(n7972)
         );
  NAND2_X1 U9599 ( .A1(n8281), .A2(n8297), .ZN(n7970) );
  MUX2_X1 U9600 ( .A(n7970), .B(n7969), .S(n7976), .Z(n7971) );
  NAND3_X1 U9601 ( .A1(n7972), .A2(n7993), .A3(n7971), .ZN(n7975) );
  INV_X1 U9602 ( .A(n8257), .ZN(n8314) );
  MUX2_X1 U9603 ( .A(n8314), .B(n8511), .S(n7976), .Z(n7973) );
  OAI21_X1 U9604 ( .B1(n8257), .B2(n8309), .A(n7973), .ZN(n7974) );
  NAND3_X1 U9605 ( .A1(n7992), .A2(n7975), .A3(n7974), .ZN(n7980) );
  MUX2_X1 U9606 ( .A(n7978), .B(n7977), .S(n7976), .Z(n7979) );
  NAND4_X1 U9607 ( .A1(n7982), .A2(n7981), .A3(n7980), .A4(n7979), .ZN(n7988)
         );
  INV_X1 U9608 ( .A(n7983), .ZN(n7985) );
  MUX2_X1 U9609 ( .A(n7986), .B(n7985), .S(n7984), .Z(n7987) );
  AOI21_X1 U9610 ( .B1(n7989), .B2(n7988), .A(n7987), .ZN(n7990) );
  INV_X1 U9611 ( .A(n8446), .ZN(n8455) );
  NAND4_X1 U9612 ( .A1(n9935), .A2(n7995), .A3(n7994), .A4(n8022), .ZN(n7998)
         );
  NOR4_X1 U9613 ( .A1(n7998), .A2(n7997), .A3(n9920), .A4(n7996), .ZN(n8000)
         );
  NAND4_X1 U9614 ( .A1(n8001), .A2(n8000), .A3(n6916), .A4(n7999), .ZN(n8002)
         );
  NOR4_X1 U9615 ( .A1(n8005), .A2(n8004), .A3(n8003), .A4(n8002), .ZN(n8006)
         );
  NAND4_X1 U9616 ( .A1(n8009), .A2(n8008), .A3(n8007), .A4(n8006), .ZN(n8010)
         );
  NOR4_X1 U9617 ( .A1(n4527), .A2(n8011), .A3(n5004), .A4(n8010), .ZN(n8012)
         );
  NAND4_X1 U9618 ( .A1(n7817), .A2(n8455), .A3(n8465), .A4(n8012), .ZN(n8013)
         );
  NOR4_X1 U9619 ( .A1(n8367), .A2(n8419), .A3(n8394), .A4(n8013), .ZN(n8014)
         );
  NAND4_X1 U9620 ( .A1(n8348), .A2(n8014), .A3(n8333), .A4(n8378), .ZN(n8015)
         );
  NOR4_X1 U9621 ( .A1(n8284), .A2(n8319), .A3(n8302), .A4(n8015), .ZN(n8016)
         );
  NAND3_X1 U9622 ( .A1(n8018), .A2(n8017), .A3(n8016), .ZN(n8019) );
  XNOR2_X1 U9623 ( .A(n8019), .B(n8340), .ZN(n8024) );
  INV_X1 U9624 ( .A(n8020), .ZN(n8021) );
  OAI22_X1 U9625 ( .A1(n8024), .A2(n8023), .B1(n8022), .B2(n8021), .ZN(n8025)
         );
  NOR4_X1 U9626 ( .A1(n9956), .A2(n8243), .A3(n8029), .A4(n8426), .ZN(n8032)
         );
  OAI21_X1 U9627 ( .B1(n8033), .B2(n8030), .A(P2_B_REG_SCAN_IN), .ZN(n8031) );
  OAI22_X1 U9628 ( .A1(n8034), .A2(n8033), .B1(n8032), .B2(n8031), .ZN(
        P2_U3244) );
  OAI222_X1 U9629 ( .A1(n9499), .A2(n10426), .B1(n8036), .B2(n8035), .C1(n4480), .C2(P1_U3084), .ZN(P1_U3325) );
  XNOR2_X1 U9630 ( .A(n8037), .B(n8038), .ZN(n8044) );
  INV_X1 U9631 ( .A(n8322), .ZN(n8040) );
  OAI22_X1 U9632 ( .A1(n8040), .A2(n8128), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8039), .ZN(n8042) );
  OAI22_X1 U9633 ( .A1(n8257), .A2(n8131), .B1(n8317), .B2(n8129), .ZN(n8041)
         );
  AOI211_X1 U9634 ( .C1(n8281), .C2(n8143), .A(n8042), .B(n8041), .ZN(n8043)
         );
  OAI21_X1 U9635 ( .B1(n8044), .B2(n8145), .A(n8043), .ZN(P2_U3216) );
  XNOR2_X1 U9636 ( .A(n8046), .B(n8045), .ZN(n8051) );
  OAI22_X1 U9637 ( .A1(n8385), .A2(n8128), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8047), .ZN(n8049) );
  OAI22_X1 U9638 ( .A1(n8149), .A2(n8131), .B1(n8150), .B2(n8129), .ZN(n8048)
         );
  AOI211_X1 U9639 ( .C1(n8538), .C2(n8143), .A(n8049), .B(n8048), .ZN(n8050)
         );
  OAI21_X1 U9640 ( .B1(n8051), .B2(n8145), .A(n8050), .ZN(P2_U3218) );
  XOR2_X1 U9641 ( .A(n8053), .B(n8052), .Z(n8054) );
  NAND2_X1 U9642 ( .A1(n8054), .A2(n8117), .ZN(n8061) );
  AOI21_X1 U9643 ( .B1(n8066), .B2(n8056), .A(n8055), .ZN(n8060) );
  OR2_X1 U9644 ( .A1(n10022), .A2(n8123), .ZN(n8059) );
  OR2_X1 U9645 ( .A1(n8128), .A2(n8057), .ZN(n8058) );
  NAND4_X1 U9646 ( .A1(n8061), .A2(n8060), .A3(n8059), .A4(n8058), .ZN(
        P2_U3219) );
  AOI21_X1 U9647 ( .B1(n8062), .B2(n8063), .A(n4554), .ZN(n8070) );
  OR2_X1 U9648 ( .A1(n8151), .A2(n8428), .ZN(n8065) );
  OR2_X1 U9649 ( .A1(n8152), .A2(n8426), .ZN(n8064) );
  NAND2_X1 U9650 ( .A1(n8065), .A2(n8064), .ZN(n8448) );
  NAND2_X1 U9651 ( .A1(n8066), .A2(n8448), .ZN(n8067) );
  NAND2_X1 U9652 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8241) );
  OAI211_X1 U9653 ( .C1(n8128), .C2(n8451), .A(n8067), .B(n8241), .ZN(n8068)
         );
  AOI21_X1 U9654 ( .B1(n8559), .B2(n8143), .A(n8068), .ZN(n8069) );
  OAI21_X1 U9655 ( .B1(n8070), .B2(n8145), .A(n8069), .ZN(P2_U3221) );
  XNOR2_X1 U9656 ( .A(n8072), .B(n8071), .ZN(n8077) );
  OAI22_X1 U9657 ( .A1(n8128), .A2(n8415), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8073), .ZN(n8075) );
  OAI22_X1 U9658 ( .A1(n8131), .A2(n8150), .B1(n8151), .B2(n8129), .ZN(n8074)
         );
  AOI211_X1 U9659 ( .C1(n8549), .C2(n8143), .A(n8075), .B(n8074), .ZN(n8076)
         );
  OAI21_X1 U9660 ( .B1(n8077), .B2(n8145), .A(n8076), .ZN(P2_U3225) );
  XNOR2_X1 U9661 ( .A(n8079), .B(n8078), .ZN(n8085) );
  NOR2_X1 U9662 ( .A1(n8149), .A2(n8426), .ZN(n8080) );
  AOI21_X1 U9663 ( .B1(n8278), .B2(n9917), .A(n8080), .ZN(n8349) );
  INV_X1 U9664 ( .A(n8081), .ZN(n8357) );
  AOI22_X1 U9665 ( .A1(n8357), .A2(n8138), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8082) );
  OAI21_X1 U9666 ( .B1(n8349), .B2(n8141), .A(n8082), .ZN(n8083) );
  AOI21_X1 U9667 ( .B1(n8529), .B2(n8143), .A(n8083), .ZN(n8084) );
  OAI21_X1 U9668 ( .B1(n8085), .B2(n8145), .A(n8084), .ZN(P2_U3227) );
  INV_X1 U9669 ( .A(n8086), .ZN(n8088) );
  NOR3_X1 U9670 ( .A1(n8089), .A2(n8088), .A3(n8087), .ZN(n8092) );
  INV_X1 U9671 ( .A(n8090), .ZN(n8091) );
  OAI21_X1 U9672 ( .B1(n8092), .B2(n8091), .A(n8117), .ZN(n8097) );
  NOR2_X1 U9673 ( .A1(n10436), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8183) );
  OAI22_X1 U9674 ( .A1(n8131), .A2(n8130), .B1(n8093), .B2(n8129), .ZN(n8094)
         );
  AOI211_X1 U9675 ( .C1(n8138), .C2(n8095), .A(n8183), .B(n8094), .ZN(n8096)
         );
  OAI211_X1 U9676 ( .C1(n8098), .C2(n8123), .A(n8097), .B(n8096), .ZN(P2_U3228) );
  XNOR2_X1 U9677 ( .A(n8100), .B(n8099), .ZN(n8105) );
  INV_X1 U9678 ( .A(n8364), .ZN(n8101) );
  OAI22_X1 U9679 ( .A1(n8101), .A2(n8128), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10253), .ZN(n8103) );
  OAI22_X1 U9680 ( .A1(n8370), .A2(n8131), .B1(n8369), .B2(n8129), .ZN(n8102)
         );
  AOI211_X1 U9681 ( .C1(n8533), .C2(n8143), .A(n8103), .B(n8102), .ZN(n8104)
         );
  OAI21_X1 U9682 ( .B1(n8105), .B2(n8145), .A(n8104), .ZN(P2_U3231) );
  XNOR2_X1 U9683 ( .A(n8108), .B(n8107), .ZN(n8113) );
  INV_X1 U9684 ( .A(n8434), .ZN(n8109) );
  OAI22_X1 U9685 ( .A1(n8128), .A2(n8109), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10318), .ZN(n8111) );
  OAI22_X1 U9686 ( .A1(n8131), .A2(n8429), .B1(n8427), .B2(n8129), .ZN(n8110)
         );
  AOI211_X1 U9687 ( .C1(n8554), .C2(n8143), .A(n8111), .B(n8110), .ZN(n8112)
         );
  OAI21_X1 U9688 ( .B1(n8113), .B2(n8145), .A(n8112), .ZN(P2_U3235) );
  INV_X1 U9689 ( .A(n8546), .ZN(n8124) );
  OAI21_X1 U9690 ( .B1(n8116), .B2(n8115), .A(n8114), .ZN(n8118) );
  NAND2_X1 U9691 ( .A1(n8118), .A2(n8117), .ZN(n8122) );
  INV_X1 U9692 ( .A(n8402), .ZN(n8120) );
  INV_X1 U9693 ( .A(n8429), .ZN(n8271) );
  AOI22_X1 U9694 ( .A1(n8273), .A2(n9917), .B1(n8271), .B2(n9915), .ZN(n8397)
         );
  OAI22_X1 U9695 ( .A1(n8397), .A2(n8141), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10424), .ZN(n8119) );
  AOI21_X1 U9696 ( .B1(n8120), .B2(n8138), .A(n8119), .ZN(n8121) );
  OAI211_X1 U9697 ( .C1(n8124), .C2(n8123), .A(n8122), .B(n8121), .ZN(P2_U3237) );
  XNOR2_X1 U9698 ( .A(n8126), .B(n8125), .ZN(n8135) );
  INV_X1 U9699 ( .A(n8127), .ZN(n8472) );
  NAND2_X1 U9700 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8219) );
  OAI21_X1 U9701 ( .B1(n8128), .B2(n8472), .A(n8219), .ZN(n8133) );
  OAI22_X1 U9702 ( .A1(n8131), .A2(n8427), .B1(n8130), .B2(n8129), .ZN(n8132)
         );
  AOI211_X1 U9703 ( .C1(n8568), .C2(n8143), .A(n8133), .B(n8132), .ZN(n8134)
         );
  OAI21_X1 U9704 ( .B1(n8135), .B2(n8145), .A(n8134), .ZN(P2_U3240) );
  XNOR2_X1 U9705 ( .A(n8136), .B(n8137), .ZN(n8146) );
  AOI22_X1 U9706 ( .A1(n8280), .A2(n9917), .B1(n9915), .B2(n8277), .ZN(n8334)
         );
  INV_X1 U9707 ( .A(n8342), .ZN(n8139) );
  AOI22_X1 U9708 ( .A1(n8139), .A2(n8138), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8140) );
  OAI21_X1 U9709 ( .B1(n8334), .B2(n8141), .A(n8140), .ZN(n8142) );
  AOI21_X1 U9710 ( .B1(n8523), .B2(n8143), .A(n8142), .ZN(n8144) );
  OAI21_X1 U9711 ( .B1(n8146), .B2(n8145), .A(n8144), .ZN(P2_U3242) );
  MUX2_X1 U9712 ( .A(n8147), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8166), .Z(
        P2_U3582) );
  MUX2_X1 U9713 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8148), .S(P2_U3966), .Z(
        P2_U3581) );
  MUX2_X1 U9714 ( .A(n8314), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8166), .Z(
        P2_U3580) );
  MUX2_X1 U9715 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8280), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U9716 ( .A(n8278), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8166), .Z(
        P2_U3578) );
  MUX2_X1 U9717 ( .A(n8277), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8166), .Z(
        P2_U3577) );
  INV_X1 U9718 ( .A(n8149), .ZN(n8380) );
  MUX2_X1 U9719 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8380), .S(P2_U3966), .Z(
        P2_U3576) );
  MUX2_X1 U9720 ( .A(n8273), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8166), .Z(
        P2_U3575) );
  INV_X1 U9721 ( .A(n8150), .ZN(n8410) );
  MUX2_X1 U9722 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8410), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9723 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8271), .S(P2_U3966), .Z(
        P2_U3573) );
  INV_X1 U9724 ( .A(n8151), .ZN(n8409) );
  MUX2_X1 U9725 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8409), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9726 ( .A(n8467), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8166), .Z(
        P2_U3571) );
  INV_X1 U9727 ( .A(n8152), .ZN(n8265) );
  MUX2_X1 U9728 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8265), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9729 ( .A(n8466), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8166), .Z(
        P2_U3569) );
  MUX2_X1 U9730 ( .A(n8260), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8166), .Z(
        P2_U3568) );
  MUX2_X1 U9731 ( .A(n8153), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8166), .Z(
        P2_U3567) );
  MUX2_X1 U9732 ( .A(n8154), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8166), .Z(
        P2_U3566) );
  MUX2_X1 U9733 ( .A(n8155), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8166), .Z(
        P2_U3565) );
  MUX2_X1 U9734 ( .A(n8156), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8166), .Z(
        P2_U3564) );
  MUX2_X1 U9735 ( .A(n8157), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8166), .Z(
        P2_U3563) );
  INV_X1 U9736 ( .A(n8158), .ZN(n8159) );
  MUX2_X1 U9737 ( .A(n8159), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8166), .Z(
        P2_U3562) );
  MUX2_X1 U9738 ( .A(n8160), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8166), .Z(
        P2_U3561) );
  MUX2_X1 U9739 ( .A(n8161), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8166), .Z(
        P2_U3560) );
  MUX2_X1 U9740 ( .A(n8162), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8166), .Z(
        P2_U3559) );
  MUX2_X1 U9741 ( .A(n8163), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8166), .Z(
        P2_U3558) );
  MUX2_X1 U9742 ( .A(n9918), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8166), .Z(
        P2_U3557) );
  MUX2_X1 U9743 ( .A(n8164), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8166), .Z(
        P2_U3556) );
  MUX2_X1 U9744 ( .A(n9916), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8166), .Z(
        P2_U3555) );
  MUX2_X1 U9745 ( .A(n8165), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8166), .Z(
        P2_U3554) );
  MUX2_X1 U9746 ( .A(n4941), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8166), .Z(
        P2_U3553) );
  MUX2_X1 U9747 ( .A(n8167), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8166), .Z(
        P2_U3552) );
  OAI21_X1 U9748 ( .B1(n8174), .B2(P2_REG2_REG_14__SCAN_IN), .A(n8168), .ZN(
        n8186) );
  OAI21_X1 U9749 ( .B1(n8169), .B2(n7571), .A(n8188), .ZN(n8178) );
  INV_X1 U9750 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8172) );
  NAND2_X1 U9751 ( .A1(n9527), .A2(n4783), .ZN(n8171) );
  OAI211_X1 U9752 ( .C1(n8172), .C2(n8242), .A(n8171), .B(n8170), .ZN(n8177)
         );
  OAI21_X1 U9753 ( .B1(n8174), .B2(P2_REG1_REG_14__SCAN_IN), .A(n8173), .ZN(
        n8180) );
  XNOR2_X1 U9754 ( .A(n8180), .B(n8187), .ZN(n8175) );
  NOR2_X1 U9755 ( .A1(n5483), .A2(n8175), .ZN(n8181) );
  AOI211_X1 U9756 ( .C1(n8175), .C2(n5483), .A(n8181), .B(n8199), .ZN(n8176)
         );
  AOI211_X1 U9757 ( .C1(n9903), .C2(n8178), .A(n8177), .B(n8176), .ZN(n8179)
         );
  INV_X1 U9758 ( .A(n8179), .ZN(P2_U3260) );
  NOR2_X1 U9759 ( .A1(n8187), .A2(n8180), .ZN(n8182) );
  NOR2_X1 U9760 ( .A1(n8182), .A2(n8181), .ZN(n8196) );
  XNOR2_X1 U9761 ( .A(n8203), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8197) );
  XNOR2_X1 U9762 ( .A(n8196), .B(n8197), .ZN(n8195) );
  INV_X1 U9763 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8185) );
  INV_X1 U9764 ( .A(n8183), .ZN(n8184) );
  OAI21_X1 U9765 ( .B1(n8242), .B2(n8185), .A(n8184), .ZN(n8193) );
  NAND2_X1 U9766 ( .A1(n8187), .A2(n8186), .ZN(n8189) );
  XNOR2_X1 U9767 ( .A(n8203), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n8190) );
  AOI211_X1 U9768 ( .C1(n8191), .C2(n8190), .A(n9907), .B(n8202), .ZN(n8192)
         );
  AOI211_X1 U9769 ( .C1(n9527), .C2(n8203), .A(n8193), .B(n8192), .ZN(n8194)
         );
  OAI21_X1 U9770 ( .B1(n8195), .B2(n8199), .A(n8194), .ZN(P2_U3261) );
  XNOR2_X1 U9771 ( .A(n8218), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8201) );
  INV_X1 U9772 ( .A(n8196), .ZN(n8198) );
  OAI22_X1 U9773 ( .A1(n8198), .A2(n8197), .B1(P2_REG1_REG_16__SCAN_IN), .B2(
        n8203), .ZN(n8200) );
  NOR2_X1 U9774 ( .A1(n8200), .A2(n8201), .ZN(n8217) );
  AOI211_X1 U9775 ( .C1(n8201), .C2(n8200), .A(n8199), .B(n8217), .ZN(n8212)
         );
  NAND2_X1 U9776 ( .A1(n8218), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8204) );
  OAI21_X1 U9777 ( .B1(n8218), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8204), .ZN(
        n8205) );
  AOI211_X1 U9778 ( .C1(n8206), .C2(n8205), .A(n9907), .B(n8213), .ZN(n8211)
         );
  INV_X1 U9779 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8209) );
  NAND2_X1 U9780 ( .A1(n9527), .A2(n8218), .ZN(n8208) );
  NAND2_X1 U9781 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3152), .ZN(n8207) );
  OAI211_X1 U9782 ( .C1(n8209), .C2(n8242), .A(n8208), .B(n8207), .ZN(n8210)
         );
  OR3_X1 U9783 ( .A1(n8212), .A2(n8211), .A3(n8210), .ZN(P2_U3262) );
  OAI21_X1 U9784 ( .B1(n8214), .B2(n8473), .A(n8228), .ZN(n8215) );
  NAND2_X1 U9785 ( .A1(n8215), .A2(n9903), .ZN(n8224) );
  INV_X1 U9786 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8216) );
  XNOR2_X1 U9787 ( .A(n8232), .B(n8216), .ZN(n8231) );
  AOI21_X1 U9788 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8218), .A(n8217), .ZN(
        n8230) );
  XNOR2_X1 U9789 ( .A(n8231), .B(n8230), .ZN(n8222) );
  INV_X1 U9790 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8220) );
  OAI21_X1 U9791 ( .B1(n8242), .B2(n8220), .A(n8219), .ZN(n8221) );
  AOI21_X1 U9792 ( .B1(n9904), .B2(n8222), .A(n8221), .ZN(n8223) );
  OAI211_X1 U9793 ( .C1(n9906), .C2(n8225), .A(n8224), .B(n8223), .ZN(P2_U3263) );
  NAND2_X1 U9794 ( .A1(n8226), .A2(n8225), .ZN(n8227) );
  NAND2_X1 U9795 ( .A1(n8228), .A2(n8227), .ZN(n8229) );
  XNOR2_X1 U9796 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8229), .ZN(n8238) );
  NAND2_X1 U9797 ( .A1(n8231), .A2(n8230), .ZN(n8234) );
  OR2_X1 U9798 ( .A1(n8232), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8233) );
  NAND2_X1 U9799 ( .A1(n8234), .A2(n8233), .ZN(n8236) );
  XNOR2_X1 U9800 ( .A(n8236), .B(n8235), .ZN(n8239) );
  INV_X1 U9801 ( .A(n8239), .ZN(n8237) );
  AOI22_X1 U9802 ( .A1(n8238), .A2(n9903), .B1(n8237), .B2(n9904), .ZN(n8240)
         );
  INV_X1 U9803 ( .A(n8281), .ZN(n8516) );
  INV_X1 U9804 ( .A(n8538), .ZN(n8388) );
  INV_X1 U9805 ( .A(n8549), .ZN(n8418) );
  INV_X1 U9806 ( .A(n8559), .ZN(n8454) );
  OR2_X1 U9807 ( .A1(n8484), .A2(n8571), .ZN(n8485) );
  NAND2_X1 U9808 ( .A1(n8418), .A2(n8433), .ZN(n8412) );
  NAND2_X1 U9809 ( .A1(n8388), .A2(n8400), .ZN(n8382) );
  OR2_X2 U9810 ( .A1(n8288), .A2(n8304), .ZN(n8287) );
  XNOR2_X1 U9811 ( .A(n8249), .B(n8246), .ZN(n8498) );
  NOR2_X1 U9812 ( .A1(n8243), .A2(n10262), .ZN(n8244) );
  OR2_X1 U9813 ( .A1(n8428), .A2(n8244), .ZN(n8255) );
  NOR2_X1 U9814 ( .A1(n8245), .A2(n8255), .ZN(n8495) );
  INV_X1 U9815 ( .A(n8495), .ZN(n8501) );
  NOR2_X1 U9816 ( .A1(n9941), .A2(n8501), .ZN(n8251) );
  NOR2_X1 U9817 ( .A1(n8246), .A2(n9951), .ZN(n8247) );
  AOI211_X1 U9818 ( .C1(n9941), .C2(P2_REG2_REG_31__SCAN_IN), .A(n8251), .B(
        n8247), .ZN(n8248) );
  OAI21_X1 U9819 ( .B1(n8498), .B2(n9948), .A(n8248), .ZN(P2_U3265) );
  INV_X1 U9820 ( .A(n8249), .ZN(n8500) );
  NAND2_X1 U9821 ( .A1(n8250), .A2(n8287), .ZN(n8499) );
  NAND3_X1 U9822 ( .A1(n8500), .A2(n8442), .A3(n8499), .ZN(n8253) );
  AOI21_X1 U9823 ( .B1(n9941), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8251), .ZN(
        n8252) );
  OAI211_X1 U9824 ( .C1(n8503), .C2(n9951), .A(n8253), .B(n8252), .ZN(P2_U3266) );
  XNOR2_X1 U9825 ( .A(n8254), .B(n8284), .ZN(n8259) );
  OAI22_X1 U9826 ( .A1(n8257), .A2(n8426), .B1(n8256), .B2(n8255), .ZN(n8258)
         );
  AOI21_X1 U9827 ( .B1(n8259), .B2(n9938), .A(n8258), .ZN(n8508) );
  NAND2_X1 U9828 ( .A1(n8578), .A2(n8260), .ZN(n8261) );
  NAND2_X1 U9829 ( .A1(n8568), .A2(n8265), .ZN(n8264) );
  NAND2_X1 U9830 ( .A1(n8463), .A2(n8264), .ZN(n8267) );
  OR2_X1 U9831 ( .A1(n8568), .A2(n8265), .ZN(n8266) );
  NAND2_X1 U9832 ( .A1(n8267), .A2(n8266), .ZN(n8456) );
  NAND2_X1 U9833 ( .A1(n8559), .A2(n8467), .ZN(n8268) );
  NAND2_X1 U9834 ( .A1(n8458), .A2(n8268), .ZN(n8439) );
  NAND2_X1 U9835 ( .A1(n8439), .A2(n8438), .ZN(n8437) );
  NAND2_X1 U9836 ( .A1(n8554), .A2(n8409), .ZN(n8269) );
  NAND2_X1 U9837 ( .A1(n8437), .A2(n8269), .ZN(n8420) );
  OR2_X1 U9838 ( .A1(n8549), .A2(n8271), .ZN(n8270) );
  NAND2_X1 U9839 ( .A1(n8549), .A2(n8271), .ZN(n8272) );
  INV_X1 U9840 ( .A(n8394), .ZN(n8396) );
  NAND2_X1 U9841 ( .A1(n8538), .A2(n8273), .ZN(n8274) );
  OR2_X1 U9842 ( .A1(n8533), .A2(n8380), .ZN(n8276) );
  INV_X1 U9843 ( .A(n8348), .ZN(n8352) );
  INV_X1 U9844 ( .A(n8333), .ZN(n8329) );
  NAND2_X1 U9845 ( .A1(n8330), .A2(n8329), .ZN(n8328) );
  OR2_X1 U9846 ( .A1(n8523), .A2(n8278), .ZN(n8279) );
  NAND2_X1 U9847 ( .A1(n8328), .A2(n8279), .ZN(n8320) );
  NAND2_X1 U9848 ( .A1(n8320), .A2(n8319), .ZN(n8318) );
  OR2_X1 U9849 ( .A1(n8281), .A2(n8280), .ZN(n8282) );
  NAND2_X1 U9850 ( .A1(n8318), .A2(n8282), .ZN(n8303) );
  NAND2_X1 U9851 ( .A1(n8303), .A2(n8302), .ZN(n8301) );
  OR2_X1 U9852 ( .A1(n8511), .A2(n8314), .ZN(n8283) );
  NAND2_X1 U9853 ( .A1(n8301), .A2(n8283), .ZN(n8285) );
  NAND2_X1 U9854 ( .A1(n8288), .A2(n8304), .ZN(n8286) );
  NAND2_X1 U9855 ( .A1(n8287), .A2(n8286), .ZN(n8505) );
  NOR2_X1 U9856 ( .A1(n8505), .A2(n9948), .ZN(n8292) );
  INV_X1 U9857 ( .A(n8288), .ZN(n8504) );
  AOI22_X1 U9858 ( .A1(n8289), .A2(n9940), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n9941), .ZN(n8290) );
  OAI21_X1 U9859 ( .B1(n8504), .B2(n9951), .A(n8290), .ZN(n8291) );
  AOI211_X1 U9860 ( .C1(n8509), .C2(n9944), .A(n8292), .B(n8291), .ZN(n8293)
         );
  OAI21_X1 U9861 ( .B1(n8508), .B2(n9941), .A(n8293), .ZN(P2_U3267) );
  INV_X1 U9862 ( .A(n8294), .ZN(n8295) );
  AOI21_X1 U9863 ( .B1(n8295), .B2(n8302), .A(n8425), .ZN(n8300) );
  OAI22_X1 U9864 ( .A1(n8297), .A2(n8426), .B1(n8296), .B2(n8428), .ZN(n8298)
         );
  AOI21_X1 U9865 ( .B1(n8300), .B2(n8299), .A(n8298), .ZN(n8514) );
  OAI21_X1 U9866 ( .B1(n8303), .B2(n8302), .A(n8301), .ZN(n8510) );
  INV_X1 U9867 ( .A(n8304), .ZN(n8305) );
  AOI21_X1 U9868 ( .B1(n8511), .B2(n8321), .A(n8305), .ZN(n8512) );
  NAND2_X1 U9869 ( .A1(n8512), .A2(n8442), .ZN(n8308) );
  AOI22_X1 U9870 ( .A1(n8306), .A2(n9940), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n9941), .ZN(n8307) );
  OAI211_X1 U9871 ( .C1(n8309), .C2(n9951), .A(n8308), .B(n8307), .ZN(n8310)
         );
  AOI21_X1 U9872 ( .B1(n8510), .B2(n9944), .A(n8310), .ZN(n8311) );
  OAI21_X1 U9873 ( .B1(n8514), .B2(n9941), .A(n8311), .ZN(P2_U3268) );
  OAI211_X1 U9874 ( .C1(n4547), .C2(n8313), .A(n8312), .B(n9938), .ZN(n8316)
         );
  NAND2_X1 U9875 ( .A1(n8314), .A2(n9917), .ZN(n8315) );
  OAI211_X1 U9876 ( .C1(n8317), .C2(n8426), .A(n8316), .B(n8315), .ZN(n8518)
         );
  INV_X1 U9877 ( .A(n8518), .ZN(n8327) );
  OAI21_X1 U9878 ( .B1(n8320), .B2(n8319), .A(n8318), .ZN(n8520) );
  OAI21_X1 U9879 ( .B1(n8516), .B2(n8339), .A(n8321), .ZN(n8517) );
  NOR2_X1 U9880 ( .A1(n8517), .A2(n9948), .ZN(n8325) );
  AOI22_X1 U9881 ( .A1(n8322), .A2(n9940), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n9941), .ZN(n8323) );
  OAI21_X1 U9882 ( .B1(n8516), .B2(n9951), .A(n8323), .ZN(n8324) );
  AOI211_X1 U9883 ( .C1(n8520), .C2(n9944), .A(n8325), .B(n8324), .ZN(n8326)
         );
  OAI21_X1 U9884 ( .B1(n8327), .B2(n9941), .A(n8326), .ZN(P2_U3269) );
  OAI21_X1 U9885 ( .B1(n8330), .B2(n8329), .A(n8328), .ZN(n8331) );
  INV_X1 U9886 ( .A(n8331), .ZN(n8526) );
  OAI21_X1 U9887 ( .B1(n4545), .B2(n8333), .A(n8332), .ZN(n8336) );
  INV_X1 U9888 ( .A(n8334), .ZN(n8335) );
  AOI21_X1 U9889 ( .B1(n8336), .B2(n9938), .A(n8335), .ZN(n8525) );
  NAND2_X1 U9890 ( .A1(n8523), .A2(n8354), .ZN(n8337) );
  NAND2_X1 U9891 ( .A1(n8337), .A2(n10003), .ZN(n8338) );
  NOR2_X1 U9892 ( .A1(n8339), .A2(n8338), .ZN(n8522) );
  NAND2_X1 U9893 ( .A1(n8522), .A2(n8340), .ZN(n8341) );
  OAI211_X1 U9894 ( .C1(n9924), .C2(n8342), .A(n8525), .B(n8341), .ZN(n8343)
         );
  NAND2_X1 U9895 ( .A1(n8343), .A2(n9927), .ZN(n8345) );
  AOI22_X1 U9896 ( .A1(n8523), .A2(n8490), .B1(n9941), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8344) );
  OAI211_X1 U9897 ( .C1(n8526), .C2(n8478), .A(n8345), .B(n8344), .ZN(P2_U3270) );
  OAI211_X1 U9898 ( .C1(n8348), .C2(n8347), .A(n8346), .B(n9938), .ZN(n8350)
         );
  OAI21_X1 U9899 ( .B1(n8353), .B2(n8352), .A(n8351), .ZN(n8527) );
  INV_X1 U9900 ( .A(n8354), .ZN(n8355) );
  AOI211_X1 U9901 ( .C1(n8529), .C2(n8363), .A(n10036), .B(n8355), .ZN(n8528)
         );
  NOR2_X1 U9902 ( .A1(n9941), .A2(n8356), .ZN(n8487) );
  NAND2_X1 U9903 ( .A1(n8528), .A2(n8487), .ZN(n8359) );
  AOI22_X1 U9904 ( .A1(n8357), .A2(n9940), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n9941), .ZN(n8358) );
  OAI211_X1 U9905 ( .C1(n4887), .C2(n9951), .A(n8359), .B(n8358), .ZN(n8360)
         );
  AOI21_X1 U9906 ( .B1(n8527), .B2(n9944), .A(n8360), .ZN(n8361) );
  OAI21_X1 U9907 ( .B1(n8531), .B2(n9941), .A(n8361), .ZN(P2_U3271) );
  XNOR2_X1 U9908 ( .A(n8362), .B(n8367), .ZN(n8537) );
  AOI21_X1 U9909 ( .B1(n8533), .B2(n8382), .A(n4888), .ZN(n8534) );
  INV_X1 U9910 ( .A(n8533), .ZN(n8366) );
  AOI22_X1 U9911 ( .A1(n8364), .A2(n9940), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n9941), .ZN(n8365) );
  OAI21_X1 U9912 ( .B1(n8366), .B2(n9951), .A(n8365), .ZN(n8375) );
  AOI21_X1 U9913 ( .B1(n8368), .B2(n8367), .A(n8425), .ZN(n8373) );
  OAI22_X1 U9914 ( .A1(n8370), .A2(n8428), .B1(n8369), .B2(n8426), .ZN(n8371)
         );
  AOI21_X1 U9915 ( .B1(n8373), .B2(n8372), .A(n8371), .ZN(n8536) );
  NOR2_X1 U9916 ( .A1(n8536), .A2(n9941), .ZN(n8374) );
  AOI211_X1 U9917 ( .C1(n8534), .C2(n8442), .A(n8375), .B(n8374), .ZN(n8376)
         );
  OAI21_X1 U9918 ( .B1(n8478), .B2(n8537), .A(n8376), .ZN(P2_U3272) );
  OAI21_X1 U9919 ( .B1(n8379), .B2(n8378), .A(n8377), .ZN(n8381) );
  AOI222_X1 U9920 ( .A1(n9938), .A2(n8381), .B1(n8410), .B2(n9915), .C1(n8380), 
        .C2(n9917), .ZN(n8541) );
  INV_X1 U9921 ( .A(n8400), .ZN(n8384) );
  INV_X1 U9922 ( .A(n8382), .ZN(n8383) );
  AOI21_X1 U9923 ( .B1(n8538), .B2(n8384), .A(n8383), .ZN(n8539) );
  INV_X1 U9924 ( .A(n8385), .ZN(n8386) );
  AOI22_X1 U9925 ( .A1(n8386), .A2(n9940), .B1(P2_REG2_REG_23__SCAN_IN), .B2(
        n9941), .ZN(n8387) );
  OAI21_X1 U9926 ( .B1(n8388), .B2(n9951), .A(n8387), .ZN(n8392) );
  OAI21_X1 U9927 ( .B1(n4511), .B2(n8390), .A(n8389), .ZN(n8542) );
  NOR2_X1 U9928 ( .A1(n8542), .A2(n8478), .ZN(n8391) );
  AOI211_X1 U9929 ( .C1(n8539), .C2(n8442), .A(n8392), .B(n8391), .ZN(n8393)
         );
  OAI21_X1 U9930 ( .B1(n9941), .B2(n8541), .A(n8393), .ZN(P2_U3273) );
  XNOR2_X1 U9931 ( .A(n8395), .B(n8394), .ZN(n8548) );
  OAI211_X1 U9932 ( .C1(n8396), .C2(n4533), .A(n4493), .B(n9938), .ZN(n8398)
         );
  NAND2_X1 U9933 ( .A1(n8398), .A2(n8397), .ZN(n8544) );
  AND2_X1 U9934 ( .A1(n8546), .A2(n8412), .ZN(n8399) );
  OR2_X1 U9935 ( .A1(n8400), .A2(n8399), .ZN(n8543) );
  INV_X1 U9936 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8401) );
  OAI22_X1 U9937 ( .A1(n8402), .A2(n9924), .B1(n9927), .B2(n8401), .ZN(n8403)
         );
  AOI21_X1 U9938 ( .B1(n8546), .B2(n8490), .A(n8403), .ZN(n8404) );
  OAI21_X1 U9939 ( .B1(n8543), .B2(n9948), .A(n8404), .ZN(n8405) );
  AOI21_X1 U9940 ( .B1(n8544), .B2(n8406), .A(n8405), .ZN(n8407) );
  OAI21_X1 U9941 ( .B1(n8478), .B2(n8548), .A(n8407), .ZN(P2_U3274) );
  XNOR2_X1 U9942 ( .A(n8408), .B(n8419), .ZN(n8411) );
  AOI222_X1 U9943 ( .A1(n9938), .A2(n8411), .B1(n8410), .B2(n9917), .C1(n8409), 
        .C2(n9915), .ZN(n8552) );
  INV_X1 U9944 ( .A(n8412), .ZN(n8413) );
  AOI21_X1 U9945 ( .B1(n8549), .B2(n8414), .A(n8413), .ZN(n8550) );
  INV_X1 U9946 ( .A(n8415), .ZN(n8416) );
  AOI22_X1 U9947 ( .A1(n9941), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8416), .B2(
        n9940), .ZN(n8417) );
  OAI21_X1 U9948 ( .B1(n8418), .B2(n9951), .A(n8417), .ZN(n8422) );
  XNOR2_X1 U9949 ( .A(n8420), .B(n8419), .ZN(n8553) );
  NOR2_X1 U9950 ( .A1(n8553), .A2(n8478), .ZN(n8421) );
  AOI211_X1 U9951 ( .C1(n8550), .C2(n8442), .A(n8422), .B(n8421), .ZN(n8423)
         );
  OAI21_X1 U9952 ( .B1(n9941), .B2(n8552), .A(n8423), .ZN(P2_U3275) );
  AOI21_X1 U9953 ( .B1(n8424), .B2(n8438), .A(n8425), .ZN(n8432) );
  OAI22_X1 U9954 ( .A1(n8429), .A2(n8428), .B1(n8427), .B2(n8426), .ZN(n8430)
         );
  AOI21_X1 U9955 ( .B1(n8432), .B2(n8431), .A(n8430), .ZN(n8557) );
  AOI21_X1 U9956 ( .B1(n8554), .B2(n8450), .A(n8433), .ZN(n8555) );
  INV_X1 U9957 ( .A(n8554), .ZN(n8436) );
  AOI22_X1 U9958 ( .A1(n9941), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8434), .B2(
        n9940), .ZN(n8435) );
  OAI21_X1 U9959 ( .B1(n8436), .B2(n9951), .A(n8435), .ZN(n8441) );
  OAI21_X1 U9960 ( .B1(n8439), .B2(n8438), .A(n8437), .ZN(n8558) );
  NOR2_X1 U9961 ( .A1(n8558), .A2(n8478), .ZN(n8440) );
  AOI211_X1 U9962 ( .C1(n8555), .C2(n8442), .A(n8441), .B(n8440), .ZN(n8443)
         );
  OAI21_X1 U9963 ( .B1(n9941), .B2(n8557), .A(n8443), .ZN(P2_U3276) );
  NAND2_X1 U9964 ( .A1(n8444), .A2(n8445), .ZN(n8447) );
  XNOR2_X1 U9965 ( .A(n8447), .B(n8446), .ZN(n8449) );
  AOI21_X1 U9966 ( .B1(n8449), .B2(n9938), .A(n8448), .ZN(n8563) );
  OAI211_X1 U9967 ( .C1(n8454), .C2(n8471), .A(n10003), .B(n8450), .ZN(n8561)
         );
  INV_X1 U9968 ( .A(n8561), .ZN(n8461) );
  INV_X1 U9969 ( .A(n8451), .ZN(n8452) );
  AOI22_X1 U9970 ( .A1(n9941), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8452), .B2(
        n9940), .ZN(n8453) );
  OAI21_X1 U9971 ( .B1(n8454), .B2(n9951), .A(n8453), .ZN(n8460) );
  NAND2_X1 U9972 ( .A1(n8456), .A2(n8455), .ZN(n8457) );
  NAND2_X1 U9973 ( .A1(n8458), .A2(n8457), .ZN(n8564) );
  NOR2_X1 U9974 ( .A1(n8564), .A2(n8478), .ZN(n8459) );
  AOI211_X1 U9975 ( .C1(n8461), .C2(n8487), .A(n8460), .B(n8459), .ZN(n8462)
         );
  OAI21_X1 U9976 ( .B1(n9941), .B2(n8563), .A(n8462), .ZN(P2_U3277) );
  XNOR2_X1 U9977 ( .A(n8463), .B(n8465), .ZN(n8570) );
  OAI211_X1 U9978 ( .C1(n8465), .C2(n8464), .A(n8444), .B(n9938), .ZN(n8469)
         );
  AOI22_X1 U9979 ( .A1(n8467), .A2(n9917), .B1(n9915), .B2(n8466), .ZN(n8468)
         );
  NAND2_X1 U9980 ( .A1(n8469), .A2(n8468), .ZN(n8566) );
  AND2_X1 U9981 ( .A1(n8568), .A2(n8485), .ZN(n8470) );
  OR2_X1 U9982 ( .A1(n8471), .A2(n8470), .ZN(n8565) );
  OAI22_X1 U9983 ( .A1(n9927), .A2(n8473), .B1(n8472), .B2(n9924), .ZN(n8474)
         );
  AOI21_X1 U9984 ( .B1(n8568), .B2(n8490), .A(n8474), .ZN(n8475) );
  OAI21_X1 U9985 ( .B1(n8565), .B2(n9948), .A(n8475), .ZN(n8476) );
  AOI21_X1 U9986 ( .B1(n8566), .B2(n9927), .A(n8476), .ZN(n8477) );
  OAI21_X1 U9987 ( .B1(n8570), .B2(n8478), .A(n8477), .ZN(P2_U3278) );
  XNOR2_X1 U9988 ( .A(n8479), .B(n4527), .ZN(n8481) );
  AOI21_X1 U9989 ( .B1(n8481), .B2(n9938), .A(n8480), .ZN(n8576) );
  OAI21_X1 U9990 ( .B1(n8483), .B2(n4527), .A(n8482), .ZN(n8575) );
  AOI21_X1 U9991 ( .B1(n8484), .B2(n8571), .A(n10036), .ZN(n8486) );
  NAND2_X1 U9992 ( .A1(n8486), .A2(n8485), .ZN(n8573) );
  INV_X1 U9993 ( .A(n8487), .ZN(n8492) );
  OAI22_X1 U9994 ( .A1(n9927), .A2(n4776), .B1(n8488), .B2(n9924), .ZN(n8489)
         );
  AOI21_X1 U9995 ( .B1(n8571), .B2(n8490), .A(n8489), .ZN(n8491) );
  OAI21_X1 U9996 ( .B1(n8573), .B2(n8492), .A(n8491), .ZN(n8493) );
  AOI21_X1 U9997 ( .B1(n8575), .B2(n9944), .A(n8493), .ZN(n8494) );
  OAI21_X1 U9998 ( .B1(n8576), .B2(n9941), .A(n8494), .ZN(P2_U3279) );
  AOI21_X1 U9999 ( .B1(n8496), .B2(n10002), .A(n8495), .ZN(n8497) );
  OAI21_X1 U10000 ( .B1(n8498), .B2(n10036), .A(n8497), .ZN(n8583) );
  MUX2_X1 U10001 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8583), .S(n10064), .Z(
        P2_U3551) );
  NAND3_X1 U10002 ( .A1(n8500), .A2(n10003), .A3(n8499), .ZN(n8502) );
  OAI211_X1 U10003 ( .C1(n8503), .C2(n10034), .A(n8502), .B(n8501), .ZN(n8584)
         );
  MUX2_X1 U10004 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8584), .S(n10064), .Z(
        P2_U3550) );
  OAI22_X1 U10005 ( .A1(n8505), .A2(n10036), .B1(n8504), .B2(n10034), .ZN(
        n8506) );
  INV_X1 U10006 ( .A(n8510), .ZN(n8515) );
  AOI22_X1 U10007 ( .A1(n8512), .A2(n10003), .B1(n10002), .B2(n8511), .ZN(
        n8513) );
  OAI211_X1 U10008 ( .C1(n9995), .C2(n8515), .A(n8514), .B(n8513), .ZN(n8587)
         );
  MUX2_X1 U10009 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8587), .S(n10064), .Z(
        P2_U3548) );
  OAI22_X1 U10010 ( .A1(n8517), .A2(n10036), .B1(n8516), .B2(n10034), .ZN(
        n8519) );
  AOI211_X1 U10011 ( .C1(n10041), .C2(n8520), .A(n8519), .B(n8518), .ZN(n8521)
         );
  INV_X1 U10012 ( .A(n8521), .ZN(n8588) );
  MUX2_X1 U10013 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8588), .S(n10064), .Z(
        P2_U3547) );
  AOI21_X1 U10014 ( .B1(n10002), .B2(n8523), .A(n8522), .ZN(n8524) );
  OAI211_X1 U10015 ( .C1(n8526), .C2(n9995), .A(n8525), .B(n8524), .ZN(n8589)
         );
  MUX2_X1 U10016 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8589), .S(n10064), .Z(
        P2_U3546) );
  INV_X1 U10017 ( .A(n8527), .ZN(n8532) );
  AOI21_X1 U10018 ( .B1(n10002), .B2(n8529), .A(n8528), .ZN(n8530) );
  OAI211_X1 U10019 ( .C1(n8532), .C2(n9995), .A(n8531), .B(n8530), .ZN(n8590)
         );
  MUX2_X1 U10020 ( .A(n8590), .B(P2_REG1_REG_25__SCAN_IN), .S(n10062), .Z(
        P2_U3545) );
  AOI22_X1 U10021 ( .A1(n8534), .A2(n10003), .B1(n10002), .B2(n8533), .ZN(
        n8535) );
  OAI211_X1 U10022 ( .C1(n8537), .C2(n9995), .A(n8536), .B(n8535), .ZN(n8591)
         );
  MUX2_X1 U10023 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8591), .S(n10064), .Z(
        P2_U3544) );
  AOI22_X1 U10024 ( .A1(n8539), .A2(n10003), .B1(n10002), .B2(n8538), .ZN(
        n8540) );
  OAI211_X1 U10025 ( .C1(n9995), .C2(n8542), .A(n8541), .B(n8540), .ZN(n8592)
         );
  MUX2_X1 U10026 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8592), .S(n10064), .Z(
        P2_U3543) );
  NOR2_X1 U10027 ( .A1(n8543), .A2(n10036), .ZN(n8545) );
  AOI211_X1 U10028 ( .C1(n10002), .C2(n8546), .A(n8545), .B(n8544), .ZN(n8547)
         );
  OAI21_X1 U10029 ( .B1(n9995), .B2(n8548), .A(n8547), .ZN(n8593) );
  MUX2_X1 U10030 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8593), .S(n10064), .Z(
        P2_U3542) );
  AOI22_X1 U10031 ( .A1(n8550), .A2(n10003), .B1(n10002), .B2(n8549), .ZN(
        n8551) );
  OAI211_X1 U10032 ( .C1(n9995), .C2(n8553), .A(n8552), .B(n8551), .ZN(n8594)
         );
  MUX2_X1 U10033 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8594), .S(n10064), .Z(
        P2_U3541) );
  AOI22_X1 U10034 ( .A1(n8555), .A2(n10003), .B1(n10002), .B2(n8554), .ZN(
        n8556) );
  OAI211_X1 U10035 ( .C1(n8558), .C2(n9995), .A(n8557), .B(n8556), .ZN(n8595)
         );
  MUX2_X1 U10036 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8595), .S(n10064), .Z(
        P2_U3540) );
  NAND2_X1 U10037 ( .A1(n8559), .A2(n10002), .ZN(n8560) );
  AND2_X1 U10038 ( .A1(n8561), .A2(n8560), .ZN(n8562) );
  OAI211_X1 U10039 ( .C1(n8564), .C2(n9995), .A(n8563), .B(n8562), .ZN(n8596)
         );
  MUX2_X1 U10040 ( .A(n8596), .B(P2_REG1_REG_19__SCAN_IN), .S(n10062), .Z(
        P2_U3539) );
  NOR2_X1 U10041 ( .A1(n8565), .A2(n10036), .ZN(n8567) );
  AOI211_X1 U10042 ( .C1(n10002), .C2(n8568), .A(n8567), .B(n8566), .ZN(n8569)
         );
  OAI21_X1 U10043 ( .B1(n9995), .B2(n8570), .A(n8569), .ZN(n8597) );
  MUX2_X1 U10044 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8597), .S(n10064), .Z(
        P2_U3538) );
  NAND2_X1 U10045 ( .A1(n8571), .A2(n10002), .ZN(n8572) );
  NAND2_X1 U10046 ( .A1(n8573), .A2(n8572), .ZN(n8574) );
  AOI21_X1 U10047 ( .B1(n8575), .B2(n10041), .A(n8574), .ZN(n8577) );
  NAND2_X1 U10048 ( .A1(n8577), .A2(n8576), .ZN(n8598) );
  MUX2_X1 U10049 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8598), .S(n10064), .Z(
        P2_U3537) );
  AOI22_X1 U10050 ( .A1(n8579), .A2(n10003), .B1(n10002), .B2(n8578), .ZN(
        n8580) );
  OAI211_X1 U10051 ( .C1(n8582), .C2(n9995), .A(n8581), .B(n8580), .ZN(n8599)
         );
  MUX2_X1 U10052 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8599), .S(n10064), .Z(
        P2_U3536) );
  MUX2_X1 U10053 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8583), .S(n10043), .Z(
        P2_U3519) );
  MUX2_X1 U10054 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8584), .S(n10043), .Z(
        P2_U3518) );
  MUX2_X1 U10055 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8587), .S(n10043), .Z(
        P2_U3516) );
  MUX2_X1 U10056 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8588), .S(n10043), .Z(
        P2_U3515) );
  MUX2_X1 U10057 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8589), .S(n10043), .Z(
        P2_U3514) );
  MUX2_X1 U10058 ( .A(n8590), .B(P2_REG0_REG_25__SCAN_IN), .S(n10042), .Z(
        P2_U3513) );
  MUX2_X1 U10059 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8591), .S(n10043), .Z(
        P2_U3512) );
  MUX2_X1 U10060 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8592), .S(n10043), .Z(
        P2_U3511) );
  MUX2_X1 U10061 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8593), .S(n10043), .Z(
        P2_U3510) );
  MUX2_X1 U10062 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8594), .S(n10043), .Z(
        P2_U3509) );
  MUX2_X1 U10063 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8595), .S(n10043), .Z(
        P2_U3508) );
  MUX2_X1 U10064 ( .A(n8596), .B(P2_REG0_REG_19__SCAN_IN), .S(n10042), .Z(
        P2_U3507) );
  MUX2_X1 U10065 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8597), .S(n10043), .Z(
        P2_U3505) );
  MUX2_X1 U10066 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8598), .S(n10043), .Z(
        P2_U3502) );
  MUX2_X1 U10067 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8599), .S(n10043), .Z(
        P2_U3499) );
  NAND3_X1 U10068 ( .A1(n8600), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n8601) );
  OAI22_X1 U10069 ( .A1(n8602), .A2(n8601), .B1(n6541), .B2(n7729), .ZN(n8603)
         );
  AOI21_X1 U10070 ( .B1(n9503), .B2(n8604), .A(n8603), .ZN(n8605) );
  INV_X1 U10071 ( .A(n8605), .ZN(P2_U3327) );
  OAI222_X1 U10072 ( .A1(n7729), .A2(n8608), .B1(n8612), .B2(n8607), .C1(n8606), .C2(P2_U3152), .ZN(P2_U3328) );
  OAI222_X1 U10073 ( .A1(n8612), .A2(n8611), .B1(P2_U3152), .B2(n8610), .C1(
        n8609), .C2(n7729), .ZN(P2_U3329) );
  MUX2_X1 U10074 ( .A(n8613), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NAND2_X1 U10075 ( .A1(n4606), .A2(n8614), .ZN(n8616) );
  XNOR2_X1 U10076 ( .A(n8616), .B(n8615), .ZN(n8621) );
  NAND2_X1 U10077 ( .A1(n9215), .A2(n8725), .ZN(n8618) );
  AOI22_X1 U10078 ( .A1(n9218), .A2(n8721), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8617) );
  OAI211_X1 U10079 ( .C1(n9397), .C2(n8723), .A(n8618), .B(n8617), .ZN(n8619)
         );
  AOI21_X1 U10080 ( .B1(n9221), .B2(n8710), .A(n8619), .ZN(n8620) );
  OAI21_X1 U10081 ( .B1(n8621), .B2(n8712), .A(n8620), .ZN(P1_U3214) );
  XOR2_X1 U10082 ( .A(n8623), .B(n8622), .Z(n8628) );
  OAI22_X1 U10083 ( .A1(n8723), .A2(n9424), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8624), .ZN(n8626) );
  INV_X1 U10084 ( .A(n9106), .ZN(n9396) );
  OAI22_X1 U10085 ( .A1(n9396), .A2(n8735), .B1(n8736), .B2(n9284), .ZN(n8625)
         );
  AOI211_X1 U10086 ( .C1(n9283), .C2(n8710), .A(n8626), .B(n8625), .ZN(n8627)
         );
  OAI21_X1 U10087 ( .B1(n8628), .B2(n8712), .A(n8627), .ZN(P1_U3217) );
  XOR2_X1 U10088 ( .A(n8630), .B(n8629), .Z(n8635) );
  NAND2_X1 U10089 ( .A1(n9254), .A2(n8725), .ZN(n8632) );
  AOI22_X1 U10090 ( .A1(n8740), .A2(n9106), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8631) );
  OAI211_X1 U10091 ( .C1(n8736), .C2(n9250), .A(n8632), .B(n8631), .ZN(n8633)
         );
  AOI21_X1 U10092 ( .B1(n9400), .B2(n8710), .A(n8633), .ZN(n8634) );
  OAI21_X1 U10093 ( .B1(n8635), .B2(n8712), .A(n8634), .ZN(P1_U3221) );
  AOI21_X1 U10094 ( .B1(n8637), .B2(n8636), .A(n8717), .ZN(n8643) );
  NAND2_X1 U10095 ( .A1(n9186), .A2(n8725), .ZN(n8640) );
  INV_X1 U10096 ( .A(n8638), .ZN(n9193) );
  AOI22_X1 U10097 ( .A1(n9193), .A2(n8721), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8639) );
  OAI211_X1 U10098 ( .C1(n9113), .C2(n8723), .A(n8640), .B(n8639), .ZN(n8641)
         );
  AOI21_X1 U10099 ( .B1(n9192), .B2(n8710), .A(n8641), .ZN(n8642) );
  OAI21_X1 U10100 ( .B1(n8643), .B2(n8712), .A(n8642), .ZN(P1_U3223) );
  INV_X1 U10101 ( .A(n8644), .ZN(n8648) );
  OAI21_X1 U10102 ( .B1(n8646), .B2(n8648), .A(n8645), .ZN(n8647) );
  OAI21_X1 U10103 ( .B1(n8649), .B2(n8648), .A(n8647), .ZN(n8650) );
  NAND2_X1 U10104 ( .A1(n8650), .A2(n8732), .ZN(n8656) );
  NOR2_X1 U10105 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8651), .ZN(n9043) );
  OAI22_X1 U10106 ( .A1(n8736), .A2(n8653), .B1(n8723), .B2(n8652), .ZN(n8654)
         );
  AOI211_X1 U10107 ( .C1(n8725), .C2(n9414), .A(n9043), .B(n8654), .ZN(n8655)
         );
  OAI211_X1 U10108 ( .C1(n4771), .C2(n8743), .A(n8656), .B(n8655), .ZN(
        P1_U3224) );
  OAI21_X1 U10109 ( .B1(n8659), .B2(n8658), .A(n8657), .ZN(n8660) );
  NAND2_X1 U10110 ( .A1(n8660), .A2(n8732), .ZN(n8664) );
  NOR2_X1 U10111 ( .A1(n8735), .A2(n9424), .ZN(n8662) );
  OAI22_X1 U10112 ( .A1(n8736), .A2(n9320), .B1(n8723), .B2(n9423), .ZN(n8661)
         );
  AOI211_X1 U10113 ( .C1(P1_REG3_REG_17__SCAN_IN), .C2(P1_U3084), .A(n8662), 
        .B(n8661), .ZN(n8663) );
  OAI211_X1 U10114 ( .C1(n4769), .C2(n8743), .A(n8664), .B(n8663), .ZN(
        P1_U3226) );
  AOI21_X1 U10115 ( .B1(n8667), .B2(n8666), .A(n8665), .ZN(n8673) );
  NAND2_X1 U10116 ( .A1(n9372), .A2(n8725), .ZN(n8670) );
  INV_X1 U10117 ( .A(n8668), .ZN(n9205) );
  AOI22_X1 U10118 ( .A1(n9205), .A2(n8721), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8669) );
  OAI211_X1 U10119 ( .C1(n9207), .C2(n8723), .A(n8670), .B(n8669), .ZN(n8671)
         );
  AOI21_X1 U10120 ( .B1(n9210), .B2(n8710), .A(n8671), .ZN(n8672) );
  OAI21_X1 U10121 ( .B1(n8673), .B2(n8712), .A(n8672), .ZN(P1_U3227) );
  NOR2_X1 U10122 ( .A1(n8675), .A2(n4988), .ZN(n8676) );
  XNOR2_X1 U10123 ( .A(n8677), .B(n8676), .ZN(n8683) );
  OAI22_X1 U10124 ( .A1(n8723), .A2(n9265), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8678), .ZN(n8679) );
  AOI21_X1 U10125 ( .B1(n9269), .B2(n8721), .A(n8679), .ZN(n8680) );
  OAI21_X1 U10126 ( .B1(n9266), .B2(n8735), .A(n8680), .ZN(n8681) );
  AOI21_X1 U10127 ( .B1(n9406), .B2(n8710), .A(n8681), .ZN(n8682) );
  OAI21_X1 U10128 ( .B1(n8683), .B2(n8712), .A(n8682), .ZN(P1_U3231) );
  NOR2_X1 U10129 ( .A1(n8685), .A2(n8684), .ZN(n8687) );
  XNOR2_X1 U10130 ( .A(n8687), .B(n8686), .ZN(n8688) );
  NAND2_X1 U10131 ( .A1(n8688), .A2(n8732), .ZN(n8693) );
  NOR2_X1 U10132 ( .A1(n9266), .A2(n8723), .ZN(n8691) );
  OAI22_X1 U10133 ( .A1(n9231), .A2(n8736), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8689), .ZN(n8690) );
  AOI211_X1 U10134 ( .C1(n9386), .C2(n8725), .A(n8691), .B(n8690), .ZN(n8692)
         );
  OAI211_X1 U10135 ( .C1(n9480), .C2(n8743), .A(n8693), .B(n8692), .ZN(
        P1_U3233) );
  OAI21_X1 U10136 ( .B1(n8696), .B2(n8695), .A(n8694), .ZN(n8697) );
  NAND2_X1 U10137 ( .A1(n8697), .A2(n8732), .ZN(n8702) );
  AOI22_X1 U10138 ( .A1(n8699), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n8710), .B2(
        n8698), .ZN(n8701) );
  AOI22_X1 U10139 ( .A1(n8740), .A2(n9794), .B1(n8725), .B2(n9773), .ZN(n8700)
         );
  NAND3_X1 U10140 ( .A1(n8702), .A2(n8701), .A3(n8700), .ZN(P1_U3235) );
  INV_X1 U10141 ( .A(n8703), .ZN(n8704) );
  NOR2_X1 U10142 ( .A1(n8705), .A2(n8704), .ZN(n8707) );
  XNOR2_X1 U10143 ( .A(n8707), .B(n8706), .ZN(n8713) );
  NAND2_X1 U10144 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9712) );
  OAI21_X1 U10145 ( .B1(n8735), .B2(n9265), .A(n9712), .ZN(n8709) );
  OAI22_X1 U10146 ( .A1(n8736), .A2(n9298), .B1(n8723), .B2(n9302), .ZN(n8708)
         );
  AOI211_X1 U10147 ( .C1(n9307), .C2(n8710), .A(n8709), .B(n8708), .ZN(n8711)
         );
  OAI21_X1 U10148 ( .B1(n8713), .B2(n8712), .A(n8711), .ZN(P1_U3236) );
  INV_X1 U10149 ( .A(n9364), .ZN(n9177) );
  INV_X1 U10150 ( .A(n8714), .ZN(n8719) );
  OAI21_X1 U10151 ( .B1(n8717), .B2(n8716), .A(n8715), .ZN(n8718) );
  NAND3_X1 U10152 ( .A1(n8719), .A2(n8732), .A3(n8718), .ZN(n8727) );
  AOI22_X1 U10153 ( .A1(n9174), .A2(n8721), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n8722) );
  OAI21_X1 U10154 ( .B1(n9204), .B2(n8723), .A(n8722), .ZN(n8724) );
  AOI21_X1 U10155 ( .B1(n9030), .B2(n8725), .A(n8724), .ZN(n8726) );
  OAI211_X1 U10156 ( .C1(n9177), .C2(n8743), .A(n8727), .B(n8726), .ZN(
        P1_U3238) );
  NAND2_X1 U10157 ( .A1(n8729), .A2(n8728), .ZN(n8731) );
  XNOR2_X1 U10158 ( .A(n8731), .B(n8730), .ZN(n8733) );
  NAND2_X1 U10159 ( .A1(n8733), .A2(n8732), .ZN(n8742) );
  INV_X1 U10160 ( .A(n8734), .ZN(n8739) );
  OAI22_X1 U10161 ( .A1(n8737), .A2(n8736), .B1(n8735), .B2(n9423), .ZN(n8738)
         );
  AOI211_X1 U10162 ( .C1(n8740), .C2(n9441), .A(n8739), .B(n8738), .ZN(n8741)
         );
  OAI211_X1 U10163 ( .C1(n8744), .C2(n8743), .A(n8742), .B(n8741), .ZN(
        P1_U3239) );
  NAND2_X1 U10164 ( .A1(n8746), .A2(n6048), .ZN(n8749) );
  OR2_X1 U10165 ( .A1(n8855), .A2(n8747), .ZN(n8748) );
  INV_X1 U10166 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9337) );
  NAND2_X1 U10167 ( .A1(n8750), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8753) );
  NAND2_X1 U10168 ( .A1(n8751), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8752) );
  OAI211_X1 U10169 ( .C1(n4479), .C2(n9337), .A(n8753), .B(n8752), .ZN(n9099)
         );
  INV_X1 U10170 ( .A(n9099), .ZN(n8940) );
  OR2_X1 U10171 ( .A1(n9070), .A2(n8940), .ZN(n8938) );
  NAND2_X1 U10172 ( .A1(n8938), .A2(n9066), .ZN(n8755) );
  INV_X1 U10173 ( .A(n9454), .ZN(n9068) );
  NAND2_X1 U10174 ( .A1(n8755), .A2(n9068), .ZN(n9012) );
  INV_X1 U10175 ( .A(n9012), .ZN(n8862) );
  INV_X1 U10176 ( .A(n8864), .ZN(n8865) );
  OAI21_X1 U10177 ( .B1(n9844), .B2(n8865), .A(n9750), .ZN(n8759) );
  NAND2_X1 U10178 ( .A1(n9844), .A2(n8865), .ZN(n8756) );
  NAND2_X1 U10179 ( .A1(n8756), .A2(n9839), .ZN(n8758) );
  AOI21_X1 U10180 ( .B1(n8759), .B2(n8758), .A(n8757), .ZN(n8762) );
  NAND3_X1 U10181 ( .A1(n9756), .A2(n8865), .A3(n8760), .ZN(n8761) );
  OAI211_X1 U10182 ( .C1(n8763), .C2(n8865), .A(n8762), .B(n8761), .ZN(n8773)
         );
  NAND2_X1 U10183 ( .A1(n8901), .A2(n8764), .ZN(n8995) );
  INV_X1 U10184 ( .A(n8995), .ZN(n8766) );
  AND2_X1 U10185 ( .A1(n8778), .A2(n9730), .ZN(n8881) );
  INV_X1 U10186 ( .A(n8881), .ZN(n8765) );
  AOI21_X1 U10187 ( .B1(n8773), .B2(n8766), .A(n8765), .ZN(n8768) );
  INV_X1 U10188 ( .A(n8767), .ZN(n8904) );
  OAI21_X1 U10189 ( .B1(n8768), .B2(n8904), .A(n8905), .ZN(n8770) );
  NAND3_X1 U10190 ( .A1(n8770), .A2(n8798), .A3(n8769), .ZN(n8783) );
  INV_X1 U10191 ( .A(n8901), .ZN(n8771) );
  AOI21_X1 U10192 ( .B1(n8773), .B2(n8772), .A(n8771), .ZN(n8776) );
  OAI21_X1 U10193 ( .B1(n8776), .B2(n8775), .A(n8774), .ZN(n8779) );
  NAND3_X1 U10194 ( .A1(n8779), .A2(n8778), .A3(n8777), .ZN(n8781) );
  NAND4_X1 U10195 ( .A1(n8784), .A2(n8971), .A3(n8796), .A4(n8969), .ZN(n8807)
         );
  NAND2_X1 U10196 ( .A1(n9032), .A2(n8865), .ZN(n8787) );
  INV_X1 U10197 ( .A(n8908), .ZN(n8785) );
  NAND4_X1 U10198 ( .A1(n8785), .A2(n8865), .A3(n8796), .A4(n8909), .ZN(n8786)
         );
  NAND2_X1 U10199 ( .A1(n9441), .A2(n8865), .ZN(n8790) );
  OAI211_X1 U10200 ( .C1(n9586), .C2(n8787), .A(n8786), .B(n8790), .ZN(n8789)
         );
  NAND2_X1 U10201 ( .A1(n8789), .A2(n8788), .ZN(n8805) );
  NAND2_X1 U10202 ( .A1(n8906), .A2(n8908), .ZN(n8794) );
  INV_X1 U10203 ( .A(n8796), .ZN(n8907) );
  AOI21_X1 U10204 ( .B1(n8907), .B2(n9568), .A(n8790), .ZN(n8793) );
  NAND2_X1 U10205 ( .A1(n8796), .A2(n9032), .ZN(n8791) );
  NAND2_X1 U10206 ( .A1(n9586), .A2(n8791), .ZN(n8792) );
  NAND3_X1 U10207 ( .A1(n8794), .A2(n8793), .A3(n8792), .ZN(n8804) );
  OR2_X1 U10208 ( .A1(n8916), .A2(n8865), .ZN(n8803) );
  AND2_X1 U10209 ( .A1(n8906), .A2(n8864), .ZN(n8801) );
  AND2_X1 U10210 ( .A1(n8796), .A2(n8795), .ZN(n8797) );
  NAND2_X1 U10211 ( .A1(n8909), .A2(n8797), .ZN(n8913) );
  INV_X1 U10212 ( .A(n8798), .ZN(n8799) );
  NAND2_X1 U10213 ( .A1(n8909), .A2(n8799), .ZN(n8800) );
  NAND4_X1 U10214 ( .A1(n8911), .A2(n8801), .A3(n8913), .A4(n8800), .ZN(n8802)
         );
  AND4_X1 U10215 ( .A1(n8805), .A2(n8804), .A3(n8803), .A4(n8802), .ZN(n8806)
         );
  NAND2_X1 U10216 ( .A1(n8809), .A2(n8808), .ZN(n8811) );
  INV_X1 U10217 ( .A(n9103), .ZN(n8976) );
  MUX2_X1 U10218 ( .A(n8919), .B(n8917), .S(n8864), .Z(n8810) );
  NAND3_X1 U10219 ( .A1(n8811), .A2(n8976), .A3(n8810), .ZN(n8813) );
  OR2_X1 U10220 ( .A1(n9317), .A2(n9302), .ZN(n9292) );
  NAND2_X1 U10221 ( .A1(n9317), .A2(n9302), .ZN(n9291) );
  MUX2_X1 U10222 ( .A(n9077), .B(n9075), .S(n8864), .Z(n8812) );
  NAND3_X1 U10223 ( .A1(n8813), .A2(n9313), .A3(n8812), .ZN(n8816) );
  NAND2_X1 U10224 ( .A1(n8953), .A2(n9292), .ZN(n9081) );
  NAND2_X1 U10225 ( .A1(n9307), .A2(n9424), .ZN(n9080) );
  NAND2_X1 U10226 ( .A1(n9080), .A2(n9291), .ZN(n9079) );
  MUX2_X1 U10227 ( .A(n9081), .B(n9079), .S(n8864), .Z(n8814) );
  INV_X1 U10228 ( .A(n8814), .ZN(n8815) );
  NAND2_X1 U10229 ( .A1(n8816), .A2(n8815), .ZN(n8819) );
  NAND2_X1 U10230 ( .A1(n9283), .A2(n9265), .ZN(n9084) );
  NAND2_X1 U10231 ( .A1(n9084), .A2(n9080), .ZN(n8924) );
  INV_X1 U10232 ( .A(n8924), .ZN(n8817) );
  NAND2_X1 U10233 ( .A1(n8819), .A2(n8817), .ZN(n8818) );
  OR2_X1 U10234 ( .A1(n9406), .A2(n9396), .ZN(n9086) );
  OR2_X1 U10235 ( .A1(n9283), .A2(n9265), .ZN(n8952) );
  AND2_X1 U10236 ( .A1(n9086), .A2(n8952), .ZN(n8922) );
  NAND3_X1 U10237 ( .A1(n8819), .A2(n8953), .A3(n8952), .ZN(n8820) );
  AND2_X1 U10238 ( .A1(n9406), .A2(n9396), .ZN(n9085) );
  INV_X1 U10239 ( .A(n9085), .ZN(n8951) );
  OR2_X1 U10240 ( .A1(n9239), .A2(n9397), .ZN(n8949) );
  AND2_X1 U10241 ( .A1(n8949), .A2(n8950), .ZN(n8923) );
  INV_X1 U10242 ( .A(n8923), .ZN(n8824) );
  NAND2_X1 U10243 ( .A1(n9221), .A2(n9207), .ZN(n9002) );
  NAND2_X1 U10244 ( .A1(n9239), .A2(n9397), .ZN(n9089) );
  NAND2_X1 U10245 ( .A1(n8950), .A2(n9085), .ZN(n8821) );
  NAND2_X1 U10246 ( .A1(n9400), .A2(n9266), .ZN(n9088) );
  AND2_X1 U10247 ( .A1(n8821), .A2(n9088), .ZN(n8822) );
  NAND2_X1 U10248 ( .A1(n9089), .A2(n8822), .ZN(n8880) );
  NAND2_X1 U10249 ( .A1(n8880), .A2(n8949), .ZN(n8926) );
  OAI211_X1 U10250 ( .C1(n8823), .C2(n8824), .A(n9002), .B(n8926), .ZN(n8827)
         );
  OR2_X1 U10251 ( .A1(n9210), .A2(n9113), .ZN(n8935) );
  NAND2_X1 U10252 ( .A1(n8825), .A2(n8935), .ZN(n8826) );
  NAND2_X1 U10253 ( .A1(n9210), .A2(n9113), .ZN(n9182) );
  NAND2_X1 U10254 ( .A1(n9182), .A2(n9091), .ZN(n8835) );
  INV_X1 U10255 ( .A(n9091), .ZN(n8828) );
  NAND2_X1 U10256 ( .A1(n9182), .A2(n8828), .ZN(n8829) );
  NAND3_X1 U10257 ( .A1(n9167), .A2(n8935), .A3(n8829), .ZN(n8832) );
  INV_X1 U10258 ( .A(n8935), .ZN(n8830) );
  OAI21_X1 U10259 ( .B1(n8830), .B2(n9002), .A(n9093), .ZN(n8831) );
  INV_X1 U10260 ( .A(n8833), .ZN(n8834) );
  NAND2_X1 U10261 ( .A1(n9167), .A2(n9153), .ZN(n8878) );
  INV_X1 U10262 ( .A(n8878), .ZN(n8836) );
  NOR2_X1 U10263 ( .A1(n9094), .A2(n8836), .ZN(n8837) );
  MUX2_X1 U10264 ( .A(n9364), .B(n8837), .S(n8864), .Z(n8838) );
  INV_X1 U10265 ( .A(n8838), .ZN(n8839) );
  NAND2_X1 U10266 ( .A1(n8840), .A2(n8839), .ZN(n8847) );
  NAND2_X1 U10267 ( .A1(n8948), .A2(n9186), .ZN(n8841) );
  NAND2_X1 U10268 ( .A1(n9096), .A2(n8841), .ZN(n8843) );
  NAND2_X1 U10269 ( .A1(n9364), .A2(n9167), .ZN(n8879) );
  NAND2_X1 U10270 ( .A1(n8875), .A2(n8879), .ZN(n8842) );
  MUX2_X1 U10271 ( .A(n8843), .B(n8842), .S(n8864), .Z(n8844) );
  OAI21_X1 U10272 ( .B1(n8845), .B2(n9155), .A(n8844), .ZN(n8846) );
  NAND2_X1 U10273 ( .A1(n8847), .A2(n8846), .ZN(n8852) );
  NAND2_X1 U10274 ( .A1(n9352), .A2(n9356), .ZN(n8876) );
  MUX2_X1 U10275 ( .A(n8875), .B(n9096), .S(n8864), .Z(n8848) );
  AND2_X1 U10276 ( .A1(n9137), .A2(n8848), .ZN(n8851) );
  MUX2_X1 U10277 ( .A(n8876), .B(n8873), .S(n8865), .Z(n8849) );
  INV_X1 U10278 ( .A(n8849), .ZN(n8850) );
  AOI21_X1 U10279 ( .B1(n8852), .B2(n8851), .A(n8850), .ZN(n8863) );
  NAND2_X1 U10280 ( .A1(n8853), .A2(n6048), .ZN(n8857) );
  OR2_X1 U10281 ( .A1(n8855), .A2(n8854), .ZN(n8856) );
  NAND3_X1 U10282 ( .A1(n9012), .A2(n8863), .A3(n9126), .ZN(n8860) );
  NAND2_X1 U10283 ( .A1(n9099), .A2(n9066), .ZN(n8858) );
  NAND2_X1 U10284 ( .A1(n9070), .A2(n8858), .ZN(n9006) );
  INV_X1 U10285 ( .A(n9066), .ZN(n8859) );
  AOI21_X1 U10286 ( .B1(n8860), .B2(n9006), .A(n8985), .ZN(n8861) );
  MUX2_X1 U10287 ( .A(n8862), .B(n8861), .S(n8865), .Z(n8870) );
  INV_X1 U10288 ( .A(n9028), .ZN(n9347) );
  INV_X1 U10289 ( .A(n9126), .ZN(n9341) );
  INV_X1 U10290 ( .A(n9006), .ZN(n8866) );
  AOI21_X1 U10291 ( .B1(n8868), .B2(n8867), .A(n8866), .ZN(n8869) );
  NAND2_X1 U10292 ( .A1(n4721), .A2(n8871), .ZN(n8946) );
  INV_X1 U10293 ( .A(n8873), .ZN(n9097) );
  AOI21_X1 U10294 ( .B1(n9341), .B2(n9028), .A(n9097), .ZN(n8988) );
  NAND2_X1 U10295 ( .A1(n9096), .A2(n9094), .ZN(n8874) );
  NAND3_X1 U10296 ( .A1(n8876), .A2(n8875), .A3(n8874), .ZN(n8877) );
  AOI22_X1 U10297 ( .A1(n8988), .A2(n8877), .B1(n9347), .B2(n9126), .ZN(n9007)
         );
  NAND2_X1 U10298 ( .A1(n8879), .A2(n8878), .ZN(n9095) );
  NOR2_X1 U10299 ( .A1(n8880), .A2(n4826), .ZN(n8928) );
  INV_X1 U10300 ( .A(n9077), .ZN(n8921) );
  INV_X1 U10301 ( .A(n8917), .ZN(n8884) );
  INV_X1 U10302 ( .A(n8913), .ZN(n8882) );
  NAND4_X1 U10303 ( .A1(n8916), .A2(n8882), .A3(n8905), .A4(n8881), .ZN(n8883)
         );
  NOR4_X1 U10304 ( .A1(n9079), .A2(n8921), .A3(n8884), .A4(n8883), .ZN(n8885)
         );
  NAND2_X1 U10305 ( .A1(n8928), .A2(n8885), .ZN(n8999) );
  INV_X1 U10306 ( .A(n8999), .ZN(n8932) );
  AND2_X1 U10307 ( .A1(n8886), .A2(n4773), .ZN(n8954) );
  INV_X1 U10308 ( .A(n8954), .ZN(n8887) );
  OAI211_X1 U10309 ( .C1(n8889), .C2(n8888), .A(n8947), .B(n8887), .ZN(n8891)
         );
  NAND2_X1 U10310 ( .A1(n8891), .A2(n8890), .ZN(n8893) );
  OAI21_X1 U10311 ( .B1(n8894), .B2(n8893), .A(n8892), .ZN(n8898) );
  AND2_X1 U10312 ( .A1(n8896), .A2(n8895), .ZN(n8992) );
  INV_X1 U10313 ( .A(n8992), .ZN(n8897) );
  AOI21_X1 U10314 ( .B1(n8898), .B2(n8989), .A(n8897), .ZN(n8902) );
  NAND2_X1 U10315 ( .A1(n8997), .A2(n8899), .ZN(n8990) );
  OAI211_X1 U10316 ( .C1(n8902), .C2(n8990), .A(n8901), .B(n8900), .ZN(n8931)
         );
  AOI21_X1 U10317 ( .B1(n8905), .B2(n8904), .A(n8903), .ZN(n8914) );
  OAI21_X1 U10318 ( .B1(n8908), .B2(n8907), .A(n8906), .ZN(n8910) );
  NAND2_X1 U10319 ( .A1(n8910), .A2(n8909), .ZN(n8912) );
  OAI211_X1 U10320 ( .C1(n8914), .C2(n8913), .A(n8912), .B(n8911), .ZN(n8915)
         );
  NAND3_X1 U10321 ( .A1(n8917), .A2(n8916), .A3(n8915), .ZN(n8918) );
  AND3_X1 U10322 ( .A1(n9075), .A2(n8919), .A3(n8918), .ZN(n8920) );
  NOR3_X1 U10323 ( .A1(n9079), .A2(n8921), .A3(n8920), .ZN(n8929) );
  INV_X1 U10324 ( .A(n9081), .ZN(n8925) );
  OAI211_X1 U10325 ( .C1(n8925), .C2(n8924), .A(n8923), .B(n8922), .ZN(n8927)
         );
  AOI22_X1 U10326 ( .A1(n8929), .A2(n8928), .B1(n8927), .B2(n8926), .ZN(n8998)
         );
  INV_X1 U10327 ( .A(n8998), .ZN(n8930) );
  AOI21_X1 U10328 ( .B1(n8932), .B2(n8931), .A(n8930), .ZN(n8934) );
  INV_X1 U10329 ( .A(n9002), .ZN(n8933) );
  NOR2_X1 U10330 ( .A1(n8934), .A2(n8933), .ZN(n8936) );
  NAND2_X1 U10331 ( .A1(n8935), .A2(n9091), .ZN(n9001) );
  OAI21_X1 U10332 ( .B1(n8936), .B2(n9001), .A(n9093), .ZN(n8937) );
  NAND4_X1 U10333 ( .A1(n8988), .A2(n9150), .A3(n9095), .A4(n8937), .ZN(n8939)
         );
  INV_X1 U10334 ( .A(n8938), .ZN(n8986) );
  AOI21_X1 U10335 ( .B1(n9007), .B2(n8939), .A(n8986), .ZN(n8944) );
  INV_X1 U10336 ( .A(n9010), .ZN(n8942) );
  NAND2_X1 U10337 ( .A1(n9070), .A2(n8940), .ZN(n8941) );
  NAND2_X1 U10338 ( .A1(n8942), .A2(n8941), .ZN(n8987) );
  INV_X1 U10339 ( .A(n8985), .ZN(n8943) );
  OAI21_X1 U10340 ( .B1(n8944), .B2(n8987), .A(n8943), .ZN(n8945) );
  XNOR2_X1 U10341 ( .A(n8945), .B(n9761), .ZN(n9021) );
  NOR2_X1 U10342 ( .A1(n8947), .A2(n8946), .ZN(n9019) );
  NAND2_X1 U10343 ( .A1(n9364), .A2(n9186), .ZN(n9118) );
  NAND2_X1 U10344 ( .A1(n9119), .A2(n9118), .ZN(n9169) );
  INV_X1 U10345 ( .A(n9181), .ZN(n9183) );
  NAND2_X1 U10346 ( .A1(n8950), .A2(n9088), .ZN(n9244) );
  INV_X1 U10347 ( .A(n9244), .ZN(n9242) );
  NAND2_X1 U10348 ( .A1(n8951), .A2(n9086), .ZN(n9262) );
  NAND2_X1 U10349 ( .A1(n8952), .A2(n9084), .ZN(n9279) );
  NAND2_X1 U10350 ( .A1(n8953), .A2(n9080), .ZN(n9296) );
  NOR2_X1 U10351 ( .A1(n8955), .A2(n8954), .ZN(n9793) );
  INV_X1 U10352 ( .A(n9771), .ZN(n8958) );
  NAND4_X1 U10353 ( .A1(n9793), .A2(n8958), .A3(n8957), .A4(n8956), .ZN(n8960)
         );
  NOR2_X1 U10354 ( .A1(n8960), .A2(n8959), .ZN(n8965) );
  INV_X1 U10355 ( .A(n8961), .ZN(n8964) );
  NAND4_X1 U10356 ( .A1(n8965), .A2(n8964), .A3(n8963), .A4(n9766), .ZN(n8968)
         );
  NOR4_X1 U10357 ( .A1(n8968), .A2(n8967), .A3(n7313), .A4(n8966), .ZN(n8970)
         );
  NAND4_X1 U10358 ( .A1(n8971), .A2(n7606), .A3(n8970), .A4(n8969), .ZN(n8972)
         );
  NOR3_X1 U10359 ( .A1(n8974), .A2(n8973), .A3(n8972), .ZN(n8975) );
  NAND3_X1 U10360 ( .A1(n9313), .A2(n8976), .A3(n8975), .ZN(n8977) );
  OR3_X1 U10361 ( .A1(n9279), .A2(n9296), .A3(n8977), .ZN(n8978) );
  NOR2_X1 U10362 ( .A1(n9262), .A2(n8978), .ZN(n8979) );
  NAND3_X1 U10363 ( .A1(n9229), .A2(n9242), .A3(n8979), .ZN(n8980) );
  NOR2_X1 U10364 ( .A1(n9220), .A2(n8980), .ZN(n8981) );
  XNOR2_X1 U10365 ( .A(n9210), .B(n9113), .ZN(n9092) );
  INV_X1 U10366 ( .A(n9092), .ZN(n9201) );
  NAND4_X1 U10367 ( .A1(n9169), .A2(n9183), .A3(n8981), .A4(n9201), .ZN(n8982)
         );
  NOR2_X1 U10368 ( .A1(n9155), .A2(n8982), .ZN(n8983) );
  NAND3_X1 U10369 ( .A1(n9123), .A2(n9137), .A3(n8983), .ZN(n8984) );
  OR4_X2 U10370 ( .A1(n8987), .A2(n8986), .A3(n8985), .A4(n8984), .ZN(n9018)
         );
  INV_X1 U10371 ( .A(n8988), .ZN(n9009) );
  INV_X1 U10372 ( .A(n8989), .ZN(n8991) );
  AOI211_X1 U10373 ( .C1(n8993), .C2(n8992), .A(n8991), .B(n8990), .ZN(n8994)
         );
  AOI211_X1 U10374 ( .C1(n8997), .C2(n8996), .A(n8995), .B(n8994), .ZN(n9000)
         );
  OAI21_X1 U10375 ( .B1(n9000), .B2(n8999), .A(n8998), .ZN(n9003) );
  AOI21_X1 U10376 ( .B1(n9003), .B2(n9002), .A(n9001), .ZN(n9005) );
  INV_X1 U10377 ( .A(n9093), .ZN(n9004) );
  OAI211_X1 U10378 ( .C1(n9005), .C2(n9004), .A(n9096), .B(n9095), .ZN(n9008)
         );
  OAI211_X1 U10379 ( .C1(n9009), .C2(n9008), .A(n9007), .B(n9006), .ZN(n9011)
         );
  NAND2_X1 U10380 ( .A1(n4721), .A2(n9761), .ZN(n9014) );
  NOR3_X1 U10381 ( .A1(n9015), .A2(n9013), .A3(n9014), .ZN(n9017) );
  NOR3_X1 U10382 ( .A1(n9015), .A2(n9014), .A3(n9018), .ZN(n9016) );
  OAI21_X1 U10383 ( .B1(n4721), .B2(n9021), .A(n9020), .ZN(n9022) );
  NOR4_X1 U10384 ( .A1(n9023), .A2(n9791), .A3(n4480), .A4(n9613), .ZN(n9026)
         );
  OAI21_X1 U10385 ( .B1(n9027), .B2(n9024), .A(P1_B_REG_SCAN_IN), .ZN(n9025)
         );
  MUX2_X1 U10386 ( .A(n9099), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9036), .Z(
        P1_U3585) );
  MUX2_X1 U10387 ( .A(n9028), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9036), .Z(
        P1_U3584) );
  MUX2_X1 U10388 ( .A(n9029), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9036), .Z(
        P1_U3583) );
  MUX2_X1 U10389 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9030), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10390 ( .A(n9186), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9036), .Z(
        P1_U3581) );
  MUX2_X1 U10391 ( .A(n9372), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9036), .Z(
        P1_U3580) );
  MUX2_X1 U10392 ( .A(n9215), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9036), .Z(
        P1_U3579) );
  MUX2_X1 U10393 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9386), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10394 ( .A(n9254), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9036), .Z(
        P1_U3577) );
  MUX2_X1 U10395 ( .A(n9385), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9036), .Z(
        P1_U3576) );
  MUX2_X1 U10396 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9106), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10397 ( .A(n9415), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9036), .Z(
        P1_U3574) );
  MUX2_X1 U10398 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9324), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10399 ( .A(n9414), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9036), .Z(
        P1_U3572) );
  MUX2_X1 U10400 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9442), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10401 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9031), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10402 ( .A(n9441), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9036), .Z(
        P1_U3569) );
  MUX2_X1 U10403 ( .A(n9032), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9036), .Z(
        P1_U3568) );
  MUX2_X1 U10404 ( .A(n9033), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9036), .Z(
        P1_U3566) );
  MUX2_X1 U10405 ( .A(n9034), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9036), .Z(
        P1_U3564) );
  MUX2_X1 U10406 ( .A(n9843), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9036), .Z(
        P1_U3562) );
  MUX2_X1 U10407 ( .A(n9855), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9036), .Z(
        P1_U3561) );
  MUX2_X1 U10408 ( .A(n9844), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9036), .Z(
        P1_U3560) );
  MUX2_X1 U10409 ( .A(n9035), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9036), .Z(
        P1_U3559) );
  MUX2_X1 U10410 ( .A(n9773), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9036), .Z(
        P1_U3558) );
  MUX2_X1 U10411 ( .A(n7151), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9036), .Z(
        P1_U3557) );
  MUX2_X1 U10412 ( .A(n9794), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9036), .Z(
        P1_U3556) );
  AOI211_X1 U10413 ( .C1(n9039), .C2(n9038), .A(n9037), .B(n9682), .ZN(n9049)
         );
  AOI211_X1 U10414 ( .C1(n9042), .C2(n9041), .A(n9040), .B(n9623), .ZN(n9048)
         );
  NAND2_X1 U10415 ( .A1(n9690), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9045) );
  INV_X1 U10416 ( .A(n9043), .ZN(n9044) );
  OAI211_X1 U10417 ( .C1(n9715), .C2(n9046), .A(n9045), .B(n9044), .ZN(n9047)
         );
  OR3_X1 U10418 ( .A1(n9049), .A2(n9048), .A3(n9047), .ZN(P1_U3257) );
  AOI211_X1 U10419 ( .C1(n9052), .C2(n9051), .A(n9050), .B(n9682), .ZN(n9061)
         );
  AOI211_X1 U10420 ( .C1(n9055), .C2(n9054), .A(n9053), .B(n9623), .ZN(n9060)
         );
  NAND2_X1 U10421 ( .A1(n9690), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9057) );
  NAND2_X1 U10422 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n9056) );
  OAI211_X1 U10423 ( .C1(n9715), .C2(n9058), .A(n9057), .B(n9056), .ZN(n9059)
         );
  OR3_X1 U10424 ( .A1(n9061), .A2(n9060), .A3(n9059), .ZN(P1_U3258) );
  NAND2_X1 U10425 ( .A1(n9173), .A2(n9466), .ZN(n9159) );
  NAND2_X1 U10426 ( .A1(n9062), .A2(n9785), .ZN(n9332) );
  NOR2_X1 U10427 ( .A1(n9222), .A2(n9063), .ZN(n9067) );
  NAND2_X1 U10428 ( .A1(n9064), .A2(P1_B_REG_SCAN_IN), .ZN(n9065) );
  AND2_X1 U10429 ( .A1(n9857), .A2(n9065), .ZN(n9100) );
  NAND2_X1 U10430 ( .A1(n9066), .A2(n9100), .ZN(n9335) );
  NOR2_X1 U10431 ( .A1(n9779), .A2(n9335), .ZN(n9073) );
  AOI211_X1 U10432 ( .C1(n9068), .C2(n9572), .A(n9067), .B(n9073), .ZN(n9069)
         );
  OAI21_X1 U10433 ( .B1(n9332), .B2(n9576), .A(n9069), .ZN(P1_U3261) );
  OAI211_X1 U10434 ( .C1(n4774), .C2(n9125), .A(n9785), .B(n9071), .ZN(n9336)
         );
  NOR2_X1 U10435 ( .A1(n4774), .A2(n9781), .ZN(n9072) );
  AOI211_X1 U10436 ( .C1(n9807), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9073), .B(
        n9072), .ZN(n9074) );
  OAI21_X1 U10437 ( .B1(n9576), .B2(n9336), .A(n9074), .ZN(P1_U3262) );
  NAND2_X1 U10438 ( .A1(n9076), .A2(n9075), .ZN(n9078) );
  NAND2_X1 U10439 ( .A1(n9078), .A2(n9077), .ZN(n9314) );
  NAND2_X1 U10440 ( .A1(n9081), .A2(n9080), .ZN(n9082) );
  NAND2_X1 U10441 ( .A1(n9228), .A2(n9229), .ZN(n9090) );
  XNOR2_X1 U10442 ( .A(n9098), .B(n9123), .ZN(n9101) );
  NOR2_X1 U10443 ( .A1(n9317), .A2(n9414), .ZN(n9105) );
  NOR2_X1 U10444 ( .A1(n9108), .A2(n9107), .ZN(n9245) );
  NAND2_X1 U10445 ( .A1(n9476), .A2(n9207), .ZN(n9111) );
  NOR2_X1 U10446 ( .A1(n9476), .A2(n9207), .ZN(n9110) );
  AOI21_X2 U10447 ( .B1(n9219), .B2(n9111), .A(n9110), .ZN(n9199) );
  NAND2_X1 U10448 ( .A1(n9210), .A2(n9215), .ZN(n9112) );
  NAND2_X1 U10449 ( .A1(n9199), .A2(n9112), .ZN(n9115) );
  NAND2_X1 U10450 ( .A1(n9375), .A2(n9113), .ZN(n9114) );
  NAND2_X1 U10451 ( .A1(n9115), .A2(n9114), .ZN(n9180) );
  NAND2_X1 U10452 ( .A1(n9180), .A2(n9181), .ZN(n9117) );
  NAND2_X1 U10453 ( .A1(n9117), .A2(n9116), .ZN(n9166) );
  INV_X1 U10454 ( .A(n9166), .ZN(n9121) );
  INV_X1 U10455 ( .A(n9118), .ZN(n9120) );
  OAI21_X2 U10456 ( .B1(n9121), .B2(n9120), .A(n9119), .ZN(n9156) );
  NAND2_X1 U10457 ( .A1(n9466), .A2(n9172), .ZN(n9122) );
  XNOR2_X1 U10458 ( .A(n9124), .B(n9123), .ZN(n9339) );
  NAND2_X1 U10459 ( .A1(n9339), .A2(n9767), .ZN(n9133) );
  AOI211_X1 U10460 ( .C1(n9126), .C2(n9143), .A(n9749), .B(n9125), .ZN(n9343)
         );
  NOR2_X1 U10461 ( .A1(n9341), .A2(n9781), .ZN(n9131) );
  INV_X1 U10462 ( .A(n9127), .ZN(n9128) );
  AOI22_X1 U10463 ( .A1(n9128), .A2(n9804), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9779), .ZN(n9129) );
  OAI21_X1 U10464 ( .B1(n9356), .B2(n9318), .A(n9129), .ZN(n9130) );
  AOI211_X1 U10465 ( .C1(n9343), .C2(n9787), .A(n9131), .B(n9130), .ZN(n9132)
         );
  OAI211_X1 U10466 ( .C1(n9340), .C2(n9779), .A(n9133), .B(n9132), .ZN(
        P1_U3355) );
  XNOR2_X1 U10467 ( .A(n9134), .B(n5076), .ZN(n9136) );
  NOR2_X1 U10468 ( .A1(n9172), .A2(n9757), .ZN(n9135) );
  AOI21_X1 U10469 ( .B1(n9136), .B2(n9427), .A(n9135), .ZN(n9346) );
  NAND2_X1 U10470 ( .A1(n9138), .A2(n9137), .ZN(n9139) );
  NAND2_X1 U10471 ( .A1(n9349), .A2(n9767), .ZN(n9148) );
  AOI22_X1 U10472 ( .A1(n9141), .A2(n9804), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9779), .ZN(n9142) );
  OAI21_X1 U10473 ( .B1(n9347), .B2(n9203), .A(n9142), .ZN(n9146) );
  INV_X1 U10474 ( .A(n9159), .ZN(n9144) );
  OAI211_X1 U10475 ( .C1(n9462), .C2(n9144), .A(n9785), .B(n9143), .ZN(n9345)
         );
  NOR2_X1 U10476 ( .A1(n9345), .A2(n9576), .ZN(n9145) );
  AOI211_X1 U10477 ( .C1(n9572), .C2(n9352), .A(n9146), .B(n9145), .ZN(n9147)
         );
  OAI211_X1 U10478 ( .C1(n9346), .C2(n9779), .A(n9148), .B(n9147), .ZN(
        P1_U3263) );
  OAI211_X1 U10479 ( .C1(n9151), .C2(n9150), .A(n9149), .B(n9427), .ZN(n9152)
         );
  INV_X1 U10480 ( .A(n9358), .ZN(n9165) );
  OAI21_X1 U10481 ( .B1(n9156), .B2(n9155), .A(n9154), .ZN(n9359) );
  NAND2_X1 U10482 ( .A1(n9359), .A2(n9767), .ZN(n9164) );
  AOI22_X1 U10483 ( .A1(n9157), .A2(n9804), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9779), .ZN(n9158) );
  OAI21_X1 U10484 ( .B1(n9356), .B2(n9203), .A(n9158), .ZN(n9161) );
  OAI211_X1 U10485 ( .C1(n9466), .C2(n9173), .A(n9785), .B(n9159), .ZN(n9355)
         );
  NOR2_X1 U10486 ( .A1(n9355), .A2(n9576), .ZN(n9160) );
  AOI211_X1 U10487 ( .C1(n9572), .C2(n9162), .A(n9161), .B(n9160), .ZN(n9163)
         );
  OAI211_X1 U10488 ( .C1(n9807), .C2(n9165), .A(n9164), .B(n9163), .ZN(
        P1_U3264) );
  XNOR2_X1 U10489 ( .A(n9166), .B(n9169), .ZN(n9366) );
  NAND2_X1 U10490 ( .A1(n9168), .A2(n9167), .ZN(n9170) );
  XNOR2_X1 U10491 ( .A(n9170), .B(n9169), .ZN(n9171) );
  OAI222_X1 U10492 ( .A1(n9735), .A2(n9172), .B1(n9757), .B2(n9204), .C1(n9171), .C2(n9862), .ZN(n9362) );
  AOI211_X1 U10493 ( .C1(n9364), .C2(n9190), .A(n9749), .B(n9173), .ZN(n9363)
         );
  NAND2_X1 U10494 ( .A1(n9363), .A2(n9787), .ZN(n9176) );
  AOI22_X1 U10495 ( .A1(n9174), .A2(n9804), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9779), .ZN(n9175) );
  OAI211_X1 U10496 ( .C1(n9177), .C2(n9781), .A(n9176), .B(n9175), .ZN(n9178)
         );
  AOI21_X1 U10497 ( .B1(n9362), .B2(n9222), .A(n9178), .ZN(n9179) );
  OAI21_X1 U10498 ( .B1(n9366), .B2(n9331), .A(n9179), .ZN(P1_U3265) );
  XNOR2_X1 U10499 ( .A(n9180), .B(n9181), .ZN(n9369) );
  INV_X1 U10500 ( .A(n9369), .ZN(n9198) );
  NAND2_X1 U10501 ( .A1(n9200), .A2(n9182), .ZN(n9184) );
  XNOR2_X1 U10502 ( .A(n9184), .B(n9183), .ZN(n9185) );
  NAND2_X1 U10503 ( .A1(n9185), .A2(n9427), .ZN(n9188) );
  AOI22_X1 U10504 ( .A1(n9186), .A2(n9857), .B1(n9856), .B2(n9215), .ZN(n9187)
         );
  NAND2_X1 U10505 ( .A1(n9188), .A2(n9187), .ZN(n9367) );
  INV_X1 U10506 ( .A(n9189), .ZN(n9202) );
  INV_X1 U10507 ( .A(n9190), .ZN(n9191) );
  AOI211_X1 U10508 ( .C1(n9192), .C2(n9202), .A(n9749), .B(n9191), .ZN(n9368)
         );
  NAND2_X1 U10509 ( .A1(n9368), .A2(n9787), .ZN(n9195) );
  AOI22_X1 U10510 ( .A1(n9193), .A2(n9804), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9779), .ZN(n9194) );
  OAI211_X1 U10511 ( .C1(n9471), .C2(n9781), .A(n9195), .B(n9194), .ZN(n9196)
         );
  AOI21_X1 U10512 ( .B1(n9367), .B2(n9222), .A(n9196), .ZN(n9197) );
  OAI21_X1 U10513 ( .B1(n9198), .B2(n9331), .A(n9197), .ZN(P1_U3266) );
  XNOR2_X1 U10514 ( .A(n9199), .B(n9201), .ZN(n9379) );
  OAI21_X1 U10515 ( .B1(n4515), .B2(n9201), .A(n9200), .ZN(n9377) );
  OAI211_X1 U10516 ( .C1(n9375), .C2(n4551), .A(n9202), .B(n9785), .ZN(n9374)
         );
  NAND2_X1 U10517 ( .A1(n9222), .A2(n9761), .ZN(n9249) );
  NOR2_X1 U10518 ( .A1(n9204), .A2(n9203), .ZN(n9209) );
  AOI22_X1 U10519 ( .A1(n9205), .A2(n9804), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9779), .ZN(n9206) );
  OAI21_X1 U10520 ( .B1(n9207), .B2(n9318), .A(n9206), .ZN(n9208) );
  AOI211_X1 U10521 ( .C1(n9210), .C2(n9572), .A(n9209), .B(n9208), .ZN(n9211)
         );
  OAI21_X1 U10522 ( .B1(n9374), .B2(n9249), .A(n9211), .ZN(n9212) );
  AOI21_X1 U10523 ( .B1(n9377), .B2(n9329), .A(n9212), .ZN(n9213) );
  OAI21_X1 U10524 ( .B1(n9379), .B2(n9331), .A(n9213), .ZN(P1_U3267) );
  OAI211_X1 U10525 ( .C1(n4519), .C2(n4824), .A(n9427), .B(n9214), .ZN(n9217)
         );
  AOI22_X1 U10526 ( .A1(n9215), .A2(n9857), .B1(n9856), .B2(n9254), .ZN(n9216)
         );
  NAND2_X1 U10527 ( .A1(n9217), .A2(n9216), .ZN(n9380) );
  AOI21_X1 U10528 ( .B1(n9218), .B2(n9804), .A(n9380), .ZN(n9227) );
  XOR2_X1 U10529 ( .A(n9219), .B(n9220), .Z(n9382) );
  NAND2_X1 U10530 ( .A1(n9382), .A2(n9767), .ZN(n9226) );
  AOI211_X1 U10531 ( .C1(n9221), .C2(n9235), .A(n9749), .B(n4551), .ZN(n9381)
         );
  INV_X1 U10532 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9223) );
  OAI22_X1 U10533 ( .A1(n9476), .A2(n9781), .B1(n9223), .B2(n9222), .ZN(n9224)
         );
  AOI21_X1 U10534 ( .B1(n9381), .B2(n9787), .A(n9224), .ZN(n9225) );
  OAI211_X1 U10535 ( .C1(n9807), .C2(n9227), .A(n9226), .B(n9225), .ZN(
        P1_U3268) );
  XOR2_X1 U10536 ( .A(n9229), .B(n9228), .Z(n9389) );
  XNOR2_X1 U10537 ( .A(n9230), .B(n9229), .ZN(n9391) );
  NAND2_X1 U10538 ( .A1(n9391), .A2(n9767), .ZN(n9241) );
  NAND2_X1 U10539 ( .A1(n9386), .A2(n9325), .ZN(n9234) );
  INV_X1 U10540 ( .A(n9231), .ZN(n9232) );
  AOI22_X1 U10541 ( .A1(n9232), .A2(n9804), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9779), .ZN(n9233) );
  OAI211_X1 U10542 ( .C1(n9266), .C2(n9318), .A(n9234), .B(n9233), .ZN(n9238)
         );
  AOI21_X1 U10543 ( .B1(n9246), .B2(n9239), .A(n9749), .ZN(n9236) );
  NAND2_X1 U10544 ( .A1(n9236), .A2(n9235), .ZN(n9387) );
  NOR2_X1 U10545 ( .A1(n9387), .A2(n9576), .ZN(n9237) );
  AOI211_X1 U10546 ( .C1(n9572), .C2(n9239), .A(n9238), .B(n9237), .ZN(n9240)
         );
  OAI211_X1 U10547 ( .C1(n9310), .C2(n9389), .A(n9241), .B(n9240), .ZN(
        P1_U3269) );
  XNOR2_X1 U10548 ( .A(n9243), .B(n9242), .ZN(n9403) );
  OR2_X1 U10549 ( .A1(n9245), .A2(n9244), .ZN(n9395) );
  NAND3_X1 U10550 ( .A1(n9395), .A2(n9394), .A3(n9767), .ZN(n9260) );
  INV_X1 U10551 ( .A(n9267), .ZN(n9248) );
  INV_X1 U10552 ( .A(n9246), .ZN(n9247) );
  AOI211_X1 U10553 ( .C1(n9400), .C2(n9248), .A(n9749), .B(n9247), .ZN(n9398)
         );
  INV_X1 U10554 ( .A(n9249), .ZN(n9258) );
  INV_X1 U10555 ( .A(n9250), .ZN(n9251) );
  AOI22_X1 U10556 ( .A1(n9251), .A2(n9804), .B1(n9807), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9252) );
  OAI21_X1 U10557 ( .B1(n9396), .B2(n9318), .A(n9252), .ZN(n9253) );
  AOI21_X1 U10558 ( .B1(n9325), .B2(n9254), .A(n9253), .ZN(n9255) );
  OAI21_X1 U10559 ( .B1(n9256), .B2(n9781), .A(n9255), .ZN(n9257) );
  AOI21_X1 U10560 ( .B1(n9398), .B2(n9258), .A(n9257), .ZN(n9259) );
  OAI211_X1 U10561 ( .C1(n9403), .C2(n9310), .A(n9260), .B(n9259), .ZN(
        P1_U3270) );
  XNOR2_X1 U10562 ( .A(n9261), .B(n9262), .ZN(n9408) );
  XNOR2_X1 U10563 ( .A(n9263), .B(n9262), .ZN(n9264) );
  OAI222_X1 U10564 ( .A1(n9735), .A2(n9266), .B1(n9757), .B2(n9265), .C1(n9264), .C2(n9862), .ZN(n9404) );
  INV_X1 U10565 ( .A(n9282), .ZN(n9268) );
  AOI211_X1 U10566 ( .C1(n9406), .C2(n9268), .A(n9749), .B(n9267), .ZN(n9405)
         );
  NAND2_X1 U10567 ( .A1(n9405), .A2(n9787), .ZN(n9271) );
  AOI22_X1 U10568 ( .A1(n9779), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9269), .B2(
        n9804), .ZN(n9270) );
  OAI211_X1 U10569 ( .C1(n9272), .C2(n9781), .A(n9271), .B(n9270), .ZN(n9273)
         );
  AOI21_X1 U10570 ( .B1(n9404), .B2(n9222), .A(n9273), .ZN(n9274) );
  OAI21_X1 U10571 ( .B1(n9408), .B2(n9331), .A(n9274), .ZN(P1_U3271) );
  INV_X1 U10572 ( .A(n9275), .ZN(n9276) );
  AOI21_X1 U10573 ( .B1(n9277), .B2(n9279), .A(n9276), .ZN(n9278) );
  OAI222_X1 U10574 ( .A1(n9735), .A2(n9396), .B1(n9757), .B2(n9424), .C1(n9862), .C2(n9278), .ZN(n9409) );
  INV_X1 U10575 ( .A(n9409), .ZN(n9290) );
  XNOR2_X1 U10576 ( .A(n9280), .B(n9279), .ZN(n9411) );
  NAND2_X1 U10577 ( .A1(n9411), .A2(n9767), .ZN(n9289) );
  INV_X1 U10578 ( .A(n9281), .ZN(n9304) );
  AOI211_X1 U10579 ( .C1(n9283), .C2(n9304), .A(n9749), .B(n9282), .ZN(n9410)
         );
  NOR2_X1 U10580 ( .A1(n9486), .A2(n9781), .ZN(n9287) );
  OAI22_X1 U10581 ( .A1(n9222), .A2(n9285), .B1(n9284), .B2(n9319), .ZN(n9286)
         );
  AOI211_X1 U10582 ( .C1(n9410), .C2(n9787), .A(n9287), .B(n9286), .ZN(n9288)
         );
  OAI211_X1 U10583 ( .C1(n9807), .C2(n9290), .A(n9289), .B(n9288), .ZN(
        P1_U3272) );
  INV_X1 U10584 ( .A(n9291), .ZN(n9293) );
  OAI21_X1 U10585 ( .B1(n9314), .B2(n9293), .A(n9292), .ZN(n9295) );
  INV_X1 U10586 ( .A(n9296), .ZN(n9294) );
  XNOR2_X1 U10587 ( .A(n9295), .B(n9294), .ZN(n9418) );
  XOR2_X1 U10588 ( .A(n9297), .B(n9296), .Z(n9420) );
  NAND2_X1 U10589 ( .A1(n9420), .A2(n9767), .ZN(n9309) );
  OAI22_X1 U10590 ( .A1(n9222), .A2(n9299), .B1(n9298), .B2(n9319), .ZN(n9300)
         );
  AOI21_X1 U10591 ( .B1(n9325), .B2(n9415), .A(n9300), .ZN(n9301) );
  OAI21_X1 U10592 ( .B1(n9302), .B2(n9318), .A(n9301), .ZN(n9306) );
  INV_X1 U10593 ( .A(n9303), .ZN(n9315) );
  OAI211_X1 U10594 ( .C1(n9490), .C2(n9315), .A(n9304), .B(n9785), .ZN(n9416)
         );
  NOR2_X1 U10595 ( .A1(n9416), .A2(n9576), .ZN(n9305) );
  AOI211_X1 U10596 ( .C1(n9572), .C2(n9307), .A(n9306), .B(n9305), .ZN(n9308)
         );
  OAI211_X1 U10597 ( .C1(n9418), .C2(n9310), .A(n9309), .B(n9308), .ZN(
        P1_U3273) );
  XNOR2_X1 U10598 ( .A(n9312), .B(n9313), .ZN(n9430) );
  XNOR2_X1 U10599 ( .A(n9314), .B(n9313), .ZN(n9428) );
  AOI211_X1 U10600 ( .C1(n9317), .C2(n9316), .A(n9749), .B(n9315), .ZN(n9425)
         );
  NAND2_X1 U10601 ( .A1(n9425), .A2(n9787), .ZN(n9327) );
  NOR2_X1 U10602 ( .A1(n9318), .A2(n9423), .ZN(n9323) );
  OAI22_X1 U10603 ( .A1(n9222), .A2(n9321), .B1(n9320), .B2(n9319), .ZN(n9322)
         );
  AOI211_X1 U10604 ( .C1(n9325), .C2(n9324), .A(n9323), .B(n9322), .ZN(n9326)
         );
  OAI211_X1 U10605 ( .C1(n4769), .C2(n9781), .A(n9327), .B(n9326), .ZN(n9328)
         );
  AOI21_X1 U10606 ( .B1(n9329), .B2(n9428), .A(n9328), .ZN(n9330) );
  OAI21_X1 U10607 ( .B1(n9430), .B2(n9331), .A(n9330), .ZN(P1_U3274) );
  INV_X1 U10608 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9333) );
  MUX2_X1 U10609 ( .A(n9333), .B(n9451), .S(n9902), .Z(n9334) );
  OAI21_X1 U10610 ( .B1(n9454), .B2(n9434), .A(n9334), .ZN(P1_U3554) );
  AND2_X1 U10611 ( .A1(n9336), .A2(n9335), .ZN(n9455) );
  MUX2_X1 U10612 ( .A(n9337), .B(n9455), .S(n9902), .Z(n9338) );
  OAI21_X1 U10613 ( .B1(n4774), .B2(n9434), .A(n9338), .ZN(P1_U3553) );
  NAND2_X1 U10614 ( .A1(n9339), .A2(n9867), .ZN(n9344) );
  OAI22_X1 U10615 ( .A1(n9341), .A2(n9869), .B1(n9356), .B2(n9757), .ZN(n9342)
         );
  MUX2_X1 U10616 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9458), .S(n9902), .Z(
        P1_U3552) );
  OAI211_X1 U10617 ( .C1(n9347), .C2(n9735), .A(n9346), .B(n9345), .ZN(n9348)
         );
  MUX2_X1 U10618 ( .A(n9350), .B(n9459), .S(n9902), .Z(n9354) );
  NAND2_X1 U10619 ( .A1(n9352), .A2(n9351), .ZN(n9353) );
  NAND2_X1 U10620 ( .A1(n9354), .A2(n9353), .ZN(P1_U3551) );
  OAI21_X1 U10621 ( .B1(n9356), .B2(n9735), .A(n9355), .ZN(n9357) );
  AOI211_X1 U10622 ( .C1(n9359), .C2(n9867), .A(n9358), .B(n9357), .ZN(n9463)
         );
  MUX2_X1 U10623 ( .A(n9360), .B(n9463), .S(n9902), .Z(n9361) );
  OAI21_X1 U10624 ( .B1(n9466), .B2(n9434), .A(n9361), .ZN(P1_U3550) );
  INV_X1 U10625 ( .A(n9867), .ZN(n9439) );
  AOI211_X1 U10626 ( .C1(n9880), .C2(n9364), .A(n9363), .B(n9362), .ZN(n9365)
         );
  OAI21_X1 U10627 ( .B1(n9366), .B2(n9439), .A(n9365), .ZN(n9467) );
  MUX2_X1 U10628 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9467), .S(n9902), .Z(
        P1_U3549) );
  AOI211_X1 U10629 ( .C1(n9369), .C2(n9867), .A(n9368), .B(n9367), .ZN(n9468)
         );
  MUX2_X1 U10630 ( .A(n9370), .B(n9468), .S(n9902), .Z(n9371) );
  OAI21_X1 U10631 ( .B1(n9471), .B2(n9434), .A(n9371), .ZN(P1_U3548) );
  AOI22_X1 U10632 ( .A1(n9372), .A2(n9857), .B1(n9856), .B2(n9386), .ZN(n9373)
         );
  OAI211_X1 U10633 ( .C1(n9375), .C2(n9869), .A(n9374), .B(n9373), .ZN(n9376)
         );
  AOI21_X1 U10634 ( .B1(n9377), .B2(n9427), .A(n9376), .ZN(n9378) );
  OAI21_X1 U10635 ( .B1(n9379), .B2(n9439), .A(n9378), .ZN(n9472) );
  MUX2_X1 U10636 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9472), .S(n9902), .Z(
        P1_U3547) );
  MUX2_X1 U10637 ( .A(n9383), .B(n9473), .S(n9902), .Z(n9384) );
  OAI21_X1 U10638 ( .B1(n9476), .B2(n9434), .A(n9384), .ZN(P1_U3546) );
  AOI22_X1 U10639 ( .A1(n9386), .A2(n9857), .B1(n9856), .B2(n9385), .ZN(n9388)
         );
  OAI211_X1 U10640 ( .C1(n9389), .C2(n9862), .A(n9388), .B(n9387), .ZN(n9390)
         );
  AOI21_X1 U10641 ( .B1(n9391), .B2(n9867), .A(n9390), .ZN(n9477) );
  MUX2_X1 U10642 ( .A(n9392), .B(n9477), .S(n9902), .Z(n9393) );
  OAI21_X1 U10643 ( .B1(n9480), .B2(n9434), .A(n9393), .ZN(P1_U3545) );
  NAND3_X1 U10644 ( .A1(n9395), .A2(n9394), .A3(n9867), .ZN(n9402) );
  OAI22_X1 U10645 ( .A1(n9397), .A2(n9735), .B1(n9396), .B2(n9757), .ZN(n9399)
         );
  AOI211_X1 U10646 ( .C1(n9880), .C2(n9400), .A(n9399), .B(n9398), .ZN(n9401)
         );
  OAI211_X1 U10647 ( .C1(n9862), .C2(n9403), .A(n9402), .B(n9401), .ZN(n9481)
         );
  MUX2_X1 U10648 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9481), .S(n9902), .Z(
        P1_U3544) );
  AOI211_X1 U10649 ( .C1(n9880), .C2(n9406), .A(n9405), .B(n9404), .ZN(n9407)
         );
  OAI21_X1 U10650 ( .B1(n9408), .B2(n9439), .A(n9407), .ZN(n9482) );
  MUX2_X1 U10651 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9482), .S(n9902), .Z(
        P1_U3543) );
  AOI211_X1 U10652 ( .C1(n9411), .C2(n9867), .A(n9410), .B(n9409), .ZN(n9483)
         );
  MUX2_X1 U10653 ( .A(n9412), .B(n9483), .S(n9902), .Z(n9413) );
  OAI21_X1 U10654 ( .B1(n9486), .B2(n9434), .A(n9413), .ZN(P1_U3542) );
  AOI22_X1 U10655 ( .A1(n9415), .A2(n9857), .B1(n9414), .B2(n9856), .ZN(n9417)
         );
  OAI211_X1 U10656 ( .C1(n9418), .C2(n9862), .A(n9417), .B(n9416), .ZN(n9419)
         );
  AOI21_X1 U10657 ( .B1(n9420), .B2(n9867), .A(n9419), .ZN(n9487) );
  MUX2_X1 U10658 ( .A(n9421), .B(n9487), .S(n9902), .Z(n9422) );
  OAI21_X1 U10659 ( .B1(n9490), .B2(n9434), .A(n9422), .ZN(P1_U3541) );
  OAI22_X1 U10660 ( .A1(n9424), .A2(n9735), .B1(n9423), .B2(n9757), .ZN(n9426)
         );
  AOI211_X1 U10661 ( .C1(n9428), .C2(n9427), .A(n9426), .B(n9425), .ZN(n9429)
         );
  OAI21_X1 U10662 ( .B1(n9430), .B2(n9439), .A(n9429), .ZN(n9491) );
  INV_X1 U10663 ( .A(n9491), .ZN(n9431) );
  MUX2_X1 U10664 ( .A(n9432), .B(n9431), .S(n9902), .Z(n9433) );
  OAI21_X1 U10665 ( .B1(n4769), .B2(n9434), .A(n9433), .ZN(P1_U3540) );
  AOI211_X1 U10666 ( .C1(n9880), .C2(n9437), .A(n9436), .B(n9435), .ZN(n9438)
         );
  OAI21_X1 U10667 ( .B1(n9440), .B2(n9439), .A(n9438), .ZN(n9495) );
  MUX2_X1 U10668 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9495), .S(n9902), .Z(
        P1_U3539) );
  AOI22_X1 U10669 ( .A1(n9442), .A2(n9857), .B1(n9856), .B2(n9441), .ZN(n9445)
         );
  NAND2_X1 U10670 ( .A1(n9443), .A2(n9880), .ZN(n9444) );
  NAND3_X1 U10671 ( .A1(n9446), .A2(n9445), .A3(n9444), .ZN(n9447) );
  AOI211_X1 U10672 ( .C1(n9449), .C2(n9867), .A(n9448), .B(n9447), .ZN(n9450)
         );
  INV_X1 U10673 ( .A(n9450), .ZN(n9496) );
  MUX2_X1 U10674 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9496), .S(n9902), .Z(
        P1_U3538) );
  MUX2_X1 U10675 ( .A(n9452), .B(n9451), .S(n9888), .Z(n9453) );
  OAI21_X1 U10676 ( .B1(n9454), .B2(n9494), .A(n9453), .ZN(P1_U3522) );
  INV_X1 U10677 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9456) );
  MUX2_X1 U10678 ( .A(n9456), .B(n9455), .S(n9888), .Z(n9457) );
  OAI21_X1 U10679 ( .B1(n4774), .B2(n9494), .A(n9457), .ZN(P1_U3521) );
  MUX2_X1 U10680 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9458), .S(n9888), .Z(
        P1_U3520) );
  INV_X1 U10681 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9460) );
  OAI21_X1 U10682 ( .B1(n9462), .B2(n9494), .A(n9461), .ZN(P1_U3519) );
  INV_X1 U10683 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9464) );
  MUX2_X1 U10684 ( .A(n9464), .B(n9463), .S(n9888), .Z(n9465) );
  OAI21_X1 U10685 ( .B1(n9466), .B2(n9494), .A(n9465), .ZN(P1_U3518) );
  MUX2_X1 U10686 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9467), .S(n9888), .Z(
        P1_U3517) );
  INV_X1 U10687 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9469) );
  MUX2_X1 U10688 ( .A(n9469), .B(n9468), .S(n9888), .Z(n9470) );
  OAI21_X1 U10689 ( .B1(n9471), .B2(n9494), .A(n9470), .ZN(P1_U3516) );
  MUX2_X1 U10690 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9472), .S(n9888), .Z(
        P1_U3515) );
  INV_X1 U10691 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9474) );
  MUX2_X1 U10692 ( .A(n9474), .B(n9473), .S(n9888), .Z(n9475) );
  OAI21_X1 U10693 ( .B1(n9476), .B2(n9494), .A(n9475), .ZN(P1_U3514) );
  INV_X1 U10694 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9478) );
  MUX2_X1 U10695 ( .A(n9478), .B(n9477), .S(n9888), .Z(n9479) );
  OAI21_X1 U10696 ( .B1(n9480), .B2(n9494), .A(n9479), .ZN(P1_U3513) );
  MUX2_X1 U10697 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9481), .S(n9888), .Z(
        P1_U3512) );
  MUX2_X1 U10698 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9482), .S(n9888), .Z(
        P1_U3511) );
  INV_X1 U10699 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9484) );
  MUX2_X1 U10700 ( .A(n9484), .B(n9483), .S(n9888), .Z(n9485) );
  OAI21_X1 U10701 ( .B1(n9486), .B2(n9494), .A(n9485), .ZN(P1_U3510) );
  INV_X1 U10702 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9488) );
  MUX2_X1 U10703 ( .A(n9488), .B(n9487), .S(n9888), .Z(n9489) );
  OAI21_X1 U10704 ( .B1(n9490), .B2(n9494), .A(n9489), .ZN(P1_U3508) );
  MUX2_X1 U10705 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9491), .S(n9888), .Z(n9492) );
  INV_X1 U10706 ( .A(n9492), .ZN(n9493) );
  OAI21_X1 U10707 ( .B1(n4769), .B2(n9494), .A(n9493), .ZN(P1_U3505) );
  MUX2_X1 U10708 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9495), .S(n9888), .Z(
        P1_U3502) );
  MUX2_X1 U10709 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9496), .S(n9888), .Z(
        P1_U3499) );
  NAND3_X1 U10710 ( .A1(n9498), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n9500) );
  OAI22_X1 U10711 ( .A1(n9497), .A2(n9500), .B1(n10261), .B2(n9499), .ZN(n9501) );
  AOI21_X1 U10712 ( .B1(n9503), .B2(n9502), .A(n9501), .ZN(n9504) );
  INV_X1 U10713 ( .A(n9504), .ZN(P1_U3322) );
  MUX2_X1 U10714 ( .A(n9505), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI22_X1 U10715 ( .A1(n9909), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n9521) );
  INV_X1 U10716 ( .A(n9506), .ZN(n9507) );
  NAND2_X1 U10717 ( .A1(n9527), .A2(n9507), .ZN(n9519) );
  NAND2_X1 U10718 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9508) );
  AND2_X1 U10719 ( .A1(n9509), .A2(n9508), .ZN(n9510) );
  OR3_X1 U10720 ( .A1(n9907), .A2(n9511), .A3(n9510), .ZN(n9518) );
  INV_X1 U10721 ( .A(n9512), .ZN(n9516) );
  NAND2_X1 U10722 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9513) );
  NAND2_X1 U10723 ( .A1(n9514), .A2(n9513), .ZN(n9515) );
  NAND3_X1 U10724 ( .A1(n9904), .A2(n9516), .A3(n9515), .ZN(n9517) );
  AND3_X1 U10725 ( .A1(n9519), .A2(n9518), .A3(n9517), .ZN(n9520) );
  NAND2_X1 U10726 ( .A1(n9521), .A2(n9520), .ZN(P2_U3246) );
  AOI22_X1 U10727 ( .A1(n9909), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9537) );
  INV_X1 U10728 ( .A(n9523), .ZN(n9524) );
  OAI21_X1 U10729 ( .B1(n9525), .B2(n4786), .A(n9524), .ZN(n9534) );
  NAND2_X1 U10730 ( .A1(n9527), .A2(n9526), .ZN(n9533) );
  AOI21_X1 U10731 ( .B1(n9530), .B2(n9529), .A(n9528), .ZN(n9531) );
  NAND2_X1 U10732 ( .A1(n9904), .A2(n9531), .ZN(n9532) );
  OAI211_X1 U10733 ( .C1(n9534), .C2(n9907), .A(n9533), .B(n9532), .ZN(n9535)
         );
  INV_X1 U10734 ( .A(n9535), .ZN(n9536) );
  NAND2_X1 U10735 ( .A1(n9537), .A2(n9536), .ZN(P2_U3247) );
  OAI22_X1 U10736 ( .A1(n9539), .A2(n10036), .B1(n9538), .B2(n10034), .ZN(
        n9541) );
  AOI211_X1 U10737 ( .C1(n10041), .C2(n9542), .A(n9541), .B(n9540), .ZN(n9555)
         );
  AOI22_X1 U10738 ( .A1(n10064), .A2(n9555), .B1(n5483), .B2(n10062), .ZN(
        P2_U3535) );
  OAI22_X1 U10739 ( .A1(n9543), .A2(n10036), .B1(n4880), .B2(n10034), .ZN(
        n9545) );
  AOI211_X1 U10740 ( .C1(n10041), .C2(n9546), .A(n9545), .B(n9544), .ZN(n9557)
         );
  AOI22_X1 U10741 ( .A1(n10064), .A2(n9557), .B1(n5453), .B2(n10062), .ZN(
        P2_U3534) );
  NOR2_X1 U10742 ( .A1(n9547), .A2(n9995), .ZN(n9553) );
  OAI22_X1 U10743 ( .A1(n9549), .A2(n10036), .B1(n9548), .B2(n10034), .ZN(
        n9551) );
  AOI211_X1 U10744 ( .C1(n9553), .C2(n9552), .A(n9551), .B(n9550), .ZN(n9559)
         );
  AOI22_X1 U10745 ( .A1(n10064), .A2(n9559), .B1(n5427), .B2(n10062), .ZN(
        P2_U3533) );
  INV_X1 U10746 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9554) );
  AOI22_X1 U10747 ( .A1(n10043), .A2(n9555), .B1(n9554), .B2(n10042), .ZN(
        P2_U3496) );
  INV_X1 U10748 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9556) );
  AOI22_X1 U10749 ( .A1(n10043), .A2(n9557), .B1(n9556), .B2(n10042), .ZN(
        P2_U3493) );
  INV_X1 U10750 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9558) );
  AOI22_X1 U10751 ( .A1(n10043), .A2(n9559), .B1(n9558), .B2(n10042), .ZN(
        P2_U3490) );
  NOR2_X1 U10752 ( .A1(n9561), .A2(n9560), .ZN(n9562) );
  OR2_X1 U10753 ( .A1(n9563), .A2(n9562), .ZN(n9578) );
  INV_X1 U10754 ( .A(n9578), .ZN(n9596) );
  NAND2_X1 U10755 ( .A1(n9565), .A2(n9564), .ZN(n9566) );
  XNOR2_X1 U10756 ( .A(n9566), .B(n7606), .ZN(n9567) );
  OAI222_X1 U10757 ( .A1(n9757), .A2(n9569), .B1(n9735), .B2(n9568), .C1(n9862), .C2(n9567), .ZN(n9595) );
  AOI21_X1 U10758 ( .B1(n9596), .B2(n9886), .A(n9595), .ZN(n9582) );
  INV_X1 U10759 ( .A(n9570), .ZN(n9571) );
  AOI222_X1 U10760 ( .A1(n9592), .A2(n9572), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n9779), .C1(n9804), .C2(n9571), .ZN(n9581) );
  AOI21_X1 U10761 ( .B1(n9573), .B2(n9592), .A(n9749), .ZN(n9575) );
  NAND2_X1 U10762 ( .A1(n9575), .A2(n9574), .ZN(n9593) );
  OAI22_X1 U10763 ( .A1(n9578), .A2(n9577), .B1(n9576), .B2(n9593), .ZN(n9579)
         );
  INV_X1 U10764 ( .A(n9579), .ZN(n9580) );
  OAI211_X1 U10765 ( .C1(n9807), .C2(n9582), .A(n9581), .B(n9580), .ZN(
        P1_U3279) );
  INV_X1 U10766 ( .A(n9589), .ZN(n9591) );
  OAI22_X1 U10767 ( .A1(n9583), .A2(n9735), .B1(n9597), .B2(n9757), .ZN(n9585)
         );
  AOI211_X1 U10768 ( .C1(n9880), .C2(n9586), .A(n9585), .B(n9584), .ZN(n9588)
         );
  OAI211_X1 U10769 ( .C1(n9589), .C2(n9883), .A(n9588), .B(n9587), .ZN(n9590)
         );
  AOI21_X1 U10770 ( .B1(n9886), .B2(n9591), .A(n9590), .ZN(n9608) );
  INV_X1 U10771 ( .A(n9902), .ZN(n9900) );
  AOI22_X1 U10772 ( .A1(n9902), .A2(n9608), .B1(n7019), .B2(n9900), .ZN(
        P1_U3536) );
  OAI21_X1 U10773 ( .B1(n4763), .B2(n9869), .A(n9593), .ZN(n9594) );
  AOI211_X1 U10774 ( .C1(n9596), .C2(n9867), .A(n9595), .B(n9594), .ZN(n9610)
         );
  AOI22_X1 U10775 ( .A1(n9902), .A2(n9610), .B1(n6889), .B2(n9900), .ZN(
        P1_U3535) );
  OAI22_X1 U10776 ( .A1(n9598), .A2(n9757), .B1(n9597), .B2(n9735), .ZN(n9600)
         );
  AOI211_X1 U10777 ( .C1(n9880), .C2(n9601), .A(n9600), .B(n9599), .ZN(n9603)
         );
  OAI211_X1 U10778 ( .C1(n9604), .C2(n9883), .A(n9603), .B(n9602), .ZN(n9605)
         );
  AOI21_X1 U10779 ( .B1(n9886), .B2(n9606), .A(n9605), .ZN(n9612) );
  AOI22_X1 U10780 ( .A1(n9902), .A2(n9612), .B1(n6894), .B2(n9900), .ZN(
        P1_U3534) );
  INV_X1 U10781 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9607) );
  AOI22_X1 U10782 ( .A1(n9888), .A2(n9608), .B1(n9607), .B2(n9887), .ZN(
        P1_U3493) );
  INV_X1 U10783 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9609) );
  AOI22_X1 U10784 ( .A1(n9888), .A2(n9610), .B1(n9609), .B2(n9887), .ZN(
        P1_U3490) );
  INV_X1 U10785 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9611) );
  AOI22_X1 U10786 ( .A1(n9888), .A2(n9612), .B1(n9611), .B2(n9887), .ZN(
        P1_U3487) );
  XNOR2_X1 U10787 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10788 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  NOR2_X1 U10789 ( .A1(n9613), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9614) );
  OR2_X1 U10790 ( .A1(n4480), .A2(n9614), .ZN(n9615) );
  INV_X1 U10791 ( .A(n9615), .ZN(n9616) );
  MUX2_X1 U10792 ( .A(n9616), .B(n9615), .S(P1_IR_REG_0__SCAN_IN), .Z(n9637)
         );
  NAND2_X1 U10793 ( .A1(n9617), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9619) );
  AOI211_X1 U10794 ( .C1(n5895), .C2(n9638), .A(n9619), .B(n9618), .ZN(n9620)
         );
  AOI22_X1 U10795 ( .A1(n9690), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(n9637), .B2(
        n9620), .ZN(n9622) );
  NAND3_X1 U10796 ( .A1(n9720), .A2(P1_IR_REG_0__SCAN_IN), .A3(n5895), .ZN(
        n9621) );
  OAI211_X1 U10797 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n5863), .A(n9622), .B(
        n9621), .ZN(P1_U3241) );
  INV_X1 U10798 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9640) );
  AOI211_X1 U10799 ( .C1(n9626), .C2(n9625), .A(n9624), .B(n9623), .ZN(n9633)
         );
  OAI21_X1 U10800 ( .B1(n9629), .B2(n9628), .A(n9627), .ZN(n9631) );
  OAI22_X1 U10801 ( .A1(n9682), .A2(n9631), .B1(n9630), .B2(n9715), .ZN(n9632)
         );
  AOI211_X1 U10802 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(P1_U3084), .A(n9633), 
        .B(n9632), .ZN(n9639) );
  OR2_X1 U10803 ( .A1(n9635), .A2(n9634), .ZN(n9636) );
  OAI211_X1 U10804 ( .C1(n9638), .C2(n9637), .A(n9636), .B(P1_U4006), .ZN(
        n9651) );
  OAI211_X1 U10805 ( .C1(n9640), .C2(n9724), .A(n9639), .B(n9651), .ZN(
        P1_U3243) );
  OAI21_X1 U10806 ( .B1(n9643), .B2(n9642), .A(n9641), .ZN(n9644) );
  AOI22_X1 U10807 ( .A1(n9695), .A2(n9645), .B1(n9720), .B2(n9644), .ZN(n9653)
         );
  AOI21_X1 U10808 ( .B1(n9647), .B2(n9646), .A(n4565), .ZN(n9648) );
  NOR2_X1 U10809 ( .A1(n9682), .A2(n9648), .ZN(n9649) );
  AOI211_X1 U10810 ( .C1(P1_ADDR_REG_4__SCAN_IN), .C2(n9690), .A(n9650), .B(
        n9649), .ZN(n9652) );
  NAND3_X1 U10811 ( .A1(n9653), .A2(n9652), .A3(n9651), .ZN(P1_U3245) );
  AOI22_X1 U10812 ( .A1(n9690), .A2(P1_ADDR_REG_6__SCAN_IN), .B1(n9695), .B2(
        n9654), .ZN(n9666) );
  INV_X1 U10813 ( .A(n9655), .ZN(n9665) );
  OAI21_X1 U10814 ( .B1(n9658), .B2(n9657), .A(n9656), .ZN(n9659) );
  NAND2_X1 U10815 ( .A1(n9659), .A2(n9720), .ZN(n9664) );
  OAI211_X1 U10816 ( .C1(n9662), .C2(n9661), .A(n9711), .B(n9660), .ZN(n9663)
         );
  NAND4_X1 U10817 ( .A1(n9666), .A2(n9665), .A3(n9664), .A4(n9663), .ZN(
        P1_U3247) );
  INV_X1 U10818 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10495) );
  AOI211_X1 U10819 ( .C1(n9669), .C2(n9668), .A(n9667), .B(n9682), .ZN(n9670)
         );
  AOI211_X1 U10820 ( .C1(n9695), .C2(n9672), .A(n9671), .B(n9670), .ZN(n9678)
         );
  OAI21_X1 U10821 ( .B1(n9675), .B2(n9674), .A(n9673), .ZN(n9676) );
  NAND2_X1 U10822 ( .A1(n9676), .A2(n9720), .ZN(n9677) );
  OAI211_X1 U10823 ( .C1(n10495), .C2(n9724), .A(n9678), .B(n9677), .ZN(
        P1_U3250) );
  OAI21_X1 U10824 ( .B1(n9681), .B2(n9680), .A(n9679), .ZN(n9688) );
  AOI211_X1 U10825 ( .C1(n9685), .C2(n9684), .A(n9683), .B(n9682), .ZN(n9686)
         );
  AOI211_X1 U10826 ( .C1(n9688), .C2(n9720), .A(n9687), .B(n9686), .ZN(n9692)
         );
  AOI22_X1 U10827 ( .A1(n9690), .A2(P1_ADDR_REG_10__SCAN_IN), .B1(n9695), .B2(
        n9689), .ZN(n9691) );
  NAND2_X1 U10828 ( .A1(n9692), .A2(n9691), .ZN(P1_U3251) );
  INV_X1 U10829 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9706) );
  AOI21_X1 U10830 ( .B1(n9695), .B2(n9694), .A(n9693), .ZN(n9705) );
  OAI21_X1 U10831 ( .B1(n9698), .B2(n9697), .A(n9696), .ZN(n9703) );
  OAI21_X1 U10832 ( .B1(n9701), .B2(n9700), .A(n9699), .ZN(n9702) );
  AOI22_X1 U10833 ( .A1(n9703), .A2(n9720), .B1(n9711), .B2(n9702), .ZN(n9704)
         );
  OAI211_X1 U10834 ( .C1(n9724), .C2(n9706), .A(n9705), .B(n9704), .ZN(
        P1_U3252) );
  INV_X1 U10835 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10506) );
  AOI21_X1 U10836 ( .B1(n9709), .B2(n9708), .A(n9707), .ZN(n9710) );
  NAND2_X1 U10837 ( .A1(n9711), .A2(n9710), .ZN(n9713) );
  OAI211_X1 U10838 ( .C1(n9715), .C2(n9714), .A(n9713), .B(n9712), .ZN(n9716)
         );
  INV_X1 U10839 ( .A(n9716), .ZN(n9723) );
  OAI21_X1 U10840 ( .B1(n9719), .B2(n9718), .A(n9717), .ZN(n9721) );
  NAND2_X1 U10841 ( .A1(n9721), .A2(n9720), .ZN(n9722) );
  OAI211_X1 U10842 ( .C1(n10506), .C2(n9724), .A(n9723), .B(n9722), .ZN(
        P1_U3259) );
  INV_X1 U10843 ( .A(n9726), .ZN(n9727) );
  AOI21_X1 U10844 ( .B1(n9729), .B2(n9725), .A(n9727), .ZN(n9874) );
  INV_X1 U10845 ( .A(n9728), .ZN(n9733) );
  AOI21_X1 U10846 ( .B1(n9731), .B2(n9730), .A(n9729), .ZN(n9732) );
  NOR3_X1 U10847 ( .A1(n9733), .A2(n9732), .A3(n9862), .ZN(n9738) );
  OAI22_X1 U10848 ( .A1(n9736), .A2(n9735), .B1(n9734), .B2(n9757), .ZN(n9737)
         );
  AOI211_X1 U10849 ( .C1(n9874), .C2(n9886), .A(n9738), .B(n9737), .ZN(n9871)
         );
  INV_X1 U10850 ( .A(n9739), .ZN(n9740) );
  AOI22_X1 U10851 ( .A1(n9779), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n9740), .B2(
        n9804), .ZN(n9741) );
  OAI21_X1 U10852 ( .B1(n9781), .B2(n9870), .A(n9741), .ZN(n9742) );
  INV_X1 U10853 ( .A(n9742), .ZN(n9748) );
  INV_X1 U10854 ( .A(n9743), .ZN(n9745) );
  OAI211_X1 U10855 ( .C1(n9745), .C2(n9870), .A(n9785), .B(n9744), .ZN(n9868)
         );
  INV_X1 U10856 ( .A(n9868), .ZN(n9746) );
  AOI22_X1 U10857 ( .A1(n9874), .A2(n9788), .B1(n9787), .B2(n9746), .ZN(n9747)
         );
  OAI211_X1 U10858 ( .C1(n9807), .C2(n9871), .A(n9748), .B(n9747), .ZN(
        P1_U3283) );
  AOI21_X1 U10859 ( .B1(n9784), .B2(n9750), .A(n9749), .ZN(n9752) );
  NAND2_X1 U10860 ( .A1(n9752), .A2(n9751), .ZN(n9838) );
  INV_X1 U10861 ( .A(n9838), .ZN(n9762) );
  NAND2_X1 U10862 ( .A1(n9855), .A2(n9857), .ZN(n9837) );
  NAND2_X1 U10863 ( .A1(n9804), .A2(n9753), .ZN(n9754) );
  OAI211_X1 U10864 ( .C1(n9839), .C2(n9755), .A(n9837), .B(n9754), .ZN(n9760)
         );
  XNOR2_X1 U10865 ( .A(n9756), .B(n9766), .ZN(n9759) );
  OAI22_X1 U10866 ( .A1(n9759), .A2(n9862), .B1(n9758), .B2(n9757), .ZN(n9840)
         );
  AOI211_X1 U10867 ( .C1(n9762), .C2(n9761), .A(n9760), .B(n9840), .ZN(n9769)
         );
  INV_X1 U10868 ( .A(n9763), .ZN(n9764) );
  AOI21_X1 U10869 ( .B1(n9766), .B2(n9765), .A(n9764), .ZN(n9842) );
  AOI22_X1 U10870 ( .A1(n9842), .A2(n9767), .B1(P1_REG2_REG_5__SCAN_IN), .B2(
        n9779), .ZN(n9768) );
  OAI21_X1 U10871 ( .B1(n9807), .B2(n9769), .A(n9768), .ZN(P1_U3286) );
  XNOR2_X1 U10872 ( .A(n9771), .B(n9770), .ZN(n9835) );
  XNOR2_X1 U10873 ( .A(n9772), .B(n9771), .ZN(n9775) );
  AOI22_X1 U10874 ( .A1(n9856), .A2(n9773), .B1(n9844), .B2(n9857), .ZN(n9774)
         );
  OAI21_X1 U10875 ( .B1(n9775), .B2(n9862), .A(n9774), .ZN(n9776) );
  AOI21_X1 U10876 ( .B1(n9886), .B2(n9835), .A(n9776), .ZN(n9832) );
  INV_X1 U10877 ( .A(n9777), .ZN(n9778) );
  AOI22_X1 U10878 ( .A1(n9779), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n9778), .B2(
        n9804), .ZN(n9780) );
  OAI21_X1 U10879 ( .B1(n9781), .B2(n9831), .A(n9780), .ZN(n9782) );
  INV_X1 U10880 ( .A(n9782), .ZN(n9790) );
  OAI211_X1 U10881 ( .C1(n4757), .C2(n9831), .A(n9785), .B(n9784), .ZN(n9830)
         );
  INV_X1 U10882 ( .A(n9830), .ZN(n9786) );
  AOI22_X1 U10883 ( .A1(n9835), .A2(n9788), .B1(n9787), .B2(n9786), .ZN(n9789)
         );
  OAI211_X1 U10884 ( .C1(n9807), .C2(n9832), .A(n9790), .B(n9789), .ZN(
        P1_U3287) );
  NAND2_X1 U10885 ( .A1(n9791), .A2(n9797), .ZN(n9792) );
  OR2_X1 U10886 ( .A1(n9793), .A2(n9792), .ZN(n9796) );
  NAND2_X1 U10887 ( .A1(n9794), .A2(n9857), .ZN(n9795) );
  AND2_X1 U10888 ( .A1(n9796), .A2(n9795), .ZN(n9801) );
  INV_X1 U10889 ( .A(n9801), .ZN(n9803) );
  INV_X1 U10890 ( .A(n9797), .ZN(n9798) );
  NAND2_X1 U10891 ( .A1(n9799), .A2(n9798), .ZN(n9800) );
  AND2_X1 U10892 ( .A1(n9801), .A2(n9800), .ZN(n9889) );
  INV_X1 U10893 ( .A(n9889), .ZN(n9802) );
  OAI21_X1 U10894 ( .B1(n9803), .B2(n9883), .A(n9802), .ZN(n9806) );
  AOI22_X1 U10895 ( .A1(n9804), .A2(P1_REG3_REG_0__SCAN_IN), .B1(
        P1_REG2_REG_0__SCAN_IN), .B2(n9807), .ZN(n9805) );
  OAI21_X1 U10896 ( .B1(n9807), .B2(n9806), .A(n9805), .ZN(P1_U3291) );
  AND2_X1 U10897 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9808), .ZN(P1_U3292) );
  AND2_X1 U10898 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9808), .ZN(P1_U3293) );
  AND2_X1 U10899 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9808), .ZN(P1_U3294) );
  AND2_X1 U10900 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9808), .ZN(P1_U3295) );
  AND2_X1 U10901 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9808), .ZN(P1_U3296) );
  AND2_X1 U10902 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9808), .ZN(P1_U3297) );
  AND2_X1 U10903 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9808), .ZN(P1_U3298) );
  AND2_X1 U10904 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9808), .ZN(P1_U3299) );
  AND2_X1 U10905 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9808), .ZN(P1_U3300) );
  AND2_X1 U10906 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9808), .ZN(P1_U3301) );
  AND2_X1 U10907 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9808), .ZN(P1_U3302) );
  AND2_X1 U10908 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9808), .ZN(P1_U3303) );
  AND2_X1 U10909 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9808), .ZN(P1_U3304) );
  AND2_X1 U10910 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9808), .ZN(P1_U3305) );
  AND2_X1 U10911 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9808), .ZN(P1_U3306) );
  AND2_X1 U10912 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9808), .ZN(P1_U3307) );
  AND2_X1 U10913 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9808), .ZN(P1_U3308) );
  AND2_X1 U10914 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9808), .ZN(P1_U3309) );
  AND2_X1 U10915 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9808), .ZN(P1_U3310) );
  AND2_X1 U10916 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9808), .ZN(P1_U3311) );
  AND2_X1 U10917 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9808), .ZN(P1_U3312) );
  AND2_X1 U10918 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9808), .ZN(P1_U3313) );
  AND2_X1 U10919 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9808), .ZN(P1_U3314) );
  AND2_X1 U10920 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9808), .ZN(P1_U3315) );
  AND2_X1 U10921 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9808), .ZN(P1_U3316) );
  AND2_X1 U10922 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9808), .ZN(P1_U3317) );
  AND2_X1 U10923 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9808), .ZN(P1_U3318) );
  AND2_X1 U10924 ( .A1(n9808), .A2(P1_D_REG_4__SCAN_IN), .ZN(P1_U3319) );
  AND2_X1 U10925 ( .A1(n9808), .A2(P1_D_REG_3__SCAN_IN), .ZN(P1_U3320) );
  AND2_X1 U10926 ( .A1(n9808), .A2(P1_D_REG_2__SCAN_IN), .ZN(P1_U3321) );
  INV_X1 U10927 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10421) );
  OAI21_X1 U10928 ( .B1(n9810), .B2(n10421), .A(n9809), .ZN(P1_U3441) );
  AOI22_X1 U10929 ( .A1(n9888), .A2(n9889), .B1(n5866), .B2(n9887), .ZN(
        P1_U3454) );
  INV_X1 U10930 ( .A(n9811), .ZN(n9816) );
  OAI21_X1 U10931 ( .B1(n9813), .B2(n9869), .A(n9812), .ZN(n9815) );
  AOI211_X1 U10932 ( .C1(n9875), .C2(n9816), .A(n9815), .B(n9814), .ZN(n9891)
         );
  AOI22_X1 U10933 ( .A1(n9888), .A2(n9891), .B1(n5914), .B2(n9887), .ZN(
        P1_U3457) );
  INV_X1 U10934 ( .A(n9817), .ZN(n9822) );
  OAI21_X1 U10935 ( .B1(n9819), .B2(n9869), .A(n9818), .ZN(n9821) );
  AOI211_X1 U10936 ( .C1(n9875), .C2(n9822), .A(n9821), .B(n9820), .ZN(n9893)
         );
  INV_X1 U10937 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9823) );
  AOI22_X1 U10938 ( .A1(n9888), .A2(n9893), .B1(n9823), .B2(n9887), .ZN(
        P1_U3460) );
  OAI21_X1 U10939 ( .B1(n9825), .B2(n9869), .A(n9824), .ZN(n9827) );
  AOI211_X1 U10940 ( .C1(n9875), .C2(n9828), .A(n9827), .B(n9826), .ZN(n9894)
         );
  INV_X1 U10941 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9829) );
  AOI22_X1 U10942 ( .A1(n9888), .A2(n9894), .B1(n9829), .B2(n9887), .ZN(
        P1_U3463) );
  OAI21_X1 U10943 ( .B1(n9831), .B2(n9869), .A(n9830), .ZN(n9834) );
  INV_X1 U10944 ( .A(n9832), .ZN(n9833) );
  AOI211_X1 U10945 ( .C1(n9875), .C2(n9835), .A(n9834), .B(n9833), .ZN(n9895)
         );
  INV_X1 U10946 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9836) );
  AOI22_X1 U10947 ( .A1(n9888), .A2(n9895), .B1(n9836), .B2(n9887), .ZN(
        P1_U3466) );
  OAI211_X1 U10948 ( .C1(n9839), .C2(n9869), .A(n9838), .B(n9837), .ZN(n9841)
         );
  AOI211_X1 U10949 ( .C1(n9842), .C2(n9867), .A(n9841), .B(n9840), .ZN(n9896)
         );
  AOI22_X1 U10950 ( .A1(n9888), .A2(n9896), .B1(n5994), .B2(n9887), .ZN(
        P1_U3469) );
  AOI22_X1 U10951 ( .A1(n9856), .A2(n9844), .B1(n9843), .B2(n9857), .ZN(n9845)
         );
  OAI211_X1 U10952 ( .C1(n9847), .C2(n9869), .A(n9846), .B(n9845), .ZN(n9852)
         );
  INV_X1 U10953 ( .A(n9853), .ZN(n9850) );
  OAI21_X1 U10954 ( .B1(n9850), .B2(n9849), .A(n9848), .ZN(n9851) );
  AOI211_X1 U10955 ( .C1(n9875), .C2(n9853), .A(n9852), .B(n9851), .ZN(n9897)
         );
  INV_X1 U10956 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9854) );
  AOI22_X1 U10957 ( .A1(n9888), .A2(n9897), .B1(n9854), .B2(n9887), .ZN(
        P1_U3472) );
  AOI22_X1 U10958 ( .A1(n9858), .A2(n9857), .B1(n9856), .B2(n9855), .ZN(n9859)
         );
  OAI211_X1 U10959 ( .C1(n9861), .C2(n9869), .A(n9860), .B(n9859), .ZN(n9865)
         );
  NOR2_X1 U10960 ( .A1(n9863), .A2(n9862), .ZN(n9864) );
  AOI211_X1 U10961 ( .C1(n9867), .C2(n9866), .A(n9865), .B(n9864), .ZN(n9898)
         );
  AOI22_X1 U10962 ( .A1(n9888), .A2(n9898), .B1(n6037), .B2(n9887), .ZN(
        P1_U3475) );
  OAI21_X1 U10963 ( .B1(n9870), .B2(n9869), .A(n9868), .ZN(n9873) );
  INV_X1 U10964 ( .A(n9871), .ZN(n9872) );
  AOI211_X1 U10965 ( .C1(n9875), .C2(n9874), .A(n9873), .B(n9872), .ZN(n9899)
         );
  INV_X1 U10966 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9876) );
  AOI22_X1 U10967 ( .A1(n9888), .A2(n9899), .B1(n9876), .B2(n9887), .ZN(
        P1_U3478) );
  INV_X1 U10968 ( .A(n9882), .ZN(n9885) );
  AOI211_X1 U10969 ( .C1(n9880), .C2(n9879), .A(n9878), .B(n9877), .ZN(n9881)
         );
  OAI21_X1 U10970 ( .B1(n9883), .B2(n9882), .A(n9881), .ZN(n9884) );
  AOI21_X1 U10971 ( .B1(n9886), .B2(n9885), .A(n9884), .ZN(n9901) );
  AOI22_X1 U10972 ( .A1(n9888), .A2(n9901), .B1(n6086), .B2(n9887), .ZN(
        P1_U3481) );
  AOI22_X1 U10973 ( .A1(n9902), .A2(n9889), .B1(n5895), .B2(n9900), .ZN(
        P1_U3523) );
  AOI22_X1 U10974 ( .A1(n9902), .A2(n9891), .B1(n9890), .B2(n9900), .ZN(
        P1_U3524) );
  AOI22_X1 U10975 ( .A1(n9902), .A2(n9893), .B1(n9892), .B2(n9900), .ZN(
        P1_U3525) );
  AOI22_X1 U10976 ( .A1(n9902), .A2(n9894), .B1(n5953), .B2(n9900), .ZN(
        P1_U3526) );
  AOI22_X1 U10977 ( .A1(n9902), .A2(n9895), .B1(n5969), .B2(n9900), .ZN(
        P1_U3527) );
  AOI22_X1 U10978 ( .A1(n9902), .A2(n9896), .B1(n5995), .B2(n9900), .ZN(
        P1_U3528) );
  AOI22_X1 U10979 ( .A1(n9902), .A2(n9897), .B1(n6013), .B2(n9900), .ZN(
        P1_U3529) );
  AOI22_X1 U10980 ( .A1(n9902), .A2(n9898), .B1(n6041), .B2(n9900), .ZN(
        P1_U3530) );
  AOI22_X1 U10981 ( .A1(n9902), .A2(n9899), .B1(n6062), .B2(n9900), .ZN(
        P1_U3531) );
  AOI22_X1 U10982 ( .A1(n9902), .A2(n9901), .B1(n6090), .B2(n9900), .ZN(
        P1_U3532) );
  AOI22_X1 U10983 ( .A1(n9903), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9904), .ZN(n9913) );
  NAND2_X1 U10984 ( .A1(n9904), .A2(n10044), .ZN(n9905) );
  OAI211_X1 U10985 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n9907), .A(n9906), .B(
        n9905), .ZN(n9908) );
  INV_X1 U10986 ( .A(n9908), .ZN(n9911) );
  AOI22_X1 U10987 ( .A1(n9909), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9910) );
  OAI221_X1 U10988 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9913), .C1(n9912), .C2(
        n9911), .A(n9910), .ZN(P2_U3245) );
  XOR2_X1 U10989 ( .A(n9920), .B(n9914), .Z(n9919) );
  AOI222_X1 U10990 ( .A1(n9938), .A2(n9919), .B1(n9918), .B2(n9917), .C1(n9916), .C2(n9915), .ZN(n9983) );
  XNOR2_X1 U10991 ( .A(n9921), .B(n9920), .ZN(n9986) );
  NAND2_X1 U10992 ( .A1(n9986), .A2(n9944), .ZN(n9931) );
  XNOR2_X1 U10993 ( .A(n9923), .B(n9922), .ZN(n9982) );
  OAI22_X1 U10994 ( .A1(n9948), .A2(n9982), .B1(n9925), .B2(n9924), .ZN(n9929)
         );
  INV_X1 U10995 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9926) );
  NOR2_X1 U10996 ( .A1(n9927), .A2(n9926), .ZN(n9928) );
  NOR2_X1 U10997 ( .A1(n9929), .A2(n9928), .ZN(n9930) );
  OAI211_X1 U10998 ( .C1(n9981), .C2(n9951), .A(n9931), .B(n9930), .ZN(n9932)
         );
  INV_X1 U10999 ( .A(n9932), .ZN(n9933) );
  OAI21_X1 U11000 ( .B1(n9941), .B2(n9983), .A(n9933), .ZN(P2_U3292) );
  OAI21_X1 U11001 ( .B1(n9936), .B2(n9935), .A(n9934), .ZN(n9939) );
  AOI21_X1 U11002 ( .B1(n9939), .B2(n9938), .A(n9937), .ZN(n9969) );
  AOI22_X1 U11003 ( .A1(P2_REG2_REG_2__SCAN_IN), .A2(n9941), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n9940), .ZN(n9954) );
  XNOR2_X1 U11004 ( .A(n9943), .B(n9942), .ZN(n9972) );
  NAND2_X1 U11005 ( .A1(n9944), .A2(n9972), .ZN(n9950) );
  OR2_X1 U11006 ( .A1(n9945), .A2(n9967), .ZN(n9946) );
  NAND2_X1 U11007 ( .A1(n9947), .A2(n9946), .ZN(n9968) );
  OR2_X1 U11008 ( .A1(n9948), .A2(n9968), .ZN(n9949) );
  OAI211_X1 U11009 ( .C1(n9967), .C2(n9951), .A(n9950), .B(n9949), .ZN(n9952)
         );
  INV_X1 U11010 ( .A(n9952), .ZN(n9953) );
  OAI211_X1 U11011 ( .C1(n9941), .C2(n9969), .A(n9954), .B(n9953), .ZN(
        P2_U3294) );
  AND2_X1 U11012 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9959), .ZN(P2_U3297) );
  AND2_X1 U11013 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9959), .ZN(P2_U3298) );
  AND2_X1 U11014 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9959), .ZN(P2_U3299) );
  AND2_X1 U11015 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9959), .ZN(P2_U3300) );
  AND2_X1 U11016 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9959), .ZN(P2_U3301) );
  AND2_X1 U11017 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9959), .ZN(P2_U3302) );
  AND2_X1 U11018 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9959), .ZN(P2_U3303) );
  AND2_X1 U11019 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9959), .ZN(P2_U3304) );
  AND2_X1 U11020 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9959), .ZN(P2_U3305) );
  AND2_X1 U11021 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9959), .ZN(P2_U3306) );
  AND2_X1 U11022 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9959), .ZN(P2_U3307) );
  AND2_X1 U11023 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9959), .ZN(P2_U3308) );
  AND2_X1 U11024 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9959), .ZN(P2_U3309) );
  AND2_X1 U11025 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9959), .ZN(P2_U3310) );
  AND2_X1 U11026 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9959), .ZN(P2_U3311) );
  AND2_X1 U11027 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9959), .ZN(P2_U3312) );
  AND2_X1 U11028 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9959), .ZN(P2_U3313) );
  AND2_X1 U11029 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9959), .ZN(P2_U3314) );
  AND2_X1 U11030 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9959), .ZN(P2_U3315) );
  AND2_X1 U11031 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9959), .ZN(P2_U3316) );
  AND2_X1 U11032 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9959), .ZN(P2_U3317) );
  AND2_X1 U11033 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9959), .ZN(P2_U3318) );
  AND2_X1 U11034 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9959), .ZN(P2_U3319) );
  AND2_X1 U11035 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9959), .ZN(P2_U3320) );
  AND2_X1 U11036 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9959), .ZN(P2_U3321) );
  AND2_X1 U11037 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9959), .ZN(P2_U3322) );
  AND2_X1 U11038 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9959), .ZN(P2_U3323) );
  AND2_X1 U11039 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9959), .ZN(P2_U3324) );
  AND2_X1 U11040 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9959), .ZN(P2_U3325) );
  AND2_X1 U11041 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9959), .ZN(P2_U3326) );
  AOI22_X1 U11042 ( .A1(n9962), .A2(n9958), .B1(n9957), .B2(n9959), .ZN(
        P2_U3437) );
  AOI22_X1 U11043 ( .A1(n9962), .A2(n9961), .B1(n9960), .B2(n9959), .ZN(
        P2_U3438) );
  AOI22_X1 U11044 ( .A1(n9964), .A2(n10041), .B1(n4940), .B2(n9963), .ZN(n9965) );
  AND2_X1 U11045 ( .A1(n9966), .A2(n9965), .ZN(n10045) );
  AOI22_X1 U11046 ( .A1(n10043), .A2(n10045), .B1(n5141), .B2(n10042), .ZN(
        P2_U3451) );
  OAI22_X1 U11047 ( .A1(n9968), .A2(n10036), .B1(n9967), .B2(n10034), .ZN(
        n9971) );
  INV_X1 U11048 ( .A(n9969), .ZN(n9970) );
  AOI211_X1 U11049 ( .C1(n10041), .C2(n9972), .A(n9971), .B(n9970), .ZN(n10047) );
  AOI22_X1 U11050 ( .A1(n10043), .A2(n10047), .B1(n5152), .B2(n10042), .ZN(
        P2_U3457) );
  OAI22_X1 U11051 ( .A1(n9973), .A2(n10036), .B1(n4879), .B2(n10034), .ZN(
        n9974) );
  NOR2_X1 U11052 ( .A1(n9975), .A2(n9974), .ZN(n9980) );
  INV_X1 U11053 ( .A(n9976), .ZN(n9977) );
  OAI21_X1 U11054 ( .B1(n10020), .B2(n9978), .A(n9977), .ZN(n9979) );
  AND2_X1 U11055 ( .A1(n9980), .A2(n9979), .ZN(n10049) );
  AOI22_X1 U11056 ( .A1(n10043), .A2(n10049), .B1(n5173), .B2(n10042), .ZN(
        P2_U3460) );
  OAI22_X1 U11057 ( .A1(n9982), .A2(n10036), .B1(n9981), .B2(n10034), .ZN(
        n9985) );
  INV_X1 U11058 ( .A(n9983), .ZN(n9984) );
  AOI211_X1 U11059 ( .C1(n10041), .C2(n9986), .A(n9985), .B(n9984), .ZN(n10050) );
  AOI22_X1 U11060 ( .A1(n10043), .A2(n10050), .B1(n5200), .B2(n10042), .ZN(
        P2_U3463) );
  OAI211_X1 U11061 ( .C1(n9989), .C2(n10034), .A(n9988), .B(n9987), .ZN(n9990)
         );
  AOI21_X1 U11062 ( .B1(n10041), .B2(n9991), .A(n9990), .ZN(n10051) );
  AOI22_X1 U11063 ( .A1(n10043), .A2(n10051), .B1(n5231), .B2(n10042), .ZN(
        P2_U3466) );
  OAI22_X1 U11064 ( .A1(n9993), .A2(n10036), .B1(n9992), .B2(n10034), .ZN(
        n9994) );
  INV_X1 U11065 ( .A(n9994), .ZN(n9998) );
  OR2_X1 U11066 ( .A1(n9996), .A2(n9995), .ZN(n9997) );
  AND3_X1 U11067 ( .A1(n9999), .A2(n9998), .A3(n9997), .ZN(n10053) );
  AOI22_X1 U11068 ( .A1(n10043), .A2(n10053), .B1(n5255), .B2(n10042), .ZN(
        P2_U3469) );
  NAND2_X1 U11069 ( .A1(n10000), .A2(n10041), .ZN(n10006) );
  AOI22_X1 U11070 ( .A1(n10004), .A2(n10003), .B1(n10002), .B2(n10001), .ZN(
        n10005) );
  AND3_X1 U11071 ( .A1(n10007), .A2(n10006), .A3(n10005), .ZN(n10055) );
  AOI22_X1 U11072 ( .A1(n10043), .A2(n10055), .B1(n5276), .B2(n10042), .ZN(
        P2_U3472) );
  OAI22_X1 U11073 ( .A1(n10008), .A2(n10036), .B1(n4883), .B2(n10034), .ZN(
        n10011) );
  INV_X1 U11074 ( .A(n10009), .ZN(n10010) );
  AOI211_X1 U11075 ( .C1(n10020), .C2(n10012), .A(n10011), .B(n10010), .ZN(
        n10057) );
  AOI22_X1 U11076 ( .A1(n10043), .A2(n10057), .B1(n5306), .B2(n10042), .ZN(
        P2_U3475) );
  INV_X1 U11077 ( .A(n10013), .ZN(n10016) );
  INV_X1 U11078 ( .A(n10014), .ZN(n10015) );
  OAI22_X1 U11079 ( .A1(n10016), .A2(n10036), .B1(n10015), .B2(n10034), .ZN(
        n10018) );
  AOI211_X1 U11080 ( .C1(n10020), .C2(n10019), .A(n10018), .B(n10017), .ZN(
        n10059) );
  AOI22_X1 U11081 ( .A1(n10043), .A2(n10059), .B1(n5326), .B2(n10042), .ZN(
        P2_U3478) );
  NAND2_X1 U11082 ( .A1(n10021), .A2(n10041), .ZN(n10026) );
  OAI22_X1 U11083 ( .A1(n10023), .A2(n10036), .B1(n10022), .B2(n10034), .ZN(
        n10024) );
  INV_X1 U11084 ( .A(n10024), .ZN(n10025) );
  AND3_X1 U11085 ( .A1(n10027), .A2(n10026), .A3(n10025), .ZN(n10060) );
  AOI22_X1 U11086 ( .A1(n10043), .A2(n10060), .B1(n5358), .B2(n10042), .ZN(
        P2_U3481) );
  INV_X1 U11087 ( .A(n10028), .ZN(n10033) );
  OAI22_X1 U11088 ( .A1(n10030), .A2(n10036), .B1(n10029), .B2(n10034), .ZN(
        n10032) );
  AOI211_X1 U11089 ( .C1(n10033), .C2(n10041), .A(n10032), .B(n10031), .ZN(
        n10061) );
  AOI22_X1 U11090 ( .A1(n10043), .A2(n10061), .B1(n5378), .B2(n10042), .ZN(
        P2_U3484) );
  OAI22_X1 U11091 ( .A1(n10037), .A2(n10036), .B1(n10035), .B2(n10034), .ZN(
        n10039) );
  AOI211_X1 U11092 ( .C1(n10041), .C2(n10040), .A(n10039), .B(n10038), .ZN(
        n10063) );
  AOI22_X1 U11093 ( .A1(n10043), .A2(n10063), .B1(n5405), .B2(n10042), .ZN(
        P2_U3487) );
  AOI22_X1 U11094 ( .A1(n10064), .A2(n10045), .B1(n10044), .B2(n10062), .ZN(
        P2_U3520) );
  INV_X1 U11095 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10046) );
  AOI22_X1 U11096 ( .A1(n10064), .A2(n10047), .B1(n10046), .B2(n10062), .ZN(
        P2_U3522) );
  INV_X1 U11097 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10048) );
  AOI22_X1 U11098 ( .A1(n10064), .A2(n10049), .B1(n10048), .B2(n10062), .ZN(
        P2_U3523) );
  AOI22_X1 U11099 ( .A1(n10064), .A2(n10050), .B1(n6588), .B2(n10062), .ZN(
        P2_U3524) );
  AOI22_X1 U11100 ( .A1(n10064), .A2(n10051), .B1(n5226), .B2(n10062), .ZN(
        P2_U3525) );
  INV_X1 U11101 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10052) );
  AOI22_X1 U11102 ( .A1(n10064), .A2(n10053), .B1(n10052), .B2(n10062), .ZN(
        P2_U3526) );
  INV_X1 U11103 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10054) );
  AOI22_X1 U11104 ( .A1(n10064), .A2(n10055), .B1(n10054), .B2(n10062), .ZN(
        P2_U3527) );
  INV_X1 U11105 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10056) );
  AOI22_X1 U11106 ( .A1(n10064), .A2(n10057), .B1(n10056), .B2(n10062), .ZN(
        P2_U3528) );
  AOI22_X1 U11107 ( .A1(n10064), .A2(n10059), .B1(n10058), .B2(n10062), .ZN(
        P2_U3529) );
  AOI22_X1 U11108 ( .A1(n10064), .A2(n10060), .B1(n6953), .B2(n10062), .ZN(
        P2_U3530) );
  AOI22_X1 U11109 ( .A1(n10064), .A2(n10061), .B1(n7051), .B2(n10062), .ZN(
        P2_U3531) );
  AOI22_X1 U11110 ( .A1(n10064), .A2(n10063), .B1(n7289), .B2(n10062), .ZN(
        P2_U3532) );
  NAND3_X1 U11111 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10072) );
  AOI21_X1 U11112 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10074) );
  INV_X1 U11113 ( .A(n10074), .ZN(n10065) );
  NAND2_X1 U11114 ( .A1(n10072), .A2(n10065), .ZN(n10066) );
  XNOR2_X1 U11115 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10066), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11116 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  NOR2_X1 U11117 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10067) );
  AOI21_X1 U11118 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10067), .ZN(n10098) );
  NOR2_X1 U11119 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10068) );
  AOI21_X1 U11120 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10068), .ZN(n10101) );
  NOR2_X1 U11121 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10069) );
  AOI21_X1 U11122 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10069), .ZN(n10104) );
  NOR2_X1 U11123 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10070) );
  AOI21_X1 U11124 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10070), .ZN(n10107) );
  NOR2_X1 U11125 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10071) );
  AOI21_X1 U11126 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10071), .ZN(n10110) );
  NOR2_X1 U11127 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10080) );
  XNOR2_X1 U11128 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10515) );
  NAND2_X1 U11129 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10078) );
  XOR2_X1 U11130 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10513) );
  NAND2_X1 U11131 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n10076) );
  XOR2_X1 U11132 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10500) );
  INV_X1 U11133 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10073) );
  OAI21_X1 U11134 ( .B1(n10074), .B2(n10073), .A(n10072), .ZN(n10499) );
  NAND2_X1 U11135 ( .A1(n10500), .A2(n10499), .ZN(n10075) );
  NAND2_X1 U11136 ( .A1(n10076), .A2(n10075), .ZN(n10512) );
  NAND2_X1 U11137 ( .A1(n10513), .A2(n10512), .ZN(n10077) );
  NAND2_X1 U11138 ( .A1(n10078), .A2(n10077), .ZN(n10514) );
  NOR2_X1 U11139 ( .A1(n10515), .A2(n10514), .ZN(n10079) );
  NOR2_X1 U11140 ( .A1(n10080), .A2(n10079), .ZN(n10081) );
  NOR2_X1 U11141 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10081), .ZN(n10502) );
  AND2_X1 U11142 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10081), .ZN(n10501) );
  NOR2_X1 U11143 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10501), .ZN(n10082) );
  NOR2_X1 U11144 ( .A1(n10502), .A2(n10082), .ZN(n10083) );
  NAND2_X1 U11145 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n10083), .ZN(n10085) );
  XOR2_X1 U11146 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n10083), .Z(n10511) );
  NAND2_X1 U11147 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10511), .ZN(n10084) );
  NAND2_X1 U11148 ( .A1(n10085), .A2(n10084), .ZN(n10086) );
  NAND2_X1 U11149 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n10086), .ZN(n10088) );
  XOR2_X1 U11150 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n10086), .Z(n10498) );
  NAND2_X1 U11151 ( .A1(n10498), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n10087) );
  NAND2_X1 U11152 ( .A1(n10088), .A2(n10087), .ZN(n10089) );
  NAND2_X1 U11153 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n10089), .ZN(n10091) );
  XOR2_X1 U11154 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n10089), .Z(n10509) );
  NAND2_X1 U11155 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10509), .ZN(n10090) );
  NAND2_X1 U11156 ( .A1(n10091), .A2(n10090), .ZN(n10092) );
  AND2_X1 U11157 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10092), .ZN(n10093) );
  XNOR2_X1 U11158 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n10092), .ZN(n10496) );
  NOR2_X1 U11159 ( .A1(n10496), .A2(n10495), .ZN(n10494) );
  NAND2_X1 U11160 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n10094) );
  OAI21_X1 U11161 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10094), .ZN(n10118) );
  AOI21_X1 U11162 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10117), .ZN(n10116) );
  NAND2_X1 U11163 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n10095) );
  OAI21_X1 U11164 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10095), .ZN(n10115) );
  NOR2_X1 U11165 ( .A1(n10116), .A2(n10115), .ZN(n10114) );
  AOI21_X1 U11166 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10114), .ZN(n10113) );
  NOR2_X1 U11167 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10096) );
  AOI21_X1 U11168 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10096), .ZN(n10112) );
  NAND2_X1 U11169 ( .A1(n10113), .A2(n10112), .ZN(n10111) );
  OAI21_X1 U11170 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10111), .ZN(n10109) );
  NAND2_X1 U11171 ( .A1(n10110), .A2(n10109), .ZN(n10108) );
  OAI21_X1 U11172 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10108), .ZN(n10106) );
  NAND2_X1 U11173 ( .A1(n10107), .A2(n10106), .ZN(n10105) );
  OAI21_X1 U11174 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10105), .ZN(n10103) );
  NAND2_X1 U11175 ( .A1(n10104), .A2(n10103), .ZN(n10102) );
  OAI21_X1 U11176 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10102), .ZN(n10100) );
  NAND2_X1 U11177 ( .A1(n10101), .A2(n10100), .ZN(n10099) );
  OAI21_X1 U11178 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10099), .ZN(n10097) );
  NAND2_X1 U11179 ( .A1(n10098), .A2(n10097), .ZN(n10488) );
  OAI21_X1 U11180 ( .B1(n10098), .B2(n10097), .A(n10488), .ZN(ADD_1071_U56) );
  OAI21_X1 U11181 ( .B1(n10101), .B2(n10100), .A(n10099), .ZN(ADD_1071_U57) );
  OAI21_X1 U11182 ( .B1(n10104), .B2(n10103), .A(n10102), .ZN(ADD_1071_U58) );
  OAI21_X1 U11183 ( .B1(n10107), .B2(n10106), .A(n10105), .ZN(ADD_1071_U59) );
  OAI21_X1 U11184 ( .B1(n10110), .B2(n10109), .A(n10108), .ZN(ADD_1071_U60) );
  OAI21_X1 U11185 ( .B1(n10113), .B2(n10112), .A(n10111), .ZN(ADD_1071_U61) );
  AOI21_X1 U11186 ( .B1(n10116), .B2(n10115), .A(n10114), .ZN(ADD_1071_U62) );
  AOI21_X1 U11187 ( .B1(n10119), .B2(n10118), .A(n10117), .ZN(ADD_1071_U63) );
  XOR2_X1 U11188 ( .A(SI_8_), .B(keyinput_g24), .Z(n10126) );
  AOI22_X1 U11189 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(keyinput_g79), .B1(
        P1_IR_REG_27__SCAN_IN), .B2(keyinput_g118), .ZN(n10120) );
  OAI221_X1 U11190 ( .B1(P2_DATAO_REG_17__SCAN_IN), .B2(keyinput_g79), .C1(
        P1_IR_REG_27__SCAN_IN), .C2(keyinput_g118), .A(n10120), .ZN(n10125) );
  AOI22_X1 U11191 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(keyinput_g116), .B1(
        P1_IR_REG_21__SCAN_IN), .B2(keyinput_g112), .ZN(n10121) );
  OAI221_X1 U11192 ( .B1(P1_IR_REG_25__SCAN_IN), .B2(keyinput_g116), .C1(
        P1_IR_REG_21__SCAN_IN), .C2(keyinput_g112), .A(n10121), .ZN(n10124) );
  AOI22_X1 U11193 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput_g45), .B1(
        SI_25_), .B2(keyinput_g7), .ZN(n10122) );
  OAI221_X1 U11194 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_g45), .C1(
        SI_25_), .C2(keyinput_g7), .A(n10122), .ZN(n10123) );
  NOR4_X1 U11195 ( .A1(n10126), .A2(n10125), .A3(n10124), .A4(n10123), .ZN(
        n10154) );
  AOI22_X1 U11196 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput_g88), .B1(
        P1_IR_REG_22__SCAN_IN), .B2(keyinput_g113), .ZN(n10127) );
  OAI221_X1 U11197 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_g88), .C1(
        P1_IR_REG_22__SCAN_IN), .C2(keyinput_g113), .A(n10127), .ZN(n10134) );
  AOI22_X1 U11198 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_g60), .B1(
        P1_IR_REG_18__SCAN_IN), .B2(keyinput_g109), .ZN(n10128) );
  OAI221_X1 U11199 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .C1(
        P1_IR_REG_18__SCAN_IN), .C2(keyinput_g109), .A(n10128), .ZN(n10133) );
  AOI22_X1 U11200 ( .A1(SI_0_), .A2(keyinput_g32), .B1(P1_D_REG_4__SCAN_IN), 
        .B2(keyinput_g127), .ZN(n10129) );
  OAI221_X1 U11201 ( .B1(SI_0_), .B2(keyinput_g32), .C1(P1_D_REG_4__SCAN_IN), 
        .C2(keyinput_g127), .A(n10129), .ZN(n10132) );
  AOI22_X1 U11202 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(keyinput_g66), .B1(
        SI_26_), .B2(keyinput_g6), .ZN(n10130) );
  OAI221_X1 U11203 ( .B1(P2_DATAO_REG_30__SCAN_IN), .B2(keyinput_g66), .C1(
        SI_26_), .C2(keyinput_g6), .A(n10130), .ZN(n10131) );
  NOR4_X1 U11204 ( .A1(n10134), .A2(n10133), .A3(n10132), .A4(n10131), .ZN(
        n10153) );
  AOI22_X1 U11205 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_g44), .B1(
        P1_D_REG_3__SCAN_IN), .B2(keyinput_g126), .ZN(n10135) );
  OAI221_X1 U11206 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_g44), .C1(
        P1_D_REG_3__SCAN_IN), .C2(keyinput_g126), .A(n10135), .ZN(n10142) );
  AOI22_X1 U11207 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_g39), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .ZN(n10136) );
  OAI221_X1 U11208 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .C1(
        P2_REG3_REG_16__SCAN_IN), .C2(keyinput_g48), .A(n10136), .ZN(n10141)
         );
  AOI22_X1 U11209 ( .A1(SI_3_), .A2(keyinput_g29), .B1(P2_RD_REG_SCAN_IN), 
        .B2(keyinput_g33), .ZN(n10137) );
  OAI221_X1 U11210 ( .B1(SI_3_), .B2(keyinput_g29), .C1(P2_RD_REG_SCAN_IN), 
        .C2(keyinput_g33), .A(n10137), .ZN(n10140) );
  AOI22_X1 U11211 ( .A1(SI_29_), .A2(keyinput_g3), .B1(P1_IR_REG_11__SCAN_IN), 
        .B2(keyinput_g102), .ZN(n10138) );
  OAI221_X1 U11212 ( .B1(SI_29_), .B2(keyinput_g3), .C1(P1_IR_REG_11__SCAN_IN), 
        .C2(keyinput_g102), .A(n10138), .ZN(n10139) );
  NOR4_X1 U11213 ( .A1(n10142), .A2(n10141), .A3(n10140), .A4(n10139), .ZN(
        n10152) );
  AOI22_X1 U11214 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_g36), .B1(
        P1_IR_REG_4__SCAN_IN), .B2(keyinput_g95), .ZN(n10143) );
  OAI221_X1 U11215 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .C1(
        P1_IR_REG_4__SCAN_IN), .C2(keyinput_g95), .A(n10143), .ZN(n10150) );
  AOI22_X1 U11216 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_g37), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(keyinput_g90), .ZN(n10144) );
  OAI221_X1 U11217 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .C1(
        P2_DATAO_REG_6__SCAN_IN), .C2(keyinput_g90), .A(n10144), .ZN(n10149)
         );
  AOI22_X1 U11218 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(keyinput_g121), .B1(SI_17_), .B2(keyinput_g15), .ZN(n10145) );
  OAI221_X1 U11219 ( .B1(P1_IR_REG_30__SCAN_IN), .B2(keyinput_g121), .C1(
        SI_17_), .C2(keyinput_g15), .A(n10145), .ZN(n10148) );
  AOI22_X1 U11220 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_g62), .B1(
        P1_IR_REG_13__SCAN_IN), .B2(keyinput_g104), .ZN(n10146) );
  OAI221_X1 U11221 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .C1(
        P1_IR_REG_13__SCAN_IN), .C2(keyinput_g104), .A(n10146), .ZN(n10147) );
  NOR4_X1 U11222 ( .A1(n10150), .A2(n10149), .A3(n10148), .A4(n10147), .ZN(
        n10151) );
  NAND4_X1 U11223 ( .A1(n10154), .A2(n10153), .A3(n10152), .A4(n10151), .ZN(
        n10289) );
  AOI22_X1 U11224 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_g0), .B1(
        P1_D_REG_0__SCAN_IN), .B2(keyinput_g123), .ZN(n10155) );
  OAI221_X1 U11225 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_g0), .C1(
        P1_D_REG_0__SCAN_IN), .C2(keyinput_g123), .A(n10155), .ZN(n10162) );
  AOI22_X1 U11226 ( .A1(SI_28_), .A2(keyinput_g4), .B1(SI_15_), .B2(
        keyinput_g17), .ZN(n10156) );
  OAI221_X1 U11227 ( .B1(SI_28_), .B2(keyinput_g4), .C1(SI_15_), .C2(
        keyinput_g17), .A(n10156), .ZN(n10161) );
  AOI22_X1 U11228 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(keyinput_g77), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_g75), .ZN(n10157) );
  OAI221_X1 U11229 ( .B1(P2_DATAO_REG_19__SCAN_IN), .B2(keyinput_g77), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput_g75), .A(n10157), .ZN(n10160)
         );
  AOI22_X1 U11230 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(keyinput_g86), .B1(
        P1_IR_REG_3__SCAN_IN), .B2(keyinput_g94), .ZN(n10158) );
  OAI221_X1 U11231 ( .B1(P2_DATAO_REG_10__SCAN_IN), .B2(keyinput_g86), .C1(
        P1_IR_REG_3__SCAN_IN), .C2(keyinput_g94), .A(n10158), .ZN(n10159) );
  NOR4_X1 U11232 ( .A1(n10162), .A2(n10161), .A3(n10160), .A4(n10159), .ZN(
        n10190) );
  AOI22_X1 U11233 ( .A1(SI_30_), .A2(keyinput_g2), .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .ZN(n10163) );
  OAI221_X1 U11234 ( .B1(SI_30_), .B2(keyinput_g2), .C1(
        P2_REG3_REG_13__SCAN_IN), .C2(keyinput_g56), .A(n10163), .ZN(n10170)
         );
  AOI22_X1 U11235 ( .A1(SI_2_), .A2(keyinput_g30), .B1(SI_27_), .B2(
        keyinput_g5), .ZN(n10164) );
  OAI221_X1 U11236 ( .B1(SI_2_), .B2(keyinput_g30), .C1(SI_27_), .C2(
        keyinput_g5), .A(n10164), .ZN(n10169) );
  AOI22_X1 U11237 ( .A1(SI_1_), .A2(keyinput_g31), .B1(SI_20_), .B2(
        keyinput_g12), .ZN(n10165) );
  OAI221_X1 U11238 ( .B1(SI_1_), .B2(keyinput_g31), .C1(SI_20_), .C2(
        keyinput_g12), .A(n10165), .ZN(n10168) );
  AOI22_X1 U11239 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_g54), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(keyinput_g81), .ZN(n10166) );
  OAI221_X1 U11240 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .C1(
        P2_DATAO_REG_15__SCAN_IN), .C2(keyinput_g81), .A(n10166), .ZN(n10167)
         );
  NOR4_X1 U11241 ( .A1(n10170), .A2(n10169), .A3(n10168), .A4(n10167), .ZN(
        n10189) );
  AOI22_X1 U11242 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(keyinput_g83), .B1(
        P1_D_REG_2__SCAN_IN), .B2(keyinput_g125), .ZN(n10171) );
  OAI221_X1 U11243 ( .B1(P2_DATAO_REG_13__SCAN_IN), .B2(keyinput_g83), .C1(
        P1_D_REG_2__SCAN_IN), .C2(keyinput_g125), .A(n10171), .ZN(n10178) );
  AOI22_X1 U11244 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_g40), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput_g34), .ZN(n10172) );
  OAI221_X1 U11245 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_g40), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput_g34), .A(n10172), .ZN(n10177) );
  AOI22_X1 U11246 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(keyinput_g67), .B1(
        P1_IR_REG_31__SCAN_IN), .B2(keyinput_g122), .ZN(n10173) );
  OAI221_X1 U11247 ( .B1(P2_DATAO_REG_29__SCAN_IN), .B2(keyinput_g67), .C1(
        P1_IR_REG_31__SCAN_IN), .C2(keyinput_g122), .A(n10173), .ZN(n10176) );
  AOI22_X1 U11248 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(keyinput_g85), .B1(
        P1_IR_REG_23__SCAN_IN), .B2(keyinput_g114), .ZN(n10174) );
  OAI221_X1 U11249 ( .B1(P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_g85), .C1(
        P1_IR_REG_23__SCAN_IN), .C2(keyinput_g114), .A(n10174), .ZN(n10175) );
  NOR4_X1 U11250 ( .A1(n10178), .A2(n10177), .A3(n10176), .A4(n10175), .ZN(
        n10188) );
  AOI22_X1 U11251 ( .A1(SI_19_), .A2(keyinput_g13), .B1(SI_21_), .B2(
        keyinput_g11), .ZN(n10179) );
  OAI221_X1 U11252 ( .B1(SI_19_), .B2(keyinput_g13), .C1(SI_21_), .C2(
        keyinput_g11), .A(n10179), .ZN(n10186) );
  AOI22_X1 U11253 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_g55), .B1(
        P1_IR_REG_12__SCAN_IN), .B2(keyinput_g103), .ZN(n10180) );
  OAI221_X1 U11254 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .C1(
        P1_IR_REG_12__SCAN_IN), .C2(keyinput_g103), .A(n10180), .ZN(n10185) );
  AOI22_X1 U11255 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput_g63), .B1(
        SI_24_), .B2(keyinput_g8), .ZN(n10181) );
  OAI221_X1 U11256 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .C1(
        SI_24_), .C2(keyinput_g8), .A(n10181), .ZN(n10184) );
  AOI22_X1 U11257 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_g50), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(keyinput_g84), .ZN(n10182) );
  OAI221_X1 U11258 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .C1(
        P2_DATAO_REG_12__SCAN_IN), .C2(keyinput_g84), .A(n10182), .ZN(n10183)
         );
  NOR4_X1 U11259 ( .A1(n10186), .A2(n10185), .A3(n10184), .A4(n10183), .ZN(
        n10187) );
  NAND4_X1 U11260 ( .A1(n10190), .A2(n10189), .A3(n10188), .A4(n10187), .ZN(
        n10288) );
  AOI22_X1 U11261 ( .A1(n10192), .A2(keyinput_g87), .B1(n10423), .B2(
        keyinput_g10), .ZN(n10191) );
  OAI221_X1 U11262 ( .B1(n10192), .B2(keyinput_g87), .C1(n10423), .C2(
        keyinput_g10), .A(n10191), .ZN(n10202) );
  INV_X1 U11263 ( .A(SI_5_), .ZN(n10195) );
  AOI22_X1 U11264 ( .A1(n10195), .A2(keyinput_g27), .B1(n10194), .B2(
        keyinput_g80), .ZN(n10193) );
  OAI221_X1 U11265 ( .B1(n10195), .B2(keyinput_g27), .C1(n10194), .C2(
        keyinput_g80), .A(n10193), .ZN(n10201) );
  AOI22_X1 U11266 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(keyinput_g119), .B1(
        P1_IR_REG_17__SCAN_IN), .B2(keyinput_g108), .ZN(n10196) );
  OAI221_X1 U11267 ( .B1(P1_IR_REG_28__SCAN_IN), .B2(keyinput_g119), .C1(
        P1_IR_REG_17__SCAN_IN), .C2(keyinput_g108), .A(n10196), .ZN(n10200) );
  XNOR2_X1 U11268 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_g98), .ZN(n10198) );
  XNOR2_X1 U11269 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_g72), .ZN(n10197) );
  NAND2_X1 U11270 ( .A1(n10198), .A2(n10197), .ZN(n10199) );
  NOR4_X1 U11271 ( .A1(n10202), .A2(n10201), .A3(n10200), .A4(n10199), .ZN(
        n10234) );
  AOI22_X1 U11272 ( .A1(n10421), .A2(keyinput_g124), .B1(keyinput_g1), .B2(
        n10204), .ZN(n10203) );
  OAI221_X1 U11273 ( .B1(n10421), .B2(keyinput_g124), .C1(n10204), .C2(
        keyinput_g1), .A(n10203), .ZN(n10212) );
  AOI22_X1 U11274 ( .A1(n10424), .A2(keyinput_g57), .B1(n10395), .B2(
        keyinput_g23), .ZN(n10205) );
  OAI221_X1 U11275 ( .B1(n10424), .B2(keyinput_g57), .C1(n10395), .C2(
        keyinput_g23), .A(n10205), .ZN(n10211) );
  XOR2_X1 U11276 ( .A(n5368), .B(keyinput_g21), .Z(n10209) );
  XNOR2_X1 U11277 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_g96), .ZN(n10208) );
  XNOR2_X1 U11278 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_g105), .ZN(n10207)
         );
  XNOR2_X1 U11279 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_g106), .ZN(n10206)
         );
  NAND4_X1 U11280 ( .A1(n10209), .A2(n10208), .A3(n10207), .A4(n10206), .ZN(
        n10210) );
  NOR3_X1 U11281 ( .A1(n10212), .A2(n10211), .A3(n10210), .ZN(n10233) );
  AOI22_X1 U11282 ( .A1(n4717), .A2(keyinput_g111), .B1(keyinput_g20), .B2(
        n10363), .ZN(n10213) );
  OAI221_X1 U11283 ( .B1(n4717), .B2(keyinput_g111), .C1(n10363), .C2(
        keyinput_g20), .A(n10213), .ZN(n10220) );
  INV_X1 U11284 ( .A(SI_18_), .ZN(n10466) );
  AOI22_X1 U11285 ( .A1(n5880), .A2(keyinput_g115), .B1(keyinput_g14), .B2(
        n10466), .ZN(n10214) );
  OAI221_X1 U11286 ( .B1(n5880), .B2(keyinput_g115), .C1(n10466), .C2(
        keyinput_g14), .A(n10214), .ZN(n10219) );
  AOI22_X1 U11287 ( .A1(n10451), .A2(keyinput_g76), .B1(keyinput_g41), .B2(
        n5573), .ZN(n10215) );
  OAI221_X1 U11288 ( .B1(n10451), .B2(keyinput_g76), .C1(n5573), .C2(
        keyinput_g41), .A(n10215), .ZN(n10218) );
  AOI22_X1 U11289 ( .A1(n5841), .A2(keyinput_g97), .B1(keyinput_g68), .B2(
        n10426), .ZN(n10216) );
  OAI221_X1 U11290 ( .B1(n5841), .B2(keyinput_g97), .C1(n10426), .C2(
        keyinput_g68), .A(n10216), .ZN(n10217) );
  NOR4_X1 U11291 ( .A1(n10220), .A2(n10219), .A3(n10218), .A4(n10217), .ZN(
        n10232) );
  AOI22_X1 U11292 ( .A1(n5278), .A2(keyinput_g35), .B1(n10455), .B2(
        keyinput_g16), .ZN(n10221) );
  OAI221_X1 U11293 ( .B1(n5278), .B2(keyinput_g35), .C1(n10455), .C2(
        keyinput_g16), .A(n10221), .ZN(n10230) );
  AOI22_X1 U11294 ( .A1(n5700), .A2(keyinput_g47), .B1(n10223), .B2(
        keyinput_g18), .ZN(n10222) );
  OAI221_X1 U11295 ( .B1(n5700), .B2(keyinput_g47), .C1(n10223), .C2(
        keyinput_g18), .A(n10222), .ZN(n10229) );
  INV_X1 U11296 ( .A(SI_6_), .ZN(n10362) );
  AOI22_X1 U11297 ( .A1(n10437), .A2(keyinput_g71), .B1(keyinput_g26), .B2(
        n10362), .ZN(n10224) );
  OAI221_X1 U11298 ( .B1(n10437), .B2(keyinput_g71), .C1(n10362), .C2(
        keyinput_g26), .A(n10224), .ZN(n10228) );
  INV_X1 U11299 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n10452) );
  XOR2_X1 U11300 ( .A(n10452), .B(keyinput_g99), .Z(n10226) );
  XNOR2_X1 U11301 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_g92), .ZN(n10225) );
  NAND2_X1 U11302 ( .A1(n10226), .A2(n10225), .ZN(n10227) );
  NOR4_X1 U11303 ( .A1(n10230), .A2(n10229), .A3(n10228), .A4(n10227), .ZN(
        n10231) );
  NAND4_X1 U11304 ( .A1(n10234), .A2(n10233), .A3(n10232), .A4(n10231), .ZN(
        n10287) );
  INV_X1 U11305 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10236) );
  AOI22_X1 U11306 ( .A1(n10236), .A2(keyinput_g52), .B1(n5328), .B2(
        keyinput_g53), .ZN(n10235) );
  OAI221_X1 U11307 ( .B1(n10236), .B2(keyinput_g52), .C1(n5328), .C2(
        keyinput_g53), .A(n10235), .ZN(n10247) );
  AOI22_X1 U11308 ( .A1(n6238), .A2(keyinput_g107), .B1(keyinput_g78), .B2(
        n10238), .ZN(n10237) );
  OAI221_X1 U11309 ( .B1(n6238), .B2(keyinput_g107), .C1(n10238), .C2(
        keyinput_g78), .A(n10237), .ZN(n10246) );
  INV_X1 U11310 ( .A(SI_4_), .ZN(n10241) );
  INV_X1 U11311 ( .A(SI_7_), .ZN(n10240) );
  AOI22_X1 U11312 ( .A1(n10241), .A2(keyinput_g28), .B1(n10240), .B2(
        keyinput_g25), .ZN(n10239) );
  OAI221_X1 U11313 ( .B1(n10241), .B2(keyinput_g28), .C1(n10240), .C2(
        keyinput_g25), .A(n10239), .ZN(n10245) );
  XNOR2_X1 U11314 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_g91), .ZN(n10243) );
  XNOR2_X1 U11315 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_g38), .ZN(n10242)
         );
  NAND2_X1 U11316 ( .A1(n10243), .A2(n10242), .ZN(n10244) );
  NOR4_X1 U11317 ( .A1(n10247), .A2(n10246), .A3(n10245), .A4(n10244), .ZN(
        n10285) );
  AOI22_X1 U11318 ( .A1(n10390), .A2(keyinput_g9), .B1(keyinput_g120), .B2(
        n5858), .ZN(n10248) );
  OAI221_X1 U11319 ( .B1(n10390), .B2(keyinput_g9), .C1(n5858), .C2(
        keyinput_g120), .A(n10248), .ZN(n10259) );
  AOI22_X1 U11320 ( .A1(n5375), .A2(keyinput_g58), .B1(keyinput_g43), .B2(
        n10250), .ZN(n10249) );
  OAI221_X1 U11321 ( .B1(n5375), .B2(keyinput_g58), .C1(n10250), .C2(
        keyinput_g43), .A(n10249), .ZN(n10258) );
  AOI22_X1 U11322 ( .A1(n10253), .A2(keyinput_g51), .B1(n10252), .B2(
        keyinput_g82), .ZN(n10251) );
  OAI221_X1 U11323 ( .B1(n10253), .B2(keyinput_g51), .C1(n10252), .C2(
        keyinput_g82), .A(n10251), .ZN(n10257) );
  XNOR2_X1 U11324 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_g110), .ZN(n10255)
         );
  XNOR2_X1 U11325 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_g74), .ZN(n10254) );
  NAND2_X1 U11326 ( .A1(n10255), .A2(n10254), .ZN(n10256) );
  NOR4_X1 U11327 ( .A1(n10259), .A2(n10258), .A3(n10257), .A4(n10256), .ZN(
        n10284) );
  AOI22_X1 U11328 ( .A1(n10262), .A2(keyinput_g64), .B1(keyinput_g65), .B2(
        n10261), .ZN(n10260) );
  OAI221_X1 U11329 ( .B1(n10262), .B2(keyinput_g64), .C1(n10261), .C2(
        keyinput_g65), .A(n10260), .ZN(n10270) );
  AOI22_X1 U11330 ( .A1(n10380), .A2(keyinput_g89), .B1(keyinput_g59), .B2(
        n10365), .ZN(n10263) );
  OAI221_X1 U11331 ( .B1(n10380), .B2(keyinput_g89), .C1(n10365), .C2(
        keyinput_g59), .A(n10263), .ZN(n10269) );
  XOR2_X1 U11332 ( .A(n5834), .B(keyinput_g42), .Z(n10267) );
  XOR2_X1 U11333 ( .A(n5228), .B(keyinput_g49), .Z(n10266) );
  XNOR2_X1 U11334 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_g101), .ZN(n10265)
         );
  XNOR2_X1 U11335 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_g93), .ZN(n10264) );
  NAND4_X1 U11336 ( .A1(n10267), .A2(n10266), .A3(n10265), .A4(n10264), .ZN(
        n10268) );
  NOR3_X1 U11337 ( .A1(n10270), .A2(n10269), .A3(n10268), .ZN(n10283) );
  AOI22_X1 U11338 ( .A1(n10272), .A2(keyinput_g69), .B1(keyinput_g46), .B2(
        n10394), .ZN(n10271) );
  OAI221_X1 U11339 ( .B1(n10272), .B2(keyinput_g69), .C1(n10394), .C2(
        keyinput_g46), .A(n10271), .ZN(n10281) );
  AOI22_X1 U11340 ( .A1(n10449), .A2(keyinput_g70), .B1(keyinput_g73), .B2(
        n10465), .ZN(n10273) );
  OAI221_X1 U11341 ( .B1(n10449), .B2(keyinput_g70), .C1(n10465), .C2(
        keyinput_g73), .A(n10273), .ZN(n10280) );
  AOI22_X1 U11342 ( .A1(n10379), .A2(keyinput_g19), .B1(keyinput_g61), .B2(
        n10275), .ZN(n10274) );
  OAI221_X1 U11343 ( .B1(n10379), .B2(keyinput_g19), .C1(n10275), .C2(
        keyinput_g61), .A(n10274), .ZN(n10279) );
  INV_X1 U11344 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n10406) );
  XOR2_X1 U11345 ( .A(n10406), .B(keyinput_g100), .Z(n10277) );
  XNOR2_X1 U11346 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_g117), .ZN(n10276)
         );
  NAND2_X1 U11347 ( .A1(n10277), .A2(n10276), .ZN(n10278) );
  NOR4_X1 U11348 ( .A1(n10281), .A2(n10280), .A3(n10279), .A4(n10278), .ZN(
        n10282) );
  NAND4_X1 U11349 ( .A1(n10285), .A2(n10284), .A3(n10283), .A4(n10282), .ZN(
        n10286) );
  NOR4_X1 U11350 ( .A1(n10289), .A2(n10288), .A3(n10287), .A4(n10286), .ZN(
        n10487) );
  OAI22_X1 U11351 ( .A1(SI_14_), .A2(keyinput_f18), .B1(
        P2_REG3_REG_21__SCAN_IN), .B2(keyinput_f45), .ZN(n10290) );
  AOI221_X1 U11352 ( .B1(SI_14_), .B2(keyinput_f18), .C1(keyinput_f45), .C2(
        P2_REG3_REG_21__SCAN_IN), .A(n10290), .ZN(n10297) );
  OAI22_X1 U11353 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(keyinput_f80), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(keyinput_f84), .ZN(n10291) );
  AOI221_X1 U11354 ( .B1(P2_DATAO_REG_16__SCAN_IN), .B2(keyinput_f80), .C1(
        keyinput_f84), .C2(P2_DATAO_REG_12__SCAN_IN), .A(n10291), .ZN(n10296)
         );
  OAI22_X1 U11355 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput_f104), .B1(SI_26_), .B2(keyinput_f6), .ZN(n10292) );
  AOI221_X1 U11356 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput_f104), .C1(
        keyinput_f6), .C2(SI_26_), .A(n10292), .ZN(n10295) );
  OAI22_X1 U11357 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(keyinput_f108), .B1(SI_11_), .B2(keyinput_f21), .ZN(n10293) );
  AOI221_X1 U11358 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(keyinput_f108), .C1(
        keyinput_f21), .C2(SI_11_), .A(n10293), .ZN(n10294) );
  NAND4_X1 U11359 ( .A1(n10297), .A2(n10296), .A3(n10295), .A4(n10294), .ZN(
        n10326) );
  OAI22_X1 U11360 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_f47), .B1(
        P2_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .ZN(n10298) );
  AOI221_X1 U11361 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .C1(
        keyinput_f39), .C2(P2_REG3_REG_10__SCAN_IN), .A(n10298), .ZN(n10305)
         );
  OAI22_X1 U11362 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(keyinput_f109), .B1(
        P1_IR_REG_10__SCAN_IN), .B2(keyinput_f101), .ZN(n10299) );
  AOI221_X1 U11363 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(keyinput_f109), .C1(
        keyinput_f101), .C2(P1_IR_REG_10__SCAN_IN), .A(n10299), .ZN(n10304) );
  OAI22_X1 U11364 ( .A1(SI_30_), .A2(keyinput_f2), .B1(P2_WR_REG_SCAN_IN), 
        .B2(keyinput_f0), .ZN(n10300) );
  AOI221_X1 U11365 ( .B1(SI_30_), .B2(keyinput_f2), .C1(keyinput_f0), .C2(
        P2_WR_REG_SCAN_IN), .A(n10300), .ZN(n10303) );
  OAI22_X1 U11366 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(keyinput_f94), .B1(
        keyinput_f119), .B2(P1_IR_REG_28__SCAN_IN), .ZN(n10301) );
  AOI221_X1 U11367 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(keyinput_f94), .C1(
        P1_IR_REG_28__SCAN_IN), .C2(keyinput_f119), .A(n10301), .ZN(n10302) );
  NAND4_X1 U11368 ( .A1(n10305), .A2(n10304), .A3(n10303), .A4(n10302), .ZN(
        n10325) );
  OAI22_X1 U11369 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(keyinput_f115), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(keyinput_f78), .ZN(n10306) );
  AOI221_X1 U11370 ( .B1(P1_IR_REG_24__SCAN_IN), .B2(keyinput_f115), .C1(
        keyinput_f78), .C2(P2_DATAO_REG_18__SCAN_IN), .A(n10306), .ZN(n10313)
         );
  OAI22_X1 U11371 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(keyinput_f118), .B1(
        P2_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .ZN(n10307) );
  AOI221_X1 U11372 ( .B1(P1_IR_REG_27__SCAN_IN), .B2(keyinput_f118), .C1(
        keyinput_f51), .C2(P2_REG3_REG_24__SCAN_IN), .A(n10307), .ZN(n10312)
         );
  OAI22_X1 U11373 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(keyinput_f122), .B1(SI_8_), 
        .B2(keyinput_f24), .ZN(n10308) );
  AOI221_X1 U11374 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(keyinput_f122), .C1(
        keyinput_f24), .C2(SI_8_), .A(n10308), .ZN(n10311) );
  OAI22_X1 U11375 ( .A1(SI_19_), .A2(keyinput_f13), .B1(keyinput_f54), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n10309) );
  AOI221_X1 U11376 ( .B1(SI_19_), .B2(keyinput_f13), .C1(
        P2_REG3_REG_0__SCAN_IN), .C2(keyinput_f54), .A(n10309), .ZN(n10310) );
  NAND4_X1 U11377 ( .A1(n10313), .A2(n10312), .A3(n10311), .A4(n10310), .ZN(
        n10324) );
  OAI22_X1 U11378 ( .A1(SI_4_), .A2(keyinput_f28), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(keyinput_f40), .ZN(n10314) );
  AOI221_X1 U11379 ( .B1(SI_4_), .B2(keyinput_f28), .C1(keyinput_f40), .C2(
        P2_REG3_REG_3__SCAN_IN), .A(n10314), .ZN(n10322) );
  OAI22_X1 U11380 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(keyinput_f93), .B1(
        P2_B_REG_SCAN_IN), .B2(keyinput_f64), .ZN(n10315) );
  AOI221_X1 U11381 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(keyinput_f93), .C1(
        keyinput_f64), .C2(P2_B_REG_SCAN_IN), .A(n10315), .ZN(n10321) );
  OAI22_X1 U11382 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput_f88), .B1(
        keyinput_f25), .B2(SI_7_), .ZN(n10316) );
  AOI221_X1 U11383 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_f88), .C1(
        SI_7_), .C2(keyinput_f25), .A(n10316), .ZN(n10320) );
  OAI22_X1 U11384 ( .A1(n10318), .A2(keyinput_f55), .B1(keyinput_f1), .B2(
        SI_31_), .ZN(n10317) );
  AOI221_X1 U11385 ( .B1(n10318), .B2(keyinput_f55), .C1(SI_31_), .C2(
        keyinput_f1), .A(n10317), .ZN(n10319) );
  NAND4_X1 U11386 ( .A1(n10322), .A2(n10321), .A3(n10320), .A4(n10319), .ZN(
        n10323) );
  NOR4_X1 U11387 ( .A1(n10326), .A2(n10325), .A3(n10324), .A4(n10323), .ZN(
        n10483) );
  OAI22_X1 U11388 ( .A1(SI_1_), .A2(keyinput_f31), .B1(keyinput_f52), .B2(
        P2_REG3_REG_4__SCAN_IN), .ZN(n10327) );
  AOI221_X1 U11389 ( .B1(SI_1_), .B2(keyinput_f31), .C1(P2_REG3_REG_4__SCAN_IN), .C2(keyinput_f52), .A(n10327), .ZN(n10334) );
  OAI22_X1 U11390 ( .A1(P1_D_REG_3__SCAN_IN), .A2(keyinput_f126), .B1(
        keyinput_f65), .B2(P2_DATAO_REG_31__SCAN_IN), .ZN(n10328) );
  AOI221_X1 U11391 ( .B1(P1_D_REG_3__SCAN_IN), .B2(keyinput_f126), .C1(
        P2_DATAO_REG_31__SCAN_IN), .C2(keyinput_f65), .A(n10328), .ZN(n10333)
         );
  OAI22_X1 U11392 ( .A1(SI_15_), .A2(keyinput_f17), .B1(keyinput_f38), .B2(
        P2_REG3_REG_23__SCAN_IN), .ZN(n10329) );
  AOI221_X1 U11393 ( .B1(SI_15_), .B2(keyinput_f17), .C1(
        P2_REG3_REG_23__SCAN_IN), .C2(keyinput_f38), .A(n10329), .ZN(n10332)
         );
  OAI22_X1 U11394 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(keyinput_f83), .B1(
        keyinput_f53), .B2(P2_REG3_REG_9__SCAN_IN), .ZN(n10330) );
  AOI221_X1 U11395 ( .B1(P2_DATAO_REG_13__SCAN_IN), .B2(keyinput_f83), .C1(
        P2_REG3_REG_9__SCAN_IN), .C2(keyinput_f53), .A(n10330), .ZN(n10331) );
  NAND4_X1 U11396 ( .A1(n10334), .A2(n10333), .A3(n10332), .A4(n10331), .ZN(
        n10481) );
  OAI22_X1 U11397 ( .A1(SI_5_), .A2(keyinput_f27), .B1(P2_REG3_REG_8__SCAN_IN), 
        .B2(keyinput_f43), .ZN(n10335) );
  AOI221_X1 U11398 ( .B1(SI_5_), .B2(keyinput_f27), .C1(keyinput_f43), .C2(
        P2_REG3_REG_8__SCAN_IN), .A(n10335), .ZN(n10360) );
  OAI22_X1 U11399 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(keyinput_f95), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(keyinput_f69), .ZN(n10336) );
  AOI221_X1 U11400 ( .B1(P1_IR_REG_4__SCAN_IN), .B2(keyinput_f95), .C1(
        keyinput_f69), .C2(P2_DATAO_REG_27__SCAN_IN), .A(n10336), .ZN(n10339)
         );
  OAI22_X1 U11401 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput_f87), .B1(
        keyinput_f41), .B2(P2_REG3_REG_19__SCAN_IN), .ZN(n10337) );
  AOI221_X1 U11402 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_f87), .C1(
        P2_REG3_REG_19__SCAN_IN), .C2(keyinput_f41), .A(n10337), .ZN(n10338)
         );
  OAI211_X1 U11403 ( .C1(n5124), .C2(keyinput_f33), .A(n10339), .B(n10338), 
        .ZN(n10340) );
  AOI21_X1 U11404 ( .B1(n5124), .B2(keyinput_f33), .A(n10340), .ZN(n10359) );
  AOI22_X1 U11405 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(keyinput_f116), .B1(
        P1_IR_REG_11__SCAN_IN), .B2(keyinput_f102), .ZN(n10341) );
  OAI221_X1 U11406 ( .B1(P1_IR_REG_25__SCAN_IN), .B2(keyinput_f116), .C1(
        P1_IR_REG_11__SCAN_IN), .C2(keyinput_f102), .A(n10341), .ZN(n10348) );
  AOI22_X1 U11407 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_f36), .B1(
        P1_D_REG_0__SCAN_IN), .B2(keyinput_f123), .ZN(n10342) );
  OAI221_X1 U11408 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .C1(
        P1_D_REG_0__SCAN_IN), .C2(keyinput_f123), .A(n10342), .ZN(n10347) );
  AOI22_X1 U11409 ( .A1(SI_25_), .A2(keyinput_f7), .B1(P1_IR_REG_12__SCAN_IN), 
        .B2(keyinput_f103), .ZN(n10343) );
  OAI221_X1 U11410 ( .B1(SI_25_), .B2(keyinput_f7), .C1(P1_IR_REG_12__SCAN_IN), 
        .C2(keyinput_f103), .A(n10343), .ZN(n10346) );
  AOI22_X1 U11411 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(keyinput_f67), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_f75), .ZN(n10344) );
  OAI221_X1 U11412 ( .B1(P2_DATAO_REG_29__SCAN_IN), .B2(keyinput_f67), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput_f75), .A(n10344), .ZN(n10345)
         );
  NOR4_X1 U11413 ( .A1(n10348), .A2(n10347), .A3(n10346), .A4(n10345), .ZN(
        n10358) );
  AOI22_X1 U11414 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(keyinput_f66), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .ZN(n10349) );
  OAI221_X1 U11415 ( .B1(P2_DATAO_REG_30__SCAN_IN), .B2(keyinput_f66), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_f62), .A(n10349), .ZN(n10356)
         );
  AOI22_X1 U11416 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_f60), .B1(
        P1_D_REG_4__SCAN_IN), .B2(keyinput_f127), .ZN(n10350) );
  OAI221_X1 U11417 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .C1(
        P1_D_REG_4__SCAN_IN), .C2(keyinput_f127), .A(n10350), .ZN(n10355) );
  AOI22_X1 U11418 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(keyinput_f120), .B1(
        P1_IR_REG_23__SCAN_IN), .B2(keyinput_f114), .ZN(n10351) );
  OAI221_X1 U11419 ( .B1(P1_IR_REG_29__SCAN_IN), .B2(keyinput_f120), .C1(
        P1_IR_REG_23__SCAN_IN), .C2(keyinput_f114), .A(n10351), .ZN(n10354) );
  AOI22_X1 U11420 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(keyinput_f82), .B1(
        P1_IR_REG_26__SCAN_IN), .B2(keyinput_f117), .ZN(n10352) );
  OAI221_X1 U11421 ( .B1(P2_DATAO_REG_14__SCAN_IN), .B2(keyinput_f82), .C1(
        P1_IR_REG_26__SCAN_IN), .C2(keyinput_f117), .A(n10352), .ZN(n10353) );
  NOR4_X1 U11422 ( .A1(n10356), .A2(n10355), .A3(n10354), .A4(n10353), .ZN(
        n10357) );
  NAND4_X1 U11423 ( .A1(n10360), .A2(n10359), .A3(n10358), .A4(n10357), .ZN(
        n10480) );
  AOI22_X1 U11424 ( .A1(n10363), .A2(keyinput_f20), .B1(keyinput_f26), .B2(
        n10362), .ZN(n10361) );
  OAI221_X1 U11425 ( .B1(n10363), .B2(keyinput_f20), .C1(n10362), .C2(
        keyinput_f26), .A(n10361), .ZN(n10375) );
  INV_X1 U11426 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10366) );
  AOI22_X1 U11427 ( .A1(n10366), .A2(keyinput_f125), .B1(keyinput_f59), .B2(
        n10365), .ZN(n10364) );
  OAI221_X1 U11428 ( .B1(n10366), .B2(keyinput_f125), .C1(n10365), .C2(
        keyinput_f59), .A(n10364), .ZN(n10374) );
  INV_X1 U11429 ( .A(SI_21_), .ZN(n10369) );
  AOI22_X1 U11430 ( .A1(n10369), .A2(keyinput_f11), .B1(n10368), .B2(
        keyinput_f72), .ZN(n10367) );
  OAI221_X1 U11431 ( .B1(n10369), .B2(keyinput_f11), .C1(n10368), .C2(
        keyinput_f72), .A(n10367), .ZN(n10373) );
  XOR2_X1 U11432 ( .A(n9498), .B(keyinput_f121), .Z(n10371) );
  XNOR2_X1 U11433 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_f110), .ZN(n10370)
         );
  NAND2_X1 U11434 ( .A1(n10371), .A2(n10370), .ZN(n10372) );
  NOR4_X1 U11435 ( .A1(n10375), .A2(n10374), .A3(n10373), .A4(n10372), .ZN(
        n10419) );
  AOI22_X1 U11436 ( .A1(n10377), .A2(keyinput_f79), .B1(n5523), .B2(
        keyinput_f15), .ZN(n10376) );
  OAI221_X1 U11437 ( .B1(n10377), .B2(keyinput_f79), .C1(n5523), .C2(
        keyinput_f15), .A(n10376), .ZN(n10387) );
  AOI22_X1 U11438 ( .A1(n10380), .A2(keyinput_f89), .B1(n10379), .B2(
        keyinput_f19), .ZN(n10378) );
  OAI221_X1 U11439 ( .B1(n10380), .B2(keyinput_f89), .C1(n10379), .C2(
        keyinput_f19), .A(n10378), .ZN(n10386) );
  XNOR2_X1 U11440 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_f98), .ZN(n10384) );
  XNOR2_X1 U11441 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_f113), .ZN(n10383)
         );
  XNOR2_X1 U11442 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_f112), .ZN(n10382)
         );
  XNOR2_X1 U11443 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_f96), .ZN(n10381) );
  NAND4_X1 U11444 ( .A1(n10384), .A2(n10383), .A3(n10382), .A4(n10381), .ZN(
        n10385) );
  NOR3_X1 U11445 ( .A1(n10387), .A2(n10386), .A3(n10385), .ZN(n10418) );
  AOI22_X1 U11446 ( .A1(n10390), .A2(keyinput_f9), .B1(keyinput_f77), .B2(
        n10389), .ZN(n10388) );
  OAI221_X1 U11447 ( .B1(n10390), .B2(keyinput_f9), .C1(n10389), .C2(
        keyinput_f77), .A(n10388), .ZN(n10402) );
  AOI22_X1 U11448 ( .A1(n10392), .A2(keyinput_f4), .B1(keyinput_f63), .B2(
        n5480), .ZN(n10391) );
  OAI221_X1 U11449 ( .B1(n10392), .B2(keyinput_f4), .C1(n5480), .C2(
        keyinput_f63), .A(n10391), .ZN(n10401) );
  AOI22_X1 U11450 ( .A1(n10395), .A2(keyinput_f23), .B1(keyinput_f46), .B2(
        n10394), .ZN(n10393) );
  OAI221_X1 U11451 ( .B1(n10395), .B2(keyinput_f23), .C1(n10394), .C2(
        keyinput_f46), .A(n10393), .ZN(n10400) );
  AOI22_X1 U11452 ( .A1(n10398), .A2(keyinput_f30), .B1(n10397), .B2(
        keyinput_f90), .ZN(n10396) );
  OAI221_X1 U11453 ( .B1(n10398), .B2(keyinput_f30), .C1(n10397), .C2(
        keyinput_f90), .A(n10396), .ZN(n10399) );
  NOR4_X1 U11454 ( .A1(n10402), .A2(n10401), .A3(n10400), .A4(n10399), .ZN(
        n10417) );
  AOI22_X1 U11455 ( .A1(n10404), .A2(keyinput_f12), .B1(keyinput_f35), .B2(
        n5278), .ZN(n10403) );
  OAI221_X1 U11456 ( .B1(n10404), .B2(keyinput_f12), .C1(n5278), .C2(
        keyinput_f35), .A(n10403), .ZN(n10415) );
  AOI22_X1 U11457 ( .A1(n10407), .A2(keyinput_f50), .B1(n10406), .B2(
        keyinput_f100), .ZN(n10405) );
  OAI221_X1 U11458 ( .B1(n10407), .B2(keyinput_f50), .C1(n10406), .C2(
        keyinput_f100), .A(n10405), .ZN(n10414) );
  AOI22_X1 U11459 ( .A1(P2_U3152), .A2(keyinput_f34), .B1(n5675), .B2(
        keyinput_f8), .ZN(n10408) );
  OAI221_X1 U11460 ( .B1(P2_U3152), .B2(keyinput_f34), .C1(n5675), .C2(
        keyinput_f8), .A(n10408), .ZN(n10413) );
  XNOR2_X1 U11461 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_f92), .ZN(n10411) );
  XNOR2_X1 U11462 ( .A(SI_3_), .B(keyinput_f29), .ZN(n10410) );
  NAND2_X1 U11463 ( .A1(n10411), .A2(n10410), .ZN(n10412) );
  NOR4_X1 U11464 ( .A1(n10415), .A2(n10414), .A3(n10413), .A4(n10412), .ZN(
        n10416) );
  NAND4_X1 U11465 ( .A1(n10419), .A2(n10418), .A3(n10417), .A4(n10416), .ZN(
        n10479) );
  AOI22_X1 U11466 ( .A1(n5228), .A2(keyinput_f49), .B1(n10421), .B2(
        keyinput_f124), .ZN(n10420) );
  OAI221_X1 U11467 ( .B1(n5228), .B2(keyinput_f49), .C1(n10421), .C2(
        keyinput_f124), .A(n10420), .ZN(n10432) );
  AOI22_X1 U11468 ( .A1(n10424), .A2(keyinput_f57), .B1(n10423), .B2(
        keyinput_f10), .ZN(n10422) );
  OAI221_X1 U11469 ( .B1(n10424), .B2(keyinput_f57), .C1(n10423), .C2(
        keyinput_f10), .A(n10422), .ZN(n10431) );
  AOI22_X1 U11470 ( .A1(n10426), .A2(keyinput_f68), .B1(keyinput_f42), .B2(
        n5834), .ZN(n10425) );
  OAI221_X1 U11471 ( .B1(n10426), .B2(keyinput_f68), .C1(n5834), .C2(
        keyinput_f42), .A(n10425), .ZN(n10430) );
  AOI22_X1 U11472 ( .A1(n10428), .A2(keyinput_f5), .B1(n6238), .B2(
        keyinput_f107), .ZN(n10427) );
  OAI221_X1 U11473 ( .B1(n10428), .B2(keyinput_f5), .C1(n6238), .C2(
        keyinput_f107), .A(n10427), .ZN(n10429) );
  NOR4_X1 U11474 ( .A1(n10432), .A2(n10431), .A3(n10430), .A4(n10429), .ZN(
        n10477) );
  AOI22_X1 U11475 ( .A1(n10434), .A2(keyinput_f74), .B1(keyinput_f58), .B2(
        n5375), .ZN(n10433) );
  OAI221_X1 U11476 ( .B1(n10434), .B2(keyinput_f74), .C1(n5375), .C2(
        keyinput_f58), .A(n10433), .ZN(n10446) );
  AOI22_X1 U11477 ( .A1(n10437), .A2(keyinput_f71), .B1(keyinput_f48), .B2(
        n10436), .ZN(n10435) );
  OAI221_X1 U11478 ( .B1(n10437), .B2(keyinput_f71), .C1(n10436), .C2(
        keyinput_f48), .A(n10435), .ZN(n10445) );
  AOI22_X1 U11479 ( .A1(n5841), .A2(keyinput_f97), .B1(keyinput_f32), .B2(
        n10439), .ZN(n10438) );
  OAI221_X1 U11480 ( .B1(n5841), .B2(keyinput_f97), .C1(n10439), .C2(
        keyinput_f32), .A(n10438), .ZN(n10444) );
  INV_X1 U11481 ( .A(SI_29_), .ZN(n10441) );
  AOI22_X1 U11482 ( .A1(n10442), .A2(keyinput_f37), .B1(keyinput_f3), .B2(
        n10441), .ZN(n10440) );
  OAI221_X1 U11483 ( .B1(n10442), .B2(keyinput_f37), .C1(n10441), .C2(
        keyinput_f3), .A(n10440), .ZN(n10443) );
  NOR4_X1 U11484 ( .A1(n10446), .A2(n10445), .A3(n10444), .A4(n10443), .ZN(
        n10476) );
  AOI22_X1 U11485 ( .A1(n10449), .A2(keyinput_f70), .B1(keyinput_f44), .B2(
        n10448), .ZN(n10447) );
  OAI221_X1 U11486 ( .B1(n10449), .B2(keyinput_f70), .C1(n10448), .C2(
        keyinput_f44), .A(n10447), .ZN(n10461) );
  AOI22_X1 U11487 ( .A1(n10452), .A2(keyinput_f99), .B1(keyinput_f76), .B2(
        n10451), .ZN(n10450) );
  OAI221_X1 U11488 ( .B1(n10452), .B2(keyinput_f99), .C1(n10451), .C2(
        keyinput_f76), .A(n10450), .ZN(n10460) );
  AOI22_X1 U11489 ( .A1(n10455), .A2(keyinput_f16), .B1(keyinput_f81), .B2(
        n10454), .ZN(n10453) );
  OAI221_X1 U11490 ( .B1(n10455), .B2(keyinput_f16), .C1(n10454), .C2(
        keyinput_f81), .A(n10453), .ZN(n10459) );
  XNOR2_X1 U11491 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_f105), .ZN(n10457)
         );
  XNOR2_X1 U11492 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_f85), .ZN(n10456) );
  NAND2_X1 U11493 ( .A1(n10457), .A2(n10456), .ZN(n10458) );
  NOR4_X1 U11494 ( .A1(n10461), .A2(n10460), .A3(n10459), .A4(n10458), .ZN(
        n10475) );
  AOI22_X1 U11495 ( .A1(n10463), .A2(keyinput_f86), .B1(keyinput_f56), .B2(
        n5428), .ZN(n10462) );
  OAI221_X1 U11496 ( .B1(n10463), .B2(keyinput_f86), .C1(n5428), .C2(
        keyinput_f56), .A(n10462), .ZN(n10473) );
  AOI22_X1 U11497 ( .A1(n4717), .A2(keyinput_f111), .B1(keyinput_f73), .B2(
        n10465), .ZN(n10464) );
  OAI221_X1 U11498 ( .B1(n4717), .B2(keyinput_f111), .C1(n10465), .C2(
        keyinput_f73), .A(n10464), .ZN(n10472) );
  XOR2_X1 U11499 ( .A(n10466), .B(keyinput_f14), .Z(n10470) );
  XNOR2_X1 U11500 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_f61), .ZN(n10469)
         );
  XNOR2_X1 U11501 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_f91), .ZN(n10468) );
  XNOR2_X1 U11502 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_f106), .ZN(n10467)
         );
  NAND4_X1 U11503 ( .A1(n10470), .A2(n10469), .A3(n10468), .A4(n10467), .ZN(
        n10471) );
  NOR3_X1 U11504 ( .A1(n10473), .A2(n10472), .A3(n10471), .ZN(n10474) );
  NAND4_X1 U11505 ( .A1(n10477), .A2(n10476), .A3(n10475), .A4(n10474), .ZN(
        n10478) );
  NOR4_X1 U11506 ( .A1(n10481), .A2(n10480), .A3(n10479), .A4(n10478), .ZN(
        n10482) );
  AOI22_X1 U11507 ( .A1(n10483), .A2(n10482), .B1(keyinput_f22), .B2(SI_10_), 
        .ZN(n10484) );
  OAI21_X1 U11508 ( .B1(keyinput_f22), .B2(SI_10_), .A(n10484), .ZN(n10485) );
  OAI21_X1 U11509 ( .B1(SI_10_), .B2(keyinput_g22), .A(n10485), .ZN(n10486) );
  AOI211_X1 U11510 ( .C1(SI_10_), .C2(keyinput_g22), .A(n10487), .B(n10486), 
        .ZN(n10493) );
  OAI21_X1 U11511 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10488), .ZN(n10505) );
  NOR2_X1 U11512 ( .A1(n10506), .A2(n10505), .ZN(n10489) );
  NAND2_X1 U11513 ( .A1(n10506), .A2(n10505), .ZN(n10504) );
  OAI21_X1 U11514 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n10489), .A(n10504), 
        .ZN(n10491) );
  XNOR2_X1 U11515 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n10490) );
  XNOR2_X1 U11516 ( .A(n10491), .B(n10490), .ZN(n10492) );
  XNOR2_X1 U11517 ( .A(n10493), .B(n10492), .ZN(ADD_1071_U4) );
  AOI21_X1 U11518 ( .B1(n10496), .B2(n10495), .A(n10494), .ZN(ADD_1071_U47) );
  XNOR2_X1 U11519 ( .A(n10498), .B(n10497), .ZN(ADD_1071_U49) );
  XOR2_X1 U11520 ( .A(n10500), .B(n10499), .Z(ADD_1071_U54) );
  NOR2_X1 U11521 ( .A1(n10502), .A2(n10501), .ZN(n10503) );
  XOR2_X1 U11522 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10503), .Z(ADD_1071_U51) );
  OAI21_X1 U11523 ( .B1(n10506), .B2(n10505), .A(n10504), .ZN(n10507) );
  XNOR2_X1 U11524 ( .A(n10507), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XNOR2_X1 U11525 ( .A(n10509), .B(n10508), .ZN(ADD_1071_U48) );
  XNOR2_X1 U11526 ( .A(n10511), .B(n10510), .ZN(ADD_1071_U50) );
  XOR2_X1 U11527 ( .A(n10513), .B(n10512), .Z(ADD_1071_U53) );
  XNOR2_X1 U11528 ( .A(n10515), .B(n10514), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U5465 ( .A(n8406), .Z(n9927) );
endmodule

