

module b21_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024;

  INV_X4 U5137 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  AND2_X4 U5138 ( .A1(n7300), .A2(n6661), .ZN(n6719) );
  CLKBUF_X2 U5139 ( .A(n6212), .Z(n5096) );
  INV_X1 U5140 ( .A(n6761), .ZN(n6706) );
  INV_X1 U5141 ( .A(n6137), .ZN(n6262) );
  NAND2_X1 U5142 ( .A1(n5724), .A2(n9918), .ZN(n6137) );
  INV_X1 U5143 ( .A(n9689), .ZN(n5358) );
  BUF_X2 U5144 ( .A(n6602), .Z(n5072) );
  INV_X1 U5145 ( .A(n5096), .ZN(n5271) );
  INV_X2 U5146 ( .A(n6261), .ZN(n6246) );
  OR2_X1 U5147 ( .A1(n9781), .A2(n9508), .ZN(n6364) );
  AND3_X1 U5148 ( .A1(n5820), .A2(n5819), .A3(n5818), .ZN(n10802) );
  OR2_X1 U5149 ( .A1(n10252), .A2(n10476), .ZN(n10243) );
  NAND2_X2 U5150 ( .A1(n7202), .A2(n7264), .ZN(n7263) );
  NAND2_X1 U5152 ( .A1(n6084), .A2(n6282), .ZN(n9742) );
  INV_X1 U5153 ( .A(n10794), .ZN(n10289) );
  INV_X1 U5154 ( .A(n9296), .ZN(n6602) );
  AOI21_X2 U5155 ( .B1(n10267), .B2(n9249), .A(n9248), .ZN(n10259) );
  AOI21_X2 U5156 ( .B1(n10280), .B2(n9247), .A(n9246), .ZN(n10267) );
  AOI21_X2 U5157 ( .B1(n9574), .B2(n6409), .A(n6408), .ZN(n9562) );
  NAND2_X2 U5158 ( .A1(n9587), .A2(n9588), .ZN(n9574) );
  XNOR2_X1 U5159 ( .A(n6678), .B(P1_IR_REG_19__SCAN_IN), .ZN(n10794) );
  XNOR2_X2 U5160 ( .A(n6676), .B(n8590), .ZN(n8630) );
  XNOR2_X1 U5161 ( .A(n6735), .B(n6736), .ZN(n9128) );
  NAND2_X1 U5162 ( .A1(n5891), .A2(n5890), .ZN(n10865) );
  OR2_X1 U5163 ( .A1(n10739), .A2(n7893), .ZN(n10776) );
  INV_X2 U5164 ( .A(n10439), .ZN(n5074) );
  INV_X2 U5165 ( .A(n7154), .ZN(n6752) );
  NAND2_X1 U5166 ( .A1(n6749), .A2(n6748), .ZN(n10720) );
  NAND2_X2 U5167 ( .A1(n7692), .A2(n7693), .ZN(n7154) );
  CLKBUF_X2 U5168 ( .A(n6754), .Z(n9196) );
  INV_X4 U5169 ( .A(n9295), .ZN(n7957) );
  NAND2_X1 U5170 ( .A1(n6723), .A2(n5094), .ZN(n6735) );
  INV_X2 U5171 ( .A(n6319), .ZN(n6417) );
  INV_X1 U5173 ( .A(n8630), .ZN(n9187) );
  CLKBUF_X2 U5174 ( .A(n6762), .Z(n8942) );
  CLKBUF_X2 U5175 ( .A(n6740), .Z(n6781) );
  NOR2_X1 U5176 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5091) );
  OR2_X1 U5177 ( .A1(n6470), .A2(n7782), .ZN(n5706) );
  OR2_X1 U5178 ( .A1(n5419), .A2(n5418), .ZN(n5417) );
  NOR4_X1 U5179 ( .A1(n9184), .A2(n9187), .A3(n9181), .A4(n9180), .ZN(n9182)
         );
  OR2_X1 U5180 ( .A1(n10189), .A2(n10195), .ZN(n5318) );
  AOI22_X1 U5181 ( .A1(n9029), .A2(n9031), .B1(n9028), .B2(n9164), .ZN(n9184)
         );
  OAI21_X1 U5182 ( .B1(n9017), .B2(n5093), .A(n9114), .ZN(n5092) );
  AND3_X1 U5183 ( .A1(n9015), .A2(n10171), .A3(n9014), .ZN(n9017) );
  NAND2_X1 U5184 ( .A1(n5480), .A2(n9220), .ZN(n10311) );
  AOI21_X1 U5185 ( .B1(n9648), .B2(n9640), .A(n6145), .ZN(n9621) );
  OAI211_X1 U5186 ( .C1(n5084), .C2(n5083), .A(n10205), .B(n9011), .ZN(n9012)
         );
  NAND2_X1 U5187 ( .A1(n9159), .A2(n9033), .ZN(n5093) );
  NAND2_X1 U5188 ( .A1(n9009), .A2(n10217), .ZN(n5083) );
  AOI21_X1 U5189 ( .B1(n5085), .B2(n9007), .A(n9010), .ZN(n5084) );
  NAND2_X1 U5190 ( .A1(n7108), .A2(n7107), .ZN(n10476) );
  NOR2_X1 U5191 ( .A1(n9768), .A2(n9769), .ZN(n5467) );
  NAND2_X1 U5192 ( .A1(n5078), .A2(n5077), .ZN(n8977) );
  NOR2_X1 U5193 ( .A1(n9236), .A2(n9235), .ZN(n10421) );
  NAND2_X1 U5194 ( .A1(n6088), .A2(n6087), .ZN(n9868) );
  OR2_X1 U5195 ( .A1(n8676), .A2(n6341), .ZN(n10921) );
  NAND2_X1 U5196 ( .A1(n6975), .A2(n6974), .ZN(n10413) );
  OR2_X1 U5197 ( .A1(n7992), .A2(n9125), .ZN(n8121) );
  AND2_X1 U5198 ( .A1(n8975), .A2(n9134), .ZN(n5077) );
  NAND2_X1 U5199 ( .A1(n6077), .A2(n5359), .ZN(n7843) );
  NAND2_X1 U5200 ( .A1(n5970), .A2(n5969), .ZN(n8857) );
  INV_X1 U5201 ( .A(n10883), .ZN(n5075) );
  NAND2_X1 U5202 ( .A1(n6937), .A2(n6936), .ZN(n9210) );
  NAND2_X1 U5203 ( .A1(n5956), .A2(n5955), .ZN(n8858) );
  NAND2_X1 U5204 ( .A1(n5877), .A2(n5876), .ZN(n10852) );
  NAND2_X1 U5205 ( .A1(n5086), .A2(n9089), .ZN(n7981) );
  NAND2_X1 U5206 ( .A1(n10742), .A2(n9123), .ZN(n5086) );
  OAI211_X1 U5207 ( .C1(n7263), .C2(n7508), .A(n6827), .B(n6826), .ZN(n8105)
         );
  AOI21_X1 U5208 ( .B1(n5920), .B2(n5919), .A(n5918), .ZN(n5925) );
  NAND2_X1 U5209 ( .A1(n5087), .A2(n9086), .ZN(n10742) );
  AND2_X2 U5210 ( .A1(n7996), .A2(n10907), .ZN(n10439) );
  AND2_X1 U5211 ( .A1(n6747), .A2(n5703), .ZN(n6748) );
  OAI21_X1 U5212 ( .B1(n5792), .B2(n5539), .A(n5102), .ZN(n5834) );
  NOR2_X1 U5213 ( .A1(n7643), .A2(n7801), .ZN(n7865) );
  NAND4_X1 U5214 ( .A1(n6804), .A2(n6803), .A3(n6802), .A4(n6801), .ZN(n10101)
         );
  NAND4_X1 U5215 ( .A1(n6745), .A2(n6744), .A3(n6743), .A4(n6742), .ZN(n7642)
         );
  NAND4_X1 U5216 ( .A1(n6766), .A2(n6765), .A3(n6764), .A4(n6763), .ZN(n10103)
         );
  OR2_X1 U5217 ( .A1(n6746), .A2(n7323), .ZN(n5478) );
  AND3_X1 U5218 ( .A1(n6725), .A2(n6724), .A3(n5095), .ZN(n5094) );
  NAND2_X1 U5219 ( .A1(n5767), .A2(n5766), .ZN(n5778) );
  CLKBUF_X1 U5220 ( .A(n6741), .Z(n8941) );
  NAND2_X2 U5221 ( .A1(n7263), .A2(n5740), .ZN(n8949) );
  XNOR2_X1 U5222 ( .A(n6284), .B(n6283), .ZN(n6286) );
  NAND2_X1 U5223 ( .A1(n10543), .A2(n9271), .ZN(n6741) );
  INV_X1 U5224 ( .A(n6667), .ZN(n10543) );
  AND2_X1 U5225 ( .A1(n5762), .A2(n5745), .ZN(n5746) );
  NAND2_X1 U5226 ( .A1(n9920), .A2(n8925), .ZN(n7372) );
  XNOR2_X1 U5227 ( .A(n5081), .B(P1_IR_REG_29__SCAN_IN), .ZN(n6667) );
  NAND2_X1 U5228 ( .A1(n6664), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5081) );
  INV_X2 U5229 ( .A(n10538), .ZN(n8088) );
  OAI21_X1 U5230 ( .B1(n6652), .B2(n6642), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5401) );
  OR2_X1 U5231 ( .A1(n5117), .A2(n6652), .ZN(n6664) );
  INV_X2 U5232 ( .A(n9910), .ZN(n5076) );
  AND2_X1 U5233 ( .A1(n5473), .A2(n5534), .ZN(n5280) );
  NOR2_X1 U5234 ( .A1(n5720), .A2(n5719), .ZN(n5473) );
  AND2_X1 U5235 ( .A1(n6461), .A2(n5721), .ZN(n5722) );
  NAND2_X1 U5236 ( .A1(n5739), .A2(n5738), .ZN(n5386) );
  AND2_X1 U5237 ( .A1(n5503), .A2(n8595), .ZN(n5082) );
  AND3_X2 U5238 ( .A1(n5582), .A2(n5583), .A3(n5580), .ZN(n6681) );
  INV_X1 U5239 ( .A(n5675), .ZN(n5535) );
  NAND2_X1 U5240 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n6643), .ZN(n6644) );
  AND2_X1 U5241 ( .A1(n6639), .A2(n6786), .ZN(n5583) );
  AND3_X1 U5242 ( .A1(n5735), .A2(n5713), .A3(n5710), .ZN(n5534) );
  NAND2_X1 U5243 ( .A1(n5306), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n5737) );
  NAND2_X1 U5244 ( .A1(n5308), .A2(n5307), .ZN(n5739) );
  AND4_X1 U5245 ( .A1(n5091), .A2(n5090), .A3(n5089), .A4(n5088), .ZN(n5582)
         );
  AND2_X1 U5246 ( .A1(n6727), .A2(n5581), .ZN(n5580) );
  NOR2_X1 U5247 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5088) );
  NOR2_X1 U5248 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5089) );
  NOR2_X1 U5249 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5090) );
  NOR2_X1 U5250 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5718) );
  INV_X1 U5251 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8590) );
  INV_X1 U5252 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8583) );
  NOR2_X2 U5253 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5735) );
  INV_X2 U5254 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X1 U5255 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n6639) );
  INV_X1 U5256 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5738) );
  NOR2_X1 U5257 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n6786) );
  NOR2_X2 U5258 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6727) );
  NAND3_X1 U5259 ( .A1(n5079), .A2(n8972), .A3(n5113), .ZN(n5078) );
  NAND3_X1 U5260 ( .A1(n5080), .A2(n8970), .A3(n9133), .ZN(n5079) );
  OAI21_X1 U5261 ( .B1(n8967), .B2(n8966), .A(n8965), .ZN(n5080) );
  NAND3_X1 U5262 ( .A1(n6681), .A2(n5622), .A3(n5082), .ZN(n6652) );
  NAND3_X1 U5263 ( .A1(n9005), .A2(n9006), .A3(n10266), .ZN(n5085) );
  NAND2_X1 U5264 ( .A1(n9088), .A2(n9127), .ZN(n5087) );
  MUX2_X1 U5265 ( .A(n5092), .B(n9019), .S(n9018), .Z(n9020) );
  NAND3_X1 U5266 ( .A1(n10543), .A2(n9271), .A3(P1_REG0_REG_1__SCAN_IN), .ZN(
        n5095) );
  INV_X2 U5267 ( .A(n6741), .ZN(n7205) );
  NOR3_X4 U5268 ( .A1(n9733), .A2(n5347), .A3(n9861), .ZN(n9682) );
  XNOR2_X2 U5269 ( .A(n6663), .B(n10534), .ZN(n9271) );
  OR2_X1 U5270 ( .A1(n10776), .A2(n10792), .ZN(n10777) );
  OAI211_X2 U5271 ( .C1(n7263), .C2(n7532), .A(n6808), .B(n6807), .ZN(n10792)
         );
  XNOR2_X2 U5272 ( .A(n5401), .B(n8382), .ZN(n7264) );
  INV_X1 U5273 ( .A(n5562), .ZN(n5380) );
  OAI21_X1 U5274 ( .B1(n5564), .B2(n5563), .A(n6022), .ZN(n5562) );
  INV_X1 U5275 ( .A(n6023), .ZN(n5563) );
  NOR2_X1 U5276 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5710) );
  AND2_X1 U5277 ( .A1(n5494), .A2(n5321), .ZN(n5320) );
  NAND2_X1 U5278 ( .A1(n5323), .A2(n5325), .ZN(n5321) );
  NAND2_X1 U5279 ( .A1(n9169), .A2(n9112), .ZN(n7693) );
  OR2_X1 U5280 ( .A1(n10449), .A2(n9016), .ZN(n9114) );
  NAND2_X1 U5281 ( .A1(n6133), .A2(n6132), .ZN(n6150) );
  AOI21_X1 U5282 ( .B1(n5555), .B2(n5557), .A(n5176), .ZN(n5554) );
  NAND2_X1 U5283 ( .A1(n5830), .A2(SI_6_), .ZN(n5846) );
  NAND2_X1 U5284 ( .A1(n7927), .A2(n6476), .ZN(n9296) );
  AND2_X1 U5285 ( .A1(n5724), .A2(n5727), .ZN(n6248) );
  NAND2_X1 U5286 ( .A1(n5206), .A2(n5683), .ZN(n8022) );
  NAND2_X1 U5287 ( .A1(n9799), .A2(n5684), .ZN(n5206) );
  AOI21_X1 U5288 ( .B1(n5684), .B2(n9798), .A(n5137), .ZN(n5683) );
  NAND2_X1 U5289 ( .A1(n6224), .A2(n6223), .ZN(n9819) );
  NAND2_X1 U5290 ( .A1(n8948), .A2(n5271), .ZN(n6224) );
  NAND2_X1 U5291 ( .A1(n6080), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6083) );
  OR2_X1 U5292 ( .A1(n7123), .A2(n7122), .ZN(n5640) );
  OAI21_X1 U5293 ( .B1(n10204), .B2(n9230), .A(n9229), .ZN(n10189) );
  AND2_X1 U5294 ( .A1(n5365), .A2(n6292), .ZN(n5364) );
  OAI21_X1 U5295 ( .B1(n10361), .B2(n5486), .A(n9217), .ZN(n5485) );
  AND2_X1 U5296 ( .A1(n9214), .A2(n9216), .ZN(n5482) );
  INV_X1 U5297 ( .A(n9918), .ZN(n5727) );
  INV_X1 U5298 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5533) );
  NOR2_X1 U5299 ( .A1(n9544), .A2(n5368), .ZN(n5367) );
  INV_X1 U5300 ( .A(n6414), .ZN(n5368) );
  OR2_X1 U5301 ( .A1(n9495), .A2(n9304), .ZN(n6293) );
  OR2_X1 U5302 ( .A1(n9839), .A2(n9518), .ZN(n6395) );
  OR2_X1 U5303 ( .A1(n9883), .A2(n9718), .ZN(n6309) );
  OR2_X1 U5304 ( .A1(n8858), .A2(n9398), .ZN(n6353) );
  OR2_X1 U5305 ( .A1(n10865), .A2(n8677), .ZN(n6338) );
  NAND2_X1 U5306 ( .A1(n7780), .A2(n6317), .ZN(n5443) );
  OR2_X1 U5307 ( .A1(n6246), .A2(n7375), .ZN(n5773) );
  OR2_X1 U5308 ( .A1(n9888), .A2(n9396), .ZN(n9736) );
  NAND2_X1 U5309 ( .A1(n6286), .A2(n9742), .ZN(n6627) );
  NAND2_X1 U5310 ( .A1(n10102), .A2(n6719), .ZN(n6790) );
  INV_X1 U5311 ( .A(n10443), .ZN(n9025) );
  OR2_X1 U5312 ( .A1(n10459), .A2(n10206), .ZN(n9256) );
  OR2_X1 U5313 ( .A1(n10464), .A2(n9971), .ZN(n9073) );
  NAND2_X1 U5314 ( .A1(n10464), .A2(n9971), .ZN(n9254) );
  NAND2_X1 U5315 ( .A1(n5430), .A2(n5428), .ZN(n10203) );
  AOI21_X1 U5316 ( .B1(n5431), .B2(n5433), .A(n5429), .ZN(n5428) );
  INV_X1 U5317 ( .A(n9253), .ZN(n5429) );
  AND2_X1 U5318 ( .A1(n10476), .A2(n9972), .ZN(n9252) );
  OR2_X1 U5319 ( .A1(n10506), .A2(n10315), .ZN(n9038) );
  NAND2_X1 U5320 ( .A1(n10506), .A2(n10315), .ZN(n9242) );
  NOR2_X1 U5321 ( .A1(n10433), .A2(n9210), .ZN(n5400) );
  NAND2_X1 U5322 ( .A1(n5329), .A2(n5115), .ZN(n5328) );
  INV_X1 U5323 ( .A(n10311), .ZN(n5329) );
  OAI21_X1 U5324 ( .B1(n6252), .B2(n8204), .A(n6251), .ZN(n6271) );
  OR2_X1 U5325 ( .A1(n6250), .A2(n6249), .ZN(n6251) );
  XNOR2_X1 U5326 ( .A(n6250), .B(n6249), .ZN(n6252) );
  NAND2_X1 U5327 ( .A1(n5110), .A2(n5380), .ZN(n5376) );
  NAND2_X1 U5328 ( .A1(n5946), .A2(n5379), .ZN(n5378) );
  NAND2_X1 U5329 ( .A1(n5921), .A2(SI_11_), .ZN(n5940) );
  AOI21_X1 U5330 ( .B1(n5100), .B2(n5542), .A(n5150), .ZN(n5541) );
  AOI21_X1 U5331 ( .B1(n5871), .B2(n5548), .A(n5547), .ZN(n5546) );
  INV_X1 U5332 ( .A(n5888), .ZN(n5547) );
  INV_X1 U5333 ( .A(n5866), .ZN(n5548) );
  NAND2_X1 U5334 ( .A1(n5868), .A2(SI_8_), .ZN(n5888) );
  INV_X1 U5335 ( .A(n5249), .ZN(n5247) );
  INV_X1 U5336 ( .A(n5515), .ZN(n5514) );
  AOI21_X1 U5337 ( .B1(n5515), .B2(n5516), .A(n5513), .ZN(n5512) );
  INV_X1 U5338 ( .A(n8661), .ZN(n5513) );
  NAND2_X1 U5339 ( .A1(n7897), .A2(n6509), .ZN(n5260) );
  NAND2_X1 U5340 ( .A1(n6286), .A2(n5106), .ZN(n9295) );
  AND4_X1 U5341 ( .A1(n6144), .A2(n6143), .A3(n6142), .A4(n6141), .ZN(n9512)
         );
  INV_X1 U5342 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5712) );
  NAND2_X1 U5343 ( .A1(n9524), .A2(n9523), .ZN(n9545) );
  NAND2_X1 U5344 ( .A1(n9561), .A2(n9393), .ZN(n6414) );
  OR2_X1 U5345 ( .A1(n9836), .A2(n9614), .ZN(n9575) );
  OR2_X1 U5346 ( .A1(n10974), .A2(n9775), .ZN(n5697) );
  OR2_X1 U5347 ( .A1(n10932), .A2(n9399), .ZN(n5699) );
  NAND2_X1 U5348 ( .A1(n8015), .A2(n8014), .ZN(n9799) );
  INV_X1 U5349 ( .A(n6278), .ZN(n6086) );
  INV_X1 U5350 ( .A(n7372), .ZN(n6085) );
  XNOR2_X1 U5351 ( .A(n5201), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5724) );
  NAND2_X1 U5352 ( .A1(n5202), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5201) );
  NAND2_X1 U5353 ( .A1(n6083), .A2(n6082), .ZN(n6282) );
  OR3_X1 U5354 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n5775) );
  NAND2_X1 U5355 ( .A1(n8099), .A2(n8100), .ZN(n5600) );
  NOR2_X1 U5356 ( .A1(n8099), .A2(n8100), .ZN(n5599) );
  NOR2_X1 U5357 ( .A1(n9996), .A2(n5639), .ZN(n5638) );
  INV_X1 U5358 ( .A(n9941), .ZN(n5639) );
  XNOR2_X1 U5359 ( .A(n7120), .B(n7154), .ZN(n7123) );
  NAND2_X1 U5360 ( .A1(n6668), .A2(n10543), .ZN(n6762) );
  NAND2_X1 U5361 ( .A1(n10190), .A2(n9263), .ZN(n10183) );
  AND2_X1 U5362 ( .A1(n9257), .A2(n9033), .ZN(n10171) );
  INV_X1 U5363 ( .A(n10174), .ZN(n10206) );
  AOI21_X1 U5364 ( .B1(n5494), .B2(n5496), .A(n5170), .ZN(n5493) );
  XNOR2_X1 U5365 ( .A(n10306), .B(n10283), .ZN(n10301) );
  NAND2_X1 U5366 ( .A1(n5412), .A2(n5410), .ZN(n10312) );
  NAND2_X1 U5367 ( .A1(n5411), .A2(n9000), .ZN(n5410) );
  INV_X1 U5368 ( .A(n5413), .ZN(n5411) );
  NOR2_X1 U5369 ( .A1(n10330), .A2(n5415), .ZN(n5414) );
  INV_X1 U5370 ( .A(n9240), .ZN(n5415) );
  INV_X1 U5371 ( .A(n6746), .ZN(n8947) );
  INV_X1 U5372 ( .A(n8949), .ZN(n7029) );
  INV_X1 U5373 ( .A(n10102), .ZN(n10783) );
  OR2_X1 U5374 ( .A1(n10454), .A2(n9232), .ZN(n9257) );
  OAI21_X1 U5375 ( .B1(n6150), .B2(n6149), .A(n6148), .ZN(n6161) );
  NAND2_X1 U5376 ( .A1(n6120), .A2(n6119), .ZN(n6133) );
  OAI21_X1 U5377 ( .B1(n6068), .B2(n5556), .A(n5554), .ZN(n6114) );
  NAND2_X1 U5378 ( .A1(n6068), .A2(n6067), .ZN(n6077) );
  NAND2_X1 U5379 ( .A1(n5568), .A2(n5564), .ZN(n6024) );
  OR2_X1 U5380 ( .A1(n5835), .A2(n5838), .ZN(n5836) );
  NAND2_X1 U5381 ( .A1(n5812), .A2(SI_5_), .ZN(n5838) );
  NAND2_X1 U5382 ( .A1(n7852), .A2(n6504), .ZN(n7898) );
  INV_X1 U5383 ( .A(n9303), .ZN(n5254) );
  NAND2_X1 U5384 ( .A1(n5355), .A2(n5354), .ZN(n5353) );
  NOR2_X1 U5385 ( .A1(n6286), .A2(n8066), .ZN(n5354) );
  XNOR2_X1 U5386 ( .A(n6452), .B(n9742), .ZN(n5355) );
  OR2_X1 U5387 ( .A1(n7408), .A2(n7407), .ZN(n5221) );
  AND2_X1 U5388 ( .A1(n5223), .A2(n5222), .ZN(n7408) );
  NAND2_X1 U5389 ( .A1(n7387), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5222) );
  AOI21_X1 U5390 ( .B1(n10195), .B2(n5317), .A(n5173), .ZN(n5316) );
  INV_X1 U5391 ( .A(n6324), .ZN(n5287) );
  NOR2_X1 U5392 ( .A1(n5300), .A2(n8049), .ZN(n5297) );
  NAND2_X1 U5393 ( .A1(n6337), .A2(n6338), .ZN(n5299) );
  INV_X1 U5394 ( .A(n5300), .ZN(n5298) );
  NOR2_X1 U5395 ( .A1(n6392), .A2(n5305), .ZN(n5304) );
  INV_X1 U5396 ( .A(n9610), .ZN(n5305) );
  NAND2_X1 U5397 ( .A1(n6396), .A2(n9607), .ZN(n6394) );
  INV_X1 U5398 ( .A(n6221), .ZN(n5576) );
  INV_X1 U5399 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5306) );
  INV_X1 U5400 ( .A(n7779), .ZN(n6317) );
  NAND2_X1 U5401 ( .A1(n10983), .A2(n5400), .ZN(n5399) );
  INV_X1 U5402 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5308) );
  INV_X1 U5403 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5307) );
  INV_X1 U5404 ( .A(n9329), .ZN(n5277) );
  INV_X1 U5405 ( .A(n6600), .ZN(n5251) );
  NOR2_X1 U5406 ( .A1(n9498), .A2(n5560), .ZN(n5559) );
  INV_X1 U5407 ( .A(n6279), .ZN(n5560) );
  AND2_X1 U5408 ( .A1(n6430), .A2(n9575), .ZN(n6409) );
  NOR2_X1 U5409 ( .A1(n9836), .A2(n5337), .ZN(n5336) );
  INV_X1 U5410 ( .A(n5338), .ZN(n5337) );
  AND2_X1 U5411 ( .A1(n9576), .A2(n5667), .ZN(n5666) );
  NAND2_X1 U5412 ( .A1(n9588), .A2(n9521), .ZN(n5667) );
  INV_X1 U5413 ( .A(n9521), .ZN(n5668) );
  NAND2_X1 U5414 ( .A1(n9830), .A2(n9565), .ZN(n6429) );
  OR2_X1 U5415 ( .A1(n9830), .A2(n9565), .ZN(n6430) );
  AND2_X1 U5416 ( .A1(n9846), .A2(n9650), .ZN(n9517) );
  OR2_X1 U5417 ( .A1(n9664), .A2(n5696), .ZN(n9624) );
  OR2_X1 U5418 ( .A1(n9851), .A2(n9512), .ZN(n6299) );
  OR2_X1 U5419 ( .A1(n9871), .A2(n9719), .ZN(n6307) );
  NOR2_X1 U5420 ( .A1(n9871), .A2(n9878), .ZN(n5348) );
  OR2_X1 U5421 ( .A1(n9878), .A2(n9395), .ZN(n6375) );
  AND2_X1 U5422 ( .A1(n5157), .A2(n10920), .ZN(n5464) );
  AND2_X1 U5423 ( .A1(n8814), .A2(n5699), .ZN(n5674) );
  NAND2_X1 U5424 ( .A1(n10932), .A2(n5344), .ZN(n5343) );
  INV_X1 U5425 ( .A(n5345), .ZN(n5344) );
  OR2_X1 U5426 ( .A1(n8811), .A2(n10865), .ZN(n5345) );
  NOR2_X1 U5427 ( .A1(n5968), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n6029) );
  INV_X1 U5428 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5677) );
  INV_X1 U5429 ( .A(n7047), .ZN(n5659) );
  XNOR2_X1 U5430 ( .A(n6753), .B(n6752), .ZN(n6755) );
  OAI21_X1 U5431 ( .B1(n8906), .B2(n5605), .A(n5601), .ZN(n6990) );
  AND2_X1 U5432 ( .A1(n5602), .A2(n10023), .ZN(n5601) );
  OR2_X1 U5433 ( .A1(n5603), .A2(n10025), .ZN(n5602) );
  NAND2_X1 U5434 ( .A1(n5103), .A2(n6950), .ZN(n5603) );
  OR2_X1 U5435 ( .A1(n9252), .A2(n9250), .ZN(n5433) );
  INV_X1 U5436 ( .A(n9251), .ZN(n5434) );
  OR2_X1 U5437 ( .A1(n10470), .A2(n10242), .ZN(n9072) );
  NAND2_X1 U5438 ( .A1(n10470), .A2(n10242), .ZN(n9253) );
  INV_X1 U5439 ( .A(n5323), .ZN(n5322) );
  AND2_X1 U5440 ( .A1(n10490), .A2(n10298), .ZN(n9246) );
  OR2_X1 U5441 ( .A1(n10490), .A2(n10298), .ZN(n8959) );
  INV_X1 U5442 ( .A(n5485), .ZN(n5484) );
  OR2_X1 U5443 ( .A1(n10356), .A2(n10371), .ZN(n9240) );
  NAND2_X1 U5444 ( .A1(n10382), .A2(n10384), .ZN(n9215) );
  NOR2_X1 U5445 ( .A1(n10420), .A2(n5491), .ZN(n5490) );
  INV_X1 U5446 ( .A(n9211), .ZN(n5491) );
  AND2_X1 U5447 ( .A1(n10885), .A2(n9048), .ZN(n9236) );
  NOR2_X1 U5448 ( .A1(n9134), .A2(n5502), .ZN(n5501) );
  INV_X1 U5449 ( .A(n8791), .ZN(n5502) );
  OR2_X1 U5450 ( .A1(n8868), .A2(n10890), .ZN(n9053) );
  NAND2_X1 U5451 ( .A1(n8174), .A2(n9100), .ZN(n9151) );
  INV_X1 U5452 ( .A(n10301), .ZN(n5327) );
  NAND2_X1 U5453 ( .A1(n8630), .A2(n5073), .ZN(n9018) );
  OAI21_X1 U5454 ( .B1(n6165), .B2(n5166), .A(n5569), .ZN(n6203) );
  INV_X1 U5455 ( .A(n5570), .ZN(n5569) );
  OAI21_X1 U5456 ( .B1(n5572), .B2(n5166), .A(n6191), .ZN(n5570) );
  NAND2_X1 U5457 ( .A1(n5624), .A2(n6641), .ZN(n5623) );
  AND2_X1 U5458 ( .A1(n5404), .A2(n5625), .ZN(n5624) );
  INV_X1 U5459 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5625) );
  AND2_X1 U5460 ( .A1(n5573), .A2(n6164), .ZN(n5572) );
  INV_X1 U5461 ( .A(n6167), .ZN(n5573) );
  INV_X1 U5462 ( .A(n6113), .ZN(n5552) );
  INV_X1 U5463 ( .A(n6076), .ZN(n5558) );
  INV_X1 U5464 ( .A(n6045), .ZN(n5372) );
  NOR2_X1 U5465 ( .A1(n5977), .A2(n5566), .ZN(n5565) );
  INV_X1 U5466 ( .A(n5966), .ZN(n5566) );
  AND2_X1 U5467 ( .A1(n5567), .A2(n5118), .ZN(n5564) );
  INV_X1 U5468 ( .A(n5980), .ZN(n5567) );
  XNOR2_X1 U5469 ( .A(n5900), .B(SI_9_), .ZN(n5902) );
  NAND2_X1 U5470 ( .A1(n9328), .A2(n9329), .ZN(n9327) );
  OR2_X1 U5471 ( .A1(n6155), .A2(n9278), .ZN(n6173) );
  NAND2_X1 U5472 ( .A1(n5520), .A2(n5519), .ZN(n8134) );
  INV_X1 U5473 ( .A(n8137), .ZN(n5520) );
  INV_X1 U5474 ( .A(n6518), .ZN(n5518) );
  AND4_X1 U5475 ( .A1(n5898), .A2(n5897), .A3(n5896), .A4(n5895), .ZN(n8677)
         );
  NAND2_X1 U5476 ( .A1(n5760), .A2(n5214), .ZN(n5213) );
  NAND2_X1 U5477 ( .A1(n6262), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5214) );
  OR2_X1 U5478 ( .A1(n6175), .A2(n10701), .ZN(n5728) );
  NAND2_X1 U5479 ( .A1(n5735), .A2(n5710), .ZN(n5798) );
  AND2_X1 U5480 ( .A1(n5238), .A2(n5237), .ZN(n7516) );
  NAND2_X1 U5481 ( .A1(n7514), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5237) );
  OR2_X1 U5482 ( .A1(n7590), .A2(n7589), .ZN(n5227) );
  AND2_X1 U5483 ( .A1(n5227), .A2(n5226), .ZN(n7711) );
  NAND2_X1 U5484 ( .A1(n7709), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5226) );
  OR2_X1 U5485 ( .A1(n7711), .A2(n7710), .ZN(n5225) );
  NAND2_X1 U5486 ( .A1(n9472), .A2(n9471), .ZN(n9478) );
  NOR2_X1 U5487 ( .A1(n9534), .A2(n9503), .ZN(n9502) );
  NAND2_X1 U5488 ( .A1(n6241), .A2(n6240), .ZN(n9495) );
  AOI21_X1 U5489 ( .B1(n5367), .B2(n9563), .A(n5136), .ZN(n5365) );
  INV_X1 U5490 ( .A(n5367), .ZN(n5366) );
  AND2_X1 U5491 ( .A1(n6293), .A2(n6292), .ZN(n9528) );
  NOR2_X1 U5492 ( .A1(n9556), .A2(n9819), .ZN(n9546) );
  XNOR2_X1 U5493 ( .A(n9819), .B(n9566), .ZN(n9544) );
  NAND2_X1 U5494 ( .A1(n9562), .A2(n9554), .ZN(n9568) );
  NAND2_X1 U5495 ( .A1(n6430), .A2(n6429), .ZN(n9576) );
  NAND2_X1 U5496 ( .A1(n9602), .A2(n9519), .ZN(n9586) );
  AND3_X1 U5497 ( .A1(n6188), .A2(n6187), .A3(n6186), .ZN(n9614) );
  OAI21_X1 U5498 ( .B1(n9675), .B2(n5114), .A(n5679), .ZN(n9602) );
  INV_X1 U5499 ( .A(n5680), .ZN(n5679) );
  OAI21_X1 U5500 ( .B1(n5114), .B2(n5682), .A(n5681), .ZN(n5680) );
  INV_X1 U5501 ( .A(n9609), .ZN(n5681) );
  OR2_X1 U5502 ( .A1(n5696), .A2(n9515), .ZN(n9626) );
  NAND2_X1 U5503 ( .A1(n5448), .A2(n6304), .ZN(n5447) );
  INV_X1 U5504 ( .A(n5451), .ZN(n5448) );
  AOI21_X1 U5505 ( .B1(n5453), .B2(n5452), .A(n9676), .ZN(n5451) );
  INV_X1 U5506 ( .A(n5454), .ZN(n5452) );
  NAND2_X1 U5507 ( .A1(n5453), .A2(n6304), .ZN(n5449) );
  AND2_X1 U5508 ( .A1(n5358), .A2(n5356), .ZN(n5454) );
  OR2_X1 U5509 ( .A1(n5357), .A2(n6075), .ZN(n5356) );
  NAND2_X1 U5510 ( .A1(n9721), .A2(n5707), .ZN(n9700) );
  AOI211_X1 U5511 ( .C1(n9757), .C2(n9736), .A(n6041), .B(n6040), .ZN(n6043)
         );
  NOR2_X1 U5512 ( .A1(n9733), .A2(n9878), .ZN(n9714) );
  AND2_X1 U5513 ( .A1(n9883), .A2(n9759), .ZN(n9509) );
  NAND2_X1 U5514 ( .A1(n6375), .A2(n6374), .ZN(n9722) );
  NAND2_X1 U5515 ( .A1(n5672), .A2(n5670), .ZN(n9721) );
  AND2_X1 U5516 ( .A1(n9722), .A2(n5671), .ZN(n5670) );
  INV_X1 U5517 ( .A(n9509), .ZN(n5671) );
  AND2_X1 U5518 ( .A1(n6309), .A2(n6308), .ZN(n9743) );
  AND2_X1 U5519 ( .A1(n9736), .A2(n6368), .ZN(n9756) );
  OAI21_X1 U5520 ( .B1(n10915), .B2(n5210), .A(n5207), .ZN(n9749) );
  INV_X1 U5521 ( .A(n5211), .ZN(n5210) );
  AND2_X1 U5522 ( .A1(n5208), .A2(n5687), .ZN(n5207) );
  NAND2_X1 U5523 ( .A1(n5688), .A2(n5691), .ZN(n5687) );
  NAND2_X1 U5524 ( .A1(n5989), .A2(n5988), .ZN(n9781) );
  AND2_X1 U5525 ( .A1(n6364), .A2(n6365), .ZN(n9766) );
  NOR2_X1 U5526 ( .A1(n9766), .A2(n5690), .ZN(n5689) );
  INV_X1 U5527 ( .A(n5697), .ZN(n5690) );
  AND2_X1 U5528 ( .A1(n8860), .A2(n8859), .ZN(n8862) );
  AND4_X1 U5529 ( .A1(n5998), .A2(n5997), .A3(n5996), .A4(n5995), .ZN(n9508)
         );
  NAND2_X1 U5530 ( .A1(n5157), .A2(n5109), .ZN(n5463) );
  NAND2_X1 U5531 ( .A1(n10921), .A2(n5464), .ZN(n5462) );
  NAND2_X1 U5532 ( .A1(n10915), .A2(n5674), .ZN(n8860) );
  AND2_X1 U5533 ( .A1(n6353), .A2(n6354), .ZN(n8817) );
  NAND2_X1 U5534 ( .A1(n10916), .A2(n10919), .ZN(n10915) );
  NOR2_X1 U5535 ( .A1(n8683), .A2(n5345), .ZN(n10931) );
  AOI21_X1 U5536 ( .B1(n8045), .B2(n5887), .A(n5469), .ZN(n5708) );
  INV_X1 U5537 ( .A(n5470), .ZN(n5469) );
  AOI21_X1 U5538 ( .B1(n8021), .B2(n5472), .A(n5471), .ZN(n5470) );
  AND4_X1 U5539 ( .A1(n5886), .A2(n5885), .A3(n5884), .A4(n5883), .ZN(n8648)
         );
  AOI21_X1 U5540 ( .B1(n7936), .B2(n5823), .A(n5141), .ZN(n9786) );
  INV_X1 U5541 ( .A(n9774), .ZN(n10924) );
  NAND2_X1 U5542 ( .A1(n7921), .A2(n7920), .ZN(n7952) );
  NAND2_X1 U5543 ( .A1(n7952), .A2(n7951), .ZN(n7950) );
  OR2_X1 U5544 ( .A1(n10729), .A2(n7781), .ZN(n7769) );
  AND2_X1 U5545 ( .A1(n5857), .A2(n5856), .ZN(n10834) );
  INV_X1 U5546 ( .A(n6458), .ZN(n5475) );
  NOR3_X1 U5547 ( .A1(n5968), .A2(n5532), .A3(P2_IR_REG_12__SCAN_IN), .ZN(
        n6052) );
  NAND2_X1 U5548 ( .A1(n5534), .A2(n5535), .ZN(n5874) );
  INV_X1 U5549 ( .A(n5600), .ZN(n5594) );
  NAND2_X1 U5550 ( .A1(n6771), .A2(n6770), .ZN(n9093) );
  AND2_X1 U5551 ( .A1(n6769), .A2(n5702), .ZN(n6770) );
  AOI21_X1 U5552 ( .B1(n5658), .B2(n5660), .A(n5657), .ZN(n5656) );
  INV_X1 U5553 ( .A(n10014), .ZN(n5657) );
  NAND2_X1 U5554 ( .A1(n7027), .A2(n10052), .ZN(n5662) );
  INV_X1 U5555 ( .A(n8886), .ZN(n5589) );
  NAND2_X1 U5556 ( .A1(n5635), .A2(n7105), .ZN(n5632) );
  INV_X1 U5557 ( .A(n9996), .ZN(n5635) );
  AND2_X1 U5558 ( .A1(n6994), .A2(n6995), .ZN(n5620) );
  NOR2_X1 U5559 ( .A1(n7106), .A2(n7104), .ZN(n9939) );
  NAND2_X1 U5560 ( .A1(n6719), .A2(n7643), .ZN(n6716) );
  AND2_X1 U5561 ( .A1(n6721), .A2(n6720), .ZN(n7583) );
  NAND2_X1 U5562 ( .A1(n6754), .A2(n7643), .ZN(n6721) );
  INV_X1 U5563 ( .A(n5661), .ZN(n5660) );
  OR2_X1 U5564 ( .A1(n10025), .A2(n5606), .ZN(n5605) );
  INV_X1 U5565 ( .A(n6950), .ZN(n5606) );
  AND2_X1 U5566 ( .A1(n6968), .A2(n6969), .ZN(n10025) );
  OR2_X1 U5567 ( .A1(n5608), .A2(n5103), .ZN(n5607) );
  AND2_X1 U5568 ( .A1(n10055), .A2(n10053), .ZN(n7026) );
  NOR2_X1 U5569 ( .A1(n7092), .A2(n7091), .ZN(n10034) );
  NAND2_X1 U5570 ( .A1(n6913), .A2(n8877), .ZN(n5590) );
  AND2_X1 U5571 ( .A1(n6912), .A2(n5592), .ZN(n5591) );
  INV_X1 U5572 ( .A(n7008), .ZN(n5617) );
  NOR2_X1 U5573 ( .A1(n9990), .A2(n6992), .ZN(n5614) );
  NAND2_X1 U5574 ( .A1(n5613), .A2(n5619), .ZN(n5612) );
  INV_X1 U5575 ( .A(n9990), .ZN(n5613) );
  XNOR2_X1 U5576 ( .A(n6830), .B(n7154), .ZN(n8099) );
  AOI21_X1 U5577 ( .B1(n5638), .B2(n7105), .A(n5148), .ZN(n5629) );
  INV_X1 U5578 ( .A(n5640), .ZN(n5636) );
  NAND2_X1 U5579 ( .A1(n5630), .A2(n5629), .ZN(n5628) );
  AND2_X1 U5580 ( .A1(n5632), .A2(n5631), .ZN(n5630) );
  INV_X1 U5581 ( .A(n5638), .ZN(n5631) );
  AOI21_X1 U5582 ( .B1(n10038), .B2(n10035), .A(n10034), .ZN(n7106) );
  OR2_X1 U5583 ( .A1(n9025), .A2(n9024), .ZN(n9179) );
  AND2_X1 U5584 ( .A1(n9112), .A2(n10289), .ZN(n7218) );
  NAND2_X1 U5585 ( .A1(n7205), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6742) );
  NAND2_X1 U5586 ( .A1(n6668), .A2(n6667), .ZN(n6740) );
  AND2_X1 U5587 ( .A1(n7274), .A2(n7275), .ZN(n7486) );
  NOR2_X1 U5588 ( .A1(n7486), .A2(n7485), .ZN(n7484) );
  OR2_X1 U5589 ( .A1(n7314), .A2(n7313), .ZN(n7284) );
  NAND2_X1 U5590 ( .A1(n7965), .A2(n5196), .ZN(n7290) );
  OR2_X1 U5591 ( .A1(n7289), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5196) );
  AND2_X1 U5592 ( .A1(n8934), .A2(n8933), .ZN(n10163) );
  AOI21_X1 U5593 ( .B1(n10203), .B2(n10205), .A(n9255), .ZN(n10196) );
  NAND2_X1 U5594 ( .A1(n5310), .A2(n5309), .ZN(n10204) );
  AOI21_X1 U5595 ( .B1(n5312), .B2(n9115), .A(n5145), .ZN(n5309) );
  NAND2_X1 U5596 ( .A1(n10234), .A2(n5312), .ZN(n5310) );
  AND2_X1 U5597 ( .A1(n9073), .A2(n9254), .ZN(n10205) );
  OR2_X1 U5598 ( .A1(n10259), .A2(n5433), .ZN(n5427) );
  INV_X1 U5599 ( .A(n5432), .ZN(n5431) );
  OAI21_X1 U5600 ( .B1(n5434), .B2(n9252), .A(n10217), .ZN(n5432) );
  INV_X1 U5601 ( .A(n10217), .ZN(n10225) );
  AND2_X1 U5602 ( .A1(n9226), .A2(n10233), .ZN(n9227) );
  AND2_X1 U5603 ( .A1(n9072), .A2(n9253), .ZN(n10217) );
  NAND2_X1 U5604 ( .A1(n10236), .A2(n9070), .ZN(n10250) );
  NAND2_X1 U5605 ( .A1(n8959), .A2(n8958), .ZN(n10281) );
  NAND2_X1 U5606 ( .A1(n5319), .A2(n5323), .ZN(n10278) );
  NAND2_X1 U5607 ( .A1(n10311), .A2(n5326), .ZN(n5319) );
  NAND2_X1 U5608 ( .A1(n10278), .A2(n10281), .ZN(n10277) );
  AND2_X1 U5609 ( .A1(n10317), .A2(n10496), .ZN(n10300) );
  AOI21_X1 U5610 ( .B1(n5414), .B2(n9241), .A(n9243), .ZN(n5413) );
  NAND2_X1 U5611 ( .A1(n9038), .A2(n9242), .ZN(n10330) );
  AND2_X1 U5612 ( .A1(n9240), .A2(n9117), .ZN(n10357) );
  NAND2_X1 U5613 ( .A1(n5438), .A2(n5436), .ZN(n10367) );
  NOR2_X1 U5614 ( .A1(n5437), .A2(n9238), .ZN(n5436) );
  INV_X1 U5615 ( .A(n9239), .ZN(n5437) );
  NAND2_X1 U5616 ( .A1(n9215), .A2(n9214), .ZN(n10362) );
  NAND2_X1 U5617 ( .A1(n6955), .A2(n6954), .ZN(n10433) );
  OAI21_X1 U5618 ( .B1(n10421), .B2(n10419), .A(n10420), .ZN(n10418) );
  AND2_X1 U5619 ( .A1(n9210), .A2(n10888), .ZN(n10419) );
  NAND2_X1 U5620 ( .A1(n9212), .A2(n5490), .ZN(n10426) );
  OAI21_X1 U5621 ( .B1(n8792), .B2(n5499), .A(n5497), .ZN(n8829) );
  INV_X1 U5622 ( .A(n5498), .ZN(n5497) );
  OAI21_X1 U5623 ( .B1(n5501), .B2(n5499), .A(n9118), .ZN(n5498) );
  NAND2_X1 U5624 ( .A1(n5500), .A2(n8827), .ZN(n5499) );
  NAND2_X1 U5625 ( .A1(n8829), .A2(n9137), .ZN(n9212) );
  NAND2_X1 U5626 ( .A1(n8792), .A2(n5501), .ZN(n8828) );
  INV_X1 U5627 ( .A(n10100), .ZN(n10786) );
  INV_X1 U5628 ( .A(n10398), .ZN(n10887) );
  NAND2_X1 U5629 ( .A1(n7162), .A2(n7161), .ZN(n10459) );
  OR2_X1 U5630 ( .A1(n10545), .A2(n6746), .ZN(n7162) );
  NAND2_X1 U5631 ( .A1(n5328), .A2(n5326), .ZN(n10495) );
  NAND2_X1 U5632 ( .A1(n5328), .A2(n9221), .ZN(n10302) );
  CLKBUF_X1 U5633 ( .A(n7692), .Z(n10895) );
  INV_X1 U5634 ( .A(n5441), .ZN(n5440) );
  XNOR2_X1 U5635 ( .A(n6239), .B(n6238), .ZN(n8948) );
  NAND2_X1 U5636 ( .A1(n6222), .A2(n6221), .ZN(n6239) );
  XNOR2_X1 U5637 ( .A(n6203), .B(n6202), .ZN(n9921) );
  XNOR2_X1 U5638 ( .A(n6193), .B(n6192), .ZN(n8841) );
  NAND2_X1 U5639 ( .A1(n6180), .A2(n6179), .ZN(n6193) );
  NAND2_X1 U5640 ( .A1(n6659), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6674) );
  NAND2_X1 U5641 ( .A1(n6077), .A2(n6076), .ZN(n6101) );
  NAND2_X1 U5642 ( .A1(n6063), .A2(n6062), .ZN(n6068) );
  OR2_X1 U5643 ( .A1(n6049), .A2(n6048), .ZN(n6063) );
  NAND2_X1 U5644 ( .A1(n5373), .A2(n5376), .ZN(n6046) );
  NAND2_X1 U5645 ( .A1(n5375), .A2(n5374), .ZN(n5373) );
  NAND2_X1 U5646 ( .A1(n5967), .A2(n5565), .ZN(n5568) );
  NAND2_X1 U5647 ( .A1(n5947), .A2(n5946), .ZN(n5967) );
  INV_X1 U5648 ( .A(n5926), .ZN(n5924) );
  AND2_X1 U5649 ( .A1(n5888), .A2(n5870), .ZN(n5871) );
  AND2_X1 U5650 ( .A1(n5866), .A2(n5850), .ZN(n5851) );
  NAND2_X1 U5651 ( .A1(n5852), .A2(n5851), .ZN(n5867) );
  NAND2_X1 U5652 ( .A1(n5537), .A2(n5536), .ZN(n5837) );
  AND2_X1 U5653 ( .A1(n5351), .A2(n5833), .ZN(n5536) );
  NAND2_X1 U5654 ( .A1(n5792), .A2(n5102), .ZN(n5537) );
  AND2_X1 U5655 ( .A1(n5846), .A2(n5832), .ZN(n5840) );
  AND2_X1 U5656 ( .A1(n5838), .A2(n5815), .ZN(n5704) );
  AND2_X1 U5657 ( .A1(n5795), .A2(n5811), .ZN(n5796) );
  NAND2_X1 U5658 ( .A1(n5746), .A2(n5747), .ZN(n5763) );
  NOR2_X1 U5659 ( .A1(n5255), .A2(n5247), .ZN(n5246) );
  NAND2_X1 U5660 ( .A1(n9301), .A2(n9391), .ZN(n5253) );
  NAND2_X1 U5661 ( .A1(n5254), .A2(n5247), .ZN(n5244) );
  NAND2_X1 U5662 ( .A1(n6124), .A2(n6123), .ZN(n9856) );
  OAI21_X1 U5663 ( .B1(n8137), .B2(n5514), .A(n5512), .ZN(n6525) );
  NAND2_X1 U5664 ( .A1(n6171), .A2(n6170), .ZN(n9839) );
  OR2_X1 U5665 ( .A1(n8773), .A2(n5096), .ZN(n6171) );
  INV_X1 U5666 ( .A(n9407), .ZN(n8148) );
  INV_X1 U5667 ( .A(n8857), .ZN(n10974) );
  AND4_X1 U5668 ( .A1(n5964), .A2(n5963), .A3(n5962), .A4(n5961), .ZN(n9398)
         );
  NAND2_X1 U5669 ( .A1(n6009), .A2(n6008), .ZN(n9888) );
  OR2_X1 U5670 ( .A1(n7613), .A2(n5096), .ZN(n6009) );
  AND4_X1 U5671 ( .A1(n5975), .A2(n5974), .A3(n5973), .A4(n5972), .ZN(n9775)
         );
  AND4_X1 U5672 ( .A1(n5939), .A2(n5938), .A3(n5937), .A4(n5936), .ZN(n9399)
         );
  NAND4_X1 U5673 ( .A1(n5810), .A2(n5809), .A3(n5808), .A4(n5807), .ZN(n9789)
         );
  AND3_X1 U5674 ( .A1(n5736), .A2(n5235), .A3(n5234), .ZN(n10648) );
  NAND2_X1 U5675 ( .A1(n5236), .A2(n5723), .ZN(n5235) );
  NAND2_X1 U5676 ( .A1(n5152), .A2(P2_IR_REG_1__SCAN_IN), .ZN(n5234) );
  OR2_X1 U5677 ( .A1(n7430), .A2(n7431), .ZN(n5223) );
  NAND2_X1 U5678 ( .A1(n7389), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5220) );
  AND2_X1 U5679 ( .A1(n5929), .A2(n5907), .ZN(n7824) );
  NAND2_X1 U5680 ( .A1(n9478), .A2(n5230), .ZN(n5229) );
  OR2_X1 U5681 ( .A1(n9479), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5230) );
  AND2_X1 U5682 ( .A1(n6214), .A2(n6213), .ZN(n9561) );
  OR2_X1 U5683 ( .A1(n10545), .A2(n5096), .ZN(n6214) );
  NAND2_X1 U5684 ( .A1(n10818), .A2(n5684), .ZN(n8050) );
  XNOR2_X1 U5685 ( .A(n5339), .B(n5732), .ZN(n8925) );
  NAND2_X1 U5686 ( .A1(n5281), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5339) );
  NOR2_X1 U5687 ( .A1(n5282), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n5279) );
  NAND2_X1 U5688 ( .A1(n6081), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n6084) );
  NAND2_X1 U5689 ( .A1(n8753), .A2(n8947), .ZN(n7094) );
  NAND3_X1 U5690 ( .A1(n5643), .A2(n5642), .A3(n5647), .ZN(n10038) );
  INV_X1 U5691 ( .A(n5648), .ZN(n5647) );
  NAND2_X1 U5692 ( .A1(n7026), .A2(n5649), .ZN(n5643) );
  NAND2_X1 U5693 ( .A1(n7027), .A2(n5645), .ZN(n5642) );
  NAND2_X1 U5694 ( .A1(n8628), .A2(n8947), .ZN(n7078) );
  INV_X1 U5695 ( .A(n10096), .ZN(n10890) );
  NAND2_X1 U5696 ( .A1(n7013), .A2(n7012), .ZN(n10506) );
  OR2_X1 U5697 ( .A1(n7843), .A2(n6746), .ZN(n7013) );
  INV_X1 U5698 ( .A(n10091), .ZN(n10242) );
  INV_X1 U5699 ( .A(n10405), .ZN(n10889) );
  NAND3_X1 U5700 ( .A1(n6785), .A2(n6784), .A3(n6783), .ZN(n10102) );
  NOR2_X1 U5701 ( .A1(n6782), .A2(n5705), .ZN(n6783) );
  XNOR2_X1 U5702 ( .A(n7290), .B(n10111), .ZN(n10106) );
  NOR2_X1 U5703 ( .A1(n10106), .A2(n10390), .ZN(n10105) );
  AND2_X1 U5704 ( .A1(n8931), .A2(n8930), .ZN(n10443) );
  NAND2_X1 U5705 ( .A1(n5318), .A2(n5317), .ZN(n10168) );
  XNOR2_X1 U5706 ( .A(n10204), .B(n10205), .ZN(n10468) );
  OR2_X1 U5707 ( .A1(n8773), .A2(n6746), .ZN(n7108) );
  NAND2_X1 U5708 ( .A1(n7049), .A2(n7048), .ZN(n10306) );
  NAND2_X1 U5709 ( .A1(n6688), .A2(n6687), .ZN(n10395) );
  OR2_X1 U5710 ( .A1(n7613), .A2(n6746), .ZN(n6688) );
  OR2_X1 U5711 ( .A1(n7576), .A2(n6746), .ZN(n6975) );
  NAND2_X1 U5712 ( .A1(n5108), .A2(n10892), .ZN(n5420) );
  AND2_X1 U5713 ( .A1(n5422), .A2(n5332), .ZN(n5419) );
  AND2_X1 U5714 ( .A1(n10451), .A2(n9262), .ZN(n5332) );
  OR2_X1 U5715 ( .A1(n10452), .A2(n10516), .ZN(n5422) );
  NAND2_X1 U5716 ( .A1(n5287), .A2(n7922), .ZN(n5286) );
  NAND2_X1 U5717 ( .A1(n6324), .A2(n5289), .ZN(n5284) );
  NAND2_X1 U5718 ( .A1(n7930), .A2(n9403), .ZN(n5289) );
  NOR2_X1 U5719 ( .A1(n5299), .A2(n5297), .ZN(n5295) );
  NAND2_X1 U5720 ( .A1(n5303), .A2(n6393), .ZN(n6396) );
  OAI21_X1 U5721 ( .B1(n6391), .B2(n9647), .A(n5304), .ZN(n5303) );
  NAND2_X1 U5722 ( .A1(n6411), .A2(n6319), .ZN(n5294) );
  NAND2_X1 U5723 ( .A1(n6412), .A2(n6417), .ZN(n5293) );
  AND2_X1 U5724 ( .A1(n10479), .A2(n10269), .ZN(n9250) );
  OAI21_X1 U5725 ( .B1(n6207), .B2(n5184), .A(n5574), .ZN(n6250) );
  INV_X1 U5726 ( .A(n5575), .ZN(n5574) );
  OAI21_X1 U5727 ( .B1(n5577), .B2(n5184), .A(n6237), .ZN(n5575) );
  INV_X1 U5728 ( .A(n6179), .ZN(n5571) );
  AND2_X1 U5729 ( .A1(n6021), .A2(n6020), .ZN(n6023) );
  INV_X1 U5730 ( .A(n5940), .ZN(n5379) );
  INV_X1 U5731 ( .A(n5902), .ZN(n5543) );
  INV_X1 U5732 ( .A(n5871), .ZN(n5542) );
  NOR2_X1 U5733 ( .A1(n5524), .A2(n5266), .ZN(n5265) );
  INV_X1 U5734 ( .A(n6571), .ZN(n5266) );
  INV_X1 U5735 ( .A(n5525), .ZN(n5524) );
  INV_X1 U5736 ( .A(n5521), .ZN(n5262) );
  AOI21_X1 U5737 ( .B1(n5525), .B2(n5523), .A(n5522), .ZN(n5521) );
  INV_X1 U5738 ( .A(n6581), .ZN(n5522) );
  INV_X1 U5739 ( .A(n9309), .ZN(n5523) );
  AND2_X1 U5740 ( .A1(n9805), .A2(n9498), .ZN(n6287) );
  AND2_X1 U5741 ( .A1(n5363), .A2(n6293), .ZN(n5362) );
  INV_X1 U5742 ( .A(n6291), .ZN(n6447) );
  INV_X1 U5743 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6027) );
  INV_X1 U5744 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6026) );
  NAND2_X1 U5745 ( .A1(n9824), .A2(n9522), .ZN(n6413) );
  NAND2_X1 U5746 ( .A1(n5348), .A2(n5456), .ZN(n5347) );
  AND2_X1 U5747 ( .A1(n5156), .A2(n8859), .ZN(n5211) );
  INV_X1 U5748 ( .A(n5689), .ZN(n5688) );
  NAND2_X1 U5749 ( .A1(n5211), .A2(n5209), .ZN(n5208) );
  INV_X1 U5750 ( .A(n5674), .ZN(n5209) );
  OR2_X1 U5751 ( .A1(n8811), .A2(n8664), .ZN(n6431) );
  INV_X1 U5752 ( .A(n6336), .ZN(n5471) );
  INV_X1 U5753 ( .A(n8004), .ZN(n5472) );
  NOR2_X1 U5754 ( .A1(n9839), .A2(n9846), .ZN(n5338) );
  NAND2_X1 U5755 ( .A1(n9642), .A2(n5336), .ZN(n9591) );
  NAND2_X1 U5756 ( .A1(n10958), .A2(n5342), .ZN(n5341) );
  INV_X1 U5757 ( .A(n5343), .ZN(n5342) );
  OR2_X1 U5758 ( .A1(n7954), .A2(n7935), .ZN(n9791) );
  OR2_X1 U5759 ( .A1(n7931), .A2(n7930), .ZN(n7954) );
  NOR2_X1 U5760 ( .A1(n10698), .A2(n8157), .ZN(n8152) );
  AND2_X1 U5761 ( .A1(n9922), .A2(n6613), .ZN(n7349) );
  NAND2_X1 U5762 ( .A1(n6051), .A2(n5531), .ZN(n5530) );
  NAND2_X1 U5763 ( .A1(n7046), .A2(n9948), .ZN(n5661) );
  NAND2_X1 U5764 ( .A1(n5656), .A2(n5653), .ZN(n5652) );
  INV_X1 U5765 ( .A(n9958), .ZN(n5653) );
  NAND2_X1 U5766 ( .A1(n10459), .A2(n10206), .ZN(n9032) );
  AND2_X1 U5767 ( .A1(n10225), .A2(n5313), .ZN(n5312) );
  NAND2_X1 U5768 ( .A1(n5314), .A2(n9228), .ZN(n5313) );
  INV_X1 U5769 ( .A(n9227), .ZN(n5314) );
  AND2_X1 U5770 ( .A1(n10476), .A2(n10260), .ZN(n9224) );
  NOR2_X1 U5771 ( .A1(n10486), .A2(n9961), .ZN(n9248) );
  INV_X1 U5772 ( .A(n9250), .ZN(n9070) );
  INV_X1 U5773 ( .A(n5495), .ZN(n5494) );
  OAI21_X1 U5774 ( .B1(n10281), .B2(n5496), .A(n9223), .ZN(n5495) );
  OR2_X1 U5775 ( .A1(n10486), .A2(n10284), .ZN(n9223) );
  INV_X1 U5776 ( .A(n9222), .ZN(n5496) );
  AND2_X1 U5777 ( .A1(n8959), .A2(n10279), .ZN(n9247) );
  INV_X1 U5778 ( .A(n9246), .ZN(n8958) );
  AOI21_X1 U5779 ( .B1(n5326), .B2(n5324), .A(n5135), .ZN(n5323) );
  INV_X1 U5780 ( .A(n5115), .ZN(n5324) );
  AND3_X1 U5781 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_REG3_REG_18__SCAN_IN), 
        .A3(n7014), .ZN(n7032) );
  OR2_X1 U5782 ( .A1(n10366), .A2(n9241), .ZN(n5416) );
  INV_X1 U5783 ( .A(n6691), .ZN(n6669) );
  OR2_X1 U5784 ( .A1(n10395), .A2(n10370), .ZN(n9239) );
  INV_X1 U5785 ( .A(n9120), .ZN(n5500) );
  AND2_X1 U5786 ( .A1(n10828), .A2(n5390), .ZN(n5389) );
  OR2_X1 U5787 ( .A1(n8929), .A2(n9186), .ZN(n7222) );
  AND2_X1 U5788 ( .A1(n5397), .A2(n11004), .ZN(n5396) );
  INV_X1 U5789 ( .A(n5399), .ZN(n5397) );
  NOR2_X1 U5790 ( .A1(n10883), .A2(n5399), .ZN(n10408) );
  NAND2_X1 U5791 ( .A1(n8128), .A2(n10828), .ZN(n8181) );
  NOR2_X1 U5792 ( .A1(n6642), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n5441) );
  AND2_X1 U5793 ( .A1(n5578), .A2(n6206), .ZN(n5577) );
  INV_X1 U5794 ( .A(n6209), .ZN(n5578) );
  INV_X1 U5795 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8591) );
  INV_X1 U5796 ( .A(n5623), .ZN(n5621) );
  INV_X1 U5797 ( .A(n5941), .ZN(n5375) );
  INV_X1 U5798 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6640) );
  NAND2_X1 U5799 ( .A1(n5942), .A2(SI_12_), .ZN(n5966) );
  NAND2_X1 U5800 ( .A1(n5796), .A2(n5538), .ZN(n5352) );
  INV_X1 U5801 ( .A(n5791), .ZN(n5538) );
  AND2_X1 U5802 ( .A1(n5704), .A2(n5840), .ZN(n5833) );
  INV_X1 U5803 ( .A(SI_6_), .ZN(n8443) );
  INV_X1 U5804 ( .A(n5796), .ZN(n5539) );
  NAND2_X1 U5805 ( .A1(n5737), .A2(n5138), .ZN(n5383) );
  NAND2_X1 U5806 ( .A1(n5579), .A2(SI_2_), .ZN(n5777) );
  OAI21_X1 U5807 ( .B1(n9355), .B2(n5264), .A(n5261), .ZN(n6584) );
  AOI21_X1 U5808 ( .B1(n5265), .B2(n5263), .A(n5262), .ZN(n5261) );
  INV_X1 U5809 ( .A(n5265), .ZN(n5264) );
  INV_X1 U5810 ( .A(n9354), .ZN(n5263) );
  AOI21_X1 U5811 ( .B1(n5506), .B2(n5107), .A(n5144), .ZN(n5276) );
  AND2_X1 U5812 ( .A1(n5250), .A2(n5179), .ZN(n5249) );
  NAND2_X1 U5813 ( .A1(n9293), .A2(n5251), .ZN(n5250) );
  OR2_X1 U5814 ( .A1(n8777), .A2(n8778), .ZN(n8775) );
  NOR2_X1 U5815 ( .A1(n9339), .A2(n5510), .ZN(n5509) );
  INV_X1 U5816 ( .A(n6555), .ZN(n5510) );
  AOI21_X1 U5817 ( .B1(n5276), .B2(n5507), .A(n5274), .ZN(n5273) );
  INV_X1 U5818 ( .A(n9284), .ZN(n5274) );
  OR2_X1 U5819 ( .A1(n6138), .A2(n9363), .ZN(n6155) );
  NOR2_X1 U5820 ( .A1(n9361), .A2(n5526), .ZN(n5525) );
  INV_X1 U5821 ( .A(n6575), .ZN(n5526) );
  NAND2_X1 U5822 ( .A1(n9310), .A2(n9309), .ZN(n5527) );
  AOI21_X1 U5823 ( .B1(n8136), .B2(n5517), .A(n5151), .ZN(n5515) );
  OR2_X1 U5824 ( .A1(n6595), .A2(n9318), .ZN(n9378) );
  OAI21_X1 U5825 ( .B1(n6427), .B2(n6426), .A(n6425), .ZN(n6468) );
  AOI21_X1 U5826 ( .B1(n5291), .B2(n5129), .A(n5290), .ZN(n6426) );
  AND3_X1 U5827 ( .A1(n6178), .A2(n6177), .A3(n6176), .ZN(n9518) );
  AND4_X1 U5828 ( .A1(n6061), .A2(n6060), .A3(n6059), .A4(n6058), .ZN(n9395)
         );
  AND4_X1 U5829 ( .A1(n6019), .A2(n6018), .A3(n6017), .A4(n6016), .ZN(n9396)
         );
  INV_X1 U5830 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5236) );
  OR2_X1 U5831 ( .A1(n7454), .A2(n7453), .ZN(n5238) );
  OR2_X1 U5832 ( .A1(n5953), .A2(n5952), .ZN(n5968) );
  NOR2_X1 U5833 ( .A1(n9468), .A2(n5231), .ZN(n9472) );
  AND2_X1 U5834 ( .A1(n9469), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5231) );
  NAND2_X1 U5835 ( .A1(n6254), .A2(n6253), .ZN(n9503) );
  AND2_X1 U5836 ( .A1(n9642), .A2(n5112), .ZN(n9580) );
  NAND2_X1 U5837 ( .A1(n5664), .A2(n5663), .ZN(n9555) );
  AOI21_X1 U5838 ( .B1(n5666), .B2(n5668), .A(n5167), .ZN(n5663) );
  NAND2_X1 U5839 ( .A1(n9586), .A2(n5666), .ZN(n5664) );
  AND2_X1 U5840 ( .A1(n6227), .A2(n6197), .ZN(n9581) );
  AND3_X1 U5841 ( .A1(n6159), .A2(n6158), .A3(n6157), .ZN(n9613) );
  AND2_X1 U5842 ( .A1(n5160), .A2(n9511), .ZN(n5682) );
  AND2_X1 U5843 ( .A1(n6395), .A2(n6294), .ZN(n9609) );
  AND2_X1 U5844 ( .A1(n9516), .A2(n9626), .ZN(n9625) );
  NAND2_X1 U5845 ( .A1(n9642), .A2(n9635), .ZN(n9630) );
  AND2_X1 U5846 ( .A1(n6300), .A2(n9610), .ZN(n9628) );
  NOR2_X1 U5847 ( .A1(n5449), .A2(n5101), .ZN(n5445) );
  OAI21_X1 U5848 ( .B1(n5447), .B2(n5101), .A(n5146), .ZN(n5444) );
  INV_X1 U5849 ( .A(n9708), .ZN(n5446) );
  NAND2_X1 U5850 ( .A1(n9675), .A2(n9511), .ZN(n9656) );
  NAND2_X1 U5851 ( .A1(n9677), .A2(n9676), .ZN(n9675) );
  OR2_X1 U5852 ( .A1(n6056), .A2(n9451), .ZN(n6091) );
  AOI21_X1 U5853 ( .B1(n9700), .B2(n9707), .A(n5698), .ZN(n9688) );
  NOR2_X1 U5854 ( .A1(n9733), .A2(n5346), .ZN(n9701) );
  INV_X1 U5855 ( .A(n5348), .ZN(n5346) );
  AND4_X1 U5856 ( .A1(n6039), .A2(n6038), .A3(n6037), .A4(n6036), .ZN(n9718)
         );
  OR2_X1 U5857 ( .A1(n9780), .A2(n9888), .ZN(n9750) );
  OR3_X1 U5858 ( .A1(n5992), .A2(n8288), .A3(n5991), .ZN(n6013) );
  NAND2_X1 U5859 ( .A1(n5958), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5992) );
  INV_X1 U5860 ( .A(n5959), .ZN(n5958) );
  NOR2_X1 U5861 ( .A1(n8853), .A2(n8857), .ZN(n9778) );
  AND2_X1 U5862 ( .A1(n5466), .A2(n5468), .ZN(n10918) );
  NAND2_X1 U5863 ( .A1(n10921), .A2(n10920), .ZN(n5466) );
  NAND2_X1 U5864 ( .A1(n5205), .A2(n5678), .ZN(n8673) );
  AOI21_X1 U5865 ( .B1(n5097), .B2(n8021), .A(n5139), .ZN(n5678) );
  NAND2_X1 U5866 ( .A1(n8022), .A2(n5097), .ZN(n5205) );
  OR2_X1 U5867 ( .A1(n5893), .A2(n8493), .ZN(n5911) );
  NAND2_X1 U5868 ( .A1(n5708), .A2(n5899), .ZN(n8651) );
  NOR2_X1 U5869 ( .A1(n9791), .A2(n9796), .ZN(n9792) );
  NAND2_X1 U5870 ( .A1(n9786), .A2(n5845), .ZN(n8045) );
  INV_X1 U5871 ( .A(n8018), .ZN(n5685) );
  INV_X1 U5872 ( .A(n6320), .ZN(n5442) );
  NAND2_X1 U5873 ( .A1(n6321), .A2(n6320), .ZN(n7779) );
  INV_X1 U5874 ( .A(n7327), .ZN(n5272) );
  AND4_X1 U5875 ( .A1(n5774), .A2(n5773), .A3(n5772), .A4(n5771), .ZN(n8147)
         );
  NAND2_X1 U5876 ( .A1(n9534), .A2(n5350), .ZN(n9816) );
  INV_X1 U5877 ( .A(n9561), .ZN(n9824) );
  INV_X1 U5878 ( .A(n10995), .ZN(n10972) );
  NAND2_X1 U5879 ( .A1(n10850), .A2(n5097), .ZN(n8670) );
  INV_X1 U5880 ( .A(n10989), .ZN(n10851) );
  INV_X1 U5881 ( .A(n8157), .ZN(n10730) );
  NAND2_X1 U5882 ( .A1(n5283), .A2(n5732), .ZN(n5695) );
  NOR2_X1 U5883 ( .A1(n5695), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U5884 ( .A1(n5733), .A2(n5283), .ZN(n5282) );
  INV_X1 U5885 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5732) );
  NAND2_X1 U5886 ( .A1(n5280), .A2(n5125), .ZN(n6458) );
  AND3_X1 U5887 ( .A1(n5217), .A2(n5216), .A3(n5215), .ZN(n6461) );
  INV_X1 U5888 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5215) );
  OAI21_X1 U5889 ( .B1(n5968), .B2(n5528), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6079) );
  NAND2_X1 U5890 ( .A1(n6028), .A2(n5529), .ZN(n5528) );
  NOR2_X1 U5891 ( .A1(n5530), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n5529) );
  NOR2_X1 U5892 ( .A1(n5798), .A2(n5676), .ZN(n5828) );
  NAND2_X1 U5893 ( .A1(n5677), .A2(n5711), .ZN(n5676) );
  OR2_X1 U5894 ( .A1(n6899), .A2(n7315), .ZN(n6920) );
  XNOR2_X1 U5895 ( .A(n6774), .B(n7154), .ZN(n6775) );
  NAND2_X1 U5896 ( .A1(n9093), .A2(n9192), .ZN(n6772) );
  OR2_X1 U5897 ( .A1(n6872), .A2(n6871), .ZN(n6899) );
  AOI21_X1 U5898 ( .B1(n8757), .B2(n6890), .A(n5140), .ZN(n10002) );
  NAND2_X1 U5899 ( .A1(n8757), .A2(n6865), .ZN(n10003) );
  AND2_X1 U5900 ( .A1(n7060), .A2(n7061), .ZN(n10013) );
  NOR2_X1 U5901 ( .A1(n5652), .A2(n5646), .ZN(n5645) );
  INV_X1 U5902 ( .A(n10052), .ZN(n5646) );
  INV_X1 U5903 ( .A(n5652), .ZN(n5649) );
  OAI21_X1 U5904 ( .B1(n5652), .B2(n5658), .A(n9956), .ZN(n5648) );
  OR2_X1 U5905 ( .A1(n6746), .A2(n7327), .ZN(n6747) );
  AND2_X1 U5906 ( .A1(n6760), .A2(n6759), .ZN(n10046) );
  AND2_X1 U5907 ( .A1(n7580), .A2(n10531), .ZN(n7200) );
  NAND2_X1 U5908 ( .A1(n9187), .A2(n9169), .ZN(n8929) );
  NOR2_X1 U5909 ( .A1(n6741), .A2(n6780), .ZN(n6782) );
  NOR2_X1 U5910 ( .A1(n10629), .A2(n10630), .ZN(n10628) );
  NOR2_X1 U5911 ( .A1(n10628), .A2(n5193), .ZN(n10666) );
  NOR2_X1 U5912 ( .A1(n10625), .A2(n7272), .ZN(n5193) );
  NOR2_X1 U5913 ( .A1(n7498), .A2(n7497), .ZN(n7496) );
  NOR2_X1 U5914 ( .A1(n7496), .A2(n5195), .ZN(n7537) );
  AND2_X1 U5915 ( .A1(n7281), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5195) );
  NAND2_X1 U5916 ( .A1(n7537), .A2(n7538), .ZN(n7536) );
  NAND2_X1 U5917 ( .A1(n7536), .A2(n5194), .ZN(n7550) );
  OR2_X1 U5918 ( .A1(n7542), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5194) );
  NOR2_X1 U5919 ( .A1(n7565), .A2(n7564), .ZN(n7563) );
  NAND2_X1 U5920 ( .A1(n7624), .A2(n7286), .ZN(n7623) );
  AND2_X1 U5921 ( .A1(n7623), .A2(n5198), .ZN(n7757) );
  NAND2_X1 U5922 ( .A1(n7636), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5198) );
  NOR2_X1 U5923 ( .A1(n7757), .A2(n7756), .ZN(n7755) );
  AND2_X1 U5924 ( .A1(n9231), .A2(n5119), .ZN(n5317) );
  NOR2_X1 U5925 ( .A1(n10209), .A2(n10459), .ZN(n10190) );
  NAND2_X1 U5926 ( .A1(n5403), .A2(n5402), .ZN(n10209) );
  OR2_X1 U5927 ( .A1(n10479), .A2(n10269), .ZN(n10236) );
  OR2_X1 U5928 ( .A1(n9115), .A2(n9224), .ZN(n10240) );
  NOR2_X1 U5929 ( .A1(n10479), .A2(n5393), .ZN(n5391) );
  NAND2_X1 U5930 ( .A1(n10317), .A2(n5104), .ZN(n10288) );
  NOR2_X1 U5931 ( .A1(n10312), .A2(n9244), .ZN(n10295) );
  AND2_X1 U5932 ( .A1(n10336), .A2(n10319), .ZN(n10317) );
  NAND2_X1 U5933 ( .A1(n10327), .A2(n10330), .ZN(n5480) );
  NOR2_X2 U5934 ( .A1(n10353), .A2(n10506), .ZN(n10336) );
  NAND2_X1 U5935 ( .A1(n5416), .A2(n9240), .ZN(n10329) );
  AND2_X1 U5936 ( .A1(n5416), .A2(n5414), .ZN(n10328) );
  INV_X1 U5937 ( .A(n6999), .ZN(n7014) );
  INV_X1 U5938 ( .A(n5488), .ZN(n5487) );
  OAI22_X1 U5939 ( .A1(n5490), .A2(n5489), .B1(n10425), .B2(n10983), .ZN(n5488) );
  NAND2_X1 U5940 ( .A1(n5134), .A2(n9213), .ZN(n5489) );
  AND2_X1 U5941 ( .A1(n5438), .A2(n9060), .ZN(n10383) );
  OR2_X1 U5942 ( .A1(n6957), .A2(n6956), .ZN(n6977) );
  INV_X1 U5943 ( .A(n5438), .ZN(n10400) );
  NOR2_X1 U5944 ( .A1(n10883), .A2(n5398), .ZN(n10428) );
  INV_X1 U5945 ( .A(n5400), .ZN(n5398) );
  INV_X1 U5946 ( .A(n10093), .ZN(n10425) );
  AND2_X1 U5947 ( .A1(n9059), .A2(n9237), .ZN(n10420) );
  NOR2_X1 U5948 ( .A1(n6920), .A2(n6919), .ZN(n6938) );
  AOI21_X1 U5949 ( .B1(n8634), .B2(n5122), .A(n5424), .ZN(n10885) );
  NAND2_X1 U5950 ( .A1(n5425), .A2(n9045), .ZN(n5424) );
  NAND2_X1 U5951 ( .A1(n9134), .A2(n8973), .ZN(n5425) );
  INV_X1 U5952 ( .A(n10094), .ZN(n10888) );
  NAND2_X1 U5953 ( .A1(n8828), .A2(n8827), .ZN(n10882) );
  AND3_X1 U5954 ( .A1(n5389), .A2(n8128), .A3(n5387), .ZN(n10884) );
  NOR2_X1 U5955 ( .A1(n8868), .A2(n8637), .ZN(n5387) );
  NAND2_X1 U5956 ( .A1(n8128), .A2(n5388), .ZN(n8640) );
  AND2_X1 U5957 ( .A1(n10843), .A2(n10828), .ZN(n5388) );
  AND2_X1 U5958 ( .A1(n9102), .A2(n8173), .ZN(n9125) );
  AND3_X1 U5959 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6819) );
  NOR2_X2 U5960 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5404) );
  AND2_X1 U5961 ( .A1(n9114), .A2(n9159), .ZN(n9258) );
  NAND2_X1 U5962 ( .A1(n8939), .A2(n8938), .ZN(n10449) );
  INV_X1 U5963 ( .A(n10413), .ZN(n10983) );
  XNOR2_X1 U5964 ( .A(n6271), .B(n6269), .ZN(n8932) );
  XNOR2_X1 U5965 ( .A(n6252), .B(SI_29_), .ZN(n9916) );
  NAND2_X1 U5966 ( .A1(n6652), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6655) );
  INV_X1 U5967 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5581) );
  NOR2_X2 U5968 ( .A1(n5623), .A2(n5116), .ZN(n5622) );
  AND2_X1 U5969 ( .A1(n6640), .A2(n8591), .ZN(n5503) );
  INV_X1 U5970 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8595) );
  NAND2_X1 U5971 ( .A1(n5557), .A2(n6113), .ZN(n5553) );
  INV_X1 U5972 ( .A(n5551), .ZN(n5550) );
  OAI21_X1 U5973 ( .B1(n5554), .B2(n5552), .A(n5174), .ZN(n5551) );
  XNOR2_X1 U5974 ( .A(n6674), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9169) );
  NAND2_X1 U5975 ( .A1(n5369), .A2(n5370), .ZN(n6049) );
  AOI21_X1 U5976 ( .B1(n5371), .B2(n5377), .A(n5177), .ZN(n5370) );
  AND2_X1 U5977 ( .A1(n6681), .A2(n6640), .ZN(n6648) );
  NAND2_X1 U5978 ( .A1(n5940), .A2(n5923), .ZN(n5926) );
  NOR2_X1 U5979 ( .A1(n5917), .A2(SI_10_), .ZN(n5918) );
  NAND2_X1 U5980 ( .A1(n5544), .A2(n5546), .ZN(n5903) );
  NAND2_X1 U5981 ( .A1(n5545), .A2(n5871), .ZN(n5544) );
  INV_X1 U5982 ( .A(n5867), .ZN(n5545) );
  NAND2_X1 U5983 ( .A1(n5779), .A2(SI_3_), .ZN(n5791) );
  NAND2_X1 U5984 ( .A1(n5778), .A2(n5777), .ZN(n5783) );
  OAI21_X1 U5985 ( .B1(n5579), .B2(SI_2_), .A(n5777), .ZN(n5765) );
  NAND2_X1 U5986 ( .A1(n5763), .A2(n5762), .ZN(n5767) );
  OR2_X1 U5987 ( .A1(n6621), .A2(n9391), .ZN(n5701) );
  XNOR2_X1 U5988 ( .A(n6584), .B(n6582), .ZN(n9277) );
  NAND2_X1 U5989 ( .A1(n8134), .A2(n6518), .ZN(n8162) );
  XNOR2_X1 U5990 ( .A(n6485), .B(n6486), .ZN(n7819) );
  NAND2_X1 U5991 ( .A1(n7820), .A2(n7819), .ZN(n7818) );
  OAI21_X1 U5992 ( .B1(n7898), .B2(n7897), .A(n6509), .ZN(n8115) );
  NAND2_X1 U5993 ( .A1(n5301), .A2(n5123), .ZN(n7771) );
  NAND2_X1 U5994 ( .A1(n5267), .A2(n6571), .ZN(n9310) );
  NAND2_X1 U5995 ( .A1(n9355), .A2(n9354), .ZN(n5267) );
  NAND2_X1 U5996 ( .A1(n5242), .A2(n7721), .ZN(n7732) );
  NAND2_X1 U5997 ( .A1(n7818), .A2(n5240), .ZN(n5242) );
  NOR2_X1 U5998 ( .A1(n7722), .A2(n5241), .ZN(n5240) );
  INV_X1 U5999 ( .A(n6488), .ZN(n5241) );
  NAND2_X1 U6000 ( .A1(n9327), .A2(n5509), .ZN(n9342) );
  NAND2_X1 U6001 ( .A1(n9327), .A2(n6555), .ZN(n9338) );
  NAND2_X1 U6002 ( .A1(n7818), .A2(n6488), .ZN(n7725) );
  OAI21_X1 U6003 ( .B1(n7898), .B2(n5259), .A(n5256), .ZN(n8137) );
  AOI21_X1 U6004 ( .B1(n5258), .B2(n5257), .A(n5143), .ZN(n5256) );
  INV_X1 U6005 ( .A(n6509), .ZN(n5257) );
  NAND2_X1 U6006 ( .A1(n5527), .A2(n6575), .ZN(n9362) );
  NAND2_X1 U6007 ( .A1(n6135), .A2(n6134), .ZN(n9851) );
  NAND2_X1 U6008 ( .A1(n5511), .A2(n5515), .ZN(n8662) );
  NAND2_X1 U6009 ( .A1(n8137), .A2(n5517), .ZN(n5511) );
  NAND2_X1 U6010 ( .A1(n9342), .A2(n9337), .ZN(n9370) );
  INV_X1 U6011 ( .A(n8147), .ZN(n9404) );
  NOR2_X1 U6012 ( .A1(n5132), .A2(n5213), .ZN(n5212) );
  NAND4_X1 U6013 ( .A1(n5731), .A2(n5730), .A3(n5729), .A4(n5728), .ZN(n9407)
         );
  NOR2_X1 U6014 ( .A1(n7463), .A2(n5169), .ZN(n7419) );
  NOR2_X1 U6015 ( .A1(n7419), .A2(n7418), .ZN(n7417) );
  NAND2_X1 U6016 ( .A1(n5233), .A2(n5232), .ZN(n7394) );
  NAND2_X1 U6017 ( .A1(n7391), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5232) );
  INV_X1 U6018 ( .A(n7417), .ZN(n5233) );
  AND2_X1 U6019 ( .A1(n7450), .A2(n5239), .ZN(n7454) );
  NAND2_X1 U6020 ( .A1(n7451), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5239) );
  INV_X1 U6021 ( .A(n5238), .ZN(n7513) );
  NOR2_X1 U6022 ( .A1(n5675), .A2(n5798), .ZN(n5854) );
  INV_X1 U6023 ( .A(n5227), .ZN(n7708) );
  INV_X1 U6024 ( .A(n5225), .ZN(n7823) );
  AND2_X1 U6025 ( .A1(n5225), .A2(n5224), .ZN(n7825) );
  NAND2_X1 U6026 ( .A1(n7824), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5224) );
  INV_X1 U6027 ( .A(n9480), .ZN(n5228) );
  INV_X1 U6028 ( .A(n9495), .ZN(n9815) );
  OAI21_X1 U6029 ( .B1(n9562), .B2(n5366), .A(n5365), .ZN(n9530) );
  NAND2_X1 U6030 ( .A1(n9568), .A2(n6414), .ZN(n9541) );
  NAND2_X1 U6031 ( .A1(n5665), .A2(n9521), .ZN(n9573) );
  NAND2_X1 U6032 ( .A1(n9586), .A2(n9520), .ZN(n5665) );
  INV_X1 U6033 ( .A(n9839), .ZN(n9607) );
  OAI21_X1 U6034 ( .B1(n9708), .B2(n5449), .A(n5447), .ZN(n9665) );
  NAND2_X1 U6035 ( .A1(n6104), .A2(n6103), .ZN(n9861) );
  NAND2_X1 U6036 ( .A1(n5450), .A2(n5453), .ZN(n9672) );
  NAND2_X1 U6037 ( .A1(n9708), .A2(n5454), .ZN(n5450) );
  AOI21_X1 U6038 ( .B1(n9708), .B2(n5357), .A(n6075), .ZN(n9690) );
  NOR2_X1 U6039 ( .A1(n9887), .A2(n9509), .ZN(n9723) );
  NAND2_X1 U6040 ( .A1(n6055), .A2(n6054), .ZN(n9878) );
  INV_X1 U6041 ( .A(n9743), .ZN(n5673) );
  NAND2_X1 U6042 ( .A1(n6032), .A2(n6031), .ZN(n9883) );
  NAND2_X1 U6043 ( .A1(n9507), .A2(n5697), .ZN(n9765) );
  NAND2_X1 U6044 ( .A1(n8862), .A2(n8861), .ZN(n9507) );
  NAND2_X1 U6045 ( .A1(n5462), .A2(n5463), .ZN(n8849) );
  NAND2_X1 U6046 ( .A1(n10915), .A2(n5699), .ZN(n8816) );
  NAND2_X1 U6047 ( .A1(n5932), .A2(n5931), .ZN(n10939) );
  NOR2_X1 U6048 ( .A1(n8683), .A2(n10865), .ZN(n8684) );
  NAND2_X1 U6049 ( .A1(n8020), .A2(n8006), .ZN(n10850) );
  INV_X1 U6050 ( .A(n8022), .ZN(n8020) );
  NAND2_X1 U6051 ( .A1(n8017), .A2(n8016), .ZN(n10818) );
  INV_X1 U6052 ( .A(n9799), .ZN(n8017) );
  NAND2_X1 U6053 ( .A1(n7950), .A2(n7922), .ZN(n8012) );
  AND3_X1 U6054 ( .A1(n5803), .A2(n5802), .A3(n5801), .ZN(n10768) );
  NAND2_X1 U6055 ( .A1(n5270), .A2(n5268), .ZN(n8157) );
  INV_X1 U6056 ( .A(n5269), .ZN(n5268) );
  NAND2_X1 U6057 ( .A1(n5272), .A2(n5271), .ZN(n5270) );
  OAI22_X1 U6058 ( .A1(n6278), .A2(n7322), .B1(n7372), .B2(n7437), .ZN(n5269)
         );
  INV_X1 U6059 ( .A(n7771), .ZN(n10711) );
  NAND2_X1 U6060 ( .A1(n6624), .A2(n7605), .ZN(n10700) );
  INV_X1 U6061 ( .A(n10705), .ZN(n9797) );
  NAND2_X1 U6062 ( .A1(n5218), .A2(n5349), .ZN(n9895) );
  AOI21_X1 U6063 ( .B1(n9814), .B2(n10995), .A(n5219), .ZN(n5218) );
  INV_X1 U6064 ( .A(n9817), .ZN(n5349) );
  OAI21_X1 U6065 ( .B1(n9816), .B2(n10991), .A(n5168), .ZN(n5219) );
  NOR2_X1 U6066 ( .A1(n6458), .A2(n5692), .ZN(n9911) );
  NAND2_X1 U6067 ( .A1(n5694), .A2(n5693), .ZN(n5692) );
  NOR2_X1 U6068 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n5694) );
  INV_X1 U6069 ( .A(n5695), .ZN(n5693) );
  XNOR2_X1 U6070 ( .A(n5199), .B(n5476), .ZN(n9918) );
  INV_X1 U6071 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5476) );
  NAND2_X1 U6072 ( .A1(n5200), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5199) );
  NAND2_X1 U6073 ( .A1(n5475), .A2(n5474), .ZN(n5200) );
  XNOR2_X1 U6074 ( .A(n5734), .B(n5733), .ZN(n9920) );
  OAI21_X1 U6075 ( .B1(n6458), .B2(P2_IR_REG_26__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5734) );
  NAND2_X1 U6076 ( .A1(n6282), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6284) );
  INV_X1 U6077 ( .A(n10648), .ZN(n7386) );
  OR3_X1 U6078 ( .A1(n10549), .A2(n8848), .A3(n8774), .ZN(n7300) );
  NAND2_X1 U6079 ( .A1(n5596), .A2(n5599), .ZN(n5595) );
  AND2_X1 U6080 ( .A1(n8089), .A2(n5600), .ZN(n5598) );
  NOR2_X1 U6081 ( .A1(n7026), .A2(n5655), .ZN(n9951) );
  INV_X1 U6082 ( .A(n5662), .ZN(n5655) );
  NAND2_X1 U6083 ( .A1(n7031), .A2(n7030), .ZN(n10503) );
  NOR2_X1 U6084 ( .A1(n7176), .A2(n5585), .ZN(n5584) );
  INV_X1 U6085 ( .A(n7159), .ZN(n5585) );
  INV_X1 U6086 ( .A(n5656), .ZN(n5651) );
  AND2_X1 U6087 ( .A1(n5644), .A2(n5662), .ZN(n5654) );
  NOR2_X1 U6088 ( .A1(n7026), .A2(n5650), .ZN(n5644) );
  AOI21_X1 U6089 ( .B1(n5591), .B2(n5590), .A(n5589), .ZN(n5588) );
  AND2_X1 U6090 ( .A1(n5637), .A2(n5640), .ZN(n5634) );
  NAND2_X1 U6091 ( .A1(n9938), .A2(n5638), .ZN(n5637) );
  NAND2_X1 U6092 ( .A1(n7125), .A2(n7124), .ZN(n10470) );
  NAND2_X1 U6093 ( .A1(n8841), .A2(n8947), .ZN(n7125) );
  AND2_X1 U6094 ( .A1(n5611), .A2(n5618), .ZN(n9989) );
  INV_X1 U6095 ( .A(n9225), .ZN(n10269) );
  AND2_X1 U6096 ( .A1(n9938), .A2(n9941), .ZN(n5633) );
  AOI21_X1 U6097 ( .B1(n9951), .B2(n7047), .A(n5660), .ZN(n10017) );
  NAND2_X1 U6098 ( .A1(n5607), .A2(n5604), .ZN(n5709) );
  INV_X1 U6099 ( .A(n5605), .ZN(n5604) );
  OR2_X1 U6100 ( .A1(n6911), .A2(n5591), .ZN(n5587) );
  NAND2_X1 U6101 ( .A1(n6918), .A2(n6917), .ZN(n8962) );
  NAND2_X1 U6102 ( .A1(n5610), .A2(n5609), .ZN(n10055) );
  AND2_X1 U6103 ( .A1(n5612), .A2(n5616), .ZN(n5609) );
  NAND2_X1 U6104 ( .A1(n5617), .A2(n7007), .ZN(n5616) );
  AND2_X1 U6105 ( .A1(n7204), .A2(n10405), .ZN(n10081) );
  INV_X1 U6106 ( .A(n9930), .ZN(n10083) );
  AOI21_X1 U6107 ( .B1(n7106), .B2(n5629), .A(n5627), .ZN(n5626) );
  NAND2_X1 U6108 ( .A1(n5628), .A2(n5641), .ZN(n5627) );
  NAND2_X1 U6109 ( .A1(n9968), .A2(n9967), .ZN(n5641) );
  NAND2_X1 U6110 ( .A1(n9921), .A2(n8947), .ZN(n7142) );
  INV_X1 U6111 ( .A(n10089), .ZN(n10069) );
  AND2_X1 U6112 ( .A1(n7204), .A2(n10398), .ZN(n10086) );
  NAND4_X1 U6113 ( .A1(n6839), .A2(n6838), .A3(n6837), .A4(n6836), .ZN(n10099)
         );
  OR2_X1 U6114 ( .A1(n6740), .A2(n10657), .ZN(n6744) );
  OR2_X1 U6115 ( .A1(n6762), .A2(n7272), .ZN(n6725) );
  OR2_X1 U6116 ( .A1(n6740), .A2(n10624), .ZN(n6724) );
  OR2_X1 U6117 ( .A1(n6740), .A2(n8622), .ZN(n6709) );
  OR2_X1 U6118 ( .A1(n6762), .A2(n6705), .ZN(n6710) );
  NOR2_X1 U6119 ( .A1(n7484), .A2(n5120), .ZN(n7675) );
  NOR2_X1 U6120 ( .A1(n7563), .A2(n5197), .ZN(n7314) );
  AND2_X1 U6121 ( .A1(n7567), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5197) );
  INV_X1 U6122 ( .A(n7284), .ZN(n7312) );
  NOR2_X1 U6123 ( .A1(n10105), .A2(n7291), .ZN(n10117) );
  INV_X1 U6124 ( .A(n10163), .ZN(n10444) );
  NAND2_X1 U6125 ( .A1(n5420), .A2(n9262), .ZN(n10448) );
  NAND2_X1 U6126 ( .A1(n8951), .A2(n8950), .ZN(n10454) );
  NAND2_X1 U6127 ( .A1(n8948), .A2(n8947), .ZN(n8951) );
  AND2_X1 U6128 ( .A1(n10176), .A2(n10175), .ZN(n10177) );
  AND2_X1 U6129 ( .A1(n10199), .A2(n10198), .ZN(n10462) );
  INV_X1 U6130 ( .A(n5504), .ZN(n10467) );
  OAI21_X1 U6131 ( .B1(n10468), .B2(n10895), .A(n5505), .ZN(n5504) );
  AOI21_X1 U6132 ( .B1(n10208), .B2(n10892), .A(n10207), .ZN(n5505) );
  NAND2_X1 U6133 ( .A1(n5427), .A2(n5431), .ZN(n10226) );
  NAND2_X1 U6134 ( .A1(n5311), .A2(n9228), .ZN(n10218) );
  NAND2_X1 U6135 ( .A1(n10234), .A2(n9227), .ZN(n5311) );
  NAND2_X1 U6136 ( .A1(n10277), .A2(n9222), .ZN(n10265) );
  NAND2_X1 U6137 ( .A1(n7065), .A2(n7064), .ZN(n10490) );
  OR2_X1 U6138 ( .A1(n8070), .A2(n6746), .ZN(n7065) );
  NAND2_X1 U6139 ( .A1(n10366), .A2(n5414), .ZN(n5409) );
  NAND2_X1 U6140 ( .A1(n6998), .A2(n6997), .ZN(n10356) );
  OR2_X1 U6141 ( .A1(n7706), .A2(n6746), .ZN(n6998) );
  NAND2_X1 U6142 ( .A1(n5483), .A2(n9216), .ZN(n10358) );
  NAND2_X1 U6143 ( .A1(n10362), .A2(n10361), .ZN(n5483) );
  NAND2_X1 U6144 ( .A1(n6651), .A2(n6650), .ZN(n10513) );
  NAND2_X1 U6145 ( .A1(n10426), .A2(n9213), .ZN(n10415) );
  OR2_X1 U6146 ( .A1(n7470), .A2(n6746), .ZN(n6937) );
  NAND2_X1 U6147 ( .A1(n8792), .A2(n8791), .ZN(n8794) );
  NAND2_X1 U6148 ( .A1(n5423), .A2(n9044), .ZN(n8830) );
  NAND2_X1 U6149 ( .A1(n8634), .A2(n5105), .ZN(n5423) );
  NAND2_X1 U6150 ( .A1(n8634), .A2(n9052), .ZN(n8784) );
  NAND2_X1 U6151 ( .A1(n5407), .A2(n9096), .ZN(n10782) );
  OAI21_X1 U6152 ( .B1(n7330), .B2(n6746), .A(n5333), .ZN(n7893) );
  NOR2_X1 U6153 ( .A1(n5128), .A2(n5334), .ZN(n5333) );
  NOR2_X1 U6154 ( .A1(n7263), .A2(n7682), .ZN(n5334) );
  OR2_X1 U6155 ( .A1(n7263), .A2(n10625), .ZN(n5477) );
  AND2_X1 U6156 ( .A1(n5074), .A2(n10791), .ZN(n10432) );
  OR3_X1 U6157 ( .A1(n10500), .A2(n10499), .A3(n10498), .ZN(n10527) );
  XNOR2_X1 U6158 ( .A(n6277), .B(n6276), .ZN(n10539) );
  NAND2_X1 U6159 ( .A1(n6274), .A2(n6273), .ZN(n6277) );
  OR2_X1 U6160 ( .A1(n10533), .A2(n6662), .ZN(n6663) );
  NAND2_X1 U6161 ( .A1(n6222), .A2(n6211), .ZN(n10545) );
  NAND2_X1 U6162 ( .A1(n6180), .A2(n6169), .ZN(n8773) );
  XNOR2_X1 U6163 ( .A(n6161), .B(n6160), .ZN(n8753) );
  NAND2_X1 U6164 ( .A1(n6675), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6676) );
  INV_X1 U6165 ( .A(n9167), .ZN(n9112) );
  NAND2_X1 U6166 ( .A1(n5360), .A2(n5555), .ZN(n5359) );
  INV_X1 U6167 ( .A(n6068), .ZN(n5360) );
  NAND2_X1 U6168 ( .A1(n6005), .A2(n6004), .ZN(n7613) );
  OR2_X1 U6169 ( .A1(n6003), .A2(n6002), .ZN(n6004) );
  NAND2_X1 U6170 ( .A1(n5568), .A2(n5118), .ZN(n5981) );
  NAND2_X1 U6171 ( .A1(n5872), .A2(n5871), .ZN(n5889) );
  AND2_X1 U6172 ( .A1(n5837), .A2(n5836), .ZN(n5847) );
  XNOR2_X1 U6173 ( .A(n5797), .B(n5796), .ZN(n7330) );
  NAND2_X1 U6174 ( .A1(n5792), .A2(n5791), .ZN(n5797) );
  NAND2_X1 U6175 ( .A1(n5254), .A2(n9293), .ZN(n5248) );
  INV_X1 U6176 ( .A(n5223), .ZN(n7429) );
  INV_X1 U6177 ( .A(n5221), .ZN(n7406) );
  XNOR2_X1 U6178 ( .A(n5229), .B(n5228), .ZN(n9494) );
  OAI211_X1 U6179 ( .C1(n5420), .C2(n5418), .A(n5417), .B(n5185), .ZN(P1_U3552) );
  INV_X1 U6180 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5421) );
  NAND2_X1 U6181 ( .A1(n5330), .A2(n5186), .ZN(P1_U3520) );
  NAND2_X1 U6182 ( .A1(n5331), .A2(n11024), .ZN(n5330) );
  NAND2_X1 U6183 ( .A1(n5419), .A2(n5420), .ZN(n5331) );
  AND2_X1 U6184 ( .A1(n8650), .A2(n8649), .ZN(n5097) );
  AND2_X1 U6185 ( .A1(n5456), .A2(n5455), .ZN(n5098) );
  OR2_X2 U6186 ( .A1(n9742), .A2(n6290), .ZN(n6319) );
  OR2_X1 U6187 ( .A1(n6990), .A2(n6989), .ZN(n5099) );
  AND2_X1 U6188 ( .A1(n5546), .A2(n5543), .ZN(n5100) );
  OR2_X1 U6189 ( .A1(n9861), .A2(n9692), .ZN(n6304) );
  AND2_X1 U6190 ( .A1(n9663), .A2(n9673), .ZN(n5101) );
  AND2_X1 U6191 ( .A1(n5352), .A2(n5811), .ZN(n5102) );
  AND2_X1 U6192 ( .A1(n8908), .A2(n6948), .ZN(n5103) );
  AND2_X1 U6193 ( .A1(n10286), .A2(n10496), .ZN(n5104) );
  NAND2_X1 U6194 ( .A1(n5634), .A2(n5124), .ZN(n9966) );
  AND2_X1 U6195 ( .A1(n9052), .A2(n5426), .ZN(n5105) );
  INV_X1 U6196 ( .A(n9798), .ZN(n8016) );
  OR2_X1 U6197 ( .A1(n10476), .A2(n10260), .ZN(n9228) );
  AND2_X1 U6198 ( .A1(n9742), .A2(n10679), .ZN(n5106) );
  INV_X1 U6199 ( .A(n8021), .ZN(n8006) );
  AND2_X1 U6200 ( .A1(n6335), .A2(n6336), .ZN(n8021) );
  OR2_X1 U6201 ( .A1(n5277), .A2(n5508), .ZN(n5107) );
  NAND2_X1 U6202 ( .A1(n6897), .A2(n6896), .ZN(n8868) );
  XOR2_X1 U6203 ( .A(n9259), .B(n9258), .Z(n5108) );
  INV_X1 U6204 ( .A(n5377), .ZN(n5374) );
  NAND2_X1 U6205 ( .A1(n5380), .A2(n5946), .ZN(n5377) );
  NAND2_X1 U6206 ( .A1(n7094), .A2(n7093), .ZN(n10479) );
  OR2_X1 U6207 ( .A1(n10919), .A2(n5465), .ZN(n5109) );
  INV_X1 U6208 ( .A(n8136), .ZN(n5519) );
  NAND2_X1 U6209 ( .A1(n5158), .A2(n5378), .ZN(n5110) );
  OR2_X1 U6210 ( .A1(n5798), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5111) );
  AND2_X1 U6211 ( .A1(n5336), .A2(n5335), .ZN(n5112) );
  INV_X1 U6212 ( .A(n10188), .ZN(n10195) );
  NAND2_X1 U6213 ( .A1(n9256), .A2(n9032), .ZN(n10188) );
  INV_X1 U6214 ( .A(n9868), .ZN(n5456) );
  NAND2_X1 U6215 ( .A1(n7139), .A2(n7138), .ZN(n9967) );
  AND2_X1 U6216 ( .A1(n6076), .A2(n6066), .ZN(n6067) );
  INV_X1 U6217 ( .A(n6067), .ZN(n5555) );
  NAND2_X1 U6218 ( .A1(n6870), .A2(n6869), .ZN(n8790) );
  INV_X1 U6219 ( .A(n8790), .ZN(n5390) );
  NAND2_X1 U6220 ( .A1(n5443), .A2(n5130), .ZN(n7936) );
  INV_X1 U6221 ( .A(n6781), .ZN(n7016) );
  NOR2_X1 U6222 ( .A1(n9051), .A2(n8973), .ZN(n5113) );
  NOR2_X1 U6223 ( .A1(n9517), .A2(n9625), .ZN(n5114) );
  NAND4_X2 U6224 ( .A1(n6707), .A2(n6710), .A3(n6709), .A4(n6708), .ZN(n7643)
         );
  NAND2_X1 U6225 ( .A1(n6991), .A2(n5099), .ZN(n9977) );
  INV_X1 U6226 ( .A(n5751), .ZN(n5878) );
  NAND2_X1 U6227 ( .A1(n7372), .A2(n5740), .ZN(n6212) );
  NAND2_X1 U6228 ( .A1(n10503), .A2(n10331), .ZN(n5115) );
  INV_X1 U6229 ( .A(n9836), .ZN(n9598) );
  NAND2_X1 U6230 ( .A1(n6182), .A2(n6181), .ZN(n9836) );
  NAND3_X1 U6231 ( .A1(n8583), .A2(n8590), .A3(n8369), .ZN(n5116) );
  XNOR2_X1 U6232 ( .A(n9868), .B(n9373), .ZN(n9689) );
  NAND2_X1 U6233 ( .A1(n5583), .A2(n6727), .ZN(n6824) );
  NAND2_X1 U6234 ( .A1(n5441), .A2(n6643), .ZN(n5117) );
  OR2_X1 U6235 ( .A1(n5976), .A2(SI_13_), .ZN(n5118) );
  NAND2_X1 U6236 ( .A1(n10193), .A2(n10206), .ZN(n5119) );
  INV_X1 U6237 ( .A(n5507), .ZN(n5506) );
  OAI21_X1 U6238 ( .B1(n5509), .B2(n5508), .A(n9369), .ZN(n5507) );
  AND2_X1 U6239 ( .A1(n7277), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5120) );
  INV_X1 U6240 ( .A(n10414), .ZN(n5439) );
  INV_X1 U6241 ( .A(n9707), .ZN(n5357) );
  INV_X1 U6242 ( .A(n9520), .ZN(n9588) );
  NAND3_X1 U6243 ( .A1(n5622), .A2(n6681), .A3(n5503), .ZN(n5121) );
  AND2_X1 U6244 ( .A1(n5105), .A2(n9134), .ZN(n5122) );
  OR2_X1 U6245 ( .A1(n5096), .A2(n7323), .ZN(n5123) );
  OR2_X1 U6246 ( .A1(n7106), .A2(n5632), .ZN(n5124) );
  AND3_X1 U6247 ( .A1(n5722), .A2(n6285), .A3(n5535), .ZN(n5125) );
  NAND2_X1 U6248 ( .A1(n6792), .A2(n6793), .ZN(n5126) );
  AND2_X1 U6249 ( .A1(n5221), .A2(n5220), .ZN(n5127) );
  NOR2_X1 U6250 ( .A1(n8949), .A2(n7329), .ZN(n5128) );
  NOR2_X1 U6251 ( .A1(n8049), .A2(n5685), .ZN(n5684) );
  AND2_X1 U6252 ( .A1(n9528), .A2(n6420), .ZN(n5129) );
  NOR2_X1 U6253 ( .A1(n7951), .A2(n5442), .ZN(n5130) );
  INV_X1 U6254 ( .A(n5403), .ZN(n10219) );
  NOR2_X1 U6255 ( .A1(n10243), .A2(n10470), .ZN(n5403) );
  NAND2_X1 U6256 ( .A1(n6152), .A2(n6151), .ZN(n9846) );
  AND2_X1 U6257 ( .A1(n5409), .A2(n5413), .ZN(n5131) );
  NOR2_X1 U6258 ( .A1(n6246), .A2(n7376), .ZN(n5132) );
  INV_X1 U6259 ( .A(n6992), .ZN(n5615) );
  INV_X1 U6260 ( .A(n7922), .ZN(n5288) );
  NAND2_X1 U6261 ( .A1(n9642), .A2(n5338), .ZN(n5133) );
  OR2_X1 U6262 ( .A1(n10413), .A2(n10093), .ZN(n5134) );
  NAND2_X1 U6263 ( .A1(n6729), .A2(n6728), .ZN(n10625) );
  AND2_X1 U6264 ( .A1(n10306), .A2(n10283), .ZN(n5135) );
  NAND2_X1 U6265 ( .A1(n6854), .A2(n6853), .ZN(n8637) );
  AND2_X1 U6266 ( .A1(n9819), .A2(n9566), .ZN(n5136) );
  AND2_X1 U6267 ( .A1(n5966), .A2(n5945), .ZN(n5946) );
  AND2_X1 U6268 ( .A1(n10834), .A2(n8019), .ZN(n5137) );
  AND2_X1 U6269 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_DATAO_REG_4__SCAN_IN), 
        .ZN(n5138) );
  NOR2_X1 U6270 ( .A1(n10865), .A2(n8669), .ZN(n5139) );
  NOR2_X1 U6271 ( .A1(n6891), .A2(n8758), .ZN(n5140) );
  NOR2_X1 U6272 ( .A1(n5822), .A2(n7937), .ZN(n5141) );
  INV_X1 U6273 ( .A(n5658), .ZN(n5650) );
  NOR2_X1 U6274 ( .A1(n10013), .A2(n5142), .ZN(n5658) );
  AND2_X1 U6275 ( .A1(n5661), .A2(n5659), .ZN(n5142) );
  AND2_X1 U6276 ( .A1(n6512), .A2(n6511), .ZN(n5143) );
  AND2_X1 U6277 ( .A1(n6562), .A2(n6561), .ZN(n5144) );
  INV_X1 U6278 ( .A(n5549), .ZN(n6120) );
  OAI21_X1 U6279 ( .B1(n6068), .B2(n5553), .A(n5550), .ZN(n5549) );
  INV_X1 U6280 ( .A(n5619), .ZN(n5618) );
  OR2_X1 U6281 ( .A1(n6993), .A2(n5620), .ZN(n5619) );
  AOI21_X1 U6282 ( .B1(n5358), .B2(n6075), .A(n5098), .ZN(n5453) );
  NOR2_X1 U6283 ( .A1(n10470), .A2(n10091), .ZN(n5145) );
  NAND2_X1 U6284 ( .A1(n9856), .A2(n9364), .ZN(n5146) );
  NAND2_X1 U6285 ( .A1(n6648), .A2(n5621), .ZN(n5147) );
  INV_X1 U6286 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5531) );
  INV_X1 U6287 ( .A(n5393), .ZN(n5392) );
  NAND2_X1 U6288 ( .A1(n5104), .A2(n5394), .ZN(n5393) );
  OR2_X1 U6289 ( .A1(n7140), .A2(n5636), .ZN(n5148) );
  NAND2_X1 U6290 ( .A1(n5318), .A2(n5119), .ZN(n5149) );
  INV_X1 U6291 ( .A(n5259), .ZN(n5258) );
  NAND2_X1 U6292 ( .A1(n8114), .A2(n5260), .ZN(n5259) );
  AND2_X1 U6293 ( .A1(n5901), .A2(n8432), .ZN(n5150) );
  AND2_X1 U6294 ( .A1(n6519), .A2(n6520), .ZN(n5151) );
  AND2_X1 U6295 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5152) );
  INV_X1 U6296 ( .A(n6028), .ZN(n5532) );
  INV_X1 U6297 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5733) );
  INV_X1 U6298 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5283) );
  INV_X1 U6299 ( .A(n5461), .ZN(n5460) );
  NAND2_X1 U6300 ( .A1(n5463), .A2(n6358), .ZN(n5461) );
  NOR2_X1 U6301 ( .A1(n5633), .A2(n9939), .ZN(n5153) );
  OR2_X1 U6302 ( .A1(n5654), .A2(n5651), .ZN(n5154) );
  NAND2_X1 U6303 ( .A1(n5793), .A2(SI_4_), .ZN(n5811) );
  AND3_X1 U6304 ( .A1(n5244), .A2(n5253), .A3(n5243), .ZN(n5155) );
  NAND2_X1 U6305 ( .A1(n6414), .A2(n6413), .ZN(n9563) );
  AND2_X1 U6306 ( .A1(n5691), .A2(n8861), .ZN(n5156) );
  NAND2_X1 U6307 ( .A1(n5909), .A2(n5908), .ZN(n8811) );
  NAND2_X1 U6308 ( .A1(n5965), .A2(n6353), .ZN(n5157) );
  AND2_X1 U6309 ( .A1(n5565), .A2(n6023), .ZN(n5158) );
  AND2_X1 U6310 ( .A1(n9000), .A2(n5414), .ZN(n5159) );
  NOR2_X1 U6311 ( .A1(n9624), .A2(n9517), .ZN(n5160) );
  AND2_X1 U6312 ( .A1(n7937), .A2(n5284), .ZN(n5161) );
  AND2_X1 U6313 ( .A1(n5439), .A2(n9237), .ZN(n5162) );
  AOI21_X1 U6314 ( .B1(n9675), .B2(n5682), .A(n5114), .ZN(n9601) );
  AND2_X1 U6315 ( .A1(n5435), .A2(n5434), .ZN(n5163) );
  INV_X1 U6316 ( .A(n9405), .ZN(n7778) );
  NAND2_X1 U6317 ( .A1(n5212), .A2(n5759), .ZN(n9405) );
  AND2_X1 U6318 ( .A1(n5836), .A2(n5846), .ZN(n5164) );
  AND2_X1 U6319 ( .A1(n5376), .A2(n5372), .ZN(n5371) );
  INV_X1 U6320 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6643) );
  NAND2_X2 U6321 ( .A1(n9271), .A2(n6667), .ZN(n6761) );
  NAND2_X1 U6322 ( .A1(n6195), .A2(n6194), .ZN(n9830) );
  INV_X1 U6323 ( .A(n9830), .ZN(n5335) );
  AND2_X1 U6324 ( .A1(n5462), .A2(n5460), .ZN(n5165) );
  INV_X1 U6325 ( .A(n9051), .ZN(n5426) );
  OR2_X1 U6326 ( .A1(n6192), .A2(n5571), .ZN(n5166) );
  INV_X1 U6327 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5384) );
  NAND2_X1 U6328 ( .A1(n5587), .A2(n5590), .ZN(n8888) );
  OAI21_X1 U6329 ( .B1(n9212), .B2(n5489), .A(n5487), .ZN(n10382) );
  AND2_X1 U6330 ( .A1(n5335), .A2(n9565), .ZN(n5167) );
  OR2_X1 U6331 ( .A1(n9815), .A2(n10989), .ZN(n5168) );
  INV_X1 U6332 ( .A(n9293), .ZN(n5252) );
  NAND2_X1 U6333 ( .A1(n5607), .A2(n6950), .ZN(n10024) );
  AND4_X1 U6334 ( .A1(n6097), .A2(n6096), .A3(n6095), .A4(n6094), .ZN(n9373)
         );
  INV_X1 U6335 ( .A(n9373), .ZN(n5455) );
  NAND2_X1 U6336 ( .A1(n7142), .A2(n7141), .ZN(n10464) );
  INV_X1 U6337 ( .A(n10464), .ZN(n5402) );
  AND2_X1 U6338 ( .A1(n7467), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5169) );
  AND2_X1 U6339 ( .A1(n10486), .A2(n10284), .ZN(n5170) );
  AND2_X1 U6340 ( .A1(n9212), .A2(n9211), .ZN(n5171) );
  NAND2_X1 U6341 ( .A1(n10317), .A2(n5392), .ZN(n5395) );
  AND2_X1 U6342 ( .A1(n5527), .A2(n5525), .ZN(n5172) );
  AND2_X1 U6343 ( .A1(n10454), .A2(n10197), .ZN(n5173) );
  INV_X1 U6344 ( .A(n5326), .ZN(n5325) );
  AND2_X1 U6345 ( .A1(n5327), .A2(n9221), .ZN(n5326) );
  INV_X1 U6346 ( .A(n5457), .ZN(n9767) );
  OAI211_X1 U6347 ( .C1(n10921), .C2(n5461), .A(n5467), .B(n5458), .ZN(n5457)
         );
  OR2_X1 U6348 ( .A1(n6112), .A2(SI_20_), .ZN(n5174) );
  INV_X1 U6349 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5711) );
  XNOR2_X1 U6350 ( .A(n7137), .B(n7154), .ZN(n9968) );
  OR3_X1 U6351 ( .A1(n5968), .A2(n5532), .A3(n5530), .ZN(n5175) );
  INV_X1 U6352 ( .A(n5672), .ZN(n9887) );
  NAND2_X1 U6353 ( .A1(n5669), .A2(n5673), .ZN(n5672) );
  INV_X1 U6354 ( .A(n5557), .ZN(n5556) );
  NOR2_X1 U6355 ( .A1(n6100), .A2(n5558), .ZN(n5557) );
  AND2_X1 U6356 ( .A1(n6099), .A2(n8222), .ZN(n5176) );
  NOR2_X1 U6357 ( .A1(n6044), .A2(SI_16_), .ZN(n5177) );
  OR2_X1 U6358 ( .A1(n9733), .A2(n5347), .ZN(n5178) );
  OR2_X1 U6359 ( .A1(n10413), .A2(n10425), .ZN(n9060) );
  INV_X1 U6360 ( .A(n9216), .ZN(n5486) );
  NAND2_X1 U6361 ( .A1(n9292), .A2(n9291), .ZN(n5179) );
  AND2_X1 U6362 ( .A1(n10850), .A2(n8649), .ZN(n5180) );
  AND2_X1 U6363 ( .A1(n9507), .A2(n5689), .ZN(n5181) );
  INV_X1 U6364 ( .A(n10919), .ZN(n5468) );
  INV_X1 U6365 ( .A(n11020), .ZN(n5418) );
  NOR2_X1 U6366 ( .A1(n6286), .A2(n6622), .ZN(n5182) );
  INV_X1 U6367 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5217) );
  NAND3_X1 U6368 ( .A1(n5389), .A2(n8128), .A3(n10843), .ZN(n5183) );
  INV_X1 U6369 ( .A(n9337), .ZN(n5508) );
  OR2_X1 U6370 ( .A1(n6238), .A2(n5576), .ZN(n5184) );
  OR2_X1 U6371 ( .A1(n11020), .A2(n5421), .ZN(n5185) );
  OR2_X1 U6372 ( .A1(n11024), .A2(n8940), .ZN(n5186) );
  NAND2_X1 U6373 ( .A1(n6818), .A2(n8089), .ZN(n8098) );
  AOI21_X1 U6374 ( .B1(n5598), .B2(n6818), .A(n5599), .ZN(n8692) );
  NAND2_X1 U6375 ( .A1(n7078), .A2(n7077), .ZN(n10486) );
  INV_X1 U6376 ( .A(n10486), .ZN(n5394) );
  NAND2_X1 U6377 ( .A1(n6648), .A2(n5622), .ZN(n5187) );
  OR2_X1 U6378 ( .A1(n8683), .A2(n5343), .ZN(n5188) );
  AND2_X1 U6379 ( .A1(n10818), .A2(n8018), .ZN(n5189) );
  INV_X1 U6380 ( .A(n5517), .ZN(n5516) );
  NOR2_X1 U6381 ( .A1(n8161), .A2(n5518), .ZN(n5517) );
  INV_X1 U6382 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5216) );
  AND2_X1 U6383 ( .A1(n5443), .A2(n6320), .ZN(n5190) );
  AND2_X1 U6384 ( .A1(n6333), .A2(n8004), .ZN(n8049) );
  INV_X1 U6385 ( .A(n8049), .ZN(n5686) );
  OR2_X1 U6386 ( .A1(n10883), .A2(n9210), .ZN(n5191) );
  NOR2_X1 U6387 ( .A1(n8683), .A2(n5341), .ZN(n5340) );
  INV_X1 U6388 ( .A(n10071), .ZN(n10078) );
  NAND2_X1 U6389 ( .A1(n6647), .A2(n6664), .ZN(n7202) );
  NOR3_X1 U6390 ( .A1(n6652), .A2(n5117), .A3(P1_IR_REG_29__SCAN_IN), .ZN(
        n10533) );
  INV_X1 U6391 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5479) );
  NAND2_X1 U6392 ( .A1(n7605), .A2(n7350), .ZN(n5192) );
  AND2_X1 U6393 ( .A1(n7371), .A2(n7355), .ZN(n7605) );
  MUX2_X1 U6394 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n7272), .S(n10625), .Z(n10629) );
  NAND2_X1 U6395 ( .A1(n7675), .A2(n7674), .ZN(n7673) );
  INV_X1 U6396 ( .A(n5724), .ZN(n5726) );
  INV_X1 U6397 ( .A(n9911), .ZN(n5202) );
  OAI21_X1 U6398 ( .B1(n7952), .B2(n5288), .A(n5203), .ZN(n8015) );
  INV_X1 U6399 ( .A(n5204), .ZN(n5203) );
  OAI21_X1 U6400 ( .B1(n5288), .B2(n7951), .A(n8011), .ZN(n5204) );
  MUX2_X1 U6401 ( .A(n5725), .B(P2_REG2_REG_1__SCAN_IN), .S(n10648), .Z(n10645) );
  NAND2_X1 U6402 ( .A1(n6484), .A2(n7742), .ZN(n7820) );
  NAND2_X1 U6403 ( .A1(n6601), .A2(n5246), .ZN(n5245) );
  NAND2_X1 U6404 ( .A1(n6601), .A2(n6600), .ZN(n9294) );
  OAI211_X1 U6405 ( .C1(n6601), .C2(n5248), .A(n5245), .B(n5155), .ZN(n9308)
         );
  NAND3_X1 U6406 ( .A1(n9302), .A2(n5249), .A3(n5252), .ZN(n5243) );
  INV_X1 U6407 ( .A(n9302), .ZN(n5255) );
  NAND2_X2 U6408 ( .A1(n7372), .A2(n7320), .ZN(n6278) );
  OAI21_X1 U6409 ( .B1(n9328), .B2(n5507), .A(n5276), .ZN(n9285) );
  NAND2_X1 U6410 ( .A1(n5275), .A2(n5273), .ZN(n6567) );
  NAND2_X1 U6411 ( .A1(n9328), .A2(n5276), .ZN(n5275) );
  NAND2_X1 U6412 ( .A1(n6311), .A2(n5278), .ZN(n6312) );
  OAI21_X1 U6413 ( .B1(n5769), .B2(n5278), .A(n6315), .ZN(n7780) );
  XNOR2_X1 U6414 ( .A(n8143), .B(n5278), .ZN(n8151) );
  NAND2_X1 U6415 ( .A1(n5757), .A2(n6434), .ZN(n5278) );
  AND3_X1 U6416 ( .A1(n5473), .A2(n5534), .A3(n5535), .ZN(n6258) );
  NAND4_X1 U6417 ( .A1(n5280), .A2(n5722), .A3(n5535), .A4(n5279), .ZN(n5281)
         );
  NAND2_X1 U6418 ( .A1(n5285), .A2(n5161), .ZN(n6328) );
  NAND3_X1 U6419 ( .A1(n6323), .A2(n6322), .A3(n5286), .ZN(n5285) );
  NAND3_X1 U6420 ( .A1(n6423), .A2(n6421), .A3(n6422), .ZN(n5290) );
  NAND3_X1 U6421 ( .A1(n5292), .A2(n6416), .A3(n6415), .ZN(n5291) );
  NAND3_X1 U6422 ( .A1(n5294), .A2(n5293), .A3(n9554), .ZN(n5292) );
  NAND3_X1 U6423 ( .A1(n6332), .A2(n6331), .A3(n5298), .ZN(n5296) );
  NAND2_X1 U6424 ( .A1(n5296), .A2(n5295), .ZN(n6343) );
  NAND2_X1 U6425 ( .A1(n8021), .A2(n6334), .ZN(n5300) );
  INV_X1 U6426 ( .A(n5302), .ZN(n5301) );
  OAI22_X1 U6427 ( .A1(n6278), .A2(n7321), .B1(n7372), .B2(n7386), .ZN(n5302)
         );
  NAND2_X4 U6428 ( .A1(n5386), .A2(n5385), .ZN(n5740) );
  NAND2_X2 U6429 ( .A1(n5737), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U6430 ( .A1(n5315), .A2(n5316), .ZN(n9234) );
  NAND2_X1 U6431 ( .A1(n10189), .A2(n5317), .ZN(n5315) );
  OAI21_X1 U6432 ( .B1(n10311), .B2(n5322), .A(n5320), .ZN(n5492) );
  NAND3_X1 U6433 ( .A1(n5677), .A2(n5711), .A3(n5712), .ZN(n5675) );
  INV_X1 U6434 ( .A(n5340), .ZN(n8853) );
  OR2_X1 U6435 ( .A1(n9546), .A2(n9815), .ZN(n5350) );
  NAND3_X1 U6436 ( .A1(n5352), .A2(n5811), .A3(n5539), .ZN(n5351) );
  NAND3_X1 U6437 ( .A1(n6471), .A2(n5706), .A3(n5353), .ZN(n6475) );
  AOI21_X2 U6438 ( .B1(n6281), .B2(n6447), .A(n6287), .ZN(n6452) );
  NAND2_X1 U6439 ( .A1(n5837), .A2(n5164), .ZN(n5852) );
  NAND2_X1 U6440 ( .A1(n5867), .A2(n5100), .ZN(n5540) );
  OAI21_X2 U6441 ( .B1(n7843), .B2(n5096), .A(n6069), .ZN(n9871) );
  NAND2_X1 U6442 ( .A1(n9562), .A2(n5364), .ZN(n5361) );
  NAND2_X1 U6443 ( .A1(n5361), .A2(n5362), .ZN(n6266) );
  NAND3_X1 U6444 ( .A1(n5365), .A2(n5366), .A3(n6292), .ZN(n5363) );
  NAND2_X1 U6445 ( .A1(n5941), .A2(n5371), .ZN(n5369) );
  NAND2_X1 U6446 ( .A1(n5941), .A2(n5940), .ZN(n5947) );
  NAND3_X1 U6447 ( .A1(n5382), .A2(n5383), .A3(n5381), .ZN(n5793) );
  NAND3_X1 U6448 ( .A1(n5739), .A2(n5738), .A3(P1_DATAO_REG_4__SCAN_IN), .ZN(
        n5381) );
  NAND3_X1 U6449 ( .A1(n5386), .A2(P2_DATAO_REG_4__SCAN_IN), .A3(n5385), .ZN(
        n5382) );
  INV_X8 U6450 ( .A(n5740), .ZN(n7320) );
  NAND2_X1 U6451 ( .A1(n10317), .A2(n5391), .ZN(n10252) );
  INV_X1 U6452 ( .A(n5395), .ZN(n10270) );
  NAND2_X1 U6453 ( .A1(n5396), .A2(n5075), .ZN(n10392) );
  NAND2_X1 U6454 ( .A1(n6996), .A2(n5404), .ZN(n6677) );
  NAND2_X1 U6455 ( .A1(n7981), .A2(n9091), .ZN(n5407) );
  NAND2_X1 U6456 ( .A1(n5407), .A2(n5405), .ZN(n5408) );
  NOR2_X1 U6457 ( .A1(n10781), .A2(n5406), .ZN(n5405) );
  INV_X1 U6458 ( .A(n9096), .ZN(n5406) );
  NAND2_X2 U6459 ( .A1(n5408), .A2(n9098), .ZN(n8963) );
  NAND2_X1 U6460 ( .A1(n10366), .A2(n5159), .ZN(n5412) );
  NAND2_X1 U6461 ( .A1(n10259), .A2(n5431), .ZN(n5430) );
  OR2_X1 U6462 ( .A1(n10259), .A2(n9250), .ZN(n5435) );
  INV_X1 U6463 ( .A(n5435), .ZN(n10238) );
  NAND2_X1 U6464 ( .A1(n10418), .A2(n5162), .ZN(n5438) );
  NAND2_X1 U6465 ( .A1(n10418), .A2(n9237), .ZN(n10401) );
  NOR2_X1 U6466 ( .A1(n6652), .A2(n5440), .ZN(n6646) );
  NAND2_X1 U6467 ( .A1(n7868), .A2(n7867), .ZN(n9088) );
  NOR2_X4 U6468 ( .A1(n10777), .A2(n8105), .ZN(n8128) );
  AOI21_X2 U6469 ( .B1(n10367), .B2(n10363), .A(n10361), .ZN(n10366) );
  NAND2_X1 U6470 ( .A1(n10295), .A2(n9245), .ZN(n10280) );
  NAND2_X1 U6471 ( .A1(n10194), .A2(n9256), .ZN(n10172) );
  NAND2_X1 U6472 ( .A1(n10172), .A2(n10171), .ZN(n10170) );
  OR2_X1 U6473 ( .A1(n6761), .A2(n7243), .ZN(n6723) );
  NAND2_X1 U6474 ( .A1(n8963), .A2(n9102), .ZN(n8174) );
  AOI21_X2 U6475 ( .B1(n5446), .B2(n5445), .A(n5444), .ZN(n9648) );
  INV_X1 U6476 ( .A(n6353), .ZN(n5465) );
  NAND2_X1 U6477 ( .A1(n5460), .A2(n5459), .ZN(n5458) );
  INV_X1 U6478 ( .A(n5464), .ZN(n5459) );
  OAI211_X2 U6479 ( .C1(n8949), .C2(n5479), .A(n5478), .B(n5477), .ZN(n6736)
         );
  NAND2_X2 U6480 ( .A1(n7263), .A2(n7320), .ZN(n6746) );
  NAND2_X1 U6481 ( .A1(n5481), .A2(n5484), .ZN(n9219) );
  NAND2_X1 U6482 ( .A1(n9215), .A2(n5482), .ZN(n5481) );
  NAND2_X1 U6483 ( .A1(n5492), .A2(n5493), .ZN(n10251) );
  NAND2_X1 U6484 ( .A1(n9405), .A2(n9295), .ZN(n6480) );
  NAND3_X1 U6485 ( .A1(n5534), .A2(n5535), .A3(n5533), .ZN(n5953) );
  NAND2_X1 U6486 ( .A1(n5540), .A2(n5541), .ZN(n5920) );
  NAND2_X1 U6487 ( .A1(n5867), .A2(n5866), .ZN(n5872) );
  NAND2_X1 U6488 ( .A1(n10539), .A2(n5271), .ZN(n5561) );
  NAND2_X1 U6489 ( .A1(n5561), .A2(n6279), .ZN(n9805) );
  NAND2_X1 U6490 ( .A1(n5561), .A2(n5559), .ZN(n6280) );
  NAND2_X1 U6491 ( .A1(n5967), .A2(n5966), .ZN(n5978) );
  NAND2_X1 U6492 ( .A1(n6165), .A2(n5572), .ZN(n6180) );
  NAND2_X1 U6493 ( .A1(n6165), .A2(n6164), .ZN(n6168) );
  NAND2_X1 U6494 ( .A1(n6207), .A2(n5577), .ZN(n6222) );
  NAND2_X1 U6495 ( .A1(n6207), .A2(n6206), .ZN(n6210) );
  MUX2_X1 U6496 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n5740), .Z(n5579) );
  NAND3_X1 U6497 ( .A1(n5582), .A2(n5583), .A3(n6727), .ZN(n6972) );
  NAND3_X1 U6498 ( .A1(n10002), .A2(n10003), .A3(n10006), .ZN(n10004) );
  NAND2_X1 U6499 ( .A1(n7178), .A2(n9208), .ZN(n7198) );
  NAND2_X1 U6500 ( .A1(n7160), .A2(n5584), .ZN(n9208) );
  NAND2_X1 U6501 ( .A1(n7160), .A2(n7159), .ZN(n7177) );
  NAND2_X1 U6502 ( .A1(n5586), .A2(n5588), .ZN(n6934) );
  NAND2_X1 U6503 ( .A1(n6911), .A2(n5590), .ZN(n5586) );
  NAND2_X1 U6504 ( .A1(n6911), .A2(n6912), .ZN(n8875) );
  OR2_X1 U6505 ( .A1(n6911), .A2(n6912), .ZN(n8876) );
  INV_X1 U6506 ( .A(n8877), .ZN(n5592) );
  NAND3_X1 U6507 ( .A1(n6818), .A2(n8089), .A3(n5593), .ZN(n5597) );
  NOR2_X1 U6508 ( .A1(n8693), .A2(n5594), .ZN(n5593) );
  NAND2_X1 U6509 ( .A1(n5597), .A2(n5595), .ZN(n6851) );
  INV_X1 U6510 ( .A(n8693), .ZN(n5596) );
  INV_X1 U6511 ( .A(n8906), .ZN(n5608) );
  NAND3_X1 U6512 ( .A1(n6991), .A2(n5614), .A3(n5099), .ZN(n5610) );
  NAND3_X1 U6513 ( .A1(n6991), .A2(n5099), .A3(n5615), .ZN(n5611) );
  AND2_X1 U6514 ( .A1(n6648), .A2(n6641), .ZN(n6996) );
  INV_X1 U6515 ( .A(n5626), .ZN(n10063) );
  NAND2_X1 U6516 ( .A1(n7106), .A2(n7104), .ZN(n9938) );
  INV_X1 U6517 ( .A(n9744), .ZN(n5669) );
  NAND2_X1 U6518 ( .A1(n10990), .A2(n9508), .ZN(n5691) );
  NAND2_X1 U6519 ( .A1(n5925), .A2(n5924), .ZN(n5941) );
  AND2_X1 U6520 ( .A1(n10183), .A2(n10182), .ZN(n10455) );
  NOR2_X2 U6521 ( .A1(n7873), .A2(n10720), .ZN(n10740) );
  NAND2_X1 U6522 ( .A1(n10169), .A2(n10168), .ZN(n10458) );
  NAND2_X1 U6523 ( .A1(n6645), .A2(n6644), .ZN(n6647) );
  NAND2_X1 U6524 ( .A1(n7989), .A2(n10781), .ZN(n7991) );
  AOI22_X1 U6525 ( .A1(n6735), .A2(n9196), .B1(n6719), .B2(n6736), .ZN(n7640)
         );
  OAI21_X1 U6526 ( .B1(n10458), .B2(n10895), .A(n10177), .ZN(n10453) );
  OR2_X1 U6527 ( .A1(n8949), .A2(n7328), .ZN(n6749) );
  INV_X1 U6528 ( .A(n9939), .ZN(n9940) );
  NAND2_X1 U6529 ( .A1(n8121), .A2(n8120), .ZN(n8170) );
  AOI21_X1 U6530 ( .B1(n8170), .B2(n8169), .A(n8168), .ZN(n8171) );
  OR2_X1 U6531 ( .A1(n6736), .A2(n7699), .ZN(n7873) );
  INV_X1 U6532 ( .A(n6258), .ZN(n6259) );
  INV_X1 U6533 ( .A(n9271), .ZN(n6668) );
  XNOR2_X1 U6534 ( .A(n7642), .B(n10720), .ZN(n9127) );
  NOR2_X1 U6535 ( .A1(n9513), .A2(n9647), .ZN(n5696) );
  INV_X1 U6536 ( .A(n8650), .ZN(n5899) );
  AND2_X1 U6537 ( .A1(n9706), .A2(n9719), .ZN(n5698) );
  OR2_X1 U6538 ( .A1(n9561), .A2(n9335), .ZN(n5700) );
  OR2_X1 U6539 ( .A1(n7263), .A2(n7495), .ZN(n5702) );
  CLKBUF_X2 U6540 ( .A(P1_U4006), .Z(n10104) );
  OR2_X1 U6541 ( .A1(n7263), .A2(n10658), .ZN(n5703) );
  NOR2_X1 U6542 ( .A1(n6781), .A2(n7888), .ZN(n5705) );
  OR2_X1 U6543 ( .A1(n9878), .A2(n9709), .ZN(n5707) );
  NAND2_X1 U6544 ( .A1(n6280), .A2(n6421), .ZN(n6291) );
  INV_X1 U6545 ( .A(n8817), .ZN(n8814) );
  INV_X1 U6546 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5713) );
  AND2_X1 U6547 ( .A1(n9380), .A2(n9378), .ZN(n6596) );
  NAND2_X1 U6548 ( .A1(n6773), .A2(n6772), .ZN(n6774) );
  INV_X1 U6549 ( .A(n6756), .ZN(n6757) );
  INV_X1 U6550 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6641) );
  OR2_X1 U6551 ( .A1(n6105), .A2(n9356), .ZN(n6126) );
  OR2_X1 U6552 ( .A1(n5934), .A2(n8663), .ZN(n5959) );
  AND2_X1 U6553 ( .A1(n6431), .A2(n10920), .ZN(n8675) );
  INV_X1 U6554 ( .A(n8860), .ZN(n8815) );
  AND2_X1 U6555 ( .A1(n9408), .A2(n10680), .ZN(n10703) );
  AOI21_X1 U6556 ( .B1(n6797), .B2(n5126), .A(n6796), .ZN(n6814) );
  AND2_X1 U6557 ( .A1(n7032), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n7051) );
  NAND2_X1 U6558 ( .A1(n10449), .A2(n9016), .ZN(n9159) );
  NOR2_X1 U6559 ( .A1(n6977), .A2(n7973), .ZN(n6978) );
  INV_X1 U6560 ( .A(n7263), .ZN(n7028) );
  INV_X1 U6561 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8369) );
  NAND2_X1 U6562 ( .A1(n5848), .A2(SI_7_), .ZN(n5866) );
  NAND2_X1 U6563 ( .A1(n8775), .A2(n6531), .ZN(n8799) );
  OR2_X1 U6564 ( .A1(n6196), .A2(n8510), .ZN(n6227) );
  NAND2_X1 U6565 ( .A1(n8672), .A2(n8671), .ZN(n8813) );
  INV_X1 U6566 ( .A(n10939), .ZN(n10932) );
  AND2_X1 U6567 ( .A1(n7784), .A2(n7783), .ZN(n9717) );
  AND2_X1 U6568 ( .A1(n7606), .A2(n7605), .ZN(n7766) );
  INV_X1 U6569 ( .A(n10081), .ZN(n10066) );
  INV_X1 U6570 ( .A(n10459), .ZN(n10193) );
  AND2_X1 U6571 ( .A1(n9053), .A2(n9045), .ZN(n9134) );
  XNOR2_X1 U6572 ( .A(n5976), .B(SI_13_), .ZN(n5977) );
  XNOR2_X1 U6573 ( .A(n5917), .B(n8431), .ZN(n5919) );
  AND2_X1 U6574 ( .A1(n5791), .A2(n5781), .ZN(n5782) );
  AND2_X1 U6575 ( .A1(n6635), .A2(n6634), .ZN(n9384) );
  INV_X1 U6576 ( .A(n9335), .ZN(n9389) );
  AND2_X1 U6577 ( .A1(n6234), .A2(n6233), .ZN(n9566) );
  AND4_X1 U6578 ( .A1(n6111), .A2(n6110), .A3(n6109), .A4(n6108), .ZN(n9692)
         );
  AND4_X1 U6579 ( .A1(n5916), .A2(n5915), .A3(n5914), .A4(n5913), .ZN(n8664)
         );
  INV_X1 U6580 ( .A(n9563), .ZN(n9554) );
  INV_X1 U6581 ( .A(n9717), .ZN(n10929) );
  AND2_X1 U6582 ( .A1(n7767), .A2(n7766), .ZN(n7926) );
  AND2_X1 U6583 ( .A1(n5987), .A2(n6006), .ZN(n9410) );
  INV_X1 U6584 ( .A(n7218), .ZN(n9186) );
  AND2_X1 U6585 ( .A1(n7252), .A2(n7251), .ZN(n7561) );
  AND2_X1 U6586 ( .A1(n7670), .A2(n7203), .ZN(n10405) );
  AND2_X1 U6587 ( .A1(n5074), .A2(n7800), .ZN(n10902) );
  OR2_X1 U6588 ( .A1(n7799), .A2(n7218), .ZN(n11015) );
  OR2_X1 U6589 ( .A1(n9018), .A2(n9167), .ZN(n10737) );
  AND2_X1 U6590 ( .A1(n10621), .A2(n7652), .ZN(n7658) );
  INV_X1 U6591 ( .A(n9781), .ZN(n10990) );
  AND2_X1 U6592 ( .A1(n6625), .A2(n10700), .ZN(n9335) );
  AND4_X1 U6593 ( .A1(n6074), .A2(n6073), .A3(n6072), .A4(n6071), .ZN(n9719)
         );
  AOI21_X1 U6594 ( .B1(n9543), .B2(n10929), .A(n9542), .ZN(n9822) );
  NAND2_X1 U6595 ( .A1(n7956), .A2(n10700), .ZN(n10947) );
  INV_X1 U6596 ( .A(n10998), .ZN(n10997) );
  INV_X1 U6597 ( .A(n11002), .ZN(n10999) );
  AND2_X1 U6598 ( .A1(n6628), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7355) );
  INV_X1 U6599 ( .A(n7387), .ZN(n7437) );
  INV_X1 U6600 ( .A(n10086), .ZN(n10065) );
  AND2_X1 U6601 ( .A1(n7199), .A2(n10907), .ZN(n10089) );
  INV_X1 U6602 ( .A(n10432), .ZN(n10905) );
  INV_X1 U6603 ( .A(n11024), .ZN(n11021) );
  CLKBUF_X1 U6604 ( .A(n10583), .Z(n10571) );
  AND2_X1 U6605 ( .A1(n6475), .A2(n6474), .ZN(P2_U3244) );
  NOR2_X1 U6606 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5717) );
  NOR2_X1 U6607 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5716) );
  NOR2_X1 U6608 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5715) );
  NOR2_X1 U6609 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5714) );
  NAND4_X1 U6610 ( .A1(n5717), .A2(n5716), .A3(n5715), .A4(n5714), .ZN(n5720)
         );
  NAND4_X1 U6611 ( .A1(n5718), .A2(n5531), .A3(n6027), .A4(n6026), .ZN(n5719)
         );
  INV_X1 U6612 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5721) );
  INV_X1 U6613 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6285) );
  INV_X1 U6614 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5723) );
  INV_X1 U6615 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9912) );
  AND2_X2 U6616 ( .A1(n5726), .A2(n9918), .ZN(n5751) );
  NAND2_X1 U6617 ( .A1(n5751), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5731) );
  NAND2_X1 U6619 ( .A1(n6261), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5730) );
  INV_X1 U6620 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n5725) );
  OR2_X1 U6621 ( .A1(n6137), .A2(n5725), .ZN(n5729) );
  INV_X1 U6622 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10701) );
  INV_X1 U6623 ( .A(n5735), .ZN(n5736) );
  INV_X1 U6624 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n7321) );
  INV_X1 U6625 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6712) );
  INV_X1 U6626 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5741) );
  MUX2_X1 U6627 ( .A(n6712), .B(n5741), .S(n5740), .Z(n5742) );
  INV_X1 U6628 ( .A(SI_0_), .ZN(n6711) );
  NOR2_X2 U6629 ( .A1(n5742), .A2(n6711), .ZN(n5743) );
  NAND2_X1 U6630 ( .A1(n5743), .A2(SI_1_), .ZN(n5762) );
  INV_X1 U6631 ( .A(n5743), .ZN(n5744) );
  INV_X1 U6632 ( .A(SI_1_), .ZN(n8454) );
  NAND2_X1 U6633 ( .A1(n5744), .A2(n8454), .ZN(n5745) );
  MUX2_X1 U6634 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n7320), .Z(n5747) );
  INV_X1 U6635 ( .A(n5746), .ZN(n5749) );
  INV_X1 U6636 ( .A(n5747), .ZN(n5748) );
  NAND2_X1 U6637 ( .A1(n5749), .A2(n5748), .ZN(n5750) );
  NAND2_X1 U6638 ( .A1(n5763), .A2(n5750), .ZN(n7323) );
  NAND2_X1 U6639 ( .A1(n8148), .A2(n7771), .ZN(n6433) );
  NAND2_X1 U6640 ( .A1(n6261), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5755) );
  NAND2_X1 U6641 ( .A1(n5751), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5754) );
  NAND2_X1 U6642 ( .A1(n6248), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U6643 ( .A1(n6262), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5752) );
  NAND4_X1 U6644 ( .A1(n5755), .A2(n5754), .A3(n5753), .A4(n5752), .ZN(n9408)
         );
  NAND2_X1 U6645 ( .A1(n5740), .A2(SI_0_), .ZN(n5756) );
  XNOR2_X1 U6646 ( .A(n5756), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9926) );
  MUX2_X1 U6647 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9926), .S(n7372), .Z(n10680)
         );
  INV_X1 U6648 ( .A(n10680), .ZN(n10699) );
  OR2_X1 U6649 ( .A1(n9408), .A2(n10699), .ZN(n10695) );
  NAND2_X1 U6650 ( .A1(n6433), .A2(n10695), .ZN(n5757) );
  NAND2_X1 U6651 ( .A1(n9407), .A2(n10711), .ZN(n6434) );
  NAND2_X1 U6652 ( .A1(n5751), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5760) );
  INV_X1 U6653 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7376) );
  INV_X1 U6654 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n8154) );
  OR2_X1 U6655 ( .A1(n6175), .A2(n8154), .ZN(n5759) );
  INV_X1 U6656 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5758) );
  OR2_X1 U6657 ( .A1(n5735), .A2(n5723), .ZN(n5761) );
  XNOR2_X1 U6658 ( .A(n5761), .B(P2_IR_REG_2__SCAN_IN), .ZN(n7387) );
  INV_X1 U6659 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n7322) );
  INV_X1 U6660 ( .A(n5767), .ZN(n5764) );
  NAND2_X1 U6661 ( .A1(n5764), .A2(n5765), .ZN(n5768) );
  INV_X1 U6662 ( .A(n5765), .ZN(n5766) );
  NAND2_X1 U6663 ( .A1(n5768), .A2(n5778), .ZN(n7327) );
  NAND2_X1 U6664 ( .A1(n9405), .A2(n10730), .ZN(n6314) );
  INV_X1 U6665 ( .A(n6314), .ZN(n5769) );
  NAND2_X1 U6666 ( .A1(n7778), .A2(n8157), .ZN(n6315) );
  NAND2_X1 U6667 ( .A1(n5751), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5774) );
  INV_X1 U6668 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7375) );
  OR2_X1 U6669 ( .A1(n6175), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5772) );
  INV_X1 U6670 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5770) );
  OR2_X1 U6671 ( .A1(n6137), .A2(n5770), .ZN(n5771) );
  NAND2_X1 U6672 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5775), .ZN(n5776) );
  XNOR2_X1 U6673 ( .A(n5776), .B(P2_IR_REG_3__SCAN_IN), .ZN(n7389) );
  INV_X1 U6674 ( .A(n7389), .ZN(n7414) );
  INV_X1 U6675 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7324) );
  OR2_X1 U6676 ( .A1(n6278), .A2(n7324), .ZN(n5786) );
  MUX2_X1 U6677 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n7320), .Z(n5779) );
  INV_X1 U6678 ( .A(n5779), .ZN(n5780) );
  INV_X1 U6679 ( .A(SI_3_), .ZN(n8444) );
  NAND2_X1 U6680 ( .A1(n5780), .A2(n8444), .ZN(n5781) );
  NAND2_X2 U6681 ( .A1(n5783), .A2(n5782), .ZN(n5792) );
  OR2_X1 U6682 ( .A1(n5783), .A2(n5782), .ZN(n5784) );
  NAND2_X1 U6683 ( .A1(n5792), .A2(n5784), .ZN(n7325) );
  OR2_X1 U6684 ( .A1(n5096), .A2(n7325), .ZN(n5785) );
  OAI211_X1 U6685 ( .C1(n7372), .C2(n7414), .A(n5786), .B(n5785), .ZN(n7790)
         );
  INV_X1 U6686 ( .A(n7790), .ZN(n8743) );
  NAND2_X1 U6687 ( .A1(n9404), .A2(n8743), .ZN(n6321) );
  NAND2_X1 U6688 ( .A1(n8147), .A2(n7790), .ZN(n6320) );
  NAND2_X1 U6689 ( .A1(n5751), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U6690 ( .A1(n6262), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U6691 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5805) );
  OAI21_X1 U6692 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5805), .ZN(n7953) );
  OR2_X1 U6693 ( .A1(n6175), .A2(n7953), .ZN(n5788) );
  INV_X1 U6694 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7378) );
  OR2_X1 U6695 ( .A1(n6246), .A2(n7378), .ZN(n5787) );
  NAND4_X1 U6696 ( .A1(n5790), .A2(n5789), .A3(n5788), .A4(n5787), .ZN(n9403)
         );
  OR2_X1 U6697 ( .A1(n6278), .A2(n5384), .ZN(n5803) );
  INV_X1 U6698 ( .A(n5793), .ZN(n5794) );
  INV_X1 U6699 ( .A(SI_4_), .ZN(n8445) );
  NAND2_X1 U6700 ( .A1(n5794), .A2(n8445), .ZN(n5795) );
  OR2_X1 U6701 ( .A1(n5096), .A2(n7330), .ZN(n5802) );
  NAND2_X1 U6702 ( .A1(n5798), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5799) );
  MUX2_X1 U6703 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5799), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5800) );
  AND2_X1 U6704 ( .A1(n5800), .A2(n5111), .ZN(n7467) );
  NAND2_X1 U6705 ( .A1(n6085), .A2(n7467), .ZN(n5801) );
  XNOR2_X1 U6706 ( .A(n9403), .B(n10768), .ZN(n7951) );
  NAND2_X1 U6707 ( .A1(n9403), .A2(n10768), .ZN(n7939) );
  INV_X1 U6708 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7374) );
  OR2_X1 U6709 ( .A1(n6246), .A2(n7374), .ZN(n5810) );
  NAND2_X1 U6710 ( .A1(n5751), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5809) );
  INV_X1 U6711 ( .A(n5805), .ZN(n5804) );
  NAND2_X1 U6712 ( .A1(n5804), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5858) );
  INV_X1 U6713 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8488) );
  NAND2_X1 U6714 ( .A1(n5805), .A2(n8488), .ZN(n5806) );
  NAND2_X1 U6715 ( .A1(n5858), .A2(n5806), .ZN(n7928) );
  OR2_X1 U6716 ( .A1(n6175), .A2(n7928), .ZN(n5808) );
  INV_X1 U6717 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7929) );
  OR2_X1 U6718 ( .A1(n6137), .A2(n7929), .ZN(n5807) );
  MUX2_X1 U6719 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n7320), .Z(n5812) );
  INV_X1 U6720 ( .A(n5812), .ZN(n5814) );
  INV_X1 U6721 ( .A(SI_5_), .ZN(n5813) );
  NAND2_X1 U6722 ( .A1(n5814), .A2(n5813), .ZN(n5815) );
  NAND2_X1 U6723 ( .A1(n5834), .A2(n5704), .ZN(n5839) );
  OR2_X1 U6724 ( .A1(n5834), .A2(n5704), .ZN(n5816) );
  NAND2_X1 U6725 ( .A1(n5839), .A2(n5816), .ZN(n7333) );
  OR2_X1 U6726 ( .A1(n5096), .A2(n7333), .ZN(n5820) );
  INV_X1 U6727 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7331) );
  OR2_X1 U6728 ( .A1(n6278), .A2(n7331), .ZN(n5819) );
  NAND2_X1 U6729 ( .A1(n5111), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5817) );
  XNOR2_X1 U6730 ( .A(n5817), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7391) );
  NAND2_X1 U6731 ( .A1(n6085), .A2(n7391), .ZN(n5818) );
  NAND2_X1 U6732 ( .A1(n9789), .A2(n10802), .ZN(n5821) );
  AND2_X1 U6733 ( .A1(n7939), .A2(n5821), .ZN(n5823) );
  INV_X1 U6734 ( .A(n5821), .ZN(n5822) );
  XNOR2_X1 U6735 ( .A(n9789), .B(n10802), .ZN(n8011) );
  INV_X1 U6736 ( .A(n8011), .ZN(n7937) );
  NAND2_X1 U6737 ( .A1(n6261), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5827) );
  NAND2_X1 U6738 ( .A1(n5751), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5826) );
  INV_X1 U6739 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8506) );
  XNOR2_X1 U6740 ( .A(n5858), .B(n8506), .ZN(n9794) );
  OR2_X1 U6741 ( .A1(n6175), .A2(n9794), .ZN(n5825) );
  INV_X1 U6742 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n9790) );
  OR2_X1 U6743 ( .A1(n6137), .A2(n9790), .ZN(n5824) );
  NAND4_X1 U6744 ( .A1(n5827), .A2(n5826), .A3(n5825), .A4(n5824), .ZN(n9402)
         );
  INV_X1 U6745 ( .A(n9402), .ZN(n8048) );
  OR2_X1 U6746 ( .A1(n5828), .A2(n5723), .ZN(n5829) );
  XNOR2_X1 U6747 ( .A(n5829), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7451) );
  AOI22_X1 U6748 ( .A1(n6086), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6085), .B2(
        n7451), .ZN(n5844) );
  MUX2_X1 U6749 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7320), .Z(n5830) );
  INV_X1 U6750 ( .A(n5830), .ZN(n5831) );
  NAND2_X1 U6751 ( .A1(n5831), .A2(n8443), .ZN(n5832) );
  INV_X1 U6752 ( .A(n5840), .ZN(n5835) );
  NAND2_X1 U6753 ( .A1(n5839), .A2(n5838), .ZN(n5841) );
  OR2_X1 U6754 ( .A1(n5841), .A2(n5840), .ZN(n5842) );
  NAND2_X1 U6755 ( .A1(n5847), .A2(n5842), .ZN(n7335) );
  OR2_X1 U6756 ( .A1(n7335), .A2(n5096), .ZN(n5843) );
  NAND2_X1 U6757 ( .A1(n5844), .A2(n5843), .ZN(n9796) );
  NAND2_X1 U6758 ( .A1(n8048), .A2(n9796), .ZN(n5845) );
  INV_X1 U6759 ( .A(n9796), .ZN(n10819) );
  NAND2_X1 U6760 ( .A1(n9402), .A2(n10819), .ZN(n8044) );
  MUX2_X1 U6761 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7320), .Z(n5848) );
  INV_X1 U6762 ( .A(n5848), .ZN(n5849) );
  INV_X1 U6763 ( .A(SI_7_), .ZN(n8234) );
  NAND2_X1 U6764 ( .A1(n5849), .A2(n8234), .ZN(n5850) );
  OR2_X1 U6765 ( .A1(n5852), .A2(n5851), .ZN(n5853) );
  NAND2_X1 U6766 ( .A1(n5867), .A2(n5853), .ZN(n7339) );
  OR2_X1 U6767 ( .A1(n7339), .A2(n5096), .ZN(n5857) );
  OR2_X1 U6768 ( .A1(n5854), .A2(n5723), .ZN(n5855) );
  XNOR2_X1 U6769 ( .A(n5855), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7514) );
  AOI22_X1 U6770 ( .A1(n6086), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6085), .B2(
        n7514), .ZN(n5856) );
  NAND2_X1 U6771 ( .A1(n6261), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5865) );
  NAND2_X1 U6772 ( .A1(n5751), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5864) );
  INV_X1 U6773 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8459) );
  OAI21_X1 U6774 ( .B1(n5858), .B2(n8506), .A(n8459), .ZN(n5861) );
  INV_X1 U6775 ( .A(n5858), .ZN(n5860) );
  AND2_X1 U6776 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n5859) );
  NAND2_X1 U6777 ( .A1(n5860), .A2(n5859), .ZN(n5881) );
  NAND2_X1 U6778 ( .A1(n5861), .A2(n5881), .ZN(n8052) );
  OR2_X1 U6779 ( .A1(n6175), .A2(n8052), .ZN(n5863) );
  INV_X1 U6780 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n8053) );
  OR2_X1 U6781 ( .A1(n6137), .A2(n8053), .ZN(n5862) );
  NAND4_X1 U6782 ( .A1(n5865), .A2(n5864), .A3(n5863), .A4(n5862), .ZN(n9788)
         );
  NAND2_X1 U6783 ( .A1(n10834), .A2(n9788), .ZN(n6333) );
  AND2_X1 U6784 ( .A1(n8044), .A2(n6333), .ZN(n8003) );
  MUX2_X1 U6785 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n7320), .Z(n5868) );
  INV_X1 U6786 ( .A(n5868), .ZN(n5869) );
  INV_X1 U6787 ( .A(SI_8_), .ZN(n8436) );
  NAND2_X1 U6788 ( .A1(n5869), .A2(n8436), .ZN(n5870) );
  OR2_X1 U6789 ( .A1(n5872), .A2(n5871), .ZN(n5873) );
  NAND2_X1 U6790 ( .A1(n5889), .A2(n5873), .ZN(n7348) );
  OR2_X1 U6791 ( .A1(n7348), .A2(n5096), .ZN(n5877) );
  NAND2_X1 U6792 ( .A1(n5874), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5875) );
  XNOR2_X1 U6793 ( .A(n5875), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7588) );
  AOI22_X1 U6794 ( .A1(n6086), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6085), .B2(
        n7588), .ZN(n5876) );
  NAND2_X1 U6795 ( .A1(n6261), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5886) );
  INV_X1 U6796 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5879) );
  OR2_X1 U6797 ( .A1(n5878), .A2(n5879), .ZN(n5885) );
  INV_X1 U6798 ( .A(n5881), .ZN(n5880) );
  NAND2_X1 U6799 ( .A1(n5880), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5893) );
  INV_X1 U6800 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8474) );
  NAND2_X1 U6801 ( .A1(n5881), .A2(n8474), .ZN(n5882) );
  NAND2_X1 U6802 ( .A1(n5893), .A2(n5882), .ZN(n8113) );
  OR2_X1 U6803 ( .A1(n6175), .A2(n8113), .ZN(n5884) );
  INV_X1 U6804 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n8023) );
  OR2_X1 U6805 ( .A1(n6137), .A2(n8023), .ZN(n5883) );
  OR2_X1 U6806 ( .A1(n10852), .A2(n8648), .ZN(n6335) );
  NAND2_X1 U6807 ( .A1(n10852), .A2(n8648), .ZN(n6336) );
  AND2_X1 U6808 ( .A1(n8003), .A2(n8021), .ZN(n5887) );
  INV_X1 U6809 ( .A(n9788), .ZN(n8019) );
  INV_X1 U6810 ( .A(n10834), .ZN(n8055) );
  NAND2_X1 U6811 ( .A1(n8019), .A2(n8055), .ZN(n8004) );
  MUX2_X1 U6812 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n7320), .Z(n5900) );
  XNOR2_X1 U6813 ( .A(n5903), .B(n5902), .ZN(n7357) );
  NAND2_X1 U6814 ( .A1(n7357), .A2(n5271), .ZN(n5891) );
  NAND2_X1 U6815 ( .A1(n5953), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5904) );
  XNOR2_X1 U6816 ( .A(n5904), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7709) );
  AOI22_X1 U6817 ( .A1(n6086), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6085), .B2(
        n7709), .ZN(n5890) );
  NAND2_X1 U6818 ( .A1(n6261), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5898) );
  INV_X1 U6819 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5892) );
  OR2_X1 U6820 ( .A1(n5878), .A2(n5892), .ZN(n5897) );
  INV_X1 U6821 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8493) );
  NAND2_X1 U6822 ( .A1(n5893), .A2(n8493), .ZN(n5894) );
  NAND2_X1 U6823 ( .A1(n5911), .A2(n5894), .ZN(n8654) );
  OR2_X1 U6824 ( .A1(n6175), .A2(n8654), .ZN(n5896) );
  INV_X1 U6825 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n8655) );
  OR2_X1 U6826 ( .A1(n6137), .A2(n8655), .ZN(n5895) );
  NAND2_X1 U6827 ( .A1(n10865), .A2(n8677), .ZN(n6345) );
  NAND2_X1 U6828 ( .A1(n6338), .A2(n6345), .ZN(n8650) );
  NAND2_X1 U6829 ( .A1(n8651), .A2(n6338), .ZN(n8676) );
  INV_X1 U6830 ( .A(n5900), .ZN(n5901) );
  INV_X1 U6831 ( .A(SI_9_), .ZN(n8432) );
  MUX2_X1 U6832 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n7320), .Z(n5917) );
  INV_X1 U6833 ( .A(SI_10_), .ZN(n8431) );
  XNOR2_X1 U6834 ( .A(n5920), .B(n5919), .ZN(n7398) );
  NAND2_X1 U6835 ( .A1(n7398), .A2(n5271), .ZN(n5909) );
  INV_X1 U6836 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5951) );
  NAND2_X1 U6837 ( .A1(n5904), .A2(n5951), .ZN(n5905) );
  NAND2_X1 U6838 ( .A1(n5905), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5906) );
  INV_X1 U6839 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5950) );
  NAND2_X1 U6840 ( .A1(n5906), .A2(n5950), .ZN(n5929) );
  OR2_X1 U6841 ( .A1(n5906), .A2(n5950), .ZN(n5907) );
  AOI22_X1 U6842 ( .A1(n6086), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6085), .B2(
        n7824), .ZN(n5908) );
  NAND2_X1 U6843 ( .A1(n5751), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5916) );
  INV_X1 U6844 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7716) );
  OR2_X1 U6845 ( .A1(n6246), .A2(n7716), .ZN(n5915) );
  INV_X1 U6846 ( .A(n5911), .ZN(n5910) );
  NAND2_X1 U6847 ( .A1(n5910), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5934) );
  INV_X1 U6848 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8463) );
  NAND2_X1 U6849 ( .A1(n5911), .A2(n8463), .ZN(n5912) );
  NAND2_X1 U6850 ( .A1(n5934), .A2(n5912), .ZN(n8686) );
  OR2_X1 U6851 ( .A1(n6175), .A2(n8686), .ZN(n5914) );
  INV_X1 U6852 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8687) );
  OR2_X1 U6853 ( .A1(n6137), .A2(n8687), .ZN(n5913) );
  INV_X1 U6854 ( .A(n6431), .ZN(n6341) );
  NAND2_X1 U6855 ( .A1(n8811), .A2(n8664), .ZN(n10920) );
  MUX2_X1 U6856 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n7320), .Z(n5921) );
  INV_X1 U6857 ( .A(n5921), .ZN(n5922) );
  INV_X1 U6858 ( .A(SI_11_), .ZN(n8238) );
  NAND2_X1 U6859 ( .A1(n5922), .A2(n8238), .ZN(n5923) );
  INV_X1 U6860 ( .A(n5925), .ZN(n5927) );
  NAND2_X1 U6861 ( .A1(n5927), .A2(n5926), .ZN(n5928) );
  NAND2_X1 U6862 ( .A1(n5941), .A2(n5928), .ZN(n7401) );
  OR2_X1 U6863 ( .A1(n7401), .A2(n5096), .ZN(n5932) );
  NAND2_X1 U6864 ( .A1(n5929), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5930) );
  XNOR2_X1 U6865 ( .A(n5930), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8038) );
  AOI22_X1 U6866 ( .A1(n6086), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6085), .B2(
        n8038), .ZN(n5931) );
  NAND2_X1 U6867 ( .A1(n5751), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5939) );
  INV_X1 U6868 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5933) );
  OR2_X1 U6869 ( .A1(n6137), .A2(n5933), .ZN(n5938) );
  INV_X1 U6870 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8663) );
  NAND2_X1 U6871 ( .A1(n5934), .A2(n8663), .ZN(n5935) );
  NAND2_X1 U6872 ( .A1(n5959), .A2(n5935), .ZN(n10936) );
  OR2_X1 U6873 ( .A1(n6175), .A2(n10936), .ZN(n5937) );
  INV_X1 U6874 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7829) );
  OR2_X1 U6875 ( .A1(n6246), .A2(n7829), .ZN(n5936) );
  OR2_X1 U6876 ( .A1(n10939), .A2(n9399), .ZN(n6352) );
  NAND2_X1 U6877 ( .A1(n10939), .A2(n9399), .ZN(n8807) );
  NAND2_X1 U6878 ( .A1(n6352), .A2(n8807), .ZN(n10919) );
  MUX2_X1 U6879 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n7320), .Z(n5942) );
  INV_X1 U6880 ( .A(n5942), .ZN(n5944) );
  INV_X1 U6881 ( .A(SI_12_), .ZN(n5943) );
  NAND2_X1 U6882 ( .A1(n5944), .A2(n5943), .ZN(n5945) );
  OR2_X1 U6883 ( .A1(n5947), .A2(n5946), .ZN(n5948) );
  NAND2_X1 U6884 ( .A1(n5967), .A2(n5948), .ZN(n7470) );
  OR2_X1 U6885 ( .A1(n7470), .A2(n5096), .ZN(n5956) );
  INV_X1 U6886 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5949) );
  NAND3_X1 U6887 ( .A1(n5951), .A2(n5950), .A3(n5949), .ZN(n5952) );
  NAND2_X1 U6888 ( .A1(n5968), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5954) );
  XNOR2_X1 U6889 ( .A(n5954), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8072) );
  AOI22_X1 U6890 ( .A1(n6086), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6085), .B2(
        n8072), .ZN(n5955) );
  NAND2_X1 U6891 ( .A1(n6261), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5964) );
  INV_X1 U6892 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n5957) );
  OR2_X1 U6893 ( .A1(n5878), .A2(n5957), .ZN(n5963) );
  INV_X1 U6894 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8481) );
  NAND2_X1 U6895 ( .A1(n5959), .A2(n8481), .ZN(n5960) );
  NAND2_X1 U6896 ( .A1(n5992), .A2(n5960), .ZN(n8820) );
  OR2_X1 U6897 ( .A1(n6175), .A2(n8820), .ZN(n5962) );
  INV_X1 U6898 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8821) );
  OR2_X1 U6899 ( .A1(n6137), .A2(n8821), .ZN(n5961) );
  NAND2_X1 U6900 ( .A1(n8858), .A2(n9398), .ZN(n6354) );
  NAND2_X1 U6901 ( .A1(n6354), .A2(n8807), .ZN(n5965) );
  MUX2_X1 U6902 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n7320), .Z(n5976) );
  XNOR2_X1 U6903 ( .A(n5978), .B(n5977), .ZN(n7558) );
  NAND2_X1 U6904 ( .A1(n7558), .A2(n5271), .ZN(n5970) );
  OR2_X1 U6905 ( .A1(n6029), .A2(n5723), .ZN(n5983) );
  XNOR2_X1 U6906 ( .A(n5983), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8192) );
  AOI22_X1 U6907 ( .A1(n6086), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6085), .B2(
        n8192), .ZN(n5969) );
  NAND2_X1 U6908 ( .A1(n5751), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5975) );
  INV_X1 U6909 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5971) );
  OR2_X1 U6910 ( .A1(n6246), .A2(n5971), .ZN(n5974) );
  INV_X1 U6911 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8288) );
  XNOR2_X1 U6912 ( .A(n5992), .B(n8288), .ZN(n8851) );
  OR2_X1 U6913 ( .A1(n6175), .A2(n8851), .ZN(n5973) );
  INV_X1 U6914 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8852) );
  OR2_X1 U6915 ( .A1(n6137), .A2(n8852), .ZN(n5972) );
  OR2_X1 U6916 ( .A1(n8857), .A2(n9775), .ZN(n6360) );
  NAND2_X1 U6917 ( .A1(n8857), .A2(n9775), .ZN(n6361) );
  NAND2_X1 U6918 ( .A1(n6360), .A2(n6361), .ZN(n8861) );
  INV_X1 U6919 ( .A(n6361), .ZN(n9769) );
  MUX2_X1 U6920 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n7320), .Z(n5979) );
  NAND2_X1 U6921 ( .A1(n5979), .A2(SI_14_), .ZN(n6021) );
  OAI21_X1 U6922 ( .B1(n5979), .B2(SI_14_), .A(n6021), .ZN(n5980) );
  NAND2_X1 U6923 ( .A1(n5981), .A2(n5980), .ZN(n5982) );
  NAND2_X1 U6924 ( .A1(n5982), .A2(n6024), .ZN(n7576) );
  OR2_X1 U6925 ( .A1(n7576), .A2(n5096), .ZN(n5989) );
  NAND2_X1 U6926 ( .A1(n5983), .A2(n6027), .ZN(n5984) );
  NAND2_X1 U6927 ( .A1(n5984), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5986) );
  INV_X1 U6928 ( .A(n5986), .ZN(n5985) );
  NAND2_X1 U6929 ( .A1(n5985), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U6930 ( .A1(n5986), .A2(n6026), .ZN(n6006) );
  AOI22_X1 U6931 ( .A1(n6086), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6085), .B2(
        n9410), .ZN(n5988) );
  NAND2_X1 U6932 ( .A1(n5751), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5998) );
  INV_X1 U6933 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5990) );
  OR2_X1 U6934 ( .A1(n6137), .A2(n5990), .ZN(n5997) );
  INV_X1 U6935 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5991) );
  OAI21_X1 U6936 ( .B1(n5992), .B2(n8288), .A(n5991), .ZN(n5993) );
  NAND2_X1 U6937 ( .A1(n5993), .A2(n6013), .ZN(n9777) );
  OR2_X1 U6938 ( .A1(n6175), .A2(n9777), .ZN(n5996) );
  INV_X1 U6939 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n5994) );
  OR2_X1 U6940 ( .A1(n6246), .A2(n5994), .ZN(n5995) );
  NAND2_X1 U6941 ( .A1(n9781), .A2(n9508), .ZN(n6365) );
  INV_X1 U6942 ( .A(n9766), .ZN(n9768) );
  INV_X1 U6943 ( .A(n6364), .ZN(n5999) );
  NOR2_X2 U6944 ( .A1(n9767), .A2(n5999), .ZN(n9757) );
  NAND2_X1 U6945 ( .A1(n6024), .A2(n6021), .ZN(n6003) );
  MUX2_X1 U6946 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n7320), .Z(n6000) );
  NAND2_X1 U6947 ( .A1(n6000), .A2(SI_15_), .ZN(n6020) );
  INV_X1 U6948 ( .A(n6000), .ZN(n6001) );
  INV_X1 U6949 ( .A(SI_15_), .ZN(n8226) );
  NAND2_X1 U6950 ( .A1(n6001), .A2(n8226), .ZN(n6022) );
  AND2_X1 U6951 ( .A1(n6020), .A2(n6022), .ZN(n6002) );
  NAND2_X1 U6952 ( .A1(n6003), .A2(n6002), .ZN(n6005) );
  NAND2_X1 U6953 ( .A1(n6006), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6007) );
  XNOR2_X1 U6954 ( .A(n6007), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9423) );
  AOI22_X1 U6955 ( .A1(n6086), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6085), .B2(
        n9423), .ZN(n6008) );
  NAND2_X1 U6956 ( .A1(n5751), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6019) );
  INV_X1 U6957 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n6010) );
  OR2_X1 U6958 ( .A1(n6246), .A2(n6010), .ZN(n6018) );
  INV_X1 U6959 ( .A(n6013), .ZN(n6011) );
  NAND2_X1 U6960 ( .A1(n6011), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6034) );
  INV_X1 U6961 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6012) );
  NAND2_X1 U6962 ( .A1(n6013), .A2(n6012), .ZN(n6014) );
  NAND2_X1 U6963 ( .A1(n6034), .A2(n6014), .ZN(n9752) );
  OR2_X1 U6964 ( .A1(n6175), .A2(n9752), .ZN(n6017) );
  INV_X1 U6965 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n6015) );
  OR2_X1 U6966 ( .A1(n6137), .A2(n6015), .ZN(n6016) );
  MUX2_X1 U6967 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n7320), .Z(n6044) );
  XNOR2_X1 U6968 ( .A(n6044), .B(SI_16_), .ZN(n6045) );
  XNOR2_X1 U6969 ( .A(n6046), .B(n6045), .ZN(n7662) );
  NAND2_X1 U6970 ( .A1(n7662), .A2(n5271), .ZN(n6032) );
  INV_X1 U6971 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6025) );
  AND3_X1 U6972 ( .A1(n6027), .A2(n6026), .A3(n6025), .ZN(n6028) );
  OR2_X1 U6973 ( .A1(n6052), .A2(n5723), .ZN(n6030) );
  XNOR2_X1 U6974 ( .A(n6030), .B(P2_IR_REG_16__SCAN_IN), .ZN(n9442) );
  AOI22_X1 U6975 ( .A1(n6086), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6085), .B2(
        n9442), .ZN(n6031) );
  NAND2_X1 U6976 ( .A1(n5751), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6039) );
  INV_X1 U6977 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9447) );
  OR2_X1 U6978 ( .A1(n6246), .A2(n9447), .ZN(n6038) );
  INV_X1 U6979 ( .A(n6034), .ZN(n6033) );
  NAND2_X1 U6980 ( .A1(n6033), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6056) );
  INV_X1 U6981 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8482) );
  NAND2_X1 U6982 ( .A1(n6034), .A2(n8482), .ZN(n6035) );
  NAND2_X1 U6983 ( .A1(n6056), .A2(n6035), .ZN(n9735) );
  OR2_X1 U6984 ( .A1(n6175), .A2(n9735), .ZN(n6037) );
  INV_X1 U6985 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9432) );
  OR2_X1 U6986 ( .A1(n6137), .A2(n9432), .ZN(n6036) );
  NAND2_X1 U6987 ( .A1(n9883), .A2(n9718), .ZN(n6308) );
  INV_X1 U6988 ( .A(n6308), .ZN(n6041) );
  NAND2_X1 U6989 ( .A1(n9888), .A2(n9396), .ZN(n6368) );
  INV_X1 U6990 ( .A(n6368), .ZN(n6040) );
  INV_X1 U6991 ( .A(n6309), .ZN(n6042) );
  NOR2_X1 U6992 ( .A1(n6043), .A2(n6042), .ZN(n9715) );
  MUX2_X1 U6993 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n7320), .Z(n6047) );
  NAND2_X1 U6994 ( .A1(n6047), .A2(SI_17_), .ZN(n6062) );
  OAI21_X1 U6995 ( .B1(n6047), .B2(SI_17_), .A(n6062), .ZN(n6048) );
  NAND2_X1 U6996 ( .A1(n6049), .A2(n6048), .ZN(n6050) );
  NAND2_X1 U6997 ( .A1(n6050), .A2(n6063), .ZN(n7706) );
  OR2_X1 U6998 ( .A1(n7706), .A2(n5096), .ZN(n6055) );
  INV_X1 U6999 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U7000 ( .A1(n5175), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6053) );
  XNOR2_X1 U7001 ( .A(n6053), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9469) );
  AOI22_X1 U7002 ( .A1(n6086), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6085), .B2(
        n9469), .ZN(n6054) );
  NAND2_X1 U7003 ( .A1(n5751), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6061) );
  INV_X1 U7004 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9460) );
  OR2_X1 U7005 ( .A1(n6246), .A2(n9460), .ZN(n6060) );
  INV_X1 U7006 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9451) );
  NAND2_X1 U7007 ( .A1(n6056), .A2(n9451), .ZN(n6057) );
  NAND2_X1 U7008 ( .A1(n6091), .A2(n6057), .ZN(n9725) );
  OR2_X1 U7009 ( .A1(n6175), .A2(n9725), .ZN(n6059) );
  INV_X1 U7010 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9726) );
  OR2_X1 U7011 ( .A1(n6137), .A2(n9726), .ZN(n6058) );
  NAND2_X1 U7012 ( .A1(n9878), .A2(n9395), .ZN(n6374) );
  OAI21_X2 U7013 ( .B1(n9715), .B2(n9722), .A(n6375), .ZN(n9708) );
  MUX2_X1 U7014 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7320), .Z(n6064) );
  NAND2_X1 U7015 ( .A1(n6064), .A2(SI_18_), .ZN(n6076) );
  INV_X1 U7016 ( .A(n6064), .ZN(n6065) );
  INV_X1 U7017 ( .A(SI_18_), .ZN(n8420) );
  NAND2_X1 U7018 ( .A1(n6065), .A2(n8420), .ZN(n6066) );
  XNOR2_X1 U7019 ( .A(n6079), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9479) );
  AOI22_X1 U7020 ( .A1(n6086), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6085), .B2(
        n9479), .ZN(n6069) );
  NAND2_X1 U7021 ( .A1(n5751), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6074) );
  INV_X1 U7022 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9461) );
  OR2_X1 U7023 ( .A1(n6246), .A2(n9461), .ZN(n6073) );
  INV_X1 U7024 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8296) );
  XNOR2_X1 U7025 ( .A(n6091), .B(n8296), .ZN(n9703) );
  OR2_X1 U7026 ( .A1(n6175), .A2(n9703), .ZN(n6072) );
  INV_X1 U7027 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n6070) );
  OR2_X1 U7028 ( .A1(n6137), .A2(n6070), .ZN(n6071) );
  NAND2_X1 U7029 ( .A1(n9871), .A2(n9719), .ZN(n6306) );
  NAND2_X1 U7030 ( .A1(n6307), .A2(n6306), .ZN(n9707) );
  INV_X1 U7031 ( .A(n6307), .ZN(n6075) );
  MUX2_X1 U7032 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n7320), .Z(n6098) );
  XNOR2_X1 U7033 ( .A(n6098), .B(SI_19_), .ZN(n6100) );
  XNOR2_X1 U7034 ( .A(n6101), .B(n6100), .ZN(n7916) );
  NAND2_X1 U7035 ( .A1(n7916), .A2(n5271), .ZN(n6088) );
  INV_X1 U7036 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6078) );
  NAND2_X1 U7037 ( .A1(n6079), .A2(n6078), .ZN(n6080) );
  INV_X1 U7038 ( .A(n6083), .ZN(n6081) );
  INV_X1 U7039 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6082) );
  INV_X1 U7040 ( .A(n9742), .ZN(n10943) );
  AOI22_X1 U7041 ( .A1(n6086), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n10943), 
        .B2(n6085), .ZN(n6087) );
  NAND2_X1 U7042 ( .A1(n5751), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6097) );
  INV_X1 U7043 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9484) );
  OR2_X1 U7044 ( .A1(n6246), .A2(n9484), .ZN(n6096) );
  INV_X1 U7045 ( .A(n6091), .ZN(n6090) );
  AND2_X1 U7046 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n6089) );
  NAND2_X1 U7047 ( .A1(n6090), .A2(n6089), .ZN(n6105) );
  INV_X1 U7048 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8265) );
  OAI21_X1 U7049 ( .B1(n6091), .B2(n8296), .A(n8265), .ZN(n6092) );
  NAND2_X1 U7050 ( .A1(n6105), .A2(n6092), .ZN(n9696) );
  OR2_X1 U7051 ( .A1(n6175), .A2(n9696), .ZN(n6095) );
  INV_X1 U7052 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6093) );
  OR2_X1 U7053 ( .A1(n6137), .A2(n6093), .ZN(n6094) );
  INV_X1 U7054 ( .A(n6098), .ZN(n6099) );
  INV_X1 U7055 ( .A(SI_19_), .ZN(n8222) );
  MUX2_X1 U7056 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n7320), .Z(n6112) );
  INV_X1 U7057 ( .A(SI_20_), .ZN(n6102) );
  XNOR2_X1 U7058 ( .A(n6112), .B(n6102), .ZN(n6113) );
  XNOR2_X1 U7059 ( .A(n6114), .B(n6113), .ZN(n8067) );
  NAND2_X1 U7060 ( .A1(n8067), .A2(n5271), .ZN(n6104) );
  INV_X1 U7061 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8068) );
  OR2_X1 U7062 ( .A1(n6278), .A2(n8068), .ZN(n6103) );
  NAND2_X1 U7063 ( .A1(n5751), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6111) );
  INV_X1 U7064 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n9679) );
  OR2_X1 U7065 ( .A1(n6137), .A2(n9679), .ZN(n6110) );
  INV_X1 U7066 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9356) );
  NAND2_X1 U7067 ( .A1(n6105), .A2(n9356), .ZN(n6106) );
  NAND2_X1 U7068 ( .A1(n6126), .A2(n6106), .ZN(n9678) );
  OR2_X1 U7069 ( .A1(n6175), .A2(n9678), .ZN(n6109) );
  INV_X1 U7070 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n6107) );
  OR2_X1 U7071 ( .A1(n6246), .A2(n6107), .ZN(n6108) );
  NAND2_X1 U7072 ( .A1(n9861), .A2(n9692), .ZN(n6305) );
  NAND2_X1 U7073 ( .A1(n6304), .A2(n6305), .ZN(n9676) );
  INV_X1 U7074 ( .A(n9676), .ZN(n6441) );
  MUX2_X1 U7075 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n7320), .Z(n6115) );
  NAND2_X1 U7076 ( .A1(n6115), .A2(SI_21_), .ZN(n6132) );
  INV_X1 U7077 ( .A(n6115), .ZN(n6117) );
  INV_X1 U7078 ( .A(SI_21_), .ZN(n6116) );
  NAND2_X1 U7079 ( .A1(n6117), .A2(n6116), .ZN(n6118) );
  NAND2_X1 U7080 ( .A1(n6132), .A2(n6118), .ZN(n6121) );
  INV_X1 U7081 ( .A(n6121), .ZN(n6119) );
  NAND2_X1 U7082 ( .A1(n5549), .A2(n6121), .ZN(n6122) );
  NAND2_X1 U7083 ( .A1(n6133), .A2(n6122), .ZN(n8070) );
  OR2_X1 U7084 ( .A1(n8070), .A2(n5096), .ZN(n6124) );
  INV_X1 U7085 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8065) );
  OR2_X1 U7086 ( .A1(n6278), .A2(n8065), .ZN(n6123) );
  INV_X1 U7087 ( .A(n9856), .ZN(n9663) );
  NAND2_X1 U7088 ( .A1(n6261), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6131) );
  NAND2_X1 U7089 ( .A1(n5751), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6130) );
  NAND2_X1 U7090 ( .A1(n6262), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6129) );
  INV_X1 U7091 ( .A(n6126), .ZN(n6125) );
  NAND2_X1 U7092 ( .A1(n6125), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6138) );
  INV_X1 U7093 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9311) );
  NAND2_X1 U7094 ( .A1(n6126), .A2(n9311), .ZN(n6127) );
  NAND2_X1 U7095 ( .A1(n6138), .A2(n6127), .ZN(n9660) );
  OR2_X1 U7096 ( .A1(n6175), .A2(n9660), .ZN(n6128) );
  NAND4_X1 U7097 ( .A1(n6131), .A2(n6130), .A3(n6129), .A4(n6128), .ZN(n9673)
         );
  INV_X1 U7098 ( .A(n9673), .ZN(n9364) );
  MUX2_X1 U7099 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n7320), .Z(n6146) );
  XNOR2_X1 U7100 ( .A(n6146), .B(SI_22_), .ZN(n6149) );
  XNOR2_X1 U7101 ( .A(n6150), .B(n6149), .ZN(n8628) );
  NAND2_X1 U7102 ( .A1(n8628), .A2(n5271), .ZN(n6135) );
  INV_X1 U7103 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8633) );
  OR2_X1 U7104 ( .A1(n6278), .A2(n8633), .ZN(n6134) );
  NAND2_X1 U7105 ( .A1(n5751), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6144) );
  INV_X1 U7106 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n6136) );
  OR2_X1 U7107 ( .A1(n6137), .A2(n6136), .ZN(n6143) );
  INV_X1 U7108 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9363) );
  NAND2_X1 U7109 ( .A1(n6138), .A2(n9363), .ZN(n6139) );
  NAND2_X1 U7110 ( .A1(n6155), .A2(n6139), .ZN(n9643) );
  OR2_X1 U7111 ( .A1(n9643), .A2(n6175), .ZN(n6142) );
  INV_X1 U7112 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n6140) );
  OR2_X1 U7113 ( .A1(n6246), .A2(n6140), .ZN(n6141) );
  NAND2_X1 U7114 ( .A1(n9851), .A2(n9512), .ZN(n6298) );
  NAND2_X1 U7115 ( .A1(n6299), .A2(n6298), .ZN(n9647) );
  INV_X1 U7116 ( .A(n9647), .ZN(n9640) );
  INV_X1 U7117 ( .A(n6299), .ZN(n6145) );
  INV_X1 U7118 ( .A(n6146), .ZN(n6147) );
  INV_X1 U7119 ( .A(SI_22_), .ZN(n8413) );
  NAND2_X1 U7120 ( .A1(n6147), .A2(n8413), .ZN(n6148) );
  MUX2_X1 U7121 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n7320), .Z(n6162) );
  INV_X1 U7122 ( .A(SI_23_), .ZN(n8215) );
  XNOR2_X1 U7123 ( .A(n6162), .B(n8215), .ZN(n6160) );
  NAND2_X1 U7124 ( .A1(n8753), .A2(n5271), .ZN(n6152) );
  OR2_X1 U7125 ( .A1(n6278), .A2(n7477), .ZN(n6151) );
  NAND2_X1 U7126 ( .A1(n6261), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6154) );
  NAND2_X1 U7127 ( .A1(n5751), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6153) );
  AND2_X1 U7128 ( .A1(n6154), .A2(n6153), .ZN(n6159) );
  INV_X1 U7129 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9278) );
  NAND2_X1 U7130 ( .A1(n6155), .A2(n9278), .ZN(n6156) );
  AND2_X1 U7131 ( .A1(n6173), .A2(n6156), .ZN(n9633) );
  NAND2_X1 U7132 ( .A1(n9633), .A2(n6248), .ZN(n6158) );
  NAND2_X1 U7133 ( .A1(n6262), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6157) );
  OR2_X1 U7134 ( .A1(n9846), .A2(n9613), .ZN(n6300) );
  NAND2_X1 U7135 ( .A1(n9846), .A2(n9613), .ZN(n9610) );
  NAND2_X1 U7136 ( .A1(n9621), .A2(n9628), .ZN(n9620) );
  NAND2_X1 U7137 ( .A1(n6161), .A2(n6160), .ZN(n6165) );
  INV_X1 U7138 ( .A(n6162), .ZN(n6163) );
  NAND2_X1 U7139 ( .A1(n6163), .A2(n8215), .ZN(n6164) );
  MUX2_X1 U7140 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n7320), .Z(n6166) );
  NAND2_X1 U7141 ( .A1(n6166), .A2(SI_24_), .ZN(n6179) );
  OAI21_X1 U7142 ( .B1(n6166), .B2(SI_24_), .A(n6179), .ZN(n6167) );
  NAND2_X1 U7143 ( .A1(n6168), .A2(n6167), .ZN(n6169) );
  INV_X1 U7144 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8770) );
  OR2_X1 U7145 ( .A1(n6278), .A2(n8770), .ZN(n6170) );
  INV_X1 U7146 ( .A(n6173), .ZN(n6172) );
  NAND2_X1 U7147 ( .A1(n6172), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6184) );
  INV_X1 U7148 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9349) );
  NAND2_X1 U7149 ( .A1(n6173), .A2(n9349), .ZN(n6174) );
  NAND2_X1 U7150 ( .A1(n6184), .A2(n6174), .ZN(n9604) );
  OR2_X1 U7151 ( .A1(n9604), .A2(n6175), .ZN(n6178) );
  AOI22_X1 U7152 ( .A1(n5751), .A2(P2_REG0_REG_24__SCAN_IN), .B1(n6262), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n6177) );
  NAND2_X1 U7153 ( .A1(n6261), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6176) );
  NAND2_X1 U7154 ( .A1(n9839), .A2(n9518), .ZN(n6294) );
  NAND3_X1 U7155 ( .A1(n9620), .A2(n9609), .A3(n9610), .ZN(n9608) );
  NAND2_X1 U7156 ( .A1(n9608), .A2(n6395), .ZN(n9587) );
  MUX2_X1 U7157 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(P2_DATAO_REG_25__SCAN_IN), 
        .S(n7320), .Z(n6189) );
  XNOR2_X1 U7158 ( .A(n6189), .B(SI_25_), .ZN(n6192) );
  NAND2_X1 U7159 ( .A1(n8841), .A2(n5271), .ZN(n6182) );
  INV_X1 U7160 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8844) );
  OR2_X1 U7161 ( .A1(n6278), .A2(n8844), .ZN(n6181) );
  INV_X1 U7162 ( .A(n6184), .ZN(n6183) );
  NAND2_X1 U7163 ( .A1(n6183), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6196) );
  INV_X1 U7164 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8483) );
  NAND2_X1 U7165 ( .A1(n6184), .A2(n8483), .ZN(n6185) );
  NAND2_X1 U7166 ( .A1(n6196), .A2(n6185), .ZN(n9594) );
  OR2_X1 U7167 ( .A1(n9594), .A2(n6175), .ZN(n6188) );
  AOI22_X1 U7168 ( .A1(n5751), .A2(P2_REG0_REG_25__SCAN_IN), .B1(n6262), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n6187) );
  NAND2_X1 U7169 ( .A1(n6261), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6186) );
  NAND2_X1 U7170 ( .A1(n9836), .A2(n9614), .ZN(n6406) );
  NAND2_X1 U7171 ( .A1(n9575), .A2(n6406), .ZN(n9520) );
  INV_X1 U7172 ( .A(n6189), .ZN(n6190) );
  INV_X1 U7173 ( .A(SI_25_), .ZN(n8409) );
  NAND2_X1 U7174 ( .A1(n6190), .A2(n8409), .ZN(n6191) );
  MUX2_X1 U7175 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .S(n7320), .Z(n6204) );
  INV_X1 U7176 ( .A(SI_26_), .ZN(n8405) );
  XNOR2_X1 U7177 ( .A(n6204), .B(n8405), .ZN(n6202) );
  NAND2_X1 U7178 ( .A1(n9921), .A2(n5271), .ZN(n6195) );
  INV_X1 U7179 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9924) );
  OR2_X1 U7180 ( .A1(n6278), .A2(n9924), .ZN(n6194) );
  INV_X1 U7181 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8510) );
  NAND2_X1 U7182 ( .A1(n6196), .A2(n8510), .ZN(n6197) );
  INV_X1 U7183 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n6200) );
  NAND2_X1 U7184 ( .A1(n5751), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6199) );
  NAND2_X1 U7185 ( .A1(n6262), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6198) );
  OAI211_X1 U7186 ( .C1(n6246), .C2(n6200), .A(n6199), .B(n6198), .ZN(n6201)
         );
  AOI21_X1 U7187 ( .B1(n9581), .B2(n6248), .A(n6201), .ZN(n9565) );
  INV_X1 U7188 ( .A(n6429), .ZN(n6408) );
  NAND2_X1 U7189 ( .A1(n6203), .A2(n6202), .ZN(n6207) );
  INV_X1 U7190 ( .A(n6204), .ZN(n6205) );
  NAND2_X1 U7191 ( .A1(n6205), .A2(n8405), .ZN(n6206) );
  MUX2_X1 U7192 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n7320), .Z(n6208) );
  NAND2_X1 U7193 ( .A1(n6208), .A2(SI_27_), .ZN(n6221) );
  OAI21_X1 U7194 ( .B1(n6208), .B2(SI_27_), .A(n6221), .ZN(n6209) );
  NAND2_X1 U7195 ( .A1(n6210), .A2(n6209), .ZN(n6211) );
  INV_X1 U7196 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9919) );
  OR2_X1 U7197 ( .A1(n6278), .A2(n9919), .ZN(n6213) );
  XNOR2_X1 U7198 ( .A(n6227), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n9559) );
  NAND2_X1 U7199 ( .A1(n9559), .A2(n6248), .ZN(n6220) );
  INV_X1 U7200 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7201 ( .A1(n5751), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U7202 ( .A1(n6262), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6215) );
  OAI211_X1 U7203 ( .C1(n6246), .C2(n6217), .A(n6216), .B(n6215), .ZN(n6218)
         );
  INV_X1 U7204 ( .A(n6218), .ZN(n6219) );
  NAND2_X1 U7205 ( .A1(n6220), .A2(n6219), .ZN(n9393) );
  INV_X1 U7206 ( .A(n9393), .ZN(n9522) );
  MUX2_X1 U7207 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7320), .Z(n6235) );
  XNOR2_X1 U7208 ( .A(n6235), .B(SI_28_), .ZN(n6238) );
  INV_X1 U7209 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8926) );
  OR2_X1 U7210 ( .A1(n6278), .A2(n8926), .ZN(n6223) );
  INV_X1 U7211 ( .A(n6227), .ZN(n6226) );
  AND2_X1 U7212 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n6225) );
  NAND2_X1 U7213 ( .A1(n6226), .A2(n6225), .ZN(n6242) );
  INV_X1 U7214 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6631) );
  INV_X1 U7215 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8473) );
  OAI21_X1 U7216 ( .B1(n6227), .B2(n6631), .A(n8473), .ZN(n6228) );
  NAND2_X1 U7217 ( .A1(n6242), .A2(n6228), .ZN(n9547) );
  OR2_X1 U7218 ( .A1(n9547), .A2(n6175), .ZN(n6234) );
  INV_X1 U7219 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6231) );
  NAND2_X1 U7220 ( .A1(n6262), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6230) );
  NAND2_X1 U7221 ( .A1(n5751), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6229) );
  OAI211_X1 U7222 ( .C1(n6246), .C2(n6231), .A(n6230), .B(n6229), .ZN(n6232)
         );
  INV_X1 U7223 ( .A(n6232), .ZN(n6233) );
  INV_X1 U7224 ( .A(n6235), .ZN(n6236) );
  INV_X1 U7225 ( .A(SI_28_), .ZN(n8205) );
  NAND2_X1 U7226 ( .A1(n6236), .A2(n8205), .ZN(n6237) );
  INV_X1 U7227 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9917) );
  INV_X1 U7228 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10541) );
  MUX2_X1 U7229 ( .A(n9917), .B(n10541), .S(n7320), .Z(n6249) );
  NAND2_X1 U7230 ( .A1(n9916), .A2(n5271), .ZN(n6241) );
  OR2_X1 U7231 ( .A1(n6278), .A2(n9917), .ZN(n6240) );
  INV_X1 U7232 ( .A(n6242), .ZN(n9535) );
  INV_X1 U7233 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U7234 ( .A1(n5751), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6244) );
  NAND2_X1 U7235 ( .A1(n6262), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6243) );
  OAI211_X1 U7236 ( .C1(n6246), .C2(n6245), .A(n6244), .B(n6243), .ZN(n6247)
         );
  AOI21_X1 U7237 ( .B1(n9535), .B2(n6248), .A(n6247), .ZN(n9304) );
  NAND2_X1 U7238 ( .A1(n9495), .A2(n9304), .ZN(n6292) );
  INV_X1 U7239 ( .A(n6266), .ZN(n6268) );
  INV_X1 U7240 ( .A(SI_29_), .ZN(n8204) );
  MUX2_X1 U7241 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n5740), .Z(n6272) );
  XNOR2_X1 U7242 ( .A(n6272), .B(SI_30_), .ZN(n6269) );
  NAND2_X1 U7243 ( .A1(n8932), .A2(n5271), .ZN(n6254) );
  INV_X1 U7244 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8927) );
  OR2_X1 U7245 ( .A1(n6278), .A2(n8927), .ZN(n6253) );
  NAND2_X1 U7246 ( .A1(n6261), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6257) );
  NAND2_X1 U7247 ( .A1(n5751), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6256) );
  NAND2_X1 U7248 ( .A1(n6262), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6255) );
  AND3_X1 U7249 ( .A1(n6257), .A2(n6256), .A3(n6255), .ZN(n9532) );
  NOR2_X1 U7250 ( .A1(n9503), .A2(n9532), .ZN(n6288) );
  NAND2_X1 U7251 ( .A1(n6259), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6260) );
  XNOR2_X1 U7252 ( .A(n6260), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7781) );
  INV_X1 U7253 ( .A(n7781), .ZN(n8066) );
  NAND2_X1 U7254 ( .A1(n6261), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6265) );
  NAND2_X1 U7255 ( .A1(n6262), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6264) );
  NAND2_X1 U7256 ( .A1(n5751), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6263) );
  NAND3_X1 U7257 ( .A1(n6265), .A2(n6264), .A3(n6263), .ZN(n7362) );
  OAI22_X1 U7258 ( .A1(n6266), .A2(n6288), .B1(n8066), .B2(n7362), .ZN(n6267)
         );
  OAI21_X1 U7259 ( .B1(n6268), .B2(n9503), .A(n6267), .ZN(n6281) );
  INV_X1 U7260 ( .A(n6269), .ZN(n6270) );
  NAND2_X1 U7261 ( .A1(n6271), .A2(n6270), .ZN(n6274) );
  NAND2_X1 U7262 ( .A1(n6272), .A2(SI_30_), .ZN(n6273) );
  MUX2_X1 U7263 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n5740), .Z(n6275) );
  XNOR2_X1 U7264 ( .A(n6275), .B(SI_31_), .ZN(n6276) );
  INV_X1 U7265 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9915) );
  OR2_X1 U7266 ( .A1(n6278), .A2(n9915), .ZN(n6279) );
  INV_X1 U7267 ( .A(n7362), .ZN(n9498) );
  NAND2_X1 U7268 ( .A1(n9503), .A2(n9532), .ZN(n6421) );
  INV_X1 U7269 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6283) );
  INV_X1 U7270 ( .A(n6286), .ZN(n7782) );
  NAND2_X1 U7271 ( .A1(n6258), .A2(n6285), .ZN(n6460) );
  NAND2_X1 U7272 ( .A1(n6460), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6453) );
  XNOR2_X1 U7273 ( .A(n6453), .B(P2_IR_REG_22__SCAN_IN), .ZN(n7776) );
  INV_X1 U7274 ( .A(n7776), .ZN(n8631) );
  AND2_X1 U7275 ( .A1(n8631), .A2(n8066), .ZN(n10679) );
  INV_X1 U7276 ( .A(n10679), .ZN(n6622) );
  INV_X1 U7277 ( .A(n6287), .ZN(n6289) );
  INV_X1 U7278 ( .A(n6288), .ZN(n6422) );
  NAND2_X1 U7279 ( .A1(n6289), .A2(n6422), .ZN(n6428) );
  OR2_X1 U7280 ( .A1(n7776), .A2(n8066), .ZN(n6290) );
  MUX2_X1 U7281 ( .A(n6291), .B(n6428), .S(n6319), .Z(n6427) );
  MUX2_X1 U7282 ( .A(n6293), .B(n6292), .S(n6319), .Z(n6423) );
  NAND2_X1 U7283 ( .A1(n6395), .A2(n6300), .ZN(n6296) );
  NAND2_X1 U7284 ( .A1(n6294), .A2(n9610), .ZN(n6295) );
  MUX2_X1 U7285 ( .A(n6296), .B(n6295), .S(n6319), .Z(n6297) );
  INV_X1 U7286 ( .A(n6297), .ZN(n6393) );
  INV_X1 U7287 ( .A(n6298), .ZN(n6302) );
  NAND2_X1 U7288 ( .A1(n6300), .A2(n6299), .ZN(n6301) );
  MUX2_X1 U7289 ( .A(n6302), .B(n6301), .S(n6319), .Z(n6392) );
  OR2_X1 U7290 ( .A1(n9856), .A2(n9673), .ZN(n9639) );
  INV_X1 U7291 ( .A(n9639), .ZN(n6390) );
  MUX2_X1 U7292 ( .A(n9673), .B(n9856), .S(n6417), .Z(n6389) );
  NAND2_X1 U7293 ( .A1(n9856), .A2(n9673), .ZN(n6303) );
  NAND2_X1 U7294 ( .A1(n6389), .A2(n6303), .ZN(n6387) );
  MUX2_X1 U7295 ( .A(n6305), .B(n6304), .S(n6319), .Z(n6386) );
  MUX2_X1 U7296 ( .A(n6307), .B(n6306), .S(n6319), .Z(n6379) );
  INV_X1 U7297 ( .A(n9722), .ZN(n6373) );
  MUX2_X1 U7298 ( .A(n6308), .B(n6309), .S(n6417), .Z(n6372) );
  NAND2_X1 U7299 ( .A1(n9408), .A2(n10699), .ZN(n6432) );
  NAND2_X1 U7300 ( .A1(n6432), .A2(n6434), .ZN(n6310) );
  AND2_X1 U7301 ( .A1(n6433), .A2(n6310), .ZN(n6313) );
  NAND3_X1 U7302 ( .A1(n6432), .A2(n6434), .A3(n7781), .ZN(n6311) );
  MUX2_X1 U7303 ( .A(n6313), .B(n6312), .S(n6319), .Z(n6318) );
  NAND2_X1 U7304 ( .A1(n6315), .A2(n6314), .ZN(n8145) );
  MUX2_X1 U7305 ( .A(n6315), .B(n6314), .S(n6319), .Z(n6316) );
  OAI211_X1 U7306 ( .C1(n6318), .C2(n8145), .A(n6317), .B(n6316), .ZN(n6323)
         );
  MUX2_X1 U7307 ( .A(n6321), .B(n6320), .S(n6319), .Z(n6322) );
  INV_X1 U7308 ( .A(n9403), .ZN(n7815) );
  NAND2_X1 U7309 ( .A1(n7815), .A2(n10768), .ZN(n7922) );
  INV_X1 U7310 ( .A(n10768), .ZN(n7930) );
  MUX2_X1 U7311 ( .A(n7930), .B(n9403), .S(n6319), .Z(n6324) );
  INV_X1 U7312 ( .A(n10802), .ZN(n7935) );
  NAND2_X1 U7313 ( .A1(n7935), .A2(n6319), .ZN(n6326) );
  NAND2_X1 U7314 ( .A1(n10802), .A2(n6417), .ZN(n6325) );
  MUX2_X1 U7315 ( .A(n6326), .B(n6325), .S(n9789), .Z(n6327) );
  NAND2_X1 U7316 ( .A1(n6328), .A2(n6327), .ZN(n6330) );
  NAND2_X1 U7317 ( .A1(n9402), .A2(n9796), .ZN(n8018) );
  MUX2_X1 U7318 ( .A(n9402), .B(n9796), .S(n6319), .Z(n6329) );
  OAI21_X1 U7319 ( .B1(n6330), .B2(n8018), .A(n6329), .ZN(n6332) );
  NAND3_X1 U7320 ( .A1(n6330), .A2(n8048), .A3(n10819), .ZN(n6331) );
  MUX2_X1 U7321 ( .A(n6333), .B(n8004), .S(n6319), .Z(n6334) );
  MUX2_X1 U7322 ( .A(n6336), .B(n6335), .S(n6319), .Z(n6337) );
  INV_X1 U7323 ( .A(n6338), .ZN(n6340) );
  NAND2_X1 U7324 ( .A1(n10920), .A2(n6345), .ZN(n6339) );
  MUX2_X1 U7325 ( .A(n6340), .B(n6339), .S(n6319), .Z(n6342) );
  NOR2_X1 U7326 ( .A1(n6342), .A2(n6341), .ZN(n6344) );
  NAND2_X1 U7327 ( .A1(n6343), .A2(n6344), .ZN(n6351) );
  NAND2_X1 U7328 ( .A1(n6352), .A2(n6431), .ZN(n6348) );
  INV_X1 U7329 ( .A(n6344), .ZN(n6346) );
  OAI211_X1 U7330 ( .C1(n6346), .C2(n6345), .A(n10920), .B(n8807), .ZN(n6347)
         );
  MUX2_X1 U7331 ( .A(n6348), .B(n6347), .S(n6417), .Z(n6349) );
  INV_X1 U7332 ( .A(n6349), .ZN(n6350) );
  NAND3_X1 U7333 ( .A1(n6351), .A2(n8817), .A3(n6350), .ZN(n6359) );
  INV_X1 U7334 ( .A(n8861), .ZN(n6358) );
  NAND2_X1 U7335 ( .A1(n6353), .A2(n6352), .ZN(n6355) );
  NAND2_X1 U7336 ( .A1(n6355), .A2(n6354), .ZN(n6356) );
  MUX2_X1 U7337 ( .A(n6356), .B(n5157), .S(n6319), .Z(n6357) );
  NAND3_X1 U7338 ( .A1(n6359), .A2(n6358), .A3(n6357), .ZN(n6363) );
  MUX2_X1 U7339 ( .A(n6361), .B(n6360), .S(n6319), .Z(n6362) );
  NAND3_X1 U7340 ( .A1(n6363), .A2(n9766), .A3(n6362), .ZN(n6367) );
  MUX2_X1 U7341 ( .A(n6365), .B(n6364), .S(n6417), .Z(n6366) );
  NAND3_X1 U7342 ( .A1(n6367), .A2(n9756), .A3(n6366), .ZN(n6370) );
  MUX2_X1 U7343 ( .A(n9736), .B(n6368), .S(n6417), .Z(n6369) );
  NAND3_X1 U7344 ( .A1(n9743), .A2(n6370), .A3(n6369), .ZN(n6371) );
  NAND3_X1 U7345 ( .A1(n6373), .A2(n6372), .A3(n6371), .ZN(n6377) );
  MUX2_X1 U7346 ( .A(n6375), .B(n6374), .S(n6417), .Z(n6376) );
  NAND3_X1 U7347 ( .A1(n5357), .A2(n6377), .A3(n6376), .ZN(n6378) );
  NAND2_X1 U7348 ( .A1(n6379), .A2(n6378), .ZN(n6380) );
  NAND2_X1 U7349 ( .A1(n5358), .A2(n6380), .ZN(n6384) );
  NAND2_X1 U7350 ( .A1(n5455), .A2(n6417), .ZN(n6382) );
  NAND2_X1 U7351 ( .A1(n9373), .A2(n6319), .ZN(n6381) );
  MUX2_X1 U7352 ( .A(n6382), .B(n6381), .S(n9868), .Z(n6383) );
  NAND3_X1 U7353 ( .A1(n6441), .A2(n6384), .A3(n6383), .ZN(n6385) );
  NAND3_X1 U7354 ( .A1(n6387), .A2(n6386), .A3(n6385), .ZN(n6388) );
  OAI21_X1 U7355 ( .B1(n6390), .B2(n6389), .A(n6388), .ZN(n6391) );
  NAND2_X1 U7356 ( .A1(n6394), .A2(n9575), .ZN(n6399) );
  NAND2_X1 U7357 ( .A1(n6399), .A2(n6417), .ZN(n6398) );
  NAND2_X1 U7358 ( .A1(n6396), .A2(n6395), .ZN(n6397) );
  NAND2_X1 U7359 ( .A1(n6398), .A2(n6397), .ZN(n6402) );
  INV_X1 U7360 ( .A(n6399), .ZN(n6400) );
  NAND3_X1 U7361 ( .A1(n6400), .A2(n6417), .A3(n9518), .ZN(n6401) );
  NAND2_X1 U7362 ( .A1(n6402), .A2(n6401), .ZN(n6407) );
  INV_X1 U7363 ( .A(n6407), .ZN(n6405) );
  AND2_X1 U7364 ( .A1(n6429), .A2(n6406), .ZN(n6404) );
  INV_X1 U7365 ( .A(n6430), .ZN(n6403) );
  AOI21_X1 U7366 ( .B1(n6405), .B2(n6404), .A(n6403), .ZN(n6412) );
  NAND2_X1 U7367 ( .A1(n6407), .A2(n6406), .ZN(n6410) );
  AOI21_X1 U7368 ( .B1(n6410), .B2(n6409), .A(n6408), .ZN(n6411) );
  INV_X1 U7369 ( .A(n9544), .ZN(n6416) );
  MUX2_X1 U7370 ( .A(n6414), .B(n6413), .S(n6319), .Z(n6415) );
  INV_X1 U7371 ( .A(n9566), .ZN(n9525) );
  NAND2_X1 U7372 ( .A1(n9525), .A2(n6319), .ZN(n6419) );
  NAND2_X1 U7373 ( .A1(n9566), .A2(n6417), .ZN(n6418) );
  MUX2_X1 U7374 ( .A(n6419), .B(n6418), .S(n9819), .Z(n6420) );
  INV_X1 U7375 ( .A(n9805), .ZN(n9499) );
  MUX2_X1 U7376 ( .A(n9805), .B(n7362), .S(n6319), .Z(n6424) );
  OAI21_X1 U7377 ( .B1(n9499), .B2(n9498), .A(n6424), .ZN(n6425) );
  INV_X1 U7378 ( .A(n6428), .ZN(n6448) );
  XNOR2_X1 U7379 ( .A(n9856), .B(n9673), .ZN(n9664) );
  INV_X1 U7380 ( .A(n9664), .ZN(n6443) );
  INV_X1 U7381 ( .A(n9756), .ZN(n9748) );
  AND2_X1 U7382 ( .A1(n10695), .A2(n6432), .ZN(n10677) );
  INV_X1 U7383 ( .A(n8145), .ZN(n8143) );
  NAND3_X1 U7384 ( .A1(n10677), .A2(n7782), .A3(n8143), .ZN(n6435) );
  NAND2_X1 U7385 ( .A1(n6434), .A2(n6433), .ZN(n10704) );
  NOR4_X1 U7386 ( .A1(n7951), .A2(n7779), .A3(n6435), .A4(n10704), .ZN(n6436)
         );
  XNOR2_X1 U7387 ( .A(n9402), .B(n9796), .ZN(n9798) );
  NAND4_X1 U7388 ( .A1(n6436), .A2(n8049), .A3(n7937), .A4(n9798), .ZN(n6437)
         );
  NOR4_X1 U7389 ( .A1(n8006), .A2(n8650), .A3(n6437), .A4(n10919), .ZN(n6438)
         );
  NAND4_X1 U7390 ( .A1(n9766), .A2(n8817), .A3(n8675), .A4(n6438), .ZN(n6439)
         );
  NOR4_X1 U7391 ( .A1(n9722), .A2(n8861), .A3(n9748), .A4(n6439), .ZN(n6440)
         );
  NAND4_X1 U7392 ( .A1(n6441), .A2(n9743), .A3(n5357), .A4(n6440), .ZN(n6442)
         );
  NOR4_X1 U7393 ( .A1(n9647), .A2(n6443), .A3(n6442), .A4(n9689), .ZN(n6444)
         );
  NAND4_X1 U7394 ( .A1(n9588), .A2(n9628), .A3(n9609), .A4(n6444), .ZN(n6445)
         );
  NOR4_X1 U7395 ( .A1(n9544), .A2(n9563), .A3(n9576), .A4(n6445), .ZN(n6446)
         );
  NAND4_X1 U7396 ( .A1(n6448), .A2(n6447), .A3(n9528), .A4(n6446), .ZN(n6449)
         );
  XNOR2_X1 U7397 ( .A(n6449), .B(n9742), .ZN(n6450) );
  AOI211_X1 U7398 ( .C1(n6286), .C2(n6468), .A(n7781), .B(n6450), .ZN(n6451)
         );
  AOI21_X1 U7399 ( .B1(n6452), .B2(n7957), .A(n6451), .ZN(n6467) );
  NAND2_X1 U7400 ( .A1(n6453), .A2(n5216), .ZN(n6454) );
  NAND2_X1 U7401 ( .A1(n6454), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6455) );
  XNOR2_X1 U7402 ( .A(n6455), .B(n5217), .ZN(n6628) );
  OR2_X1 U7403 ( .A1(n6628), .A2(P2_U3152), .ZN(n8754) );
  INV_X1 U7404 ( .A(n6627), .ZN(n6634) );
  NAND2_X1 U7405 ( .A1(n6455), .A2(n5217), .ZN(n6456) );
  NAND2_X1 U7406 ( .A1(n6456), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6457) );
  XNOR2_X1 U7407 ( .A(n6457), .B(P2_IR_REG_24__SCAN_IN), .ZN(n6616) );
  NAND2_X1 U7408 ( .A1(n6458), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6459) );
  XNOR2_X1 U7409 ( .A(n6459), .B(P2_IR_REG_26__SCAN_IN), .ZN(n9922) );
  INV_X1 U7410 ( .A(n6460), .ZN(n6462) );
  NAND2_X1 U7411 ( .A1(n6462), .A2(n6461), .ZN(n6463) );
  NAND2_X1 U7412 ( .A1(n6463), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6464) );
  XNOR2_X1 U7413 ( .A(n6464), .B(P2_IR_REG_25__SCAN_IN), .ZN(n8842) );
  AND2_X1 U7414 ( .A1(n9922), .A2(n8842), .ZN(n6465) );
  NAND2_X1 U7415 ( .A1(n6616), .A2(n6465), .ZN(n7371) );
  INV_X1 U7416 ( .A(n9920), .ZN(n9496) );
  INV_X1 U7417 ( .A(n8925), .ZN(n7392) );
  AND2_X1 U7418 ( .A1(n7776), .A2(n7781), .ZN(n7341) );
  NAND2_X1 U7419 ( .A1(n7392), .A2(n7341), .ZN(n9774) );
  NAND4_X1 U7420 ( .A1(n6634), .A2(n7605), .A3(n9496), .A4(n10924), .ZN(n6466)
         );
  OAI211_X1 U7421 ( .C1(n7776), .C2(n8754), .A(n6466), .B(P2_B_REG_SCAN_IN), 
        .ZN(n6472) );
  AND2_X1 U7422 ( .A1(n6467), .A2(n6472), .ZN(n6471) );
  OR2_X1 U7423 ( .A1(n9742), .A2(n8631), .ZN(n7783) );
  NAND2_X1 U7424 ( .A1(n7783), .A2(n6622), .ZN(n6469) );
  MUX2_X1 U7425 ( .A(n7783), .B(n6469), .S(n6468), .Z(n6470) );
  INV_X1 U7426 ( .A(n6472), .ZN(n6473) );
  INV_X1 U7427 ( .A(n8754), .ZN(n7343) );
  OR2_X1 U7428 ( .A1(n6473), .A2(n7343), .ZN(n6474) );
  AND2_X1 U7429 ( .A1(n9407), .A2(n9295), .ZN(n7743) );
  NAND2_X1 U7430 ( .A1(n10703), .A2(n9295), .ZN(n7614) );
  NAND2_X1 U7431 ( .A1(n6286), .A2(n7781), .ZN(n7927) );
  NAND2_X1 U7432 ( .A1(n9742), .A2(n7776), .ZN(n6476) );
  OR2_X1 U7433 ( .A1(n10680), .A2(n9296), .ZN(n6477) );
  NAND2_X1 U7434 ( .A1(n7614), .A2(n6477), .ZN(n7602) );
  NAND2_X1 U7435 ( .A1(n7602), .A2(n7743), .ZN(n6478) );
  XNOR2_X1 U7436 ( .A(n10711), .B(n9296), .ZN(n7746) );
  NAND2_X1 U7437 ( .A1(n6478), .A2(n7746), .ZN(n6479) );
  XNOR2_X1 U7438 ( .A(n10730), .B(n9296), .ZN(n6481) );
  NAND2_X1 U7439 ( .A1(n6480), .A2(n6481), .ZN(n7741) );
  OAI211_X1 U7440 ( .C1(n7743), .C2(n7602), .A(n6479), .B(n7741), .ZN(n6484)
         );
  INV_X1 U7441 ( .A(n6480), .ZN(n6483) );
  INV_X1 U7442 ( .A(n6481), .ZN(n6482) );
  NAND2_X1 U7443 ( .A1(n6483), .A2(n6482), .ZN(n7742) );
  OR2_X1 U7444 ( .A1(n8147), .A2(n7957), .ZN(n6485) );
  XNOR2_X1 U7445 ( .A(n9296), .B(n7790), .ZN(n6486) );
  INV_X1 U7446 ( .A(n6485), .ZN(n6487) );
  NAND2_X1 U7447 ( .A1(n6487), .A2(n6486), .ZN(n6488) );
  AND2_X1 U7448 ( .A1(n9403), .A2(n9295), .ZN(n6490) );
  XNOR2_X1 U7449 ( .A(n5072), .B(n10768), .ZN(n6489) );
  AND2_X1 U7450 ( .A1(n6490), .A2(n6489), .ZN(n7722) );
  INV_X1 U7451 ( .A(n6489), .ZN(n6492) );
  INV_X1 U7452 ( .A(n6490), .ZN(n6491) );
  NAND2_X1 U7453 ( .A1(n6492), .A2(n6491), .ZN(n7721) );
  XNOR2_X1 U7454 ( .A(n5072), .B(n10802), .ZN(n6493) );
  AND2_X1 U7455 ( .A1(n9789), .A2(n9295), .ZN(n6494) );
  NAND2_X1 U7456 ( .A1(n6493), .A2(n6494), .ZN(n6497) );
  INV_X1 U7457 ( .A(n6493), .ZN(n6496) );
  INV_X1 U7458 ( .A(n6494), .ZN(n6495) );
  NAND2_X1 U7459 ( .A1(n6496), .A2(n6495), .ZN(n6498) );
  AND2_X1 U7460 ( .A1(n6497), .A2(n6498), .ZN(n7733) );
  NAND2_X1 U7461 ( .A1(n7732), .A2(n7733), .ZN(n7731) );
  NAND2_X1 U7462 ( .A1(n7731), .A2(n6498), .ZN(n7853) );
  XNOR2_X1 U7463 ( .A(n5072), .B(n9796), .ZN(n6500) );
  NAND2_X1 U7464 ( .A1(n9402), .A2(n9295), .ZN(n6499) );
  NAND2_X1 U7465 ( .A1(n6500), .A2(n6499), .ZN(n6504) );
  INV_X1 U7466 ( .A(n6499), .ZN(n6502) );
  INV_X1 U7467 ( .A(n6500), .ZN(n6501) );
  NAND2_X1 U7468 ( .A1(n6502), .A2(n6501), .ZN(n6503) );
  AND2_X1 U7469 ( .A1(n6504), .A2(n6503), .ZN(n7854) );
  NAND2_X1 U7470 ( .A1(n7853), .A2(n7854), .ZN(n7852) );
  XNOR2_X1 U7471 ( .A(n10834), .B(n9296), .ZN(n6505) );
  NAND2_X1 U7472 ( .A1(n9788), .A2(n9295), .ZN(n6506) );
  XNOR2_X1 U7473 ( .A(n6505), .B(n6506), .ZN(n7897) );
  INV_X1 U7474 ( .A(n6505), .ZN(n6508) );
  INV_X1 U7475 ( .A(n6506), .ZN(n6507) );
  NAND2_X1 U7476 ( .A1(n6508), .A2(n6507), .ZN(n6509) );
  XNOR2_X1 U7477 ( .A(n10852), .B(n5072), .ZN(n6510) );
  NOR2_X1 U7478 ( .A1(n8648), .A2(n7957), .ZN(n6511) );
  XNOR2_X1 U7479 ( .A(n6510), .B(n6511), .ZN(n8114) );
  INV_X1 U7480 ( .A(n6510), .ZN(n6512) );
  XNOR2_X1 U7481 ( .A(n10865), .B(n5072), .ZN(n6513) );
  OR2_X1 U7482 ( .A1(n8677), .A2(n7957), .ZN(n6514) );
  NAND2_X1 U7483 ( .A1(n6513), .A2(n6514), .ZN(n6518) );
  INV_X1 U7484 ( .A(n6513), .ZN(n6516) );
  INV_X1 U7485 ( .A(n6514), .ZN(n6515) );
  NAND2_X1 U7486 ( .A1(n6516), .A2(n6515), .ZN(n6517) );
  NAND2_X1 U7487 ( .A1(n6518), .A2(n6517), .ZN(n8136) );
  XNOR2_X1 U7488 ( .A(n8811), .B(n9296), .ZN(n6519) );
  NOR2_X1 U7489 ( .A1(n8664), .A2(n7957), .ZN(n6520) );
  XNOR2_X1 U7490 ( .A(n6519), .B(n6520), .ZN(n8161) );
  XNOR2_X1 U7491 ( .A(n10939), .B(n5072), .ZN(n6521) );
  NOR2_X1 U7492 ( .A1(n9399), .A2(n7957), .ZN(n6522) );
  XNOR2_X1 U7493 ( .A(n6521), .B(n6522), .ZN(n8661) );
  INV_X1 U7494 ( .A(n6521), .ZN(n6523) );
  NAND2_X1 U7495 ( .A1(n6523), .A2(n6522), .ZN(n6524) );
  NAND2_X1 U7496 ( .A1(n6525), .A2(n6524), .ZN(n8777) );
  XNOR2_X1 U7497 ( .A(n8858), .B(n5072), .ZN(n6526) );
  OR2_X1 U7498 ( .A1(n9398), .A2(n7957), .ZN(n6527) );
  NAND2_X1 U7499 ( .A1(n6526), .A2(n6527), .ZN(n6531) );
  INV_X1 U7500 ( .A(n6526), .ZN(n6529) );
  INV_X1 U7501 ( .A(n6527), .ZN(n6528) );
  NAND2_X1 U7502 ( .A1(n6529), .A2(n6528), .ZN(n6530) );
  NAND2_X1 U7503 ( .A1(n6531), .A2(n6530), .ZN(n8778) );
  XNOR2_X1 U7504 ( .A(n8857), .B(n5072), .ZN(n6532) );
  OR2_X1 U7505 ( .A1(n9775), .A2(n7957), .ZN(n6533) );
  NAND2_X1 U7506 ( .A1(n6532), .A2(n6533), .ZN(n6537) );
  INV_X1 U7507 ( .A(n6532), .ZN(n6535) );
  INV_X1 U7508 ( .A(n6533), .ZN(n6534) );
  NAND2_X1 U7509 ( .A1(n6535), .A2(n6534), .ZN(n6536) );
  AND2_X1 U7510 ( .A1(n6537), .A2(n6536), .ZN(n8800) );
  NAND2_X1 U7511 ( .A1(n8799), .A2(n8800), .ZN(n8798) );
  NAND2_X1 U7512 ( .A1(n8798), .A2(n6537), .ZN(n8897) );
  XNOR2_X1 U7513 ( .A(n9781), .B(n5072), .ZN(n6538) );
  OR2_X1 U7514 ( .A1(n9508), .A2(n7957), .ZN(n6539) );
  NAND2_X1 U7515 ( .A1(n6538), .A2(n6539), .ZN(n6543) );
  INV_X1 U7516 ( .A(n6538), .ZN(n6541) );
  INV_X1 U7517 ( .A(n6539), .ZN(n6540) );
  NAND2_X1 U7518 ( .A1(n6541), .A2(n6540), .ZN(n6542) );
  AND2_X1 U7519 ( .A1(n6543), .A2(n6542), .ZN(n8898) );
  NAND2_X1 U7520 ( .A1(n8897), .A2(n8898), .ZN(n8896) );
  NAND2_X1 U7521 ( .A1(n8896), .A2(n6543), .ZN(n8918) );
  XNOR2_X1 U7522 ( .A(n9888), .B(n5072), .ZN(n6544) );
  OR2_X1 U7523 ( .A1(n9396), .A2(n7957), .ZN(n6545) );
  NAND2_X1 U7524 ( .A1(n6544), .A2(n6545), .ZN(n6549) );
  INV_X1 U7525 ( .A(n6544), .ZN(n6547) );
  INV_X1 U7526 ( .A(n6545), .ZN(n6546) );
  NAND2_X1 U7527 ( .A1(n6547), .A2(n6546), .ZN(n6548) );
  AND2_X1 U7528 ( .A1(n6549), .A2(n6548), .ZN(n8919) );
  NAND2_X1 U7529 ( .A1(n8918), .A2(n8919), .ZN(n8917) );
  NAND2_X1 U7530 ( .A1(n8917), .A2(n6549), .ZN(n9328) );
  XNOR2_X1 U7531 ( .A(n9883), .B(n5072), .ZN(n6550) );
  OR2_X1 U7532 ( .A1(n9718), .A2(n7957), .ZN(n6551) );
  NAND2_X1 U7533 ( .A1(n6550), .A2(n6551), .ZN(n6555) );
  INV_X1 U7534 ( .A(n6550), .ZN(n6553) );
  INV_X1 U7535 ( .A(n6551), .ZN(n6552) );
  NAND2_X1 U7536 ( .A1(n6553), .A2(n6552), .ZN(n6554) );
  AND2_X1 U7537 ( .A1(n6555), .A2(n6554), .ZN(n9329) );
  XNOR2_X1 U7538 ( .A(n9878), .B(n5072), .ZN(n6556) );
  OR2_X1 U7539 ( .A1(n9395), .A2(n7957), .ZN(n6557) );
  AND2_X1 U7540 ( .A1(n6556), .A2(n6557), .ZN(n9339) );
  INV_X1 U7541 ( .A(n6556), .ZN(n6559) );
  INV_X1 U7542 ( .A(n6557), .ZN(n6558) );
  NAND2_X1 U7543 ( .A1(n6559), .A2(n6558), .ZN(n9337) );
  XNOR2_X1 U7544 ( .A(n9871), .B(n5072), .ZN(n6560) );
  NOR2_X1 U7545 ( .A1(n9719), .A2(n7957), .ZN(n6561) );
  XNOR2_X1 U7546 ( .A(n6560), .B(n6561), .ZN(n9369) );
  INV_X1 U7547 ( .A(n6560), .ZN(n6562) );
  XNOR2_X1 U7548 ( .A(n9868), .B(n5072), .ZN(n6563) );
  NOR2_X1 U7549 ( .A1(n9373), .A2(n7957), .ZN(n6564) );
  XNOR2_X1 U7550 ( .A(n6563), .B(n6564), .ZN(n9284) );
  INV_X1 U7551 ( .A(n6563), .ZN(n6565) );
  NAND2_X1 U7552 ( .A1(n6565), .A2(n6564), .ZN(n6566) );
  NAND2_X1 U7553 ( .A1(n6567), .A2(n6566), .ZN(n9355) );
  XNOR2_X1 U7554 ( .A(n9861), .B(n5072), .ZN(n6568) );
  NOR2_X1 U7555 ( .A1(n9692), .A2(n7957), .ZN(n6569) );
  XNOR2_X1 U7556 ( .A(n6568), .B(n6569), .ZN(n9354) );
  INV_X1 U7557 ( .A(n6568), .ZN(n6570) );
  NAND2_X1 U7558 ( .A1(n6570), .A2(n6569), .ZN(n6571) );
  XNOR2_X1 U7559 ( .A(n9856), .B(n9296), .ZN(n6574) );
  NAND2_X1 U7560 ( .A1(n9673), .A2(n9295), .ZN(n6572) );
  XNOR2_X1 U7561 ( .A(n6574), .B(n6572), .ZN(n9309) );
  INV_X1 U7562 ( .A(n6572), .ZN(n6573) );
  NAND2_X1 U7563 ( .A1(n6574), .A2(n6573), .ZN(n6575) );
  XNOR2_X1 U7564 ( .A(n9851), .B(n5072), .ZN(n6576) );
  INV_X1 U7565 ( .A(n9512), .ZN(n9667) );
  NAND2_X1 U7566 ( .A1(n9667), .A2(n9295), .ZN(n6577) );
  NAND2_X1 U7567 ( .A1(n6576), .A2(n6577), .ZN(n6581) );
  INV_X1 U7568 ( .A(n6576), .ZN(n6579) );
  INV_X1 U7569 ( .A(n6577), .ZN(n6578) );
  NAND2_X1 U7570 ( .A1(n6579), .A2(n6578), .ZN(n6580) );
  NAND2_X1 U7571 ( .A1(n6581), .A2(n6580), .ZN(n9361) );
  XNOR2_X1 U7572 ( .A(n9846), .B(n9296), .ZN(n6582) );
  NOR2_X1 U7573 ( .A1(n9613), .A2(n7957), .ZN(n9276) );
  NAND2_X1 U7574 ( .A1(n9277), .A2(n9276), .ZN(n6586) );
  INV_X1 U7575 ( .A(n6582), .ZN(n6583) );
  OR2_X1 U7576 ( .A1(n6584), .A2(n6583), .ZN(n6585) );
  NAND2_X1 U7577 ( .A1(n6586), .A2(n6585), .ZN(n6589) );
  XNOR2_X1 U7578 ( .A(n9839), .B(n5072), .ZN(n6587) );
  XNOR2_X1 U7579 ( .A(n6589), .B(n6587), .ZN(n9348) );
  NOR2_X1 U7580 ( .A1(n9518), .A2(n7957), .ZN(n9347) );
  NAND2_X1 U7581 ( .A1(n9348), .A2(n9347), .ZN(n9317) );
  INV_X1 U7582 ( .A(n6587), .ZN(n6588) );
  NAND2_X1 U7583 ( .A1(n6589), .A2(n6588), .ZN(n9316) );
  XNOR2_X1 U7584 ( .A(n9836), .B(n5072), .ZN(n6594) );
  INV_X1 U7585 ( .A(n6594), .ZN(n6590) );
  NOR2_X1 U7586 ( .A1(n9614), .A2(n7957), .ZN(n6593) );
  NAND2_X1 U7587 ( .A1(n6590), .A2(n6593), .ZN(n6592) );
  AND2_X1 U7588 ( .A1(n9316), .A2(n6592), .ZN(n6591) );
  NAND2_X1 U7589 ( .A1(n9317), .A2(n6591), .ZN(n9379) );
  XNOR2_X1 U7590 ( .A(n9830), .B(n5072), .ZN(n6597) );
  NOR2_X1 U7591 ( .A1(n9565), .A2(n7957), .ZN(n6598) );
  XNOR2_X1 U7592 ( .A(n6597), .B(n6598), .ZN(n9380) );
  INV_X1 U7593 ( .A(n6592), .ZN(n6595) );
  XNOR2_X1 U7594 ( .A(n6594), .B(n6593), .ZN(n9318) );
  NAND2_X1 U7595 ( .A1(n9379), .A2(n6596), .ZN(n6601) );
  INV_X1 U7596 ( .A(n6597), .ZN(n6599) );
  NAND2_X1 U7597 ( .A1(n6599), .A2(n6598), .ZN(n6600) );
  XNOR2_X1 U7598 ( .A(n9561), .B(n5072), .ZN(n9292) );
  NAND2_X1 U7599 ( .A1(n9393), .A2(n9295), .ZN(n9290) );
  XNOR2_X1 U7600 ( .A(n9292), .B(n9290), .ZN(n9293) );
  XNOR2_X1 U7601 ( .A(n9294), .B(n9293), .ZN(n6621) );
  NOR4_X1 U7602 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6606) );
  NOR4_X1 U7603 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6605) );
  NOR4_X1 U7604 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6604) );
  NOR4_X1 U7605 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6603) );
  NAND4_X1 U7606 ( .A1(n6606), .A2(n6605), .A3(n6604), .A4(n6603), .ZN(n6615)
         );
  NOR2_X1 U7607 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6610) );
  NOR4_X1 U7608 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6609) );
  NOR4_X1 U7609 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6608) );
  NOR4_X1 U7610 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6607) );
  NAND4_X1 U7611 ( .A1(n6610), .A2(n6609), .A3(n6608), .A4(n6607), .ZN(n6614)
         );
  INV_X1 U7612 ( .A(P2_B_REG_SCAN_IN), .ZN(n6611) );
  INV_X1 U7613 ( .A(n6616), .ZN(n8771) );
  AOI221_X1 U7614 ( .B1(P2_B_REG_SCAN_IN), .B2(n6616), .C1(n6611), .C2(n8771), 
        .A(n8842), .ZN(n6612) );
  INV_X1 U7615 ( .A(n6612), .ZN(n6613) );
  OAI21_X1 U7616 ( .B1(n6615), .B2(n6614), .A(n7349), .ZN(n7767) );
  OR2_X1 U7617 ( .A1(n6616), .A2(n9922), .ZN(n7353) );
  INV_X1 U7618 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n7356) );
  NAND2_X1 U7619 ( .A1(n7349), .A2(n7356), .ZN(n6617) );
  NAND2_X1 U7620 ( .A1(n7353), .A2(n6617), .ZN(n7924) );
  INV_X1 U7621 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n7352) );
  NOR2_X1 U7622 ( .A1(n9922), .A2(n8842), .ZN(n7351) );
  AOI21_X1 U7623 ( .B1(n7349), .B2(n7352), .A(n7351), .ZN(n7923) );
  INV_X1 U7624 ( .A(n7923), .ZN(n7768) );
  NOR2_X1 U7625 ( .A1(n7924), .A2(n7768), .ZN(n6618) );
  NAND2_X1 U7626 ( .A1(n7767), .A2(n6618), .ZN(n6626) );
  INV_X1 U7627 ( .A(n7605), .ZN(n6619) );
  NOR2_X1 U7628 ( .A1(n6626), .A2(n6619), .ZN(n6635) );
  NAND2_X1 U7629 ( .A1(n6627), .A2(n10679), .ZN(n10989) );
  INV_X1 U7630 ( .A(n7341), .ZN(n7369) );
  AND2_X1 U7631 ( .A1(n10989), .A2(n7369), .ZN(n6620) );
  NAND2_X1 U7632 ( .A1(n6635), .A2(n6620), .ZN(n9391) );
  NAND2_X1 U7633 ( .A1(n6635), .A2(n5182), .ZN(n6625) );
  NOR2_X1 U7634 ( .A1(n9742), .A2(n7776), .ZN(n6623) );
  NAND2_X1 U7635 ( .A1(n6286), .A2(n6623), .ZN(n10729) );
  INV_X1 U7636 ( .A(n7769), .ZN(n6624) );
  INV_X1 U7637 ( .A(n9559), .ZN(n6632) );
  NAND2_X1 U7638 ( .A1(n6626), .A2(n7769), .ZN(n7607) );
  NAND2_X1 U7639 ( .A1(n6627), .A2(n7341), .ZN(n7606) );
  AND3_X1 U7640 ( .A1(n7606), .A2(n7371), .A3(n6628), .ZN(n6629) );
  NAND2_X1 U7641 ( .A1(n7607), .A2(n6629), .ZN(n6630) );
  NAND2_X1 U7642 ( .A1(n6630), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9386) );
  OAI22_X1 U7643 ( .A1(n6632), .A2(n9386), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6631), .ZN(n6633) );
  INV_X1 U7644 ( .A(n6633), .ZN(n6638) );
  AND2_X1 U7645 ( .A1(n8925), .A2(n7341), .ZN(n10926) );
  NAND2_X1 U7646 ( .A1(n9384), .A2(n10926), .ZN(n9372) );
  NAND2_X1 U7647 ( .A1(n9384), .A2(n10924), .ZN(n9371) );
  OAI22_X1 U7648 ( .A1(n9566), .A2(n9372), .B1(n9371), .B2(n9565), .ZN(n6636)
         );
  INV_X1 U7649 ( .A(n6636), .ZN(n6637) );
  NAND4_X1 U7650 ( .A1(n5701), .A2(n5700), .A3(n6638), .A4(n6637), .ZN(
        P2_U3216) );
  INV_X1 U7651 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n8599) );
  INV_X1 U7652 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6654) );
  NAND2_X1 U7653 ( .A1(n8599), .A2(n6654), .ZN(n6642) );
  OAI21_X1 U7654 ( .B1(n6646), .B2(n6662), .A(P1_IR_REG_28__SCAN_IN), .ZN(
        n6645) );
  INV_X1 U7655 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8382) );
  NAND2_X1 U7656 ( .A1(n7662), .A2(n8947), .ZN(n6651) );
  OR2_X1 U7657 ( .A1(n6648), .A2(n6662), .ZN(n6649) );
  XNOR2_X1 U7658 ( .A(n6649), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7293) );
  AOI22_X1 U7659 ( .A1(n7029), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7028), .B2(
        n7293), .ZN(n6650) );
  NAND2_X1 U7660 ( .A1(n6655), .A2(n6654), .ZN(n6657) );
  NAND2_X1 U7661 ( .A1(n6657), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6653) );
  XNOR2_X1 U7662 ( .A(n6653), .B(n8599), .ZN(n10549) );
  OR2_X1 U7663 ( .A1(n6655), .A2(n6654), .ZN(n6656) );
  NAND2_X1 U7664 ( .A1(n6657), .A2(n6656), .ZN(n8848) );
  NAND2_X1 U7665 ( .A1(n5121), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6658) );
  XNOR2_X1 U7666 ( .A(n6658), .B(n8595), .ZN(n8774) );
  NAND2_X1 U7667 ( .A1(n5147), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6660) );
  NAND2_X1 U7668 ( .A1(n6660), .A2(n8583), .ZN(n6659) );
  XNOR2_X1 U7669 ( .A(n6660), .B(P1_IR_REG_20__SCAN_IN), .ZN(n9167) );
  INV_X1 U7670 ( .A(n7693), .ZN(n6661) );
  INV_X1 U7671 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6662) );
  INV_X1 U7672 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10534) );
  NAND2_X1 U7673 ( .A1(n6706), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6673) );
  INV_X1 U7674 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n6665) );
  OR2_X1 U7675 ( .A1(n8941), .A2(n6665), .ZN(n6672) );
  INV_X1 U7676 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n6666) );
  OR2_X1 U7677 ( .A1(n8942), .A2(n6666), .ZN(n6671) );
  NAND2_X1 U7678 ( .A1(n6819), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6834) );
  INV_X1 U7679 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6833) );
  NOR2_X1 U7680 ( .A1(n6834), .A2(n6833), .ZN(n6855) );
  NAND2_X1 U7681 ( .A1(n6855), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6872) );
  INV_X1 U7682 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6871) );
  INV_X1 U7683 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7315) );
  INV_X1 U7684 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6919) );
  NAND2_X1 U7685 ( .A1(n6938), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6957) );
  INV_X1 U7686 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6956) );
  INV_X1 U7687 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7973) );
  NAND2_X1 U7688 ( .A1(n6978), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6691) );
  NAND2_X1 U7689 ( .A1(n6669), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6999) );
  OAI21_X1 U7690 ( .B1(n6669), .B2(P1_REG3_REG_16__SCAN_IN), .A(n6999), .ZN(
        n10374) );
  OR2_X1 U7691 ( .A1(n6781), .A2(n10374), .ZN(n6670) );
  NAND4_X1 U7692 ( .A1(n6673), .A2(n6672), .A3(n6671), .A4(n6670), .ZN(n10349)
         );
  NAND2_X1 U7693 ( .A1(n7300), .A2(n7693), .ZN(n6689) );
  NAND2_X1 U7694 ( .A1(n6674), .A2(n8369), .ZN(n6675) );
  NAND2_X1 U7695 ( .A1(n6677), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6678) );
  AND2_X1 U7696 ( .A1(n8630), .A2(n7218), .ZN(n6679) );
  NOR2_X1 U7697 ( .A1(n6689), .A2(n6679), .ZN(n6754) );
  AND2_X1 U7698 ( .A1(n10349), .A2(n9196), .ZN(n6680) );
  AOI21_X1 U7699 ( .B1(n10513), .B2(n6719), .A(n6680), .ZN(n6995) );
  NOR2_X1 U7700 ( .A1(n6681), .A2(n6662), .ZN(n6682) );
  MUX2_X1 U7701 ( .A(n6662), .B(n6682), .S(P1_IR_REG_15__SCAN_IN), .Z(n6683)
         );
  INV_X1 U7702 ( .A(n6683), .ZN(n6685) );
  INV_X1 U7703 ( .A(n6648), .ZN(n6684) );
  NAND2_X1 U7704 ( .A1(n6685), .A2(n6684), .ZN(n10111) );
  INV_X1 U7705 ( .A(n10111), .ZN(n6686) );
  AOI22_X1 U7706 ( .A1(n7029), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7028), .B2(
        n6686), .ZN(n6687) );
  INV_X2 U7707 ( .A(n6689), .ZN(n9192) );
  NAND2_X1 U7708 ( .A1(n10395), .A2(n9192), .ZN(n6698) );
  NAND2_X1 U7709 ( .A1(n7205), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6696) );
  INV_X1 U7710 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n6690) );
  OR2_X1 U7711 ( .A1(n6761), .A2(n6690), .ZN(n6695) );
  OR2_X1 U7712 ( .A1(n6978), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6692) );
  NAND2_X1 U7713 ( .A1(n6692), .A2(n6691), .ZN(n10389) );
  OR2_X1 U7714 ( .A1(n6781), .A2(n10389), .ZN(n6694) );
  INV_X1 U7715 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10390) );
  OR2_X1 U7716 ( .A1(n8942), .A2(n10390), .ZN(n6693) );
  NAND4_X1 U7717 ( .A1(n6696), .A2(n6695), .A3(n6694), .A4(n6693), .ZN(n10399)
         );
  NAND2_X1 U7718 ( .A1(n10399), .A2(n6719), .ZN(n6697) );
  NAND2_X1 U7719 ( .A1(n6698), .A2(n6697), .ZN(n6700) );
  AOI21_X1 U7720 ( .B1(n8630), .B2(n7693), .A(n5073), .ZN(n6699) );
  NAND2_X1 U7721 ( .A1(n7222), .A2(n6699), .ZN(n7692) );
  XNOR2_X1 U7722 ( .A(n6700), .B(n6752), .ZN(n9978) );
  AND2_X1 U7723 ( .A1(n10399), .A2(n9196), .ZN(n6701) );
  AOI21_X1 U7724 ( .B1(n10395), .B2(n6719), .A(n6701), .ZN(n10073) );
  NAND2_X1 U7725 ( .A1(n9978), .A2(n10073), .ZN(n6704) );
  INV_X1 U7726 ( .A(n6704), .ZN(n6994) );
  INV_X1 U7727 ( .A(n6995), .ZN(n9981) );
  AOI22_X1 U7728 ( .A1(n10513), .A2(n9192), .B1(n6719), .B2(n10349), .ZN(n6702) );
  XNOR2_X1 U7729 ( .A(n6702), .B(n7154), .ZN(n9982) );
  INV_X1 U7730 ( .A(n9982), .ZN(n6703) );
  AOI21_X1 U7731 ( .B1(n9981), .B2(n6704), .A(n6703), .ZN(n6993) );
  INV_X1 U7732 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6705) );
  INV_X1 U7733 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n8622) );
  NAND2_X1 U7734 ( .A1(n7205), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6708) );
  NAND2_X1 U7735 ( .A1(n6706), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6707) );
  NOR2_X1 U7736 ( .A1(n5740), .A2(n6711), .ZN(n6713) );
  XNOR2_X1 U7737 ( .A(n6713), .B(n6712), .ZN(n10550) );
  MUX2_X1 U7738 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10550), .S(n7263), .Z(n7699)
         );
  INV_X1 U7739 ( .A(n7300), .ZN(n6714) );
  AOI22_X1 U7740 ( .A1(n7699), .A2(n9192), .B1(n6714), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n6715) );
  NAND2_X1 U7741 ( .A1(n6716), .A2(n6715), .ZN(n7581) );
  INV_X1 U7742 ( .A(n7581), .ZN(n6717) );
  NAND2_X1 U7743 ( .A1(n6717), .A2(n7154), .ZN(n6722) );
  INV_X1 U7744 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10633) );
  NOR2_X1 U7745 ( .A1(n7300), .A2(n10633), .ZN(n6718) );
  AOI21_X1 U7746 ( .B1(n7699), .B2(n6719), .A(n6718), .ZN(n6720) );
  NAND2_X1 U7747 ( .A1(n7583), .A2(n7581), .ZN(n7582) );
  NAND2_X1 U7748 ( .A1(n6722), .A2(n7582), .ZN(n6738) );
  INV_X1 U7749 ( .A(n6738), .ZN(n6734) );
  INV_X1 U7750 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10624) );
  INV_X1 U7751 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7243) );
  NAND2_X1 U7752 ( .A1(n6735), .A2(n6719), .ZN(n6731) );
  NAND2_X1 U7753 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6726) );
  MUX2_X1 U7754 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6726), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n6729) );
  INV_X1 U7755 ( .A(n6727), .ZN(n6728) );
  NAND2_X1 U7756 ( .A1(n6736), .A2(n9192), .ZN(n6730) );
  NAND2_X1 U7757 ( .A1(n6731), .A2(n6730), .ZN(n6732) );
  XNOR2_X1 U7758 ( .A(n6732), .B(n6752), .ZN(n6737) );
  INV_X1 U7759 ( .A(n6737), .ZN(n6733) );
  NAND2_X1 U7760 ( .A1(n6734), .A2(n6733), .ZN(n7638) );
  NAND2_X1 U7761 ( .A1(n7638), .A2(n7640), .ZN(n6739) );
  NAND2_X1 U7762 ( .A1(n6738), .A2(n6737), .ZN(n7639) );
  NAND2_X1 U7763 ( .A1(n6739), .A2(n7639), .ZN(n10045) );
  INV_X1 U7764 ( .A(n6762), .ZN(n6898) );
  NAND2_X1 U7765 ( .A1(n6898), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6745) );
  INV_X1 U7766 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10657) );
  INV_X1 U7767 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n7242) );
  OR2_X1 U7768 ( .A1(n6761), .A2(n7242), .ZN(n6743) );
  NAND2_X1 U7769 ( .A1(n7642), .A2(n6719), .ZN(n6751) );
  INV_X1 U7770 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7328) );
  OR2_X1 U7771 ( .A1(n6727), .A2(n6662), .ZN(n6788) );
  INV_X1 U7772 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8556) );
  NAND2_X1 U7773 ( .A1(n6788), .A2(n8556), .ZN(n6767) );
  OAI21_X1 U7774 ( .B1(n6788), .B2(n8556), .A(n6767), .ZN(n10658) );
  NAND2_X1 U7775 ( .A1(n10720), .A2(n9192), .ZN(n6750) );
  NAND2_X1 U7776 ( .A1(n6751), .A2(n6750), .ZN(n6753) );
  AOI22_X1 U7777 ( .A1(n7642), .A2(n6754), .B1(n6719), .B2(n10720), .ZN(n6756)
         );
  NAND2_X1 U7778 ( .A1(n6755), .A2(n6756), .ZN(n6760) );
  INV_X1 U7779 ( .A(n6755), .ZN(n6758) );
  NAND2_X1 U7780 ( .A1(n6758), .A2(n6757), .ZN(n6759) );
  NAND2_X1 U7781 ( .A1(n10045), .A2(n10046), .ZN(n10044) );
  NAND2_X1 U7782 ( .A1(n10044), .A2(n6760), .ZN(n7807) );
  NAND2_X1 U7783 ( .A1(n7205), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6766) );
  INV_X1 U7784 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7241) );
  OR2_X1 U7785 ( .A1(n6761), .A2(n7241), .ZN(n6765) );
  INV_X1 U7786 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10756) );
  OR2_X1 U7787 ( .A1(n6762), .A2(n10756), .ZN(n6764) );
  OR2_X1 U7788 ( .A1(n6781), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6763) );
  NAND2_X1 U7789 ( .A1(n10103), .A2(n6719), .ZN(n6773) );
  OR2_X1 U7790 ( .A1(n6746), .A2(n7325), .ZN(n6771) );
  INV_X1 U7791 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7326) );
  OR2_X1 U7792 ( .A1(n8949), .A2(n7326), .ZN(n6769) );
  NAND2_X1 U7793 ( .A1(n6767), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6768) );
  XNOR2_X1 U7794 ( .A(n6768), .B(P1_IR_REG_3__SCAN_IN), .ZN(n7277) );
  INV_X1 U7795 ( .A(n7277), .ZN(n7495) );
  AOI22_X1 U7796 ( .A1(n10103), .A2(n9196), .B1(n6719), .B2(n9093), .ZN(n6776)
         );
  XNOR2_X1 U7797 ( .A(n6775), .B(n6776), .ZN(n7808) );
  NAND2_X1 U7798 ( .A1(n7807), .A2(n7808), .ZN(n7806) );
  INV_X1 U7799 ( .A(n6775), .ZN(n6777) );
  NAND2_X1 U7800 ( .A1(n6777), .A2(n6776), .ZN(n6778) );
  NAND2_X1 U7801 ( .A1(n7806), .A2(n6778), .ZN(n7846) );
  INV_X1 U7802 ( .A(n7846), .ZN(n6797) );
  INV_X1 U7803 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6779) );
  OR2_X1 U7804 ( .A1(n6761), .A2(n6779), .ZN(n6785) );
  INV_X1 U7805 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7889) );
  OR2_X1 U7806 ( .A1(n8942), .A2(n7889), .ZN(n6784) );
  INV_X1 U7807 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6780) );
  XNOR2_X1 U7808 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n7888) );
  OR2_X1 U7809 ( .A1(n6786), .A2(n6662), .ZN(n6787) );
  NAND2_X1 U7810 ( .A1(n6788), .A2(n6787), .ZN(n6805) );
  INV_X1 U7811 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8555) );
  XNOR2_X1 U7812 ( .A(n6805), .B(n8555), .ZN(n7278) );
  INV_X1 U7813 ( .A(n7278), .ZN(n7682) );
  INV_X1 U7814 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7329) );
  NAND2_X1 U7815 ( .A1(n7893), .A2(n9192), .ZN(n6789) );
  NAND2_X1 U7816 ( .A1(n6790), .A2(n6789), .ZN(n6791) );
  XOR2_X1 U7817 ( .A(n6791), .B(n6752), .Z(n6795) );
  INV_X1 U7818 ( .A(n6795), .ZN(n6792) );
  AOI22_X1 U7819 ( .A1(n10102), .A2(n9196), .B1(n6719), .B2(n7893), .ZN(n6793)
         );
  INV_X1 U7820 ( .A(n6793), .ZN(n6794) );
  NAND2_X1 U7821 ( .A1(n6795), .A2(n6794), .ZN(n7844) );
  INV_X1 U7822 ( .A(n7844), .ZN(n6796) );
  AOI21_X1 U7823 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6798) );
  NOR2_X1 U7824 ( .A1(n6798), .A2(n6819), .ZN(n10789) );
  NAND2_X1 U7825 ( .A1(n7016), .A2(n10789), .ZN(n6804) );
  INV_X1 U7826 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7240) );
  OR2_X1 U7827 ( .A1(n6761), .A2(n7240), .ZN(n6803) );
  INV_X1 U7828 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6799) );
  OR2_X1 U7829 ( .A1(n8941), .A2(n6799), .ZN(n6802) );
  INV_X1 U7830 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6800) );
  OR2_X1 U7831 ( .A1(n8942), .A2(n6800), .ZN(n6801) );
  NAND2_X1 U7832 ( .A1(n10101), .A2(n6719), .ZN(n6810) );
  OAI21_X1 U7833 ( .B1(n6805), .B2(P1_IR_REG_4__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6806) );
  XNOR2_X1 U7834 ( .A(n6806), .B(P1_IR_REG_5__SCAN_IN), .ZN(n7280) );
  INV_X1 U7835 ( .A(n7280), .ZN(n7532) );
  OR2_X1 U7836 ( .A1(n6746), .A2(n7333), .ZN(n6808) );
  INV_X1 U7837 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7332) );
  OR2_X1 U7838 ( .A1(n8949), .A2(n7332), .ZN(n6807) );
  NAND2_X1 U7839 ( .A1(n10792), .A2(n9192), .ZN(n6809) );
  NAND2_X1 U7840 ( .A1(n6810), .A2(n6809), .ZN(n6811) );
  XNOR2_X1 U7841 ( .A(n6811), .B(n6752), .ZN(n6815) );
  NAND2_X1 U7842 ( .A1(n6814), .A2(n6815), .ZN(n8090) );
  NAND2_X1 U7843 ( .A1(n10101), .A2(n9196), .ZN(n6813) );
  NAND2_X1 U7844 ( .A1(n10792), .A2(n6719), .ZN(n6812) );
  NAND2_X1 U7845 ( .A1(n6813), .A2(n6812), .ZN(n8092) );
  NAND2_X1 U7846 ( .A1(n8090), .A2(n8092), .ZN(n6818) );
  INV_X1 U7847 ( .A(n6814), .ZN(n6817) );
  INV_X1 U7848 ( .A(n6815), .ZN(n6816) );
  NAND2_X1 U7849 ( .A1(n6817), .A2(n6816), .ZN(n8089) );
  NAND2_X1 U7850 ( .A1(n7205), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6823) );
  INV_X1 U7851 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7239) );
  OR2_X1 U7852 ( .A1(n6761), .A2(n7239), .ZN(n6822) );
  OAI21_X1 U7853 ( .B1(n6819), .B2(P1_REG3_REG_6__SCAN_IN), .A(n6834), .ZN(
        n8102) );
  OR2_X1 U7854 ( .A1(n6781), .A2(n8102), .ZN(n6821) );
  INV_X1 U7855 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7997) );
  OR2_X1 U7856 ( .A1(n8942), .A2(n7997), .ZN(n6820) );
  NAND4_X1 U7857 ( .A1(n6823), .A2(n6822), .A3(n6821), .A4(n6820), .ZN(n10100)
         );
  NAND2_X1 U7858 ( .A1(n10100), .A2(n6719), .ZN(n6829) );
  NAND2_X1 U7859 ( .A1(n6824), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6825) );
  XNOR2_X1 U7860 ( .A(n6825), .B(P1_IR_REG_6__SCAN_IN), .ZN(n7281) );
  INV_X1 U7861 ( .A(n7281), .ZN(n7508) );
  INV_X1 U7862 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7336) );
  OR2_X1 U7863 ( .A1(n8949), .A2(n7336), .ZN(n6827) );
  OR2_X1 U7864 ( .A1(n6746), .A2(n7335), .ZN(n6826) );
  NAND2_X1 U7865 ( .A1(n8105), .A2(n9192), .ZN(n6828) );
  NAND2_X1 U7866 ( .A1(n6829), .A2(n6828), .ZN(n6830) );
  NAND2_X1 U7867 ( .A1(n10100), .A2(n9196), .ZN(n6832) );
  NAND2_X1 U7868 ( .A1(n8105), .A2(n6719), .ZN(n6831) );
  NAND2_X1 U7869 ( .A1(n6832), .A2(n6831), .ZN(n8100) );
  NAND2_X1 U7870 ( .A1(n7205), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6839) );
  INV_X1 U7871 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7248) );
  OR2_X1 U7872 ( .A1(n6761), .A2(n7248), .ZN(n6838) );
  AND2_X1 U7873 ( .A1(n6834), .A2(n6833), .ZN(n6835) );
  OR2_X1 U7874 ( .A1(n6835), .A2(n6855), .ZN(n8694) );
  OR2_X1 U7875 ( .A1(n6781), .A2(n8694), .ZN(n6837) );
  INV_X1 U7876 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n8127) );
  OR2_X1 U7877 ( .A1(n8942), .A2(n8127), .ZN(n6836) );
  NAND2_X1 U7878 ( .A1(n10099), .A2(n6719), .ZN(n6844) );
  OR2_X1 U7879 ( .A1(n6824), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n6852) );
  NAND2_X1 U7880 ( .A1(n6852), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6840) );
  XNOR2_X1 U7881 ( .A(n6840), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7542) );
  INV_X1 U7882 ( .A(n7542), .ZN(n7338) );
  OR2_X1 U7883 ( .A1(n7339), .A2(n6746), .ZN(n6842) );
  INV_X1 U7884 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7340) );
  OR2_X1 U7885 ( .A1(n8949), .A2(n7340), .ZN(n6841) );
  OAI211_X1 U7886 ( .C1(n7263), .C2(n7338), .A(n6842), .B(n6841), .ZN(n8697)
         );
  NAND2_X1 U7887 ( .A1(n8697), .A2(n9192), .ZN(n6843) );
  NAND2_X1 U7888 ( .A1(n6844), .A2(n6843), .ZN(n6845) );
  XNOR2_X1 U7889 ( .A(n6845), .B(n6752), .ZN(n6846) );
  AOI22_X1 U7890 ( .A1(n10099), .A2(n9196), .B1(n6719), .B2(n8697), .ZN(n6847)
         );
  NAND2_X1 U7891 ( .A1(n6846), .A2(n6847), .ZN(n8756) );
  INV_X1 U7892 ( .A(n6846), .ZN(n6849) );
  INV_X1 U7893 ( .A(n6847), .ZN(n6848) );
  NAND2_X1 U7894 ( .A1(n6849), .A2(n6848), .ZN(n6850) );
  NAND2_X1 U7895 ( .A1(n8756), .A2(n6850), .ZN(n8693) );
  INV_X1 U7896 ( .A(n6851), .ZN(n8757) );
  OR2_X1 U7897 ( .A1(n7348), .A2(n6746), .ZN(n6854) );
  NOR2_X1 U7898 ( .A1(n6852), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n6894) );
  OR2_X1 U7899 ( .A1(n6894), .A2(n6662), .ZN(n6866) );
  XNOR2_X1 U7900 ( .A(n6866), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7553) );
  AOI22_X1 U7901 ( .A1(n7029), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7028), .B2(
        n7553), .ZN(n6853) );
  NAND2_X1 U7902 ( .A1(n8637), .A2(n6719), .ZN(n6863) );
  NAND2_X1 U7903 ( .A1(n6898), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6861) );
  INV_X1 U7904 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7250) );
  OR2_X1 U7905 ( .A1(n6761), .A2(n7250), .ZN(n6860) );
  OR2_X1 U7906 ( .A1(n6855), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6856) );
  NAND2_X1 U7907 ( .A1(n6872), .A2(n6856), .ZN(n8764) );
  OR2_X1 U7908 ( .A1(n6781), .A2(n8764), .ZN(n6859) );
  INV_X1 U7909 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n6857) );
  OR2_X1 U7910 ( .A1(n8941), .A2(n6857), .ZN(n6858) );
  NAND4_X1 U7911 ( .A1(n6861), .A2(n6860), .A3(n6859), .A4(n6858), .ZN(n10098)
         );
  NAND2_X1 U7912 ( .A1(n10098), .A2(n9196), .ZN(n6862) );
  AND2_X1 U7913 ( .A1(n6863), .A2(n6862), .ZN(n8758) );
  INV_X1 U7914 ( .A(n8758), .ZN(n6864) );
  AND2_X1 U7915 ( .A1(n8756), .A2(n6864), .ZN(n6865) );
  NAND2_X1 U7916 ( .A1(n7357), .A2(n8947), .ZN(n6870) );
  INV_X1 U7917 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8567) );
  NAND2_X1 U7918 ( .A1(n6866), .A2(n8567), .ZN(n6867) );
  NAND2_X1 U7919 ( .A1(n6867), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6868) );
  XNOR2_X1 U7920 ( .A(n6868), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7567) );
  AOI22_X1 U7921 ( .A1(n7029), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7028), .B2(
        n7567), .ZN(n6869) );
  NAND2_X1 U7922 ( .A1(n8790), .A2(n9192), .ZN(n6879) );
  NAND2_X1 U7923 ( .A1(n7205), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6877) );
  INV_X1 U7924 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7253) );
  OR2_X1 U7925 ( .A1(n6761), .A2(n7253), .ZN(n6876) );
  NAND2_X1 U7926 ( .A1(n6872), .A2(n6871), .ZN(n6873) );
  NAND2_X1 U7927 ( .A1(n6899), .A2(n6873), .ZN(n10008) );
  OR2_X1 U7928 ( .A1(n6781), .A2(n10008), .ZN(n6875) );
  INV_X1 U7929 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n8642) );
  OR2_X1 U7930 ( .A1(n8942), .A2(n8642), .ZN(n6874) );
  NAND4_X1 U7931 ( .A1(n6877), .A2(n6876), .A3(n6875), .A4(n6874), .ZN(n10097)
         );
  NAND2_X1 U7932 ( .A1(n10097), .A2(n6719), .ZN(n6878) );
  NAND2_X1 U7933 ( .A1(n6879), .A2(n6878), .ZN(n6880) );
  XNOR2_X1 U7934 ( .A(n6880), .B(n6752), .ZN(n6882) );
  AND2_X1 U7935 ( .A1(n10097), .A2(n9196), .ZN(n6881) );
  AOI21_X1 U7936 ( .B1(n8790), .B2(n6719), .A(n6881), .ZN(n6883) );
  NAND2_X1 U7937 ( .A1(n6882), .A2(n6883), .ZN(n6892) );
  INV_X1 U7938 ( .A(n6882), .ZN(n6885) );
  INV_X1 U7939 ( .A(n6883), .ZN(n6884) );
  NAND2_X1 U7940 ( .A1(n6885), .A2(n6884), .ZN(n6886) );
  AND2_X1 U7941 ( .A1(n6892), .A2(n6886), .ZN(n10006) );
  NAND2_X1 U7942 ( .A1(n8637), .A2(n9192), .ZN(n6888) );
  NAND2_X1 U7943 ( .A1(n10098), .A2(n6719), .ZN(n6887) );
  NAND2_X1 U7944 ( .A1(n6888), .A2(n6887), .ZN(n6889) );
  XNOR2_X1 U7945 ( .A(n6889), .B(n7154), .ZN(n8761) );
  AND2_X1 U7946 ( .A1(n8756), .A2(n8761), .ZN(n6890) );
  INV_X1 U7947 ( .A(n8761), .ZN(n6891) );
  NAND2_X1 U7948 ( .A1(n10004), .A2(n6892), .ZN(n6911) );
  NAND2_X1 U7949 ( .A1(n7398), .A2(n8947), .ZN(n6897) );
  NOR2_X1 U7950 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n6893) );
  NAND2_X1 U7951 ( .A1(n6894), .A2(n6893), .ZN(n6914) );
  NAND2_X1 U7952 ( .A1(n6914), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6895) );
  XNOR2_X1 U7953 ( .A(n6895), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7283) );
  AOI22_X1 U7954 ( .A1(n7029), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7028), .B2(
        n7283), .ZN(n6896) );
  NAND2_X1 U7955 ( .A1(n8868), .A2(n9192), .ZN(n6907) );
  NAND2_X1 U7956 ( .A1(n6898), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6905) );
  INV_X1 U7957 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7254) );
  OR2_X1 U7958 ( .A1(n6761), .A2(n7254), .ZN(n6904) );
  NAND2_X1 U7959 ( .A1(n6899), .A2(n7315), .ZN(n6900) );
  NAND2_X1 U7960 ( .A1(n6920), .A2(n6900), .ZN(n8880) );
  OR2_X1 U7961 ( .A1(n6781), .A2(n8880), .ZN(n6903) );
  INV_X1 U7962 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n6901) );
  OR2_X1 U7963 ( .A1(n8941), .A2(n6901), .ZN(n6902) );
  NAND4_X1 U7964 ( .A1(n6905), .A2(n6904), .A3(n6903), .A4(n6902), .ZN(n10096)
         );
  NAND2_X1 U7965 ( .A1(n10096), .A2(n6719), .ZN(n6906) );
  NAND2_X1 U7966 ( .A1(n6907), .A2(n6906), .ZN(n6908) );
  XNOR2_X1 U7967 ( .A(n6908), .B(n6752), .ZN(n6912) );
  NAND2_X1 U7968 ( .A1(n8868), .A2(n6719), .ZN(n6910) );
  NAND2_X1 U7969 ( .A1(n10096), .A2(n9196), .ZN(n6909) );
  NAND2_X1 U7970 ( .A1(n6910), .A2(n6909), .ZN(n8877) );
  INV_X1 U7971 ( .A(n6912), .ZN(n6913) );
  OR2_X1 U7972 ( .A1(n7401), .A2(n6746), .ZN(n6918) );
  OR2_X1 U7973 ( .A1(n6914), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6935) );
  NAND2_X1 U7974 ( .A1(n6935), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6916) );
  INV_X1 U7975 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6915) );
  XNOR2_X1 U7976 ( .A(n6916), .B(n6915), .ZN(n7629) );
  INV_X1 U7977 ( .A(n7629), .ZN(n7636) );
  AOI22_X1 U7978 ( .A1(n7029), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7028), .B2(
        n7636), .ZN(n6917) );
  NAND2_X1 U7979 ( .A1(n8962), .A2(n9192), .ZN(n6927) );
  NAND2_X1 U7980 ( .A1(n7205), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6925) );
  INV_X1 U7981 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7255) );
  OR2_X1 U7982 ( .A1(n6761), .A2(n7255), .ZN(n6924) );
  AND2_X1 U7983 ( .A1(n6920), .A2(n6919), .ZN(n6921) );
  OR2_X1 U7984 ( .A1(n6921), .A2(n6938), .ZN(n10908) );
  OR2_X1 U7985 ( .A1(n6781), .A2(n10908), .ZN(n6923) );
  INV_X1 U7986 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10909) );
  OR2_X1 U7987 ( .A1(n8942), .A2(n10909), .ZN(n6922) );
  NAND4_X1 U7988 ( .A1(n6925), .A2(n6924), .A3(n6923), .A4(n6922), .ZN(n10095)
         );
  NAND2_X1 U7989 ( .A1(n10095), .A2(n6719), .ZN(n6926) );
  NAND2_X1 U7990 ( .A1(n6927), .A2(n6926), .ZN(n6928) );
  XNOR2_X1 U7991 ( .A(n6928), .B(n6752), .ZN(n6930) );
  AND2_X1 U7992 ( .A1(n10095), .A2(n9196), .ZN(n6929) );
  AOI21_X1 U7993 ( .B1(n8962), .B2(n6719), .A(n6929), .ZN(n6931) );
  NAND2_X1 U7994 ( .A1(n6930), .A2(n6931), .ZN(n8886) );
  INV_X1 U7995 ( .A(n6930), .ZN(n6933) );
  INV_X1 U7996 ( .A(n6931), .ZN(n6932) );
  NAND2_X1 U7997 ( .A1(n6933), .A2(n6932), .ZN(n8887) );
  NAND2_X1 U7998 ( .A1(n6934), .A2(n8887), .ZN(n8906) );
  OAI21_X1 U7999 ( .B1(n6935), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6951) );
  INV_X1 U8000 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8571) );
  XNOR2_X1 U8001 ( .A(n6951), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7763) );
  AOI22_X1 U8002 ( .A1(n7029), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7028), .B2(
        n7763), .ZN(n6936) );
  NAND2_X1 U8003 ( .A1(n9210), .A2(n9192), .ZN(n6945) );
  NAND2_X1 U8004 ( .A1(n7205), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6943) );
  INV_X1 U8005 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7238) );
  OR2_X1 U8006 ( .A1(n6761), .A2(n7238), .ZN(n6942) );
  OR2_X1 U8007 ( .A1(n6938), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6939) );
  NAND2_X1 U8008 ( .A1(n6957), .A2(n6939), .ZN(n8910) );
  OR2_X1 U8009 ( .A1(n6781), .A2(n8910), .ZN(n6941) );
  INV_X1 U8010 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n8836) );
  OR2_X1 U8011 ( .A1(n8942), .A2(n8836), .ZN(n6940) );
  NAND4_X1 U8012 ( .A1(n6943), .A2(n6942), .A3(n6941), .A4(n6940), .ZN(n10094)
         );
  NAND2_X1 U8013 ( .A1(n10094), .A2(n6719), .ZN(n6944) );
  NAND2_X1 U8014 ( .A1(n6945), .A2(n6944), .ZN(n6946) );
  XNOR2_X1 U8015 ( .A(n6946), .B(n6752), .ZN(n8908) );
  AND2_X1 U8016 ( .A1(n10094), .A2(n9196), .ZN(n6947) );
  AOI21_X1 U8017 ( .B1(n9210), .B2(n6719), .A(n6947), .ZN(n6948) );
  INV_X1 U8018 ( .A(n8908), .ZN(n6949) );
  INV_X1 U8019 ( .A(n6948), .ZN(n8907) );
  NAND2_X1 U8020 ( .A1(n6949), .A2(n8907), .ZN(n6950) );
  NAND2_X1 U8021 ( .A1(n7558), .A2(n8947), .ZN(n6955) );
  NAND2_X1 U8022 ( .A1(n6951), .A2(n8571), .ZN(n6952) );
  NAND2_X1 U8023 ( .A1(n6952), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6953) );
  XNOR2_X1 U8024 ( .A(n6953), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7913) );
  AOI22_X1 U8025 ( .A1(n7029), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7028), .B2(
        n7913), .ZN(n6954) );
  NAND2_X1 U8026 ( .A1(n10433), .A2(n9192), .ZN(n6964) );
  NAND2_X1 U8027 ( .A1(n7205), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6962) );
  INV_X1 U8028 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7237) );
  OR2_X1 U8029 ( .A1(n6761), .A2(n7237), .ZN(n6961) );
  INV_X1 U8030 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7288) );
  OR2_X1 U8031 ( .A1(n8942), .A2(n7288), .ZN(n6960) );
  NAND2_X1 U8032 ( .A1(n6957), .A2(n6956), .ZN(n6958) );
  NAND2_X1 U8033 ( .A1(n6977), .A2(n6958), .ZN(n10430) );
  OR2_X1 U8034 ( .A1(n6781), .A2(n10430), .ZN(n6959) );
  NAND4_X1 U8035 ( .A1(n6962), .A2(n6961), .A3(n6960), .A4(n6959), .ZN(n10404)
         );
  NAND2_X1 U8036 ( .A1(n10404), .A2(n6719), .ZN(n6963) );
  NAND2_X1 U8037 ( .A1(n6964), .A2(n6963), .ZN(n6965) );
  XNOR2_X1 U8038 ( .A(n6965), .B(n7154), .ZN(n6968) );
  NAND2_X1 U8039 ( .A1(n10433), .A2(n6719), .ZN(n6967) );
  NAND2_X1 U8040 ( .A1(n10404), .A2(n9196), .ZN(n6966) );
  NAND2_X1 U8041 ( .A1(n6967), .A2(n6966), .ZN(n6969) );
  INV_X1 U8042 ( .A(n6968), .ZN(n6971) );
  INV_X1 U8043 ( .A(n6969), .ZN(n6970) );
  NAND2_X1 U8044 ( .A1(n6971), .A2(n6970), .ZN(n10023) );
  NAND2_X1 U8045 ( .A1(n6972), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6973) );
  XNOR2_X1 U8046 ( .A(n6973), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7289) );
  AOI22_X1 U8047 ( .A1(n7029), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7028), .B2(
        n7289), .ZN(n6974) );
  NAND2_X1 U8048 ( .A1(n10413), .A2(n9192), .ZN(n6985) );
  NAND2_X1 U8049 ( .A1(n7205), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6983) );
  INV_X1 U8050 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6976) );
  OR2_X1 U8051 ( .A1(n6761), .A2(n6976), .ZN(n6982) );
  INV_X1 U8052 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10407) );
  OR2_X1 U8053 ( .A1(n8942), .A2(n10407), .ZN(n6981) );
  AND2_X1 U8054 ( .A1(n6977), .A2(n7973), .ZN(n6979) );
  OR2_X1 U8055 ( .A1(n6979), .A2(n6978), .ZN(n10406) );
  OR2_X1 U8056 ( .A1(n6781), .A2(n10406), .ZN(n6980) );
  NAND4_X1 U8057 ( .A1(n6983), .A2(n6982), .A3(n6981), .A4(n6980), .ZN(n10093)
         );
  NAND2_X1 U8058 ( .A1(n10093), .A2(n6719), .ZN(n6984) );
  NAND2_X1 U8059 ( .A1(n6985), .A2(n6984), .ZN(n6986) );
  XNOR2_X1 U8060 ( .A(n6986), .B(n6752), .ZN(n6989) );
  NAND2_X1 U8061 ( .A1(n6990), .A2(n6989), .ZN(n9927) );
  NAND2_X1 U8062 ( .A1(n10413), .A2(n6719), .ZN(n6988) );
  NAND2_X1 U8063 ( .A1(n10093), .A2(n9196), .ZN(n6987) );
  NAND2_X1 U8064 ( .A1(n6988), .A2(n6987), .ZN(n9929) );
  NAND2_X1 U8065 ( .A1(n9927), .A2(n9929), .ZN(n6991) );
  OAI22_X1 U8066 ( .A1(n9982), .A2(n6995), .B1(n10073), .B2(n9978), .ZN(n6992)
         );
  OR2_X1 U8067 ( .A1(n6996), .A2(n6662), .ZN(n7009) );
  XNOR2_X1 U8068 ( .A(n7009), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10136) );
  AOI22_X1 U8069 ( .A1(n7029), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7028), .B2(
        n10136), .ZN(n6997) );
  NAND2_X1 U8070 ( .A1(n7205), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n7003) );
  INV_X1 U8071 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n7235) );
  OR2_X1 U8072 ( .A1(n6761), .A2(n7235), .ZN(n7002) );
  XNOR2_X1 U8073 ( .A(P1_REG3_REG_17__SCAN_IN), .B(n7014), .ZN(n10350) );
  OR2_X1 U8074 ( .A1(n6781), .A2(n10350), .ZN(n7001) );
  INV_X1 U8075 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10351) );
  OR2_X1 U8076 ( .A1(n8942), .A2(n10351), .ZN(n7000) );
  NAND4_X1 U8077 ( .A1(n7003), .A2(n7002), .A3(n7001), .A4(n7000), .ZN(n10332)
         );
  AOI22_X1 U8078 ( .A1(n10356), .A2(n6719), .B1(n9196), .B2(n10332), .ZN(n7007) );
  NAND2_X1 U8079 ( .A1(n10356), .A2(n9192), .ZN(n7005) );
  NAND2_X1 U8080 ( .A1(n10332), .A2(n6719), .ZN(n7004) );
  NAND2_X1 U8081 ( .A1(n7005), .A2(n7004), .ZN(n7006) );
  XNOR2_X1 U8082 ( .A(n7006), .B(n7154), .ZN(n7008) );
  XOR2_X1 U8083 ( .A(n7007), .B(n7008), .Z(n9990) );
  INV_X1 U8084 ( .A(n10055), .ZN(n7024) );
  INV_X1 U8085 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8364) );
  NAND2_X1 U8086 ( .A1(n7009), .A2(n8364), .ZN(n7010) );
  NAND2_X1 U8087 ( .A1(n7010), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7011) );
  XNOR2_X1 U8088 ( .A(n7011), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10146) );
  AOI22_X1 U8089 ( .A1(n7029), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7028), .B2(
        n10146), .ZN(n7012) );
  AOI21_X1 U8090 ( .B1(P1_REG3_REG_17__SCAN_IN), .B2(n7014), .A(
        P1_REG3_REG_18__SCAN_IN), .ZN(n7015) );
  NOR2_X1 U8091 ( .A1(n7015), .A2(n7032), .ZN(n10337) );
  NAND2_X1 U8092 ( .A1(n7016), .A2(n10337), .ZN(n7022) );
  INV_X1 U8093 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10134) );
  OR2_X1 U8094 ( .A1(n6761), .A2(n10134), .ZN(n7021) );
  INV_X1 U8095 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n7017) );
  OR2_X1 U8096 ( .A1(n8941), .A2(n7017), .ZN(n7020) );
  INV_X1 U8097 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n7018) );
  OR2_X1 U8098 ( .A1(n8942), .A2(n7018), .ZN(n7019) );
  NAND4_X1 U8099 ( .A1(n7022), .A2(n7021), .A3(n7020), .A4(n7019), .ZN(n10348)
         );
  AOI22_X1 U8100 ( .A1(n10506), .A2(n9192), .B1(n6719), .B2(n10348), .ZN(n7023) );
  XOR2_X1 U8101 ( .A(n7154), .B(n7023), .Z(n7025) );
  NAND2_X1 U8102 ( .A1(n7024), .A2(n7025), .ZN(n7027) );
  AOI22_X1 U8103 ( .A1(n10506), .A2(n6719), .B1(n9196), .B2(n10348), .ZN(
        n10052) );
  INV_X1 U8104 ( .A(n7025), .ZN(n10053) );
  NAND2_X1 U8105 ( .A1(n7916), .A2(n8947), .ZN(n7031) );
  AOI22_X1 U8106 ( .A1(n7029), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5073), .B2(
        n7028), .ZN(n7030) );
  NAND2_X1 U8107 ( .A1(n10503), .A2(n9192), .ZN(n7042) );
  NAND2_X1 U8108 ( .A1(n7205), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n7040) );
  INV_X1 U8109 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10147) );
  OR2_X1 U8110 ( .A1(n6761), .A2(n10147), .ZN(n7039) );
  INV_X1 U8111 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n10321) );
  OR2_X1 U8112 ( .A1(n8942), .A2(n10321), .ZN(n7038) );
  INV_X1 U8113 ( .A(n7051), .ZN(n7036) );
  INV_X1 U8114 ( .A(n7032), .ZN(n7034) );
  INV_X1 U8115 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n7033) );
  NAND2_X1 U8116 ( .A1(n7034), .A2(n7033), .ZN(n7035) );
  NAND2_X1 U8117 ( .A1(n7036), .A2(n7035), .ZN(n10320) );
  OR2_X1 U8118 ( .A1(n6781), .A2(n10320), .ZN(n7037) );
  NAND4_X1 U8119 ( .A1(n7040), .A2(n7039), .A3(n7038), .A4(n7037), .ZN(n10331)
         );
  NAND2_X1 U8120 ( .A1(n10331), .A2(n6719), .ZN(n7041) );
  NAND2_X1 U8121 ( .A1(n7042), .A2(n7041), .ZN(n7043) );
  XNOR2_X1 U8122 ( .A(n7043), .B(n6752), .ZN(n9949) );
  AND2_X1 U8123 ( .A1(n10331), .A2(n9196), .ZN(n7044) );
  AOI21_X1 U8124 ( .B1(n10503), .B2(n6719), .A(n7044), .ZN(n7045) );
  NAND2_X1 U8125 ( .A1(n9949), .A2(n7045), .ZN(n7047) );
  INV_X1 U8126 ( .A(n9949), .ZN(n7046) );
  INV_X1 U8127 ( .A(n7045), .ZN(n9948) );
  NAND2_X1 U8128 ( .A1(n8067), .A2(n8947), .ZN(n7049) );
  INV_X1 U8129 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8086) );
  OR2_X1 U8130 ( .A1(n8949), .A2(n8086), .ZN(n7048) );
  NAND2_X1 U8131 ( .A1(n10306), .A2(n9192), .ZN(n7057) );
  NAND2_X1 U8132 ( .A1(n6706), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n7055) );
  INV_X1 U8133 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n7050) );
  OR2_X1 U8134 ( .A1(n8941), .A2(n7050), .ZN(n7054) );
  NAND2_X1 U8135 ( .A1(n7051), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n7066) );
  OAI21_X1 U8136 ( .B1(n7051), .B2(P1_REG3_REG_20__SCAN_IN), .A(n7066), .ZN(
        n10303) );
  OR2_X1 U8137 ( .A1(n6781), .A2(n10303), .ZN(n7053) );
  INV_X1 U8138 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n10304) );
  OR2_X1 U8139 ( .A1(n8942), .A2(n10304), .ZN(n7052) );
  NAND4_X1 U8140 ( .A1(n7055), .A2(n7054), .A3(n7053), .A4(n7052), .ZN(n10283)
         );
  NAND2_X1 U8141 ( .A1(n10283), .A2(n6719), .ZN(n7056) );
  NAND2_X1 U8142 ( .A1(n7057), .A2(n7056), .ZN(n7058) );
  XNOR2_X1 U8143 ( .A(n7058), .B(n6752), .ZN(n7060) );
  AND2_X1 U8144 ( .A1(n10283), .A2(n9196), .ZN(n7059) );
  AOI21_X1 U8145 ( .B1(n10306), .B2(n6719), .A(n7059), .ZN(n7061) );
  INV_X1 U8146 ( .A(n7060), .ZN(n7063) );
  INV_X1 U8147 ( .A(n7061), .ZN(n7062) );
  NAND2_X1 U8148 ( .A1(n7063), .A2(n7062), .ZN(n10014) );
  INV_X1 U8149 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8069) );
  OR2_X1 U8150 ( .A1(n8949), .A2(n8069), .ZN(n7064) );
  NAND2_X1 U8151 ( .A1(n6706), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n7073) );
  INV_X1 U8152 ( .A(n7066), .ZN(n7067) );
  NAND2_X1 U8153 ( .A1(n7067), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n7079) );
  OAI21_X1 U8154 ( .B1(n7067), .B2(P1_REG3_REG_21__SCAN_IN), .A(n7079), .ZN(
        n10291) );
  OR2_X1 U8155 ( .A1(n6781), .A2(n10291), .ZN(n7072) );
  INV_X1 U8156 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n7068) );
  OR2_X1 U8157 ( .A1(n8942), .A2(n7068), .ZN(n7071) );
  INV_X1 U8158 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n7069) );
  OR2_X1 U8159 ( .A1(n8941), .A2(n7069), .ZN(n7070) );
  NAND4_X1 U8160 ( .A1(n7073), .A2(n7072), .A3(n7071), .A4(n7070), .ZN(n10092)
         );
  AOI22_X1 U8161 ( .A1(n10490), .A2(n9192), .B1(n6719), .B2(n10092), .ZN(n7074) );
  XNOR2_X1 U8162 ( .A(n7074), .B(n7154), .ZN(n7076) );
  AOI22_X1 U8163 ( .A1(n10490), .A2(n6719), .B1(n9196), .B2(n10092), .ZN(n7075) );
  NOR2_X1 U8164 ( .A1(n7076), .A2(n7075), .ZN(n9958) );
  NAND2_X1 U8165 ( .A1(n7076), .A2(n7075), .ZN(n9956) );
  INV_X1 U8166 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8629) );
  OR2_X1 U8167 ( .A1(n8949), .A2(n8629), .ZN(n7077) );
  NAND2_X1 U8168 ( .A1(n10486), .A2(n9192), .ZN(n7087) );
  NAND2_X1 U8169 ( .A1(n6706), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n7085) );
  INV_X1 U8170 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n10272) );
  OR2_X1 U8171 ( .A1(n8942), .A2(n10272), .ZN(n7084) );
  INV_X1 U8172 ( .A(n7079), .ZN(n7080) );
  NAND2_X1 U8173 ( .A1(n7080), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n7096) );
  OAI21_X1 U8174 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n7080), .A(n7096), .ZN(
        n10271) );
  OR2_X1 U8175 ( .A1(n6781), .A2(n10271), .ZN(n7083) );
  INV_X1 U8176 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n7081) );
  OR2_X1 U8177 ( .A1(n8941), .A2(n7081), .ZN(n7082) );
  NAND4_X1 U8178 ( .A1(n7085), .A2(n7084), .A3(n7083), .A4(n7082), .ZN(n10284)
         );
  NAND2_X1 U8179 ( .A1(n10284), .A2(n6719), .ZN(n7086) );
  NAND2_X1 U8180 ( .A1(n7087), .A2(n7086), .ZN(n7088) );
  XNOR2_X1 U8181 ( .A(n7088), .B(n7154), .ZN(n7092) );
  NAND2_X1 U8182 ( .A1(n10486), .A2(n6719), .ZN(n7090) );
  NAND2_X1 U8183 ( .A1(n10284), .A2(n9196), .ZN(n7089) );
  NAND2_X1 U8184 ( .A1(n7090), .A2(n7089), .ZN(n7091) );
  NAND2_X1 U8185 ( .A1(n7092), .A2(n7091), .ZN(n10035) );
  INV_X1 U8186 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8752) );
  OR2_X1 U8187 ( .A1(n8949), .A2(n8752), .ZN(n7093) );
  NAND2_X1 U8188 ( .A1(n7205), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n7102) );
  INV_X1 U8189 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n7095) );
  OR2_X1 U8190 ( .A1(n6761), .A2(n7095), .ZN(n7101) );
  INV_X1 U8191 ( .A(n7096), .ZN(n7097) );
  NAND2_X1 U8192 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(n7097), .ZN(n7111) );
  OAI21_X1 U8193 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n7097), .A(n7111), .ZN(
        n10254) );
  OR2_X1 U8194 ( .A1(n6781), .A2(n10254), .ZN(n7100) );
  INV_X1 U8195 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n7098) );
  OR2_X1 U8196 ( .A1(n8942), .A2(n7098), .ZN(n7099) );
  NAND4_X1 U8197 ( .A1(n7102), .A2(n7101), .A3(n7100), .A4(n7099), .ZN(n9225)
         );
  AOI22_X1 U8198 ( .A1(n10479), .A2(n9192), .B1(n6719), .B2(n9225), .ZN(n7103)
         );
  XOR2_X1 U8199 ( .A(n7154), .B(n7103), .Z(n7104) );
  AOI22_X1 U8200 ( .A1(n10479), .A2(n6719), .B1(n9196), .B2(n9225), .ZN(n9941)
         );
  INV_X1 U8201 ( .A(n7104), .ZN(n7105) );
  INV_X1 U8202 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8772) );
  OR2_X1 U8203 ( .A1(n8949), .A2(n8772), .ZN(n7107) );
  NAND2_X1 U8204 ( .A1(n7205), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n7117) );
  INV_X1 U8205 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n7109) );
  OR2_X1 U8206 ( .A1(n6761), .A2(n7109), .ZN(n7116) );
  INV_X1 U8207 ( .A(n7111), .ZN(n7110) );
  NAND2_X1 U8208 ( .A1(n7110), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n7128) );
  INV_X1 U8209 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9997) );
  NAND2_X1 U8210 ( .A1(n7111), .A2(n9997), .ZN(n7112) );
  NAND2_X1 U8211 ( .A1(n7128), .A2(n7112), .ZN(n10245) );
  OR2_X1 U8212 ( .A1(n6781), .A2(n10245), .ZN(n7115) );
  INV_X1 U8213 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n7113) );
  OR2_X1 U8214 ( .A1(n8942), .A2(n7113), .ZN(n7114) );
  NAND4_X1 U8215 ( .A1(n7117), .A2(n7116), .A3(n7115), .A4(n7114), .ZN(n10260)
         );
  AOI22_X1 U8216 ( .A1(n10476), .A2(n6719), .B1(n9196), .B2(n10260), .ZN(n7121) );
  NAND2_X1 U8217 ( .A1(n10476), .A2(n9192), .ZN(n7119) );
  NAND2_X1 U8218 ( .A1(n10260), .A2(n6719), .ZN(n7118) );
  NAND2_X1 U8219 ( .A1(n7119), .A2(n7118), .ZN(n7120) );
  XOR2_X1 U8220 ( .A(n7121), .B(n7123), .Z(n9996) );
  INV_X1 U8221 ( .A(n7121), .ZN(n7122) );
  INV_X1 U8222 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8846) );
  OR2_X1 U8223 ( .A1(n8949), .A2(n8846), .ZN(n7124) );
  NAND2_X1 U8224 ( .A1(n10470), .A2(n9192), .ZN(n7136) );
  NAND2_X1 U8225 ( .A1(n7205), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n7134) );
  INV_X1 U8226 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n7126) );
  OR2_X1 U8227 ( .A1(n6761), .A2(n7126), .ZN(n7133) );
  INV_X1 U8228 ( .A(n7128), .ZN(n7127) );
  NAND2_X1 U8229 ( .A1(n7127), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n7145) );
  INV_X1 U8230 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9970) );
  NAND2_X1 U8231 ( .A1(n7128), .A2(n9970), .ZN(n7129) );
  NAND2_X1 U8232 ( .A1(n7145), .A2(n7129), .ZN(n10220) );
  OR2_X1 U8233 ( .A1(n6781), .A2(n10220), .ZN(n7132) );
  INV_X1 U8234 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n7130) );
  OR2_X1 U8235 ( .A1(n8942), .A2(n7130), .ZN(n7131) );
  NAND4_X1 U8236 ( .A1(n7134), .A2(n7133), .A3(n7132), .A4(n7131), .ZN(n10091)
         );
  NAND2_X1 U8237 ( .A1(n10091), .A2(n6719), .ZN(n7135) );
  NAND2_X1 U8238 ( .A1(n7136), .A2(n7135), .ZN(n7137) );
  NAND2_X1 U8239 ( .A1(n10470), .A2(n6719), .ZN(n7139) );
  NAND2_X1 U8240 ( .A1(n10091), .A2(n9196), .ZN(n7138) );
  NOR2_X1 U8241 ( .A1(n9968), .A2(n9967), .ZN(n7140) );
  INV_X1 U8242 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10547) );
  OR2_X1 U8243 ( .A1(n8949), .A2(n10547), .ZN(n7141) );
  NAND2_X1 U8244 ( .A1(n10464), .A2(n9192), .ZN(n7153) );
  NAND2_X1 U8245 ( .A1(n7205), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n7151) );
  INV_X1 U8246 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n7143) );
  OR2_X1 U8247 ( .A1(n6761), .A2(n7143), .ZN(n7150) );
  INV_X1 U8248 ( .A(n7145), .ZN(n7144) );
  NAND2_X1 U8249 ( .A1(n7144), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n7209) );
  INV_X1 U8250 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n10064) );
  NAND2_X1 U8251 ( .A1(n7145), .A2(n10064), .ZN(n7146) );
  NAND2_X1 U8252 ( .A1(n7209), .A2(n7146), .ZN(n10211) );
  OR2_X1 U8253 ( .A1(n6781), .A2(n10211), .ZN(n7149) );
  INV_X1 U8254 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n7147) );
  OR2_X1 U8255 ( .A1(n8942), .A2(n7147), .ZN(n7148) );
  NAND4_X1 U8256 ( .A1(n7151), .A2(n7150), .A3(n7149), .A4(n7148), .ZN(n10228)
         );
  NAND2_X1 U8257 ( .A1(n10228), .A2(n6719), .ZN(n7152) );
  NAND2_X1 U8258 ( .A1(n7153), .A2(n7152), .ZN(n7155) );
  XNOR2_X1 U8259 ( .A(n7155), .B(n7154), .ZN(n7158) );
  AOI22_X1 U8260 ( .A1(n10464), .A2(n6719), .B1(n9196), .B2(n10228), .ZN(n7156) );
  XNOR2_X1 U8261 ( .A(n7158), .B(n7156), .ZN(n10062) );
  NAND2_X1 U8262 ( .A1(n10063), .A2(n10062), .ZN(n7160) );
  INV_X1 U8263 ( .A(n7156), .ZN(n7157) );
  NAND2_X1 U8264 ( .A1(n7158), .A2(n7157), .ZN(n7159) );
  INV_X1 U8265 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10544) );
  OR2_X1 U8266 ( .A1(n8949), .A2(n10544), .ZN(n7161) );
  NAND2_X1 U8267 ( .A1(n10459), .A2(n9192), .ZN(n7170) );
  NAND2_X1 U8268 ( .A1(n6706), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n7168) );
  INV_X1 U8269 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n7163) );
  OR2_X1 U8270 ( .A1(n8941), .A2(n7163), .ZN(n7167) );
  INV_X1 U8271 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n7208) );
  XNOR2_X1 U8272 ( .A(n7209), .B(n7208), .ZN(n7217) );
  OR2_X1 U8273 ( .A1(n6781), .A2(n7217), .ZN(n7166) );
  INV_X1 U8274 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n7164) );
  OR2_X1 U8275 ( .A1(n8942), .A2(n7164), .ZN(n7165) );
  NAND4_X1 U8276 ( .A1(n7168), .A2(n7167), .A3(n7166), .A4(n7165), .ZN(n10174)
         );
  NAND2_X1 U8277 ( .A1(n10174), .A2(n6719), .ZN(n7169) );
  NAND2_X1 U8278 ( .A1(n7170), .A2(n7169), .ZN(n7171) );
  XNOR2_X1 U8279 ( .A(n7171), .B(n6752), .ZN(n7175) );
  AND2_X1 U8280 ( .A1(n10174), .A2(n9196), .ZN(n7172) );
  AOI21_X1 U8281 ( .B1(n10459), .B2(n6719), .A(n7172), .ZN(n7174) );
  NAND2_X1 U8282 ( .A1(n7175), .A2(n7174), .ZN(n9202) );
  OAI21_X1 U8283 ( .B1(n7175), .B2(n7174), .A(n9202), .ZN(n7176) );
  NAND2_X1 U8284 ( .A1(n7177), .A2(n7176), .ZN(n7178) );
  INV_X1 U8285 ( .A(n10549), .ZN(n7182) );
  NAND2_X1 U8286 ( .A1(n8848), .A2(P1_B_REG_SCAN_IN), .ZN(n7179) );
  MUX2_X1 U8287 ( .A(P1_B_REG_SCAN_IN), .B(n7179), .S(n8774), .Z(n7180) );
  NAND2_X1 U8288 ( .A1(n7182), .A2(n7180), .ZN(n7194) );
  INV_X1 U8289 ( .A(n8848), .ZN(n7181) );
  OAI22_X1 U8290 ( .A1(n7194), .A2(P1_D_REG_1__SCAN_IN), .B1(n7182), .B2(n7181), .ZN(n7647) );
  NOR4_X1 U8291 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n7186) );
  NOR4_X1 U8292 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n7185) );
  NOR4_X1 U8293 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n7184) );
  NOR4_X1 U8294 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n7183) );
  NAND4_X1 U8295 ( .A1(n7186), .A2(n7185), .A3(n7184), .A4(n7183), .ZN(n7192)
         );
  NOR2_X1 U8296 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .ZN(
        n7190) );
  NOR4_X1 U8297 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_30__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n7189) );
  NOR4_X1 U8298 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n7188) );
  NOR4_X1 U8299 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n7187) );
  NAND4_X1 U8300 ( .A1(n7190), .A2(n7189), .A3(n7188), .A4(n7187), .ZN(n7191)
         );
  NOR2_X1 U8301 ( .A1(n7192), .A2(n7191), .ZN(n7193) );
  NOR2_X1 U8302 ( .A1(n7194), .A2(n7193), .ZN(n7651) );
  OR2_X1 U8303 ( .A1(n7647), .A2(n7651), .ZN(n7687) );
  INV_X1 U8304 ( .A(n7194), .ZN(n10551) );
  INV_X1 U8305 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n8608) );
  NAND2_X1 U8306 ( .A1(n10551), .A2(n8608), .ZN(n7196) );
  NAND2_X1 U8307 ( .A1(n10549), .A2(n8774), .ZN(n7195) );
  NAND2_X1 U8308 ( .A1(n7196), .A2(n7195), .ZN(n7689) );
  NOR2_X1 U8309 ( .A1(n7687), .A2(n7689), .ZN(n7580) );
  NAND2_X1 U8310 ( .A1(n5187), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7197) );
  XNOR2_X1 U8311 ( .A(n7197), .B(n8591), .ZN(n8750) );
  AND2_X1 U8312 ( .A1(n8750), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7230) );
  NAND2_X1 U8313 ( .A1(n7300), .A2(n7230), .ZN(n10623) );
  INV_X1 U8314 ( .A(n10623), .ZN(n10531) );
  INV_X1 U8315 ( .A(n9169), .ZN(n9172) );
  NAND2_X1 U8316 ( .A1(n8630), .A2(n9172), .ZN(n7799) );
  AND2_X1 U8317 ( .A1(n11015), .A2(n8929), .ZN(n7220) );
  NAND2_X1 U8318 ( .A1(n7200), .A2(n7220), .ZN(n10071) );
  NAND2_X1 U8319 ( .A1(n7198), .A2(n10078), .ZN(n7229) );
  INV_X1 U8320 ( .A(n7799), .ZN(n7654) );
  AND2_X1 U8321 ( .A1(n7654), .A2(n9167), .ZN(n10791) );
  NAND2_X1 U8322 ( .A1(n7200), .A2(n10791), .ZN(n7199) );
  OR2_X1 U8323 ( .A1(n10737), .A2(n9169), .ZN(n7649) );
  OR2_X2 U8324 ( .A1(n10623), .A2(n7649), .ZN(n10907) );
  INV_X1 U8325 ( .A(n7200), .ZN(n7201) );
  NOR2_X1 U8326 ( .A1(n7201), .A2(n9186), .ZN(n7204) );
  INV_X1 U8327 ( .A(n7202), .ZN(n7670) );
  INV_X1 U8328 ( .A(n8929), .ZN(n7203) );
  AOI22_X1 U8329 ( .A1(n10081), .A2(n10228), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3084), .ZN(n7226) );
  AND2_X1 U8330 ( .A1(n7202), .A2(n7203), .ZN(n10398) );
  NAND2_X1 U8331 ( .A1(n7205), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7216) );
  INV_X1 U8332 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7206) );
  OR2_X1 U8333 ( .A1(n6761), .A2(n7206), .ZN(n7215) );
  INV_X1 U8334 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7207) );
  OAI21_X1 U8335 ( .B1(n7209), .B2(n7208), .A(n7207), .ZN(n7212) );
  INV_X1 U8336 ( .A(n7209), .ZN(n7211) );
  AND2_X1 U8337 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .ZN(n7210) );
  NAND2_X1 U8338 ( .A1(n7211), .A2(n7210), .ZN(n9265) );
  NAND2_X1 U8339 ( .A1(n7212), .A2(n9265), .ZN(n10178) );
  OR2_X1 U8340 ( .A1(n6781), .A2(n10178), .ZN(n7214) );
  INV_X1 U8341 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n10179) );
  OR2_X1 U8342 ( .A1(n8942), .A2(n10179), .ZN(n7213) );
  NAND4_X1 U8343 ( .A1(n7216), .A2(n7215), .A3(n7214), .A4(n7213), .ZN(n10197)
         );
  INV_X1 U8344 ( .A(n7217), .ZN(n10191) );
  INV_X1 U8345 ( .A(n7580), .ZN(n7223) );
  OR2_X1 U8346 ( .A1(n8929), .A2(n7218), .ZN(n7648) );
  NAND3_X1 U8347 ( .A1(n7300), .A2(n8750), .A3(n7648), .ZN(n7219) );
  AOI21_X1 U8348 ( .B1(n7223), .B2(n7220), .A(n7219), .ZN(n7221) );
  OR2_X1 U8349 ( .A1(n7221), .A2(P1_U3084), .ZN(n7224) );
  INV_X1 U8350 ( .A(n7222), .ZN(n7655) );
  OAI211_X1 U8351 ( .C1(n7655), .C2(n10791), .A(n7223), .B(n10531), .ZN(n7579)
         );
  NAND2_X1 U8352 ( .A1(n7224), .A2(n7579), .ZN(n9930) );
  AOI22_X1 U8353 ( .A1(n10086), .A2(n10197), .B1(n10191), .B2(n9930), .ZN(
        n7225) );
  OAI211_X1 U8354 ( .C1(n10193), .C2(n10089), .A(n7226), .B(n7225), .ZN(n7227)
         );
  INV_X1 U8355 ( .A(n7227), .ZN(n7228) );
  NAND2_X1 U8356 ( .A1(n7229), .A2(n7228), .ZN(P1_U3212) );
  INV_X1 U8357 ( .A(n7230), .ZN(n7231) );
  NOR2_X1 U8358 ( .A1(n7300), .A2(n7231), .ZN(P1_U4006) );
  INV_X1 U8359 ( .A(n7355), .ZN(n7232) );
  OR2_X2 U8360 ( .A1(n7371), .A2(n7232), .ZN(n9406) );
  INV_X1 U8361 ( .A(n9406), .ZN(P2_U3966) );
  NAND2_X1 U8362 ( .A1(n7300), .A2(n8929), .ZN(n7233) );
  NAND2_X1 U8363 ( .A1(n7233), .A2(n8750), .ZN(n7262) );
  NAND2_X1 U8364 ( .A1(n7262), .A2(n7263), .ZN(n7234) );
  NAND2_X1 U8365 ( .A1(n7234), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NOR2_X1 U8366 ( .A1(n10136), .A2(n7235), .ZN(n7236) );
  AOI21_X1 U8367 ( .B1(n10136), .B2(n7235), .A(n7236), .ZN(n7266) );
  INV_X1 U8368 ( .A(n7289), .ZN(n7972) );
  AOI22_X1 U8369 ( .A1(n7289), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n6976), .B2(
        n7972), .ZN(n7971) );
  MUX2_X1 U8370 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7237), .S(n7913), .Z(n7911)
         );
  OR2_X1 U8371 ( .A1(n7763), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7258) );
  MUX2_X1 U8372 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7238), .S(n7763), .Z(n7760)
         );
  NOR2_X1 U8373 ( .A1(n7255), .A2(n7629), .ZN(n7628) );
  INV_X1 U8374 ( .A(n7283), .ZN(n7402) );
  INV_X1 U8375 ( .A(n7567), .ZN(n7358) );
  OR2_X1 U8376 ( .A1(n7553), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7252) );
  NOR2_X1 U8377 ( .A1(n7542), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7249) );
  NAND2_X1 U8378 ( .A1(n7281), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7247) );
  MUX2_X1 U8379 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n7239), .S(n7281), .Z(n7504)
         );
  NAND2_X1 U8380 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n7280), .ZN(n7246) );
  MUX2_X1 U8381 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n7240), .S(n7280), .Z(n7528)
         );
  AOI22_X1 U8382 ( .A1(n7278), .A2(n6779), .B1(P1_REG1_REG_4__SCAN_IN), .B2(
        n7682), .ZN(n7680) );
  NAND2_X1 U8383 ( .A1(P1_REG1_REG_3__SCAN_IN), .A2(n7277), .ZN(n7244) );
  MUX2_X1 U8384 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n7241), .S(n7277), .Z(n7492)
         );
  MUX2_X1 U8385 ( .A(n7242), .B(P1_REG1_REG_2__SCAN_IN), .S(n10658), .Z(n10663) );
  MUX2_X1 U8386 ( .A(n7243), .B(P1_REG1_REG_1__SCAN_IN), .S(n10625), .Z(n10635) );
  NAND3_X1 U8387 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .A3(n10635), .ZN(n10634) );
  OAI21_X1 U8388 ( .B1(n10625), .B2(n7243), .A(n10634), .ZN(n10664) );
  NAND2_X1 U8389 ( .A1(n10663), .A2(n10664), .ZN(n10661) );
  OAI21_X1 U8390 ( .B1(n10658), .B2(n7242), .A(n10661), .ZN(n7491) );
  NAND2_X1 U8391 ( .A1(n7492), .A2(n7491), .ZN(n7490) );
  NAND2_X1 U8392 ( .A1(n7244), .A2(n7490), .ZN(n7679) );
  NOR2_X1 U8393 ( .A1(n7680), .A2(n7679), .ZN(n7678) );
  NOR2_X1 U8394 ( .A1(n7278), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7245) );
  NOR2_X1 U8395 ( .A1(n7678), .A2(n7245), .ZN(n7529) );
  NAND2_X1 U8396 ( .A1(n7528), .A2(n7529), .ZN(n7527) );
  NAND2_X1 U8397 ( .A1(n7246), .A2(n7527), .ZN(n7505) );
  NAND2_X1 U8398 ( .A1(n7504), .A2(n7505), .ZN(n7503) );
  NAND2_X1 U8399 ( .A1(n7247), .A2(n7503), .ZN(n7535) );
  MUX2_X1 U8400 ( .A(n7248), .B(P1_REG1_REG_7__SCAN_IN), .S(n7542), .Z(n7534)
         );
  NOR2_X1 U8401 ( .A1(n7535), .A2(n7534), .ZN(n7533) );
  NOR2_X1 U8402 ( .A1(n7249), .A2(n7533), .ZN(n7548) );
  MUX2_X1 U8403 ( .A(n7250), .B(P1_REG1_REG_8__SCAN_IN), .S(n7553), .Z(n7547)
         );
  NOR2_X1 U8404 ( .A1(n7548), .A2(n7547), .ZN(n7546) );
  INV_X1 U8405 ( .A(n7546), .ZN(n7251) );
  MUX2_X1 U8406 ( .A(n7253), .B(P1_REG1_REG_9__SCAN_IN), .S(n7567), .Z(n7562)
         );
  NOR2_X1 U8407 ( .A1(n7561), .A2(n7562), .ZN(n7560) );
  AOI21_X1 U8408 ( .B1(n7358), .B2(n7253), .A(n7560), .ZN(n7310) );
  MUX2_X1 U8409 ( .A(n7254), .B(P1_REG1_REG_10__SCAN_IN), .S(n7283), .Z(n7309)
         );
  NOR2_X1 U8410 ( .A1(n7310), .A2(n7309), .ZN(n7308) );
  AOI21_X1 U8411 ( .B1(n7254), .B2(n7402), .A(n7308), .ZN(n7631) );
  OR2_X1 U8412 ( .A1(n7628), .A2(n7631), .ZN(n7257) );
  NAND2_X1 U8413 ( .A1(n7629), .A2(n7255), .ZN(n7256) );
  NAND2_X1 U8414 ( .A1(n7257), .A2(n7256), .ZN(n7761) );
  NAND2_X1 U8415 ( .A1(n7760), .A2(n7761), .ZN(n7759) );
  NAND2_X1 U8416 ( .A1(n7258), .A2(n7759), .ZN(n7910) );
  NAND2_X1 U8417 ( .A1(n7911), .A2(n7910), .ZN(n7909) );
  OAI21_X1 U8418 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n7913), .A(n7909), .ZN(
        n7970) );
  NAND2_X1 U8419 ( .A1(n7971), .A2(n7970), .ZN(n7969) );
  OAI21_X1 U8420 ( .B1(n7289), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7969), .ZN(
        n7259) );
  NOR2_X1 U8421 ( .A1(n10111), .A2(n7259), .ZN(n7260) );
  XNOR2_X1 U8422 ( .A(n7259), .B(n10111), .ZN(n10108) );
  NOR2_X1 U8423 ( .A1(n6690), .A2(n10108), .ZN(n10107) );
  NOR2_X1 U8424 ( .A1(n7260), .A2(n10107), .ZN(n10121) );
  INV_X1 U8425 ( .A(n7293), .ZN(n10124) );
  NOR2_X1 U8426 ( .A1(n10124), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7261) );
  AOI21_X1 U8427 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n10124), .A(n7261), .ZN(
        n10120) );
  NOR2_X1 U8428 ( .A1(n10121), .A2(n10120), .ZN(n10119) );
  AOI21_X1 U8429 ( .B1(n7293), .B2(P1_REG1_REG_16__SCAN_IN), .A(n10119), .ZN(
        n7265) );
  AND2_X1 U8430 ( .A1(n7262), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7295) );
  NAND2_X1 U8431 ( .A1(n7295), .A2(n7263), .ZN(n8623) );
  INV_X1 U8432 ( .A(n7264), .ZN(n8620) );
  OR2_X1 U8433 ( .A1(n8623), .A2(n8620), .ZN(n10118) );
  NOR2_X1 U8434 ( .A1(n7265), .A2(n7266), .ZN(n10135) );
  AOI211_X1 U8435 ( .C1(n7266), .C2(n7265), .A(n10118), .B(n10135), .ZN(n7307)
         );
  NOR2_X1 U8436 ( .A1(n7289), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7267) );
  AOI21_X1 U8437 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n7289), .A(n7267), .ZN(
        n7967) );
  NAND2_X1 U8438 ( .A1(n7629), .A2(n10909), .ZN(n7286) );
  NAND2_X1 U8439 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n7283), .ZN(n7285) );
  NAND2_X1 U8440 ( .A1(n7567), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7268) );
  OAI21_X1 U8441 ( .B1(n7567), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7268), .ZN(
        n7564) );
  NOR2_X1 U8442 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n7553), .ZN(n7269) );
  AOI21_X1 U8443 ( .B1(n7553), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7269), .ZN(
        n7551) );
  NAND2_X1 U8444 ( .A1(n7281), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7270) );
  OAI21_X1 U8445 ( .B1(n7281), .B2(P1_REG2_REG_6__SCAN_IN), .A(n7270), .ZN(
        n7497) );
  NOR2_X1 U8446 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n7280), .ZN(n7271) );
  AOI21_X1 U8447 ( .B1(n7280), .B2(P1_REG2_REG_5__SCAN_IN), .A(n7271), .ZN(
        n7522) );
  INV_X1 U8448 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7273) );
  OR2_X1 U8449 ( .A1(n10658), .A2(n7273), .ZN(n7275) );
  NAND2_X1 U8450 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10630) );
  INV_X1 U8451 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7272) );
  MUX2_X1 U8452 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n7273), .S(n10658), .Z(n10667) );
  NOR2_X1 U8453 ( .A1(n10666), .A2(n10667), .ZN(n10665) );
  INV_X1 U8454 ( .A(n10665), .ZN(n7274) );
  NAND2_X1 U8455 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(n7277), .ZN(n7276) );
  OAI21_X1 U8456 ( .B1(n7277), .B2(P1_REG2_REG_3__SCAN_IN), .A(n7276), .ZN(
        n7485) );
  AOI22_X1 U8457 ( .A1(n7278), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7889), .B2(
        n7682), .ZN(n7674) );
  OR2_X1 U8458 ( .A1(n7278), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7279) );
  NAND2_X1 U8459 ( .A1(n7673), .A2(n7279), .ZN(n7523) );
  NAND2_X1 U8460 ( .A1(n7522), .A2(n7523), .ZN(n7521) );
  OAI21_X1 U8461 ( .B1(n7280), .B2(P1_REG2_REG_5__SCAN_IN), .A(n7521), .ZN(
        n7498) );
  NOR2_X1 U8462 ( .A1(n7542), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7282) );
  AOI21_X1 U8463 ( .B1(n7542), .B2(P1_REG2_REG_7__SCAN_IN), .A(n7282), .ZN(
        n7538) );
  NAND2_X1 U8464 ( .A1(n7551), .A2(n7550), .ZN(n7549) );
  OAI21_X1 U8465 ( .B1(n7553), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7549), .ZN(
        n7565) );
  OAI21_X1 U8466 ( .B1(n7283), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7285), .ZN(
        n7313) );
  NAND2_X1 U8467 ( .A1(n7285), .A2(n7284), .ZN(n7624) );
  NAND2_X1 U8468 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7763), .ZN(n7287) );
  OAI21_X1 U8469 ( .B1(n7763), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7287), .ZN(
        n7756) );
  AOI21_X1 U8470 ( .B1(n7763), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7755), .ZN(
        n7907) );
  MUX2_X1 U8471 ( .A(n7288), .B(P1_REG2_REG_13__SCAN_IN), .S(n7913), .Z(n7906)
         );
  NOR2_X1 U8472 ( .A1(n7907), .A2(n7906), .ZN(n7905) );
  AOI21_X1 U8473 ( .B1(n7913), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7905), .ZN(
        n7966) );
  NAND2_X1 U8474 ( .A1(n7967), .A2(n7966), .ZN(n7965) );
  NOR2_X1 U8475 ( .A1(n10111), .A2(n7290), .ZN(n7291) );
  NAND2_X1 U8476 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n7293), .ZN(n7292) );
  OAI21_X1 U8477 ( .B1(n7293), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7292), .ZN(
        n10116) );
  NOR2_X1 U8478 ( .A1(n10117), .A2(n10116), .ZN(n10115) );
  AOI21_X1 U8479 ( .B1(n7293), .B2(P1_REG2_REG_16__SCAN_IN), .A(n10115), .ZN(
        n7297) );
  NAND2_X1 U8480 ( .A1(n10136), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7294) );
  OAI21_X1 U8481 ( .B1(n10136), .B2(P1_REG2_REG_17__SCAN_IN), .A(n7294), .ZN(
        n7296) );
  NAND2_X1 U8482 ( .A1(n7295), .A2(n8620), .ZN(n7622) );
  OR2_X1 U8483 ( .A1(n7622), .A2(n7202), .ZN(n10627) );
  NOR2_X1 U8484 ( .A1(n7297), .A2(n7296), .ZN(n10128) );
  AOI211_X1 U8485 ( .C1(n7297), .C2(n7296), .A(n10627), .B(n10128), .ZN(n7306)
         );
  OR2_X1 U8486 ( .A1(n7622), .A2(n7670), .ZN(n10659) );
  INV_X1 U8487 ( .A(n10136), .ZN(n7298) );
  NOR2_X1 U8488 ( .A1(n10659), .A2(n7298), .ZN(n7305) );
  INV_X1 U8489 ( .A(n8750), .ZN(n7299) );
  NOR2_X1 U8490 ( .A1(n7300), .A2(n7299), .ZN(n7301) );
  OR2_X1 U8491 ( .A1(P1_U3083), .A2(n7301), .ZN(n7975) );
  INV_X1 U8492 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7303) );
  NAND2_X1 U8493 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n7302) );
  OAI21_X1 U8494 ( .B1(n7975), .B2(n7303), .A(n7302), .ZN(n7304) );
  OR4_X1 U8495 ( .A1(n7307), .A2(n7306), .A3(n7305), .A4(n7304), .ZN(P1_U3258)
         );
  AOI21_X1 U8496 ( .B1(n7310), .B2(n7309), .A(n7308), .ZN(n7311) );
  OAI22_X1 U8497 ( .A1(n7402), .A2(n10659), .B1(n10118), .B2(n7311), .ZN(n7319) );
  AOI211_X1 U8498 ( .C1(n7314), .C2(n7313), .A(n10627), .B(n7312), .ZN(n7318)
         );
  NOR2_X1 U8499 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7315), .ZN(n8882) );
  INV_X1 U8500 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7316) );
  NOR2_X1 U8501 ( .A1(n7975), .A2(n7316), .ZN(n7317) );
  OR4_X1 U8502 ( .A1(n7319), .A2(n7318), .A3(n8882), .A4(n7317), .ZN(P1_U3251)
         );
  AND2_X1 U8503 ( .A1(n7320), .A2(P2_U3152), .ZN(n7841) );
  INV_X2 U8504 ( .A(n7841), .ZN(n9923) );
  AND2_X1 U8505 ( .A1(n5740), .A2(P2_U3152), .ZN(n9910) );
  OAI222_X1 U8506 ( .A1(n9923), .A2(n7321), .B1(n7386), .B2(P2_U3152), .C1(
        n5076), .C2(n7323), .ZN(P2_U3357) );
  OAI222_X1 U8507 ( .A1(n9923), .A2(n7322), .B1(n7437), .B2(P2_U3152), .C1(
        n5076), .C2(n7327), .ZN(P2_U3356) );
  NOR2_X1 U8508 ( .A1(n5740), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10538) );
  NAND2_X1 U8509 ( .A1(n5740), .A2(P1_U3084), .ZN(n10546) );
  OAI222_X1 U8510 ( .A1(P1_U3084), .A2(n10625), .B1(n8088), .B2(n7323), .C1(
        n5479), .C2(n10546), .ZN(P1_U3352) );
  OAI222_X1 U8511 ( .A1(n9923), .A2(n7324), .B1(n7414), .B2(P2_U3152), .C1(
        n5076), .C2(n7325), .ZN(P2_U3355) );
  INV_X1 U8512 ( .A(n10546), .ZN(n7839) );
  INV_X1 U8513 ( .A(n7839), .ZN(n8845) );
  OAI222_X1 U8514 ( .A1(n8845), .A2(n7326), .B1(n8088), .B2(n7325), .C1(
        P1_U3084), .C2(n7495), .ZN(P1_U3350) );
  OAI222_X1 U8515 ( .A1(n8845), .A2(n7328), .B1(n8088), .B2(n7327), .C1(
        P1_U3084), .C2(n10658), .ZN(P1_U3351) );
  OAI222_X1 U8516 ( .A1(n8845), .A2(n7329), .B1(P1_U3084), .B2(n7682), .C1(
        n7330), .C2(n8088), .ZN(P1_U3349) );
  INV_X1 U8517 ( .A(n7467), .ZN(n7379) );
  OAI222_X1 U8518 ( .A1(n9923), .A2(n5384), .B1(n7379), .B2(P2_U3152), .C1(
        n5076), .C2(n7330), .ZN(P2_U3354) );
  INV_X1 U8519 ( .A(n7391), .ZN(n7426) );
  OAI222_X1 U8520 ( .A1(n5076), .A2(n7333), .B1(n7426), .B2(P2_U3152), .C1(
        n7331), .C2(n9923), .ZN(P2_U3353) );
  OAI222_X1 U8521 ( .A1(P1_U3084), .A2(n7532), .B1(n8088), .B2(n7333), .C1(
        n7332), .C2(n10546), .ZN(P1_U3348) );
  INV_X1 U8522 ( .A(n7451), .ZN(n7441) );
  INV_X1 U8523 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7334) );
  OAI222_X1 U8524 ( .A1(n5076), .A2(n7335), .B1(n7441), .B2(P2_U3152), .C1(
        n7334), .C2(n9923), .ZN(P2_U3352) );
  OAI222_X1 U8525 ( .A1(n8845), .A2(n7336), .B1(n8088), .B2(n7335), .C1(
        P1_U3084), .C2(n7508), .ZN(P1_U3347) );
  INV_X1 U8526 ( .A(n7514), .ZN(n7452) );
  INV_X1 U8527 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7337) );
  OAI222_X1 U8528 ( .A1(n5076), .A2(n7339), .B1(n7452), .B2(P2_U3152), .C1(
        n7337), .C2(n9923), .ZN(P2_U3351) );
  OAI222_X1 U8529 ( .A1(n8845), .A2(n7340), .B1(n8088), .B2(n7339), .C1(
        P1_U3084), .C2(n7338), .ZN(P1_U3346) );
  NAND2_X1 U8530 ( .A1(n7605), .A2(n7341), .ZN(n7342) );
  NAND2_X1 U8531 ( .A1(n7342), .A2(n7372), .ZN(n7345) );
  OR2_X1 U8532 ( .A1(n7605), .A2(n7343), .ZN(n7344) );
  AND2_X1 U8533 ( .A1(n7345), .A2(n7344), .ZN(n9487) );
  NOR2_X1 U8534 ( .A1(n9487), .A2(P2_U3966), .ZN(P2_U3151) );
  AOI22_X1 U8535 ( .A1(n7553), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n7839), .ZN(n7346) );
  OAI21_X1 U8536 ( .B1(n7348), .B2(n8088), .A(n7346), .ZN(P1_U3345) );
  INV_X1 U8537 ( .A(n7588), .ZN(n7593) );
  INV_X1 U8538 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7347) );
  OAI222_X1 U8539 ( .A1(n5076), .A2(n7348), .B1(n7593), .B2(P2_U3152), .C1(
        n7347), .C2(n9923), .ZN(P2_U3350) );
  INV_X1 U8540 ( .A(n7349), .ZN(n7350) );
  NAND2_X1 U8541 ( .A1(n7605), .A2(n7350), .ZN(n10584) );
  AOI22_X1 U8542 ( .A1(n5192), .A2(n7352), .B1(n7355), .B2(n7351), .ZN(
        P2_U3438) );
  INV_X1 U8543 ( .A(n7353), .ZN(n7354) );
  AOI22_X1 U8544 ( .A1(n5192), .A2(n7356), .B1(n7355), .B2(n7354), .ZN(
        P2_U3437) );
  INV_X1 U8545 ( .A(n7357), .ZN(n7359) );
  INV_X1 U8546 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7367) );
  OAI222_X1 U8547 ( .A1(n7358), .A2(P1_U3084), .B1(n8088), .B2(n7359), .C1(
        n8845), .C2(n7367), .ZN(P1_U3344) );
  INV_X1 U8548 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7360) );
  INV_X1 U8549 ( .A(n7709), .ZN(n7715) );
  OAI222_X1 U8550 ( .A1(n9923), .A2(n7360), .B1(n5076), .B2(n7359), .C1(
        P2_U3152), .C2(n7715), .ZN(P2_U3349) );
  NAND2_X1 U8551 ( .A1(n9406), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7361) );
  OAI21_X1 U8552 ( .B1(n9532), .B2(n9406), .A(n7361), .ZN(P2_U3582) );
  INV_X1 U8553 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7364) );
  NAND2_X1 U8554 ( .A1(n7362), .A2(P2_U3966), .ZN(n7363) );
  OAI21_X1 U8555 ( .B1(P2_U3966), .B2(n7364), .A(n7363), .ZN(P2_U3583) );
  NAND2_X1 U8556 ( .A1(n9406), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n7365) );
  OAI21_X1 U8557 ( .B1(n9719), .B2(n9406), .A(n7365), .ZN(P2_U3570) );
  INV_X1 U8558 ( .A(n8677), .ZN(n8669) );
  NAND2_X1 U8559 ( .A1(n8669), .A2(P2_U3966), .ZN(n7366) );
  OAI21_X1 U8560 ( .B1(P2_U3966), .B2(n7367), .A(n7366), .ZN(P2_U3561) );
  INV_X1 U8561 ( .A(n8038), .ZN(n7835) );
  INV_X1 U8562 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7368) );
  OAI222_X1 U8563 ( .A1(n5076), .A2(n7401), .B1(n7835), .B2(P2_U3152), .C1(
        n7368), .C2(n9923), .ZN(P2_U3347) );
  NAND2_X1 U8564 ( .A1(n7605), .A2(n7369), .ZN(n7370) );
  OAI211_X1 U8565 ( .C1(P2_U3152), .C2(n7371), .A(n7370), .B(n8754), .ZN(n7373) );
  NAND2_X1 U8566 ( .A1(n7373), .A2(n7372), .ZN(n7381) );
  NAND2_X1 U8567 ( .A1(n7381), .A2(n9406), .ZN(n7393) );
  NAND2_X1 U8568 ( .A1(n7393), .A2(n8925), .ZN(n9490) );
  NAND2_X1 U8569 ( .A1(P2_U3152), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7855) );
  INV_X1 U8570 ( .A(n7855), .ZN(n7385) );
  NAND2_X1 U8571 ( .A1(n7391), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7380) );
  MUX2_X1 U8572 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n7374), .S(n7391), .Z(n7422)
         );
  NAND2_X1 U8573 ( .A1(n7389), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7377) );
  MUX2_X1 U8574 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n7375), .S(n7389), .Z(n7411)
         );
  MUX2_X1 U8575 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n7376), .S(n7387), .Z(n7433)
         );
  INV_X1 U8576 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10717) );
  MUX2_X1 U8577 ( .A(n10717), .B(P2_REG1_REG_1__SCAN_IN), .S(n7386), .Z(n10653) );
  NAND3_X1 U8578 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n10653), .ZN(n10651) );
  OAI21_X1 U8579 ( .B1(n7386), .B2(n10717), .A(n10651), .ZN(n7434) );
  NAND2_X1 U8580 ( .A1(n7433), .A2(n7434), .ZN(n7432) );
  OAI21_X1 U8581 ( .B1(n7437), .B2(n7376), .A(n7432), .ZN(n7410) );
  NAND2_X1 U8582 ( .A1(n7411), .A2(n7410), .ZN(n7409) );
  NAND2_X1 U8583 ( .A1(n7377), .A2(n7409), .ZN(n7460) );
  MUX2_X1 U8584 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n7378), .S(n7467), .Z(n7459)
         );
  NAND2_X1 U8585 ( .A1(n7460), .A2(n7459), .ZN(n7458) );
  OAI21_X1 U8586 ( .B1(n7379), .B2(n7378), .A(n7458), .ZN(n7421) );
  NAND2_X1 U8587 ( .A1(n7422), .A2(n7421), .ZN(n7420) );
  AND2_X1 U8588 ( .A1(n7380), .A2(n7420), .ZN(n7383) );
  INV_X1 U8589 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10824) );
  MUX2_X1 U8590 ( .A(n10824), .B(P2_REG1_REG_6__SCAN_IN), .S(n7451), .Z(n7382)
         );
  NOR2_X1 U8591 ( .A1(n7383), .A2(n7382), .ZN(n7447) );
  OR2_X1 U8592 ( .A1(n7381), .A2(n9496), .ZN(n9464) );
  AOI211_X1 U8593 ( .C1(n7383), .C2(n7382), .A(n7447), .B(n9464), .ZN(n7384)
         );
  AOI211_X1 U8594 ( .C1(n9487), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n7385), .B(
        n7384), .ZN(n7397) );
  MUX2_X1 U8595 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n9790), .S(n7451), .Z(n7395)
         );
  XNOR2_X1 U8596 ( .A(n7467), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n7464) );
  NAND2_X1 U8597 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10644) );
  NOR2_X1 U8598 ( .A1(n10645), .A2(n10644), .ZN(n10643) );
  AOI21_X1 U8599 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n10648), .A(n10643), .ZN(
        n7430) );
  AOI22_X1 U8600 ( .A1(n7387), .A2(n5758), .B1(P2_REG2_REG_2__SCAN_IN), .B2(
        n7437), .ZN(n7431) );
  NAND2_X1 U8601 ( .A1(n7389), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7388) );
  OAI21_X1 U8602 ( .B1(n7389), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7388), .ZN(
        n7407) );
  NOR2_X1 U8603 ( .A1(n7464), .A2(n5127), .ZN(n7463) );
  NAND2_X1 U8604 ( .A1(n7391), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7390) );
  OAI21_X1 U8605 ( .B1(n7391), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7390), .ZN(
        n7418) );
  NAND3_X1 U8606 ( .A1(n7393), .A2(n7392), .A3(n9496), .ZN(n10642) );
  INV_X1 U8607 ( .A(n10642), .ZN(n9474) );
  NAND2_X1 U8608 ( .A1(n7395), .A2(n7394), .ZN(n7450) );
  OAI211_X1 U8609 ( .C1(n7395), .C2(n7394), .A(n9474), .B(n7450), .ZN(n7396)
         );
  OAI211_X1 U8610 ( .C1(n9490), .C2(n7441), .A(n7397), .B(n7396), .ZN(P2_U3251) );
  INV_X1 U8611 ( .A(n7398), .ZN(n7403) );
  INV_X1 U8612 ( .A(n7824), .ZN(n7828) );
  INV_X1 U8613 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7399) );
  OAI222_X1 U8614 ( .A1(n5076), .A2(n7403), .B1(n7828), .B2(P2_U3152), .C1(
        n7399), .C2(n9923), .ZN(P2_U3348) );
  INV_X1 U8615 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n7400) );
  OAI222_X1 U8616 ( .A1(P1_U3084), .A2(n7629), .B1(n8088), .B2(n7401), .C1(
        n7400), .C2(n8845), .ZN(P1_U3342) );
  INV_X1 U8617 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7404) );
  OAI222_X1 U8618 ( .A1(n8845), .A2(n7404), .B1(n8088), .B2(n7403), .C1(
        P1_U3084), .C2(n7402), .ZN(P1_U3343) );
  INV_X1 U8619 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7577) );
  INV_X1 U8620 ( .A(n9508), .ZN(n9758) );
  NAND2_X1 U8621 ( .A1(n9758), .A2(P2_U3966), .ZN(n7405) );
  OAI21_X1 U8622 ( .B1(P2_U3966), .B2(n7577), .A(n7405), .ZN(P2_U3566) );
  AOI211_X1 U8623 ( .C1(n7408), .C2(n7407), .A(n7406), .B(n10642), .ZN(n7416)
         );
  INV_X1 U8624 ( .A(n9464), .ZN(n10652) );
  OAI211_X1 U8625 ( .C1(n7411), .C2(n7410), .A(n10652), .B(n7409), .ZN(n7413)
         );
  AOI22_X1 U8626 ( .A1(n9487), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(P2_U3152), .ZN(n7412) );
  OAI211_X1 U8627 ( .C1(n9490), .C2(n7414), .A(n7413), .B(n7412), .ZN(n7415)
         );
  OR2_X1 U8628 ( .A1(n7416), .A2(n7415), .ZN(P2_U3248) );
  AOI211_X1 U8629 ( .C1(n7419), .C2(n7418), .A(n7417), .B(n10642), .ZN(n7428)
         );
  OAI211_X1 U8630 ( .C1(n7422), .C2(n7421), .A(n10652), .B(n7420), .ZN(n7425)
         );
  NOR2_X1 U8631 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8488), .ZN(n7423) );
  AOI21_X1 U8632 ( .B1(n9487), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n7423), .ZN(
        n7424) );
  OAI211_X1 U8633 ( .C1(n9490), .C2(n7426), .A(n7425), .B(n7424), .ZN(n7427)
         );
  OR2_X1 U8634 ( .A1(n7428), .A2(n7427), .ZN(P2_U3250) );
  AOI211_X1 U8635 ( .C1(n7431), .C2(n7430), .A(n7429), .B(n10642), .ZN(n7439)
         );
  OAI211_X1 U8636 ( .C1(n7434), .C2(n7433), .A(n10652), .B(n7432), .ZN(n7436)
         );
  AOI22_X1 U8637 ( .A1(n9487), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n7435) );
  OAI211_X1 U8638 ( .C1(n9490), .C2(n7437), .A(n7436), .B(n7435), .ZN(n7438)
         );
  OR2_X1 U8639 ( .A1(n7439), .A2(n7438), .ZN(P2_U3247) );
  AOI22_X1 U8640 ( .A1(n7763), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n7839), .ZN(n7440) );
  OAI21_X1 U8641 ( .B1(n7470), .B2(n8088), .A(n7440), .ZN(P1_U3341) );
  INV_X1 U8642 ( .A(n9490), .ZN(n10649) );
  INV_X1 U8643 ( .A(n9487), .ZN(n10641) );
  INV_X1 U8644 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7449) );
  INV_X1 U8645 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10839) );
  MUX2_X1 U8646 ( .A(n10839), .B(P2_REG1_REG_7__SCAN_IN), .S(n7514), .Z(n7443)
         );
  NOR2_X1 U8647 ( .A1(n7441), .A2(n10824), .ZN(n7445) );
  INV_X1 U8648 ( .A(n7445), .ZN(n7442) );
  NAND2_X1 U8649 ( .A1(n7443), .A2(n7442), .ZN(n7446) );
  MUX2_X1 U8650 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10839), .S(n7514), .Z(n7444)
         );
  OAI21_X1 U8651 ( .B1(n7447), .B2(n7445), .A(n7444), .ZN(n7511) );
  OAI211_X1 U8652 ( .C1(n7447), .C2(n7446), .A(n7511), .B(n10652), .ZN(n7448)
         );
  NAND2_X1 U8653 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7899) );
  OAI211_X1 U8654 ( .C1(n10641), .C2(n7449), .A(n7448), .B(n7899), .ZN(n7456)
         );
  AOI22_X1 U8655 ( .A1(n7514), .A2(n8053), .B1(P2_REG2_REG_7__SCAN_IN), .B2(
        n7452), .ZN(n7453) );
  AOI211_X1 U8656 ( .C1(n7454), .C2(n7453), .A(n7513), .B(n10642), .ZN(n7455)
         );
  AOI211_X1 U8657 ( .C1(n10649), .C2(n7514), .A(n7456), .B(n7455), .ZN(n7457)
         );
  INV_X1 U8658 ( .A(n7457), .ZN(P2_U3252) );
  INV_X1 U8659 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7462) );
  OAI211_X1 U8660 ( .C1(n7460), .C2(n7459), .A(n10652), .B(n7458), .ZN(n7461)
         );
  NAND2_X1 U8661 ( .A1(P2_U3152), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7726) );
  OAI211_X1 U8662 ( .C1(n10641), .C2(n7462), .A(n7461), .B(n7726), .ZN(n7466)
         );
  AOI211_X1 U8663 ( .C1(n5127), .C2(n7464), .A(n7463), .B(n10642), .ZN(n7465)
         );
  AOI211_X1 U8664 ( .C1(n10649), .C2(n7467), .A(n7466), .B(n7465), .ZN(n7468)
         );
  INV_X1 U8665 ( .A(n7468), .ZN(P2_U3249) );
  INV_X1 U8666 ( .A(n8072), .ZN(n8077) );
  INV_X1 U8667 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7469) );
  OAI222_X1 U8668 ( .A1(n5076), .A2(n7470), .B1(n8077), .B2(P2_U3152), .C1(
        n7469), .C2(n9923), .ZN(P2_U3346) );
  INV_X1 U8669 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n7474) );
  NAND2_X1 U8670 ( .A1(n6706), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n7473) );
  INV_X1 U8671 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n7471) );
  OR2_X1 U8672 ( .A1(n8941), .A2(n7471), .ZN(n7472) );
  OAI211_X1 U8673 ( .C1(n8942), .C2(n7474), .A(n7473), .B(n7472), .ZN(n10159)
         );
  NAND2_X1 U8674 ( .A1(n10159), .A2(n10104), .ZN(n7475) );
  OAI21_X1 U8675 ( .B1(n10104), .B2(n9915), .A(n7475), .ZN(P1_U3586) );
  INV_X1 U8676 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7477) );
  NAND2_X1 U8677 ( .A1(n9225), .A2(n10104), .ZN(n7476) );
  OAI21_X1 U8678 ( .B1(n10104), .B2(n7477), .A(n7476), .ZN(P1_U3578) );
  AOI22_X1 U8679 ( .A1(n9474), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10652), .ZN(n7481) );
  INV_X1 U8680 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7479) );
  OAI21_X1 U8681 ( .B1(n9464), .B2(P2_REG1_REG_0__SCAN_IN), .A(n9490), .ZN(
        n7478) );
  AOI21_X1 U8682 ( .B1(n9474), .B2(n7479), .A(n7478), .ZN(n7480) );
  MUX2_X1 U8683 ( .A(n7481), .B(n7480), .S(P2_IR_REG_0__SCAN_IN), .Z(n7483) );
  AOI22_X1 U8684 ( .A1(n9487), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n7482) );
  NAND2_X1 U8685 ( .A1(n7483), .A2(n7482), .ZN(P2_U3245) );
  AOI211_X1 U8686 ( .C1(n7486), .C2(n7485), .A(n10627), .B(n7484), .ZN(n7489)
         );
  AND2_X1 U8687 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7809) );
  INV_X1 U8688 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7487) );
  NOR2_X1 U8689 ( .A1(n7975), .A2(n7487), .ZN(n7488) );
  NOR3_X1 U8690 ( .A1(n7489), .A2(n7809), .A3(n7488), .ZN(n7494) );
  INV_X1 U8691 ( .A(n10118), .ZN(n10662) );
  OAI211_X1 U8692 ( .C1(n7492), .C2(n7491), .A(n10662), .B(n7490), .ZN(n7493)
         );
  OAI211_X1 U8693 ( .C1(n10659), .C2(n7495), .A(n7494), .B(n7493), .ZN(
        P1_U3244) );
  AOI211_X1 U8694 ( .C1(n7498), .C2(n7497), .A(n10627), .B(n7496), .ZN(n7502)
         );
  INV_X1 U8695 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7499) );
  NOR2_X1 U8696 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7499), .ZN(n8104) );
  INV_X1 U8697 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n7500) );
  NOR2_X1 U8698 ( .A1(n7975), .A2(n7500), .ZN(n7501) );
  NOR3_X1 U8699 ( .A1(n7502), .A2(n8104), .A3(n7501), .ZN(n7507) );
  OAI211_X1 U8700 ( .C1(n7505), .C2(n7504), .A(n10662), .B(n7503), .ZN(n7506)
         );
  OAI211_X1 U8701 ( .C1(n10659), .C2(n7508), .A(n7507), .B(n7506), .ZN(
        P1_U3247) );
  NAND2_X1 U8702 ( .A1(n7514), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7510) );
  INV_X1 U8703 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10857) );
  MUX2_X1 U8704 ( .A(n10857), .B(P2_REG1_REG_8__SCAN_IN), .S(n7588), .Z(n7509)
         );
  AOI21_X1 U8705 ( .B1(n7511), .B2(n7510), .A(n7509), .ZN(n7599) );
  AND3_X1 U8706 ( .A1(n7511), .A2(n7510), .A3(n7509), .ZN(n7512) );
  NOR3_X1 U8707 ( .A1(n7599), .A2(n7512), .A3(n9464), .ZN(n7518) );
  XNOR2_X1 U8708 ( .A(n7588), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n7515) );
  NOR2_X1 U8709 ( .A1(n7515), .A2(n7516), .ZN(n7587) );
  AOI211_X1 U8710 ( .C1(n7516), .C2(n7515), .A(n7587), .B(n10642), .ZN(n7517)
         );
  NOR2_X1 U8711 ( .A1(n7518), .A2(n7517), .ZN(n7520) );
  NOR2_X1 U8712 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8474), .ZN(n8110) );
  AOI21_X1 U8713 ( .B1(n9487), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n8110), .ZN(
        n7519) );
  OAI211_X1 U8714 ( .C1(n7593), .C2(n9490), .A(n7520), .B(n7519), .ZN(P2_U3253) );
  INV_X1 U8715 ( .A(n10627), .ZN(n10669) );
  OAI21_X1 U8716 ( .B1(n7523), .B2(n7522), .A(n7521), .ZN(n7526) );
  AND2_X1 U8717 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n8094) );
  INV_X1 U8718 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7524) );
  NOR2_X1 U8719 ( .A1(n7975), .A2(n7524), .ZN(n7525) );
  AOI211_X1 U8720 ( .C1(n10669), .C2(n7526), .A(n8094), .B(n7525), .ZN(n7531)
         );
  OAI211_X1 U8721 ( .C1(n7529), .C2(n7528), .A(n10662), .B(n7527), .ZN(n7530)
         );
  OAI211_X1 U8722 ( .C1(n10659), .C2(n7532), .A(n7531), .B(n7530), .ZN(
        P1_U3246) );
  AOI21_X1 U8723 ( .B1(n7535), .B2(n7534), .A(n7533), .ZN(n7545) );
  OAI21_X1 U8724 ( .B1(n7538), .B2(n7537), .A(n7536), .ZN(n7541) );
  AND2_X1 U8725 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8696) );
  INV_X1 U8726 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7539) );
  NOR2_X1 U8727 ( .A1(n7975), .A2(n7539), .ZN(n7540) );
  AOI211_X1 U8728 ( .C1(n10669), .C2(n7541), .A(n8696), .B(n7540), .ZN(n7544)
         );
  INV_X1 U8729 ( .A(n10659), .ZN(n10151) );
  NAND2_X1 U8730 ( .A1(n10151), .A2(n7542), .ZN(n7543) );
  OAI211_X1 U8731 ( .C1(n7545), .C2(n10118), .A(n7544), .B(n7543), .ZN(
        P1_U3248) );
  AOI21_X1 U8732 ( .B1(n7548), .B2(n7547), .A(n7546), .ZN(n7557) );
  OAI21_X1 U8733 ( .B1(n7551), .B2(n7550), .A(n7549), .ZN(n7552) );
  AOI22_X1 U8734 ( .A1(n7553), .A2(n10151), .B1(n10669), .B2(n7552), .ZN(n7556) );
  INV_X1 U8735 ( .A(n7975), .ZN(n10670) );
  INV_X1 U8736 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7554) );
  NOR2_X1 U8737 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7554), .ZN(n8767) );
  AOI21_X1 U8738 ( .B1(n10670), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n8767), .ZN(
        n7555) );
  OAI211_X1 U8739 ( .C1(n7557), .C2(n10118), .A(n7556), .B(n7555), .ZN(
        P1_U3249) );
  INV_X1 U8740 ( .A(n7558), .ZN(n7571) );
  AOI22_X1 U8741 ( .A1(n7913), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n7839), .ZN(n7559) );
  OAI21_X1 U8742 ( .B1(n7571), .B2(n8088), .A(n7559), .ZN(P1_U3340) );
  AOI21_X1 U8743 ( .B1(n7562), .B2(n7561), .A(n7560), .ZN(n7570) );
  AND2_X1 U8744 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n10010) );
  AOI211_X1 U8745 ( .C1(n7565), .C2(n7564), .A(n10627), .B(n7563), .ZN(n7566)
         );
  AOI211_X1 U8746 ( .C1(n10670), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n10010), .B(
        n7566), .ZN(n7569) );
  NAND2_X1 U8747 ( .A1(n10151), .A2(n7567), .ZN(n7568) );
  OAI211_X1 U8748 ( .C1(n7570), .C2(n10118), .A(n7569), .B(n7568), .ZN(
        P1_U3250) );
  INV_X1 U8749 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7572) );
  INV_X1 U8750 ( .A(n8192), .ZN(n8188) );
  OAI222_X1 U8751 ( .A1(n9923), .A2(n7572), .B1(n5076), .B2(n7571), .C1(
        P2_U3152), .C2(n8188), .ZN(P2_U3345) );
  NAND2_X1 U8752 ( .A1(n9406), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7573) );
  OAI21_X1 U8753 ( .B1(n9304), .B2(n9406), .A(n7573), .ZN(P2_U3581) );
  NAND2_X1 U8754 ( .A1(n9406), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7574) );
  OAI21_X1 U8755 ( .B1(n9565), .B2(n9406), .A(n7574), .ZN(P2_U3578) );
  INV_X1 U8756 ( .A(n9410), .ZN(n9417) );
  INV_X1 U8757 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7575) );
  OAI222_X1 U8758 ( .A1(n5076), .A2(n7576), .B1(n9417), .B2(P2_U3152), .C1(
        n7575), .C2(n9923), .ZN(P2_U3344) );
  OAI222_X1 U8759 ( .A1(n7972), .A2(P1_U3084), .B1(n8845), .B2(n7577), .C1(
        n7576), .C2(n8088), .ZN(P1_U3339) );
  INV_X1 U8760 ( .A(n6735), .ZN(n7866) );
  INV_X1 U8761 ( .A(n11015), .ZN(n10721) );
  INV_X1 U8762 ( .A(n7648), .ZN(n7578) );
  NOR2_X1 U8763 ( .A1(n10623), .A2(n7578), .ZN(n7688) );
  OAI211_X1 U8764 ( .C1(n7580), .C2(n10721), .A(n7688), .B(n7579), .ZN(n10048)
         );
  AOI22_X1 U8765 ( .A1(n10069), .A2(n7699), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n10048), .ZN(n7585) );
  OAI21_X1 U8766 ( .B1(n7583), .B2(n7581), .A(n7582), .ZN(n7667) );
  NAND2_X1 U8767 ( .A1(n7667), .A2(n10078), .ZN(n7584) );
  OAI211_X1 U8768 ( .C1(n7866), .C2(n10065), .A(n7585), .B(n7584), .ZN(
        P1_U3230) );
  INV_X1 U8769 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7586) );
  NAND2_X1 U8770 ( .A1(P2_U3152), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8138) );
  OAI21_X1 U8771 ( .B1(n10641), .B2(n7586), .A(n8138), .ZN(n7592) );
  AOI21_X1 U8772 ( .B1(n7588), .B2(P2_REG2_REG_8__SCAN_IN), .A(n7587), .ZN(
        n7590) );
  AOI22_X1 U8773 ( .A1(n7709), .A2(n8655), .B1(P2_REG2_REG_9__SCAN_IN), .B2(
        n7715), .ZN(n7589) );
  AOI211_X1 U8774 ( .C1(n7590), .C2(n7589), .A(n7708), .B(n10642), .ZN(n7591)
         );
  AOI211_X1 U8775 ( .C1(n10649), .C2(n7709), .A(n7592), .B(n7591), .ZN(n7601)
         );
  INV_X1 U8776 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10871) );
  MUX2_X1 U8777 ( .A(n10871), .B(P2_REG1_REG_9__SCAN_IN), .S(n7709), .Z(n7595)
         );
  NOR2_X1 U8778 ( .A1(n7593), .A2(n10857), .ZN(n7597) );
  INV_X1 U8779 ( .A(n7597), .ZN(n7594) );
  NAND2_X1 U8780 ( .A1(n7595), .A2(n7594), .ZN(n7598) );
  MUX2_X1 U8781 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10871), .S(n7709), .Z(n7596)
         );
  OAI21_X1 U8782 ( .B1(n7599), .B2(n7597), .A(n7596), .ZN(n7714) );
  OAI211_X1 U8783 ( .C1(n7599), .C2(n7598), .A(n7714), .B(n10652), .ZN(n7600)
         );
  NAND2_X1 U8784 ( .A1(n7601), .A2(n7600), .ZN(P2_U3254) );
  XOR2_X1 U8785 ( .A(n7746), .B(n7743), .Z(n7603) );
  NOR2_X1 U8786 ( .A1(n7603), .A2(n7602), .ZN(n7744) );
  AOI21_X1 U8787 ( .B1(n7603), .B2(n7602), .A(n7744), .ZN(n7610) );
  INV_X1 U8788 ( .A(n9408), .ZN(n7604) );
  INV_X1 U8789 ( .A(n10926), .ZN(n9720) );
  OAI22_X1 U8790 ( .A1(n7604), .A2(n9774), .B1(n7778), .B2(n9720), .ZN(n10696)
         );
  NAND2_X1 U8791 ( .A1(n7607), .A2(n7766), .ZN(n7751) );
  AOI22_X1 U8792 ( .A1(n9384), .A2(n10696), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n7751), .ZN(n7609) );
  NAND2_X1 U8793 ( .A1(n9389), .A2(n7771), .ZN(n7608) );
  OAI211_X1 U8794 ( .C1(n7610), .C2(n9391), .A(n7609), .B(n7608), .ZN(P2_U3224) );
  INV_X1 U8795 ( .A(n9423), .ZN(n9429) );
  INV_X1 U8796 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7611) );
  OAI222_X1 U8797 ( .A1(n5076), .A2(n7613), .B1(n9429), .B2(P2_U3152), .C1(
        n7611), .C2(n9923), .ZN(P2_U3343) );
  INV_X1 U8798 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7612) );
  OAI222_X1 U8799 ( .A1(P1_U3084), .A2(n10111), .B1(n8088), .B2(n7613), .C1(
        n7612), .C2(n10546), .ZN(P1_U3338) );
  NAND2_X1 U8800 ( .A1(n7751), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7618) );
  INV_X1 U8801 ( .A(n7614), .ZN(n7616) );
  AOI21_X1 U8802 ( .B1(n9408), .B2(n9295), .A(n10680), .ZN(n7615) );
  OR3_X1 U8803 ( .A1(n9391), .A2(n7616), .A3(n7615), .ZN(n7617) );
  OAI211_X1 U8804 ( .C1(n9335), .C2(n10699), .A(n7618), .B(n7617), .ZN(n7619)
         );
  INV_X1 U8805 ( .A(n7619), .ZN(n7620) );
  OAI21_X1 U8806 ( .B1(n8148), .B2(n9372), .A(n7620), .ZN(P2_U3234) );
  NAND2_X1 U8807 ( .A1(n7624), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7621) );
  OAI21_X1 U8808 ( .B1(n7622), .B2(n7621), .A(n10659), .ZN(n7635) );
  MUX2_X1 U8809 ( .A(n10909), .B(P1_REG2_REG_11__SCAN_IN), .S(n7629), .Z(n7625) );
  OAI21_X1 U8810 ( .B1(n7625), .B2(n7624), .A(n7623), .ZN(n7627) );
  NAND2_X1 U8811 ( .A1(n10670), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n7626) );
  NAND2_X1 U8812 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8891) );
  OAI211_X1 U8813 ( .C1(n10627), .C2(n7627), .A(n7626), .B(n8891), .ZN(n7634)
         );
  AOI21_X1 U8814 ( .B1(n7255), .B2(n7629), .A(n7628), .ZN(n7630) );
  XNOR2_X1 U8815 ( .A(n7631), .B(n7630), .ZN(n7632) );
  NOR2_X1 U8816 ( .A1(n7632), .A2(n10118), .ZN(n7633) );
  AOI211_X1 U8817 ( .C1(n7636), .C2(n7635), .A(n7634), .B(n7633), .ZN(n7637)
         );
  INV_X1 U8818 ( .A(n7637), .ZN(P1_U3252) );
  NAND2_X1 U8819 ( .A1(n7638), .A2(n7639), .ZN(n7641) );
  XNOR2_X1 U8820 ( .A(n7641), .B(n7640), .ZN(n7646) );
  AOI22_X1 U8821 ( .A1(n10069), .A2(n6736), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n10048), .ZN(n7645) );
  AOI22_X1 U8822 ( .A1(n10086), .A2(n7642), .B1(n10081), .B2(n7643), .ZN(n7644) );
  OAI211_X1 U8823 ( .C1(n7646), .C2(n10071), .A(n7645), .B(n7644), .ZN(
        P1_U3220) );
  AND2_X1 U8824 ( .A1(n7647), .A2(n10531), .ZN(n10621) );
  NAND2_X1 U8825 ( .A1(n7649), .A2(n7648), .ZN(n7650) );
  NOR2_X1 U8826 ( .A1(n7651), .A2(n7650), .ZN(n7652) );
  INV_X1 U8827 ( .A(n7689), .ZN(n10532) );
  AND2_X2 U8828 ( .A1(n7658), .A2(n10532), .ZN(n11020) );
  INV_X1 U8829 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10632) );
  INV_X1 U8830 ( .A(n7699), .ZN(n7801) );
  NAND2_X1 U8831 ( .A1(n7643), .A2(n7801), .ZN(n9084) );
  INV_X1 U8832 ( .A(n9084), .ZN(n7653) );
  OR2_X1 U8833 ( .A1(n7653), .A2(n7865), .ZN(n9121) );
  NOR2_X1 U8834 ( .A1(n7655), .A2(n7654), .ZN(n7656) );
  AOI22_X1 U8835 ( .A1(n9121), .A2(n7656), .B1(n10398), .B2(n6735), .ZN(n7805)
         );
  OAI21_X1 U8836 ( .B1(n7801), .B2(n7799), .A(n7805), .ZN(n7659) );
  NAND2_X1 U8837 ( .A1(n7659), .A2(n11020), .ZN(n7657) );
  OAI21_X1 U8838 ( .B1(n11020), .B2(n10632), .A(n7657), .ZN(P1_U3523) );
  AND2_X2 U8839 ( .A1(n7658), .A2(n7689), .ZN(n11024) );
  INV_X1 U8840 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7661) );
  NAND2_X1 U8841 ( .A1(n7659), .A2(n11024), .ZN(n7660) );
  OAI21_X1 U8842 ( .B1(n11024), .B2(n7661), .A(n7660), .ZN(P1_U3454) );
  INV_X1 U8843 ( .A(n7662), .ZN(n7664) );
  INV_X1 U8844 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7663) );
  OAI222_X1 U8845 ( .A1(n10124), .A2(P1_U3084), .B1(n8088), .B2(n7664), .C1(
        n7663), .C2(n10546), .ZN(P1_U3337) );
  INV_X1 U8846 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7665) );
  INV_X1 U8847 ( .A(n9442), .ZN(n9448) );
  OAI222_X1 U8848 ( .A1(n9923), .A2(n7665), .B1(n5076), .B2(n7664), .C1(
        P2_U3152), .C2(n9448), .ZN(P2_U3342) );
  AOI22_X1 U8849 ( .A1(n10136), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n7839), .ZN(n7666) );
  OAI21_X1 U8850 ( .B1(n7706), .B2(n8088), .A(n7666), .ZN(P1_U3336) );
  AOI21_X1 U8851 ( .B1(n8620), .B2(n6705), .A(n7202), .ZN(n8619) );
  INV_X1 U8852 ( .A(n10630), .ZN(n7669) );
  INV_X1 U8853 ( .A(n7667), .ZN(n7668) );
  MUX2_X1 U8854 ( .A(n7669), .B(n7668), .S(n7264), .Z(n7671) );
  NAND2_X1 U8855 ( .A1(n7671), .A2(n7670), .ZN(n7672) );
  OAI211_X1 U8856 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n8619), .A(n7672), .B(
        n10104), .ZN(n10674) );
  OAI21_X1 U8857 ( .B1(n7675), .B2(n7674), .A(n7673), .ZN(n7685) );
  INV_X1 U8858 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7677) );
  AND2_X1 U8859 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7848) );
  INV_X1 U8860 ( .A(n7848), .ZN(n7676) );
  OAI21_X1 U8861 ( .B1(n7975), .B2(n7677), .A(n7676), .ZN(n7684) );
  AOI21_X1 U8862 ( .B1(n7680), .B2(n7679), .A(n7678), .ZN(n7681) );
  OAI22_X1 U8863 ( .A1(n7682), .A2(n10659), .B1(n10118), .B2(n7681), .ZN(n7683) );
  AOI211_X1 U8864 ( .C1(n10669), .C2(n7685), .A(n7684), .B(n7683), .ZN(n7686)
         );
  NAND2_X1 U8865 ( .A1(n10674), .A2(n7686), .ZN(P1_U3245) );
  INV_X1 U8866 ( .A(n7687), .ZN(n7691) );
  AND2_X1 U8867 ( .A1(n7689), .A2(n7688), .ZN(n7690) );
  NAND2_X1 U8868 ( .A1(n7691), .A2(n7690), .ZN(n7996) );
  NOR2_X1 U8869 ( .A1(n7693), .A2(n10289), .ZN(n7864) );
  INV_X1 U8870 ( .A(n7864), .ZN(n7694) );
  NAND2_X1 U8871 ( .A1(n10895), .A2(n7694), .ZN(n10799) );
  NAND2_X1 U8872 ( .A1(n5074), .A2(n10799), .ZN(n10381) );
  NAND2_X1 U8873 ( .A1(n7643), .A2(n7699), .ZN(n7695) );
  XNOR2_X1 U8874 ( .A(n9128), .B(n7695), .ZN(n10687) );
  INV_X1 U8875 ( .A(n7642), .ZN(n10743) );
  XOR2_X1 U8876 ( .A(n7865), .B(n9128), .Z(n7698) );
  OR2_X1 U8877 ( .A1(n8630), .A2(n10289), .ZN(n7696) );
  NAND2_X1 U8878 ( .A1(n9169), .A2(n9167), .ZN(n9180) );
  NAND2_X1 U8879 ( .A1(n7696), .A2(n9180), .ZN(n10892) );
  INV_X1 U8880 ( .A(n10892), .ZN(n10784) );
  INV_X1 U8881 ( .A(n7643), .ZN(n7697) );
  OAI222_X1 U8882 ( .A1(n10887), .A2(n10743), .B1(n7698), .B2(n10784), .C1(
        n10889), .C2(n7697), .ZN(n10692) );
  INV_X1 U8883 ( .A(n7873), .ZN(n7700) );
  AND2_X1 U8884 ( .A1(n6736), .A2(n7699), .ZN(n7861) );
  OR2_X1 U8885 ( .A1(n7799), .A2(n9167), .ZN(n11005) );
  NOR3_X1 U8886 ( .A1(n7700), .A2(n7861), .A3(n11005), .ZN(n10689) );
  INV_X1 U8887 ( .A(n10689), .ZN(n7701) );
  OAI22_X1 U8888 ( .A1(n7701), .A2(n5073), .B1(n10907), .B2(n10624), .ZN(n7702) );
  OAI21_X1 U8889 ( .B1(n10692), .B2(n7702), .A(n5074), .ZN(n7704) );
  AOI22_X1 U8890 ( .A1(n10432), .A2(n6736), .B1(n10439), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7703) );
  OAI211_X1 U8891 ( .C1(n10381), .C2(n10687), .A(n7704), .B(n7703), .ZN(
        P1_U3290) );
  INV_X1 U8892 ( .A(n9469), .ZN(n9459) );
  INV_X1 U8893 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7705) );
  OAI222_X1 U8894 ( .A1(n5076), .A2(n7706), .B1(n9459), .B2(P2_U3152), .C1(
        n7705), .C2(n9923), .ZN(P2_U3341) );
  INV_X1 U8895 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7707) );
  NAND2_X1 U8896 ( .A1(P2_U3152), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8163) );
  OAI21_X1 U8897 ( .B1(n10641), .B2(n7707), .A(n8163), .ZN(n7713) );
  AOI22_X1 U8898 ( .A1(n7824), .A2(n8687), .B1(P2_REG2_REG_10__SCAN_IN), .B2(
        n7828), .ZN(n7710) );
  AOI211_X1 U8899 ( .C1(n7711), .C2(n7710), .A(n7823), .B(n10642), .ZN(n7712)
         );
  AOI211_X1 U8900 ( .C1(n10649), .C2(n7824), .A(n7713), .B(n7712), .ZN(n7720)
         );
  OAI21_X1 U8901 ( .B1(n10871), .B2(n7715), .A(n7714), .ZN(n7718) );
  MUX2_X1 U8902 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7716), .S(n7824), .Z(n7717)
         );
  NAND2_X1 U8903 ( .A1(n7717), .A2(n7718), .ZN(n7827) );
  OAI211_X1 U8904 ( .C1(n7718), .C2(n7717), .A(n10652), .B(n7827), .ZN(n7719)
         );
  NAND2_X1 U8905 ( .A1(n7720), .A2(n7719), .ZN(P2_U3255) );
  INV_X1 U8906 ( .A(n7721), .ZN(n7723) );
  NOR2_X1 U8907 ( .A1(n7723), .A2(n7722), .ZN(n7724) );
  XNOR2_X1 U8908 ( .A(n7725), .B(n7724), .ZN(n7730) );
  INV_X1 U8909 ( .A(n9371), .ZN(n7902) );
  OAI21_X1 U8910 ( .B1(n9386), .B2(n7953), .A(n7726), .ZN(n7728) );
  INV_X1 U8911 ( .A(n9789), .ZN(n8013) );
  OAI22_X1 U8912 ( .A1(n8013), .A2(n9372), .B1(n9335), .B2(n10768), .ZN(n7727)
         );
  AOI211_X1 U8913 ( .C1(n7902), .C2(n9404), .A(n7728), .B(n7727), .ZN(n7729)
         );
  OAI21_X1 U8914 ( .B1(n7730), .B2(n9391), .A(n7729), .ZN(P2_U3232) );
  OAI21_X1 U8915 ( .B1(n7733), .B2(n7732), .A(n7731), .ZN(n7739) );
  INV_X1 U8916 ( .A(n9391), .ZN(n9341) );
  INV_X1 U8917 ( .A(n9384), .ZN(n7736) );
  NAND2_X1 U8918 ( .A1(n9402), .A2(n10926), .ZN(n7735) );
  NAND2_X1 U8919 ( .A1(n9403), .A2(n10924), .ZN(n7734) );
  AND2_X1 U8920 ( .A1(n7735), .A2(n7734), .ZN(n7942) );
  OAI22_X1 U8921 ( .A1(n7736), .A2(n7942), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8488), .ZN(n7738) );
  OAI22_X1 U8922 ( .A1(n9335), .A2(n10802), .B1(n7928), .B2(n9386), .ZN(n7737)
         );
  AOI211_X1 U8923 ( .C1(n7739), .C2(n9341), .A(n7738), .B(n7737), .ZN(n7740)
         );
  INV_X1 U8924 ( .A(n7740), .ZN(P2_U3229) );
  NAND2_X1 U8925 ( .A1(n7742), .A2(n7741), .ZN(n7748) );
  INV_X1 U8926 ( .A(n7743), .ZN(n7745) );
  AOI21_X1 U8927 ( .B1(n7746), .B2(n7745), .A(n7744), .ZN(n7747) );
  XOR2_X1 U8928 ( .A(n7748), .B(n7747), .Z(n7753) );
  NOR2_X1 U8929 ( .A1(n9335), .A2(n10730), .ZN(n7750) );
  OAI22_X1 U8930 ( .A1(n8147), .A2(n9372), .B1(n9371), .B2(n8148), .ZN(n7749)
         );
  AOI211_X1 U8931 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(n7751), .A(n7750), .B(
        n7749), .ZN(n7752) );
  OAI21_X1 U8932 ( .B1(n7753), .B2(n9391), .A(n7752), .ZN(P2_U3239) );
  INV_X1 U8933 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7754) );
  NOR2_X1 U8934 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7754), .ZN(n8913) );
  AOI211_X1 U8935 ( .C1(n7757), .C2(n7756), .A(n10627), .B(n7755), .ZN(n7758)
         );
  AOI211_X1 U8936 ( .C1(n10670), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n8913), .B(
        n7758), .ZN(n7765) );
  OAI21_X1 U8937 ( .B1(n7761), .B2(n7760), .A(n7759), .ZN(n7762) );
  AOI22_X1 U8938 ( .A1(n7763), .A2(n10151), .B1(n10662), .B2(n7762), .ZN(n7764) );
  NAND2_X1 U8939 ( .A1(n7765), .A2(n7764), .ZN(P1_U3253) );
  NAND2_X1 U8940 ( .A1(n7769), .A2(n7768), .ZN(n7794) );
  NOR2_X1 U8941 ( .A1(n7794), .A2(n7924), .ZN(n7770) );
  AND2_X2 U8942 ( .A1(n7926), .A2(n7770), .ZN(n10998) );
  OAI21_X1 U8943 ( .B1(n9407), .B2(n7771), .A(n10703), .ZN(n7773) );
  NAND2_X1 U8944 ( .A1(n9407), .A2(n7771), .ZN(n7772) );
  AND2_X1 U8945 ( .A1(n7773), .A2(n7772), .ZN(n8146) );
  NAND2_X1 U8946 ( .A1(n8146), .A2(n8145), .ZN(n8144) );
  NAND2_X1 U8947 ( .A1(n7778), .A2(n10730), .ZN(n7774) );
  NAND2_X1 U8948 ( .A1(n8144), .A2(n7774), .ZN(n7775) );
  NAND2_X1 U8949 ( .A1(n7775), .A2(n7779), .ZN(n7921) );
  OAI21_X1 U8950 ( .B1(n7775), .B2(n7779), .A(n7921), .ZN(n7788) );
  INV_X1 U8951 ( .A(n7788), .ZN(n8745) );
  XNOR2_X1 U8952 ( .A(n7927), .B(n7776), .ZN(n7777) );
  NAND2_X1 U8953 ( .A1(n7777), .A2(n9742), .ZN(n9813) );
  INV_X1 U8954 ( .A(n9813), .ZN(n8682) );
  OAI22_X1 U8955 ( .A1(n7815), .A2(n9720), .B1(n7778), .B2(n9774), .ZN(n7787)
         );
  XNOR2_X1 U8956 ( .A(n7780), .B(n7779), .ZN(n7785) );
  NAND2_X1 U8957 ( .A1(n7782), .A2(n7781), .ZN(n7784) );
  NOR2_X1 U8958 ( .A1(n7785), .A2(n9717), .ZN(n7786) );
  AOI211_X1 U8959 ( .C1(n8682), .C2(n7788), .A(n7787), .B(n7786), .ZN(n8749)
         );
  NAND2_X1 U8960 ( .A1(n10711), .A2(n10699), .ZN(n10698) );
  INV_X1 U8961 ( .A(n8152), .ZN(n7789) );
  NAND2_X1 U8962 ( .A1(n8152), .A2(n8743), .ZN(n7931) );
  INV_X1 U8963 ( .A(n7931), .ZN(n7955) );
  AOI21_X1 U8964 ( .B1(n7790), .B2(n7789), .A(n7955), .ZN(n8741) );
  NAND2_X1 U8965 ( .A1(n6286), .A2(n10679), .ZN(n10991) );
  INV_X1 U8966 ( .A(n10991), .ZN(n10930) );
  AOI22_X1 U8967 ( .A1(n8741), .A2(n10930), .B1(n10851), .B2(n7790), .ZN(n7791) );
  OAI211_X1 U8968 ( .C1(n8745), .C2(n10729), .A(n8749), .B(n7791), .ZN(n7796)
         );
  NAND2_X1 U8969 ( .A1(n7796), .A2(n10998), .ZN(n7792) );
  OAI21_X1 U8970 ( .B1(n10998), .B2(n7375), .A(n7792), .ZN(P2_U3523) );
  INV_X1 U8971 ( .A(n7924), .ZN(n7793) );
  NOR2_X1 U8972 ( .A1(n7794), .A2(n7793), .ZN(n7795) );
  AND2_X2 U8973 ( .A1(n7926), .A2(n7795), .ZN(n11002) );
  INV_X1 U8974 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7798) );
  NAND2_X1 U8975 ( .A1(n7796), .A2(n11002), .ZN(n7797) );
  OAI21_X1 U8976 ( .B1(n11002), .B2(n7798), .A(n7797), .ZN(P2_U3460) );
  NOR2_X1 U8977 ( .A1(n7799), .A2(n9186), .ZN(n7800) );
  INV_X1 U8978 ( .A(n10902), .ZN(n10435) );
  AOI21_X1 U8979 ( .B1(n10435), .B2(n10905), .A(n7801), .ZN(n7803) );
  OAI22_X1 U8980 ( .A1(n5074), .A2(n6705), .B1(n8622), .B2(n10907), .ZN(n7802)
         );
  NOR2_X1 U8981 ( .A1(n7803), .A2(n7802), .ZN(n7804) );
  OAI21_X1 U8982 ( .B1(n10439), .B2(n7805), .A(n7804), .ZN(P1_U3291) );
  OAI21_X1 U8983 ( .B1(n7808), .B2(n7807), .A(n7806), .ZN(n7813) );
  AOI22_X1 U8984 ( .A1(n10081), .A2(n7642), .B1(n10086), .B2(n10102), .ZN(
        n7811) );
  AOI21_X1 U8985 ( .B1(n10069), .B2(n9093), .A(n7809), .ZN(n7810) );
  OAI211_X1 U8986 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n10083), .A(n7811), .B(
        n7810), .ZN(n7812) );
  AOI21_X1 U8987 ( .B1(n7813), .B2(n10078), .A(n7812), .ZN(n7814) );
  INV_X1 U8988 ( .A(n7814), .ZN(P1_U3216) );
  INV_X1 U8989 ( .A(n9386), .ZN(n8903) );
  MUX2_X1 U8990 ( .A(n8903), .B(P2_U3152), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n7817) );
  OAI22_X1 U8991 ( .A1(n7815), .A2(n9372), .B1(n9335), .B2(n8743), .ZN(n7816)
         );
  AOI211_X1 U8992 ( .C1(n7902), .C2(n9405), .A(n7817), .B(n7816), .ZN(n7822)
         );
  OAI211_X1 U8993 ( .C1(n7820), .C2(n7819), .A(n7818), .B(n9341), .ZN(n7821)
         );
  NAND2_X1 U8994 ( .A1(n7822), .A2(n7821), .ZN(P2_U3220) );
  AOI22_X1 U8995 ( .A1(n8038), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n5933), .B2(
        n7835), .ZN(n7826) );
  NAND2_X1 U8996 ( .A1(n7825), .A2(n7826), .ZN(n8037) );
  OAI21_X1 U8997 ( .B1(n7826), .B2(n7825), .A(n8037), .ZN(n7837) );
  OAI21_X1 U8998 ( .B1(n7828), .B2(n7716), .A(n7827), .ZN(n7831) );
  MUX2_X1 U8999 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n7829), .S(n8038), .Z(n7830)
         );
  NAND2_X1 U9000 ( .A1(n7830), .A2(n7831), .ZN(n8030) );
  OAI211_X1 U9001 ( .C1(n7831), .C2(n7830), .A(n10652), .B(n8030), .ZN(n7834)
         );
  NOR2_X1 U9002 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8663), .ZN(n7832) );
  AOI21_X1 U9003 ( .B1(n9487), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7832), .ZN(
        n7833) );
  OAI211_X1 U9004 ( .C1(n9490), .C2(n7835), .A(n7834), .B(n7833), .ZN(n7836)
         );
  AOI21_X1 U9005 ( .B1(n9474), .B2(n7837), .A(n7836), .ZN(n7838) );
  INV_X1 U9006 ( .A(n7838), .ZN(P2_U3256) );
  AOI22_X1 U9007 ( .A1(n10146), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n7839), .ZN(n7840) );
  OAI21_X1 U9008 ( .B1(n7843), .B2(n8088), .A(n7840), .ZN(P1_U3335) );
  AOI22_X1 U9009 ( .A1(n9479), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n7841), .ZN(n7842) );
  OAI21_X1 U9010 ( .B1(n7843), .B2(n5076), .A(n7842), .ZN(P2_U3340) );
  NAND2_X1 U9011 ( .A1(n5126), .A2(n7844), .ZN(n7845) );
  XNOR2_X1 U9012 ( .A(n7846), .B(n7845), .ZN(n7851) );
  AOI22_X1 U9013 ( .A1(n10081), .A2(n10103), .B1(n10086), .B2(n10101), .ZN(
        n7850) );
  NOR2_X1 U9014 ( .A1(n10083), .A2(n7888), .ZN(n7847) );
  AOI211_X1 U9015 ( .C1(n7893), .C2(n10069), .A(n7848), .B(n7847), .ZN(n7849)
         );
  OAI211_X1 U9016 ( .C1(n7851), .C2(n10071), .A(n7850), .B(n7849), .ZN(
        P1_U3228) );
  OAI21_X1 U9017 ( .B1(n7854), .B2(n7853), .A(n7852), .ZN(n7859) );
  OAI22_X1 U9018 ( .A1(n8019), .A2(n9372), .B1(n9335), .B2(n10819), .ZN(n7858)
         );
  NAND2_X1 U9019 ( .A1(n7902), .A2(n9789), .ZN(n7856) );
  OAI211_X1 U9020 ( .C1(n9386), .C2(n9794), .A(n7856), .B(n7855), .ZN(n7857)
         );
  AOI211_X1 U9021 ( .C1(n7859), .C2(n9341), .A(n7858), .B(n7857), .ZN(n7860)
         );
  INV_X1 U9022 ( .A(n7860), .ZN(P2_U3241) );
  NAND2_X1 U9023 ( .A1(n7861), .A2(n7643), .ZN(n7862) );
  NAND2_X1 U9024 ( .A1(n7862), .A2(n7866), .ZN(n7863) );
  OAI211_X1 U9025 ( .C1(n7643), .C2(n6736), .A(n7863), .B(n7873), .ZN(n7879)
         );
  XNOR2_X1 U9026 ( .A(n7879), .B(n9127), .ZN(n10724) );
  NAND2_X1 U9027 ( .A1(n5074), .A2(n7864), .ZN(n10751) );
  NAND2_X1 U9028 ( .A1(n9128), .A2(n7865), .ZN(n7868) );
  NAND2_X1 U9029 ( .A1(n7866), .A2(n6736), .ZN(n7867) );
  XNOR2_X1 U9030 ( .A(n9088), .B(n9127), .ZN(n7869) );
  NAND2_X1 U9031 ( .A1(n7869), .A2(n10892), .ZN(n7871) );
  AOI22_X1 U9032 ( .A1(n10405), .A2(n6735), .B1(n10103), .B2(n10398), .ZN(
        n7870) );
  OAI211_X1 U9033 ( .C1(n10724), .C2(n10895), .A(n7871), .B(n7870), .ZN(n10726) );
  MUX2_X1 U9034 ( .A(n10726), .B(P1_REG2_REG_2__SCAN_IN), .S(n10439), .Z(n7872) );
  INV_X1 U9035 ( .A(n7872), .ZN(n7877) );
  AND2_X1 U9036 ( .A1(n7873), .A2(n10720), .ZN(n7874) );
  NOR2_X1 U9037 ( .A1(n10740), .A2(n7874), .ZN(n10722) );
  INV_X1 U9038 ( .A(n10720), .ZN(n7880) );
  OAI22_X1 U9039 ( .A1(n10905), .A2(n7880), .B1(n10907), .B2(n10657), .ZN(
        n7875) );
  AOI21_X1 U9040 ( .B1(n10902), .B2(n10722), .A(n7875), .ZN(n7876) );
  OAI211_X1 U9041 ( .C1(n10724), .C2(n10751), .A(n7877), .B(n7876), .ZN(
        P1_U3289) );
  INV_X1 U9042 ( .A(n9127), .ZN(n7878) );
  NAND2_X1 U9043 ( .A1(n7879), .A2(n7878), .ZN(n7882) );
  NAND2_X1 U9044 ( .A1(n10743), .A2(n7880), .ZN(n7881) );
  NAND2_X1 U9045 ( .A1(n7882), .A2(n7881), .ZN(n10738) );
  XNOR2_X1 U9046 ( .A(n10103), .B(n9093), .ZN(n9123) );
  INV_X1 U9047 ( .A(n9123), .ZN(n10741) );
  NAND2_X1 U9048 ( .A1(n10738), .A2(n10741), .ZN(n7884) );
  INV_X1 U9049 ( .A(n10103), .ZN(n9094) );
  INV_X1 U9050 ( .A(n9093), .ZN(n10755) );
  NAND2_X1 U9051 ( .A1(n9094), .A2(n10755), .ZN(n7883) );
  NAND2_X1 U9052 ( .A1(n7884), .A2(n7883), .ZN(n7986) );
  NAND2_X1 U9053 ( .A1(n10783), .A2(n7893), .ZN(n9096) );
  INV_X1 U9054 ( .A(n7893), .ZN(n10762) );
  NAND2_X1 U9055 ( .A1(n10102), .A2(n10762), .ZN(n9091) );
  NAND2_X1 U9056 ( .A1(n9096), .A2(n9091), .ZN(n9122) );
  XNOR2_X1 U9057 ( .A(n7986), .B(n9122), .ZN(n10766) );
  INV_X1 U9058 ( .A(n10766), .ZN(n7896) );
  NAND2_X1 U9059 ( .A1(n10743), .A2(n10720), .ZN(n9086) );
  NAND2_X1 U9060 ( .A1(n9094), .A2(n9093), .ZN(n9089) );
  XNOR2_X1 U9061 ( .A(n9122), .B(n7981), .ZN(n7887) );
  INV_X1 U9062 ( .A(n10895), .ZN(n10745) );
  INV_X1 U9063 ( .A(n10101), .ZN(n7982) );
  OAI22_X1 U9064 ( .A1(n7982), .A2(n10887), .B1(n9094), .B2(n10889), .ZN(n7885) );
  AOI21_X1 U9065 ( .B1(n10766), .B2(n10745), .A(n7885), .ZN(n7886) );
  OAI21_X1 U9066 ( .B1(n7887), .B2(n10784), .A(n7886), .ZN(n10764) );
  NAND2_X1 U9067 ( .A1(n10764), .A2(n5074), .ZN(n7895) );
  OAI22_X1 U9068 ( .A1(n5074), .A2(n7889), .B1(n7888), .B2(n10907), .ZN(n7892)
         );
  NAND2_X1 U9069 ( .A1(n10740), .A2(n10755), .ZN(n10739) );
  NAND2_X1 U9070 ( .A1(n10739), .A2(n7893), .ZN(n7890) );
  NAND2_X1 U9071 ( .A1(n10776), .A2(n7890), .ZN(n10763) );
  NOR2_X1 U9072 ( .A1(n10763), .A2(n10435), .ZN(n7891) );
  AOI211_X1 U9073 ( .C1(n10432), .C2(n7893), .A(n7892), .B(n7891), .ZN(n7894)
         );
  OAI211_X1 U9074 ( .C1(n7896), .C2(n10751), .A(n7895), .B(n7894), .ZN(
        P1_U3287) );
  XNOR2_X1 U9075 ( .A(n7898), .B(n7897), .ZN(n7904) );
  OAI21_X1 U9076 ( .B1(n9386), .B2(n8052), .A(n7899), .ZN(n7901) );
  OAI22_X1 U9077 ( .A1(n8648), .A2(n9372), .B1(n9335), .B2(n10834), .ZN(n7900)
         );
  AOI211_X1 U9078 ( .C1(n7902), .C2(n9402), .A(n7901), .B(n7900), .ZN(n7903)
         );
  OAI21_X1 U9079 ( .B1(n7904), .B2(n9391), .A(n7903), .ZN(P2_U3215) );
  AND2_X1 U9080 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10031) );
  AOI211_X1 U9081 ( .C1(n7907), .C2(n7906), .A(n10627), .B(n7905), .ZN(n7908)
         );
  AOI211_X1 U9082 ( .C1(n10670), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n10031), .B(
        n7908), .ZN(n7915) );
  OAI21_X1 U9083 ( .B1(n7911), .B2(n7910), .A(n7909), .ZN(n7912) );
  AOI22_X1 U9084 ( .A1(n7913), .A2(n10151), .B1(n10662), .B2(n7912), .ZN(n7914) );
  NAND2_X1 U9085 ( .A1(n7915), .A2(n7914), .ZN(P1_U3254) );
  INV_X1 U9086 ( .A(n7916), .ZN(n7918) );
  INV_X1 U9087 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7917) );
  OAI222_X1 U9088 ( .A1(n10289), .A2(P1_U3084), .B1(n8088), .B2(n7918), .C1(
        n7917), .C2(n10546), .ZN(P1_U3334) );
  INV_X1 U9089 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7919) );
  OAI222_X1 U9090 ( .A1(n9923), .A2(n7919), .B1(n5076), .B2(n7918), .C1(n9742), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  NAND2_X1 U9091 ( .A1(n8147), .A2(n8743), .ZN(n7920) );
  XNOR2_X1 U9092 ( .A(n8011), .B(n8012), .ZN(n10805) );
  INV_X1 U9093 ( .A(n10805), .ZN(n7946) );
  AND2_X1 U9094 ( .A1(n7924), .A2(n7923), .ZN(n7925) );
  NAND2_X1 U9095 ( .A1(n7926), .A2(n7925), .ZN(n7956) );
  OR2_X1 U9096 ( .A1(n7927), .A2(n9742), .ZN(n8156) );
  NAND2_X1 U9097 ( .A1(n9813), .A2(n8156), .ZN(n10945) );
  NAND2_X1 U9098 ( .A1(n10947), .A2(n10945), .ZN(n10706) );
  NAND2_X1 U9099 ( .A1(n10947), .A2(n5182), .ZN(n10705) );
  OAI22_X1 U9100 ( .A1(n10947), .A2(n7929), .B1(n7928), .B2(n10700), .ZN(n7934) );
  AND2_X1 U9101 ( .A1(n10947), .A2(n9742), .ZN(n9593) );
  INV_X1 U9102 ( .A(n9593), .ZN(n8027) );
  AOI21_X1 U9103 ( .B1(n7954), .B2(n7935), .A(n10991), .ZN(n7932) );
  NAND2_X1 U9104 ( .A1(n7932), .A2(n9791), .ZN(n10801) );
  NOR2_X1 U9105 ( .A1(n8027), .A2(n10801), .ZN(n7933) );
  AOI211_X1 U9106 ( .C1(n9797), .C2(n7935), .A(n7934), .B(n7933), .ZN(n7945)
         );
  NAND2_X1 U9107 ( .A1(n7936), .A2(n7939), .ZN(n7938) );
  NAND2_X1 U9108 ( .A1(n7938), .A2(n7937), .ZN(n7941) );
  NAND3_X1 U9109 ( .A1(n7936), .A2(n8011), .A3(n7939), .ZN(n7940) );
  NAND3_X1 U9110 ( .A1(n7941), .A2(n10929), .A3(n7940), .ZN(n7943) );
  NAND2_X1 U9111 ( .A1(n7943), .A2(n7942), .ZN(n10803) );
  NAND2_X1 U9112 ( .A1(n10803), .A2(n10947), .ZN(n7944) );
  OAI211_X1 U9113 ( .C1(n7946), .C2(n10706), .A(n7945), .B(n7944), .ZN(
        P2_U3291) );
  INV_X2 U9114 ( .A(n10947), .ZN(n10949) );
  INV_X1 U9115 ( .A(n7951), .ZN(n7947) );
  OAI211_X1 U9116 ( .C1(n5190), .C2(n7947), .A(n7936), .B(n10929), .ZN(n7949)
         );
  AOI22_X1 U9117 ( .A1(n9404), .A2(n10924), .B1(n10926), .B2(n9789), .ZN(n7948) );
  NAND2_X1 U9118 ( .A1(n7949), .A2(n7948), .ZN(n10770) );
  INV_X1 U9119 ( .A(n10770), .ZN(n7964) );
  INV_X1 U9120 ( .A(n10706), .ZN(n9800) );
  OAI21_X1 U9121 ( .B1(n7952), .B2(n7951), .A(n7950), .ZN(n10772) );
  NOR2_X1 U9122 ( .A1(n7953), .A2(n10700), .ZN(n7960) );
  OAI21_X1 U9123 ( .B1(n7955), .B2(n10768), .A(n7954), .ZN(n10769) );
  INV_X1 U9124 ( .A(n7956), .ZN(n7958) );
  NAND2_X1 U9125 ( .A1(n7958), .A2(n7957), .ZN(n10702) );
  NOR2_X1 U9126 ( .A1(n10769), .A2(n10702), .ZN(n7959) );
  AOI211_X1 U9127 ( .C1(n10949), .C2(P2_REG2_REG_4__SCAN_IN), .A(n7960), .B(
        n7959), .ZN(n7961) );
  OAI21_X1 U9128 ( .B1(n10768), .B2(n10705), .A(n7961), .ZN(n7962) );
  AOI21_X1 U9129 ( .B1(n9800), .B2(n10772), .A(n7962), .ZN(n7963) );
  OAI21_X1 U9130 ( .B1(n10949), .B2(n7964), .A(n7963), .ZN(P2_U3292) );
  OAI21_X1 U9131 ( .B1(n7967), .B2(n7966), .A(n7965), .ZN(n7968) );
  INV_X1 U9132 ( .A(n7968), .ZN(n7980) );
  OAI21_X1 U9133 ( .B1(n7971), .B2(n7970), .A(n7969), .ZN(n7978) );
  NOR2_X1 U9134 ( .A1(n10659), .A2(n7972), .ZN(n7977) );
  INV_X1 U9135 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7974) );
  OR2_X1 U9136 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7973), .ZN(n9932) );
  OAI21_X1 U9137 ( .B1(n7975), .B2(n7974), .A(n9932), .ZN(n7976) );
  AOI211_X1 U9138 ( .C1(n7978), .C2(n10662), .A(n7977), .B(n7976), .ZN(n7979)
         );
  OAI21_X1 U9139 ( .B1(n7980), .B2(n10627), .A(n7979), .ZN(P1_U3255) );
  NAND2_X1 U9140 ( .A1(n7982), .A2(n10792), .ZN(n9095) );
  INV_X1 U9141 ( .A(n10792), .ZN(n10780) );
  NAND2_X1 U9142 ( .A1(n10101), .A2(n10780), .ZN(n9098) );
  NAND2_X1 U9143 ( .A1(n9095), .A2(n9098), .ZN(n10781) );
  NAND2_X1 U9144 ( .A1(n10786), .A2(n8105), .ZN(n9102) );
  INV_X1 U9145 ( .A(n8105), .ZN(n10811) );
  NAND2_X1 U9146 ( .A1(n10100), .A2(n10811), .ZN(n8173) );
  INV_X1 U9147 ( .A(n9125), .ZN(n8966) );
  XNOR2_X1 U9148 ( .A(n8963), .B(n8966), .ZN(n7983) );
  NAND2_X1 U9149 ( .A1(n7983), .A2(n10892), .ZN(n7985) );
  AOI22_X1 U9150 ( .A1(n10405), .A2(n10101), .B1(n10099), .B2(n10398), .ZN(
        n7984) );
  NAND2_X1 U9151 ( .A1(n7985), .A2(n7984), .ZN(n10813) );
  INV_X1 U9152 ( .A(n10813), .ZN(n8002) );
  NAND2_X1 U9153 ( .A1(n7986), .A2(n9122), .ZN(n7988) );
  NAND2_X1 U9154 ( .A1(n10783), .A2(n10762), .ZN(n7987) );
  NAND2_X1 U9155 ( .A1(n7988), .A2(n7987), .ZN(n10775) );
  INV_X1 U9156 ( .A(n10775), .ZN(n7989) );
  NAND2_X1 U9157 ( .A1(n10101), .A2(n10792), .ZN(n7990) );
  NAND2_X1 U9158 ( .A1(n7991), .A2(n7990), .ZN(n7992) );
  NAND2_X1 U9159 ( .A1(n7992), .A2(n9125), .ZN(n7993) );
  NAND2_X1 U9160 ( .A1(n8121), .A2(n7993), .ZN(n10808) );
  INV_X1 U9161 ( .A(n10381), .ZN(n10437) );
  INV_X1 U9162 ( .A(n8128), .ZN(n7995) );
  AOI21_X1 U9163 ( .B1(n10777), .B2(n8105), .A(n11005), .ZN(n7994) );
  NAND2_X1 U9164 ( .A1(n7995), .A2(n7994), .ZN(n10809) );
  NOR2_X1 U9165 ( .A1(n7996), .A2(n5073), .ZN(n10373) );
  INV_X1 U9166 ( .A(n10373), .ZN(n10410) );
  OAI22_X1 U9167 ( .A1(n5074), .A2(n7997), .B1(n8102), .B2(n10907), .ZN(n7998)
         );
  AOI21_X1 U9168 ( .B1(n10432), .B2(n8105), .A(n7998), .ZN(n7999) );
  OAI21_X1 U9169 ( .B1(n10809), .B2(n10410), .A(n7999), .ZN(n8000) );
  AOI21_X1 U9170 ( .B1(n10808), .B2(n10437), .A(n8000), .ZN(n8001) );
  OAI21_X1 U9171 ( .B1(n8002), .B2(n10439), .A(n8001), .ZN(P1_U3285) );
  NAND2_X1 U9172 ( .A1(n8045), .A2(n8003), .ZN(n8005) );
  AND2_X1 U9173 ( .A1(n8005), .A2(n8004), .ZN(n8007) );
  XNOR2_X1 U9174 ( .A(n8007), .B(n8006), .ZN(n8009) );
  NAND2_X1 U9175 ( .A1(n9788), .A2(n10924), .ZN(n8008) );
  OAI21_X1 U9176 ( .B1(n8677), .B2(n9720), .A(n8008), .ZN(n8109) );
  AOI21_X1 U9177 ( .B1(n8009), .B2(n10929), .A(n8109), .ZN(n10856) );
  NAND2_X1 U9178 ( .A1(n9792), .A2(n10834), .ZN(n8051) );
  AOI21_X1 U9179 ( .B1(n8051), .B2(n10852), .A(n10991), .ZN(n8010) );
  OR2_X2 U9180 ( .A1(n8051), .A2(n10852), .ZN(n8683) );
  NAND2_X1 U9181 ( .A1(n8010), .A2(n8683), .ZN(n10854) );
  NAND2_X1 U9182 ( .A1(n8013), .A2(n10802), .ZN(n8014) );
  NAND2_X1 U9183 ( .A1(n8022), .A2(n8021), .ZN(n10849) );
  NAND3_X1 U9184 ( .A1(n10850), .A2(n10849), .A3(n9800), .ZN(n8026) );
  OAI22_X1 U9185 ( .A1(n10947), .A2(n8023), .B1(n8113), .B2(n10700), .ZN(n8024) );
  AOI21_X1 U9186 ( .B1(n9797), .B2(n10852), .A(n8024), .ZN(n8025) );
  OAI211_X1 U9187 ( .C1(n8027), .C2(n10854), .A(n8026), .B(n8025), .ZN(n8028)
         );
  INV_X1 U9188 ( .A(n8028), .ZN(n8029) );
  OAI21_X1 U9189 ( .B1(n10856), .B2(n10949), .A(n8029), .ZN(P2_U3288) );
  INV_X1 U9190 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n8036) );
  INV_X1 U9191 ( .A(n8030), .ZN(n8031) );
  AOI21_X1 U9192 ( .B1(n8038), .B2(P2_REG1_REG_11__SCAN_IN), .A(n8031), .ZN(
        n8033) );
  INV_X1 U9193 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10963) );
  MUX2_X1 U9194 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n10963), .S(n8072), .Z(n8032) );
  AND2_X1 U9195 ( .A1(n8033), .A2(n8032), .ZN(n8076) );
  NOR2_X1 U9196 ( .A1(n8033), .A2(n8032), .ZN(n8034) );
  OAI21_X1 U9197 ( .B1(n8076), .B2(n8034), .A(n10652), .ZN(n8035) );
  NAND2_X1 U9198 ( .A1(P2_U3152), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8779) );
  OAI211_X1 U9199 ( .C1(n10641), .C2(n8036), .A(n8035), .B(n8779), .ZN(n8042)
         );
  OAI21_X1 U9200 ( .B1(n8038), .B2(P2_REG2_REG_11__SCAN_IN), .A(n8037), .ZN(
        n8040) );
  XNOR2_X1 U9201 ( .A(n8072), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n8039) );
  NOR2_X1 U9202 ( .A1(n8039), .A2(n8040), .ZN(n8071) );
  AOI211_X1 U9203 ( .C1(n8040), .C2(n8039), .A(n8071), .B(n10642), .ZN(n8041)
         );
  AOI211_X1 U9204 ( .C1(n10649), .C2(n8072), .A(n8042), .B(n8041), .ZN(n8043)
         );
  INV_X1 U9205 ( .A(n8043), .ZN(P2_U3257) );
  NAND2_X1 U9206 ( .A1(n8045), .A2(n8044), .ZN(n8046) );
  XNOR2_X1 U9207 ( .A(n8046), .B(n8049), .ZN(n8047) );
  OAI222_X1 U9208 ( .A1(n9720), .A2(n8648), .B1(n9774), .B2(n8048), .C1(n9717), 
        .C2(n8047), .ZN(n10836) );
  INV_X1 U9209 ( .A(n10836), .ZN(n8059) );
  OAI21_X1 U9210 ( .B1(n5189), .B2(n5686), .A(n8050), .ZN(n10838) );
  OAI21_X1 U9211 ( .B1(n9792), .B2(n10834), .A(n8051), .ZN(n10835) );
  OAI22_X1 U9212 ( .A1(n10947), .A2(n8053), .B1(n8052), .B2(n10700), .ZN(n8054) );
  AOI21_X1 U9213 ( .B1(n9797), .B2(n8055), .A(n8054), .ZN(n8056) );
  OAI21_X1 U9214 ( .B1(n10835), .B2(n10702), .A(n8056), .ZN(n8057) );
  AOI21_X1 U9215 ( .B1(n10838), .B2(n9800), .A(n8057), .ZN(n8058) );
  OAI21_X1 U9216 ( .B1(n8059), .B2(n10949), .A(n8058), .ZN(P2_U3289) );
  OAI22_X1 U9217 ( .A1(n10677), .A2(n9717), .B1(n8148), .B2(n9720), .ZN(n8060)
         );
  INV_X1 U9218 ( .A(n8060), .ZN(n10683) );
  INV_X1 U9219 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n8061) );
  OAI22_X1 U9220 ( .A1(n10683), .A2(n10949), .B1(n8061), .B2(n10700), .ZN(
        n8062) );
  AOI21_X1 U9221 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n10949), .A(n8062), .ZN(
        n8064) );
  INV_X1 U9222 ( .A(n10702), .ZN(n9763) );
  OAI21_X1 U9223 ( .B1(n9797), .B2(n9763), .A(n10680), .ZN(n8063) );
  OAI211_X1 U9224 ( .C1(n10677), .C2(n10706), .A(n8064), .B(n8063), .ZN(
        P2_U3296) );
  OAI222_X1 U9225 ( .A1(n5076), .A2(n8070), .B1(n8066), .B2(P2_U3152), .C1(
        n8065), .C2(n9923), .ZN(P2_U3337) );
  INV_X1 U9226 ( .A(n8067), .ZN(n8087) );
  OAI222_X1 U9227 ( .A1(n5076), .A2(n8087), .B1(P2_U3152), .B2(n6286), .C1(
        n8068), .C2(n9923), .ZN(P2_U3338) );
  OAI222_X1 U9228 ( .A1(P1_U3084), .A2(n9172), .B1(n8088), .B2(n8070), .C1(
        n8069), .C2(n10546), .ZN(P1_U3332) );
  AOI21_X1 U9229 ( .B1(n8072), .B2(P2_REG2_REG_12__SCAN_IN), .A(n8071), .ZN(
        n8074) );
  AOI22_X1 U9230 ( .A1(n8192), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8852), .B2(
        n8188), .ZN(n8073) );
  NAND2_X1 U9231 ( .A1(n8074), .A2(n8073), .ZN(n8191) );
  OAI21_X1 U9232 ( .B1(n8074), .B2(n8073), .A(n8191), .ZN(n8075) );
  NAND2_X1 U9233 ( .A1(n8075), .A2(n9474), .ZN(n8085) );
  AOI21_X1 U9234 ( .B1(n10963), .B2(n8077), .A(n8076), .ZN(n8079) );
  AOI22_X1 U9235 ( .A1(n8192), .A2(n5971), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n8188), .ZN(n8078) );
  NOR2_X1 U9236 ( .A1(n8079), .A2(n8078), .ZN(n8187) );
  AOI21_X1 U9237 ( .B1(n8079), .B2(n8078), .A(n8187), .ZN(n8080) );
  NOR2_X1 U9238 ( .A1(n8080), .A2(n9464), .ZN(n8083) );
  INV_X1 U9239 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8081) );
  NOR2_X1 U9240 ( .A1(n10641), .A2(n8081), .ZN(n8082) );
  AND2_X1 U9241 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8803) );
  NOR3_X1 U9242 ( .A1(n8083), .A2(n8082), .A3(n8803), .ZN(n8084) );
  OAI211_X1 U9243 ( .C1(n9490), .C2(n8188), .A(n8085), .B(n8084), .ZN(P2_U3258) );
  OAI222_X1 U9244 ( .A1(P1_U3084), .A2(n9112), .B1(n8088), .B2(n8087), .C1(
        n8086), .C2(n8845), .ZN(P1_U3333) );
  NAND2_X1 U9245 ( .A1(n8090), .A2(n8089), .ZN(n8091) );
  XOR2_X1 U9246 ( .A(n8092), .B(n8091), .Z(n8097) );
  AOI22_X1 U9247 ( .A1(n10081), .A2(n10102), .B1(n10086), .B2(n10100), .ZN(
        n8096) );
  NOR2_X1 U9248 ( .A1(n10089), .A2(n10780), .ZN(n8093) );
  AOI211_X1 U9249 ( .C1(n10789), .C2(n9930), .A(n8094), .B(n8093), .ZN(n8095)
         );
  OAI211_X1 U9250 ( .C1(n8097), .C2(n10071), .A(n8096), .B(n8095), .ZN(
        P1_U3225) );
  XOR2_X1 U9251 ( .A(n8100), .B(n8099), .Z(n8101) );
  XNOR2_X1 U9252 ( .A(n8098), .B(n8101), .ZN(n8108) );
  AOI22_X1 U9253 ( .A1(n10081), .A2(n10101), .B1(n10086), .B2(n10099), .ZN(
        n8107) );
  NOR2_X1 U9254 ( .A1(n10083), .A2(n8102), .ZN(n8103) );
  AOI211_X1 U9255 ( .C1(n8105), .C2(n10069), .A(n8104), .B(n8103), .ZN(n8106)
         );
  OAI211_X1 U9256 ( .C1(n8108), .C2(n10071), .A(n8107), .B(n8106), .ZN(
        P1_U3237) );
  NAND2_X1 U9257 ( .A1(n9384), .A2(n8109), .ZN(n8112) );
  INV_X1 U9258 ( .A(n8110), .ZN(n8111) );
  OAI211_X1 U9259 ( .C1(n9386), .C2(n8113), .A(n8112), .B(n8111), .ZN(n8118)
         );
  XNOR2_X1 U9260 ( .A(n8115), .B(n8114), .ZN(n8116) );
  NOR2_X1 U9261 ( .A1(n8116), .A2(n9391), .ZN(n8117) );
  AOI211_X1 U9262 ( .C1(n10852), .C2(n9389), .A(n8118), .B(n8117), .ZN(n8119)
         );
  INV_X1 U9263 ( .A(n8119), .ZN(P2_U3223) );
  NAND2_X1 U9264 ( .A1(n10786), .A2(n10811), .ZN(n8120) );
  INV_X1 U9265 ( .A(n10099), .ZN(n8122) );
  NAND2_X1 U9266 ( .A1(n8122), .A2(n8697), .ZN(n8969) );
  INV_X1 U9267 ( .A(n8697), .ZN(n10828) );
  NAND2_X1 U9268 ( .A1(n10099), .A2(n10828), .ZN(n8968) );
  NAND2_X1 U9269 ( .A1(n8969), .A2(n8968), .ZN(n8169) );
  XNOR2_X1 U9270 ( .A(n8170), .B(n8169), .ZN(n10831) );
  INV_X1 U9271 ( .A(n10831), .ZN(n8133) );
  NAND2_X1 U9272 ( .A1(n8174), .A2(n8173), .ZN(n8123) );
  INV_X1 U9273 ( .A(n8169), .ZN(n9129) );
  XNOR2_X1 U9274 ( .A(n8123), .B(n9129), .ZN(n8126) );
  INV_X1 U9275 ( .A(n10098), .ZN(n8636) );
  OAI22_X1 U9276 ( .A1(n10786), .A2(n10889), .B1(n8636), .B2(n10887), .ZN(
        n8124) );
  AOI21_X1 U9277 ( .B1(n10831), .B2(n10745), .A(n8124), .ZN(n8125) );
  OAI21_X1 U9278 ( .B1(n10784), .B2(n8126), .A(n8125), .ZN(n10829) );
  NAND2_X1 U9279 ( .A1(n10829), .A2(n5074), .ZN(n8132) );
  OAI22_X1 U9280 ( .A1(n5074), .A2(n8127), .B1(n8694), .B2(n10907), .ZN(n8130)
         );
  INV_X1 U9281 ( .A(n11005), .ZN(n10778) );
  OAI211_X1 U9282 ( .C1(n8128), .C2(n10828), .A(n8181), .B(n10778), .ZN(n10827) );
  NOR2_X1 U9283 ( .A1(n10827), .A2(n10410), .ZN(n8129) );
  AOI211_X1 U9284 ( .C1(n10432), .C2(n8697), .A(n8130), .B(n8129), .ZN(n8131)
         );
  OAI211_X1 U9285 ( .C1(n8133), .C2(n10751), .A(n8132), .B(n8131), .ZN(
        P1_U3284) );
  INV_X1 U9286 ( .A(n8134), .ZN(n8135) );
  AOI21_X1 U9287 ( .B1(n8137), .B2(n8136), .A(n8135), .ZN(n8142) );
  OAI21_X1 U9288 ( .B1(n9386), .B2(n8654), .A(n8138), .ZN(n8140) );
  OAI22_X1 U9289 ( .A1(n8648), .A2(n9371), .B1(n9372), .B2(n8664), .ZN(n8139)
         );
  AOI211_X1 U9290 ( .C1(n10865), .C2(n9389), .A(n8140), .B(n8139), .ZN(n8141)
         );
  OAI21_X1 U9291 ( .B1(n8142), .B2(n9391), .A(n8141), .ZN(P2_U3233) );
  OAI21_X1 U9292 ( .B1(n8146), .B2(n8145), .A(n8144), .ZN(n10734) );
  OAI22_X1 U9293 ( .A1(n8148), .A2(n9774), .B1(n8147), .B2(n9720), .ZN(n8149)
         );
  AOI21_X1 U9294 ( .B1(n10734), .B2(n8682), .A(n8149), .ZN(n8150) );
  OAI21_X1 U9295 ( .B1(n9717), .B2(n8151), .A(n8150), .ZN(n10732) );
  INV_X1 U9296 ( .A(n10732), .ZN(n8160) );
  AND2_X1 U9297 ( .A1(n10698), .A2(n8157), .ZN(n8153) );
  OR2_X1 U9298 ( .A1(n8153), .A2(n8152), .ZN(n10731) );
  OAI22_X1 U9299 ( .A1(n10702), .A2(n10731), .B1(n8154), .B2(n10700), .ZN(
        n8155) );
  AOI21_X1 U9300 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n10949), .A(n8155), .ZN(
        n8159) );
  NOR2_X1 U9301 ( .A1(n10949), .A2(n8156), .ZN(n9728) );
  AOI22_X1 U9302 ( .A1(n9728), .A2(n10734), .B1(n9797), .B2(n8157), .ZN(n8158)
         );
  OAI211_X1 U9303 ( .C1(n8160), .C2(n10949), .A(n8159), .B(n8158), .ZN(
        P2_U3294) );
  XNOR2_X1 U9304 ( .A(n8162), .B(n8161), .ZN(n8167) );
  OAI21_X1 U9305 ( .B1(n9386), .B2(n8686), .A(n8163), .ZN(n8165) );
  OAI22_X1 U9306 ( .A1(n8677), .A2(n9371), .B1(n9372), .B2(n9399), .ZN(n8164)
         );
  AOI211_X1 U9307 ( .C1(n8811), .C2(n9389), .A(n8165), .B(n8164), .ZN(n8166)
         );
  OAI21_X1 U9308 ( .B1(n8167), .B2(n9391), .A(n8166), .ZN(P2_U3219) );
  NOR2_X1 U9309 ( .A1(n10099), .A2(n8697), .ZN(n8168) );
  INV_X1 U9310 ( .A(n8637), .ZN(n10843) );
  NAND2_X1 U9311 ( .A1(n10843), .A2(n10098), .ZN(n9052) );
  NAND2_X1 U9312 ( .A1(n8636), .A2(n8637), .ZN(n8971) );
  NAND2_X1 U9313 ( .A1(n9052), .A2(n8971), .ZN(n8175) );
  NAND2_X1 U9314 ( .A1(n8171), .A2(n8175), .ZN(n8639) );
  OR2_X1 U9315 ( .A1(n8171), .A2(n8175), .ZN(n8172) );
  NAND2_X1 U9316 ( .A1(n8639), .A2(n8172), .ZN(n10842) );
  AOI22_X1 U9317 ( .A1(n10405), .A2(n10099), .B1(n10097), .B2(n10398), .ZN(
        n8179) );
  AND2_X1 U9318 ( .A1(n8968), .A2(n8173), .ZN(n9100) );
  NAND2_X1 U9319 ( .A1(n9151), .A2(n8969), .ZN(n8176) );
  INV_X1 U9320 ( .A(n8175), .ZN(n9133) );
  XNOR2_X1 U9321 ( .A(n8176), .B(n9133), .ZN(n8177) );
  NAND2_X1 U9322 ( .A1(n8177), .A2(n10892), .ZN(n8178) );
  OAI211_X1 U9323 ( .C1(n10842), .C2(n10895), .A(n8179), .B(n8178), .ZN(n10845) );
  NAND2_X1 U9324 ( .A1(n10845), .A2(n5074), .ZN(n8186) );
  INV_X1 U9325 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n8180) );
  OAI22_X1 U9326 ( .A1(n5074), .A2(n8180), .B1(n8764), .B2(n10907), .ZN(n8184)
         );
  NAND2_X1 U9327 ( .A1(n8181), .A2(n8637), .ZN(n8182) );
  NAND2_X1 U9328 ( .A1(n8640), .A2(n8182), .ZN(n10844) );
  NOR2_X1 U9329 ( .A1(n10844), .A2(n10435), .ZN(n8183) );
  AOI211_X1 U9330 ( .C1(n10432), .C2(n8637), .A(n8184), .B(n8183), .ZN(n8185)
         );
  OAI211_X1 U9331 ( .C1(n10842), .C2(n10751), .A(n8186), .B(n8185), .ZN(
        P1_U3283) );
  AOI21_X1 U9332 ( .B1(n8188), .B2(n5971), .A(n8187), .ZN(n8190) );
  AOI22_X1 U9333 ( .A1(n9410), .A2(n5994), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n9417), .ZN(n8189) );
  NOR2_X1 U9334 ( .A1(n8190), .A2(n8189), .ZN(n9416) );
  AOI21_X1 U9335 ( .B1(n8190), .B2(n8189), .A(n9416), .ZN(n8200) );
  AOI22_X1 U9336 ( .A1(n9410), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n5990), .B2(
        n9417), .ZN(n8194) );
  OAI21_X1 U9337 ( .B1(n8192), .B2(P2_REG2_REG_13__SCAN_IN), .A(n8191), .ZN(
        n8193) );
  NAND2_X1 U9338 ( .A1(n8194), .A2(n8193), .ZN(n9409) );
  OAI21_X1 U9339 ( .B1(n8194), .B2(n8193), .A(n9409), .ZN(n8195) );
  NAND2_X1 U9340 ( .A1(n8195), .A2(n9474), .ZN(n8199) );
  AND2_X1 U9341 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8901) );
  INV_X1 U9342 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8196) );
  NOR2_X1 U9343 ( .A1(n10641), .A2(n8196), .ZN(n8197) );
  AOI211_X1 U9344 ( .C1(n9410), .C2(n10649), .A(n8901), .B(n8197), .ZN(n8198)
         );
  OAI211_X1 U9345 ( .C1(n8200), .C2(n9464), .A(n8199), .B(n8198), .ZN(P2_U3259) );
  XOR2_X1 U9346 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_0), .Z(n8203) );
  XOR2_X1 U9347 ( .A(SI_31_), .B(keyinput_1), .Z(n8202) );
  XOR2_X1 U9348 ( .A(SI_30_), .B(keyinput_2), .Z(n8201) );
  AOI21_X1 U9349 ( .B1(n8203), .B2(n8202), .A(n8201), .ZN(n8208) );
  XNOR2_X1 U9350 ( .A(n8204), .B(keyinput_3), .ZN(n8207) );
  XNOR2_X1 U9351 ( .A(n8205), .B(keyinput_4), .ZN(n8206) );
  NOR3_X1 U9352 ( .A1(n8208), .A2(n8207), .A3(n8206), .ZN(n8211) );
  XNOR2_X1 U9353 ( .A(SI_27_), .B(keyinput_5), .ZN(n8210) );
  XNOR2_X1 U9354 ( .A(n8405), .B(keyinput_6), .ZN(n8209) );
  OAI21_X1 U9355 ( .B1(n8211), .B2(n8210), .A(n8209), .ZN(n8214) );
  XOR2_X1 U9356 ( .A(SI_24_), .B(keyinput_8), .Z(n8213) );
  XNOR2_X1 U9357 ( .A(SI_25_), .B(keyinput_7), .ZN(n8212) );
  NAND3_X1 U9358 ( .A1(n8214), .A2(n8213), .A3(n8212), .ZN(n8218) );
  XNOR2_X1 U9359 ( .A(n8215), .B(keyinput_9), .ZN(n8217) );
  XNOR2_X1 U9360 ( .A(SI_22_), .B(keyinput_10), .ZN(n8216) );
  AOI21_X1 U9361 ( .B1(n8218), .B2(n8217), .A(n8216), .ZN(n8221) );
  XNOR2_X1 U9362 ( .A(SI_21_), .B(keyinput_11), .ZN(n8220) );
  XNOR2_X1 U9363 ( .A(SI_20_), .B(keyinput_12), .ZN(n8219) );
  OAI21_X1 U9364 ( .B1(n8221), .B2(n8220), .A(n8219), .ZN(n8225) );
  XNOR2_X1 U9365 ( .A(n8222), .B(keyinput_13), .ZN(n8224) );
  XNOR2_X1 U9366 ( .A(SI_18_), .B(keyinput_14), .ZN(n8223) );
  AOI21_X1 U9367 ( .B1(n8225), .B2(n8224), .A(n8223), .ZN(n8230) );
  XNOR2_X1 U9368 ( .A(n8226), .B(keyinput_17), .ZN(n8229) );
  XOR2_X1 U9369 ( .A(SI_16_), .B(keyinput_16), .Z(n8228) );
  XOR2_X1 U9370 ( .A(SI_17_), .B(keyinput_15), .Z(n8227) );
  NOR4_X1 U9371 ( .A1(n8230), .A2(n8229), .A3(n8228), .A4(n8227), .ZN(n8233)
         );
  XNOR2_X1 U9372 ( .A(SI_14_), .B(keyinput_18), .ZN(n8232) );
  XOR2_X1 U9373 ( .A(SI_13_), .B(keyinput_19), .Z(n8231) );
  OAI21_X1 U9374 ( .B1(n8233), .B2(n8232), .A(n8231), .ZN(n8244) );
  XNOR2_X1 U9375 ( .A(SI_12_), .B(keyinput_20), .ZN(n8243) );
  XNOR2_X1 U9376 ( .A(n8436), .B(keyinput_24), .ZN(n8237) );
  XNOR2_X1 U9377 ( .A(n8234), .B(keyinput_25), .ZN(n8236) );
  XNOR2_X1 U9378 ( .A(SI_9_), .B(keyinput_23), .ZN(n8235) );
  NOR3_X1 U9379 ( .A1(n8237), .A2(n8236), .A3(n8235), .ZN(n8241) );
  XNOR2_X1 U9380 ( .A(n8431), .B(keyinput_22), .ZN(n8240) );
  XNOR2_X1 U9381 ( .A(n8238), .B(keyinput_21), .ZN(n8239) );
  NAND3_X1 U9382 ( .A1(n8241), .A2(n8240), .A3(n8239), .ZN(n8242) );
  AOI21_X1 U9383 ( .B1(n8244), .B2(n8243), .A(n8242), .ZN(n8251) );
  XNOR2_X1 U9384 ( .A(n8443), .B(keyinput_26), .ZN(n8248) );
  XNOR2_X1 U9385 ( .A(n8444), .B(keyinput_29), .ZN(n8247) );
  XNOR2_X1 U9386 ( .A(SI_4_), .B(keyinput_28), .ZN(n8246) );
  XNOR2_X1 U9387 ( .A(SI_5_), .B(keyinput_27), .ZN(n8245) );
  NAND4_X1 U9388 ( .A1(n8248), .A2(n8247), .A3(n8246), .A4(n8245), .ZN(n8250)
         );
  XNOR2_X1 U9389 ( .A(SI_2_), .B(keyinput_30), .ZN(n8249) );
  OAI21_X1 U9390 ( .B1(n8251), .B2(n8250), .A(n8249), .ZN(n8258) );
  XNOR2_X1 U9391 ( .A(P2_U3152), .B(keyinput_34), .ZN(n8255) );
  XNOR2_X1 U9392 ( .A(n8454), .B(keyinput_31), .ZN(n8254) );
  XNOR2_X1 U9393 ( .A(SI_0_), .B(keyinput_32), .ZN(n8253) );
  XNOR2_X1 U9394 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_33), .ZN(n8252) );
  NOR4_X1 U9395 ( .A1(n8255), .A2(n8254), .A3(n8253), .A4(n8252), .ZN(n8257)
         );
  XNOR2_X1 U9396 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_35), .ZN(n8256) );
  AOI21_X1 U9397 ( .B1(n8258), .B2(n8257), .A(n8256), .ZN(n8264) );
  XOR2_X1 U9398 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_36), .Z(n8263) );
  XNOR2_X1 U9399 ( .A(n8463), .B(keyinput_39), .ZN(n8261) );
  XNOR2_X1 U9400 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_38), .ZN(n8260) );
  XNOR2_X1 U9401 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_37), .ZN(n8259) );
  NOR3_X1 U9402 ( .A1(n8261), .A2(n8260), .A3(n8259), .ZN(n8262) );
  OAI21_X1 U9403 ( .B1(n8264), .B2(n8263), .A(n8262), .ZN(n8268) );
  XOR2_X1 U9404 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_40), .Z(n8267) );
  XNOR2_X1 U9405 ( .A(n8265), .B(keyinput_41), .ZN(n8266) );
  AOI21_X1 U9406 ( .B1(n8268), .B2(n8267), .A(n8266), .ZN(n8271) );
  XNOR2_X1 U9407 ( .A(n8473), .B(keyinput_42), .ZN(n8270) );
  XNOR2_X1 U9408 ( .A(n8474), .B(keyinput_43), .ZN(n8269) );
  NOR3_X1 U9409 ( .A1(n8271), .A2(n8270), .A3(n8269), .ZN(n8274) );
  XOR2_X1 U9410 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_44), .Z(n8273) );
  XNOR2_X1 U9411 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_45), .ZN(n8272) );
  NOR3_X1 U9412 ( .A1(n8274), .A2(n8273), .A3(n8272), .ZN(n8278) );
  XNOR2_X1 U9413 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_46), .ZN(n8277) );
  XNOR2_X1 U9414 ( .A(n8482), .B(keyinput_48), .ZN(n8276) );
  XNOR2_X1 U9415 ( .A(n8483), .B(keyinput_47), .ZN(n8275) );
  OAI211_X1 U9416 ( .C1(n8278), .C2(n8277), .A(n8276), .B(n8275), .ZN(n8285)
         );
  XNOR2_X1 U9417 ( .A(n8488), .B(keyinput_49), .ZN(n8282) );
  XNOR2_X1 U9418 ( .A(P2_REG3_REG_24__SCAN_IN), .B(keyinput_51), .ZN(n8281) );
  XNOR2_X1 U9419 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_52), .ZN(n8280) );
  XNOR2_X1 U9420 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_50), .ZN(n8279) );
  NOR4_X1 U9421 ( .A1(n8282), .A2(n8281), .A3(n8280), .A4(n8279), .ZN(n8284)
         );
  XNOR2_X1 U9422 ( .A(n8493), .B(keyinput_53), .ZN(n8283) );
  AOI21_X1 U9423 ( .B1(n8285), .B2(n8284), .A(n8283), .ZN(n8292) );
  XOR2_X1 U9424 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_54), .Z(n8291) );
  OAI22_X1 U9425 ( .A1(n8288), .A2(keyinput_56), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(keyinput_57), .ZN(n8287) );
  AND2_X1 U9426 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_57), .ZN(n8286)
         );
  AOI211_X1 U9427 ( .C1(keyinput_56), .C2(n8288), .A(n8287), .B(n8286), .ZN(
        n8290) );
  XNOR2_X1 U9428 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_55), .ZN(n8289) );
  OAI211_X1 U9429 ( .C1(n8292), .C2(n8291), .A(n8290), .B(n8289), .ZN(n8295)
         );
  XOR2_X1 U9430 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_59), .Z(n8294) );
  XNOR2_X1 U9431 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_58), .ZN(n8293) );
  NAND3_X1 U9432 ( .A1(n8295), .A2(n8294), .A3(n8293), .ZN(n8299) );
  XNOR2_X1 U9433 ( .A(n8296), .B(keyinput_60), .ZN(n8298) );
  XNOR2_X1 U9434 ( .A(n8506), .B(keyinput_61), .ZN(n8297) );
  AOI21_X1 U9435 ( .B1(n8299), .B2(n8298), .A(n8297), .ZN(n8306) );
  XOR2_X1 U9436 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_65), .Z(n8303) );
  XOR2_X1 U9437 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_64), .Z(n8302) );
  XNOR2_X1 U9438 ( .A(n8510), .B(keyinput_62), .ZN(n8301) );
  XNOR2_X1 U9439 ( .A(P2_REG3_REG_15__SCAN_IN), .B(keyinput_63), .ZN(n8300) );
  NAND4_X1 U9440 ( .A1(n8303), .A2(n8302), .A3(n8301), .A4(n8300), .ZN(n8305)
         );
  XOR2_X1 U9441 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(keyinput_66), .Z(n8304) );
  OAI21_X1 U9442 ( .B1(n8306), .B2(n8305), .A(n8304), .ZN(n8309) );
  XOR2_X1 U9443 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_68), .Z(n8308) );
  XNOR2_X1 U9444 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput_67), .ZN(n8307)
         );
  NAND3_X1 U9445 ( .A1(n8309), .A2(n8308), .A3(n8307), .ZN(n8312) );
  XNOR2_X1 U9446 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput_69), .ZN(n8311)
         );
  XOR2_X1 U9447 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(keyinput_70), .Z(n8310) );
  AOI21_X1 U9448 ( .B1(n8312), .B2(n8311), .A(n8310), .ZN(n8318) );
  XOR2_X1 U9449 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_71), .Z(n8317) );
  XOR2_X1 U9450 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput_73), .Z(n8315) );
  XOR2_X1 U9451 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_72), .Z(n8314) );
  XNOR2_X1 U9452 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_74), .ZN(n8313)
         );
  NOR3_X1 U9453 ( .A1(n8315), .A2(n8314), .A3(n8313), .ZN(n8316) );
  OAI21_X1 U9454 ( .B1(n8318), .B2(n8317), .A(n8316), .ZN(n8321) );
  XOR2_X1 U9455 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_75), .Z(n8320) );
  XNOR2_X1 U9456 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput_76), .ZN(n8319)
         );
  AOI21_X1 U9457 ( .B1(n8321), .B2(n8320), .A(n8319), .ZN(n8324) );
  XOR2_X1 U9458 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_77), .Z(n8323) );
  XOR2_X1 U9459 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_78), .Z(n8322) );
  OAI21_X1 U9460 ( .B1(n8324), .B2(n8323), .A(n8322), .ZN(n8327) );
  XOR2_X1 U9461 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(keyinput_80), .Z(n8326) );
  XNOR2_X1 U9462 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_79), .ZN(n8325)
         );
  NAND3_X1 U9463 ( .A1(n8327), .A2(n8326), .A3(n8325), .ZN(n8333) );
  XNOR2_X1 U9464 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_81), .ZN(n8332)
         );
  XOR2_X1 U9465 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput_82), .Z(n8330) );
  XNOR2_X1 U9466 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_84), .ZN(n8329)
         );
  XNOR2_X1 U9467 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_83), .ZN(n8328)
         );
  NAND3_X1 U9468 ( .A1(n8330), .A2(n8329), .A3(n8328), .ZN(n8331) );
  AOI21_X1 U9469 ( .B1(n8333), .B2(n8332), .A(n8331), .ZN(n8336) );
  XNOR2_X1 U9470 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_85), .ZN(n8335)
         );
  XNOR2_X1 U9471 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_86), .ZN(n8334)
         );
  OAI21_X1 U9472 ( .B1(n8336), .B2(n8335), .A(n8334), .ZN(n8343) );
  XNOR2_X1 U9473 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput_87), .ZN(n8342) );
  XNOR2_X1 U9474 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_91), .ZN(n8340) );
  XNOR2_X1 U9475 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_88), .ZN(n8339) );
  XNOR2_X1 U9476 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_89), .ZN(n8338) );
  XNOR2_X1 U9477 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput_90), .ZN(n8337) );
  NAND4_X1 U9478 ( .A1(n8340), .A2(n8339), .A3(n8338), .A4(n8337), .ZN(n8341)
         );
  AOI21_X1 U9479 ( .B1(n8343), .B2(n8342), .A(n8341), .ZN(n8345) );
  XNOR2_X1 U9480 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_92), .ZN(n8344) );
  NOR2_X1 U9481 ( .A1(n8345), .A2(n8344), .ZN(n8349) );
  XNOR2_X1 U9482 ( .A(n8555), .B(keyinput_95), .ZN(n8348) );
  XNOR2_X1 U9483 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_94), .ZN(n8347) );
  XNOR2_X1 U9484 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_93), .ZN(n8346) );
  NOR4_X1 U9485 ( .A1(n8349), .A2(n8348), .A3(n8347), .A4(n8346), .ZN(n8353)
         );
  XOR2_X1 U9486 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_97), .Z(n8352) );
  XOR2_X1 U9487 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_96), .Z(n8351) );
  XNOR2_X1 U9488 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_98), .ZN(n8350) );
  NOR4_X1 U9489 ( .A1(n8353), .A2(n8352), .A3(n8351), .A4(n8350), .ZN(n8356)
         );
  XNOR2_X1 U9490 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_99), .ZN(n8355) );
  XOR2_X1 U9491 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_100), .Z(n8354) );
  OAI21_X1 U9492 ( .B1(n8356), .B2(n8355), .A(n8354), .ZN(n8360) );
  XOR2_X1 U9493 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_101), .Z(n8359) );
  XNOR2_X1 U9494 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_103), .ZN(n8358) );
  XNOR2_X1 U9495 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_102), .ZN(n8357) );
  NAND4_X1 U9496 ( .A1(n8360), .A2(n8359), .A3(n8358), .A4(n8357), .ZN(n8363)
         );
  XOR2_X1 U9497 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_104), .Z(n8362) );
  XNOR2_X1 U9498 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_105), .ZN(n8361) );
  AOI21_X1 U9499 ( .B1(n8363), .B2(n8362), .A(n8361), .ZN(n8368) );
  XNOR2_X1 U9500 ( .A(n8364), .B(keyinput_108), .ZN(n8367) );
  XNOR2_X1 U9501 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_107), .ZN(n8366) );
  XNOR2_X1 U9502 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_106), .ZN(n8365) );
  NOR4_X1 U9503 ( .A1(n8368), .A2(n8367), .A3(n8366), .A4(n8365), .ZN(n8375)
         );
  XOR2_X1 U9504 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_109), .Z(n8374) );
  XNOR2_X1 U9505 ( .A(n8369), .B(keyinput_112), .ZN(n8372) );
  XNOR2_X1 U9506 ( .A(n8583), .B(keyinput_111), .ZN(n8371) );
  XNOR2_X1 U9507 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_110), .ZN(n8370) );
  NOR3_X1 U9508 ( .A1(n8372), .A2(n8371), .A3(n8370), .ZN(n8373) );
  OAI21_X1 U9509 ( .B1(n8375), .B2(n8374), .A(n8373), .ZN(n8378) );
  XNOR2_X1 U9510 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_113), .ZN(n8377) );
  XNOR2_X1 U9511 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_114), .ZN(n8376) );
  AOI21_X1 U9512 ( .B1(n8378), .B2(n8377), .A(n8376), .ZN(n8381) );
  XNOR2_X1 U9513 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_115), .ZN(n8380) );
  XNOR2_X1 U9514 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_116), .ZN(n8379) );
  OAI21_X1 U9515 ( .B1(n8381), .B2(n8380), .A(n8379), .ZN(n8385) );
  XNOR2_X1 U9516 ( .A(n8382), .B(keyinput_118), .ZN(n8384) );
  XNOR2_X1 U9517 ( .A(n8599), .B(keyinput_117), .ZN(n8383) );
  NAND3_X1 U9518 ( .A1(n8385), .A2(n8384), .A3(n8383), .ZN(n8388) );
  XNOR2_X1 U9519 ( .A(n6643), .B(keyinput_119), .ZN(n8387) );
  XNOR2_X1 U9520 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_120), .ZN(n8386) );
  NAND3_X1 U9521 ( .A1(n8388), .A2(n8387), .A3(n8386), .ZN(n8394) );
  XNOR2_X1 U9522 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_121), .ZN(n8393) );
  XOR2_X1 U9523 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_122), .Z(n8391) );
  XOR2_X1 U9524 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_124), .Z(n8390) );
  XNOR2_X1 U9525 ( .A(n8608), .B(keyinput_123), .ZN(n8389) );
  NAND3_X1 U9526 ( .A1(n8391), .A2(n8390), .A3(n8389), .ZN(n8392) );
  AOI21_X1 U9527 ( .B1(n8394), .B2(n8393), .A(n8392), .ZN(n8398) );
  INV_X1 U9528 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10552) );
  XNOR2_X1 U9529 ( .A(n10552), .B(keyinput_125), .ZN(n8397) );
  XOR2_X1 U9530 ( .A(P1_D_REG_3__SCAN_IN), .B(keyinput_126), .Z(n8396) );
  XOR2_X1 U9531 ( .A(P1_D_REG_4__SCAN_IN), .B(keyinput_127), .Z(n8395) );
  OAI211_X1 U9532 ( .C1(n8398), .C2(n8397), .A(n8396), .B(n8395), .ZN(n8618)
         );
  XOR2_X1 U9533 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_128), .Z(n8401) );
  XOR2_X1 U9534 ( .A(SI_31_), .B(keyinput_129), .Z(n8400) );
  XOR2_X1 U9535 ( .A(SI_30_), .B(keyinput_130), .Z(n8399) );
  AOI21_X1 U9536 ( .B1(n8401), .B2(n8400), .A(n8399), .ZN(n8404) );
  XNOR2_X1 U9537 ( .A(SI_29_), .B(keyinput_131), .ZN(n8403) );
  XNOR2_X1 U9538 ( .A(SI_28_), .B(keyinput_132), .ZN(n8402) );
  NOR3_X1 U9539 ( .A1(n8404), .A2(n8403), .A3(n8402), .ZN(n8408) );
  XOR2_X1 U9540 ( .A(SI_27_), .B(keyinput_133), .Z(n8407) );
  XNOR2_X1 U9541 ( .A(n8405), .B(keyinput_134), .ZN(n8406) );
  OAI21_X1 U9542 ( .B1(n8408), .B2(n8407), .A(n8406), .ZN(n8412) );
  XNOR2_X1 U9543 ( .A(n8409), .B(keyinput_135), .ZN(n8411) );
  XNOR2_X1 U9544 ( .A(SI_24_), .B(keyinput_136), .ZN(n8410) );
  NAND3_X1 U9545 ( .A1(n8412), .A2(n8411), .A3(n8410), .ZN(n8416) );
  XNOR2_X1 U9546 ( .A(SI_23_), .B(keyinput_137), .ZN(n8415) );
  XNOR2_X1 U9547 ( .A(n8413), .B(keyinput_138), .ZN(n8414) );
  AOI21_X1 U9548 ( .B1(n8416), .B2(n8415), .A(n8414), .ZN(n8419) );
  XNOR2_X1 U9549 ( .A(SI_21_), .B(keyinput_139), .ZN(n8418) );
  XNOR2_X1 U9550 ( .A(SI_20_), .B(keyinput_140), .ZN(n8417) );
  OAI21_X1 U9551 ( .B1(n8419), .B2(n8418), .A(n8417), .ZN(n8423) );
  XNOR2_X1 U9552 ( .A(SI_19_), .B(keyinput_141), .ZN(n8422) );
  XNOR2_X1 U9553 ( .A(n8420), .B(keyinput_142), .ZN(n8421) );
  AOI21_X1 U9554 ( .B1(n8423), .B2(n8422), .A(n8421), .ZN(n8427) );
  XOR2_X1 U9555 ( .A(SI_16_), .B(keyinput_144), .Z(n8426) );
  XNOR2_X1 U9556 ( .A(SI_15_), .B(keyinput_145), .ZN(n8425) );
  XNOR2_X1 U9557 ( .A(SI_17_), .B(keyinput_143), .ZN(n8424) );
  NOR4_X1 U9558 ( .A1(n8427), .A2(n8426), .A3(n8425), .A4(n8424), .ZN(n8430)
         );
  XOR2_X1 U9559 ( .A(SI_14_), .B(keyinput_146), .Z(n8429) );
  XOR2_X1 U9560 ( .A(SI_13_), .B(keyinput_147), .Z(n8428) );
  OAI21_X1 U9561 ( .B1(n8430), .B2(n8429), .A(n8428), .ZN(n8442) );
  XNOR2_X1 U9562 ( .A(SI_12_), .B(keyinput_148), .ZN(n8441) );
  XNOR2_X1 U9563 ( .A(n8431), .B(keyinput_150), .ZN(n8435) );
  XNOR2_X1 U9564 ( .A(n8432), .B(keyinput_151), .ZN(n8434) );
  XNOR2_X1 U9565 ( .A(SI_7_), .B(keyinput_153), .ZN(n8433) );
  NOR3_X1 U9566 ( .A1(n8435), .A2(n8434), .A3(n8433), .ZN(n8439) );
  XNOR2_X1 U9567 ( .A(n8436), .B(keyinput_152), .ZN(n8438) );
  XNOR2_X1 U9568 ( .A(SI_11_), .B(keyinput_149), .ZN(n8437) );
  NAND3_X1 U9569 ( .A1(n8439), .A2(n8438), .A3(n8437), .ZN(n8440) );
  AOI21_X1 U9570 ( .B1(n8442), .B2(n8441), .A(n8440), .ZN(n8452) );
  XNOR2_X1 U9571 ( .A(n8443), .B(keyinput_154), .ZN(n8449) );
  XNOR2_X1 U9572 ( .A(n8444), .B(keyinput_157), .ZN(n8448) );
  XNOR2_X1 U9573 ( .A(n8445), .B(keyinput_156), .ZN(n8447) );
  XNOR2_X1 U9574 ( .A(SI_5_), .B(keyinput_155), .ZN(n8446) );
  NAND4_X1 U9575 ( .A1(n8449), .A2(n8448), .A3(n8447), .A4(n8446), .ZN(n8451)
         );
  XOR2_X1 U9576 ( .A(SI_2_), .B(keyinput_158), .Z(n8450) );
  OAI21_X1 U9577 ( .B1(n8452), .B2(n8451), .A(n8450), .ZN(n8462) );
  XNOR2_X1 U9578 ( .A(n5306), .B(keyinput_161), .ZN(n8458) );
  XNOR2_X1 U9579 ( .A(P2_U3152), .B(keyinput_162), .ZN(n8457) );
  XNOR2_X1 U9580 ( .A(n8454), .B(keyinput_159), .ZN(n8456) );
  XNOR2_X1 U9581 ( .A(SI_0_), .B(keyinput_160), .ZN(n8455) );
  NOR4_X1 U9582 ( .A1(n8458), .A2(n8457), .A3(n8456), .A4(n8455), .ZN(n8461)
         );
  XNOR2_X1 U9583 ( .A(n8459), .B(keyinput_163), .ZN(n8460) );
  AOI21_X1 U9584 ( .B1(n8462), .B2(n8461), .A(n8460), .ZN(n8469) );
  XNOR2_X1 U9585 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_164), .ZN(n8468)
         );
  XNOR2_X1 U9586 ( .A(n8463), .B(keyinput_167), .ZN(n8466) );
  XNOR2_X1 U9587 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_165), .ZN(n8465)
         );
  XNOR2_X1 U9588 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_166), .ZN(n8464)
         );
  NOR3_X1 U9589 ( .A1(n8466), .A2(n8465), .A3(n8464), .ZN(n8467) );
  OAI21_X1 U9590 ( .B1(n8469), .B2(n8468), .A(n8467), .ZN(n8472) );
  XNOR2_X1 U9591 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_168), .ZN(n8471) );
  XNOR2_X1 U9592 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput_169), .ZN(n8470)
         );
  AOI21_X1 U9593 ( .B1(n8472), .B2(n8471), .A(n8470), .ZN(n8477) );
  XNOR2_X1 U9594 ( .A(n8473), .B(keyinput_170), .ZN(n8476) );
  XNOR2_X1 U9595 ( .A(n8474), .B(keyinput_171), .ZN(n8475) );
  NOR3_X1 U9596 ( .A1(n8477), .A2(n8476), .A3(n8475), .ZN(n8480) );
  XOR2_X1 U9597 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_172), .Z(n8479) );
  XNOR2_X1 U9598 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_173), .ZN(n8478)
         );
  NOR3_X1 U9599 ( .A1(n8480), .A2(n8479), .A3(n8478), .ZN(n8487) );
  XNOR2_X1 U9600 ( .A(n8481), .B(keyinput_174), .ZN(n8486) );
  XNOR2_X1 U9601 ( .A(n8482), .B(keyinput_176), .ZN(n8485) );
  XNOR2_X1 U9602 ( .A(n8483), .B(keyinput_175), .ZN(n8484) );
  OAI211_X1 U9603 ( .C1(n8487), .C2(n8486), .A(n8485), .B(n8484), .ZN(n8496)
         );
  XNOR2_X1 U9604 ( .A(n8488), .B(keyinput_177), .ZN(n8492) );
  XNOR2_X1 U9605 ( .A(P2_REG3_REG_24__SCAN_IN), .B(keyinput_179), .ZN(n8491)
         );
  XNOR2_X1 U9606 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_180), .ZN(n8490) );
  XNOR2_X1 U9607 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_178), .ZN(n8489)
         );
  NOR4_X1 U9608 ( .A1(n8492), .A2(n8491), .A3(n8490), .A4(n8489), .ZN(n8495)
         );
  XNOR2_X1 U9609 ( .A(n8493), .B(keyinput_181), .ZN(n8494) );
  AOI21_X1 U9610 ( .B1(n8496), .B2(n8495), .A(n8494), .ZN(n8502) );
  XNOR2_X1 U9611 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_182), .ZN(n8501) );
  OAI22_X1 U9612 ( .A1(n9363), .A2(keyinput_185), .B1(P2_REG3_REG_13__SCAN_IN), 
        .B2(keyinput_184), .ZN(n8498) );
  AND2_X1 U9613 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput_184), .ZN(n8497)
         );
  AOI211_X1 U9614 ( .C1(keyinput_185), .C2(n9363), .A(n8498), .B(n8497), .ZN(
        n8500) );
  XNOR2_X1 U9615 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_183), .ZN(n8499)
         );
  OAI211_X1 U9616 ( .C1(n8502), .C2(n8501), .A(n8500), .B(n8499), .ZN(n8505)
         );
  XNOR2_X1 U9617 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_186), .ZN(n8504)
         );
  XNOR2_X1 U9618 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_187), .ZN(n8503) );
  NAND3_X1 U9619 ( .A1(n8505), .A2(n8504), .A3(n8503), .ZN(n8509) );
  XNOR2_X1 U9620 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_188), .ZN(n8508)
         );
  XNOR2_X1 U9621 ( .A(n8506), .B(keyinput_189), .ZN(n8507) );
  AOI21_X1 U9622 ( .B1(n8509), .B2(n8508), .A(n8507), .ZN(n8517) );
  XOR2_X1 U9623 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_193), .Z(n8514) );
  XNOR2_X1 U9624 ( .A(n8510), .B(keyinput_190), .ZN(n8513) );
  XNOR2_X1 U9625 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_192), .ZN(n8512) );
  XNOR2_X1 U9626 ( .A(P2_REG3_REG_15__SCAN_IN), .B(keyinput_191), .ZN(n8511)
         );
  NAND4_X1 U9627 ( .A1(n8514), .A2(n8513), .A3(n8512), .A4(n8511), .ZN(n8516)
         );
  XNOR2_X1 U9628 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(keyinput_194), .ZN(n8515)
         );
  OAI21_X1 U9629 ( .B1(n8517), .B2(n8516), .A(n8515), .ZN(n8520) );
  XNOR2_X1 U9630 ( .A(n10541), .B(keyinput_195), .ZN(n8519) );
  XNOR2_X1 U9631 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_196), .ZN(n8518)
         );
  NAND3_X1 U9632 ( .A1(n8520), .A2(n8519), .A3(n8518), .ZN(n8523) );
  XOR2_X1 U9633 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput_197), .Z(n8522) );
  XOR2_X1 U9634 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(keyinput_198), .Z(n8521) );
  AOI21_X1 U9635 ( .B1(n8523), .B2(n8522), .A(n8521), .ZN(n8529) );
  XNOR2_X1 U9636 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_199), .ZN(n8528)
         );
  XOR2_X1 U9637 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_200), .Z(n8526) );
  XOR2_X1 U9638 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput_201), .Z(n8525) );
  XNOR2_X1 U9639 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_202), .ZN(n8524)
         );
  NOR3_X1 U9640 ( .A1(n8526), .A2(n8525), .A3(n8524), .ZN(n8527) );
  OAI21_X1 U9641 ( .B1(n8529), .B2(n8528), .A(n8527), .ZN(n8532) );
  XNOR2_X1 U9642 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_203), .ZN(n8531)
         );
  XNOR2_X1 U9643 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput_204), .ZN(n8530)
         );
  AOI21_X1 U9644 ( .B1(n8532), .B2(n8531), .A(n8530), .ZN(n8535) );
  XNOR2_X1 U9645 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_205), .ZN(n8534)
         );
  XNOR2_X1 U9646 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_206), .ZN(n8533)
         );
  OAI21_X1 U9647 ( .B1(n8535), .B2(n8534), .A(n8533), .ZN(n8538) );
  XOR2_X1 U9648 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_207), .Z(n8537) );
  XNOR2_X1 U9649 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(keyinput_208), .ZN(n8536)
         );
  NAND3_X1 U9650 ( .A1(n8538), .A2(n8537), .A3(n8536), .ZN(n8544) );
  XNOR2_X1 U9651 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_209), .ZN(n8543)
         );
  XOR2_X1 U9652 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput_210), .Z(n8541) );
  XNOR2_X1 U9653 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_212), .ZN(n8540)
         );
  XNOR2_X1 U9654 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_211), .ZN(n8539)
         );
  NAND3_X1 U9655 ( .A1(n8541), .A2(n8540), .A3(n8539), .ZN(n8542) );
  AOI21_X1 U9656 ( .B1(n8544), .B2(n8543), .A(n8542), .ZN(n8547) );
  XOR2_X1 U9657 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_213), .Z(n8546) );
  XNOR2_X1 U9658 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_214), .ZN(n8545)
         );
  OAI21_X1 U9659 ( .B1(n8547), .B2(n8546), .A(n8545), .ZN(n8554) );
  XNOR2_X1 U9660 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput_215), .ZN(n8553)
         );
  XOR2_X1 U9661 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_217), .Z(n8551) );
  XNOR2_X1 U9662 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput_218), .ZN(n8550)
         );
  XNOR2_X1 U9663 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_216), .ZN(n8549)
         );
  XNOR2_X1 U9664 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_219), .ZN(n8548) );
  NAND4_X1 U9665 ( .A1(n8551), .A2(n8550), .A3(n8549), .A4(n8548), .ZN(n8552)
         );
  AOI21_X1 U9666 ( .B1(n8554), .B2(n8553), .A(n8552), .ZN(n8562) );
  XNOR2_X1 U9667 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_220), .ZN(n8561) );
  XOR2_X1 U9668 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_222), .Z(n8559) );
  XNOR2_X1 U9669 ( .A(n8555), .B(keyinput_223), .ZN(n8558) );
  XNOR2_X1 U9670 ( .A(n8556), .B(keyinput_221), .ZN(n8557) );
  NOR3_X1 U9671 ( .A1(n8559), .A2(n8558), .A3(n8557), .ZN(n8560) );
  OAI21_X1 U9672 ( .B1(n8562), .B2(n8561), .A(n8560), .ZN(n8566) );
  XNOR2_X1 U9673 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_226), .ZN(n8565) );
  XNOR2_X1 U9674 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_225), .ZN(n8564) );
  XNOR2_X1 U9675 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_224), .ZN(n8563) );
  NAND4_X1 U9676 ( .A1(n8566), .A2(n8565), .A3(n8564), .A4(n8563), .ZN(n8570)
         );
  XNOR2_X1 U9677 ( .A(n8567), .B(keyinput_227), .ZN(n8569) );
  XNOR2_X1 U9678 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_228), .ZN(n8568) );
  AOI21_X1 U9679 ( .B1(n8570), .B2(n8569), .A(n8568), .ZN(n8575) );
  XNOR2_X1 U9680 ( .A(n8571), .B(keyinput_231), .ZN(n8574) );
  XOR2_X1 U9681 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_229), .Z(n8573) );
  XNOR2_X1 U9682 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_230), .ZN(n8572) );
  NOR4_X1 U9683 ( .A1(n8575), .A2(n8574), .A3(n8573), .A4(n8572), .ZN(n8578)
         );
  XNOR2_X1 U9684 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_232), .ZN(n8577) );
  XNOR2_X1 U9685 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_233), .ZN(n8576) );
  OAI21_X1 U9686 ( .B1(n8578), .B2(n8577), .A(n8576), .ZN(n8582) );
  XNOR2_X1 U9687 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_235), .ZN(n8581) );
  XNOR2_X1 U9688 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_236), .ZN(n8580) );
  XNOR2_X1 U9689 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_234), .ZN(n8579) );
  NAND4_X1 U9690 ( .A1(n8582), .A2(n8581), .A3(n8580), .A4(n8579), .ZN(n8589)
         );
  XNOR2_X1 U9691 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_237), .ZN(n8588) );
  XOR2_X1 U9692 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_238), .Z(n8586) );
  XNOR2_X1 U9693 ( .A(n8583), .B(keyinput_239), .ZN(n8585) );
  XNOR2_X1 U9694 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_240), .ZN(n8584) );
  NAND3_X1 U9695 ( .A1(n8586), .A2(n8585), .A3(n8584), .ZN(n8587) );
  AOI21_X1 U9696 ( .B1(n8589), .B2(n8588), .A(n8587), .ZN(n8594) );
  XNOR2_X1 U9697 ( .A(n8590), .B(keyinput_241), .ZN(n8593) );
  XNOR2_X1 U9698 ( .A(n8591), .B(keyinput_242), .ZN(n8592) );
  OAI21_X1 U9699 ( .B1(n8594), .B2(n8593), .A(n8592), .ZN(n8598) );
  XNOR2_X1 U9700 ( .A(n8595), .B(keyinput_243), .ZN(n8597) );
  XNOR2_X1 U9701 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_244), .ZN(n8596) );
  AOI21_X1 U9702 ( .B1(n8598), .B2(n8597), .A(n8596), .ZN(n8602) );
  XNOR2_X1 U9703 ( .A(n8599), .B(keyinput_245), .ZN(n8601) );
  XNOR2_X1 U9704 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_246), .ZN(n8600) );
  NOR3_X1 U9705 ( .A1(n8602), .A2(n8601), .A3(n8600), .ZN(n8605) );
  XNOR2_X1 U9706 ( .A(n6643), .B(keyinput_247), .ZN(n8604) );
  XOR2_X1 U9707 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_248), .Z(n8603) );
  NOR3_X1 U9708 ( .A1(n8605), .A2(n8604), .A3(n8603), .ZN(n8612) );
  XNOR2_X1 U9709 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_249), .ZN(n8611) );
  XOR2_X1 U9710 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_252), .Z(n8610) );
  OAI22_X1 U9711 ( .A1(n8608), .A2(keyinput_251), .B1(keyinput_250), .B2(
        P1_IR_REG_31__SCAN_IN), .ZN(n8607) );
  AND2_X1 U9712 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(keyinput_250), .ZN(n8606) );
  AOI211_X1 U9713 ( .C1(keyinput_251), .C2(n8608), .A(n8607), .B(n8606), .ZN(
        n8609) );
  OAI211_X1 U9714 ( .C1(n8612), .C2(n8611), .A(n8610), .B(n8609), .ZN(n8616)
         );
  XNOR2_X1 U9715 ( .A(P1_D_REG_2__SCAN_IN), .B(keyinput_253), .ZN(n8615) );
  XNOR2_X1 U9716 ( .A(keyinput_254), .B(P1_D_REG_3__SCAN_IN), .ZN(n8614) );
  XNOR2_X1 U9717 ( .A(keyinput_255), .B(P1_D_REG_4__SCAN_IN), .ZN(n8613) );
  AOI211_X1 U9718 ( .C1(n8616), .C2(n8615), .A(n8614), .B(n8613), .ZN(n8617)
         );
  NOR2_X1 U9719 ( .A1(n8618), .A2(n8617), .ZN(n8627) );
  OAI21_X1 U9720 ( .B1(n8620), .B2(P1_REG1_REG_0__SCAN_IN), .A(n8619), .ZN(
        n8621) );
  XOR2_X1 U9721 ( .A(P1_IR_REG_0__SCAN_IN), .B(n8621), .Z(n8624) );
  OAI22_X1 U9722 ( .A1(n8624), .A2(n8623), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8622), .ZN(n8625) );
  AOI21_X1 U9723 ( .B1(n10670), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n8625), .ZN(
        n8626) );
  XNOR2_X1 U9724 ( .A(n8627), .B(n8626), .ZN(P1_U3241) );
  INV_X1 U9725 ( .A(n8628), .ZN(n8632) );
  OAI222_X1 U9726 ( .A1(n8630), .A2(P1_U3084), .B1(n8088), .B2(n8632), .C1(
        n8629), .C2(n10546), .ZN(P1_U3331) );
  OAI222_X1 U9727 ( .A1(n9923), .A2(n8633), .B1(n5076), .B2(n8632), .C1(
        P2_U3152), .C2(n8631), .ZN(P2_U3336) );
  AND2_X1 U9728 ( .A1(n8969), .A2(n8971), .ZN(n9076) );
  NAND2_X1 U9729 ( .A1(n9151), .A2(n9076), .ZN(n8634) );
  INV_X1 U9730 ( .A(n10097), .ZN(n8765) );
  NOR2_X1 U9731 ( .A1(n8790), .A2(n8765), .ZN(n9051) );
  NAND2_X1 U9732 ( .A1(n8790), .A2(n8765), .ZN(n9044) );
  INV_X1 U9733 ( .A(n9044), .ZN(n8973) );
  XNOR2_X1 U9734 ( .A(n8784), .B(n5113), .ZN(n8635) );
  OAI222_X1 U9735 ( .A1(n10887), .A2(n10890), .B1(n10889), .B2(n8636), .C1(
        n10784), .C2(n8635), .ZN(n10860) );
  INV_X1 U9736 ( .A(n10860), .ZN(n8647) );
  NAND2_X1 U9737 ( .A1(n8637), .A2(n10098), .ZN(n8638) );
  NAND2_X1 U9738 ( .A1(n8639), .A2(n8638), .ZN(n8789) );
  XNOR2_X1 U9739 ( .A(n8789), .B(n5113), .ZN(n10862) );
  INV_X1 U9740 ( .A(n8640), .ZN(n8641) );
  OAI21_X1 U9741 ( .B1(n5390), .B2(n8641), .A(n5183), .ZN(n10859) );
  OAI22_X1 U9742 ( .A1(n5074), .A2(n8642), .B1(n10008), .B2(n10907), .ZN(n8643) );
  AOI21_X1 U9743 ( .B1(n10432), .B2(n8790), .A(n8643), .ZN(n8644) );
  OAI21_X1 U9744 ( .B1(n10859), .B2(n10435), .A(n8644), .ZN(n8645) );
  AOI21_X1 U9745 ( .B1(n10862), .B2(n10437), .A(n8645), .ZN(n8646) );
  OAI21_X1 U9746 ( .B1(n8647), .B2(n10439), .A(n8646), .ZN(P1_U3282) );
  INV_X1 U9747 ( .A(n8648), .ZN(n9401) );
  NAND2_X1 U9748 ( .A1(n10852), .A2(n9401), .ZN(n8649) );
  OAI21_X1 U9749 ( .B1(n5180), .B2(n8650), .A(n8670), .ZN(n10870) );
  INV_X1 U9750 ( .A(n10870), .ZN(n8660) );
  INV_X1 U9751 ( .A(n9728), .ZN(n8744) );
  INV_X1 U9752 ( .A(n8664), .ZN(n10925) );
  AOI22_X1 U9753 ( .A1(n10924), .A2(n9401), .B1(n10925), .B2(n10926), .ZN(
        n8653) );
  OAI211_X1 U9754 ( .C1(n5708), .C2(n5899), .A(n10929), .B(n8651), .ZN(n8652)
         );
  OAI211_X1 U9755 ( .C1(n8660), .C2(n9813), .A(n8653), .B(n8652), .ZN(n10868)
         );
  NAND2_X1 U9756 ( .A1(n10868), .A2(n10947), .ZN(n8659) );
  OAI22_X1 U9757 ( .A1(n10947), .A2(n8655), .B1(n8654), .B2(n10700), .ZN(n8657) );
  XNOR2_X1 U9758 ( .A(n8683), .B(n10865), .ZN(n10867) );
  NOR2_X1 U9759 ( .A1(n10867), .A2(n10702), .ZN(n8656) );
  AOI211_X1 U9760 ( .C1(n9797), .C2(n10865), .A(n8657), .B(n8656), .ZN(n8658)
         );
  OAI211_X1 U9761 ( .C1(n8660), .C2(n8744), .A(n8659), .B(n8658), .ZN(P2_U3287) );
  XNOR2_X1 U9762 ( .A(n8662), .B(n8661), .ZN(n8668) );
  OAI22_X1 U9763 ( .A1(n9386), .A2(n10936), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8663), .ZN(n8666) );
  OAI22_X1 U9764 ( .A1(n9398), .A2(n9372), .B1(n9371), .B2(n8664), .ZN(n8665)
         );
  AOI211_X1 U9765 ( .C1(n10939), .C2(n9389), .A(n8666), .B(n8665), .ZN(n8667)
         );
  OAI21_X1 U9766 ( .B1(n8668), .B2(n9391), .A(n8667), .ZN(P2_U3238) );
  INV_X1 U9767 ( .A(n8673), .ZN(n8672) );
  INV_X1 U9768 ( .A(n8675), .ZN(n8671) );
  NAND2_X1 U9769 ( .A1(n8673), .A2(n8675), .ZN(n8674) );
  AND2_X1 U9770 ( .A1(n8813), .A2(n8674), .ZN(n10877) );
  XNOR2_X1 U9771 ( .A(n8676), .B(n8675), .ZN(n8680) );
  OAI22_X1 U9772 ( .A1(n9399), .A2(n9720), .B1(n8677), .B2(n9774), .ZN(n8678)
         );
  INV_X1 U9773 ( .A(n8678), .ZN(n8679) );
  OAI21_X1 U9774 ( .B1(n8680), .B2(n9717), .A(n8679), .ZN(n8681) );
  AOI21_X1 U9775 ( .B1(n10877), .B2(n8682), .A(n8681), .ZN(n10879) );
  INV_X1 U9776 ( .A(n8811), .ZN(n10873) );
  NOR2_X1 U9777 ( .A1(n8684), .A2(n10873), .ZN(n8685) );
  OR2_X1 U9778 ( .A1(n10931), .A2(n8685), .ZN(n10874) );
  OAI22_X1 U9779 ( .A1(n10947), .A2(n8687), .B1(n8686), .B2(n10700), .ZN(n8688) );
  AOI21_X1 U9780 ( .B1(n9797), .B2(n8811), .A(n8688), .ZN(n8689) );
  OAI21_X1 U9781 ( .B1(n10874), .B2(n10702), .A(n8689), .ZN(n8690) );
  AOI21_X1 U9782 ( .B1(n10877), .B2(n9728), .A(n8690), .ZN(n8691) );
  OAI21_X1 U9783 ( .B1(n10879), .B2(n10949), .A(n8691), .ZN(P2_U3286) );
  AOI21_X1 U9784 ( .B1(n8693), .B2(n8692), .A(n6851), .ZN(n8700) );
  AOI22_X1 U9785 ( .A1(n10086), .A2(n10098), .B1(n10081), .B2(n10100), .ZN(
        n8699) );
  NOR2_X1 U9786 ( .A1(n10083), .A2(n8694), .ZN(n8695) );
  AOI211_X1 U9787 ( .C1(n8697), .C2(n10069), .A(n8696), .B(n8695), .ZN(n8698)
         );
  OAI211_X1 U9788 ( .C1(n8700), .C2(n10071), .A(n8699), .B(n8698), .ZN(
        P1_U3211) );
  NOR2_X1 U9789 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n8736) );
  NOR2_X1 U9790 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n8734) );
  NOR2_X1 U9791 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n8732) );
  NOR2_X1 U9792 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n8730) );
  NOR2_X1 U9793 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n8728) );
  NOR2_X1 U9794 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n8726) );
  NAND2_X1 U9795 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n8724) );
  XOR2_X1 U9796 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n10605) );
  NAND2_X1 U9797 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n8722) );
  XOR2_X1 U9798 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n10603) );
  NOR2_X1 U9799 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n8706) );
  XNOR2_X1 U9800 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10594) );
  NAND2_X1 U9801 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n8704) );
  XOR2_X1 U9802 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(P1_ADDR_REG_3__SCAN_IN), .Z(
        n10592) );
  NAND2_X1 U9803 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n8702) );
  XOR2_X1 U9804 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10590) );
  AOI21_X1 U9805 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10585) );
  INV_X1 U9806 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10640) );
  NAND3_X1 U9807 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_1__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10587) );
  OAI21_X1 U9808 ( .B1(n10585), .B2(n10640), .A(n10587), .ZN(n10589) );
  NAND2_X1 U9809 ( .A1(n10590), .A2(n10589), .ZN(n8701) );
  NAND2_X1 U9810 ( .A1(n8702), .A2(n8701), .ZN(n10591) );
  NAND2_X1 U9811 ( .A1(n10592), .A2(n10591), .ZN(n8703) );
  NAND2_X1 U9812 ( .A1(n8704), .A2(n8703), .ZN(n10593) );
  NOR2_X1 U9813 ( .A1(n10594), .A2(n10593), .ZN(n8705) );
  NOR2_X1 U9814 ( .A1(n8706), .A2(n8705), .ZN(n8707) );
  NOR2_X1 U9815 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n8707), .ZN(n10596) );
  AND2_X1 U9816 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n8707), .ZN(n10595) );
  NOR2_X1 U9817 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10595), .ZN(n8708) );
  NOR2_X1 U9818 ( .A1(n10596), .A2(n8708), .ZN(n8709) );
  NAND2_X1 U9819 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n8709), .ZN(n8711) );
  XOR2_X1 U9820 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n8709), .Z(n10598) );
  NAND2_X1 U9821 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10598), .ZN(n8710) );
  NAND2_X1 U9822 ( .A1(n8711), .A2(n8710), .ZN(n8712) );
  NAND2_X1 U9823 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n8712), .ZN(n8714) );
  XOR2_X1 U9824 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n8712), .Z(n10599) );
  NAND2_X1 U9825 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10599), .ZN(n8713) );
  NAND2_X1 U9826 ( .A1(n8714), .A2(n8713), .ZN(n8715) );
  NAND2_X1 U9827 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n8715), .ZN(n8717) );
  XOR2_X1 U9828 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n8715), .Z(n10600) );
  NAND2_X1 U9829 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10600), .ZN(n8716) );
  NAND2_X1 U9830 ( .A1(n8717), .A2(n8716), .ZN(n8718) );
  NAND2_X1 U9831 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n8718), .ZN(n8720) );
  XOR2_X1 U9832 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n8718), .Z(n10601) );
  NAND2_X1 U9833 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10601), .ZN(n8719) );
  NAND2_X1 U9834 ( .A1(n8720), .A2(n8719), .ZN(n10602) );
  NAND2_X1 U9835 ( .A1(n10603), .A2(n10602), .ZN(n8721) );
  NAND2_X1 U9836 ( .A1(n8722), .A2(n8721), .ZN(n10604) );
  NAND2_X1 U9837 ( .A1(n10605), .A2(n10604), .ZN(n8723) );
  NAND2_X1 U9838 ( .A1(n8724), .A2(n8723), .ZN(n10607) );
  XNOR2_X1 U9839 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10606) );
  NOR2_X1 U9840 ( .A1(n10607), .A2(n10606), .ZN(n8725) );
  NOR2_X1 U9841 ( .A1(n8726), .A2(n8725), .ZN(n10609) );
  XNOR2_X1 U9842 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10608) );
  NOR2_X1 U9843 ( .A1(n10609), .A2(n10608), .ZN(n8727) );
  NOR2_X1 U9844 ( .A1(n8728), .A2(n8727), .ZN(n10611) );
  XNOR2_X1 U9845 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10610) );
  NOR2_X1 U9846 ( .A1(n10611), .A2(n10610), .ZN(n8729) );
  NOR2_X1 U9847 ( .A1(n8730), .A2(n8729), .ZN(n10613) );
  XNOR2_X1 U9848 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10612) );
  NOR2_X1 U9849 ( .A1(n10613), .A2(n10612), .ZN(n8731) );
  NOR2_X1 U9850 ( .A1(n8732), .A2(n8731), .ZN(n10615) );
  XNOR2_X1 U9851 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10614) );
  NOR2_X1 U9852 ( .A1(n10615), .A2(n10614), .ZN(n8733) );
  NOR2_X1 U9853 ( .A1(n8734), .A2(n8733), .ZN(n10617) );
  XNOR2_X1 U9854 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10616) );
  NOR2_X1 U9855 ( .A1(n10617), .A2(n10616), .ZN(n8735) );
  NOR2_X1 U9856 ( .A1(n8736), .A2(n8735), .ZN(n8737) );
  AND2_X1 U9857 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n8737), .ZN(n10618) );
  NOR2_X1 U9858 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10618), .ZN(n8738) );
  NOR2_X1 U9859 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n8737), .ZN(n10619) );
  NOR2_X1 U9860 ( .A1(n8738), .A2(n10619), .ZN(n8740) );
  XNOR2_X1 U9861 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n8739) );
  XNOR2_X1 U9862 ( .A(n8740), .B(n8739), .ZN(ADD_1071_U4) );
  INV_X1 U9863 ( .A(n8741), .ZN(n8742) );
  OAI22_X1 U9864 ( .A1(n8742), .A2(n10702), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n10700), .ZN(n8747) );
  OAI22_X1 U9865 ( .A1(n8745), .A2(n8744), .B1(n8743), .B2(n10705), .ZN(n8746)
         );
  AOI211_X1 U9866 ( .C1(P2_REG2_REG_3__SCAN_IN), .C2(n10949), .A(n8747), .B(
        n8746), .ZN(n8748) );
  OAI21_X1 U9867 ( .B1(n8749), .B2(n10949), .A(n8748), .ZN(P2_U3293) );
  NAND2_X1 U9868 ( .A1(n8753), .A2(n10538), .ZN(n8751) );
  OR2_X1 U9869 ( .A1(n8750), .A2(P1_U3084), .ZN(n9190) );
  OAI211_X1 U9870 ( .C1(n8752), .C2(n8845), .A(n8751), .B(n9190), .ZN(P1_U3330) );
  NAND2_X1 U9871 ( .A1(n8753), .A2(n9910), .ZN(n8755) );
  OAI211_X1 U9872 ( .C1(n7477), .C2(n9923), .A(n8755), .B(n8754), .ZN(P2_U3335) );
  NAND2_X1 U9873 ( .A1(n8757), .A2(n8756), .ZN(n8759) );
  NAND2_X1 U9874 ( .A1(n8759), .A2(n8758), .ZN(n8760) );
  NAND2_X1 U9875 ( .A1(n10003), .A2(n8760), .ZN(n8762) );
  XNOR2_X1 U9876 ( .A(n8762), .B(n8761), .ZN(n8763) );
  NAND2_X1 U9877 ( .A1(n8763), .A2(n10078), .ZN(n8769) );
  OAI22_X1 U9878 ( .A1(n10065), .A2(n8765), .B1(n10083), .B2(n8764), .ZN(n8766) );
  AOI211_X1 U9879 ( .C1(n10081), .C2(n10099), .A(n8767), .B(n8766), .ZN(n8768)
         );
  OAI211_X1 U9880 ( .C1(n10843), .C2(n10089), .A(n8769), .B(n8768), .ZN(
        P1_U3219) );
  OAI222_X1 U9881 ( .A1(n5076), .A2(n8773), .B1(P2_U3152), .B2(n8771), .C1(
        n8770), .C2(n9923), .ZN(P2_U3334) );
  OAI222_X1 U9882 ( .A1(n8774), .A2(P1_U3084), .B1(n8088), .B2(n8773), .C1(
        n8772), .C2(n10546), .ZN(P1_U3329) );
  INV_X1 U9883 ( .A(n8775), .ZN(n8776) );
  AOI21_X1 U9884 ( .B1(n8778), .B2(n8777), .A(n8776), .ZN(n8783) );
  OAI21_X1 U9885 ( .B1(n9386), .B2(n8820), .A(n8779), .ZN(n8781) );
  OAI22_X1 U9886 ( .A1(n9775), .A2(n9372), .B1(n9371), .B2(n9399), .ZN(n8780)
         );
  AOI211_X1 U9887 ( .C1(n8858), .C2(n9389), .A(n8781), .B(n8780), .ZN(n8782)
         );
  OAI21_X1 U9888 ( .B1(n8783), .B2(n9391), .A(n8782), .ZN(P2_U3226) );
  NAND2_X1 U9889 ( .A1(n8868), .A2(n10890), .ZN(n9045) );
  XNOR2_X1 U9890 ( .A(n8830), .B(n9134), .ZN(n8785) );
  AOI222_X1 U9891 ( .A1(n10097), .A2(n10405), .B1(n10095), .B2(n10398), .C1(
        n10892), .C2(n8785), .ZN(n8870) );
  INV_X1 U9892 ( .A(n8868), .ZN(n8885) );
  AOI211_X1 U9893 ( .C1(n8868), .C2(n5183), .A(n11005), .B(n10884), .ZN(n8867)
         );
  INV_X1 U9894 ( .A(n8880), .ZN(n8786) );
  INV_X1 U9895 ( .A(n10907), .ZN(n10790) );
  AOI22_X1 U9896 ( .A1(n10439), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n8786), .B2(
        n10790), .ZN(n8787) );
  OAI21_X1 U9897 ( .B1(n8885), .B2(n10905), .A(n8787), .ZN(n8796) );
  OR2_X1 U9898 ( .A1(n8790), .A2(n10097), .ZN(n8788) );
  NAND2_X1 U9899 ( .A1(n8789), .A2(n8788), .ZN(n8792) );
  NAND2_X1 U9900 ( .A1(n8790), .A2(n10097), .ZN(n8791) );
  INV_X1 U9901 ( .A(n8828), .ZN(n8793) );
  AOI21_X1 U9902 ( .B1(n9134), .B2(n8794), .A(n8793), .ZN(n8871) );
  NOR2_X1 U9903 ( .A1(n8871), .A2(n10381), .ZN(n8795) );
  AOI211_X1 U9904 ( .C1(n8867), .C2(n10373), .A(n8796), .B(n8795), .ZN(n8797)
         );
  OAI21_X1 U9905 ( .B1(n10439), .B2(n8870), .A(n8797), .ZN(P1_U3281) );
  OAI21_X1 U9906 ( .B1(n8800), .B2(n8799), .A(n8798), .ZN(n8801) );
  NAND2_X1 U9907 ( .A1(n8801), .A2(n9341), .ZN(n8806) );
  INV_X1 U9908 ( .A(n8851), .ZN(n8804) );
  OAI22_X1 U9909 ( .A1(n9508), .A2(n9372), .B1(n9371), .B2(n9398), .ZN(n8802)
         );
  AOI211_X1 U9910 ( .C1(n8903), .C2(n8804), .A(n8803), .B(n8802), .ZN(n8805)
         );
  OAI211_X1 U9911 ( .C1(n10974), .C2(n9335), .A(n8806), .B(n8805), .ZN(
        P2_U3236) );
  INV_X1 U9912 ( .A(n8807), .ZN(n8808) );
  NOR2_X1 U9913 ( .A1(n10918), .A2(n8808), .ZN(n8809) );
  XNOR2_X1 U9914 ( .A(n8809), .B(n8817), .ZN(n8810) );
  OAI222_X1 U9915 ( .A1(n9720), .A2(n9775), .B1(n8810), .B2(n9717), .C1(n9774), 
        .C2(n9399), .ZN(n10960) );
  INV_X1 U9916 ( .A(n10960), .ZN(n8826) );
  NAND2_X1 U9917 ( .A1(n8811), .A2(n10925), .ZN(n8812) );
  NAND2_X1 U9918 ( .A1(n8813), .A2(n8812), .ZN(n10916) );
  AOI21_X1 U9919 ( .B1(n8817), .B2(n8816), .A(n8815), .ZN(n8818) );
  INV_X1 U9920 ( .A(n8818), .ZN(n10962) );
  NAND2_X1 U9921 ( .A1(n5188), .A2(n8858), .ZN(n8819) );
  NAND2_X1 U9922 ( .A1(n8853), .A2(n8819), .ZN(n10959) );
  OAI22_X1 U9923 ( .A1(n10947), .A2(n8821), .B1(n8820), .B2(n10700), .ZN(n8822) );
  AOI21_X1 U9924 ( .B1(n8858), .B2(n9797), .A(n8822), .ZN(n8823) );
  OAI21_X1 U9925 ( .B1(n10959), .B2(n10702), .A(n8823), .ZN(n8824) );
  AOI21_X1 U9926 ( .B1(n10962), .B2(n9800), .A(n8824), .ZN(n8825) );
  OAI21_X1 U9927 ( .B1(n10949), .B2(n8826), .A(n8825), .ZN(P2_U3284) );
  OR2_X1 U9928 ( .A1(n8868), .A2(n10096), .ZN(n8827) );
  NOR2_X1 U9929 ( .A1(n8962), .A2(n10095), .ZN(n9120) );
  NAND2_X1 U9930 ( .A1(n8962), .A2(n10095), .ZN(n9118) );
  OR2_X1 U9931 ( .A1(n9210), .A2(n10888), .ZN(n9056) );
  INV_X1 U9932 ( .A(n10419), .ZN(n9057) );
  NAND2_X1 U9933 ( .A1(n9056), .A2(n9057), .ZN(n9137) );
  OAI21_X1 U9934 ( .B1(n8829), .B2(n9137), .A(n9212), .ZN(n10950) );
  INV_X1 U9935 ( .A(n10095), .ZN(n8911) );
  NAND2_X1 U9936 ( .A1(n8962), .A2(n8911), .ZN(n9048) );
  OR2_X1 U9937 ( .A1(n8962), .A2(n8911), .ZN(n9055) );
  INV_X1 U9938 ( .A(n9055), .ZN(n8831) );
  OR2_X1 U9939 ( .A1(n9236), .A2(n8831), .ZN(n8832) );
  XNOR2_X1 U9940 ( .A(n8832), .B(n9137), .ZN(n8833) );
  NAND2_X1 U9941 ( .A1(n8833), .A2(n10892), .ZN(n8835) );
  AOI22_X1 U9942 ( .A1(n10405), .A2(n10095), .B1(n10404), .B2(n10398), .ZN(
        n8834) );
  NAND2_X1 U9943 ( .A1(n8835), .A2(n8834), .ZN(n10953) );
  NAND2_X1 U9944 ( .A1(n10953), .A2(n5074), .ZN(n8840) );
  OAI22_X1 U9945 ( .A1(n5074), .A2(n8836), .B1(n8910), .B2(n10907), .ZN(n8838)
         );
  INV_X1 U9946 ( .A(n8962), .ZN(n10906) );
  NAND2_X1 U9947 ( .A1(n10884), .A2(n10906), .ZN(n10883) );
  INV_X1 U9948 ( .A(n9210), .ZN(n10952) );
  OAI211_X1 U9949 ( .C1(n5075), .C2(n10952), .A(n10778), .B(n5191), .ZN(n10951) );
  NOR2_X1 U9950 ( .A1(n10951), .A2(n10410), .ZN(n8837) );
  AOI211_X1 U9951 ( .C1(n10432), .C2(n9210), .A(n8838), .B(n8837), .ZN(n8839)
         );
  OAI211_X1 U9952 ( .C1(n10381), .C2(n10950), .A(n8840), .B(n8839), .ZN(
        P1_U3279) );
  INV_X1 U9953 ( .A(n8841), .ZN(n8847) );
  INV_X1 U9954 ( .A(n8842), .ZN(n8843) );
  OAI222_X1 U9955 ( .A1(n9923), .A2(n8844), .B1(n5076), .B2(n8847), .C1(n8843), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  OAI222_X1 U9956 ( .A1(P1_U3084), .A2(n8848), .B1(n8088), .B2(n8847), .C1(
        n8846), .C2(n8845), .ZN(P1_U3328) );
  AOI21_X1 U9957 ( .B1(n8849), .B2(n8861), .A(n5165), .ZN(n8850) );
  OAI222_X1 U9958 ( .A1(n9720), .A2(n9508), .B1(n9774), .B2(n9398), .C1(n9717), 
        .C2(n8850), .ZN(n10976) );
  INV_X1 U9959 ( .A(n10976), .ZN(n8866) );
  OAI22_X1 U9960 ( .A1(n10947), .A2(n8852), .B1(n8851), .B2(n10700), .ZN(n8856) );
  INV_X1 U9961 ( .A(n9778), .ZN(n8854) );
  OAI21_X1 U9962 ( .B1(n10974), .B2(n5340), .A(n8854), .ZN(n10975) );
  NOR2_X1 U9963 ( .A1(n10975), .A2(n10702), .ZN(n8855) );
  AOI211_X1 U9964 ( .C1(n9797), .C2(n8857), .A(n8856), .B(n8855), .ZN(n8865)
         );
  INV_X1 U9965 ( .A(n8858), .ZN(n10958) );
  NAND2_X1 U9966 ( .A1(n10958), .A2(n9398), .ZN(n8859) );
  NOR2_X1 U9967 ( .A1(n8862), .A2(n8861), .ZN(n10973) );
  INV_X1 U9968 ( .A(n10973), .ZN(n8863) );
  NAND3_X1 U9969 ( .A1(n8863), .A2(n9800), .A3(n9507), .ZN(n8864) );
  OAI211_X1 U9970 ( .C1(n8866), .C2(n10949), .A(n8865), .B(n8864), .ZN(
        P2_U3283) );
  AND2_X1 U9971 ( .A1(n10895), .A2(n10737), .ZN(n10516) );
  AOI21_X1 U9972 ( .B1(n10721), .B2(n8868), .A(n8867), .ZN(n8869) );
  OAI211_X1 U9973 ( .C1(n10516), .C2(n8871), .A(n8870), .B(n8869), .ZN(n8873)
         );
  NAND2_X1 U9974 ( .A1(n8873), .A2(n11020), .ZN(n8872) );
  OAI21_X1 U9975 ( .B1(n11020), .B2(n7254), .A(n8872), .ZN(P1_U3533) );
  NAND2_X1 U9976 ( .A1(n8873), .A2(n11024), .ZN(n8874) );
  OAI21_X1 U9977 ( .B1(n11024), .B2(n6901), .A(n8874), .ZN(P1_U3484) );
  NAND2_X1 U9978 ( .A1(n8876), .A2(n8875), .ZN(n8878) );
  XNOR2_X1 U9979 ( .A(n8878), .B(n8877), .ZN(n8879) );
  NAND2_X1 U9980 ( .A1(n8879), .A2(n10078), .ZN(n8884) );
  OAI22_X1 U9981 ( .A1(n10065), .A2(n8911), .B1(n10083), .B2(n8880), .ZN(n8881) );
  AOI211_X1 U9982 ( .C1(n10081), .C2(n10097), .A(n8882), .B(n8881), .ZN(n8883)
         );
  OAI211_X1 U9983 ( .C1(n8885), .C2(n10089), .A(n8884), .B(n8883), .ZN(
        P1_U3215) );
  NAND2_X1 U9984 ( .A1(n8887), .A2(n8886), .ZN(n8889) );
  XOR2_X1 U9985 ( .A(n8889), .B(n8888), .Z(n8895) );
  INV_X1 U9986 ( .A(n10908), .ZN(n8890) );
  AOI22_X1 U9987 ( .A1(n10086), .A2(n10094), .B1(n8890), .B2(n9930), .ZN(n8892) );
  OAI211_X1 U9988 ( .C1(n10890), .C2(n10066), .A(n8892), .B(n8891), .ZN(n8893)
         );
  AOI21_X1 U9989 ( .B1(n8962), .B2(n10069), .A(n8893), .ZN(n8894) );
  OAI21_X1 U9990 ( .B1(n8895), .B2(n10071), .A(n8894), .ZN(P1_U3234) );
  OAI21_X1 U9991 ( .B1(n8898), .B2(n8897), .A(n8896), .ZN(n8899) );
  NAND2_X1 U9992 ( .A1(n8899), .A2(n9341), .ZN(n8905) );
  INV_X1 U9993 ( .A(n9777), .ZN(n8902) );
  OAI22_X1 U9994 ( .A1(n9396), .A2(n9372), .B1(n9371), .B2(n9775), .ZN(n8900)
         );
  AOI211_X1 U9995 ( .C1(n8903), .C2(n8902), .A(n8901), .B(n8900), .ZN(n8904)
         );
  OAI211_X1 U9996 ( .C1(n10990), .C2(n9335), .A(n8905), .B(n8904), .ZN(
        P2_U3217) );
  XNOR2_X1 U9997 ( .A(n8908), .B(n8907), .ZN(n8909) );
  XNOR2_X1 U9998 ( .A(n8906), .B(n8909), .ZN(n8916) );
  OAI22_X1 U9999 ( .A1(n10066), .A2(n8911), .B1(n10083), .B2(n8910), .ZN(n8912) );
  AOI211_X1 U10000 ( .C1(n10086), .C2(n10404), .A(n8913), .B(n8912), .ZN(n8915) );
  NAND2_X1 U10001 ( .A1(n9210), .A2(n10069), .ZN(n8914) );
  OAI211_X1 U10002 ( .C1(n8916), .C2(n10071), .A(n8915), .B(n8914), .ZN(
        P1_U3222) );
  OAI21_X1 U10003 ( .B1(n8919), .B2(n8918), .A(n8917), .ZN(n8920) );
  NAND2_X1 U10004 ( .A1(n8920), .A2(n9341), .ZN(n8924) );
  NAND2_X1 U10005 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9413) );
  OAI21_X1 U10006 ( .B1(n9386), .B2(n9752), .A(n9413), .ZN(n8922) );
  OAI22_X1 U10007 ( .A1(n9508), .A2(n9371), .B1(n9372), .B2(n9718), .ZN(n8921)
         );
  AOI211_X1 U10008 ( .C1(n9888), .C2(n9389), .A(n8922), .B(n8921), .ZN(n8923)
         );
  NAND2_X1 U10009 ( .A1(n8924), .A2(n8923), .ZN(P2_U3243) );
  INV_X1 U10010 ( .A(n8948), .ZN(n9275) );
  OAI222_X1 U10011 ( .A1(n9923), .A2(n8926), .B1(n5076), .B2(n9275), .C1(
        P2_U3152), .C2(n8925), .ZN(P2_U3330) );
  INV_X1 U10012 ( .A(n8932), .ZN(n9273) );
  OAI222_X1 U10013 ( .A1(n9923), .A2(n8927), .B1(n5076), .B2(n9273), .C1(
        P2_U3152), .C2(n5726), .ZN(P2_U3328) );
  AND2_X1 U10014 ( .A1(n9167), .A2(n5073), .ZN(n9173) );
  INV_X1 U10015 ( .A(n9173), .ZN(n8928) );
  NOR2_X1 U10016 ( .A1(n8929), .A2(n8928), .ZN(n9185) );
  INV_X1 U10017 ( .A(n9018), .ZN(n9028) );
  NAND2_X1 U10018 ( .A1(n10539), .A2(n8947), .ZN(n8931) );
  OR2_X1 U10019 ( .A1(n8949), .A2(n7364), .ZN(n8930) );
  NAND2_X1 U10020 ( .A1(n8932), .A2(n8947), .ZN(n8934) );
  INV_X1 U10021 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9272) );
  OR2_X1 U10022 ( .A1(n8949), .A2(n9272), .ZN(n8933) );
  INV_X1 U10023 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n10164) );
  NAND2_X1 U10024 ( .A1(n6706), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8937) );
  INV_X1 U10025 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n8935) );
  OR2_X1 U10026 ( .A1(n8941), .A2(n8935), .ZN(n8936) );
  OAI211_X1 U10027 ( .C1(n8942), .C2(n10164), .A(n8937), .B(n8936), .ZN(n10090) );
  NAND2_X1 U10028 ( .A1(n10163), .A2(n10090), .ZN(n9030) );
  NAND2_X1 U10029 ( .A1(n9916), .A2(n8947), .ZN(n8939) );
  OR2_X1 U10030 ( .A1(n8949), .A2(n10541), .ZN(n8938) );
  NAND2_X1 U10031 ( .A1(n6706), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8946) );
  INV_X1 U10032 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8940) );
  OR2_X1 U10033 ( .A1(n8941), .A2(n8940), .ZN(n8945) );
  OR2_X1 U10034 ( .A1(n6781), .A2(n9265), .ZN(n8944) );
  INV_X1 U10035 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9266) );
  OR2_X1 U10036 ( .A1(n8942), .A2(n9266), .ZN(n8943) );
  NAND4_X1 U10037 ( .A1(n8946), .A2(n8945), .A3(n8944), .A4(n8943), .ZN(n10173) );
  INV_X1 U10038 ( .A(n10173), .ZN(n9016) );
  MUX2_X1 U10039 ( .A(n9256), .B(n9032), .S(n9018), .Z(n9015) );
  INV_X1 U10040 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9274) );
  OR2_X1 U10041 ( .A1(n8949), .A2(n9274), .ZN(n8950) );
  INV_X1 U10042 ( .A(n10197), .ZN(n9232) );
  NAND2_X1 U10043 ( .A1(n10454), .A2(n9232), .ZN(n9033) );
  INV_X1 U10044 ( .A(n10228), .ZN(n9971) );
  MUX2_X1 U10045 ( .A(n9254), .B(n9073), .S(n9018), .Z(n9013) );
  MUX2_X1 U10046 ( .A(n9253), .B(n9072), .S(n9028), .Z(n9011) );
  INV_X1 U10047 ( .A(n10260), .ZN(n9972) );
  OR2_X1 U10048 ( .A1(n10476), .A2(n9972), .ZN(n9008) );
  NAND2_X1 U10049 ( .A1(n9008), .A2(n10236), .ZN(n9251) );
  OR2_X1 U10050 ( .A1(n9252), .A2(n9250), .ZN(n8952) );
  MUX2_X1 U10051 ( .A(n9251), .B(n8952), .S(n9018), .Z(n9010) );
  INV_X1 U10052 ( .A(n10284), .ZN(n9961) );
  NAND2_X1 U10053 ( .A1(n10486), .A2(n9961), .ZN(n9249) );
  INV_X1 U10054 ( .A(n9249), .ZN(n8953) );
  MUX2_X1 U10055 ( .A(n8953), .B(n9248), .S(n9018), .Z(n8954) );
  NOR2_X1 U10056 ( .A1(n10250), .A2(n8954), .ZN(n9007) );
  INV_X1 U10057 ( .A(n10092), .ZN(n10298) );
  INV_X1 U10058 ( .A(n10283), .ZN(n10316) );
  OR2_X1 U10059 ( .A1(n10306), .A2(n10316), .ZN(n10279) );
  OR2_X1 U10060 ( .A1(n9247), .A2(n9246), .ZN(n8957) );
  NAND2_X1 U10061 ( .A1(n10306), .A2(n10316), .ZN(n9245) );
  INV_X1 U10062 ( .A(n9245), .ZN(n8955) );
  NAND2_X1 U10063 ( .A1(n8959), .A2(n8955), .ZN(n8956) );
  AND2_X1 U10064 ( .A1(n8958), .A2(n8956), .ZN(n9035) );
  MUX2_X1 U10065 ( .A(n8957), .B(n9035), .S(n9018), .Z(n9006) );
  XNOR2_X1 U10066 ( .A(n10486), .B(n10284), .ZN(n10266) );
  INV_X1 U10067 ( .A(n10281), .ZN(n9143) );
  INV_X1 U10068 ( .A(n10331), .ZN(n10297) );
  NAND2_X1 U10069 ( .A1(n10503), .A2(n10297), .ZN(n9036) );
  OR2_X1 U10070 ( .A1(n10503), .A2(n10297), .ZN(n9041) );
  MUX2_X1 U10071 ( .A(n9036), .B(n9041), .S(n9018), .Z(n9004) );
  INV_X1 U10072 ( .A(n10332), .ZN(n10371) );
  INV_X1 U10073 ( .A(n10348), .ZN(n10315) );
  INV_X1 U10074 ( .A(n10330), .ZN(n10326) );
  INV_X1 U10075 ( .A(n10349), .ZN(n10385) );
  NAND2_X1 U10076 ( .A1(n10513), .A2(n10385), .ZN(n10344) );
  INV_X1 U10077 ( .A(n10399), .ZN(n10370) );
  NAND2_X1 U10078 ( .A1(n10395), .A2(n10370), .ZN(n10363) );
  NAND2_X1 U10079 ( .A1(n10344), .A2(n10363), .ZN(n8960) );
  OR2_X1 U10080 ( .A1(n10513), .A2(n10385), .ZN(n9116) );
  NAND4_X1 U10081 ( .A1(n9240), .A2(n9028), .A3(n8960), .A4(n9116), .ZN(n8961)
         );
  OAI211_X1 U10082 ( .C1(n9028), .C2(n9240), .A(n10326), .B(n8961), .ZN(n9002)
         );
  MUX2_X1 U10083 ( .A(n10095), .B(n8962), .S(n9028), .Z(n8978) );
  XNOR2_X1 U10084 ( .A(n8963), .B(n9018), .ZN(n8967) );
  AND2_X1 U10085 ( .A1(n9102), .A2(n8969), .ZN(n8964) );
  MUX2_X1 U10086 ( .A(n8964), .B(n9100), .S(n9028), .Z(n8965) );
  MUX2_X1 U10087 ( .A(n8969), .B(n8968), .S(n9018), .Z(n8970) );
  MUX2_X1 U10088 ( .A(n9052), .B(n8971), .S(n9018), .Z(n8972) );
  MUX2_X1 U10089 ( .A(n8973), .B(n9051), .S(n9018), .Z(n8974) );
  INV_X1 U10090 ( .A(n8974), .ZN(n8975) );
  MUX2_X1 U10091 ( .A(n9045), .B(n9053), .S(n9028), .Z(n8976) );
  OAI211_X1 U10092 ( .C1(n9120), .C2(n8978), .A(n8977), .B(n8976), .ZN(n8981)
         );
  INV_X1 U10093 ( .A(n9137), .ZN(n8980) );
  NAND2_X1 U10094 ( .A1(n8978), .A2(n9118), .ZN(n8979) );
  NAND3_X1 U10095 ( .A1(n8981), .A2(n8980), .A3(n8979), .ZN(n8985) );
  NAND2_X1 U10096 ( .A1(n10413), .A2(n10425), .ZN(n9075) );
  NAND2_X1 U10097 ( .A1(n9060), .A2(n9075), .ZN(n10414) );
  AND2_X1 U10098 ( .A1(n10094), .A2(n9028), .ZN(n8983) );
  OAI21_X1 U10099 ( .B1(n9028), .B2(n10094), .A(n9210), .ZN(n8982) );
  OAI21_X1 U10100 ( .B1(n8983), .B2(n9210), .A(n8982), .ZN(n8984) );
  NAND3_X1 U10101 ( .A1(n8985), .A2(n5439), .A3(n8984), .ZN(n8987) );
  INV_X1 U10102 ( .A(n10404), .ZN(n9934) );
  OR2_X1 U10103 ( .A1(n10433), .A2(n9934), .ZN(n9059) );
  NAND2_X1 U10104 ( .A1(n10433), .A2(n9934), .ZN(n9237) );
  OR2_X1 U10105 ( .A1(n10414), .A2(n10420), .ZN(n8986) );
  NAND2_X1 U10106 ( .A1(n8987), .A2(n8986), .ZN(n8994) );
  INV_X1 U10107 ( .A(n9060), .ZN(n9238) );
  AOI21_X1 U10108 ( .B1(n8994), .B2(n9237), .A(n9238), .ZN(n8998) );
  NAND2_X1 U10109 ( .A1(n10356), .A2(n10371), .ZN(n9117) );
  NAND4_X1 U10110 ( .A1(n9117), .A2(n9018), .A3(n10363), .A4(n10344), .ZN(
        n8997) );
  NAND2_X1 U10111 ( .A1(n9116), .A2(n9239), .ZN(n9064) );
  NAND3_X1 U10112 ( .A1(n9064), .A2(n9018), .A3(n10344), .ZN(n8988) );
  NAND2_X1 U10113 ( .A1(n8988), .A2(n9117), .ZN(n8989) );
  OAI21_X1 U10114 ( .B1(n9028), .B2(n9117), .A(n8989), .ZN(n8996) );
  INV_X1 U10115 ( .A(n9075), .ZN(n8993) );
  INV_X1 U10116 ( .A(n9059), .ZN(n8990) );
  AOI21_X1 U10117 ( .B1(n9075), .B2(n8990), .A(n9018), .ZN(n8991) );
  AND4_X1 U10118 ( .A1(n9240), .A2(n8991), .A3(n9116), .A4(n9239), .ZN(n8992)
         );
  OAI21_X1 U10119 ( .B1(n8994), .B2(n8993), .A(n8992), .ZN(n8995) );
  OAI211_X1 U10120 ( .C1(n8998), .C2(n8997), .A(n8996), .B(n8995), .ZN(n9001)
         );
  NAND2_X1 U10121 ( .A1(n9041), .A2(n9036), .ZN(n10313) );
  INV_X1 U10122 ( .A(n10313), .ZN(n9000) );
  MUX2_X1 U10123 ( .A(n9038), .B(n9242), .S(n9018), .Z(n8999) );
  OAI211_X1 U10124 ( .C1(n9002), .C2(n9001), .A(n9000), .B(n8999), .ZN(n9003)
         );
  NAND4_X1 U10125 ( .A1(n9143), .A2(n10301), .A3(n9004), .A4(n9003), .ZN(n9005) );
  INV_X1 U10126 ( .A(n9252), .ZN(n10224) );
  MUX2_X1 U10127 ( .A(n9008), .B(n10224), .S(n9028), .Z(n9009) );
  NAND3_X1 U10128 ( .A1(n10195), .A2(n9013), .A3(n9012), .ZN(n9014) );
  NAND2_X1 U10129 ( .A1(n9114), .A2(n9257), .ZN(n9161) );
  OAI21_X1 U10130 ( .B1(n9161), .B2(n9017), .A(n9159), .ZN(n9019) );
  OAI21_X1 U10131 ( .B1(n10443), .B2(n9030), .A(n9020), .ZN(n9022) );
  NAND2_X1 U10132 ( .A1(n10159), .A2(n10090), .ZN(n9021) );
  NAND2_X1 U10133 ( .A1(n10444), .A2(n9021), .ZN(n9158) );
  MUX2_X1 U10134 ( .A(n9028), .B(n9022), .S(n9158), .Z(n9023) );
  INV_X1 U10135 ( .A(n10159), .ZN(n9024) );
  NAND2_X1 U10136 ( .A1(n9023), .A2(n9179), .ZN(n9029) );
  NAND2_X1 U10137 ( .A1(n9025), .A2(n9024), .ZN(n9031) );
  INV_X1 U10138 ( .A(n9030), .ZN(n9026) );
  NAND2_X1 U10139 ( .A1(n9026), .A2(n10159), .ZN(n9027) );
  NAND2_X1 U10140 ( .A1(n9027), .A2(n9031), .ZN(n9164) );
  NAND2_X1 U10141 ( .A1(n9031), .A2(n9030), .ZN(n9149) );
  INV_X1 U10142 ( .A(n9256), .ZN(n9034) );
  OAI211_X1 U10143 ( .C1(n9034), .C2(n9254), .A(n9033), .B(n9032), .ZN(n9157)
         );
  AND2_X1 U10144 ( .A1(n9035), .A2(n9249), .ZN(n9043) );
  INV_X1 U10145 ( .A(n9043), .ZN(n9037) );
  INV_X1 U10146 ( .A(n9036), .ZN(n9244) );
  OR2_X1 U10147 ( .A1(n9037), .A2(n9244), .ZN(n9081) );
  NAND2_X1 U10148 ( .A1(n9038), .A2(n9240), .ZN(n9039) );
  NAND2_X1 U10149 ( .A1(n9039), .A2(n9242), .ZN(n9040) );
  AND2_X1 U10150 ( .A1(n9041), .A2(n9040), .ZN(n9069) );
  INV_X1 U10151 ( .A(n9247), .ZN(n9042) );
  AOI21_X1 U10152 ( .B1(n9043), .B2(n9042), .A(n9248), .ZN(n9068) );
  NAND2_X1 U10153 ( .A1(n9045), .A2(n9044), .ZN(n9046) );
  NAND2_X1 U10154 ( .A1(n9046), .A2(n9053), .ZN(n9047) );
  NAND2_X1 U10155 ( .A1(n9048), .A2(n9047), .ZN(n9049) );
  NOR2_X1 U10156 ( .A1(n10419), .A2(n9049), .ZN(n9050) );
  AND2_X1 U10157 ( .A1(n9237), .A2(n9050), .ZN(n9077) );
  NAND3_X1 U10158 ( .A1(n5426), .A2(n9053), .A3(n9052), .ZN(n9054) );
  NAND2_X1 U10159 ( .A1(n9077), .A2(n9054), .ZN(n9061) );
  NAND2_X1 U10160 ( .A1(n9056), .A2(n9055), .ZN(n9235) );
  NAND3_X1 U10161 ( .A1(n9237), .A2(n9057), .A3(n9235), .ZN(n9058) );
  NAND4_X1 U10162 ( .A1(n9061), .A2(n9060), .A3(n9059), .A4(n9058), .ZN(n9062)
         );
  AND3_X1 U10163 ( .A1(n10363), .A2(n9075), .A3(n9062), .ZN(n9063) );
  NOR2_X1 U10164 ( .A1(n9064), .A2(n9063), .ZN(n9066) );
  AND2_X1 U10165 ( .A1(n9117), .A2(n10344), .ZN(n9065) );
  NAND2_X1 U10166 ( .A1(n9242), .A2(n9065), .ZN(n9079) );
  OR3_X1 U10167 ( .A1(n9081), .A2(n9066), .A3(n9079), .ZN(n9067) );
  OAI211_X1 U10168 ( .C1(n9081), .C2(n9069), .A(n9068), .B(n9067), .ZN(n9071)
         );
  AOI21_X1 U10169 ( .B1(n9071), .B2(n9070), .A(n9251), .ZN(n9074) );
  NAND2_X1 U10170 ( .A1(n9253), .A2(n10224), .ZN(n9082) );
  OAI211_X1 U10171 ( .C1(n9074), .C2(n9082), .A(n9073), .B(n9072), .ZN(n9154)
         );
  NAND4_X1 U10172 ( .A1(n10363), .A2(n9077), .A3(n9076), .A4(n9075), .ZN(n9078) );
  OR3_X1 U10173 ( .A1(n9250), .A2(n9079), .A3(n9078), .ZN(n9080) );
  OR3_X1 U10174 ( .A1(n9082), .A2(n9081), .A3(n9080), .ZN(n9152) );
  INV_X1 U10175 ( .A(n6736), .ZN(n10688) );
  NAND2_X1 U10176 ( .A1(n6735), .A2(n10688), .ZN(n9083) );
  NAND3_X1 U10177 ( .A1(n9084), .A2(n9169), .A3(n9083), .ZN(n9085) );
  NAND2_X1 U10178 ( .A1(n9086), .A2(n9085), .ZN(n9087) );
  OAI22_X1 U10179 ( .A1(n9088), .A2(n9087), .B1(n10743), .B2(n10720), .ZN(
        n9090) );
  NAND2_X1 U10180 ( .A1(n9090), .A2(n9089), .ZN(n9092) );
  OAI211_X1 U10181 ( .C1(n9094), .C2(n9093), .A(n9092), .B(n9091), .ZN(n9097)
         );
  NAND3_X1 U10182 ( .A1(n9097), .A2(n9096), .A3(n9095), .ZN(n9099) );
  NAND2_X1 U10183 ( .A1(n9099), .A2(n9098), .ZN(n9103) );
  INV_X1 U10184 ( .A(n9100), .ZN(n9101) );
  AOI21_X1 U10185 ( .B1(n9103), .B2(n9102), .A(n9101), .ZN(n9104) );
  NOR2_X1 U10186 ( .A1(n9152), .A2(n9104), .ZN(n9105) );
  NOR3_X1 U10187 ( .A1(n10188), .A2(n9154), .A3(n9105), .ZN(n9106) );
  NOR2_X1 U10188 ( .A1(n9157), .A2(n9106), .ZN(n9108) );
  INV_X1 U10189 ( .A(n10090), .ZN(n9107) );
  NAND2_X1 U10190 ( .A1(n10444), .A2(n9107), .ZN(n9147) );
  OAI211_X1 U10191 ( .C1(n9161), .C2(n9108), .A(n9159), .B(n9147), .ZN(n9109)
         );
  INV_X1 U10192 ( .A(n9109), .ZN(n9110) );
  OAI21_X1 U10193 ( .B1(n9149), .B2(n9110), .A(n9179), .ZN(n9111) );
  XNOR2_X1 U10194 ( .A(n9111), .B(n10289), .ZN(n9113) );
  NAND2_X1 U10195 ( .A1(n9113), .A2(n9112), .ZN(n9178) );
  INV_X1 U10196 ( .A(n10250), .ZN(n10258) );
  INV_X1 U10197 ( .A(n9228), .ZN(n9115) );
  NAND2_X1 U10198 ( .A1(n9116), .A2(n10344), .ZN(n10361) );
  INV_X1 U10199 ( .A(n10361), .ZN(n10365) );
  NAND2_X1 U10200 ( .A1(n9239), .A2(n10363), .ZN(n10384) );
  INV_X1 U10201 ( .A(n9118), .ZN(n9119) );
  OR2_X1 U10202 ( .A1(n9120), .A2(n9119), .ZN(n10886) );
  NOR2_X1 U10203 ( .A1(n9121), .A2(n10781), .ZN(n9126) );
  INV_X1 U10204 ( .A(n9122), .ZN(n9124) );
  NAND4_X1 U10205 ( .A1(n9126), .A2(n9125), .A3(n9124), .A4(n9123), .ZN(n9131)
         );
  NAND3_X1 U10206 ( .A1(n9129), .A2(n9128), .A3(n9127), .ZN(n9130) );
  NOR2_X1 U10207 ( .A1(n9131), .A2(n9130), .ZN(n9132) );
  NAND4_X1 U10208 ( .A1(n10886), .A2(n5113), .A3(n9133), .A4(n9132), .ZN(n9136) );
  INV_X1 U10209 ( .A(n9134), .ZN(n9135) );
  OR3_X1 U10210 ( .A1(n9137), .A2(n9136), .A3(n9135), .ZN(n9138) );
  INV_X1 U10211 ( .A(n10420), .ZN(n10427) );
  OR3_X1 U10212 ( .A1(n9138), .A2(n10414), .A3(n10427), .ZN(n9139) );
  NOR2_X1 U10213 ( .A1(n10384), .A2(n9139), .ZN(n9140) );
  NAND4_X1 U10214 ( .A1(n10326), .A2(n10365), .A3(n10357), .A4(n9140), .ZN(
        n9141) );
  NOR2_X1 U10215 ( .A1(n10313), .A2(n9141), .ZN(n9142) );
  AND4_X1 U10216 ( .A1(n10240), .A2(n9143), .A3(n9142), .A4(n10301), .ZN(n9144) );
  NAND4_X1 U10217 ( .A1(n10217), .A2(n10258), .A3(n9144), .A4(n10266), .ZN(
        n9145) );
  NOR2_X1 U10218 ( .A1(n10188), .A2(n9145), .ZN(n9146) );
  AND4_X1 U10219 ( .A1(n9258), .A2(n10171), .A3(n10205), .A4(n9146), .ZN(n9148) );
  NAND3_X1 U10220 ( .A1(n9148), .A2(n9179), .A3(n9147), .ZN(n9150) );
  NOR2_X1 U10221 ( .A1(n9150), .A2(n9149), .ZN(n9171) );
  INV_X1 U10222 ( .A(n9151), .ZN(n9153) );
  OAI21_X1 U10223 ( .B1(n9153), .B2(n9152), .A(n9256), .ZN(n9155) );
  NOR2_X1 U10224 ( .A1(n9155), .A2(n9154), .ZN(n9156) );
  NOR2_X1 U10225 ( .A1(n9157), .A2(n9156), .ZN(n9160) );
  OAI211_X1 U10226 ( .C1(n9161), .C2(n9160), .A(n9159), .B(n9158), .ZN(n9162)
         );
  INV_X1 U10227 ( .A(n9162), .ZN(n9163) );
  OR2_X1 U10228 ( .A1(n9164), .A2(n9163), .ZN(n9166) );
  AND2_X1 U10229 ( .A1(n9179), .A2(n9169), .ZN(n9165) );
  NAND2_X1 U10230 ( .A1(n9166), .A2(n9165), .ZN(n9170) );
  AND2_X1 U10231 ( .A1(n9167), .A2(n10289), .ZN(n9168) );
  NAND3_X1 U10232 ( .A1(n9171), .A2(n9170), .A3(n9168), .ZN(n9177) );
  NAND3_X1 U10233 ( .A1(n9170), .A2(n9169), .A3(n9168), .ZN(n9176) );
  INV_X1 U10234 ( .A(n9171), .ZN(n9174) );
  NAND3_X1 U10235 ( .A1(n9174), .A2(n9173), .A3(n9172), .ZN(n9175) );
  NAND4_X1 U10236 ( .A1(n9178), .A2(n9177), .A3(n9176), .A4(n9175), .ZN(n9183)
         );
  INV_X1 U10237 ( .A(n9179), .ZN(n9181) );
  AOI211_X1 U10238 ( .C1(n9185), .C2(n9184), .A(n9183), .B(n9182), .ZN(n9191)
         );
  NOR4_X1 U10239 ( .A1(n10889), .A2(n10623), .A3(n9186), .A4(n7264), .ZN(n9189) );
  OAI21_X1 U10240 ( .B1(n9187), .B2(n9190), .A(P1_B_REG_SCAN_IN), .ZN(n9188)
         );
  OAI22_X1 U10241 ( .A1(n9191), .A2(n9190), .B1(n9189), .B2(n9188), .ZN(
        P1_U3240) );
  NAND2_X1 U10242 ( .A1(n10454), .A2(n9192), .ZN(n9194) );
  NAND2_X1 U10243 ( .A1(n10197), .A2(n6719), .ZN(n9193) );
  NAND2_X1 U10244 ( .A1(n9194), .A2(n9193), .ZN(n9195) );
  XNOR2_X1 U10245 ( .A(n9195), .B(n6752), .ZN(n9198) );
  INV_X1 U10246 ( .A(n10454), .ZN(n9263) );
  AOI22_X1 U10247 ( .A1(n10454), .A2(n6719), .B1(n9196), .B2(n10197), .ZN(
        n9197) );
  XNOR2_X1 U10248 ( .A(n9198), .B(n9197), .ZN(n9203) );
  INV_X1 U10249 ( .A(n9203), .ZN(n9199) );
  NAND2_X1 U10250 ( .A1(n9199), .A2(n10078), .ZN(n9209) );
  NAND4_X1 U10251 ( .A1(n9208), .A2(n10078), .A3(n9202), .A4(n9203), .ZN(n9207) );
  AOI22_X1 U10252 ( .A1(n10081), .A2(n10174), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9201) );
  NAND2_X1 U10253 ( .A1(n10086), .A2(n10173), .ZN(n9200) );
  OAI211_X1 U10254 ( .C1(n10083), .C2(n10178), .A(n9201), .B(n9200), .ZN(n9205) );
  NOR3_X1 U10255 ( .A1(n9203), .A2(n10071), .A3(n9202), .ZN(n9204) );
  AOI211_X1 U10256 ( .C1(n10454), .C2(n10069), .A(n9205), .B(n9204), .ZN(n9206) );
  OAI211_X1 U10257 ( .C1(n9209), .C2(n9208), .A(n9207), .B(n9206), .ZN(
        P1_U3218) );
  NAND2_X1 U10258 ( .A1(n9210), .A2(n10094), .ZN(n9211) );
  OR2_X1 U10259 ( .A1(n10433), .A2(n10404), .ZN(n9213) );
  NAND2_X1 U10260 ( .A1(n10395), .A2(n10399), .ZN(n9214) );
  NAND2_X1 U10261 ( .A1(n10513), .A2(n10349), .ZN(n9216) );
  OR2_X1 U10262 ( .A1(n10356), .A2(n10332), .ZN(n9217) );
  NAND2_X1 U10263 ( .A1(n10356), .A2(n10332), .ZN(n9218) );
  NAND2_X1 U10264 ( .A1(n9219), .A2(n9218), .ZN(n10327) );
  NAND2_X1 U10265 ( .A1(n10506), .A2(n10348), .ZN(n9220) );
  OR2_X1 U10266 ( .A1(n10503), .A2(n10331), .ZN(n9221) );
  NAND2_X1 U10267 ( .A1(n10490), .A2(n10092), .ZN(n9222) );
  NAND2_X1 U10268 ( .A1(n10251), .A2(n10250), .ZN(n10234) );
  INV_X1 U10269 ( .A(n9224), .ZN(n9226) );
  NAND2_X1 U10270 ( .A1(n10479), .A2(n9225), .ZN(n10233) );
  NOR2_X1 U10271 ( .A1(n10464), .A2(n10228), .ZN(n9230) );
  NAND2_X1 U10272 ( .A1(n10464), .A2(n10228), .ZN(n9229) );
  INV_X1 U10273 ( .A(n10171), .ZN(n9231) );
  INV_X1 U10274 ( .A(n9258), .ZN(n9233) );
  XNOR2_X1 U10275 ( .A(n9234), .B(n9233), .ZN(n10452) );
  NAND2_X1 U10276 ( .A1(n10357), .A2(n10344), .ZN(n9241) );
  INV_X1 U10277 ( .A(n9242), .ZN(n9243) );
  INV_X1 U10278 ( .A(n9254), .ZN(n9255) );
  NAND2_X1 U10279 ( .A1(n10196), .A2(n10195), .ZN(n10194) );
  NAND2_X1 U10280 ( .A1(n10170), .A2(n9257), .ZN(n9259) );
  INV_X1 U10281 ( .A(P1_B_REG_SCAN_IN), .ZN(n9260) );
  OR2_X1 U10282 ( .A1(n7264), .A2(n9260), .ZN(n9261) );
  AND2_X1 U10283 ( .A1(n10398), .A2(n9261), .ZN(n10158) );
  AOI22_X1 U10284 ( .A1(n10405), .A2(n10197), .B1(n10090), .B2(n10158), .ZN(
        n9262) );
  NAND2_X1 U10285 ( .A1(n10448), .A2(n5074), .ZN(n9270) );
  INV_X1 U10286 ( .A(n10479), .ZN(n10257) );
  INV_X1 U10287 ( .A(n10490), .ZN(n10286) );
  INV_X1 U10288 ( .A(n10395), .ZN(n11004) );
  OR2_X2 U10289 ( .A1(n10392), .A2(n10513), .ZN(n10352) );
  OR2_X2 U10290 ( .A1(n10352), .A2(n10356), .ZN(n10353) );
  INV_X1 U10291 ( .A(n10503), .ZN(n10319) );
  INV_X1 U10292 ( .A(n10306), .ZN(n10496) );
  NOR2_X2 U10293 ( .A1(n10449), .A2(n10183), .ZN(n10162) );
  AOI21_X1 U10294 ( .B1(n10449), .B2(n10183), .A(n10162), .ZN(n10450) );
  INV_X1 U10295 ( .A(n10449), .ZN(n9264) );
  NOR2_X1 U10296 ( .A1(n9264), .A2(n10905), .ZN(n9268) );
  OAI22_X1 U10297 ( .A1(n5074), .A2(n9266), .B1(n9265), .B2(n10907), .ZN(n9267) );
  AOI211_X1 U10298 ( .C1(n10450), .C2(n10902), .A(n9268), .B(n9267), .ZN(n9269) );
  OAI211_X1 U10299 ( .C1(n10381), .C2(n10452), .A(n9270), .B(n9269), .ZN(
        P1_U3355) );
  OAI222_X1 U10300 ( .A1(n9271), .A2(P1_U3084), .B1(n8088), .B2(n9273), .C1(
        n9272), .C2(n10546), .ZN(P1_U3323) );
  OAI222_X1 U10301 ( .A1(n7202), .A2(P1_U3084), .B1(n8088), .B2(n9275), .C1(
        n9274), .C2(n10546), .ZN(P1_U3325) );
  XNOR2_X1 U10302 ( .A(n9277), .B(n9276), .ZN(n9283) );
  INV_X1 U10303 ( .A(n9633), .ZN(n9279) );
  OAI22_X1 U10304 ( .A1(n9386), .A2(n9279), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9278), .ZN(n9281) );
  OAI22_X1 U10305 ( .A1(n9512), .A2(n9371), .B1(n9372), .B2(n9518), .ZN(n9280)
         );
  AOI211_X1 U10306 ( .C1(n9846), .C2(n9389), .A(n9281), .B(n9280), .ZN(n9282)
         );
  OAI21_X1 U10307 ( .B1(n9283), .B2(n9391), .A(n9282), .ZN(P2_U3218) );
  XNOR2_X1 U10308 ( .A(n9285), .B(n9284), .ZN(n9289) );
  NAND2_X1 U10309 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9489) );
  OAI21_X1 U10310 ( .B1(n9386), .B2(n9696), .A(n9489), .ZN(n9287) );
  OAI22_X1 U10311 ( .A1(n9719), .A2(n9371), .B1(n9372), .B2(n9692), .ZN(n9286)
         );
  AOI211_X1 U10312 ( .C1(n9868), .C2(n9389), .A(n9287), .B(n9286), .ZN(n9288)
         );
  OAI21_X1 U10313 ( .B1(n9289), .B2(n9391), .A(n9288), .ZN(P2_U3221) );
  INV_X1 U10314 ( .A(n9290), .ZN(n9291) );
  INV_X1 U10315 ( .A(n9819), .ZN(n9550) );
  NAND2_X1 U10316 ( .A1(n9525), .A2(n9295), .ZN(n9297) );
  MUX2_X1 U10317 ( .A(n9297), .B(n9525), .S(n9296), .Z(n9300) );
  NOR3_X1 U10318 ( .A1(n9550), .A2(n9300), .A3(n9389), .ZN(n9298) );
  AOI21_X1 U10319 ( .B1(n9550), .B2(n9300), .A(n9298), .ZN(n9303) );
  NAND3_X1 U10320 ( .A1(n9819), .A2(n9335), .A3(n9300), .ZN(n9299) );
  OAI21_X1 U10321 ( .B1(n9300), .B2(n9819), .A(n9299), .ZN(n9302) );
  NAND2_X1 U10322 ( .A1(n9819), .A2(n9389), .ZN(n9301) );
  OR2_X1 U10323 ( .A1(n9304), .A2(n9720), .ZN(n9306) );
  NAND2_X1 U10324 ( .A1(n9393), .A2(n10924), .ZN(n9305) );
  NAND2_X1 U10325 ( .A1(n9306), .A2(n9305), .ZN(n9542) );
  AOI22_X1 U10326 ( .A1(n9542), .A2(n9384), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n9307) );
  OAI211_X1 U10327 ( .C1(n9547), .C2(n9386), .A(n9308), .B(n9307), .ZN(
        P2_U3222) );
  XNOR2_X1 U10328 ( .A(n9310), .B(n9309), .ZN(n9315) );
  OAI22_X1 U10329 ( .A1(n9386), .A2(n9660), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9311), .ZN(n9313) );
  OAI22_X1 U10330 ( .A1(n9692), .A2(n9371), .B1(n9372), .B2(n9512), .ZN(n9312)
         );
  AOI211_X1 U10331 ( .C1(n9856), .C2(n9389), .A(n9313), .B(n9312), .ZN(n9314)
         );
  OAI21_X1 U10332 ( .B1(n9315), .B2(n9391), .A(n9314), .ZN(P2_U3225) );
  NAND2_X1 U10333 ( .A1(n9317), .A2(n9316), .ZN(n9319) );
  XNOR2_X1 U10334 ( .A(n9319), .B(n9318), .ZN(n9326) );
  OR2_X1 U10335 ( .A1(n9565), .A2(n9720), .ZN(n9321) );
  INV_X1 U10336 ( .A(n9518), .ZN(n9622) );
  NAND2_X1 U10337 ( .A1(n9622), .A2(n10924), .ZN(n9320) );
  AND2_X1 U10338 ( .A1(n9321), .A2(n9320), .ZN(n9589) );
  INV_X1 U10339 ( .A(n9589), .ZN(n9322) );
  AOI22_X1 U10340 ( .A1(n9322), .A2(n9384), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n9323) );
  OAI21_X1 U10341 ( .B1(n9594), .B2(n9386), .A(n9323), .ZN(n9324) );
  AOI21_X1 U10342 ( .B1(n9836), .B2(n9389), .A(n9324), .ZN(n9325) );
  OAI21_X1 U10343 ( .B1(n9326), .B2(n9391), .A(n9325), .ZN(P2_U3227) );
  INV_X1 U10344 ( .A(n9883), .ZN(n9336) );
  OAI21_X1 U10345 ( .B1(n9329), .B2(n9328), .A(n9327), .ZN(n9330) );
  NAND2_X1 U10346 ( .A1(n9330), .A2(n9341), .ZN(n9334) );
  OR2_X1 U10347 ( .A1(n9395), .A2(n9720), .ZN(n9331) );
  OAI21_X1 U10348 ( .B1(n9396), .B2(n9774), .A(n9331), .ZN(n9738) );
  AND2_X1 U10349 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9437) );
  NOR2_X1 U10350 ( .A1(n9386), .A2(n9735), .ZN(n9332) );
  AOI211_X1 U10351 ( .C1(n9384), .C2(n9738), .A(n9437), .B(n9332), .ZN(n9333)
         );
  OAI211_X1 U10352 ( .C1(n9336), .C2(n9335), .A(n9334), .B(n9333), .ZN(
        P2_U3228) );
  OAI21_X1 U10353 ( .B1(n5508), .B2(n9339), .A(n9338), .ZN(n9340) );
  OAI211_X1 U10354 ( .C1(n9342), .C2(n5508), .A(n9341), .B(n9340), .ZN(n9346)
         );
  OAI22_X1 U10355 ( .A1(n9386), .A2(n9725), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9451), .ZN(n9344) );
  OAI22_X1 U10356 ( .A1(n9719), .A2(n9372), .B1(n9371), .B2(n9718), .ZN(n9343)
         );
  AOI211_X1 U10357 ( .C1(n9878), .C2(n9389), .A(n9344), .B(n9343), .ZN(n9345)
         );
  NAND2_X1 U10358 ( .A1(n9346), .A2(n9345), .ZN(P2_U3230) );
  XNOR2_X1 U10359 ( .A(n9348), .B(n9347), .ZN(n9353) );
  OAI22_X1 U10360 ( .A1(n9386), .A2(n9604), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9349), .ZN(n9351) );
  OAI22_X1 U10361 ( .A1(n9613), .A2(n9371), .B1(n9372), .B2(n9614), .ZN(n9350)
         );
  AOI211_X1 U10362 ( .C1(n9839), .C2(n9389), .A(n9351), .B(n9350), .ZN(n9352)
         );
  OAI21_X1 U10363 ( .B1(n9353), .B2(n9391), .A(n9352), .ZN(P2_U3231) );
  XNOR2_X1 U10364 ( .A(n9355), .B(n9354), .ZN(n9360) );
  OAI22_X1 U10365 ( .A1(n9386), .A2(n9678), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9356), .ZN(n9358) );
  OAI22_X1 U10366 ( .A1(n9373), .A2(n9371), .B1(n9372), .B2(n9364), .ZN(n9357)
         );
  AOI211_X1 U10367 ( .C1(n9861), .C2(n9389), .A(n9358), .B(n9357), .ZN(n9359)
         );
  OAI21_X1 U10368 ( .B1(n9360), .B2(n9391), .A(n9359), .ZN(P2_U3235) );
  AOI21_X1 U10369 ( .B1(n9362), .B2(n9361), .A(n5172), .ZN(n9368) );
  OAI22_X1 U10370 ( .A1(n9386), .A2(n9643), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9363), .ZN(n9366) );
  OAI22_X1 U10371 ( .A1(n9364), .A2(n9371), .B1(n9372), .B2(n9613), .ZN(n9365)
         );
  AOI211_X1 U10372 ( .C1(n9851), .C2(n9389), .A(n9366), .B(n9365), .ZN(n9367)
         );
  OAI21_X1 U10373 ( .B1(n9368), .B2(n9391), .A(n9367), .ZN(P2_U3237) );
  XNOR2_X1 U10374 ( .A(n9370), .B(n9369), .ZN(n9377) );
  NAND2_X1 U10375 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9457) );
  OAI21_X1 U10376 ( .B1(n9386), .B2(n9703), .A(n9457), .ZN(n9375) );
  OAI22_X1 U10377 ( .A1(n9373), .A2(n9372), .B1(n9371), .B2(n9395), .ZN(n9374)
         );
  AOI211_X1 U10378 ( .C1(n9871), .C2(n9389), .A(n9375), .B(n9374), .ZN(n9376)
         );
  OAI21_X1 U10379 ( .B1(n9377), .B2(n9391), .A(n9376), .ZN(P2_U3240) );
  AND2_X1 U10380 ( .A1(n9379), .A2(n9378), .ZN(n9381) );
  XNOR2_X1 U10381 ( .A(n9381), .B(n9380), .ZN(n9392) );
  INV_X1 U10382 ( .A(n9581), .ZN(n9387) );
  NAND2_X1 U10383 ( .A1(n9393), .A2(n10926), .ZN(n9383) );
  INV_X1 U10384 ( .A(n9614), .ZN(n9394) );
  NAND2_X1 U10385 ( .A1(n9394), .A2(n10924), .ZN(n9382) );
  NAND2_X1 U10386 ( .A1(n9383), .A2(n9382), .ZN(n9578) );
  AOI22_X1 U10387 ( .A1(n9578), .A2(n9384), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n9385) );
  OAI21_X1 U10388 ( .B1(n9387), .B2(n9386), .A(n9385), .ZN(n9388) );
  AOI21_X1 U10389 ( .B1(n9830), .B2(n9389), .A(n9388), .ZN(n9390) );
  OAI21_X1 U10390 ( .B1(n9392), .B2(n9391), .A(n9390), .ZN(P2_U3242) );
  MUX2_X1 U10391 ( .A(n9525), .B(P2_DATAO_REG_28__SCAN_IN), .S(n9406), .Z(
        P2_U3580) );
  MUX2_X1 U10392 ( .A(n9393), .B(P2_DATAO_REG_27__SCAN_IN), .S(n9406), .Z(
        P2_U3579) );
  MUX2_X1 U10393 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n9394), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U10394 ( .A(n9622), .B(P2_DATAO_REG_24__SCAN_IN), .S(n9406), .Z(
        P2_U3576) );
  INV_X1 U10395 ( .A(n9613), .ZN(n9650) );
  MUX2_X1 U10396 ( .A(n9650), .B(P2_DATAO_REG_23__SCAN_IN), .S(n9406), .Z(
        P2_U3575) );
  MUX2_X1 U10397 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9667), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U10398 ( .A(n9673), .B(P2_DATAO_REG_21__SCAN_IN), .S(n9406), .Z(
        P2_U3573) );
  INV_X1 U10399 ( .A(n9692), .ZN(n9668) );
  MUX2_X1 U10400 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9668), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U10401 ( .A(n5455), .B(P2_DATAO_REG_19__SCAN_IN), .S(n9406), .Z(
        P2_U3571) );
  INV_X1 U10402 ( .A(n9395), .ZN(n9709) );
  MUX2_X1 U10403 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9709), .S(P2_U3966), .Z(
        P2_U3569) );
  INV_X1 U10404 ( .A(n9718), .ZN(n9759) );
  MUX2_X1 U10405 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9759), .S(P2_U3966), .Z(
        P2_U3568) );
  INV_X1 U10406 ( .A(n9396), .ZN(n9771) );
  MUX2_X1 U10407 ( .A(n9771), .B(P2_DATAO_REG_15__SCAN_IN), .S(n9406), .Z(
        P2_U3567) );
  INV_X1 U10408 ( .A(n9775), .ZN(n9397) );
  MUX2_X1 U10409 ( .A(n9397), .B(P2_DATAO_REG_13__SCAN_IN), .S(n9406), .Z(
        P2_U3565) );
  INV_X1 U10410 ( .A(n9398), .ZN(n10927) );
  MUX2_X1 U10411 ( .A(n10927), .B(P2_DATAO_REG_12__SCAN_IN), .S(n9406), .Z(
        P2_U3564) );
  INV_X1 U10412 ( .A(n9399), .ZN(n9400) );
  MUX2_X1 U10413 ( .A(n9400), .B(P2_DATAO_REG_11__SCAN_IN), .S(n9406), .Z(
        P2_U3563) );
  MUX2_X1 U10414 ( .A(n10925), .B(P2_DATAO_REG_10__SCAN_IN), .S(n9406), .Z(
        P2_U3562) );
  MUX2_X1 U10415 ( .A(n9401), .B(P2_DATAO_REG_8__SCAN_IN), .S(n9406), .Z(
        P2_U3560) );
  MUX2_X1 U10416 ( .A(n9788), .B(P2_DATAO_REG_7__SCAN_IN), .S(n9406), .Z(
        P2_U3559) );
  MUX2_X1 U10417 ( .A(n9402), .B(P2_DATAO_REG_6__SCAN_IN), .S(n9406), .Z(
        P2_U3558) );
  MUX2_X1 U10418 ( .A(n9789), .B(P2_DATAO_REG_5__SCAN_IN), .S(n9406), .Z(
        P2_U3557) );
  MUX2_X1 U10419 ( .A(n9403), .B(P2_DATAO_REG_4__SCAN_IN), .S(n9406), .Z(
        P2_U3556) );
  MUX2_X1 U10420 ( .A(n9404), .B(P2_DATAO_REG_3__SCAN_IN), .S(n9406), .Z(
        P2_U3555) );
  MUX2_X1 U10421 ( .A(n9405), .B(P2_DATAO_REG_2__SCAN_IN), .S(n9406), .Z(
        P2_U3554) );
  MUX2_X1 U10422 ( .A(n9407), .B(P2_DATAO_REG_1__SCAN_IN), .S(n9406), .Z(
        P2_U3553) );
  MUX2_X1 U10423 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n9408), .S(P2_U3966), .Z(
        P2_U3552) );
  OAI21_X1 U10424 ( .B1(n9410), .B2(P2_REG2_REG_14__SCAN_IN), .A(n9409), .ZN(
        n9428) );
  XOR2_X1 U10425 ( .A(n9429), .B(n9428), .Z(n9411) );
  NAND2_X1 U10426 ( .A1(n9411), .A2(n6015), .ZN(n9430) );
  OAI21_X1 U10427 ( .B1(n9411), .B2(n6015), .A(n9430), .ZN(n9412) );
  INV_X1 U10428 ( .A(n9412), .ZN(n9421) );
  INV_X1 U10429 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n9414) );
  OAI21_X1 U10430 ( .B1(n10641), .B2(n9414), .A(n9413), .ZN(n9415) );
  AOI21_X1 U10431 ( .B1(n9423), .B2(n10649), .A(n9415), .ZN(n9420) );
  AOI21_X1 U10432 ( .B1(n9417), .B2(n5994), .A(n9416), .ZN(n9422) );
  XNOR2_X1 U10433 ( .A(n9422), .B(n9429), .ZN(n9418) );
  NAND2_X1 U10434 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n9418), .ZN(n9424) );
  OAI211_X1 U10435 ( .C1(n9418), .C2(P2_REG1_REG_15__SCAN_IN), .A(n10652), .B(
        n9424), .ZN(n9419) );
  OAI211_X1 U10436 ( .C1(n9421), .C2(n10642), .A(n9420), .B(n9419), .ZN(
        P2_U3260) );
  NAND2_X1 U10437 ( .A1(n9423), .A2(n9422), .ZN(n9425) );
  NAND2_X1 U10438 ( .A1(n9425), .A2(n9424), .ZN(n9427) );
  XNOR2_X1 U10439 ( .A(n9442), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n9426) );
  NOR2_X1 U10440 ( .A1(n9427), .A2(n9426), .ZN(n9446) );
  AOI21_X1 U10441 ( .B1(n9427), .B2(n9426), .A(n9446), .ZN(n9440) );
  NAND2_X1 U10442 ( .A1(n9429), .A2(n9428), .ZN(n9431) );
  NAND2_X1 U10443 ( .A1(n9431), .A2(n9430), .ZN(n9434) );
  AOI22_X1 U10444 ( .A1(n9442), .A2(n9432), .B1(P2_REG2_REG_16__SCAN_IN), .B2(
        n9448), .ZN(n9433) );
  NOR2_X1 U10445 ( .A1(n9434), .A2(n9433), .ZN(n9441) );
  AOI211_X1 U10446 ( .C1(n9434), .C2(n9433), .A(n9441), .B(n10642), .ZN(n9435)
         );
  INV_X1 U10447 ( .A(n9435), .ZN(n9439) );
  NOR2_X1 U10448 ( .A1(n9490), .A2(n9448), .ZN(n9436) );
  AOI211_X1 U10449 ( .C1(n9487), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n9437), .B(
        n9436), .ZN(n9438) );
  OAI211_X1 U10450 ( .C1(n9440), .C2(n9464), .A(n9439), .B(n9438), .ZN(
        P2_U3261) );
  AOI21_X1 U10451 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n9442), .A(n9441), .ZN(
        n9445) );
  NAND2_X1 U10452 ( .A1(n9469), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n9443) );
  OAI21_X1 U10453 ( .B1(n9469), .B2(P2_REG2_REG_17__SCAN_IN), .A(n9443), .ZN(
        n9444) );
  NOR2_X1 U10454 ( .A1(n9445), .A2(n9444), .ZN(n9468) );
  AOI211_X1 U10455 ( .C1(n9445), .C2(n9444), .A(n9468), .B(n10642), .ZN(n9456)
         );
  XNOR2_X1 U10456 ( .A(n9459), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n9450) );
  AOI21_X1 U10457 ( .B1(n9448), .B2(n9447), .A(n9446), .ZN(n9449) );
  NAND2_X1 U10458 ( .A1(n9450), .A2(n9449), .ZN(n9458) );
  OAI211_X1 U10459 ( .C1(n9450), .C2(n9449), .A(n10652), .B(n9458), .ZN(n9454)
         );
  NOR2_X1 U10460 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9451), .ZN(n9452) );
  AOI21_X1 U10461 ( .B1(n9487), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n9452), .ZN(
        n9453) );
  OAI211_X1 U10462 ( .C1(n9490), .C2(n9459), .A(n9454), .B(n9453), .ZN(n9455)
         );
  OR2_X1 U10463 ( .A1(n9456), .A2(n9455), .ZN(P2_U3262) );
  INV_X1 U10464 ( .A(n9479), .ZN(n9477) );
  INV_X1 U10465 ( .A(n9457), .ZN(n9467) );
  OAI21_X1 U10466 ( .B1(n9460), .B2(n9459), .A(n9458), .ZN(n9463) );
  NAND2_X1 U10467 ( .A1(n9477), .A2(n9461), .ZN(n9481) );
  OAI21_X1 U10468 ( .B1(n9477), .B2(n9461), .A(n9481), .ZN(n9462) );
  NOR2_X1 U10469 ( .A1(n9462), .A2(n9463), .ZN(n9483) );
  AOI21_X1 U10470 ( .B1(n9463), .B2(n9462), .A(n9483), .ZN(n9465) );
  NOR2_X1 U10471 ( .A1(n9465), .A2(n9464), .ZN(n9466) );
  AOI211_X1 U10472 ( .C1(n9487), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n9467), .B(
        n9466), .ZN(n9476) );
  MUX2_X1 U10473 ( .A(n6070), .B(P2_REG2_REG_18__SCAN_IN), .S(n9479), .Z(n9470) );
  INV_X1 U10474 ( .A(n9470), .ZN(n9471) );
  OAI21_X1 U10475 ( .B1(n9472), .B2(n9471), .A(n9478), .ZN(n9473) );
  NAND2_X1 U10476 ( .A1(n9474), .A2(n9473), .ZN(n9475) );
  OAI211_X1 U10477 ( .C1(n9490), .C2(n9477), .A(n9476), .B(n9475), .ZN(
        P2_U3263) );
  MUX2_X1 U10478 ( .A(n6093), .B(P2_REG2_REG_19__SCAN_IN), .S(n9742), .Z(n9480) );
  INV_X1 U10479 ( .A(n9481), .ZN(n9482) );
  NOR2_X1 U10480 ( .A1(n9483), .A2(n9482), .ZN(n9486) );
  XNOR2_X1 U10481 ( .A(n9742), .B(n9484), .ZN(n9485) );
  XNOR2_X1 U10482 ( .A(n9486), .B(n9485), .ZN(n9492) );
  NAND2_X1 U10483 ( .A1(n9487), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n9488) );
  OAI211_X1 U10484 ( .C1(n9490), .C2(n9742), .A(n9489), .B(n9488), .ZN(n9491)
         );
  AOI21_X1 U10485 ( .B1(n9492), .B2(n10652), .A(n9491), .ZN(n9493) );
  OAI21_X1 U10486 ( .B1(n10642), .B2(n9494), .A(n9493), .ZN(P2_U3264) );
  INV_X1 U10487 ( .A(n9846), .ZN(n9635) );
  INV_X1 U10488 ( .A(n9871), .ZN(n9706) );
  NAND2_X1 U10489 ( .A1(n9778), .A2(n10990), .ZN(n9780) );
  OR2_X2 U10490 ( .A1(n9750), .A2(n9883), .ZN(n9733) );
  NAND2_X1 U10491 ( .A1(n9663), .A2(n9682), .ZN(n9657) );
  NOR2_X2 U10492 ( .A1(n9657), .A2(n9851), .ZN(n9642) );
  NAND2_X1 U10493 ( .A1(n9561), .A2(n9580), .ZN(n9556) );
  NAND2_X1 U10494 ( .A1(n9815), .A2(n9546), .ZN(n9534) );
  XNOR2_X1 U10495 ( .A(n9502), .B(n9499), .ZN(n9807) );
  NAND2_X1 U10496 ( .A1(n9496), .A2(P2_B_REG_SCAN_IN), .ZN(n9497) );
  NAND2_X1 U10497 ( .A1(n10926), .A2(n9497), .ZN(n9533) );
  NOR2_X1 U10498 ( .A1(n9498), .A2(n9533), .ZN(n9804) );
  INV_X1 U10499 ( .A(n9804), .ZN(n9810) );
  NOR2_X1 U10500 ( .A1(n10949), .A2(n9810), .ZN(n9504) );
  NOR2_X1 U10501 ( .A1(n9499), .A2(n10705), .ZN(n9500) );
  AOI211_X1 U10502 ( .C1(n10949), .C2(P2_REG2_REG_31__SCAN_IN), .A(n9504), .B(
        n9500), .ZN(n9501) );
  OAI21_X1 U10503 ( .B1(n9807), .B2(n10702), .A(n9501), .ZN(P2_U3265) );
  INV_X1 U10504 ( .A(n9503), .ZN(n9812) );
  INV_X1 U10505 ( .A(n9502), .ZN(n9809) );
  NAND2_X1 U10506 ( .A1(n9534), .A2(n9503), .ZN(n9808) );
  NAND3_X1 U10507 ( .A1(n9809), .A2(n9763), .A3(n9808), .ZN(n9506) );
  AOI21_X1 U10508 ( .B1(n10949), .B2(P2_REG2_REG_30__SCAN_IN), .A(n9504), .ZN(
        n9505) );
  OAI211_X1 U10509 ( .C1(n9812), .C2(n10705), .A(n9506), .B(n9505), .ZN(
        P2_U3266) );
  OAI22_X1 U10510 ( .A1(n9749), .A2(n9756), .B1(n9771), .B2(n9888), .ZN(n9744)
         );
  NAND2_X1 U10511 ( .A1(n9688), .A2(n9689), .ZN(n9687) );
  NAND2_X1 U10512 ( .A1(n9868), .A2(n5455), .ZN(n9510) );
  NAND2_X1 U10513 ( .A1(n9687), .A2(n9510), .ZN(n9677) );
  NAND2_X1 U10514 ( .A1(n9861), .A2(n9668), .ZN(n9511) );
  INV_X1 U10515 ( .A(n9851), .ZN(n9646) );
  NAND2_X1 U10516 ( .A1(n9646), .A2(n9512), .ZN(n9514) );
  INV_X1 U10517 ( .A(n9514), .ZN(n9513) );
  INV_X1 U10518 ( .A(n9628), .ZN(n9516) );
  AND2_X1 U10519 ( .A1(n9639), .A2(n9514), .ZN(n9515) );
  NAND2_X1 U10520 ( .A1(n9607), .A2(n9518), .ZN(n9519) );
  NAND2_X1 U10521 ( .A1(n9598), .A2(n9614), .ZN(n9521) );
  NAND2_X1 U10522 ( .A1(n9555), .A2(n9563), .ZN(n9524) );
  NAND2_X1 U10523 ( .A1(n9561), .A2(n9522), .ZN(n9523) );
  NOR2_X1 U10524 ( .A1(n9819), .A2(n9525), .ZN(n9526) );
  AOI21_X1 U10525 ( .B1(n9545), .B2(n9544), .A(n9526), .ZN(n9527) );
  XNOR2_X1 U10526 ( .A(n9527), .B(n9528), .ZN(n9814) );
  INV_X1 U10527 ( .A(n9814), .ZN(n9540) );
  INV_X1 U10528 ( .A(n9528), .ZN(n9529) );
  XNOR2_X1 U10529 ( .A(n9530), .B(n9529), .ZN(n9531) );
  OAI222_X1 U10530 ( .A1(n9533), .A2(n9532), .B1(n9531), .B2(n9717), .C1(n9774), .C2(n9566), .ZN(n9817) );
  NOR2_X1 U10531 ( .A1(n9816), .A2(n10702), .ZN(n9538) );
  INV_X1 U10532 ( .A(n10700), .ZN(n10938) );
  AOI22_X1 U10533 ( .A1(n10949), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n9535), 
        .B2(n10938), .ZN(n9536) );
  OAI21_X1 U10534 ( .B1(n9815), .B2(n10705), .A(n9536), .ZN(n9537) );
  AOI211_X1 U10535 ( .C1(n9817), .C2(n10947), .A(n9538), .B(n9537), .ZN(n9539)
         );
  OAI21_X1 U10536 ( .B1(n9540), .B2(n10706), .A(n9539), .ZN(P2_U3267) );
  XNOR2_X1 U10537 ( .A(n9541), .B(n9544), .ZN(n9543) );
  XNOR2_X1 U10538 ( .A(n9545), .B(n9544), .ZN(n9818) );
  NAND2_X1 U10539 ( .A1(n9818), .A2(n9800), .ZN(n9553) );
  AOI21_X1 U10540 ( .B1(n9819), .B2(n9556), .A(n9546), .ZN(n9820) );
  INV_X1 U10541 ( .A(n9547), .ZN(n9548) );
  AOI22_X1 U10542 ( .A1(n10949), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n9548), 
        .B2(n10938), .ZN(n9549) );
  OAI21_X1 U10543 ( .B1(n9550), .B2(n10705), .A(n9549), .ZN(n9551) );
  AOI21_X1 U10544 ( .B1(n9820), .B2(n9763), .A(n9551), .ZN(n9552) );
  OAI211_X1 U10545 ( .C1(n9822), .C2(n10949), .A(n9553), .B(n9552), .ZN(
        P2_U3268) );
  XNOR2_X1 U10546 ( .A(n9555), .B(n9554), .ZN(n9828) );
  INV_X1 U10547 ( .A(n9580), .ZN(n9558) );
  INV_X1 U10548 ( .A(n9556), .ZN(n9557) );
  AOI21_X1 U10549 ( .B1(n9824), .B2(n9558), .A(n9557), .ZN(n9825) );
  AOI22_X1 U10550 ( .A1(n10949), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n9559), 
        .B2(n10938), .ZN(n9560) );
  OAI21_X1 U10551 ( .B1(n9561), .B2(n10705), .A(n9560), .ZN(n9571) );
  INV_X1 U10552 ( .A(n9562), .ZN(n9564) );
  AOI21_X1 U10553 ( .B1(n9564), .B2(n9563), .A(n9717), .ZN(n9569) );
  OAI22_X1 U10554 ( .A1(n9566), .A2(n9720), .B1(n9565), .B2(n9774), .ZN(n9567)
         );
  AOI21_X1 U10555 ( .B1(n9569), .B2(n9568), .A(n9567), .ZN(n9827) );
  NOR2_X1 U10556 ( .A1(n9827), .A2(n10949), .ZN(n9570) );
  AOI211_X1 U10557 ( .C1(n9825), .C2(n9763), .A(n9571), .B(n9570), .ZN(n9572)
         );
  OAI21_X1 U10558 ( .B1(n9828), .B2(n10706), .A(n9572), .ZN(P2_U3269) );
  XOR2_X1 U10559 ( .A(n9576), .B(n9573), .Z(n9833) );
  NOR2_X1 U10560 ( .A1(n5335), .A2(n10705), .ZN(n9584) );
  NAND2_X1 U10561 ( .A1(n9574), .A2(n9575), .ZN(n9577) );
  XNOR2_X1 U10562 ( .A(n9577), .B(n9576), .ZN(n9579) );
  AOI21_X1 U10563 ( .B1(n9579), .B2(n10929), .A(n9578), .ZN(n9832) );
  AOI211_X1 U10564 ( .C1(n9830), .C2(n9591), .A(n10991), .B(n9580), .ZN(n9829)
         );
  AOI22_X1 U10565 ( .A1(n9829), .A2(n9742), .B1(n10938), .B2(n9581), .ZN(n9582) );
  AOI21_X1 U10566 ( .B1(n9832), .B2(n9582), .A(n10949), .ZN(n9583) );
  AOI211_X1 U10567 ( .C1(n10949), .C2(P2_REG2_REG_26__SCAN_IN), .A(n9584), .B(
        n9583), .ZN(n9585) );
  OAI21_X1 U10568 ( .B1(n9833), .B2(n10706), .A(n9585), .ZN(P2_U3270) );
  XNOR2_X1 U10569 ( .A(n9586), .B(n9588), .ZN(n9838) );
  OAI211_X1 U10570 ( .C1(n9588), .C2(n9587), .A(n9574), .B(n10929), .ZN(n9590)
         );
  NAND2_X1 U10571 ( .A1(n9590), .A2(n9589), .ZN(n9834) );
  INV_X1 U10572 ( .A(n9591), .ZN(n9592) );
  AOI211_X1 U10573 ( .C1(n9836), .C2(n5133), .A(n10991), .B(n9592), .ZN(n9835)
         );
  NAND2_X1 U10574 ( .A1(n9835), .A2(n9593), .ZN(n9597) );
  INV_X1 U10575 ( .A(n9594), .ZN(n9595) );
  AOI22_X1 U10576 ( .A1(n10949), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n9595), 
        .B2(n10938), .ZN(n9596) );
  OAI211_X1 U10577 ( .C1(n9598), .C2(n10705), .A(n9597), .B(n9596), .ZN(n9599)
         );
  AOI21_X1 U10578 ( .B1(n9834), .B2(n10947), .A(n9599), .ZN(n9600) );
  OAI21_X1 U10579 ( .B1(n9838), .B2(n10706), .A(n9600), .ZN(P2_U3271) );
  INV_X1 U10580 ( .A(n9602), .ZN(n9603) );
  AOI21_X1 U10581 ( .B1(n9609), .B2(n9601), .A(n9603), .ZN(n9843) );
  XNOR2_X1 U10582 ( .A(n9607), .B(n9630), .ZN(n9840) );
  INV_X1 U10583 ( .A(n9604), .ZN(n9605) );
  AOI22_X1 U10584 ( .A1(n10949), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n9605), 
        .B2(n10938), .ZN(n9606) );
  OAI21_X1 U10585 ( .B1(n9607), .B2(n10705), .A(n9606), .ZN(n9618) );
  INV_X1 U10586 ( .A(n9608), .ZN(n9612) );
  AOI21_X1 U10587 ( .B1(n9620), .B2(n9610), .A(n9609), .ZN(n9611) );
  NOR3_X1 U10588 ( .A1(n9612), .A2(n9611), .A3(n9717), .ZN(n9616) );
  OAI22_X1 U10589 ( .A1(n9614), .A2(n9720), .B1(n9613), .B2(n9774), .ZN(n9615)
         );
  NOR2_X1 U10590 ( .A1(n9616), .A2(n9615), .ZN(n9842) );
  NOR2_X1 U10591 ( .A1(n9842), .A2(n10949), .ZN(n9617) );
  AOI211_X1 U10592 ( .C1(n9840), .C2(n9763), .A(n9618), .B(n9617), .ZN(n9619)
         );
  OAI21_X1 U10593 ( .B1(n9843), .B2(n10706), .A(n9619), .ZN(P2_U3272) );
  OAI21_X1 U10594 ( .B1(n9621), .B2(n9628), .A(n9620), .ZN(n9623) );
  AOI222_X1 U10595 ( .A1(n10929), .A2(n9623), .B1(n9622), .B2(n10926), .C1(
        n9667), .C2(n10924), .ZN(n9849) );
  OR2_X1 U10596 ( .A1(n9656), .A2(n9624), .ZN(n9627) );
  NAND2_X1 U10597 ( .A1(n9627), .A2(n9625), .ZN(n9845) );
  NAND2_X1 U10598 ( .A1(n9627), .A2(n9626), .ZN(n9629) );
  NAND2_X1 U10599 ( .A1(n9629), .A2(n9628), .ZN(n9844) );
  NAND3_X1 U10600 ( .A1(n9845), .A2(n9844), .A3(n9800), .ZN(n9638) );
  INV_X1 U10601 ( .A(n9642), .ZN(n9632) );
  INV_X1 U10602 ( .A(n9630), .ZN(n9631) );
  AOI21_X1 U10603 ( .B1(n9846), .B2(n9632), .A(n9631), .ZN(n9847) );
  AOI22_X1 U10604 ( .A1(n10949), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n9633), 
        .B2(n10938), .ZN(n9634) );
  OAI21_X1 U10605 ( .B1(n9635), .B2(n10705), .A(n9634), .ZN(n9636) );
  AOI21_X1 U10606 ( .B1(n9847), .B2(n9763), .A(n9636), .ZN(n9637) );
  OAI211_X1 U10607 ( .C1(n10949), .C2(n9849), .A(n9638), .B(n9637), .ZN(
        P2_U3273) );
  OR2_X1 U10608 ( .A1(n9656), .A2(n9664), .ZN(n9654) );
  NAND2_X1 U10609 ( .A1(n9654), .A2(n9639), .ZN(n9641) );
  XNOR2_X1 U10610 ( .A(n9641), .B(n9640), .ZN(n9855) );
  AOI21_X1 U10611 ( .B1(n9851), .B2(n9657), .A(n9642), .ZN(n9852) );
  INV_X1 U10612 ( .A(n9643), .ZN(n9644) );
  AOI22_X1 U10613 ( .A1(n10949), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9644), 
        .B2(n10938), .ZN(n9645) );
  OAI21_X1 U10614 ( .B1(n9646), .B2(n10705), .A(n9645), .ZN(n9652) );
  XNOR2_X1 U10615 ( .A(n9648), .B(n9647), .ZN(n9649) );
  AOI222_X1 U10616 ( .A1(n9673), .A2(n10924), .B1(n9650), .B2(n10926), .C1(
        n10929), .C2(n9649), .ZN(n9854) );
  NOR2_X1 U10617 ( .A1(n9854), .A2(n10949), .ZN(n9651) );
  AOI211_X1 U10618 ( .C1(n9852), .C2(n9763), .A(n9652), .B(n9651), .ZN(n9653)
         );
  OAI21_X1 U10619 ( .B1(n9855), .B2(n10706), .A(n9653), .ZN(P2_U3274) );
  INV_X1 U10620 ( .A(n9654), .ZN(n9655) );
  AOI21_X1 U10621 ( .B1(n9664), .B2(n9656), .A(n9655), .ZN(n9860) );
  INV_X1 U10622 ( .A(n9682), .ZN(n9659) );
  INV_X1 U10623 ( .A(n9657), .ZN(n9658) );
  AOI21_X1 U10624 ( .B1(n9856), .B2(n9659), .A(n9658), .ZN(n9857) );
  INV_X1 U10625 ( .A(n9660), .ZN(n9661) );
  AOI22_X1 U10626 ( .A1(n10949), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9661), 
        .B2(n10938), .ZN(n9662) );
  OAI21_X1 U10627 ( .B1(n9663), .B2(n10705), .A(n9662), .ZN(n9670) );
  XNOR2_X1 U10628 ( .A(n9665), .B(n9664), .ZN(n9666) );
  AOI222_X1 U10629 ( .A1(n9668), .A2(n10924), .B1(n9667), .B2(n10926), .C1(
        n10929), .C2(n9666), .ZN(n9859) );
  NOR2_X1 U10630 ( .A1(n9859), .A2(n10949), .ZN(n9669) );
  AOI211_X1 U10631 ( .C1(n9857), .C2(n9763), .A(n9670), .B(n9669), .ZN(n9671)
         );
  OAI21_X1 U10632 ( .B1(n9860), .B2(n10706), .A(n9671), .ZN(P2_U3275) );
  XNOR2_X1 U10633 ( .A(n9672), .B(n9676), .ZN(n9674) );
  AOI222_X1 U10634 ( .A1(n10929), .A2(n9674), .B1(n9673), .B2(n10926), .C1(
        n5455), .C2(n10924), .ZN(n9864) );
  OAI21_X1 U10635 ( .B1(n9677), .B2(n9676), .A(n9675), .ZN(n9865) );
  OAI22_X1 U10636 ( .A1(n10947), .A2(n9679), .B1(n9678), .B2(n10700), .ZN(
        n9680) );
  AOI21_X1 U10637 ( .B1(n9861), .B2(n9797), .A(n9680), .ZN(n9684) );
  AND2_X1 U10638 ( .A1(n9861), .A2(n5178), .ZN(n9681) );
  NOR2_X1 U10639 ( .A1(n9682), .A2(n9681), .ZN(n9862) );
  NAND2_X1 U10640 ( .A1(n9862), .A2(n9763), .ZN(n9683) );
  OAI211_X1 U10641 ( .C1(n9865), .C2(n10706), .A(n9684), .B(n9683), .ZN(n9685)
         );
  INV_X1 U10642 ( .A(n9685), .ZN(n9686) );
  OAI21_X1 U10643 ( .B1(n10949), .B2(n9864), .A(n9686), .ZN(P2_U3276) );
  OAI21_X1 U10644 ( .B1(n9688), .B2(n9689), .A(n9687), .ZN(n9870) );
  AOI22_X1 U10645 ( .A1(n9868), .A2(n9797), .B1(P2_REG2_REG_19__SCAN_IN), .B2(
        n10949), .ZN(n9699) );
  XNOR2_X1 U10646 ( .A(n9690), .B(n9689), .ZN(n9691) );
  OAI222_X1 U10647 ( .A1(n9720), .A2(n9692), .B1(n9691), .B2(n9717), .C1(n9774), .C2(n9719), .ZN(n9866) );
  INV_X1 U10648 ( .A(n9701), .ZN(n9693) );
  NAND2_X1 U10649 ( .A1(n9693), .A2(n9868), .ZN(n9694) );
  AND3_X1 U10650 ( .A1(n5178), .A2(n9694), .A3(n10930), .ZN(n9867) );
  NAND2_X1 U10651 ( .A1(n9867), .A2(n9742), .ZN(n9695) );
  OAI21_X1 U10652 ( .B1(n10700), .B2(n9696), .A(n9695), .ZN(n9697) );
  OAI21_X1 U10653 ( .B1(n9866), .B2(n9697), .A(n10947), .ZN(n9698) );
  OAI211_X1 U10654 ( .C1(n9870), .C2(n10706), .A(n9699), .B(n9698), .ZN(
        P2_U3277) );
  XNOR2_X1 U10655 ( .A(n9700), .B(n5357), .ZN(n9875) );
  INV_X1 U10656 ( .A(n9714), .ZN(n9702) );
  AOI21_X1 U10657 ( .B1(n9871), .B2(n9702), .A(n9701), .ZN(n9872) );
  INV_X1 U10658 ( .A(n9703), .ZN(n9704) );
  AOI22_X1 U10659 ( .A1(n10949), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9704), 
        .B2(n10938), .ZN(n9705) );
  OAI21_X1 U10660 ( .B1(n9706), .B2(n10705), .A(n9705), .ZN(n9712) );
  XNOR2_X1 U10661 ( .A(n9708), .B(n9707), .ZN(n9710) );
  AOI222_X1 U10662 ( .A1(n10929), .A2(n9710), .B1(n5455), .B2(n10926), .C1(
        n9709), .C2(n10924), .ZN(n9874) );
  NOR2_X1 U10663 ( .A1(n9874), .A2(n10949), .ZN(n9711) );
  AOI211_X1 U10664 ( .C1(n9872), .C2(n9763), .A(n9712), .B(n9711), .ZN(n9713)
         );
  OAI21_X1 U10665 ( .B1(n9875), .B2(n10706), .A(n9713), .ZN(P2_U3278) );
  AOI211_X1 U10666 ( .C1(n9878), .C2(n9733), .A(n10991), .B(n9714), .ZN(n9877)
         );
  XNOR2_X1 U10667 ( .A(n9715), .B(n9722), .ZN(n9716) );
  OAI222_X1 U10668 ( .A1(n9720), .A2(n9719), .B1(n9774), .B2(n9718), .C1(n9717), .C2(n9716), .ZN(n9876) );
  OAI21_X1 U10669 ( .B1(n9723), .B2(n9722), .A(n9721), .ZN(n9729) );
  INV_X1 U10670 ( .A(n9729), .ZN(n9880) );
  NOR2_X1 U10671 ( .A1(n9880), .A2(n9813), .ZN(n9724) );
  AOI211_X1 U10672 ( .C1(n9877), .C2(n9742), .A(n9876), .B(n9724), .ZN(n9732)
         );
  OAI22_X1 U10673 ( .A1(n10947), .A2(n9726), .B1(n9725), .B2(n10700), .ZN(
        n9727) );
  AOI21_X1 U10674 ( .B1(n9878), .B2(n9797), .A(n9727), .ZN(n9731) );
  NAND2_X1 U10675 ( .A1(n9729), .A2(n9728), .ZN(n9730) );
  OAI211_X1 U10676 ( .C1(n9732), .C2(n10949), .A(n9731), .B(n9730), .ZN(
        P2_U3279) );
  INV_X1 U10677 ( .A(n9733), .ZN(n9734) );
  AOI211_X1 U10678 ( .C1(n9883), .C2(n9750), .A(n10991), .B(n9734), .ZN(n9882)
         );
  NOR2_X1 U10679 ( .A1(n10700), .A2(n9735), .ZN(n9741) );
  OAI21_X1 U10680 ( .B1(n9757), .B2(n9748), .A(n9736), .ZN(n9737) );
  XOR2_X1 U10681 ( .A(n9743), .B(n9737), .Z(n9739) );
  AOI21_X1 U10682 ( .B1(n9739), .B2(n10929), .A(n9738), .ZN(n9885) );
  INV_X1 U10683 ( .A(n9885), .ZN(n9740) );
  AOI211_X1 U10684 ( .C1(n9882), .C2(n9742), .A(n9741), .B(n9740), .ZN(n9747)
         );
  AOI22_X1 U10685 ( .A1(n9883), .A2(n9797), .B1(n10949), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n9746) );
  NAND2_X1 U10686 ( .A1(n9744), .A2(n9743), .ZN(n9881) );
  NAND3_X1 U10687 ( .A1(n5672), .A2(n9800), .A3(n9881), .ZN(n9745) );
  OAI211_X1 U10688 ( .C1(n9747), .C2(n10949), .A(n9746), .B(n9745), .ZN(
        P2_U3280) );
  XNOR2_X1 U10689 ( .A(n9749), .B(n9748), .ZN(n9892) );
  INV_X1 U10690 ( .A(n9750), .ZN(n9751) );
  AOI21_X1 U10691 ( .B1(n9888), .B2(n9780), .A(n9751), .ZN(n9889) );
  INV_X1 U10692 ( .A(n9888), .ZN(n9755) );
  INV_X1 U10693 ( .A(n9752), .ZN(n9753) );
  AOI22_X1 U10694 ( .A1(n10949), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n9753), 
        .B2(n10938), .ZN(n9754) );
  OAI21_X1 U10695 ( .B1(n9755), .B2(n10705), .A(n9754), .ZN(n9762) );
  XNOR2_X1 U10696 ( .A(n9757), .B(n9756), .ZN(n9760) );
  AOI222_X1 U10697 ( .A1(n10929), .A2(n9760), .B1(n9759), .B2(n10926), .C1(
        n9758), .C2(n10924), .ZN(n9891) );
  NOR2_X1 U10698 ( .A1(n9891), .A2(n10949), .ZN(n9761) );
  AOI211_X1 U10699 ( .C1(n9889), .C2(n9763), .A(n9762), .B(n9761), .ZN(n9764)
         );
  OAI21_X1 U10700 ( .B1(n9892), .B2(n10706), .A(n9764), .ZN(P2_U3281) );
  AOI21_X1 U10701 ( .B1(n9766), .B2(n9765), .A(n5181), .ZN(n10988) );
  OAI21_X1 U10702 ( .B1(n5165), .B2(n9769), .A(n9768), .ZN(n9770) );
  NAND3_X1 U10703 ( .A1(n5457), .A2(n10929), .A3(n9770), .ZN(n9773) );
  NAND2_X1 U10704 ( .A1(n9771), .A2(n10926), .ZN(n9772) );
  OAI211_X1 U10705 ( .C1(n9775), .C2(n9774), .A(n9773), .B(n9772), .ZN(n10994)
         );
  INV_X1 U10706 ( .A(n10994), .ZN(n9776) );
  OAI21_X1 U10707 ( .B1(n9777), .B2(n10700), .A(n9776), .ZN(n9784) );
  OR2_X1 U10708 ( .A1(n9778), .A2(n10990), .ZN(n9779) );
  NAND2_X1 U10709 ( .A1(n9780), .A2(n9779), .ZN(n10992) );
  AOI22_X1 U10710 ( .A1(n9781), .A2(n9797), .B1(n10949), .B2(
        P2_REG2_REG_14__SCAN_IN), .ZN(n9782) );
  OAI21_X1 U10711 ( .B1(n10992), .B2(n10702), .A(n9782), .ZN(n9783) );
  AOI21_X1 U10712 ( .B1(n9784), .B2(n10947), .A(n9783), .ZN(n9785) );
  OAI21_X1 U10713 ( .B1(n10988), .B2(n10706), .A(n9785), .ZN(P2_U3282) );
  XOR2_X1 U10714 ( .A(n9786), .B(n9798), .Z(n9787) );
  AOI222_X1 U10715 ( .A1(n9789), .A2(n10924), .B1(n9788), .B2(n10926), .C1(
        n10929), .C2(n9787), .ZN(n10816) );
  MUX2_X1 U10716 ( .A(n9790), .B(n10816), .S(n10947), .Z(n9803) );
  AND2_X1 U10717 ( .A1(n9791), .A2(n9796), .ZN(n9793) );
  OR2_X1 U10718 ( .A1(n9793), .A2(n9792), .ZN(n10820) );
  OAI22_X1 U10719 ( .A1(n10820), .A2(n10702), .B1(n9794), .B2(n10700), .ZN(
        n9795) );
  AOI21_X1 U10720 ( .B1(n9797), .B2(n9796), .A(n9795), .ZN(n9802) );
  NAND2_X1 U10721 ( .A1(n9799), .A2(n9798), .ZN(n10817) );
  NAND3_X1 U10722 ( .A1(n10818), .A2(n10817), .A3(n9800), .ZN(n9801) );
  NAND3_X1 U10723 ( .A1(n9803), .A2(n9802), .A3(n9801), .ZN(P2_U3290) );
  AOI21_X1 U10724 ( .B1(n9805), .B2(n10851), .A(n9804), .ZN(n9806) );
  OAI21_X1 U10725 ( .B1(n9807), .B2(n10991), .A(n9806), .ZN(n9893) );
  MUX2_X1 U10726 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9893), .S(n10998), .Z(
        P2_U3551) );
  NAND3_X1 U10727 ( .A1(n9809), .A2(n10930), .A3(n9808), .ZN(n9811) );
  OAI211_X1 U10728 ( .C1(n9812), .C2(n10989), .A(n9811), .B(n9810), .ZN(n9894)
         );
  MUX2_X1 U10729 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9894), .S(n10998), .Z(
        P2_U3550) );
  NAND2_X1 U10730 ( .A1(n9813), .A2(n10729), .ZN(n10995) );
  MUX2_X1 U10731 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9895), .S(n10998), .Z(
        P2_U3549) );
  NAND2_X1 U10732 ( .A1(n9818), .A2(n10995), .ZN(n9823) );
  AOI22_X1 U10733 ( .A1(n9820), .A2(n10930), .B1(n10851), .B2(n9819), .ZN(
        n9821) );
  NAND3_X1 U10734 ( .A1(n9823), .A2(n9822), .A3(n9821), .ZN(n9896) );
  MUX2_X1 U10735 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9896), .S(n10998), .Z(
        P2_U3548) );
  AOI22_X1 U10736 ( .A1(n9825), .A2(n10930), .B1(n10851), .B2(n9824), .ZN(
        n9826) );
  OAI211_X1 U10737 ( .C1(n9828), .C2(n10972), .A(n9827), .B(n9826), .ZN(n9897)
         );
  MUX2_X1 U10738 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9897), .S(n10998), .Z(
        P2_U3547) );
  AOI21_X1 U10739 ( .B1(n10851), .B2(n9830), .A(n9829), .ZN(n9831) );
  OAI211_X1 U10740 ( .C1(n9833), .C2(n10972), .A(n9832), .B(n9831), .ZN(n9898)
         );
  MUX2_X1 U10741 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9898), .S(n10998), .Z(
        P2_U3546) );
  AOI211_X1 U10742 ( .C1(n10851), .C2(n9836), .A(n9835), .B(n9834), .ZN(n9837)
         );
  OAI21_X1 U10743 ( .B1(n9838), .B2(n10972), .A(n9837), .ZN(n9899) );
  MUX2_X1 U10744 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9899), .S(n10998), .Z(
        P2_U3545) );
  AOI22_X1 U10745 ( .A1(n9840), .A2(n10930), .B1(n10851), .B2(n9839), .ZN(
        n9841) );
  OAI211_X1 U10746 ( .C1(n9843), .C2(n10972), .A(n9842), .B(n9841), .ZN(n9900)
         );
  MUX2_X1 U10747 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9900), .S(n10998), .Z(
        P2_U3544) );
  NAND3_X1 U10748 ( .A1(n9845), .A2(n9844), .A3(n10995), .ZN(n9850) );
  AOI22_X1 U10749 ( .A1(n9847), .A2(n10930), .B1(n10851), .B2(n9846), .ZN(
        n9848) );
  NAND3_X1 U10750 ( .A1(n9850), .A2(n9849), .A3(n9848), .ZN(n9901) );
  MUX2_X1 U10751 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9901), .S(n10998), .Z(
        P2_U3543) );
  AOI22_X1 U10752 ( .A1(n9852), .A2(n10930), .B1(n10851), .B2(n9851), .ZN(
        n9853) );
  OAI211_X1 U10753 ( .C1(n9855), .C2(n10972), .A(n9854), .B(n9853), .ZN(n9902)
         );
  MUX2_X1 U10754 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9902), .S(n10998), .Z(
        P2_U3542) );
  AOI22_X1 U10755 ( .A1(n9857), .A2(n10930), .B1(n10851), .B2(n9856), .ZN(
        n9858) );
  OAI211_X1 U10756 ( .C1(n9860), .C2(n10972), .A(n9859), .B(n9858), .ZN(n9903)
         );
  MUX2_X1 U10757 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9903), .S(n10998), .Z(
        P2_U3541) );
  AOI22_X1 U10758 ( .A1(n9862), .A2(n10930), .B1(n10851), .B2(n9861), .ZN(
        n9863) );
  OAI211_X1 U10759 ( .C1(n9865), .C2(n10972), .A(n9864), .B(n9863), .ZN(n9904)
         );
  MUX2_X1 U10760 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9904), .S(n10998), .Z(
        P2_U3540) );
  AOI211_X1 U10761 ( .C1(n10851), .C2(n9868), .A(n9867), .B(n9866), .ZN(n9869)
         );
  OAI21_X1 U10762 ( .B1(n9870), .B2(n10972), .A(n9869), .ZN(n9905) );
  MUX2_X1 U10763 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9905), .S(n10998), .Z(
        P2_U3539) );
  AOI22_X1 U10764 ( .A1(n9872), .A2(n10930), .B1(n10851), .B2(n9871), .ZN(
        n9873) );
  OAI211_X1 U10765 ( .C1(n9875), .C2(n10972), .A(n9874), .B(n9873), .ZN(n9906)
         );
  MUX2_X1 U10766 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9906), .S(n10998), .Z(
        P2_U3538) );
  AOI211_X1 U10767 ( .C1(n10851), .C2(n9878), .A(n9877), .B(n9876), .ZN(n9879)
         );
  OAI21_X1 U10768 ( .B1(n9880), .B2(n10972), .A(n9879), .ZN(n9907) );
  MUX2_X1 U10769 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9907), .S(n10998), .Z(
        P2_U3537) );
  NAND2_X1 U10770 ( .A1(n9881), .A2(n10995), .ZN(n9886) );
  AOI21_X1 U10771 ( .B1(n10851), .B2(n9883), .A(n9882), .ZN(n9884) );
  OAI211_X1 U10772 ( .C1(n9887), .C2(n9886), .A(n9885), .B(n9884), .ZN(n9908)
         );
  MUX2_X1 U10773 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9908), .S(n10998), .Z(
        P2_U3536) );
  AOI22_X1 U10774 ( .A1(n9889), .A2(n10930), .B1(n10851), .B2(n9888), .ZN(
        n9890) );
  OAI211_X1 U10775 ( .C1(n9892), .C2(n10972), .A(n9891), .B(n9890), .ZN(n9909)
         );
  MUX2_X1 U10776 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9909), .S(n10998), .Z(
        P2_U3535) );
  MUX2_X1 U10777 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9893), .S(n11002), .Z(
        P2_U3519) );
  MUX2_X1 U10778 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9894), .S(n11002), .Z(
        P2_U3518) );
  MUX2_X1 U10779 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9895), .S(n11002), .Z(
        P2_U3517) );
  MUX2_X1 U10780 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9896), .S(n11002), .Z(
        P2_U3516) );
  MUX2_X1 U10781 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9897), .S(n11002), .Z(
        P2_U3515) );
  MUX2_X1 U10782 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9898), .S(n11002), .Z(
        P2_U3514) );
  MUX2_X1 U10783 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9899), .S(n11002), .Z(
        P2_U3513) );
  MUX2_X1 U10784 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9900), .S(n11002), .Z(
        P2_U3512) );
  MUX2_X1 U10785 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9901), .S(n11002), .Z(
        P2_U3511) );
  MUX2_X1 U10786 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9902), .S(n11002), .Z(
        P2_U3510) );
  MUX2_X1 U10787 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9903), .S(n11002), .Z(
        P2_U3509) );
  MUX2_X1 U10788 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9904), .S(n11002), .Z(
        P2_U3508) );
  MUX2_X1 U10789 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9905), .S(n11002), .Z(
        P2_U3507) );
  MUX2_X1 U10790 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9906), .S(n11002), .Z(
        P2_U3505) );
  MUX2_X1 U10791 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9907), .S(n11002), .Z(
        P2_U3502) );
  MUX2_X1 U10792 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9908), .S(n11002), .Z(
        P2_U3499) );
  MUX2_X1 U10793 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9909), .S(n11002), .Z(
        P2_U3496) );
  NAND2_X1 U10794 ( .A1(n10539), .A2(n9910), .ZN(n9914) );
  NAND4_X1 U10795 ( .A1(n9911), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .A4(n9912), .ZN(n9913) );
  OAI211_X1 U10796 ( .C1(n9915), .C2(n9923), .A(n9914), .B(n9913), .ZN(
        P2_U3327) );
  INV_X1 U10797 ( .A(n9916), .ZN(n10542) );
  OAI222_X1 U10798 ( .A1(n5076), .A2(n10542), .B1(n9918), .B2(P2_U3152), .C1(
        n9917), .C2(n9923), .ZN(P2_U3329) );
  OAI222_X1 U10799 ( .A1(n5076), .A2(n10545), .B1(n9920), .B2(P2_U3152), .C1(
        n9919), .C2(n9923), .ZN(P2_U3331) );
  INV_X1 U10800 ( .A(n9921), .ZN(n10548) );
  INV_X1 U10801 ( .A(n9922), .ZN(n9925) );
  OAI222_X1 U10802 ( .A1(n5076), .A2(n10548), .B1(P2_U3152), .B2(n9925), .C1(
        n9924), .C2(n9923), .ZN(P2_U3332) );
  MUX2_X1 U10803 ( .A(n9926), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NAND2_X1 U10804 ( .A1(n5099), .A2(n9927), .ZN(n9928) );
  XOR2_X1 U10805 ( .A(n9929), .B(n9928), .Z(n9937) );
  INV_X1 U10806 ( .A(n10406), .ZN(n9931) );
  AOI22_X1 U10807 ( .A1(n10086), .A2(n10399), .B1(n9931), .B2(n9930), .ZN(
        n9933) );
  OAI211_X1 U10808 ( .C1(n9934), .C2(n10066), .A(n9933), .B(n9932), .ZN(n9935)
         );
  AOI21_X1 U10809 ( .B1(n10413), .B2(n10069), .A(n9935), .ZN(n9936) );
  OAI21_X1 U10810 ( .B1(n9937), .B2(n10071), .A(n9936), .ZN(P1_U3213) );
  NAND2_X1 U10811 ( .A1(n9938), .A2(n9940), .ZN(n9942) );
  XNOR2_X1 U10812 ( .A(n9942), .B(n9941), .ZN(n9947) );
  INV_X1 U10813 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9943) );
  OAI22_X1 U10814 ( .A1(n10065), .A2(n9972), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9943), .ZN(n9945) );
  OAI22_X1 U10815 ( .A1(n10066), .A2(n9961), .B1(n10083), .B2(n10254), .ZN(
        n9944) );
  AOI211_X1 U10816 ( .C1(n10479), .C2(n10069), .A(n9945), .B(n9944), .ZN(n9946) );
  OAI21_X1 U10817 ( .B1(n9947), .B2(n10071), .A(n9946), .ZN(P1_U3214) );
  XNOR2_X1 U10818 ( .A(n9949), .B(n9948), .ZN(n9950) );
  XNOR2_X1 U10819 ( .A(n9951), .B(n9950), .ZN(n9955) );
  NAND2_X1 U10820 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n10152)
         );
  OAI21_X1 U10821 ( .B1(n10066), .B2(n10315), .A(n10152), .ZN(n9953) );
  OAI22_X1 U10822 ( .A1(n10065), .A2(n10316), .B1(n10083), .B2(n10320), .ZN(
        n9952) );
  AOI211_X1 U10823 ( .C1(n10503), .C2(n10069), .A(n9953), .B(n9952), .ZN(n9954) );
  OAI21_X1 U10824 ( .B1(n9955), .B2(n10071), .A(n9954), .ZN(P1_U3217) );
  INV_X1 U10825 ( .A(n9956), .ZN(n9957) );
  NOR2_X1 U10826 ( .A1(n9958), .A2(n9957), .ZN(n9959) );
  XNOR2_X1 U10827 ( .A(n5154), .B(n9959), .ZN(n9965) );
  INV_X1 U10828 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9960) );
  OAI22_X1 U10829 ( .A1(n10065), .A2(n9961), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9960), .ZN(n9963) );
  OAI22_X1 U10830 ( .A1(n10066), .A2(n10316), .B1(n10291), .B2(n10083), .ZN(
        n9962) );
  AOI211_X1 U10831 ( .C1(n10490), .C2(n10069), .A(n9963), .B(n9962), .ZN(n9964) );
  OAI21_X1 U10832 ( .B1(n9965), .B2(n10071), .A(n9964), .ZN(P1_U3221) );
  XNOR2_X1 U10833 ( .A(n9968), .B(n9967), .ZN(n9969) );
  XNOR2_X1 U10834 ( .A(n9966), .B(n9969), .ZN(n9976) );
  OAI22_X1 U10835 ( .A1(n10065), .A2(n9971), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9970), .ZN(n9974) );
  OAI22_X1 U10836 ( .A1(n10066), .A2(n9972), .B1(n10083), .B2(n10220), .ZN(
        n9973) );
  AOI211_X1 U10837 ( .C1(n10470), .C2(n10069), .A(n9974), .B(n9973), .ZN(n9975) );
  OAI21_X1 U10838 ( .B1(n9976), .B2(n10071), .A(n9975), .ZN(P1_U3223) );
  INV_X1 U10839 ( .A(n9978), .ZN(n9979) );
  NOR2_X1 U10840 ( .A1(n9977), .A2(n9979), .ZN(n10076) );
  NOR2_X1 U10841 ( .A1(n10076), .A2(n10073), .ZN(n10075) );
  INV_X1 U10842 ( .A(n10075), .ZN(n9980) );
  NAND2_X1 U10843 ( .A1(n9977), .A2(n9979), .ZN(n10074) );
  NAND2_X1 U10844 ( .A1(n9980), .A2(n10074), .ZN(n10077) );
  XNOR2_X1 U10845 ( .A(n9982), .B(n9981), .ZN(n9983) );
  XNOR2_X1 U10846 ( .A(n10077), .B(n9983), .ZN(n9988) );
  INV_X1 U10847 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9984) );
  OAI22_X1 U10848 ( .A1(n10065), .A2(n10371), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9984), .ZN(n9986) );
  OAI22_X1 U10849 ( .A1(n10066), .A2(n10370), .B1(n10374), .B2(n10083), .ZN(
        n9985) );
  AOI211_X1 U10850 ( .C1(n10513), .C2(n10069), .A(n9986), .B(n9985), .ZN(n9987) );
  OAI21_X1 U10851 ( .B1(n9988), .B2(n10071), .A(n9987), .ZN(P1_U3224) );
  XOR2_X1 U10852 ( .A(n9990), .B(n9989), .Z(n9995) );
  INV_X1 U10853 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9991) );
  OAI22_X1 U10854 ( .A1(n10065), .A2(n10315), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9991), .ZN(n9993) );
  OAI22_X1 U10855 ( .A1(n10066), .A2(n10385), .B1(n10350), .B2(n10083), .ZN(
        n9992) );
  AOI211_X1 U10856 ( .C1(n10356), .C2(n10069), .A(n9993), .B(n9992), .ZN(n9994) );
  OAI21_X1 U10857 ( .B1(n9995), .B2(n10071), .A(n9994), .ZN(P1_U3226) );
  XOR2_X1 U10858 ( .A(n9996), .B(n5153), .Z(n10001) );
  OAI22_X1 U10859 ( .A1(n10065), .A2(n10242), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9997), .ZN(n9999) );
  OAI22_X1 U10860 ( .A1(n10066), .A2(n10269), .B1(n10083), .B2(n10245), .ZN(
        n9998) );
  AOI211_X1 U10861 ( .C1(n10476), .C2(n10069), .A(n9999), .B(n9998), .ZN(
        n10000) );
  OAI21_X1 U10862 ( .B1(n10001), .B2(n10071), .A(n10000), .ZN(P1_U3227) );
  AND2_X1 U10863 ( .A1(n10003), .A2(n10002), .ZN(n10005) );
  OAI21_X1 U10864 ( .B1(n10006), .B2(n10005), .A(n10004), .ZN(n10007) );
  NAND2_X1 U10865 ( .A1(n10007), .A2(n10078), .ZN(n10012) );
  OAI22_X1 U10866 ( .A1(n10065), .A2(n10890), .B1(n10083), .B2(n10008), .ZN(
        n10009) );
  AOI211_X1 U10867 ( .C1(n10081), .C2(n10098), .A(n10010), .B(n10009), .ZN(
        n10011) );
  OAI211_X1 U10868 ( .C1(n5390), .C2(n10089), .A(n10012), .B(n10011), .ZN(
        P1_U3229) );
  INV_X1 U10869 ( .A(n10013), .ZN(n10015) );
  NAND2_X1 U10870 ( .A1(n10015), .A2(n10014), .ZN(n10016) );
  XNOR2_X1 U10871 ( .A(n10017), .B(n10016), .ZN(n10022) );
  INV_X1 U10872 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n10018) );
  OAI22_X1 U10873 ( .A1(n10066), .A2(n10297), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10018), .ZN(n10020) );
  OAI22_X1 U10874 ( .A1(n10065), .A2(n10298), .B1(n10083), .B2(n10303), .ZN(
        n10019) );
  AOI211_X1 U10875 ( .C1(n10306), .C2(n10069), .A(n10020), .B(n10019), .ZN(
        n10021) );
  OAI21_X1 U10876 ( .B1(n10022), .B2(n10071), .A(n10021), .ZN(P1_U3231) );
  INV_X1 U10877 ( .A(n10433), .ZN(n10965) );
  INV_X1 U10878 ( .A(n10023), .ZN(n10027) );
  OAI21_X1 U10879 ( .B1(n10027), .B2(n10025), .A(n10024), .ZN(n10026) );
  OAI21_X1 U10880 ( .B1(n5709), .B2(n10027), .A(n10026), .ZN(n10028) );
  NAND2_X1 U10881 ( .A1(n10028), .A2(n10078), .ZN(n10033) );
  NAND2_X1 U10882 ( .A1(n10081), .A2(n10094), .ZN(n10029) );
  OAI21_X1 U10883 ( .B1(n10083), .B2(n10430), .A(n10029), .ZN(n10030) );
  AOI211_X1 U10884 ( .C1(n10086), .C2(n10093), .A(n10031), .B(n10030), .ZN(
        n10032) );
  OAI211_X1 U10885 ( .C1(n10965), .C2(n10089), .A(n10033), .B(n10032), .ZN(
        P1_U3232) );
  INV_X1 U10886 ( .A(n10034), .ZN(n10036) );
  NAND2_X1 U10887 ( .A1(n10036), .A2(n10035), .ZN(n10037) );
  XNOR2_X1 U10888 ( .A(n10038), .B(n10037), .ZN(n10043) );
  INV_X1 U10889 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n10039) );
  OAI22_X1 U10890 ( .A1(n10065), .A2(n10269), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10039), .ZN(n10041) );
  OAI22_X1 U10891 ( .A1(n10066), .A2(n10298), .B1(n10083), .B2(n10271), .ZN(
        n10040) );
  AOI211_X1 U10892 ( .C1(n10486), .C2(n10069), .A(n10041), .B(n10040), .ZN(
        n10042) );
  OAI21_X1 U10893 ( .B1(n10043), .B2(n10071), .A(n10042), .ZN(P1_U3233) );
  OAI21_X1 U10894 ( .B1(n10046), .B2(n10045), .A(n10044), .ZN(n10047) );
  NAND2_X1 U10895 ( .A1(n10047), .A2(n10078), .ZN(n10051) );
  AOI22_X1 U10896 ( .A1(n10069), .A2(n10720), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n10048), .ZN(n10050) );
  AOI22_X1 U10897 ( .A1(n10086), .A2(n10103), .B1(n10081), .B2(n6735), .ZN(
        n10049) );
  NAND3_X1 U10898 ( .A1(n10051), .A2(n10050), .A3(n10049), .ZN(P1_U3235) );
  XNOR2_X1 U10899 ( .A(n10053), .B(n10052), .ZN(n10054) );
  XNOR2_X1 U10900 ( .A(n10055), .B(n10054), .ZN(n10061) );
  INV_X1 U10901 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n10056) );
  OAI22_X1 U10902 ( .A1(n10066), .A2(n10371), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10056), .ZN(n10059) );
  INV_X1 U10903 ( .A(n10337), .ZN(n10057) );
  OAI22_X1 U10904 ( .A1(n10065), .A2(n10297), .B1(n10083), .B2(n10057), .ZN(
        n10058) );
  AOI211_X1 U10905 ( .C1(n10506), .C2(n10069), .A(n10059), .B(n10058), .ZN(
        n10060) );
  OAI21_X1 U10906 ( .B1(n10061), .B2(n10071), .A(n10060), .ZN(P1_U3236) );
  XNOR2_X1 U10907 ( .A(n10063), .B(n10062), .ZN(n10072) );
  OAI22_X1 U10908 ( .A1(n10065), .A2(n10206), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10064), .ZN(n10068) );
  OAI22_X1 U10909 ( .A1(n10066), .A2(n10242), .B1(n10083), .B2(n10211), .ZN(
        n10067) );
  AOI211_X1 U10910 ( .C1(n10464), .C2(n10069), .A(n10068), .B(n10067), .ZN(
        n10070) );
  OAI21_X1 U10911 ( .B1(n10072), .B2(n10071), .A(n10070), .ZN(P1_U3238) );
  AOI21_X1 U10912 ( .B1(n10075), .B2(n10074), .A(n10073), .ZN(n10080) );
  NOR2_X1 U10913 ( .A1(n10077), .A2(n10076), .ZN(n10079) );
  OAI21_X1 U10914 ( .B1(n10080), .B2(n10079), .A(n10078), .ZN(n10088) );
  NAND2_X1 U10915 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10109)
         );
  INV_X1 U10916 ( .A(n10109), .ZN(n10085) );
  NAND2_X1 U10917 ( .A1(n10081), .A2(n10093), .ZN(n10082) );
  OAI21_X1 U10918 ( .B1(n10083), .B2(n10389), .A(n10082), .ZN(n10084) );
  AOI211_X1 U10919 ( .C1(n10086), .C2(n10349), .A(n10085), .B(n10084), .ZN(
        n10087) );
  OAI211_X1 U10920 ( .C1(n11004), .C2(n10089), .A(n10088), .B(n10087), .ZN(
        P1_U3239) );
  MUX2_X1 U10921 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n10090), .S(n10104), .Z(
        P1_U3585) );
  MUX2_X1 U10922 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n10173), .S(n10104), .Z(
        P1_U3584) );
  MUX2_X1 U10923 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n10197), .S(n10104), .Z(
        P1_U3583) );
  MUX2_X1 U10924 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n10174), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10925 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n10228), .S(n10104), .Z(
        P1_U3581) );
  MUX2_X1 U10926 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n10091), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10927 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n10260), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10928 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n10284), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10929 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n10092), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10930 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n10283), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10931 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n10331), .S(n10104), .Z(
        P1_U3574) );
  MUX2_X1 U10932 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n10348), .S(n10104), .Z(
        P1_U3573) );
  MUX2_X1 U10933 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n10332), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10934 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n10349), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10935 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n10399), .S(n10104), .Z(
        P1_U3570) );
  MUX2_X1 U10936 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n10093), .S(n10104), .Z(
        P1_U3569) );
  MUX2_X1 U10937 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n10404), .S(n10104), .Z(
        P1_U3568) );
  MUX2_X1 U10938 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n10094), .S(n10104), .Z(
        P1_U3567) );
  MUX2_X1 U10939 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n10095), .S(n10104), .Z(
        P1_U3566) );
  MUX2_X1 U10940 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n10096), .S(n10104), .Z(
        P1_U3565) );
  MUX2_X1 U10941 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n10097), .S(n10104), .Z(
        P1_U3564) );
  MUX2_X1 U10942 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n10098), .S(n10104), .Z(
        P1_U3563) );
  MUX2_X1 U10943 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n10099), .S(n10104), .Z(
        P1_U3562) );
  MUX2_X1 U10944 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n10100), .S(n10104), .Z(
        P1_U3561) );
  MUX2_X1 U10945 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n10101), .S(n10104), .Z(
        P1_U3560) );
  MUX2_X1 U10946 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n10102), .S(n10104), .Z(
        P1_U3559) );
  MUX2_X1 U10947 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n10103), .S(n10104), .Z(
        P1_U3558) );
  MUX2_X1 U10948 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n7642), .S(n10104), .Z(
        P1_U3557) );
  MUX2_X1 U10949 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6735), .S(n10104), .Z(
        P1_U3556) );
  MUX2_X1 U10950 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n7643), .S(n10104), .Z(
        P1_U3555) );
  AOI211_X1 U10951 ( .C1(n10106), .C2(n10390), .A(n10105), .B(n10627), .ZN(
        n10114) );
  AOI211_X1 U10952 ( .C1(n10108), .C2(n6690), .A(n10107), .B(n10118), .ZN(
        n10113) );
  NAND2_X1 U10953 ( .A1(n10670), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n10110) );
  OAI211_X1 U10954 ( .C1(n10659), .C2(n10111), .A(n10110), .B(n10109), .ZN(
        n10112) );
  OR3_X1 U10955 ( .A1(n10114), .A2(n10113), .A3(n10112), .ZN(P1_U3256) );
  AOI211_X1 U10956 ( .C1(n10117), .C2(n10116), .A(n10115), .B(n10627), .ZN(
        n10127) );
  AOI211_X1 U10957 ( .C1(n10121), .C2(n10120), .A(n10119), .B(n10118), .ZN(
        n10126) );
  NAND2_X1 U10958 ( .A1(n10670), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n10123) );
  NAND2_X1 U10959 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n10122)
         );
  OAI211_X1 U10960 ( .C1(n10659), .C2(n10124), .A(n10123), .B(n10122), .ZN(
        n10125) );
  OR3_X1 U10961 ( .A1(n10127), .A2(n10126), .A3(n10125), .ZN(P1_U3257) );
  AND2_X1 U10962 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3084), .ZN(n10133) );
  AOI21_X1 U10963 ( .B1(n10136), .B2(P1_REG2_REG_17__SCAN_IN), .A(n10128), 
        .ZN(n10131) );
  NAND2_X1 U10964 ( .A1(n10146), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n10129) );
  OAI21_X1 U10965 ( .B1(n10146), .B2(P1_REG2_REG_18__SCAN_IN), .A(n10129), 
        .ZN(n10130) );
  NOR2_X1 U10966 ( .A1(n10131), .A2(n10130), .ZN(n10142) );
  AOI211_X1 U10967 ( .C1(n10131), .C2(n10130), .A(n10142), .B(n10627), .ZN(
        n10132) );
  AOI211_X1 U10968 ( .C1(n10670), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n10133), 
        .B(n10132), .ZN(n10141) );
  XNOR2_X1 U10969 ( .A(n10146), .B(n10134), .ZN(n10138) );
  AOI21_X1 U10970 ( .B1(n10136), .B2(P1_REG1_REG_17__SCAN_IN), .A(n10135), 
        .ZN(n10137) );
  NAND2_X1 U10971 ( .A1(n10137), .A2(n10138), .ZN(n10145) );
  OAI21_X1 U10972 ( .B1(n10138), .B2(n10137), .A(n10145), .ZN(n10139) );
  AOI22_X1 U10973 ( .A1(n10146), .A2(n10151), .B1(n10662), .B2(n10139), .ZN(
        n10140) );
  NAND2_X1 U10974 ( .A1(n10141), .A2(n10140), .ZN(P1_U3259) );
  MUX2_X1 U10975 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n10321), .S(n5073), .Z(
        n10144) );
  AOI21_X1 U10976 ( .B1(n10146), .B2(P1_REG2_REG_18__SCAN_IN), .A(n10142), 
        .ZN(n10143) );
  XOR2_X1 U10977 ( .A(n10144), .B(n10143), .Z(n10156) );
  OAI21_X1 U10978 ( .B1(n10146), .B2(P1_REG1_REG_18__SCAN_IN), .A(n10145), 
        .ZN(n10149) );
  XNOR2_X1 U10979 ( .A(n5073), .B(n10147), .ZN(n10148) );
  XNOR2_X1 U10980 ( .A(n10149), .B(n10148), .ZN(n10150) );
  AOI22_X1 U10981 ( .A1(n5073), .A2(n10151), .B1(n10662), .B2(n10150), .ZN(
        n10155) );
  INV_X1 U10982 ( .A(n10152), .ZN(n10153) );
  AOI21_X1 U10983 ( .B1(n10670), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n10153), 
        .ZN(n10154) );
  OAI211_X1 U10984 ( .C1(n10156), .C2(n10627), .A(n10155), .B(n10154), .ZN(
        P1_U3260) );
  NAND2_X1 U10985 ( .A1(n10163), .A2(n10162), .ZN(n10157) );
  XNOR2_X1 U10986 ( .A(n10443), .B(n10157), .ZN(n10441) );
  NAND2_X1 U10987 ( .A1(n10441), .A2(n10902), .ZN(n10161) );
  NAND2_X1 U10988 ( .A1(n10159), .A2(n10158), .ZN(n10446) );
  NOR2_X1 U10989 ( .A1(n10439), .A2(n10446), .ZN(n10165) );
  AOI21_X1 U10990 ( .B1(n10439), .B2(P1_REG2_REG_31__SCAN_IN), .A(n10165), 
        .ZN(n10160) );
  OAI211_X1 U10991 ( .C1(n10443), .C2(n10905), .A(n10161), .B(n10160), .ZN(
        P1_U3261) );
  XNOR2_X1 U10992 ( .A(n10163), .B(n10162), .ZN(n10447) );
  NOR2_X1 U10993 ( .A1(n5074), .A2(n10164), .ZN(n10166) );
  AOI211_X1 U10994 ( .C1(n10444), .C2(n10432), .A(n10166), .B(n10165), .ZN(
        n10167) );
  OAI21_X1 U10995 ( .B1(n10447), .B2(n10435), .A(n10167), .ZN(P1_U3262) );
  NAND2_X1 U10996 ( .A1(n5149), .A2(n10171), .ZN(n10169) );
  OAI211_X1 U10997 ( .C1(n10172), .C2(n10171), .A(n10170), .B(n10892), .ZN(
        n10176) );
  AOI22_X1 U10998 ( .A1(n10405), .A2(n10174), .B1(n10173), .B2(n10398), .ZN(
        n10175) );
  OAI22_X1 U10999 ( .A1(n5074), .A2(n10179), .B1(n10178), .B2(n10907), .ZN(
        n10180) );
  AOI21_X1 U11000 ( .B1(n10454), .B2(n10432), .A(n10180), .ZN(n10185) );
  INV_X1 U11001 ( .A(n10190), .ZN(n10181) );
  NAND2_X1 U11002 ( .A1(n10454), .A2(n10181), .ZN(n10182) );
  NAND2_X1 U11003 ( .A1(n10455), .A2(n10902), .ZN(n10184) );
  OAI211_X1 U11004 ( .C1(n10458), .C2(n10751), .A(n10185), .B(n10184), .ZN(
        n10186) );
  AOI21_X1 U11005 ( .B1(n10453), .B2(n5074), .A(n10186), .ZN(n10187) );
  INV_X1 U11006 ( .A(n10187), .ZN(P1_U3263) );
  XNOR2_X1 U11007 ( .A(n10189), .B(n10188), .ZN(n10463) );
  AOI21_X1 U11008 ( .B1(n10459), .B2(n10209), .A(n10190), .ZN(n10460) );
  AOI22_X1 U11009 ( .A1(n10439), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n10191), 
        .B2(n10790), .ZN(n10192) );
  OAI21_X1 U11010 ( .B1(n10193), .B2(n10905), .A(n10192), .ZN(n10201) );
  OAI211_X1 U11011 ( .C1(n10196), .C2(n10195), .A(n10194), .B(n10892), .ZN(
        n10199) );
  AOI22_X1 U11012 ( .A1(n10405), .A2(n10228), .B1(n10197), .B2(n10398), .ZN(
        n10198) );
  NOR2_X1 U11013 ( .A1(n10462), .A2(n10439), .ZN(n10200) );
  AOI211_X1 U11014 ( .C1(n10460), .C2(n10902), .A(n10201), .B(n10200), .ZN(
        n10202) );
  OAI21_X1 U11015 ( .B1(n10381), .B2(n10463), .A(n10202), .ZN(P1_U3264) );
  XNOR2_X1 U11016 ( .A(n10203), .B(n10205), .ZN(n10208) );
  OAI22_X1 U11017 ( .A1(n10206), .A2(n10887), .B1(n10242), .B2(n10889), .ZN(
        n10207) );
  INV_X1 U11018 ( .A(n10209), .ZN(n10210) );
  AOI21_X1 U11019 ( .B1(n10464), .B2(n10219), .A(n10210), .ZN(n10465) );
  INV_X1 U11020 ( .A(n10211), .ZN(n10212) );
  AOI22_X1 U11021 ( .A1(n10439), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n10212), 
        .B2(n10790), .ZN(n10213) );
  OAI21_X1 U11022 ( .B1(n5402), .B2(n10905), .A(n10213), .ZN(n10215) );
  NOR2_X1 U11023 ( .A1(n10468), .A2(n10751), .ZN(n10214) );
  AOI211_X1 U11024 ( .C1(n10465), .C2(n10902), .A(n10215), .B(n10214), .ZN(
        n10216) );
  OAI21_X1 U11025 ( .B1(n10467), .B2(n10439), .A(n10216), .ZN(P1_U3265) );
  XNOR2_X1 U11026 ( .A(n10218), .B(n10217), .ZN(n10473) );
  AOI211_X1 U11027 ( .C1(n10470), .C2(n10243), .A(n11005), .B(n5403), .ZN(
        n10469) );
  INV_X1 U11028 ( .A(n10470), .ZN(n10223) );
  INV_X1 U11029 ( .A(n10220), .ZN(n10221) );
  AOI22_X1 U11030 ( .A1(n10439), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n10221), 
        .B2(n10790), .ZN(n10222) );
  OAI21_X1 U11031 ( .B1(n10223), .B2(n10905), .A(n10222), .ZN(n10231) );
  NAND2_X1 U11032 ( .A1(n10225), .A2(n10224), .ZN(n10227) );
  OAI21_X1 U11033 ( .B1(n5163), .B2(n10227), .A(n10226), .ZN(n10229) );
  AOI222_X1 U11034 ( .A1(n10892), .A2(n10229), .B1(n10228), .B2(n10398), .C1(
        n10260), .C2(n10405), .ZN(n10472) );
  NOR2_X1 U11035 ( .A1(n10472), .A2(n10439), .ZN(n10230) );
  AOI211_X1 U11036 ( .C1(n10469), .C2(n10373), .A(n10231), .B(n10230), .ZN(
        n10232) );
  OAI21_X1 U11037 ( .B1(n10473), .B2(n10381), .A(n10232), .ZN(P1_U3266) );
  NAND2_X1 U11038 ( .A1(n10234), .A2(n10233), .ZN(n10235) );
  XOR2_X1 U11039 ( .A(n10240), .B(n10235), .Z(n10478) );
  INV_X1 U11040 ( .A(n10236), .ZN(n10237) );
  NOR2_X1 U11041 ( .A1(n10238), .A2(n10237), .ZN(n10239) );
  XOR2_X1 U11042 ( .A(n10240), .B(n10239), .Z(n10241) );
  OAI222_X1 U11043 ( .A1(n10887), .A2(n10242), .B1(n10241), .B2(n10784), .C1(
        n10889), .C2(n10269), .ZN(n10474) );
  INV_X1 U11044 ( .A(n10243), .ZN(n10244) );
  AOI211_X1 U11045 ( .C1(n10476), .C2(n10252), .A(n11005), .B(n10244), .ZN(
        n10475) );
  INV_X1 U11046 ( .A(n10475), .ZN(n10246) );
  OAI22_X1 U11047 ( .A1(n10246), .A2(n5073), .B1(n10907), .B2(n10245), .ZN(
        n10247) );
  OAI21_X1 U11048 ( .B1(n10474), .B2(n10247), .A(n5074), .ZN(n10249) );
  AOI22_X1 U11049 ( .A1(n10476), .A2(n10432), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10439), .ZN(n10248) );
  OAI211_X1 U11050 ( .C1(n10478), .C2(n10381), .A(n10249), .B(n10248), .ZN(
        P1_U3267) );
  XNOR2_X1 U11051 ( .A(n10251), .B(n10250), .ZN(n10483) );
  INV_X1 U11052 ( .A(n10252), .ZN(n10253) );
  AOI21_X1 U11053 ( .B1(n10479), .B2(n5395), .A(n10253), .ZN(n10480) );
  INV_X1 U11054 ( .A(n10254), .ZN(n10255) );
  AOI22_X1 U11055 ( .A1(n10439), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n10255), 
        .B2(n10790), .ZN(n10256) );
  OAI21_X1 U11056 ( .B1(n10257), .B2(n10905), .A(n10256), .ZN(n10263) );
  XNOR2_X1 U11057 ( .A(n10259), .B(n10258), .ZN(n10261) );
  AOI222_X1 U11058 ( .A1(n10892), .A2(n10261), .B1(n10260), .B2(n10398), .C1(
        n10284), .C2(n10405), .ZN(n10482) );
  NOR2_X1 U11059 ( .A1(n10482), .A2(n10439), .ZN(n10262) );
  AOI211_X1 U11060 ( .C1(n10480), .C2(n10902), .A(n10263), .B(n10262), .ZN(
        n10264) );
  OAI21_X1 U11061 ( .B1(n10381), .B2(n10483), .A(n10264), .ZN(P1_U3268) );
  XOR2_X1 U11062 ( .A(n10265), .B(n10266), .Z(n10488) );
  XNOR2_X1 U11063 ( .A(n10267), .B(n10266), .ZN(n10268) );
  OAI222_X1 U11064 ( .A1(n10887), .A2(n10269), .B1(n10889), .B2(n10298), .C1(
        n10784), .C2(n10268), .ZN(n10484) );
  NAND2_X1 U11065 ( .A1(n10484), .A2(n5074), .ZN(n10276) );
  AOI211_X1 U11066 ( .C1(n10486), .C2(n10288), .A(n11005), .B(n10270), .ZN(
        n10485) );
  NOR2_X1 U11067 ( .A1(n5394), .A2(n10905), .ZN(n10274) );
  OAI22_X1 U11068 ( .A1(n5074), .A2(n10272), .B1(n10271), .B2(n10907), .ZN(
        n10273) );
  AOI211_X1 U11069 ( .C1(n10485), .C2(n10373), .A(n10274), .B(n10273), .ZN(
        n10275) );
  OAI211_X1 U11070 ( .C1(n10488), .C2(n10381), .A(n10276), .B(n10275), .ZN(
        P1_U3269) );
  OAI21_X1 U11071 ( .B1(n10278), .B2(n10281), .A(n10277), .ZN(n10493) );
  NAND2_X1 U11072 ( .A1(n10280), .A2(n10279), .ZN(n10282) );
  XNOR2_X1 U11073 ( .A(n10282), .B(n10281), .ZN(n10285) );
  AOI222_X1 U11074 ( .A1(n10892), .A2(n10285), .B1(n10284), .B2(n10398), .C1(
        n10283), .C2(n10405), .ZN(n10492) );
  OR2_X1 U11075 ( .A1(n10300), .A2(n10286), .ZN(n10287) );
  AND3_X1 U11076 ( .A1(n10288), .A2(n10287), .A3(n10778), .ZN(n10489) );
  NAND2_X1 U11077 ( .A1(n10489), .A2(n10289), .ZN(n10290) );
  OAI211_X1 U11078 ( .C1(n10291), .C2(n10907), .A(n10492), .B(n10290), .ZN(
        n10292) );
  NAND2_X1 U11079 ( .A1(n10292), .A2(n5074), .ZN(n10294) );
  AOI22_X1 U11080 ( .A1(n10490), .A2(n10432), .B1(n10439), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n10293) );
  OAI211_X1 U11081 ( .C1(n10493), .C2(n10381), .A(n10294), .B(n10293), .ZN(
        P1_U3270) );
  XNOR2_X1 U11082 ( .A(n10295), .B(n10301), .ZN(n10296) );
  OAI222_X1 U11083 ( .A1(n10887), .A2(n10298), .B1(n10889), .B2(n10297), .C1(
        n10784), .C2(n10296), .ZN(n10500) );
  NOR2_X1 U11084 ( .A1(n10317), .A2(n10496), .ZN(n10299) );
  OR2_X1 U11085 ( .A1(n10300), .A2(n10299), .ZN(n10497) );
  NAND2_X1 U11086 ( .A1(n10302), .A2(n10301), .ZN(n10494) );
  NAND3_X1 U11087 ( .A1(n10495), .A2(n10494), .A3(n10437), .ZN(n10308) );
  OAI22_X1 U11088 ( .A1(n5074), .A2(n10304), .B1(n10303), .B2(n10907), .ZN(
        n10305) );
  AOI21_X1 U11089 ( .B1(n10306), .B2(n10432), .A(n10305), .ZN(n10307) );
  OAI211_X1 U11090 ( .C1(n10497), .C2(n10435), .A(n10308), .B(n10307), .ZN(
        n10309) );
  AOI21_X1 U11091 ( .B1(n10500), .B2(n5074), .A(n10309), .ZN(n10310) );
  INV_X1 U11092 ( .A(n10310), .ZN(P1_U3271) );
  XNOR2_X1 U11093 ( .A(n10311), .B(n10313), .ZN(n10505) );
  AOI21_X1 U11094 ( .B1(n5131), .B2(n10313), .A(n10312), .ZN(n10314) );
  OAI222_X1 U11095 ( .A1(n10887), .A2(n10316), .B1(n10889), .B2(n10315), .C1(
        n10784), .C2(n10314), .ZN(n10501) );
  NAND2_X1 U11096 ( .A1(n10501), .A2(n5074), .ZN(n10325) );
  INV_X1 U11097 ( .A(n10336), .ZN(n10318) );
  AOI211_X1 U11098 ( .C1(n10503), .C2(n10318), .A(n11005), .B(n10317), .ZN(
        n10502) );
  NOR2_X1 U11099 ( .A1(n10319), .A2(n10905), .ZN(n10323) );
  OAI22_X1 U11100 ( .A1(n5074), .A2(n10321), .B1(n10320), .B2(n10907), .ZN(
        n10322) );
  AOI211_X1 U11101 ( .C1(n10502), .C2(n10373), .A(n10323), .B(n10322), .ZN(
        n10324) );
  OAI211_X1 U11102 ( .C1(n10505), .C2(n10381), .A(n10325), .B(n10324), .ZN(
        P1_U3272) );
  XNOR2_X1 U11103 ( .A(n10327), .B(n10326), .ZN(n10340) );
  AOI21_X1 U11104 ( .B1(n10330), .B2(n10329), .A(n10328), .ZN(n10334) );
  AOI22_X1 U11105 ( .A1(n10405), .A2(n10332), .B1(n10331), .B2(n10398), .ZN(
        n10333) );
  OAI21_X1 U11106 ( .B1(n10334), .B2(n10784), .A(n10333), .ZN(n10335) );
  AOI21_X1 U11107 ( .B1(n10745), .B2(n10340), .A(n10335), .ZN(n10509) );
  AOI21_X1 U11108 ( .B1(n10506), .B2(n10353), .A(n10336), .ZN(n10507) );
  INV_X1 U11109 ( .A(n10506), .ZN(n10339) );
  AOI22_X1 U11110 ( .A1(n10439), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n10337), 
        .B2(n10790), .ZN(n10338) );
  OAI21_X1 U11111 ( .B1(n10339), .B2(n10905), .A(n10338), .ZN(n10342) );
  INV_X1 U11112 ( .A(n10340), .ZN(n10510) );
  NOR2_X1 U11113 ( .A1(n10510), .A2(n10751), .ZN(n10341) );
  AOI211_X1 U11114 ( .C1(n10507), .C2(n10902), .A(n10342), .B(n10341), .ZN(
        n10343) );
  OAI21_X1 U11115 ( .B1(n10509), .B2(n10439), .A(n10343), .ZN(P1_U3273) );
  INV_X1 U11116 ( .A(n10344), .ZN(n10345) );
  NOR2_X1 U11117 ( .A1(n10366), .A2(n10345), .ZN(n10346) );
  XOR2_X1 U11118 ( .A(n10357), .B(n10346), .Z(n10347) );
  AOI222_X1 U11119 ( .A1(n10349), .A2(n10405), .B1(n10348), .B2(n10398), .C1(
        n10892), .C2(n10347), .ZN(n11014) );
  OAI22_X1 U11120 ( .A1(n5074), .A2(n10351), .B1(n10350), .B2(n10907), .ZN(
        n10355) );
  INV_X1 U11121 ( .A(n10352), .ZN(n10372) );
  INV_X1 U11122 ( .A(n10356), .ZN(n11016) );
  OAI211_X1 U11123 ( .C1(n10372), .C2(n11016), .A(n10778), .B(n10353), .ZN(
        n11013) );
  NOR2_X1 U11124 ( .A1(n11013), .A2(n10410), .ZN(n10354) );
  AOI211_X1 U11125 ( .C1(n10432), .C2(n10356), .A(n10355), .B(n10354), .ZN(
        n10360) );
  XNOR2_X1 U11126 ( .A(n10358), .B(n10357), .ZN(n11019) );
  NAND2_X1 U11127 ( .A1(n11019), .A2(n10437), .ZN(n10359) );
  OAI211_X1 U11128 ( .C1(n11014), .C2(n10439), .A(n10360), .B(n10359), .ZN(
        P1_U3274) );
  XNOR2_X1 U11129 ( .A(n10362), .B(n10361), .ZN(n10515) );
  INV_X1 U11130 ( .A(n10363), .ZN(n10364) );
  NOR2_X1 U11131 ( .A1(n10365), .A2(n10364), .ZN(n10368) );
  AOI21_X1 U11132 ( .B1(n10368), .B2(n10367), .A(n10366), .ZN(n10369) );
  OAI222_X1 U11133 ( .A1(n10887), .A2(n10371), .B1(n10889), .B2(n10370), .C1(
        n10784), .C2(n10369), .ZN(n10511) );
  INV_X1 U11134 ( .A(n10513), .ZN(n10378) );
  AOI211_X1 U11135 ( .C1(n10513), .C2(n10392), .A(n11005), .B(n10372), .ZN(
        n10512) );
  NAND2_X1 U11136 ( .A1(n10512), .A2(n10373), .ZN(n10377) );
  NOR2_X1 U11137 ( .A1(n10907), .A2(n10374), .ZN(n10375) );
  AOI21_X1 U11138 ( .B1(n10439), .B2(P1_REG2_REG_16__SCAN_IN), .A(n10375), 
        .ZN(n10376) );
  OAI211_X1 U11139 ( .C1(n10378), .C2(n10905), .A(n10377), .B(n10376), .ZN(
        n10379) );
  AOI21_X1 U11140 ( .B1(n10511), .B2(n5074), .A(n10379), .ZN(n10380) );
  OAI21_X1 U11141 ( .B1(n10381), .B2(n10515), .A(n10380), .ZN(P1_U3275) );
  XNOR2_X1 U11142 ( .A(n10382), .B(n10384), .ZN(n11003) );
  XOR2_X1 U11143 ( .A(n10384), .B(n10383), .Z(n10387) );
  OAI22_X1 U11144 ( .A1(n10385), .A2(n10887), .B1(n10425), .B2(n10889), .ZN(
        n10386) );
  AOI21_X1 U11145 ( .B1(n10387), .B2(n10892), .A(n10386), .ZN(n10388) );
  OAI21_X1 U11146 ( .B1(n10895), .B2(n11003), .A(n10388), .ZN(n11007) );
  NAND2_X1 U11147 ( .A1(n11007), .A2(n5074), .ZN(n10397) );
  OAI22_X1 U11148 ( .A1(n5074), .A2(n10390), .B1(n10389), .B2(n10907), .ZN(
        n10394) );
  OR2_X1 U11149 ( .A1(n10408), .A2(n11004), .ZN(n10391) );
  NAND2_X1 U11150 ( .A1(n10392), .A2(n10391), .ZN(n11006) );
  NOR2_X1 U11151 ( .A1(n11006), .A2(n10435), .ZN(n10393) );
  AOI211_X1 U11152 ( .C1(n10432), .C2(n10395), .A(n10394), .B(n10393), .ZN(
        n10396) );
  OAI211_X1 U11153 ( .C1(n11003), .C2(n10751), .A(n10397), .B(n10396), .ZN(
        P1_U3276) );
  AND2_X1 U11154 ( .A1(n10399), .A2(n10398), .ZN(n10403) );
  AOI211_X1 U11155 ( .C1(n10414), .C2(n10401), .A(n10784), .B(n10400), .ZN(
        n10402) );
  AOI211_X1 U11156 ( .C1(n10405), .C2(n10404), .A(n10403), .B(n10402), .ZN(
        n10982) );
  OAI22_X1 U11157 ( .A1(n5074), .A2(n10407), .B1(n10406), .B2(n10907), .ZN(
        n10412) );
  INV_X1 U11158 ( .A(n10408), .ZN(n10409) );
  OAI211_X1 U11159 ( .C1(n10983), .C2(n10428), .A(n10409), .B(n10778), .ZN(
        n10981) );
  NOR2_X1 U11160 ( .A1(n10981), .A2(n10410), .ZN(n10411) );
  AOI211_X1 U11161 ( .C1(n10432), .C2(n10413), .A(n10412), .B(n10411), .ZN(
        n10417) );
  XNOR2_X1 U11162 ( .A(n10415), .B(n10414), .ZN(n10985) );
  NAND2_X1 U11163 ( .A1(n10985), .A2(n10437), .ZN(n10416) );
  OAI211_X1 U11164 ( .C1(n10982), .C2(n10439), .A(n10417), .B(n10416), .ZN(
        P1_U3277) );
  INV_X1 U11165 ( .A(n10418), .ZN(n10423) );
  NOR3_X1 U11166 ( .A1(n10421), .A2(n10420), .A3(n10419), .ZN(n10422) );
  NOR2_X1 U11167 ( .A1(n10423), .A2(n10422), .ZN(n10424) );
  OAI222_X1 U11168 ( .A1(n10887), .A2(n10425), .B1(n10889), .B2(n10888), .C1(
        n10784), .C2(n10424), .ZN(n10967) );
  INV_X1 U11169 ( .A(n10967), .ZN(n10440) );
  OAI21_X1 U11170 ( .B1(n5171), .B2(n10427), .A(n10426), .ZN(n10969) );
  AND2_X1 U11171 ( .A1(n5191), .A2(n10433), .ZN(n10429) );
  OR2_X1 U11172 ( .A1(n10429), .A2(n10428), .ZN(n10966) );
  OAI22_X1 U11173 ( .A1(n5074), .A2(n7288), .B1(n10430), .B2(n10907), .ZN(
        n10431) );
  AOI21_X1 U11174 ( .B1(n10433), .B2(n10432), .A(n10431), .ZN(n10434) );
  OAI21_X1 U11175 ( .B1(n10966), .B2(n10435), .A(n10434), .ZN(n10436) );
  AOI21_X1 U11176 ( .B1(n10969), .B2(n10437), .A(n10436), .ZN(n10438) );
  OAI21_X1 U11177 ( .B1(n10440), .B2(n10439), .A(n10438), .ZN(P1_U3278) );
  NAND2_X1 U11178 ( .A1(n10441), .A2(n10778), .ZN(n10442) );
  OAI211_X1 U11179 ( .C1(n10443), .C2(n11015), .A(n10442), .B(n10446), .ZN(
        n10517) );
  MUX2_X1 U11180 ( .A(n10517), .B(P1_REG1_REG_31__SCAN_IN), .S(n5418), .Z(
        P1_U3554) );
  NAND2_X1 U11181 ( .A1(n10444), .A2(n10721), .ZN(n10445) );
  OAI211_X1 U11182 ( .C1(n10447), .C2(n11005), .A(n10446), .B(n10445), .ZN(
        n10518) );
  MUX2_X1 U11183 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10518), .S(n11020), .Z(
        P1_U3553) );
  AOI22_X1 U11184 ( .A1(n10450), .A2(n10778), .B1(n10721), .B2(n10449), .ZN(
        n10451) );
  INV_X1 U11185 ( .A(n10453), .ZN(n10457) );
  AOI22_X1 U11186 ( .A1(n10455), .A2(n10778), .B1(n10721), .B2(n10454), .ZN(
        n10456) );
  OAI211_X1 U11187 ( .C1(n10737), .C2(n10458), .A(n10457), .B(n10456), .ZN(
        n10519) );
  MUX2_X1 U11188 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n10519), .S(n11020), .Z(
        P1_U3551) );
  AOI22_X1 U11189 ( .A1(n10460), .A2(n10778), .B1(n10721), .B2(n10459), .ZN(
        n10461) );
  OAI211_X1 U11190 ( .C1(n10516), .C2(n10463), .A(n10462), .B(n10461), .ZN(
        n10520) );
  MUX2_X1 U11191 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10520), .S(n11020), .Z(
        P1_U3550) );
  AOI22_X1 U11192 ( .A1(n10465), .A2(n10778), .B1(n10721), .B2(n10464), .ZN(
        n10466) );
  OAI211_X1 U11193 ( .C1(n10468), .C2(n10737), .A(n10467), .B(n10466), .ZN(
        n10521) );
  MUX2_X1 U11194 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10521), .S(n11020), .Z(
        P1_U3549) );
  AOI21_X1 U11195 ( .B1(n10721), .B2(n10470), .A(n10469), .ZN(n10471) );
  OAI211_X1 U11196 ( .C1(n10516), .C2(n10473), .A(n10472), .B(n10471), .ZN(
        n10522) );
  MUX2_X1 U11197 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10522), .S(n11020), .Z(
        P1_U3548) );
  AOI211_X1 U11198 ( .C1(n10721), .C2(n10476), .A(n10475), .B(n10474), .ZN(
        n10477) );
  OAI21_X1 U11199 ( .B1(n10516), .B2(n10478), .A(n10477), .ZN(n10523) );
  MUX2_X1 U11200 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10523), .S(n11020), .Z(
        P1_U3547) );
  AOI22_X1 U11201 ( .A1(n10480), .A2(n10778), .B1(n10721), .B2(n10479), .ZN(
        n10481) );
  OAI211_X1 U11202 ( .C1(n10516), .C2(n10483), .A(n10482), .B(n10481), .ZN(
        n10524) );
  MUX2_X1 U11203 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10524), .S(n11020), .Z(
        P1_U3546) );
  AOI211_X1 U11204 ( .C1(n10721), .C2(n10486), .A(n10485), .B(n10484), .ZN(
        n10487) );
  OAI21_X1 U11205 ( .B1(n10516), .B2(n10488), .A(n10487), .ZN(n10525) );
  MUX2_X1 U11206 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10525), .S(n11020), .Z(
        P1_U3545) );
  AOI21_X1 U11207 ( .B1(n10721), .B2(n10490), .A(n10489), .ZN(n10491) );
  OAI211_X1 U11208 ( .C1(n10516), .C2(n10493), .A(n10492), .B(n10491), .ZN(
        n10526) );
  MUX2_X1 U11209 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10526), .S(n11020), .Z(
        P1_U3544) );
  INV_X1 U11210 ( .A(n10516), .ZN(n11018) );
  AND3_X1 U11211 ( .A1(n10495), .A2(n11018), .A3(n10494), .ZN(n10499) );
  OAI22_X1 U11212 ( .A1(n10497), .A2(n11005), .B1(n10496), .B2(n11015), .ZN(
        n10498) );
  MUX2_X1 U11213 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10527), .S(n11020), .Z(
        P1_U3543) );
  AOI211_X1 U11214 ( .C1(n10721), .C2(n10503), .A(n10502), .B(n10501), .ZN(
        n10504) );
  OAI21_X1 U11215 ( .B1(n10516), .B2(n10505), .A(n10504), .ZN(n10528) );
  MUX2_X1 U11216 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10528), .S(n11020), .Z(
        P1_U3542) );
  AOI22_X1 U11217 ( .A1(n10507), .A2(n10778), .B1(n10721), .B2(n10506), .ZN(
        n10508) );
  OAI211_X1 U11218 ( .C1(n10737), .C2(n10510), .A(n10509), .B(n10508), .ZN(
        n10529) );
  MUX2_X1 U11219 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10529), .S(n11020), .Z(
        P1_U3541) );
  AOI211_X1 U11220 ( .C1(n10721), .C2(n10513), .A(n10512), .B(n10511), .ZN(
        n10514) );
  OAI21_X1 U11221 ( .B1(n10516), .B2(n10515), .A(n10514), .ZN(n10530) );
  MUX2_X1 U11222 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10530), .S(n11020), .Z(
        P1_U3539) );
  MUX2_X1 U11223 ( .A(n10517), .B(P1_REG0_REG_31__SCAN_IN), .S(n11021), .Z(
        P1_U3522) );
  MUX2_X1 U11224 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10518), .S(n11024), .Z(
        P1_U3521) );
  MUX2_X1 U11225 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10519), .S(n11024), .Z(
        P1_U3519) );
  MUX2_X1 U11226 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10520), .S(n11024), .Z(
        P1_U3518) );
  MUX2_X1 U11227 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10521), .S(n11024), .Z(
        P1_U3517) );
  MUX2_X1 U11228 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10522), .S(n11024), .Z(
        P1_U3516) );
  MUX2_X1 U11229 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10523), .S(n11024), .Z(
        P1_U3515) );
  MUX2_X1 U11230 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10524), .S(n11024), .Z(
        P1_U3514) );
  MUX2_X1 U11231 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10525), .S(n11024), .Z(
        P1_U3513) );
  MUX2_X1 U11232 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10526), .S(n11024), .Z(
        P1_U3512) );
  MUX2_X1 U11233 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10527), .S(n11024), .Z(
        P1_U3511) );
  MUX2_X1 U11234 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10528), .S(n11024), .Z(
        P1_U3510) );
  MUX2_X1 U11235 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10529), .S(n11024), .Z(
        P1_U3508) );
  MUX2_X1 U11236 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10530), .S(n11024), .Z(
        P1_U3502) );
  MUX2_X1 U11237 ( .A(P1_D_REG_0__SCAN_IN), .B(n10532), .S(n10531), .Z(
        P1_U3440) );
  INV_X1 U11238 ( .A(n10533), .ZN(n10536) );
  NAND3_X1 U11239 ( .A1(n10534), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n10535) );
  OAI22_X1 U11240 ( .A1(n10536), .A2(n10535), .B1(n7364), .B2(n10546), .ZN(
        n10537) );
  AOI21_X1 U11241 ( .B1(n10539), .B2(n10538), .A(n10537), .ZN(n10540) );
  INV_X1 U11242 ( .A(n10540), .ZN(P1_U3322) );
  OAI222_X1 U11243 ( .A1(P1_U3084), .A2(n10543), .B1(n8088), .B2(n10542), .C1(
        n10541), .C2(n10546), .ZN(P1_U3324) );
  OAI222_X1 U11244 ( .A1(P1_U3084), .A2(n7264), .B1(n8088), .B2(n10545), .C1(
        n10544), .C2(n10546), .ZN(P1_U3326) );
  OAI222_X1 U11245 ( .A1(n10549), .A2(P1_U3084), .B1(n8088), .B2(n10548), .C1(
        n10547), .C2(n10546), .ZN(P1_U3327) );
  MUX2_X1 U11246 ( .A(n10550), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NOR2_X1 U11247 ( .A1(n10551), .A2(n10623), .ZN(n10583) );
  NOR2_X1 U11248 ( .A1(n10571), .A2(n10552), .ZN(P1_U3321) );
  INV_X1 U11249 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10553) );
  NOR2_X1 U11250 ( .A1(n10571), .A2(n10553), .ZN(P1_U3320) );
  INV_X1 U11251 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10554) );
  NOR2_X1 U11252 ( .A1(n10571), .A2(n10554), .ZN(P1_U3319) );
  INV_X1 U11253 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10555) );
  NOR2_X1 U11254 ( .A1(n10571), .A2(n10555), .ZN(P1_U3318) );
  INV_X1 U11255 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10556) );
  NOR2_X1 U11256 ( .A1(n10571), .A2(n10556), .ZN(P1_U3317) );
  INV_X1 U11257 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10557) );
  NOR2_X1 U11258 ( .A1(n10571), .A2(n10557), .ZN(P1_U3316) );
  INV_X1 U11259 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10558) );
  NOR2_X1 U11260 ( .A1(n10571), .A2(n10558), .ZN(P1_U3315) );
  INV_X1 U11261 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10559) );
  NOR2_X1 U11262 ( .A1(n10571), .A2(n10559), .ZN(P1_U3314) );
  INV_X1 U11263 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10560) );
  NOR2_X1 U11264 ( .A1(n10571), .A2(n10560), .ZN(P1_U3313) );
  INV_X1 U11265 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10561) );
  NOR2_X1 U11266 ( .A1(n10571), .A2(n10561), .ZN(P1_U3312) );
  INV_X1 U11267 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10562) );
  NOR2_X1 U11268 ( .A1(n10571), .A2(n10562), .ZN(P1_U3311) );
  INV_X1 U11269 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10563) );
  NOR2_X1 U11270 ( .A1(n10571), .A2(n10563), .ZN(P1_U3310) );
  INV_X1 U11271 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10564) );
  NOR2_X1 U11272 ( .A1(n10571), .A2(n10564), .ZN(P1_U3309) );
  INV_X1 U11273 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10565) );
  NOR2_X1 U11274 ( .A1(n10571), .A2(n10565), .ZN(P1_U3308) );
  INV_X1 U11275 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10566) );
  NOR2_X1 U11276 ( .A1(n10571), .A2(n10566), .ZN(P1_U3307) );
  INV_X1 U11277 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10567) );
  NOR2_X1 U11278 ( .A1(n10571), .A2(n10567), .ZN(P1_U3306) );
  INV_X1 U11279 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10568) );
  NOR2_X1 U11280 ( .A1(n10571), .A2(n10568), .ZN(P1_U3305) );
  INV_X1 U11281 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10569) );
  NOR2_X1 U11282 ( .A1(n10571), .A2(n10569), .ZN(P1_U3304) );
  INV_X1 U11283 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10570) );
  NOR2_X1 U11284 ( .A1(n10571), .A2(n10570), .ZN(P1_U3303) );
  INV_X1 U11285 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10572) );
  NOR2_X1 U11286 ( .A1(n10583), .A2(n10572), .ZN(P1_U3302) );
  INV_X1 U11287 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10573) );
  NOR2_X1 U11288 ( .A1(n10583), .A2(n10573), .ZN(P1_U3301) );
  INV_X1 U11289 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10574) );
  NOR2_X1 U11290 ( .A1(n10583), .A2(n10574), .ZN(P1_U3300) );
  INV_X1 U11291 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10575) );
  NOR2_X1 U11292 ( .A1(n10583), .A2(n10575), .ZN(P1_U3299) );
  INV_X1 U11293 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10576) );
  NOR2_X1 U11294 ( .A1(n10583), .A2(n10576), .ZN(P1_U3298) );
  INV_X1 U11295 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10577) );
  NOR2_X1 U11296 ( .A1(n10583), .A2(n10577), .ZN(P1_U3297) );
  INV_X1 U11297 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10578) );
  NOR2_X1 U11298 ( .A1(n10583), .A2(n10578), .ZN(P1_U3296) );
  INV_X1 U11299 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10579) );
  NOR2_X1 U11300 ( .A1(n10583), .A2(n10579), .ZN(P1_U3295) );
  INV_X1 U11301 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10580) );
  NOR2_X1 U11302 ( .A1(n10583), .A2(n10580), .ZN(P1_U3294) );
  INV_X1 U11303 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10581) );
  NOR2_X1 U11304 ( .A1(n10583), .A2(n10581), .ZN(P1_U3293) );
  INV_X1 U11305 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10582) );
  NOR2_X1 U11306 ( .A1(n10583), .A2(n10582), .ZN(P1_U3292) );
  AND2_X1 U11307 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10584), .ZN(P2_U3326) );
  AND2_X1 U11308 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10584), .ZN(P2_U3325) );
  AND2_X1 U11309 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10584), .ZN(P2_U3324) );
  AND2_X1 U11310 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10584), .ZN(P2_U3323) );
  AND2_X1 U11311 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10584), .ZN(P2_U3322) );
  AND2_X1 U11312 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10584), .ZN(P2_U3321) );
  AND2_X1 U11313 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10584), .ZN(P2_U3320) );
  AND2_X1 U11314 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10584), .ZN(P2_U3319) );
  AND2_X1 U11315 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10584), .ZN(P2_U3318) );
  AND2_X1 U11316 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10584), .ZN(P2_U3317) );
  AND2_X1 U11317 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10584), .ZN(P2_U3316) );
  AND2_X1 U11318 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10584), .ZN(P2_U3315) );
  AND2_X1 U11319 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10584), .ZN(P2_U3314) );
  AND2_X1 U11320 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10584), .ZN(P2_U3313) );
  AND2_X1 U11321 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10584), .ZN(P2_U3312) );
  AND2_X1 U11322 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10584), .ZN(P2_U3311) );
  AND2_X1 U11323 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n5192), .ZN(P2_U3310) );
  AND2_X1 U11324 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n5192), .ZN(P2_U3309) );
  AND2_X1 U11325 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n5192), .ZN(P2_U3308) );
  AND2_X1 U11326 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n5192), .ZN(P2_U3307) );
  AND2_X1 U11327 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n5192), .ZN(P2_U3306) );
  AND2_X1 U11328 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n5192), .ZN(P2_U3305) );
  AND2_X1 U11329 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n5192), .ZN(P2_U3304) );
  AND2_X1 U11330 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n5192), .ZN(P2_U3303) );
  AND2_X1 U11331 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n5192), .ZN(P2_U3302) );
  AND2_X1 U11332 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n5192), .ZN(P2_U3301) );
  AND2_X1 U11333 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n5192), .ZN(P2_U3300) );
  AND2_X1 U11334 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n5192), .ZN(P2_U3299) );
  AND2_X1 U11335 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n5192), .ZN(P2_U3298) );
  AND2_X1 U11336 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n5192), .ZN(P2_U3297) );
  XOR2_X1 U11337 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  INV_X1 U11338 ( .A(n10585), .ZN(n10586) );
  NAND2_X1 U11339 ( .A1(n10587), .A2(n10586), .ZN(n10588) );
  XNOR2_X1 U11340 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10588), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11341 ( .A(n10590), .B(n10589), .Z(ADD_1071_U54) );
  XOR2_X1 U11342 ( .A(n10592), .B(n10591), .Z(ADD_1071_U53) );
  XNOR2_X1 U11343 ( .A(n10594), .B(n10593), .ZN(ADD_1071_U52) );
  NOR2_X1 U11344 ( .A1(n10596), .A2(n10595), .ZN(n10597) );
  XOR2_X1 U11345 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n10597), .Z(ADD_1071_U51) );
  XOR2_X1 U11346 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10598), .Z(ADD_1071_U50) );
  XOR2_X1 U11347 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10599), .Z(ADD_1071_U49) );
  XOR2_X1 U11348 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10600), .Z(ADD_1071_U48) );
  XOR2_X1 U11349 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n10601), .Z(ADD_1071_U47) );
  XOR2_X1 U11350 ( .A(n10603), .B(n10602), .Z(ADD_1071_U63) );
  XOR2_X1 U11351 ( .A(n10605), .B(n10604), .Z(ADD_1071_U62) );
  XNOR2_X1 U11352 ( .A(n10607), .B(n10606), .ZN(ADD_1071_U61) );
  XNOR2_X1 U11353 ( .A(n10609), .B(n10608), .ZN(ADD_1071_U60) );
  XNOR2_X1 U11354 ( .A(n10611), .B(n10610), .ZN(ADD_1071_U59) );
  XNOR2_X1 U11355 ( .A(n10613), .B(n10612), .ZN(ADD_1071_U58) );
  XNOR2_X1 U11356 ( .A(n10615), .B(n10614), .ZN(ADD_1071_U57) );
  XNOR2_X1 U11357 ( .A(n10617), .B(n10616), .ZN(ADD_1071_U56) );
  NOR2_X1 U11358 ( .A1(n10619), .A2(n10618), .ZN(n10620) );
  XOR2_X1 U11359 ( .A(P1_ADDR_REG_18__SCAN_IN), .B(n10620), .Z(ADD_1071_U55)
         );
  INV_X1 U11360 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10622) );
  AOI21_X1 U11361 ( .B1(n10623), .B2(n10622), .A(n10621), .ZN(P1_U3441) );
  OAI22_X1 U11362 ( .A1(n10659), .A2(n10625), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10624), .ZN(n10626) );
  INV_X1 U11363 ( .A(n10626), .ZN(n10639) );
  AOI211_X1 U11364 ( .C1(n10630), .C2(n10629), .A(n10628), .B(n10627), .ZN(
        n10631) );
  AOI21_X1 U11365 ( .B1(n10670), .B2(P1_ADDR_REG_1__SCAN_IN), .A(n10631), .ZN(
        n10638) );
  NOR2_X1 U11366 ( .A1(n10633), .A2(n10632), .ZN(n10636) );
  OAI211_X1 U11367 ( .C1(n10636), .C2(n10635), .A(n10662), .B(n10634), .ZN(
        n10637) );
  NAND3_X1 U11368 ( .A1(n10639), .A2(n10638), .A3(n10637), .ZN(P1_U3242) );
  OAI22_X1 U11369 ( .A1(n10641), .A2(n10640), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10701), .ZN(n10647) );
  AOI211_X1 U11370 ( .C1(n10645), .C2(n10644), .A(n10643), .B(n10642), .ZN(
        n10646) );
  AOI211_X1 U11371 ( .C1(n10649), .C2(n10648), .A(n10647), .B(n10646), .ZN(
        n10656) );
  INV_X1 U11372 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10650) );
  INV_X1 U11373 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10684) );
  NOR2_X1 U11374 ( .A1(n10650), .A2(n10684), .ZN(n10654) );
  OAI211_X1 U11375 ( .C1(n10654), .C2(n10653), .A(n10652), .B(n10651), .ZN(
        n10655) );
  NAND2_X1 U11376 ( .A1(n10656), .A2(n10655), .ZN(P2_U3246) );
  XNOR2_X1 U11377 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  OAI22_X1 U11378 ( .A1(n10659), .A2(n10658), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10657), .ZN(n10660) );
  INV_X1 U11379 ( .A(n10660), .ZN(n10676) );
  OAI211_X1 U11380 ( .C1(n10664), .C2(n10663), .A(n10662), .B(n10661), .ZN(
        n10673) );
  AOI21_X1 U11381 ( .B1(n10667), .B2(n10666), .A(n10665), .ZN(n10668) );
  NAND2_X1 U11382 ( .A1(n10669), .A2(n10668), .ZN(n10672) );
  NAND2_X1 U11383 ( .A1(n10670), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n10671) );
  AND3_X1 U11384 ( .A1(n10673), .A2(n10672), .A3(n10671), .ZN(n10675) );
  NAND3_X1 U11385 ( .A1(n10676), .A2(n10675), .A3(n10674), .ZN(P1_U3243) );
  INV_X1 U11386 ( .A(n10677), .ZN(n10678) );
  NAND2_X1 U11387 ( .A1(n10678), .A2(n10995), .ZN(n10682) );
  NAND2_X1 U11388 ( .A1(n10680), .A2(n10679), .ZN(n10681) );
  AND3_X1 U11389 ( .A1(n10683), .A2(n10682), .A3(n10681), .ZN(n10686) );
  AOI22_X1 U11390 ( .A1(n10998), .A2(n10686), .B1(n10684), .B2(n10997), .ZN(
        P2_U3520) );
  INV_X1 U11391 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10685) );
  AOI22_X1 U11392 ( .A1(n11002), .A2(n10686), .B1(n10685), .B2(n10999), .ZN(
        P2_U3451) );
  AOI21_X1 U11393 ( .B1(n10737), .B2(n10895), .A(n10687), .ZN(n10691) );
  NOR2_X1 U11394 ( .A1(n10688), .A2(n11015), .ZN(n10690) );
  NOR4_X1 U11395 ( .A1(n10692), .A2(n10691), .A3(n10690), .A4(n10689), .ZN(
        n10694) );
  AOI22_X1 U11396 ( .A1(n11020), .A2(n10694), .B1(n7243), .B2(n5418), .ZN(
        P1_U3524) );
  INV_X1 U11397 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10693) );
  AOI22_X1 U11398 ( .A1(n11024), .A2(n10694), .B1(n10693), .B2(n11021), .ZN(
        P1_U3457) );
  XNOR2_X1 U11399 ( .A(n10704), .B(n10695), .ZN(n10697) );
  AOI21_X1 U11400 ( .B1(n10697), .B2(n10929), .A(n10696), .ZN(n10713) );
  OAI21_X1 U11401 ( .B1(n10711), .B2(n10699), .A(n10698), .ZN(n10712) );
  OAI22_X1 U11402 ( .A1(n10702), .A2(n10712), .B1(n10701), .B2(n10700), .ZN(
        n10708) );
  XNOR2_X1 U11403 ( .A(n10704), .B(n10703), .ZN(n10710) );
  OAI22_X1 U11404 ( .A1(n10710), .A2(n10706), .B1(n10705), .B2(n10711), .ZN(
        n10707) );
  AOI211_X1 U11405 ( .C1(n10949), .C2(P2_REG2_REG_1__SCAN_IN), .A(n10708), .B(
        n10707), .ZN(n10709) );
  OAI21_X1 U11406 ( .B1(n10949), .B2(n10713), .A(n10709), .ZN(P2_U3295) );
  INV_X1 U11407 ( .A(n10710), .ZN(n10716) );
  OAI22_X1 U11408 ( .A1(n10712), .A2(n10991), .B1(n10711), .B2(n10989), .ZN(
        n10715) );
  INV_X1 U11409 ( .A(n10713), .ZN(n10714) );
  AOI211_X1 U11410 ( .C1(n10995), .C2(n10716), .A(n10715), .B(n10714), .ZN(
        n10719) );
  AOI22_X1 U11411 ( .A1(n10998), .A2(n10719), .B1(n10717), .B2(n10997), .ZN(
        P2_U3521) );
  INV_X1 U11412 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10718) );
  AOI22_X1 U11413 ( .A1(n11002), .A2(n10719), .B1(n10718), .B2(n10999), .ZN(
        P2_U3454) );
  AOI22_X1 U11414 ( .A1(n10722), .A2(n10778), .B1(n10721), .B2(n10720), .ZN(
        n10723) );
  OAI21_X1 U11415 ( .B1(n10724), .B2(n10737), .A(n10723), .ZN(n10725) );
  NOR2_X1 U11416 ( .A1(n10726), .A2(n10725), .ZN(n10728) );
  AOI22_X1 U11417 ( .A1(n11020), .A2(n10728), .B1(n7242), .B2(n5418), .ZN(
        P1_U3525) );
  INV_X1 U11418 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10727) );
  AOI22_X1 U11419 ( .A1(n11024), .A2(n10728), .B1(n10727), .B2(n11021), .ZN(
        P1_U3460) );
  INV_X1 U11420 ( .A(n10729), .ZN(n10876) );
  OAI22_X1 U11421 ( .A1(n10731), .A2(n10991), .B1(n10730), .B2(n10989), .ZN(
        n10733) );
  AOI211_X1 U11422 ( .C1(n10876), .C2(n10734), .A(n10733), .B(n10732), .ZN(
        n10736) );
  AOI22_X1 U11423 ( .A1(n10998), .A2(n10736), .B1(n7376), .B2(n10997), .ZN(
        P2_U3522) );
  INV_X1 U11424 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10735) );
  AOI22_X1 U11425 ( .A1(n11002), .A2(n10736), .B1(n10735), .B2(n10999), .ZN(
        P2_U3457) );
  INV_X1 U11426 ( .A(n10737), .ZN(n11010) );
  XNOR2_X1 U11427 ( .A(n10738), .B(n10741), .ZN(n10754) );
  OAI21_X1 U11428 ( .B1(n10740), .B2(n10755), .A(n10739), .ZN(n10752) );
  OAI22_X1 U11429 ( .A1(n10752), .A2(n11005), .B1(n10755), .B2(n11015), .ZN(
        n10748) );
  XNOR2_X1 U11430 ( .A(n10742), .B(n10741), .ZN(n10747) );
  OAI22_X1 U11431 ( .A1(n10783), .A2(n10887), .B1(n10743), .B2(n10889), .ZN(
        n10744) );
  AOI21_X1 U11432 ( .B1(n10754), .B2(n10745), .A(n10744), .ZN(n10746) );
  OAI21_X1 U11433 ( .B1(n10747), .B2(n10784), .A(n10746), .ZN(n10759) );
  AOI211_X1 U11434 ( .C1(n11010), .C2(n10754), .A(n10748), .B(n10759), .ZN(
        n10750) );
  AOI22_X1 U11435 ( .A1(n11020), .A2(n10750), .B1(n7241), .B2(n5418), .ZN(
        P1_U3526) );
  INV_X1 U11436 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10749) );
  AOI22_X1 U11437 ( .A1(n11024), .A2(n10750), .B1(n10749), .B2(n11021), .ZN(
        P1_U3463) );
  INV_X1 U11438 ( .A(n10751), .ZN(n10903) );
  INV_X1 U11439 ( .A(n10752), .ZN(n10753) );
  AOI22_X1 U11440 ( .A1(n10754), .A2(n10903), .B1(n10902), .B2(n10753), .ZN(
        n10761) );
  NOR2_X1 U11441 ( .A1(n10905), .A2(n10755), .ZN(n10758) );
  OAI22_X1 U11442 ( .A1(n5074), .A2(n10756), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10907), .ZN(n10757) );
  AOI211_X1 U11443 ( .C1(n10759), .C2(n5074), .A(n10758), .B(n10757), .ZN(
        n10760) );
  NAND2_X1 U11444 ( .A1(n10761), .A2(n10760), .ZN(P1_U3288) );
  OAI22_X1 U11445 ( .A1(n10763), .A2(n11005), .B1(n10762), .B2(n11015), .ZN(
        n10765) );
  AOI211_X1 U11446 ( .C1(n11010), .C2(n10766), .A(n10765), .B(n10764), .ZN(
        n10767) );
  AOI22_X1 U11447 ( .A1(n11020), .A2(n10767), .B1(n6779), .B2(n5418), .ZN(
        P1_U3527) );
  AOI22_X1 U11448 ( .A1(n11024), .A2(n10767), .B1(n6780), .B2(n11021), .ZN(
        P1_U3466) );
  OAI22_X1 U11449 ( .A1(n10769), .A2(n10991), .B1(n10768), .B2(n10989), .ZN(
        n10771) );
  AOI211_X1 U11450 ( .C1(n10995), .C2(n10772), .A(n10771), .B(n10770), .ZN(
        n10774) );
  AOI22_X1 U11451 ( .A1(n10998), .A2(n10774), .B1(n7378), .B2(n10997), .ZN(
        P2_U3524) );
  INV_X1 U11452 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U11453 ( .A1(n11002), .A2(n10774), .B1(n10773), .B2(n10999), .ZN(
        P2_U3463) );
  XNOR2_X1 U11454 ( .A(n10775), .B(n10781), .ZN(n10798) );
  INV_X1 U11455 ( .A(n10776), .ZN(n10779) );
  OAI211_X1 U11456 ( .C1(n10779), .C2(n10780), .A(n10778), .B(n10777), .ZN(
        n10795) );
  OAI21_X1 U11457 ( .B1(n10780), .B2(n11015), .A(n10795), .ZN(n10787) );
  XNOR2_X1 U11458 ( .A(n10782), .B(n10781), .ZN(n10785) );
  OAI222_X1 U11459 ( .A1(n10887), .A2(n10786), .B1(n10785), .B2(n10784), .C1(
        n10889), .C2(n10783), .ZN(n10796) );
  AOI211_X1 U11460 ( .C1(n11018), .C2(n10798), .A(n10787), .B(n10796), .ZN(
        n10788) );
  AOI22_X1 U11461 ( .A1(n11020), .A2(n10788), .B1(n7240), .B2(n5418), .ZN(
        P1_U3528) );
  AOI22_X1 U11462 ( .A1(n11024), .A2(n10788), .B1(n6799), .B2(n11021), .ZN(
        P1_U3469) );
  AOI22_X1 U11463 ( .A1(n10792), .A2(n10791), .B1(n10790), .B2(n10789), .ZN(
        n10793) );
  OAI21_X1 U11464 ( .B1(n10795), .B2(n5073), .A(n10793), .ZN(n10797) );
  AOI211_X1 U11465 ( .C1(n10799), .C2(n10798), .A(n10797), .B(n10796), .ZN(
        n10800) );
  AOI22_X1 U11466 ( .A1(n10439), .A2(n6800), .B1(n10800), .B2(n5074), .ZN(
        P1_U3286) );
  OAI21_X1 U11467 ( .B1(n10802), .B2(n10989), .A(n10801), .ZN(n10804) );
  AOI211_X1 U11468 ( .C1(n10805), .C2(n10995), .A(n10804), .B(n10803), .ZN(
        n10807) );
  AOI22_X1 U11469 ( .A1(n10998), .A2(n10807), .B1(n7374), .B2(n10997), .ZN(
        P2_U3525) );
  INV_X1 U11470 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10806) );
  AOI22_X1 U11471 ( .A1(n11002), .A2(n10807), .B1(n10806), .B2(n10999), .ZN(
        P2_U3466) );
  NAND2_X1 U11472 ( .A1(n10808), .A2(n11018), .ZN(n10810) );
  OAI211_X1 U11473 ( .C1(n10811), .C2(n11015), .A(n10810), .B(n10809), .ZN(
        n10812) );
  NOR2_X1 U11474 ( .A1(n10813), .A2(n10812), .ZN(n10815) );
  AOI22_X1 U11475 ( .A1(n11020), .A2(n10815), .B1(n7239), .B2(n5418), .ZN(
        P1_U3529) );
  INV_X1 U11476 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10814) );
  AOI22_X1 U11477 ( .A1(n11024), .A2(n10815), .B1(n10814), .B2(n11021), .ZN(
        P1_U3472) );
  INV_X1 U11478 ( .A(n10816), .ZN(n10823) );
  AND3_X1 U11479 ( .A1(n10818), .A2(n10995), .A3(n10817), .ZN(n10822) );
  OAI22_X1 U11480 ( .A1(n10820), .A2(n10991), .B1(n10819), .B2(n10989), .ZN(
        n10821) );
  NOR3_X1 U11481 ( .A1(n10823), .A2(n10822), .A3(n10821), .ZN(n10826) );
  AOI22_X1 U11482 ( .A1(n10998), .A2(n10826), .B1(n10824), .B2(n10997), .ZN(
        P2_U3526) );
  INV_X1 U11483 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10825) );
  AOI22_X1 U11484 ( .A1(n11002), .A2(n10826), .B1(n10825), .B2(n10999), .ZN(
        P2_U3469) );
  OAI21_X1 U11485 ( .B1(n10828), .B2(n11015), .A(n10827), .ZN(n10830) );
  AOI211_X1 U11486 ( .C1(n11010), .C2(n10831), .A(n10830), .B(n10829), .ZN(
        n10833) );
  AOI22_X1 U11487 ( .A1(n11020), .A2(n10833), .B1(n7248), .B2(n5418), .ZN(
        P1_U3530) );
  INV_X1 U11488 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10832) );
  AOI22_X1 U11489 ( .A1(n11024), .A2(n10833), .B1(n10832), .B2(n11021), .ZN(
        P1_U3475) );
  OAI22_X1 U11490 ( .A1(n10835), .A2(n10991), .B1(n10834), .B2(n10989), .ZN(
        n10837) );
  AOI211_X1 U11491 ( .C1(n10995), .C2(n10838), .A(n10837), .B(n10836), .ZN(
        n10841) );
  AOI22_X1 U11492 ( .A1(n10998), .A2(n10841), .B1(n10839), .B2(n10997), .ZN(
        P2_U3527) );
  INV_X1 U11493 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10840) );
  AOI22_X1 U11494 ( .A1(n11002), .A2(n10841), .B1(n10840), .B2(n10999), .ZN(
        P2_U3472) );
  INV_X1 U11495 ( .A(n10842), .ZN(n10847) );
  OAI22_X1 U11496 ( .A1(n10844), .A2(n11005), .B1(n10843), .B2(n11015), .ZN(
        n10846) );
  AOI211_X1 U11497 ( .C1(n11010), .C2(n10847), .A(n10846), .B(n10845), .ZN(
        n10848) );
  AOI22_X1 U11498 ( .A1(n11020), .A2(n10848), .B1(n7250), .B2(n5418), .ZN(
        P1_U3531) );
  AOI22_X1 U11499 ( .A1(n11024), .A2(n10848), .B1(n6857), .B2(n11021), .ZN(
        P1_U3478) );
  NAND3_X1 U11500 ( .A1(n10850), .A2(n10849), .A3(n10995), .ZN(n10855) );
  NAND2_X1 U11501 ( .A1(n10852), .A2(n10851), .ZN(n10853) );
  AND4_X1 U11502 ( .A1(n10856), .A2(n10855), .A3(n10854), .A4(n10853), .ZN(
        n10858) );
  AOI22_X1 U11503 ( .A1(n10998), .A2(n10858), .B1(n10857), .B2(n10997), .ZN(
        P2_U3528) );
  AOI22_X1 U11504 ( .A1(n11002), .A2(n10858), .B1(n5879), .B2(n10999), .ZN(
        P2_U3475) );
  OAI22_X1 U11505 ( .A1(n10859), .A2(n11005), .B1(n5390), .B2(n11015), .ZN(
        n10861) );
  AOI211_X1 U11506 ( .C1(n10862), .C2(n11018), .A(n10861), .B(n10860), .ZN(
        n10864) );
  AOI22_X1 U11507 ( .A1(n11020), .A2(n10864), .B1(n7253), .B2(n5418), .ZN(
        P1_U3532) );
  INV_X1 U11508 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10863) );
  AOI22_X1 U11509 ( .A1(n11024), .A2(n10864), .B1(n10863), .B2(n11021), .ZN(
        P1_U3481) );
  INV_X1 U11510 ( .A(n10865), .ZN(n10866) );
  OAI22_X1 U11511 ( .A1(n10867), .A2(n10991), .B1(n10866), .B2(n10989), .ZN(
        n10869) );
  AOI211_X1 U11512 ( .C1(n10876), .C2(n10870), .A(n10869), .B(n10868), .ZN(
        n10872) );
  AOI22_X1 U11513 ( .A1(n10998), .A2(n10872), .B1(n10871), .B2(n10997), .ZN(
        P2_U3529) );
  AOI22_X1 U11514 ( .A1(n11002), .A2(n10872), .B1(n5892), .B2(n10999), .ZN(
        P2_U3478) );
  OAI22_X1 U11515 ( .A1(n10874), .A2(n10991), .B1(n10873), .B2(n10989), .ZN(
        n10875) );
  AOI21_X1 U11516 ( .B1(n10877), .B2(n10876), .A(n10875), .ZN(n10878) );
  AND2_X1 U11517 ( .A1(n10879), .A2(n10878), .ZN(n10881) );
  AOI22_X1 U11518 ( .A1(n10998), .A2(n10881), .B1(n7716), .B2(n10997), .ZN(
        P2_U3530) );
  INV_X1 U11519 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10880) );
  AOI22_X1 U11520 ( .A1(n11002), .A2(n10881), .B1(n10880), .B2(n10999), .ZN(
        P2_U3481) );
  XNOR2_X1 U11521 ( .A(n10882), .B(n10886), .ZN(n10896) );
  INV_X1 U11522 ( .A(n10896), .ZN(n10904) );
  OAI21_X1 U11523 ( .B1(n10884), .B2(n10906), .A(n10883), .ZN(n10900) );
  OAI22_X1 U11524 ( .A1(n10900), .A2(n11005), .B1(n10906), .B2(n11015), .ZN(
        n10897) );
  XOR2_X1 U11525 ( .A(n10886), .B(n10885), .Z(n10893) );
  OAI22_X1 U11526 ( .A1(n10890), .A2(n10889), .B1(n10888), .B2(n10887), .ZN(
        n10891) );
  AOI21_X1 U11527 ( .B1(n10893), .B2(n10892), .A(n10891), .ZN(n10894) );
  OAI21_X1 U11528 ( .B1(n10896), .B2(n10895), .A(n10894), .ZN(n10912) );
  AOI211_X1 U11529 ( .C1(n11010), .C2(n10904), .A(n10897), .B(n10912), .ZN(
        n10899) );
  AOI22_X1 U11530 ( .A1(n11020), .A2(n10899), .B1(n7255), .B2(n5418), .ZN(
        P1_U3534) );
  INV_X1 U11531 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10898) );
  AOI22_X1 U11532 ( .A1(n11024), .A2(n10899), .B1(n10898), .B2(n11021), .ZN(
        P1_U3487) );
  INV_X1 U11533 ( .A(n10900), .ZN(n10901) );
  AOI22_X1 U11534 ( .A1(n10904), .A2(n10903), .B1(n10902), .B2(n10901), .ZN(
        n10914) );
  NOR2_X1 U11535 ( .A1(n10906), .A2(n10905), .ZN(n10911) );
  OAI22_X1 U11536 ( .A1(n5074), .A2(n10909), .B1(n10908), .B2(n10907), .ZN(
        n10910) );
  AOI211_X1 U11537 ( .C1(n10912), .C2(n5074), .A(n10911), .B(n10910), .ZN(
        n10913) );
  NAND2_X1 U11538 ( .A1(n10914), .A2(n10913), .ZN(P1_U3280) );
  OAI21_X1 U11539 ( .B1(n10916), .B2(n10919), .A(n10915), .ZN(n10917) );
  INV_X1 U11540 ( .A(n10917), .ZN(n10946) );
  INV_X1 U11541 ( .A(n10918), .ZN(n10923) );
  NAND3_X1 U11542 ( .A1(n10921), .A2(n10920), .A3(n10919), .ZN(n10922) );
  NAND2_X1 U11543 ( .A1(n10923), .A2(n10922), .ZN(n10928) );
  AOI222_X1 U11544 ( .A1(n10929), .A2(n10928), .B1(n10927), .B2(n10926), .C1(
        n10925), .C2(n10924), .ZN(n10941) );
  OAI211_X1 U11545 ( .C1(n10931), .C2(n10932), .A(n10930), .B(n5188), .ZN(
        n10942) );
  OAI211_X1 U11546 ( .C1(n10932), .C2(n10989), .A(n10941), .B(n10942), .ZN(
        n10933) );
  AOI21_X1 U11547 ( .B1(n10946), .B2(n10995), .A(n10933), .ZN(n10935) );
  AOI22_X1 U11548 ( .A1(n10998), .A2(n10935), .B1(n7829), .B2(n10997), .ZN(
        P2_U3531) );
  INV_X1 U11549 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10934) );
  AOI22_X1 U11550 ( .A1(n11002), .A2(n10935), .B1(n10934), .B2(n10999), .ZN(
        P2_U3484) );
  INV_X1 U11551 ( .A(n10936), .ZN(n10937) );
  AOI22_X1 U11552 ( .A1(n10939), .A2(n5182), .B1(n10938), .B2(n10937), .ZN(
        n10940) );
  OAI211_X1 U11553 ( .C1(n10943), .C2(n10942), .A(n10941), .B(n10940), .ZN(
        n10944) );
  AOI21_X1 U11554 ( .B1(n10946), .B2(n10945), .A(n10944), .ZN(n10948) );
  AOI22_X1 U11555 ( .A1(n10949), .A2(n5933), .B1(n10948), .B2(n10947), .ZN(
        P2_U3285) );
  INV_X1 U11556 ( .A(n10950), .ZN(n10955) );
  OAI21_X1 U11557 ( .B1(n10952), .B2(n11015), .A(n10951), .ZN(n10954) );
  AOI211_X1 U11558 ( .C1(n10955), .C2(n11018), .A(n10954), .B(n10953), .ZN(
        n10957) );
  AOI22_X1 U11559 ( .A1(n11020), .A2(n10957), .B1(n7238), .B2(n5418), .ZN(
        P1_U3535) );
  INV_X1 U11560 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10956) );
  AOI22_X1 U11561 ( .A1(n11024), .A2(n10957), .B1(n10956), .B2(n11021), .ZN(
        P1_U3490) );
  OAI22_X1 U11562 ( .A1(n10959), .A2(n10991), .B1(n10958), .B2(n10989), .ZN(
        n10961) );
  AOI211_X1 U11563 ( .C1(n10962), .C2(n10995), .A(n10961), .B(n10960), .ZN(
        n10964) );
  AOI22_X1 U11564 ( .A1(n10998), .A2(n10964), .B1(n10963), .B2(n10997), .ZN(
        P2_U3532) );
  AOI22_X1 U11565 ( .A1(n11002), .A2(n10964), .B1(n5957), .B2(n10999), .ZN(
        P2_U3487) );
  OAI22_X1 U11566 ( .A1(n10966), .A2(n11005), .B1(n10965), .B2(n11015), .ZN(
        n10968) );
  AOI211_X1 U11567 ( .C1(n11018), .C2(n10969), .A(n10968), .B(n10967), .ZN(
        n10971) );
  AOI22_X1 U11568 ( .A1(n11020), .A2(n10971), .B1(n7237), .B2(n5418), .ZN(
        P1_U3536) );
  INV_X1 U11569 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10970) );
  AOI22_X1 U11570 ( .A1(n11024), .A2(n10971), .B1(n10970), .B2(n11021), .ZN(
        P1_U3493) );
  NOR2_X1 U11571 ( .A1(n10973), .A2(n10972), .ZN(n10978) );
  OAI22_X1 U11572 ( .A1(n10975), .A2(n10991), .B1(n10974), .B2(n10989), .ZN(
        n10977) );
  AOI211_X1 U11573 ( .C1(n10978), .C2(n9507), .A(n10977), .B(n10976), .ZN(
        n10980) );
  AOI22_X1 U11574 ( .A1(n10998), .A2(n10980), .B1(n5971), .B2(n10997), .ZN(
        P2_U3533) );
  INV_X1 U11575 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10979) );
  AOI22_X1 U11576 ( .A1(n11002), .A2(n10980), .B1(n10979), .B2(n10999), .ZN(
        P2_U3490) );
  OAI211_X1 U11577 ( .C1(n10983), .C2(n11015), .A(n10982), .B(n10981), .ZN(
        n10984) );
  AOI21_X1 U11578 ( .B1(n11018), .B2(n10985), .A(n10984), .ZN(n10987) );
  AOI22_X1 U11579 ( .A1(n11020), .A2(n10987), .B1(n6976), .B2(n5418), .ZN(
        P1_U3537) );
  INV_X1 U11580 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10986) );
  AOI22_X1 U11581 ( .A1(n11024), .A2(n10987), .B1(n10986), .B2(n11021), .ZN(
        P1_U3496) );
  INV_X1 U11582 ( .A(n10988), .ZN(n10996) );
  OAI22_X1 U11583 ( .A1(n10992), .A2(n10991), .B1(n10990), .B2(n10989), .ZN(
        n10993) );
  AOI211_X1 U11584 ( .C1(n10996), .C2(n10995), .A(n10994), .B(n10993), .ZN(
        n11001) );
  AOI22_X1 U11585 ( .A1(n10998), .A2(n11001), .B1(n5994), .B2(n10997), .ZN(
        P2_U3534) );
  INV_X1 U11586 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n11000) );
  AOI22_X1 U11587 ( .A1(n11002), .A2(n11001), .B1(n11000), .B2(n10999), .ZN(
        P2_U3493) );
  INV_X1 U11588 ( .A(n11003), .ZN(n11009) );
  OAI22_X1 U11589 ( .A1(n11006), .A2(n11005), .B1(n11004), .B2(n11015), .ZN(
        n11008) );
  AOI211_X1 U11590 ( .C1(n11010), .C2(n11009), .A(n11008), .B(n11007), .ZN(
        n11012) );
  AOI22_X1 U11591 ( .A1(n11020), .A2(n11012), .B1(n6690), .B2(n5418), .ZN(
        P1_U3538) );
  INV_X1 U11592 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n11011) );
  AOI22_X1 U11593 ( .A1(n11024), .A2(n11012), .B1(n11011), .B2(n11021), .ZN(
        P1_U3499) );
  OAI211_X1 U11594 ( .C1(n11016), .C2(n11015), .A(n11014), .B(n11013), .ZN(
        n11017) );
  AOI21_X1 U11595 ( .B1(n11019), .B2(n11018), .A(n11017), .ZN(n11023) );
  AOI22_X1 U11596 ( .A1(n11020), .A2(n11023), .B1(n7235), .B2(n5418), .ZN(
        P1_U3540) );
  INV_X1 U11597 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n11022) );
  AOI22_X1 U11598 ( .A1(n11024), .A2(n11023), .B1(n11022), .B2(n11021), .ZN(
        P1_U3505) );
  XNOR2_X1 U11599 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  AND2_X1 U6618 ( .A1(n5726), .A2(n5727), .ZN(n6261) );
  INV_X2 U5151 ( .A(n6248), .ZN(n6175) );
  CLKBUF_X1 U5172 ( .A(n10794), .Z(n5073) );
endmodule

