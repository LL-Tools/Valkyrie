

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, keyinput58, 
        keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, keyinput52, 
        keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, keyinput46, 
        keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, keyinput40, 
        keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, keyinput34, 
        keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, keyinput28, 
        keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, keyinput22, 
        keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, keyinput16, 
        keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, 
        keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, 
        keyinput3, keyinput2, keyinput1, keyinput0 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput63,
         keyinput62, keyinput61, keyinput60, keyinput59, keyinput58,
         keyinput57, keyinput56, keyinput55, keyinput54, keyinput53,
         keyinput52, keyinput51, keyinput50, keyinput49, keyinput48,
         keyinput47, keyinput46, keyinput45, keyinput44, keyinput43,
         keyinput42, keyinput41, keyinput40, keyinput39, keyinput38,
         keyinput37, keyinput36, keyinput35, keyinput34, keyinput33,
         keyinput32, keyinput31, keyinput30, keyinput29, keyinput28,
         keyinput27, keyinput26, keyinput25, keyinput24, keyinput23,
         keyinput22, keyinput21, keyinput20, keyinput19, keyinput18,
         keyinput17, keyinput16, keyinput15, keyinput14, keyinput13,
         keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, keyinput7,
         keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, keyinput1,
         keyinput0;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6433, n6436, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185;

  NAND2_X1 U7181 ( .A1(n10885), .A2(n10884), .ZN(n11936) );
  INV_X2 U7182 ( .A(n12153), .ZN(n12180) );
  BUF_X1 U7184 ( .A(n8753), .Z(n12346) );
  INV_X2 U7185 ( .A(n8130), .ZN(n8086) );
  INV_X2 U7186 ( .A(n11873), .ZN(n6911) );
  CLKBUF_X1 U7187 ( .A(n8748), .Z(n6452) );
  CLKBUF_X2 U7188 ( .A(n8756), .Z(n12333) );
  INV_X1 U7189 ( .A(n8186), .ZN(n8124) );
  INV_X1 U7190 ( .A(n12023), .ZN(n11627) );
  OR2_X1 U7191 ( .A1(n6440), .A2(n8730), .ZN(n8732) );
  AND2_X1 U7192 ( .A1(n11501), .A2(n8715), .ZN(n8753) );
  AND2_X1 U7194 ( .A1(n11887), .A2(n14741), .ZN(n12034) );
  INV_X1 U7195 ( .A(n8487), .ZN(n7582) );
  CLKBUF_X2 U7196 ( .A(n9600), .Z(n11872) );
  INV_X1 U7197 ( .A(n11816), .ZN(n11846) );
  NAND2_X2 U7198 ( .A1(n11680), .A2(n9354), .ZN(n11610) );
  CLKBUF_X1 U7199 ( .A(n9281), .Z(n6453) );
  NOR2_X1 U7200 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n6737) );
  CLKBUF_X1 U7201 ( .A(n13662), .Z(n6433) );
  NOR2_X1 U7202 ( .A1(n9706), .A2(n9707), .ZN(n13662) );
  NOR2_X1 U7203 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n6736) );
  AND2_X1 U7204 ( .A1(n6809), .A2(n6814), .ZN(n6806) );
  NOR2_X1 U7205 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n9211) );
  NOR2_X1 U7206 ( .A1(n9845), .A2(n9829), .ZN(n9915) );
  INV_X1 U7207 ( .A(n10514), .ZN(n10517) );
  NAND4_X1 U7208 ( .A1(n6737), .A2(n6736), .A3(n8591), .A4(n8942), .ZN(n8676)
         );
  INV_X2 U7209 ( .A(n10161), .ZN(n11775) );
  INV_X1 U7210 ( .A(n11680), .ZN(n11626) );
  AND3_X1 U7211 ( .A1(n13888), .A2(n13887), .A3(n14756), .ZN(n14114) );
  NAND2_X1 U7212 ( .A1(n9130), .A2(n10517), .ZN(n9834) );
  NAND2_X1 U7213 ( .A1(n7520), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7519) );
  AND4_X1 U7214 ( .A1(n6473), .A2(n6908), .A3(n6902), .A4(n6560), .ZN(n7458)
         );
  INV_X1 U7215 ( .A(n11818), .ZN(n11845) );
  NAND2_X1 U7216 ( .A1(n13903), .A2(n13886), .ZN(n13888) );
  OR2_X1 U7217 ( .A1(n12023), .A2(n7509), .ZN(n9597) );
  INV_X1 U7218 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n14216) );
  XNOR2_X1 U7219 ( .A(n8210), .B(n14264), .ZN(n8253) );
  AND3_X1 U7220 ( .A1(n8763), .A2(n8762), .A3(n8761), .ZN(n10595) );
  XNOR2_X1 U7221 ( .A(n10536), .B(n10550), .ZN(n14972) );
  NAND2_X1 U7222 ( .A1(n13271), .A2(n13270), .ZN(n13442) );
  NAND2_X1 U7223 ( .A1(n8010), .A2(n8009), .ZN(n13465) );
  NAND2_X1 U7224 ( .A1(n11700), .A2(n11699), .ZN(n14144) );
  NAND2_X1 U7225 ( .A1(n10845), .A2(n10844), .ZN(n11927) );
  NAND2_X1 U7226 ( .A1(n10139), .A2(n7190), .ZN(n11895) );
  INV_X2 U7227 ( .A(n11814), .ZN(n11839) );
  NOR2_X1 U7228 ( .A1(n13888), .A2(n14109), .ZN(n6968) );
  OAI211_X1 U7229 ( .C1(n11680), .C2(n9762), .A(n9761), .B(n9760), .ZN(n10695)
         );
  AND2_X1 U7230 ( .A1(n14392), .A2(n8286), .ZN(n8288) );
  INV_X1 U7231 ( .A(n9998), .ZN(n13226) );
  INV_X1 U7232 ( .A(n13700), .ZN(n9671) );
  INV_X1 U7233 ( .A(n9519), .ZN(n14370) );
  XNOR2_X1 U7234 ( .A(n9274), .B(n9244), .ZN(n9281) );
  NAND2_X2 U7235 ( .A1(n7290), .A2(n7291), .ZN(n10312) );
  NOR2_X4 U7236 ( .A1(n9209), .A2(n9285), .ZN(n7291) );
  NAND2_X2 U7241 ( .A1(n6489), .A2(n8755), .ZN(n12556) );
  OR4_X2 U7242 ( .A1(n13276), .A2(n13347), .A3(n13328), .A4(n8568), .ZN(n8569)
         );
  AND2_X2 U7243 ( .A1(n13347), .A2(n6504), .ZN(n7231) );
  XNOR2_X2 U7244 ( .A(n13472), .B(n12987), .ZN(n13347) );
  XNOR2_X2 U7245 ( .A(n8638), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8911) );
  NAND2_X2 U7246 ( .A1(n8637), .A2(n8636), .ZN(n8638) );
  OR4_X2 U7247 ( .A1(n13858), .A2(n13992), .A3(n13850), .A4(n12055), .ZN(
        n12056) );
  XNOR2_X2 U7248 ( .A(n14149), .B(n13851), .ZN(n13850) );
  BUF_X8 U7249 ( .A(n8340), .Z(n8541) );
  INV_X2 U7250 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n6720) );
  XNOR2_X2 U7251 ( .A(n13095), .B(n8319), .ZN(n9630) );
  NAND4_X2 U7252 ( .A1(n7555), .A2(n7554), .A3(n7553), .A4(n7552), .ZN(n13095)
         );
  NAND2_X2 U7253 ( .A1(n8686), .A2(n8685), .ZN(n12670) );
  AND2_X2 U7255 ( .A1(n14950), .A2(n10535), .ZN(n10536) );
  NAND2_X1 U7256 ( .A1(n9130), .A2(n10517), .ZN(n6438) );
  NAND2_X1 U7257 ( .A1(n9130), .A2(n10517), .ZN(n6439) );
  XOR2_X2 U7258 ( .A(n8269), .B(n8268), .Z(n15172) );
  AND2_X2 U7259 ( .A1(n7116), .A2(n6559), .ZN(n8210) );
  NOR2_X2 U7260 ( .A1(n15009), .A2(n15010), .ZN(n15008) );
  XNOR2_X2 U7261 ( .A(n12564), .B(n15014), .ZN(n15009) );
  AOI21_X2 U7262 ( .B1(n8547), .B2(n8546), .A(n8545), .ZN(n8552) );
  XOR2_X2 U7263 ( .A(n8260), .B(n8259), .Z(n8262) );
  NAND2_X1 U7264 ( .A1(n11501), .A2(n12935), .ZN(n6440) );
  BUF_X4 U7265 ( .A(n8749), .Z(n6445) );
  NOR2_X2 U7266 ( .A1(n10952), .A2(n8806), .ZN(n10953) );
  XNOR2_X2 U7267 ( .A(n6884), .B(n10963), .ZN(n10952) );
  NOR2_X2 U7268 ( .A1(n8207), .A2(n8208), .ZN(n8209) );
  XOR2_X2 U7269 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n8254), .Z(n8255) );
  OAI21_X2 U7270 ( .B1(n8259), .B2(n8260), .A(n6551), .ZN(n7126) );
  XNOR2_X2 U7271 ( .A(n6720), .B(P1_ADDR_REG_1__SCAN_IN), .ZN(n8259) );
  XNOR2_X2 U7272 ( .A(n7519), .B(P2_IR_REG_29__SCAN_IN), .ZN(n7522) );
  OAI21_X2 U7273 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n8265), .A(n14382), .ZN(
        n15181) );
  XNOR2_X1 U7274 ( .A(n8471), .B(n8470), .ZN(n11850) );
  NAND2_X1 U7275 ( .A1(n7096), .A2(n7097), .ZN(n12155) );
  INV_X1 U7276 ( .A(n13969), .ZN(n6441) );
  AOI21_X1 U7277 ( .B1(n13653), .B2(n13654), .A(n6537), .ZN(n13588) );
  NAND2_X1 U7278 ( .A1(n7067), .A2(n7064), .ZN(n12467) );
  CLKBUF_X1 U7279 ( .A(n11473), .Z(n6721) );
  NOR2_X1 U7280 ( .A1(n8290), .A2(n8289), .ZN(n14565) );
  OAI21_X1 U7281 ( .B1(n10319), .B2(n10318), .A(n10317), .ZN(n10330) );
  NAND2_X1 U7282 ( .A1(n10392), .A2(n10391), .ZN(n10395) );
  INV_X1 U7283 ( .A(n13933), .ZN(n13900) );
  NAND2_X1 U7284 ( .A1(n7747), .A2(n7746), .ZN(n12126) );
  OR2_X1 U7285 ( .A1(n10843), .A2(n7908), .ZN(n7730) );
  INV_X1 U7286 ( .A(n14734), .ZN(n14785) );
  NAND2_X1 U7287 ( .A1(n7636), .A2(n7635), .ZN(n10274) );
  NOR2_X1 U7288 ( .A1(n6442), .A2(n10643), .ZN(n14697) );
  OAI21_X1 U7289 ( .B1(n15175), .B2(n15176), .A(n7115), .ZN(n7114) );
  NAND2_X1 U7290 ( .A1(n10687), .A2(n14753), .ZN(n11891) );
  INV_X1 U7291 ( .A(n14753), .ZN(n14773) );
  XNOR2_X1 U7292 ( .A(n9983), .B(n10006), .ZN(n9721) );
  INV_X2 U7293 ( .A(n13094), .ZN(n9983) );
  INV_X1 U7294 ( .A(n14723), .ZN(n13697) );
  INV_X1 U7295 ( .A(n13696), .ZN(n10793) );
  AND4_X1 U7296 ( .A1(n8783), .A2(n8782), .A3(n8781), .A4(n8780), .ZN(n10834)
         );
  CLKBUF_X1 U7297 ( .A(n7610), .Z(n7908) );
  AND2_X1 U7298 ( .A1(n7523), .A2(n13546), .ZN(n7570) );
  INV_X2 U7299 ( .A(n7610), .ZN(n8509) );
  CLKBUF_X2 U7300 ( .A(n8729), .Z(n12350) );
  INV_X2 U7301 ( .A(n7771), .ZN(n9428) );
  OAI211_X1 U7302 ( .C1(n8146), .C2(n7505), .A(n7504), .B(n7503), .ZN(n13548)
         );
  AND3_X1 U7303 ( .A1(n7468), .A2(n7163), .A3(n7679), .ZN(n7478) );
  NOR2_X1 U7305 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n7041) );
  NOR2_X1 U7306 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n7040) );
  INV_X1 U7307 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10137) );
  AND2_X1 U7308 ( .A1(n14116), .A2(n6695), .ZN(n6694) );
  MUX2_X1 U7309 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n12827), .S(n15166), .Z(
        n12828) );
  MUX2_X1 U7310 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n12827), .S(n15158), .Z(
        n12088) );
  NOR2_X1 U7311 ( .A1(n7388), .A2(n7386), .ZN(n7385) );
  AOI21_X1 U7312 ( .B1(n13554), .B2(n13555), .A(n6536), .ZN(n11813) );
  AND2_X1 U7313 ( .A1(n11516), .A2(n11515), .ZN(n12087) );
  AOI21_X1 U7314 ( .B1(n7315), .B2(n14685), .A(n7312), .ZN(n14117) );
  MUX2_X1 U7315 ( .A(P3_REG1_REG_29__SCAN_IN), .B(n9203), .S(n15166), .Z(n9204) );
  MUX2_X1 U7316 ( .A(P3_REG0_REG_29__SCAN_IN), .B(n9203), .S(n15158), .Z(n9200) );
  NAND2_X1 U7317 ( .A1(n6616), .A2(n11779), .ZN(n13554) );
  NOR2_X1 U7318 ( .A1(n13902), .A2(n13901), .ZN(n6804) );
  NAND2_X1 U7319 ( .A1(n6773), .A2(n8525), .ZN(n8530) );
  NAND2_X1 U7320 ( .A1(n7075), .A2(n7074), .ZN(n12510) );
  NAND2_X1 U7321 ( .A1(n12995), .A2(n12994), .ZN(n8080) );
  AND2_X1 U7322 ( .A1(n7335), .A2(n7338), .ZN(n13435) );
  NAND2_X1 U7323 ( .A1(n12345), .A2(n12344), .ZN(n12878) );
  AND2_X1 U7324 ( .A1(n6654), .A2(n6656), .ZN(n6653) );
  NAND2_X1 U7325 ( .A1(n8512), .A2(n8511), .ZN(n13427) );
  INV_X1 U7326 ( .A(n14103), .ZN(n13812) );
  AND2_X1 U7327 ( .A1(n6628), .A2(n11559), .ZN(n13271) );
  OR2_X1 U7328 ( .A1(n13275), .A2(n11557), .ZN(n6628) );
  AOI21_X1 U7329 ( .B1(n12491), .B2(n12747), .A(n12157), .ZN(n12160) );
  NOR2_X1 U7330 ( .A1(n12057), .A2(n13837), .ZN(n6907) );
  NAND2_X1 U7331 ( .A1(n6807), .A2(n6806), .ZN(n13935) );
  OAI211_X1 U7332 ( .C1(n8508), .C2(n8507), .A(n8506), .B(n8505), .ZN(n14222)
         );
  AND2_X1 U7333 ( .A1(n6610), .A2(n11714), .ZN(n6609) );
  AND2_X1 U7334 ( .A1(n7186), .A2(n6810), .ZN(n6809) );
  NAND2_X1 U7335 ( .A1(n8489), .A2(n8488), .ZN(n13434) );
  OAI21_X1 U7336 ( .B1(n11552), .B2(n7219), .A(n7217), .ZN(n6629) );
  NAND2_X1 U7337 ( .A1(n6776), .A2(n6775), .ZN(n8506) );
  XNOR2_X1 U7338 ( .A(n12155), .B(n12154), .ZN(n12491) );
  OR2_X1 U7339 ( .A1(n13320), .A2(n11550), .ZN(n11552) );
  OR2_X1 U7340 ( .A1(n14378), .A2(n14379), .ZN(n7120) );
  NAND2_X1 U7341 ( .A1(n6441), .A2(n13957), .ZN(n13953) );
  NAND2_X1 U7342 ( .A1(n11795), .A2(n11794), .ZN(n14115) );
  NAND2_X1 U7343 ( .A1(n13586), .A2(n11646), .ZN(n13636) );
  OR3_X1 U7344 ( .A1(n8411), .A2(n7383), .A3(n8414), .ZN(n7381) );
  XNOR2_X1 U7345 ( .A(n8486), .B(n8485), .ZN(n13544) );
  NAND2_X1 U7346 ( .A1(n8486), .A2(n8485), .ZN(n8504) );
  NAND2_X1 U7347 ( .A1(n8466), .A2(n8465), .ZN(n8486) );
  NAND2_X1 U7348 ( .A1(n6633), .A2(n6498), .ZN(n11548) );
  NAND2_X1 U7349 ( .A1(n13588), .A2(n13587), .ZN(n13586) );
  OAI21_X1 U7350 ( .B1(n6677), .B2(n6676), .A(n13020), .ZN(n12985) );
  NAND2_X1 U7351 ( .A1(n13356), .A2(n13355), .ZN(n13354) );
  NAND2_X1 U7352 ( .A1(n7170), .A2(n6464), .ZN(n14159) );
  OR2_X1 U7353 ( .A1(n8177), .A2(n8176), .ZN(n8466) );
  NAND2_X1 U7354 ( .A1(n14013), .A2(n13822), .ZN(n13993) );
  NAND2_X1 U7355 ( .A1(n6634), .A2(n11546), .ZN(n13375) );
  XNOR2_X1 U7356 ( .A(n8106), .B(n8168), .ZN(n13547) );
  OR2_X1 U7357 ( .A1(n14044), .A2(n7173), .ZN(n7170) );
  INV_X1 U7358 ( .A(n13282), .ZN(n13451) );
  NAND2_X1 U7359 ( .A1(n11762), .A2(n11761), .ZN(n14126) );
  XNOR2_X1 U7360 ( .A(n8008), .B(n8007), .ZN(n11697) );
  NAND2_X1 U7361 ( .A1(n14574), .A2(n14572), .ZN(n14579) );
  OR2_X1 U7362 ( .A1(n13419), .A2(n13420), .ZN(n13417) );
  AND2_X2 U7363 ( .A1(n11650), .A2(n11649), .ZN(n14161) );
  NAND2_X1 U7364 ( .A1(n7950), .A2(n7949), .ZN(n13481) );
  NOR2_X2 U7365 ( .A1(n14027), .A2(n14045), .ZN(n14030) );
  OR2_X1 U7366 ( .A1(n14027), .A2(n14054), .ZN(n11975) );
  NAND2_X1 U7367 ( .A1(n11740), .A2(n11739), .ZN(n14133) );
  XNOR2_X1 U7368 ( .A(n8102), .B(n8100), .ZN(n11759) );
  NAND2_X1 U7369 ( .A1(n11629), .A2(n11628), .ZN(n14027) );
  XNOR2_X1 U7370 ( .A(n8103), .B(SI_26_), .ZN(n8102) );
  NOR2_X1 U7371 ( .A1(n7275), .A2(n13612), .ZN(n7274) );
  AND2_X1 U7372 ( .A1(n7201), .A2(n7200), .ZN(n11211) );
  NAND2_X1 U7373 ( .A1(n8040), .A2(n8039), .ZN(n13462) );
  NAND2_X1 U7374 ( .A1(n7279), .A2(n6461), .ZN(n11452) );
  OAI21_X1 U7375 ( .B1(n8082), .B2(n8081), .A(n8083), .ZN(n8103) );
  XNOR2_X1 U7376 ( .A(n7948), .B(n7947), .ZN(n11647) );
  AOI21_X1 U7377 ( .B1(n7278), .B2(n13563), .A(n6555), .ZN(n7277) );
  NAND2_X1 U7378 ( .A1(n11613), .A2(n11612), .ZN(n14174) );
  NAND2_X1 U7379 ( .A1(n7252), .A2(n7251), .ZN(n7946) );
  NAND2_X1 U7380 ( .A1(n7911), .A2(n7910), .ZN(n13493) );
  AND2_X1 U7381 ( .A1(n7927), .A2(n7945), .ZN(n7252) );
  NAND2_X1 U7382 ( .A1(n6759), .A2(n7968), .ZN(n8025) );
  AOI21_X1 U7383 ( .B1(n7207), .B2(n7205), .A(n7204), .ZN(n7203) );
  OR2_X1 U7384 ( .A1(n15062), .A2(n15061), .ZN(n15059) );
  AND2_X1 U7385 ( .A1(n7109), .A2(n14560), .ZN(n8290) );
  NAND2_X1 U7386 ( .A1(n7716), .A2(n10202), .ZN(n10208) );
  OAI21_X1 U7387 ( .B1(n14562), .B2(n14561), .A(n7110), .ZN(n7109) );
  NAND3_X1 U7388 ( .A1(n7925), .A2(n7262), .A3(n7261), .ZN(n7926) );
  AND2_X1 U7389 ( .A1(n7925), .A2(n6590), .ZN(n6764) );
  NAND2_X1 U7390 ( .A1(n6627), .A2(SI_18_), .ZN(n7925) );
  AOI21_X1 U7391 ( .B1(n7361), .B2(n7359), .A(n6542), .ZN(n7358) );
  AND2_X1 U7392 ( .A1(n6997), .A2(n6994), .ZN(n15043) );
  NAND2_X1 U7393 ( .A1(n8652), .A2(n8651), .ZN(n8991) );
  NAND2_X1 U7394 ( .A1(n8945), .A2(n8944), .ZN(n12925) );
  AOI21_X1 U7395 ( .B1(n7309), .B2(n7307), .A(n6541), .ZN(n7306) );
  AND2_X1 U7396 ( .A1(n15024), .A2(n12567), .ZN(n12568) );
  NAND2_X1 U7397 ( .A1(n7821), .A2(n7820), .ZN(n14508) );
  NAND2_X1 U7398 ( .A1(n14397), .A2(n14395), .ZN(n14558) );
  NAND2_X1 U7399 ( .A1(n11283), .A2(n11282), .ZN(n14194) );
  NAND2_X1 U7400 ( .A1(n11054), .A2(n11053), .ZN(n11179) );
  NAND2_X1 U7401 ( .A1(n10023), .A2(n10022), .ZN(n10291) );
  NAND2_X1 U7402 ( .A1(n6625), .A2(n7876), .ZN(n7899) );
  NAND2_X1 U7403 ( .A1(n11092), .A2(n12237), .ZN(n11065) );
  AND2_X1 U7404 ( .A1(n10427), .A2(n8556), .ZN(n10396) );
  NAND2_X1 U7405 ( .A1(n7795), .A2(n7794), .ZN(n7817) );
  OAI21_X1 U7406 ( .B1(n7795), .B2(n7241), .A(n7239), .ZN(n7853) );
  XNOR2_X1 U7407 ( .A(n7763), .B(n7762), .ZN(n10883) );
  NAND2_X1 U7408 ( .A1(n6624), .A2(n6623), .ZN(n7874) );
  OAI21_X1 U7409 ( .B1(n9928), .B2(n9927), .A(n9929), .ZN(n9931) );
  NAND2_X1 U7410 ( .A1(n7685), .A2(n7684), .ZN(n12975) );
  NAND2_X1 U7411 ( .A1(n10728), .A2(n10727), .ZN(n11923) );
  NAND2_X1 U7412 ( .A1(n8640), .A2(n8639), .ZN(n8926) );
  NAND2_X1 U7413 ( .A1(n7790), .A2(n7789), .ZN(n7797) );
  NAND2_X1 U7414 ( .A1(n9790), .A2(n9789), .ZN(n9928) );
  NAND2_X1 U7415 ( .A1(n7660), .A2(n7659), .ZN(n10289) );
  NAND2_X1 U7416 ( .A1(n7722), .A2(n7721), .ZN(n7725) );
  NAND2_X1 U7417 ( .A1(n10443), .A2(n10442), .ZN(n10441) );
  OAI21_X1 U7418 ( .B1(n7673), .B2(n7675), .A(n6768), .ZN(n7704) );
  NAND2_X1 U7419 ( .A1(n10302), .A2(n9100), .ZN(n10443) );
  NAND2_X1 U7420 ( .A1(n8908), .A2(n8634), .ZN(n8637) );
  OAI21_X1 U7421 ( .B1(n14723), .B2(n11895), .A(n14725), .ZN(n12036) );
  AND2_X2 U7422 ( .A1(n10003), .A2(n13377), .ZN(n13426) );
  AOI21_X1 U7423 ( .B1(n15118), .B2(n12200), .A(n6486), .ZN(n10304) );
  INV_X2 U7424 ( .A(n14691), .ZN(n6442) );
  INV_X2 U7425 ( .A(n14928), .ZN(n6443) );
  AND2_X1 U7426 ( .A1(n12216), .A2(n12215), .ZN(n12358) );
  NAND2_X1 U7427 ( .A1(n10591), .A2(n12816), .ZN(n12818) );
  NAND2_X1 U7428 ( .A1(n7589), .A2(n7588), .ZN(n10073) );
  INV_X1 U7429 ( .A(n8845), .ZN(n8631) );
  AND2_X1 U7430 ( .A1(n8867), .A2(n8628), .ZN(n8845) );
  NAND2_X1 U7431 ( .A1(n15170), .A2(n8270), .ZN(n8275) );
  OR2_X1 U7432 ( .A1(n8865), .A2(n8864), .ZN(n8867) );
  AND3_X1 U7433 ( .A1(n8821), .A2(n8820), .A3(n8819), .ZN(n10924) );
  AND4_X1 U7434 ( .A1(n8813), .A2(n8812), .A3(n8811), .A4(n8810), .ZN(n11081)
         );
  AND4_X1 U7435 ( .A1(n8769), .A2(n8768), .A3(n8767), .A4(n8766), .ZN(n10710)
         );
  NAND2_X1 U7436 ( .A1(n6873), .A2(n6986), .ZN(n14949) );
  NAND4_X1 U7437 ( .A1(n7530), .A2(n7529), .A3(n7531), .A4(n7532), .ZN(n9465)
         );
  AND3_X1 U7438 ( .A1(n8777), .A2(n8776), .A3(n8775), .ZN(n10494) );
  AND3_X1 U7439 ( .A1(n8793), .A2(n8792), .A3(n8791), .ZN(n10712) );
  OAI21_X1 U7440 ( .B1(n9395), .B2(P3_D_REG_0__SCAN_IN), .A(n9422), .ZN(n10040) );
  NAND2_X1 U7441 ( .A1(n9231), .A2(n11334), .ZN(n10182) );
  OR2_X2 U7442 ( .A1(n11867), .A2(n11843), .ZN(n14090) );
  AND2_X1 U7443 ( .A1(n7633), .A2(n6774), .ZN(n6724) );
  AND2_X2 U7444 ( .A1(n12415), .A2(n12195), .ZN(n12327) );
  INV_X2 U7445 ( .A(n8753), .ZN(n9127) );
  OAI21_X1 U7446 ( .B1(n8803), .B2(n7028), .A(n7026), .ZN(n8835) );
  AND2_X1 U7447 ( .A1(n13546), .A2(n11576), .ZN(n7571) );
  NAND2_X2 U7448 ( .A1(n7166), .A2(n7165), .ZN(n8050) );
  INV_X1 U7449 ( .A(n7523), .ZN(n11576) );
  INV_X2 U7450 ( .A(n8729), .ZN(n9188) );
  OR2_X1 U7451 ( .A1(n6901), .A2(n7607), .ZN(n6774) );
  NAND2_X1 U7452 ( .A1(n8620), .A2(n8619), .ZN(n8803) );
  NAND2_X1 U7453 ( .A1(n6989), .A2(n6988), .ZN(n6987) );
  XNOR2_X1 U7454 ( .A(n7235), .B(P2_IR_REG_30__SCAN_IN), .ZN(n7523) );
  NAND2_X1 U7455 ( .A1(n8157), .A2(n7474), .ZN(n11264) );
  NAND2_X1 U7456 ( .A1(n13539), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7235) );
  OAI21_X1 U7457 ( .B1(n8758), .B2(n7015), .A(n7013), .ZN(n8785) );
  NAND2_X1 U7458 ( .A1(n7472), .A2(n7471), .ZN(n8157) );
  MUX2_X1 U7459 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7473), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n7474) );
  NAND2_X1 U7460 ( .A1(n9265), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9266) );
  NAND2_X1 U7461 ( .A1(n6647), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9249) );
  NAND2_X1 U7462 ( .A1(n9273), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9274) );
  XNOR2_X1 U7463 ( .A(n8713), .B(P3_IR_REG_29__SCAN_IN), .ZN(n8715) );
  NAND2_X1 U7464 ( .A1(n14217), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9248) );
  NAND2_X1 U7465 ( .A1(n7499), .A2(n7452), .ZN(n8146) );
  INV_X1 U7466 ( .A(n7476), .ZN(n7472) );
  NAND2_X1 U7467 ( .A1(n7483), .A2(n6650), .ZN(n11102) );
  AND2_X1 U7468 ( .A1(n7567), .A2(n7584), .ZN(n13110) );
  AND3_X1 U7469 ( .A1(n7477), .A2(n6576), .A3(n7476), .ZN(n7517) );
  NAND2_X1 U7470 ( .A1(n6741), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6740) );
  XNOR2_X1 U7471 ( .A(n9496), .B(P1_IR_REG_19__SCAN_IN), .ZN(n12058) );
  NOR2_X1 U7472 ( .A1(n9495), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n9261) );
  NAND2_X2 U7473 ( .A1(n6450), .A2(P2_U3088), .ZN(n13549) );
  AND2_X1 U7474 ( .A1(n8617), .A2(n7017), .ZN(n7016) );
  AND2_X1 U7475 ( .A1(n7442), .A2(n7063), .ZN(n7062) );
  AND4_X1 U7476 ( .A1(n7494), .A2(n7493), .A3(n7492), .A4(n8158), .ZN(n7452)
         );
  NAND2_X1 U7477 ( .A1(n8739), .A2(n8738), .ZN(n9844) );
  CLKBUF_X2 U7478 ( .A(n7563), .Z(n6448) );
  AND2_X1 U7479 ( .A1(n6491), .A2(n8681), .ZN(n7442) );
  AND4_X1 U7480 ( .A1(n8586), .A2(n8585), .A3(n8830), .A4(n8817), .ZN(n8587)
         );
  AND4_X2 U7481 ( .A1(n7041), .A2(n7040), .A3(n7428), .A4(n7039), .ZN(n8786)
         );
  NOR2_X1 U7482 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n9212) );
  INV_X1 U7483 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9243) );
  INV_X1 U7484 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9218) );
  NOR2_X1 U7485 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n9208) );
  INV_X4 U7486 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7487 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9291) );
  INV_X1 U7488 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8830) );
  NOR2_X1 U7489 ( .A1(P3_IR_REG_26__SCAN_IN), .A2(P3_IR_REG_25__SCAN_IN), .ZN(
        n7063) );
  INV_X4 U7490 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X1 U7491 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n7856) );
  NOR2_X1 U7492 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n7464) );
  INV_X4 U7493 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7494 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n7471) );
  INV_X1 U7495 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8942) );
  INV_X1 U7496 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8591) );
  INV_X1 U7497 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8588) );
  NOR2_X1 U7498 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8585) );
  OAI21_X1 U7499 ( .B1(n14579), .B2(n14578), .A(n7112), .ZN(n6730) );
  OAI21_X2 U7500 ( .B1(n6479), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8590) );
  XNOR2_X1 U7501 ( .A(n12966), .B(n13087), .ZN(n10429) );
  NAND2_X1 U7502 ( .A1(n9281), .A2(n11492), .ZN(n6444) );
  NAND2_X2 U7503 ( .A1(n9281), .A2(n11492), .ZN(n11680) );
  NAND2_X2 U7504 ( .A1(n12557), .A2(n10052), .ZN(n12196) );
  INV_X2 U7505 ( .A(n6448), .ZN(n9354) );
  OAI21_X1 U7506 ( .B1(n8712), .B2(P3_IR_REG_28__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8713) );
  OAI222_X1 U7507 ( .A1(P3_U3151), .A2(n11501), .B1(n11500), .B2(n11499), .C1(
        n12332), .C2(n12939), .ZN(P3_U3265) );
  NOR2_X2 U7508 ( .A1(n15078), .A2(n12626), .ZN(n15077) );
  AOI21_X2 U7509 ( .B1(n13369), .B2(n13376), .A(n11529), .ZN(n13356) );
  OAI21_X2 U7510 ( .B1(n13391), .B2(n13392), .A(n11528), .ZN(n13369) );
  XNOR2_X2 U7511 ( .A(n14693), .B(n14703), .ZN(n14686) );
  NAND2_X2 U7512 ( .A1(n9293), .A2(n9206), .ZN(n9285) );
  NOR2_X4 U7513 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9293) );
  AOI211_X2 U7514 ( .C1(n13513), .C2(n13451), .A(n13450), .B(n13449), .ZN(
        n13452) );
  INV_X1 U7515 ( .A(n9097), .ZN(n12557) );
  NAND2_X1 U7518 ( .A1(n8749), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8721) );
  INV_X1 U7519 ( .A(n8731), .ZN(n8749) );
  AND2_X1 U7520 ( .A1(n11576), .A2(n7522), .ZN(n6446) );
  AND2_X1 U7521 ( .A1(n11576), .A2(n7522), .ZN(n6447) );
  NAND2_X2 U7522 ( .A1(n12196), .A2(n12191), .ZN(n10043) );
  INV_X4 U7523 ( .A(n8344), .ZN(n8340) );
  XNOR2_X2 U7524 ( .A(n7498), .B(n7518), .ZN(n8192) );
  OAI21_X2 U7525 ( .B1(n10831), .B2(n7402), .A(n7399), .ZN(n11093) );
  NAND2_X2 U7526 ( .A1(n10833), .A2(n10832), .ZN(n10831) );
  AND2_X1 U7527 ( .A1(n7522), .A2(n7523), .ZN(n7591) );
  NAND2_X2 U7528 ( .A1(n12768), .A2(n12774), .ZN(n12767) );
  AOI21_X2 U7529 ( .B1(n12914), .B2(n12800), .A(n12781), .ZN(n12768) );
  NOR2_X2 U7530 ( .A1(n12782), .A2(n12783), .ZN(n12781) );
  NOR2_X2 U7531 ( .A1(n6958), .A2(n14693), .ZN(n14688) );
  NAND2_X2 U7532 ( .A1(n14736), .A2(n6954), .ZN(n6958) );
  OAI22_X2 U7533 ( .A1(n12796), .A2(n12801), .B1(n12812), .B2(n12918), .ZN(
        n12782) );
  AOI21_X2 U7534 ( .B1(n11439), .B2(n6503), .A(n7433), .ZN(n12796) );
  BUF_X4 U7535 ( .A(n7563), .Z(n6450) );
  AND2_X2 U7536 ( .A1(n7260), .A2(n7259), .ZN(n7563) );
  INV_X2 U7537 ( .A(n10602), .ZN(n10052) );
  OAI211_X2 U7538 ( .C1(n8888), .C2(n9347), .A(n7427), .B(n7426), .ZN(n10602)
         );
  OAI222_X1 U7539 ( .A1(P3_U3151), .A2(n9130), .B1(n11500), .B2(n12941), .C1(
        n12940), .C2(n12939), .ZN(P3_U3267) );
  NAND2_X1 U7540 ( .A1(n8714), .A2(n8715), .ZN(n8748) );
  INV_X2 U7541 ( .A(n12026), .ZN(n6454) );
  NAND2_X1 U7543 ( .A1(n9671), .A2(n11876), .ZN(n11879) );
  OAI22_X4 U7544 ( .A1(n11376), .A2(n12372), .B1(n14482), .B2(n11441), .ZN(
        n11439) );
  AOI22_X2 U7545 ( .A1(n11217), .A2(n12370), .B1(n12548), .B2(n14487), .ZN(
        n11376) );
  NAND2_X1 U7546 ( .A1(n8530), .A2(n8517), .ZN(n8524) );
  AND2_X1 U7547 ( .A1(n7245), .A2(n6916), .ZN(n6915) );
  OR2_X1 U7548 ( .A1(n7703), .A2(n6917), .ZN(n6916) );
  OAI21_X1 U7549 ( .B1(n12654), .B2(n12195), .A(n10196), .ZN(n10042) );
  NAND2_X1 U7550 ( .A1(n9924), .A2(n9923), .ZN(n9926) );
  AND2_X1 U7551 ( .A1(n14039), .A2(n7175), .ZN(n7174) );
  NAND2_X1 U7552 ( .A1(n13847), .A2(n13846), .ZN(n7175) );
  OR2_X1 U7553 ( .A1(n13686), .A2(n14085), .ZN(n11954) );
  NAND2_X1 U7554 ( .A1(n6438), .A2(n6450), .ZN(n8756) );
  AND2_X1 U7555 ( .A1(n11562), .A2(n8553), .ZN(n13249) );
  NAND2_X1 U7556 ( .A1(n7478), .A2(n7470), .ZN(n7476) );
  INV_X1 U7557 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7470) );
  CLKBUF_X1 U7558 ( .A(n10328), .Z(n11808) );
  NAND3_X1 U7559 ( .A1(n7168), .A2(n6535), .A3(n7167), .ZN(n6789) );
  NAND2_X1 U7560 ( .A1(n6789), .A2(n6788), .ZN(n11024) );
  AND2_X1 U7561 ( .A1(n12045), .A2(n6790), .ZN(n6788) );
  AND2_X1 U7562 ( .A1(n10420), .A2(n9999), .ZN(n8308) );
  INV_X1 U7563 ( .A(n11897), .ZN(n6947) );
  AND2_X1 U7564 ( .A1(n6824), .A2(n6823), .ZN(n8333) );
  NAND2_X1 U7565 ( .A1(n13094), .A2(n8344), .ZN(n6824) );
  NAND2_X1 U7566 ( .A1(n10006), .A2(n8340), .ZN(n6823) );
  NAND2_X1 U7567 ( .A1(n11985), .A2(n11987), .ZN(n6939) );
  XNOR2_X1 U7568 ( .A(n13427), .B(n13231), .ZN(n8525) );
  NAND2_X1 U7569 ( .A1(n6912), .A2(n6910), .ZN(n12068) );
  NAND2_X1 U7570 ( .A1(n12064), .A2(n12026), .ZN(n6910) );
  NAND2_X1 U7571 ( .A1(n12063), .A2(n6454), .ZN(n6912) );
  OR2_X1 U7572 ( .A1(n14194), .A2(n11585), .ZN(n11951) );
  NAND2_X1 U7573 ( .A1(n8105), .A2(n8104), .ZN(n8170) );
  NAND2_X1 U7574 ( .A1(n8102), .A2(n8101), .ZN(n8105) );
  OR2_X1 U7575 ( .A1(n10040), .A2(n12392), .ZN(n10041) );
  INV_X1 U7576 ( .A(n6755), .ZN(n6754) );
  AOI21_X1 U7577 ( .B1(n6756), .B2(n6478), .A(n12636), .ZN(n6755) );
  OR2_X1 U7578 ( .A1(n12170), .A2(n12676), .ZN(n9095) );
  NOR2_X1 U7579 ( .A1(n12705), .A2(n6854), .ZN(n6853) );
  INV_X1 U7580 ( .A(n12312), .ZN(n6854) );
  OR2_X1 U7581 ( .A1(n12736), .A2(n12747), .ZN(n12302) );
  OR2_X1 U7582 ( .A1(n12750), .A2(n12758), .ZN(n12295) );
  OR2_X1 U7583 ( .A1(n12482), .A2(n12746), .ZN(n12292) );
  OR2_X1 U7584 ( .A1(n12439), .A2(n12785), .ZN(n12288) );
  NAND2_X1 U7585 ( .A1(n8663), .A2(n8662), .ZN(n8664) );
  NAND2_X1 U7586 ( .A1(n9037), .A2(n9036), .ZN(n8663) );
  OR2_X1 U7587 ( .A1(n8119), .A2(n8118), .ZN(n7143) );
  OR2_X1 U7588 ( .A1(n12943), .A2(n7145), .ZN(n7144) );
  NAND2_X1 U7589 ( .A1(n7149), .A2(n8099), .ZN(n7145) );
  INV_X1 U7590 ( .A(n8524), .ZN(n6772) );
  OAI21_X1 U7591 ( .B1(n6484), .B2(n7219), .A(n11555), .ZN(n7218) );
  INV_X1 U7592 ( .A(n11102), .ZN(n9462) );
  INV_X1 U7593 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8141) );
  NAND2_X1 U7594 ( .A1(n11352), .A2(n13814), .ZN(n7298) );
  AND2_X1 U7595 ( .A1(n6795), .A2(n6485), .ZN(n6793) );
  NAND2_X1 U7596 ( .A1(n14027), .A2(n14054), .ZN(n13821) );
  NAND2_X1 U7597 ( .A1(n6642), .A2(n6641), .ZN(n6640) );
  INV_X1 U7598 ( .A(n14039), .ZN(n6641) );
  INV_X1 U7599 ( .A(n14038), .ZN(n6642) );
  NAND2_X1 U7600 ( .A1(n14544), .A2(n11947), .ZN(n7185) );
  INV_X1 U7601 ( .A(n10312), .ZN(n9247) );
  AOI21_X1 U7602 ( .B1(n7237), .B2(n7240), .A(n6550), .ZN(n6623) );
  NAND2_X1 U7603 ( .A1(n7797), .A2(n7237), .ZN(n6624) );
  XNOR2_X1 U7604 ( .A(n7875), .B(SI_16_), .ZN(n7873) );
  AOI21_X1 U7605 ( .B1(n7245), .B2(n7247), .A(n7244), .ZN(n7243) );
  INV_X1 U7606 ( .A(n7786), .ZN(n7244) );
  AND2_X1 U7607 ( .A1(n6915), .A2(n6767), .ZN(n6766) );
  NAND2_X1 U7608 ( .A1(n6768), .A2(n7675), .ZN(n6767) );
  XNOR2_X1 U7609 ( .A(n7788), .B(SI_12_), .ZN(n7786) );
  NAND2_X1 U7610 ( .A1(n6630), .A2(SI_10_), .ZN(n7741) );
  NOR2_X1 U7611 ( .A1(n9388), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n10211) );
  NAND2_X1 U7612 ( .A1(n8216), .A2(n8215), .ZN(n8279) );
  OR2_X1 U7613 ( .A1(n8277), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n8215) );
  OR2_X1 U7614 ( .A1(n8946), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8959) );
  NAND2_X1 U7615 ( .A1(n11420), .A2(n11419), .ZN(n11473) );
  AOI21_X1 U7616 ( .B1(n6455), .B2(n12483), .A(n6514), .ZN(n7097) );
  NAND2_X1 U7617 ( .A1(n12313), .A2(n12680), .ZN(n12689) );
  INV_X1 U7618 ( .A(n12689), .ZN(n12696) );
  OR2_X1 U7619 ( .A1(n12725), .A2(n12733), .ZN(n12312) );
  NOR2_X1 U7620 ( .A1(n7049), .A2(n8923), .ZN(n7048) );
  OR2_X1 U7621 ( .A1(n8855), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8896) );
  NAND2_X1 U7622 ( .A1(n9166), .A2(n12406), .ZN(n12766) );
  OR2_X1 U7623 ( .A1(n9834), .A2(n9844), .ZN(n7426) );
  INV_X1 U7624 ( .A(n10196), .ZN(n9165) );
  INV_X1 U7625 ( .A(n12654), .ZN(n12404) );
  NAND2_X2 U7626 ( .A1(n6439), .A2(n9354), .ZN(n8888) );
  INV_X1 U7627 ( .A(n8888), .ZN(n12343) );
  XNOR2_X1 U7628 ( .A(n9142), .B(P3_IR_REG_26__SCAN_IN), .ZN(n9159) );
  AND2_X1 U7629 ( .A1(n8601), .A2(n9160), .ZN(n12195) );
  NAND2_X1 U7630 ( .A1(n7018), .A2(n7019), .ZN(n9016) );
  AOI21_X1 U7631 ( .B1(n7021), .B2(n8653), .A(n7020), .ZN(n7019) );
  INV_X1 U7632 ( .A(n8657), .ZN(n7020) );
  INV_X1 U7633 ( .A(n8991), .ZN(n7025) );
  NAND2_X1 U7634 ( .A1(n8593), .A2(n8592), .ZN(n8599) );
  INV_X1 U7635 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8592) );
  INV_X1 U7636 ( .A(n8595), .ZN(n8593) );
  NAND2_X1 U7637 ( .A1(n7030), .A2(n7031), .ZN(n8954) );
  AOI21_X1 U7638 ( .B1(n7033), .B2(n8641), .A(n7032), .ZN(n7031) );
  INV_X1 U7639 ( .A(n8644), .ZN(n7032) );
  NAND2_X1 U7640 ( .A1(n8631), .A2(n8630), .ZN(n8846) );
  INV_X1 U7641 ( .A(n14500), .ZN(n7158) );
  NAND2_X1 U7642 ( .A1(n13031), .A2(n7815), .ZN(n14501) );
  NAND2_X1 U7643 ( .A1(n7771), .A2(n6436), .ZN(n7610) );
  NAND2_X2 U7644 ( .A1(n13548), .A2(n8192), .ZN(n7771) );
  NAND2_X1 U7645 ( .A1(n12115), .A2(n7944), .ZN(n6677) );
  NOR2_X1 U7646 ( .A1(n8464), .A2(n8463), .ZN(n7386) );
  NAND2_X1 U7647 ( .A1(n8538), .A2(n7389), .ZN(n7388) );
  NAND2_X1 U7648 ( .A1(n7391), .A2(n7390), .ZN(n7389) );
  NAND2_X1 U7649 ( .A1(n8464), .A2(n8463), .ZN(n7387) );
  NAND2_X1 U7650 ( .A1(n7591), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7531) );
  NAND2_X1 U7651 ( .A1(n7570), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7530) );
  AOI21_X1 U7652 ( .B1(n7203), .B2(n7208), .A(n6540), .ZN(n7200) );
  NAND2_X1 U7653 ( .A1(n11275), .A2(n11200), .ZN(n11387) );
  INV_X1 U7654 ( .A(n10483), .ZN(n7228) );
  NAND2_X1 U7655 ( .A1(n10283), .A2(n10282), .ZN(n10286) );
  BUF_X1 U7656 ( .A(n7582), .Z(n8510) );
  XNOR2_X1 U7657 ( .A(n7197), .B(n11564), .ZN(n13436) );
  INV_X1 U7658 ( .A(n11563), .ZN(n11564) );
  AND2_X1 U7659 ( .A1(n14906), .A2(n8162), .ZN(n9994) );
  INV_X1 U7660 ( .A(n7879), .ZN(n6841) );
  NOR2_X1 U7661 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(n7491), .ZN(n7163) );
  NOR2_X1 U7662 ( .A1(n7273), .A2(n6614), .ZN(n6613) );
  INV_X1 U7663 ( .A(n11582), .ZN(n6614) );
  INV_X1 U7664 ( .A(n7274), .ZN(n7273) );
  NAND2_X1 U7665 ( .A1(n10165), .A2(n10164), .ZN(n10166) );
  NAND2_X1 U7666 ( .A1(n9280), .A2(n9691), .ZN(n9693) );
  INV_X1 U7667 ( .A(n7265), .ZN(n7264) );
  OAI21_X1 U7668 ( .B1(n7267), .B2(n7266), .A(n13644), .ZN(n7265) );
  INV_X1 U7669 ( .A(n11677), .ZN(n7266) );
  NAND2_X2 U7670 ( .A1(n14367), .A2(n9519), .ZN(n11818) );
  NAND2_X1 U7671 ( .A1(n13903), .A2(n6965), .ZN(n13808) );
  NOR2_X1 U7672 ( .A1(n13812), .A2(n6966), .ZN(n6965) );
  NAND2_X1 U7673 ( .A1(n6967), .A2(n13886), .ZN(n6966) );
  INV_X1 U7674 ( .A(n14109), .ZN(n6967) );
  NAND2_X1 U7675 ( .A1(n13905), .A2(n13832), .ZN(n7180) );
  INV_X1 U7676 ( .A(n7187), .ZN(n7186) );
  OAI21_X1 U7677 ( .B1(n7188), .B2(n6458), .A(n13856), .ZN(n7187) );
  AOI21_X1 U7678 ( .B1(n7174), .B2(n7172), .A(n6534), .ZN(n7171) );
  INV_X1 U7679 ( .A(n13846), .ZN(n7172) );
  INV_X1 U7680 ( .A(n7174), .ZN(n7173) );
  NAND2_X1 U7681 ( .A1(n7184), .A2(n6508), .ZN(n11341) );
  INV_X2 U7682 ( .A(n11610), .ZN(n12022) );
  NAND2_X1 U7683 ( .A1(n11035), .A2(n11034), .ZN(n11301) );
  INV_X1 U7684 ( .A(n10890), .ZN(n7168) );
  INV_X1 U7685 ( .A(n14720), .ZN(n14702) );
  NAND2_X1 U7686 ( .A1(n11891), .A2(n14741), .ZN(n6637) );
  NAND2_X1 U7687 ( .A1(n14742), .A2(n11891), .ZN(n6636) );
  NAND2_X1 U7688 ( .A1(n10656), .A2(n10655), .ZN(n6781) );
  NAND2_X1 U7689 ( .A1(n11879), .A2(n6517), .ZN(n6643) );
  INV_X1 U7690 ( .A(n14685), .ZN(n14744) );
  INV_X1 U7691 ( .A(n14118), .ZN(n6696) );
  AOI21_X1 U7692 ( .B1(n13912), .B2(n13858), .A(n6582), .ZN(n13894) );
  NAND2_X1 U7693 ( .A1(n13894), .A2(n13896), .ZN(n13893) );
  NAND2_X1 U7694 ( .A1(n13660), .A2(n13661), .ZN(n6616) );
  NAND2_X1 U7695 ( .A1(n8334), .A2(n8333), .ZN(n7380) );
  INV_X1 U7696 ( .A(n11925), .ZN(n6934) );
  NAND2_X1 U7697 ( .A1(n11930), .A2(n11931), .ZN(n11929) );
  NAND2_X1 U7698 ( .A1(n7461), .A2(n8375), .ZN(n7393) );
  NOR2_X1 U7699 ( .A1(n14082), .A2(n6944), .ZN(n6943) );
  NOR2_X1 U7700 ( .A1(n11948), .A2(n11949), .ZN(n6944) );
  AND2_X1 U7701 ( .A1(n8423), .A2(n8424), .ZN(n6837) );
  INV_X1 U7702 ( .A(n8418), .ZN(n7382) );
  NAND2_X1 U7703 ( .A1(n6836), .A2(n6835), .ZN(n6834) );
  INV_X1 U7704 ( .A(n8424), .ZN(n6836) );
  INV_X1 U7705 ( .A(n8423), .ZN(n6835) );
  NAND2_X1 U7706 ( .A1(n6931), .A2(n11995), .ZN(n6929) );
  OAI21_X1 U7707 ( .B1(n8441), .B2(n8440), .A(n6524), .ZN(n6816) );
  NAND2_X1 U7708 ( .A1(n12007), .A2(n12009), .ZN(n7256) );
  INV_X1 U7709 ( .A(n11472), .ZN(n7072) );
  OR2_X1 U7710 ( .A1(n8873), .A2(n8872), .ZN(n8875) );
  INV_X1 U7711 ( .A(n6761), .ZN(n6760) );
  OAI21_X1 U7712 ( .B1(n7965), .B2(n6762), .A(n8024), .ZN(n6761) );
  INV_X1 U7713 ( .A(n7721), .ZN(n6917) );
  INV_X1 U7714 ( .A(n6861), .ZN(n6860) );
  INV_X1 U7715 ( .A(n12395), .ZN(n6865) );
  NAND2_X1 U7716 ( .A1(n14990), .A2(n10539), .ZN(n6884) );
  OAI21_X1 U7717 ( .B1(n12623), .B2(n14491), .A(n15063), .ZN(n12591) );
  NAND2_X1 U7718 ( .A1(n6712), .A2(n6600), .ZN(n12594) );
  NAND2_X1 U7719 ( .A1(n15098), .A2(n6713), .ZN(n6712) );
  NAND2_X1 U7720 ( .A1(n6746), .A2(n6745), .ZN(n6744) );
  NAND2_X1 U7721 ( .A1(n12644), .A2(n12643), .ZN(n6745) );
  INV_X1 U7722 ( .A(n14441), .ZN(n6746) );
  INV_X1 U7723 ( .A(n12324), .ZN(n6867) );
  NOR2_X1 U7724 ( .A1(n9119), .A2(n6864), .ZN(n6863) );
  INV_X1 U7725 ( .A(n12318), .ZN(n6864) );
  OR2_X1 U7726 ( .A1(n9086), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9088) );
  INV_X1 U7727 ( .A(n9111), .ZN(n7406) );
  NAND2_X1 U7728 ( .A1(n7412), .A2(n9111), .ZN(n7408) );
  INV_X1 U7729 ( .A(n12279), .ZN(n6872) );
  OR2_X1 U7730 ( .A1(n12918), .A2(n12544), .ZN(n12275) );
  NAND2_X1 U7731 ( .A1(n8936), .A2(n12262), .ZN(n7060) );
  INV_X1 U7732 ( .A(n9110), .ZN(n7421) );
  NAND2_X1 U7733 ( .A1(n7423), .A2(n7420), .ZN(n7418) );
  NAND2_X1 U7734 ( .A1(n7422), .A2(n7424), .ZN(n7416) );
  INV_X1 U7735 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n8635) );
  INV_X1 U7736 ( .A(n7011), .ZN(n7010) );
  OAI21_X1 U7737 ( .B1(n8630), .B2(n7012), .A(n8633), .ZN(n7011) );
  INV_X1 U7738 ( .A(n8632), .ZN(n7012) );
  INV_X1 U7739 ( .A(n8623), .ZN(n7027) );
  NAND2_X1 U7740 ( .A1(n8615), .A2(n8616), .ZN(n7017) );
  INV_X1 U7741 ( .A(n8616), .ZN(n7014) );
  NOR2_X1 U7742 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n8584) );
  INV_X1 U7743 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8158) );
  INV_X1 U7744 ( .A(n8132), .ZN(n6660) );
  XNOR2_X1 U7745 ( .A(n12975), .B(n8086), .ZN(n7696) );
  INV_X1 U7746 ( .A(n13065), .ZN(n7150) );
  NOR2_X1 U7747 ( .A1(n7802), .A2(n14854), .ZN(n7822) );
  INV_X1 U7748 ( .A(n7328), .ZN(n7326) );
  NAND2_X1 U7749 ( .A1(n13289), .A2(n6480), .ZN(n7327) );
  INV_X1 U7750 ( .A(n11554), .ZN(n7219) );
  OR2_X1 U7751 ( .A1(n11201), .A2(n7223), .ZN(n7222) );
  INV_X1 U7752 ( .A(n11382), .ZN(n7223) );
  INV_X1 U7753 ( .A(n11523), .ZN(n7346) );
  OR2_X1 U7754 ( .A1(n13498), .A2(n14517), .ZN(n11523) );
  OR2_X1 U7755 ( .A1(n7210), .A2(n11209), .ZN(n7209) );
  NAND2_X1 U7756 ( .A1(n7213), .A2(n11143), .ZN(n7210) );
  INV_X1 U7757 ( .A(n10427), .ZN(n7342) );
  INV_X1 U7758 ( .A(n10394), .ZN(n7344) );
  INV_X1 U7759 ( .A(n7590), .ZN(n8130) );
  NAND2_X1 U7760 ( .A1(n13579), .A2(n10160), .ZN(n10165) );
  NOR2_X1 U7761 ( .A1(n13596), .A2(n7268), .ZN(n7267) );
  INV_X1 U7762 ( .A(n11658), .ZN(n7268) );
  NAND2_X1 U7763 ( .A1(n6904), .A2(n6903), .ZN(n6902) );
  INV_X1 U7764 ( .A(n12059), .ZN(n6903) );
  XNOR2_X1 U7765 ( .A(n6905), .B(n12058), .ZN(n6904) );
  OR2_X1 U7766 ( .A1(n14154), .A2(n14017), .ZN(n13849) );
  AND2_X1 U7767 ( .A1(n6964), .A2(n14544), .ZN(n6963) );
  INV_X1 U7768 ( .A(n14194), .ZN(n6964) );
  INV_X1 U7769 ( .A(n10886), .ZN(n7307) );
  NOR2_X1 U7770 ( .A1(n10758), .A2(n11136), .ZN(n10852) );
  INV_X1 U7771 ( .A(n14743), .ZN(n6639) );
  NOR2_X1 U7772 ( .A1(n9514), .A2(n9515), .ZN(n10225) );
  INV_X1 U7773 ( .A(n11876), .ZN(n9600) );
  AND3_X1 U7774 ( .A1(n9245), .A2(n7453), .A3(n9269), .ZN(n9246) );
  XNOR2_X1 U7775 ( .A(n8170), .B(n11332), .ZN(n8169) );
  NAND2_X1 U7776 ( .A1(n6777), .A2(n8059), .ZN(n8082) );
  NAND2_X1 U7777 ( .A1(n8057), .A2(n8056), .ZN(n6777) );
  NOR2_X1 U7778 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n9224) );
  INV_X1 U7779 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9216) );
  INV_X1 U7780 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9215) );
  INV_X1 U7781 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9207) );
  INV_X1 U7782 ( .A(n7796), .ZN(n7794) );
  INV_X1 U7783 ( .A(n7797), .ZN(n7795) );
  INV_X1 U7784 ( .A(n7246), .ZN(n7245) );
  OAI21_X1 U7785 ( .B1(n7247), .B2(n7724), .A(n7761), .ZN(n7246) );
  INV_X1 U7786 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n8205) );
  OR2_X1 U7787 ( .A1(n8254), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n7116) );
  AOI22_X1 U7788 ( .A1(n8272), .A2(n8213), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n15007), .ZN(n8214) );
  OAI21_X1 U7789 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n8218), .A(n8217), .ZN(
        n8252) );
  AOI21_X1 U7790 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n14311), .A(n8227), .ZN(
        n8245) );
  INV_X1 U7791 ( .A(n10451), .ZN(n7086) );
  NAND2_X1 U7792 ( .A1(n12169), .A2(n12168), .ZN(n12179) );
  NAND2_X1 U7793 ( .A1(n8698), .A2(n8697), .ZN(n8972) );
  INV_X1 U7794 ( .A(n10450), .ZN(n7085) );
  NOR2_X1 U7795 ( .A1(n7083), .A2(n10453), .ZN(n7082) );
  INV_X1 U7796 ( .A(n7089), .ZN(n7083) );
  NAND2_X1 U7797 ( .A1(n11255), .A2(n7107), .ZN(n7104) );
  INV_X1 U7798 ( .A(n11253), .ZN(n7107) );
  NAND2_X1 U7799 ( .A1(n11418), .A2(n11412), .ZN(n7102) );
  INV_X1 U7800 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11430) );
  AND2_X1 U7801 ( .A1(n11413), .A2(n11412), .ZN(n11481) );
  NAND2_X1 U7802 ( .A1(n9097), .A2(n7095), .ZN(n10098) );
  NAND2_X1 U7803 ( .A1(n7092), .A2(n7091), .ZN(n7095) );
  INV_X1 U7804 ( .A(n7065), .ZN(n7064) );
  NAND2_X1 U7805 ( .A1(n11473), .A2(n7068), .ZN(n7067) );
  OAI22_X1 U7806 ( .A1(n12458), .A2(n7066), .B1(n12545), .B2(n12138), .ZN(
        n7065) );
  AND2_X1 U7807 ( .A1(n12450), .A2(n7078), .ZN(n7077) );
  OR2_X1 U7808 ( .A1(n12476), .A2(n7079), .ZN(n7078) );
  INV_X1 U7809 ( .A(n12164), .ZN(n7079) );
  OR2_X1 U7810 ( .A1(n9201), .A2(n12185), .ZN(n12397) );
  NOR2_X1 U7811 ( .A1(n9915), .A2(n6875), .ZN(n9916) );
  AND2_X1 U7812 ( .A1(n8737), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n6875) );
  XNOR2_X1 U7813 ( .A(n10521), .B(n6874), .ZN(n9917) );
  OR2_X1 U7814 ( .A1(n9916), .A2(n9917), .ZN(n6989) );
  OR2_X1 U7815 ( .A1(n14971), .A2(n10537), .ZN(n6993) );
  NAND2_X1 U7816 ( .A1(n6993), .A2(n6992), .ZN(n14990) );
  INV_X1 U7817 ( .A(n14992), .ZN(n6992) );
  OR2_X1 U7818 ( .A1(n10957), .A2(n10956), .ZN(n12561) );
  INV_X1 U7819 ( .A(n6601), .ZN(n6752) );
  NAND2_X1 U7820 ( .A1(n6749), .A2(n6752), .ZN(n6748) );
  INV_X1 U7821 ( .A(n15035), .ZN(n6749) );
  NAND2_X1 U7822 ( .A1(n15013), .A2(n6750), .ZN(n6747) );
  NOR2_X1 U7823 ( .A1(n15035), .A2(n6751), .ZN(n6750) );
  INV_X1 U7824 ( .A(n15011), .ZN(n6751) );
  NAND2_X1 U7825 ( .A1(n7000), .A2(n15049), .ZN(n6999) );
  INV_X1 U7826 ( .A(n12567), .ZN(n7000) );
  NAND2_X1 U7827 ( .A1(n6877), .A2(n6583), .ZN(n6997) );
  XNOR2_X1 U7828 ( .A(n12591), .B(n12629), .ZN(n15080) );
  NAND2_X1 U7829 ( .A1(n15080), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n15079) );
  AND2_X1 U7830 ( .A1(n15071), .A2(n12625), .ZN(n15088) );
  NAND2_X1 U7831 ( .A1(n15059), .A2(n12570), .ZN(n6985) );
  NAND2_X1 U7832 ( .A1(n15088), .A2(n15089), .ZN(n15087) );
  NAND2_X1 U7833 ( .A1(n6984), .A2(n12635), .ZN(n12574) );
  NOR2_X1 U7834 ( .A1(n8941), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n8955) );
  XNOR2_X1 U7835 ( .A(n6744), .B(n6743), .ZN(n14458) );
  NAND2_X1 U7836 ( .A1(n6879), .A2(n6519), .ZN(n6991) );
  INV_X1 U7837 ( .A(n14449), .ZN(n6879) );
  NAND2_X1 U7838 ( .A1(n6991), .A2(n6990), .ZN(n14464) );
  INV_X1 U7839 ( .A(n14465), .ZN(n6990) );
  NOR2_X1 U7840 ( .A1(n6744), .A2(n6743), .ZN(n6742) );
  NAND2_X1 U7841 ( .A1(n6867), .A2(n6862), .ZN(n6861) );
  INV_X1 U7842 ( .A(n12325), .ZN(n6862) );
  INV_X1 U7843 ( .A(n9196), .ZN(n12384) );
  AOI21_X1 U7844 ( .B1(n9122), .B2(n12320), .A(n6546), .ZN(n7430) );
  AND2_X1 U7845 ( .A1(n12397), .A2(n12393), .ZN(n9196) );
  OR2_X1 U7846 ( .A1(n12516), .A2(n12453), .ZN(n12318) );
  NAND2_X1 U7847 ( .A1(n6851), .A2(n12310), .ZN(n6850) );
  NAND2_X1 U7848 ( .A1(n9045), .A2(n6853), .ZN(n12710) );
  NAND2_X1 U7849 ( .A1(n7038), .A2(n12302), .ZN(n12723) );
  AOI21_X1 U7850 ( .B1(n7412), .B2(n7410), .A(n6545), .ZN(n7409) );
  INV_X1 U7851 ( .A(n12760), .ZN(n7410) );
  AND4_X1 U7852 ( .A1(n9013), .A2(n9012), .A3(n9011), .A4(n9010), .ZN(n12746)
         );
  NAND2_X1 U7853 ( .A1(n12756), .A2(n12760), .ZN(n7413) );
  AND2_X1 U7854 ( .A1(n7413), .A2(n6505), .ZN(n12743) );
  NAND2_X1 U7855 ( .A1(n9014), .A2(n12292), .ZN(n12749) );
  OR2_X1 U7856 ( .A1(n12759), .A2(n12760), .ZN(n9014) );
  AND3_X1 U7857 ( .A1(n9025), .A2(n9024), .A3(n9023), .ZN(n12758) );
  OAI21_X1 U7858 ( .B1(n7435), .B2(n7434), .A(n6544), .ZN(n7433) );
  NOR2_X1 U7859 ( .A1(n12373), .A2(n12258), .ZN(n7437) );
  INV_X1 U7860 ( .A(n7436), .ZN(n7435) );
  OAI21_X1 U7861 ( .B1(n12373), .B2(n7441), .A(n7439), .ZN(n7436) );
  NAND2_X1 U7862 ( .A1(n7440), .A2(n12546), .ZN(n7439) );
  INV_X1 U7863 ( .A(n12925), .ZN(n7440) );
  INV_X1 U7864 ( .A(n12545), .ZN(n12798) );
  INV_X1 U7865 ( .A(n8917), .ZN(n8694) );
  AOI21_X1 U7866 ( .B1(n11222), .B2(n7053), .A(n7052), .ZN(n7051) );
  INV_X1 U7867 ( .A(n12250), .ZN(n7052) );
  INV_X1 U7868 ( .A(n12247), .ZN(n7053) );
  NOR2_X1 U7869 ( .A1(n12370), .A2(n6856), .ZN(n6855) );
  INV_X1 U7870 ( .A(n12374), .ZN(n6856) );
  AND4_X1 U7871 ( .A1(n8901), .A2(n8900), .A3(n8899), .A4(n8898), .ZN(n11423)
         );
  AND4_X1 U7872 ( .A1(n8843), .A2(n8842), .A3(n8841), .A4(n8840), .ZN(n11245)
         );
  NAND2_X1 U7873 ( .A1(n11246), .A2(n12374), .ZN(n11247) );
  NAND2_X1 U7874 ( .A1(n11065), .A2(n12243), .ZN(n11064) );
  NAND2_X1 U7875 ( .A1(n8691), .A2(n11183), .ZN(n8855) );
  INV_X1 U7876 ( .A(n8853), .ZN(n8691) );
  NAND2_X1 U7877 ( .A1(n10830), .A2(n12362), .ZN(n10829) );
  INV_X1 U7878 ( .A(n12766), .ZN(n15128) );
  NOR2_X2 U7879 ( .A1(n12559), .A2(n11836), .ZN(n12193) );
  NAND2_X1 U7880 ( .A1(n9006), .A2(n9005), .ZN(n12482) );
  INV_X1 U7881 ( .A(n12333), .ZN(n8993) );
  INV_X1 U7882 ( .A(n12769), .ZN(n15122) );
  NAND2_X1 U7883 ( .A1(n9143), .A2(n9159), .ZN(n9395) );
  NAND2_X1 U7884 ( .A1(n9183), .A2(n9182), .ZN(n11494) );
  NAND2_X1 U7885 ( .A1(n7001), .A2(n8670), .ZN(n9083) );
  NAND2_X1 U7886 ( .A1(n9058), .A2(n8667), .ZN(n9069) );
  INV_X1 U7887 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7061) );
  NAND2_X1 U7888 ( .A1(n7003), .A2(n7002), .ZN(n9037) );
  AOI21_X1 U7889 ( .B1(n7005), .B2(n7007), .A(n6597), .ZN(n7002) );
  NAND2_X1 U7890 ( .A1(n8659), .A2(n7005), .ZN(n7003) );
  XNOR2_X1 U7891 ( .A(n9162), .B(n9161), .ZN(n9885) );
  INV_X1 U7892 ( .A(n9016), .ZN(n8659) );
  OR2_X1 U7893 ( .A1(n7444), .A2(n8676), .ZN(n8595) );
  NAND2_X1 U7894 ( .A1(n8979), .A2(n8650), .ZN(n8652) );
  AND2_X1 U7895 ( .A1(n8646), .A2(n8645), .ZN(n8953) );
  NAND2_X1 U7896 ( .A1(n8954), .A2(n8953), .ZN(n8952) );
  NAND2_X1 U7897 ( .A1(n7037), .A2(n7036), .ZN(n7035) );
  INV_X1 U7898 ( .A(n8926), .ZN(n7037) );
  INV_X1 U7899 ( .A(n8642), .ZN(n7034) );
  NAND2_X1 U7900 ( .A1(n8902), .A2(n6491), .ZN(n7444) );
  NAND2_X1 U7901 ( .A1(n8626), .A2(n8625), .ZN(n8865) );
  NAND2_X1 U7902 ( .A1(n8835), .A2(n8624), .ZN(n8626) );
  NAND2_X1 U7903 ( .A1(n9373), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8623) );
  INV_X1 U7904 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8816) );
  INV_X1 U7905 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7428) );
  INV_X1 U7906 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7039) );
  AND2_X1 U7907 ( .A1(n6481), .A2(n6660), .ZN(n6659) );
  OAI21_X1 U7908 ( .B1(n6481), .B2(n8132), .A(n6657), .ZN(n6656) );
  NAND2_X1 U7909 ( .A1(n6481), .A2(n6658), .ZN(n6657) );
  NAND2_X1 U7910 ( .A1(n7146), .A2(n6660), .ZN(n6658) );
  NAND2_X1 U7911 ( .A1(n6662), .A2(n8132), .ZN(n6661) );
  INV_X1 U7912 ( .A(n7146), .ZN(n6662) );
  NOR2_X1 U7913 ( .A1(n12962), .A2(n7161), .ZN(n7160) );
  INV_X1 U7914 ( .A(n7720), .ZN(n7161) );
  OAI21_X1 U7915 ( .B1(n6668), .B2(n6665), .A(n6549), .ZN(n14514) );
  INV_X1 U7916 ( .A(n6666), .ZN(n6665) );
  NAND2_X1 U7917 ( .A1(n7154), .A2(n7851), .ZN(n7153) );
  XNOR2_X1 U7918 ( .A(n10073), .B(n7590), .ZN(n9969) );
  NOR2_X1 U7919 ( .A1(n11264), .A2(n11099), .ZN(n9431) );
  XNOR2_X1 U7920 ( .A(n7696), .B(n7697), .ZN(n12978) );
  NAND2_X1 U7921 ( .A1(n12985), .A2(n12984), .ZN(n7982) );
  XNOR2_X1 U7922 ( .A(n12966), .B(n8086), .ZN(n12120) );
  NAND2_X1 U7923 ( .A1(n13012), .A2(n7151), .ZN(n12107) );
  NOR2_X1 U7924 ( .A1(n13058), .A2(n7152), .ZN(n7151) );
  INV_X1 U7925 ( .A(n7897), .ZN(n7152) );
  OR2_X1 U7926 ( .A1(n7886), .A2(n7885), .ZN(n7913) );
  NAND2_X1 U7927 ( .A1(n9979), .A2(n7162), .ZN(n10089) );
  AND2_X1 U7928 ( .A1(n7648), .A2(n7628), .ZN(n7162) );
  NAND2_X1 U7929 ( .A1(n7822), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7842) );
  NOR2_X1 U7930 ( .A1(n9234), .A2(n7157), .ZN(n7156) );
  INV_X1 U7931 ( .A(n7831), .ZN(n7157) );
  NAND2_X1 U7932 ( .A1(n6772), .A2(n6771), .ZN(n8533) );
  AND2_X1 U7933 ( .A1(n8093), .A2(n8092), .ZN(n11558) );
  NAND2_X1 U7934 ( .A1(n7570), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7525) );
  XNOR2_X1 U7935 ( .A(n9526), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n9427) );
  OR2_X1 U7936 ( .A1(n13117), .A2(n13116), .ZN(n6972) );
  AND2_X1 U7937 ( .A1(n6972), .A2(n6971), .ZN(n13132) );
  NAND2_X1 U7938 ( .A1(n13125), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6971) );
  OR2_X1 U7939 ( .A1(n13132), .A2(n13131), .ZN(n6970) );
  NOR2_X1 U7940 ( .A1(n13241), .A2(n13434), .ZN(n7127) );
  AND2_X1 U7941 ( .A1(n13235), .A2(n11571), .ZN(n13433) );
  NAND2_X1 U7942 ( .A1(n13292), .A2(n7322), .ZN(n7321) );
  NAND2_X1 U7943 ( .A1(n11552), .A2(n6484), .ZN(n13309) );
  OAI21_X1 U7944 ( .B1(n7230), .B2(n11548), .A(n6632), .ZN(n13320) );
  AOI21_X1 U7945 ( .B1(n7234), .B2(n7231), .A(n6468), .ZN(n6632) );
  NAND2_X1 U7946 ( .A1(n7356), .A2(n7354), .ZN(n13329) );
  NAND2_X1 U7947 ( .A1(n13354), .A2(n6518), .ZN(n7356) );
  INV_X1 U7948 ( .A(n7460), .ZN(n7355) );
  NAND2_X1 U7949 ( .A1(n11548), .A2(n7233), .ZN(n7232) );
  NOR2_X1 U7950 ( .A1(n11389), .A2(n7350), .ZN(n7349) );
  INV_X1 U7951 ( .A(n11388), .ZN(n7350) );
  NAND2_X1 U7952 ( .A1(n11387), .A2(n11386), .ZN(n7351) );
  NAND2_X1 U7953 ( .A1(n7840), .A2(n7839), .ZN(n11273) );
  NOR2_X1 U7954 ( .A1(n11209), .A2(n7212), .ZN(n7211) );
  INV_X1 U7955 ( .A(n7213), .ZN(n7212) );
  INV_X1 U7956 ( .A(n7361), .ZN(n7360) );
  AOI21_X1 U7957 ( .B1(n10673), .B2(n10902), .A(n6527), .ZN(n7361) );
  NAND2_X1 U7958 ( .A1(n11146), .A2(n13084), .ZN(n7213) );
  OR2_X1 U7959 ( .A1(n10674), .A2(n10673), .ZN(n10903) );
  AOI21_X1 U7960 ( .B1(n6456), .B2(n10482), .A(n6462), .ZN(n7225) );
  NAND2_X1 U7961 ( .A1(n14923), .A2(n10476), .ZN(n7229) );
  INV_X1 U7962 ( .A(n10475), .ZN(n10669) );
  NAND2_X1 U7963 ( .A1(n10426), .A2(n10425), .ZN(n10483) );
  OAI21_X1 U7964 ( .B1(n9926), .B2(n7216), .A(n7214), .ZN(n10283) );
  INV_X1 U7965 ( .A(n7215), .ZN(n7214) );
  INV_X1 U7966 ( .A(n10014), .ZN(n7216) );
  NAND2_X1 U7967 ( .A1(n9926), .A2(n9930), .ZN(n10015) );
  INV_X1 U7968 ( .A(n13406), .ZN(n13294) );
  NAND2_X1 U7969 ( .A1(n9575), .A2(n9574), .ZN(n9577) );
  NOR2_X1 U7970 ( .A1(n9999), .A2(n11264), .ZN(n7489) );
  XNOR2_X1 U7971 ( .A(n13434), .B(n13073), .ZN(n11563) );
  AND2_X1 U7972 ( .A1(n7196), .A2(n7195), .ZN(n7334) );
  AOI21_X1 U7973 ( .B1(n13434), .B2(n13513), .A(n11541), .ZN(n7195) );
  INV_X1 U7974 ( .A(n13433), .ZN(n7196) );
  NAND2_X1 U7975 ( .A1(n7864), .A2(n7863), .ZN(n13504) );
  OR2_X1 U7976 ( .A1(n10320), .A2(n7908), .ZN(n7636) );
  INV_X1 U7977 ( .A(n14922), .ZN(n13513) );
  AND2_X1 U7978 ( .A1(n9456), .A2(n9455), .ZN(n9996) );
  NAND2_X1 U7979 ( .A1(n11264), .A2(n8182), .ZN(n10420) );
  NOR2_X1 U7980 ( .A1(n11338), .A2(n8154), .ZN(n14873) );
  AND2_X1 U7981 ( .A1(n11170), .A2(n8153), .ZN(n8154) );
  NOR2_X1 U7982 ( .A1(n7497), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n6839) );
  NAND2_X1 U7983 ( .A1(n8146), .A2(n7455), .ZN(n7504) );
  NAND2_X1 U7984 ( .A1(n8142), .A2(n8141), .ZN(n8148) );
  INV_X1 U7985 ( .A(n8146), .ZN(n8142) );
  NOR2_X1 U7986 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7363) );
  NOR2_X1 U7987 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n7362) );
  INV_X1 U7988 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8608) );
  NAND2_X1 U7989 ( .A1(n11614), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n11631) );
  NAND2_X1 U7990 ( .A1(n13570), .A2(n6611), .ZN(n6610) );
  INV_X1 U7991 ( .A(n11696), .ZN(n6611) );
  NAND2_X1 U7992 ( .A1(n10166), .A2(n7271), .ZN(n7270) );
  INV_X1 U7993 ( .A(n10168), .ZN(n7271) );
  AND2_X1 U7994 ( .A1(n7263), .A2(n9276), .ZN(n9280) );
  OAI211_X1 U7995 ( .C1(n9766), .C2(n6617), .A(n9279), .B(n6543), .ZN(n9691)
         );
  NAND2_X1 U7996 ( .A1(n13634), .A2(n7267), .ZN(n13593) );
  OAI21_X1 U7997 ( .B1(n11131), .B2(n6608), .A(n6605), .ZN(n7279) );
  INV_X1 U7998 ( .A(n11134), .ZN(n6608) );
  AND2_X1 U7999 ( .A1(n7280), .A2(n6606), .ZN(n6605) );
  NOR2_X1 U8000 ( .A1(n11234), .A2(n7281), .ZN(n7280) );
  AND4_X1 U8001 ( .A1(n11043), .A2(n11042), .A3(n11041), .A4(n11040), .ZN(
        n11585) );
  NAND2_X1 U8002 ( .A1(n6471), .A2(n14367), .ZN(n6924) );
  NAND2_X1 U8003 ( .A1(n6927), .A2(n14370), .ZN(n6925) );
  AND2_X1 U8004 ( .A1(n9521), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6927) );
  NAND2_X1 U8005 ( .A1(n13708), .A2(n6686), .ZN(n9322) );
  NOR2_X1 U8006 ( .A1(n9318), .A2(n6893), .ZN(n13720) );
  AND2_X1 U8007 ( .A1(n9307), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6893) );
  OR2_X1 U8008 ( .A1(n13720), .A2(n13719), .ZN(n6892) );
  NOR2_X1 U8009 ( .A1(n14592), .A2(n6895), .ZN(n10351) );
  AND2_X1 U8010 ( .A1(n14597), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6895) );
  NAND2_X1 U8011 ( .A1(n14614), .A2(n6887), .ZN(n13784) );
  OR2_X1 U8012 ( .A1(n13783), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6887) );
  NAND2_X1 U8013 ( .A1(n12025), .A2(n12024), .ZN(n14109) );
  INV_X1 U8014 ( .A(n13837), .ZN(n13861) );
  NAND2_X1 U8015 ( .A1(n13935), .A2(n7449), .ZN(n13912) );
  OR2_X1 U8016 ( .A1(n13857), .A2(n13960), .ZN(n7449) );
  NAND2_X1 U8017 ( .A1(n6808), .A2(n6812), .ZN(n6807) );
  AND2_X1 U8018 ( .A1(n13938), .A2(n13830), .ZN(n7317) );
  NAND2_X1 U8019 ( .A1(n13972), .A2(n13828), .ZN(n13959) );
  OR2_X1 U8020 ( .A1(n13959), .A2(n13958), .ZN(n13963) );
  NOR2_X1 U8021 ( .A1(n13855), .A2(n7189), .ZN(n7188) );
  INV_X1 U8022 ( .A(n13853), .ZN(n7189) );
  INV_X1 U8023 ( .A(n13827), .ZN(n13973) );
  NAND2_X1 U8024 ( .A1(n13982), .A2(n13850), .ZN(n13854) );
  NAND2_X1 U8025 ( .A1(n13997), .A2(n13849), .ZN(n13982) );
  AOI21_X1 U8026 ( .B1(n13993), .B2(n13999), .A(n13824), .ZN(n13979) );
  AND2_X1 U8027 ( .A1(n14050), .A2(n7294), .ZN(n7293) );
  OR2_X1 U8028 ( .A1(n14174), .A2(n14065), .ZN(n13846) );
  NOR2_X1 U8029 ( .A1(n13818), .A2(n7300), .ZN(n7299) );
  INV_X1 U8030 ( .A(n13814), .ZN(n7300) );
  NAND2_X1 U8031 ( .A1(n11603), .A2(n11602), .ZN(n14070) );
  AOI21_X1 U8032 ( .B1(n7450), .B2(n6796), .A(n6539), .ZN(n6795) );
  INV_X1 U8033 ( .A(n11340), .ZN(n6796) );
  INV_X1 U8034 ( .A(n7450), .ZN(n6797) );
  OR2_X1 U8035 ( .A1(n11353), .A2(n11352), .ZN(n13815) );
  INV_X1 U8036 ( .A(n12051), .ZN(n11352) );
  OR2_X1 U8037 ( .A1(n13686), .A2(n13690), .ZN(n11340) );
  NAND2_X1 U8038 ( .A1(n14194), .A2(n13691), .ZN(n7183) );
  NOR2_X1 U8039 ( .A1(n14078), .A2(n7182), .ZN(n7181) );
  INV_X1 U8040 ( .A(n7185), .ZN(n7182) );
  NAND2_X1 U8041 ( .A1(n11936), .A2(n13693), .ZN(n6790) );
  NAND2_X1 U8042 ( .A1(n7311), .A2(n7310), .ZN(n10887) );
  INV_X1 U8043 ( .A(n12043), .ZN(n7310) );
  INV_X1 U8044 ( .A(n10849), .ZN(n7311) );
  INV_X1 U8045 ( .A(n6787), .ZN(n6783) );
  NAND2_X1 U8046 ( .A1(n14687), .A2(n6529), .ZN(n6782) );
  NOR2_X1 U8047 ( .A1(n10757), .A2(n6785), .ZN(n6784) );
  INV_X1 U8048 ( .A(n10755), .ZN(n6785) );
  INV_X1 U8049 ( .A(n13694), .ZN(n10888) );
  NAND2_X1 U8050 ( .A1(n10770), .A2(n10769), .ZN(n14681) );
  INV_X1 U8051 ( .A(n14090), .ZN(n14756) );
  NAND2_X1 U8052 ( .A1(n6640), .A2(n13821), .ZN(n14015) );
  NAND2_X1 U8053 ( .A1(n11001), .A2(n11000), .ZN(n11939) );
  INV_X1 U8054 ( .A(n14792), .ZN(n14821) );
  AND3_X1 U8055 ( .A1(n9243), .A2(n9242), .A3(n9241), .ZN(n9271) );
  INV_X1 U8056 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9242) );
  INV_X1 U8057 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9241) );
  NAND2_X1 U8058 ( .A1(n9261), .A2(n7284), .ZN(n9265) );
  NOR2_X1 U8059 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n7284) );
  INV_X1 U8060 ( .A(n9265), .ZN(n9257) );
  NOR2_X1 U8061 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n9256) );
  INV_X1 U8062 ( .A(n7905), .ZN(n7261) );
  NAND2_X1 U8063 ( .A1(n7742), .A2(n7741), .ZN(n7763) );
  AND2_X1 U8064 ( .A1(n10211), .A2(n9401), .ZN(n9416) );
  INV_X1 U8065 ( .A(n7632), .ZN(n7633) );
  INV_X1 U8066 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n8204) );
  XNOR2_X1 U8067 ( .A(n8206), .B(n7123), .ZN(n8256) );
  NAND2_X1 U8068 ( .A1(n14389), .A2(n8282), .ZN(n8285) );
  NAND2_X1 U8069 ( .A1(n8223), .A2(n8222), .ZN(n8249) );
  INV_X1 U8070 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7112) );
  AND3_X1 U8071 ( .A1(n8851), .A2(n8850), .A3(n8849), .ZN(n15153) );
  INV_X1 U8072 ( .A(n12540), .ZN(n12747) );
  NAND2_X1 U8073 ( .A1(n12485), .A2(n12151), .ZN(n12442) );
  NAND2_X1 U8074 ( .A1(n9060), .A2(n9059), .ZN(n12698) );
  OR2_X1 U8075 ( .A1(n12333), .A2(n11830), .ZN(n9059) );
  OR2_X1 U8076 ( .A1(n11831), .A2(n8888), .ZN(n9060) );
  INV_X1 U8077 ( .A(n12922), .ZN(n12463) );
  AND4_X1 U8078 ( .A1(n8800), .A2(n8799), .A3(n8798), .A4(n8797), .ZN(n10921)
         );
  AND2_X1 U8079 ( .A1(n9067), .A2(n9066), .ZN(n12677) );
  NAND2_X1 U8080 ( .A1(n9048), .A2(n9047), .ZN(n12712) );
  OR2_X1 U8081 ( .A1(n12333), .A2(n10928), .ZN(n9047) );
  AND4_X1 U8082 ( .A1(n9001), .A2(n9000), .A3(n8999), .A4(n8998), .ZN(n12785)
         );
  AND3_X1 U8083 ( .A1(n9044), .A2(n9043), .A3(n9042), .ZN(n12733) );
  NAND2_X1 U8084 ( .A1(n9031), .A2(n9030), .ZN(n12736) );
  INV_X1 U8085 ( .A(n12884), .ZN(n12516) );
  NOR2_X1 U8086 ( .A1(n12403), .A2(n12402), .ZN(n12405) );
  AND2_X1 U8087 ( .A1(n12353), .A2(n9192), .ZN(n12354) );
  NAND2_X1 U8088 ( .A1(n8720), .A2(n8719), .ZN(n12537) );
  INV_X1 U8089 ( .A(n11245), .ZN(n12550) );
  NOR2_X1 U8090 ( .A1(n9832), .A2(n9872), .ZN(n9903) );
  NAND2_X1 U8091 ( .A1(n9864), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9872) );
  NOR2_X1 U8092 ( .A1(n14972), .A2(n10633), .ZN(n14971) );
  OAI21_X1 U8093 ( .B1(n14976), .B2(n14973), .A(n10529), .ZN(n14989) );
  NAND2_X1 U8094 ( .A1(n14989), .A2(n14988), .ZN(n14987) );
  XNOR2_X1 U8095 ( .A(n6985), .B(n15084), .ZN(n15078) );
  INV_X1 U8096 ( .A(n11514), .ZN(n11515) );
  OAI21_X1 U8097 ( .B1(n12086), .B2(n11513), .A(n11512), .ZN(n11514) );
  INV_X1 U8098 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8682) );
  NAND2_X1 U8099 ( .A1(n8712), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8683) );
  XNOR2_X1 U8100 ( .A(n8594), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12415) );
  OR3_X1 U8101 ( .A1(n11087), .A2(n11170), .A3(n11338), .ZN(n9432) );
  NAND2_X1 U8102 ( .A1(n7159), .A2(n7158), .ZN(n14504) );
  NAND2_X1 U8103 ( .A1(n12107), .A2(n7940), .ZN(n12115) );
  AND2_X1 U8104 ( .A1(n12109), .A2(n7939), .ZN(n7940) );
  NAND2_X1 U8105 ( .A1(n6663), .A2(n14515), .ZN(n8185) );
  OAI211_X1 U8106 ( .C1(n8080), .C2(n6655), .A(n6652), .B(n14523), .ZN(n6663)
         );
  NAND2_X1 U8107 ( .A1(n6656), .A2(n6661), .ZN(n6655) );
  NAND2_X1 U8108 ( .A1(n8080), .A2(n6653), .ZN(n6652) );
  NAND2_X1 U8109 ( .A1(n6709), .A2(n6722), .ZN(n9990) );
  NAND2_X1 U8110 ( .A1(n9733), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14528) );
  NAND2_X1 U8111 ( .A1(n8129), .A2(n8128), .ZN(n13074) );
  INV_X1 U8112 ( .A(n11558), .ZN(n13076) );
  NAND2_X1 U8113 ( .A1(n8075), .A2(n8074), .ZN(n13077) );
  NOR2_X1 U8114 ( .A1(n9659), .A2(n9658), .ZN(n9802) );
  NOR2_X1 U8115 ( .A1(n9656), .A2(n6977), .ZN(n9659) );
  AND2_X1 U8116 ( .A1(n9660), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6977) );
  INV_X1 U8117 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n6622) );
  OAI21_X1 U8118 ( .B1(n13222), .B2(n14856), .A(n6983), .ZN(n6982) );
  AOI21_X1 U8119 ( .B1(n13221), .B2(n13224), .A(n14862), .ZN(n6983) );
  NAND2_X1 U8120 ( .A1(n7339), .A2(n13406), .ZN(n7335) );
  NAND2_X1 U8121 ( .A1(n7970), .A2(n7969), .ZN(n13477) );
  INV_X1 U8122 ( .A(n9758), .ZN(n7544) );
  AND2_X1 U8123 ( .A1(n14933), .A2(n13406), .ZN(n7333) );
  OR2_X1 U8124 ( .A1(n7334), .A2(n14931), .ZN(n7332) );
  OAI211_X1 U8125 ( .C1(n13516), .C2(n13436), .A(n7335), .B(n7334), .ZN(n6635)
         );
  NAND2_X1 U8126 ( .A1(n11131), .A2(n11130), .ZN(n11135) );
  NAND2_X1 U8127 ( .A1(n9700), .A2(n9768), .ZN(n9701) );
  OR2_X1 U8128 ( .A1(n9699), .A2(n9698), .ZN(n9700) );
  NAND2_X1 U8129 ( .A1(n13626), .A2(n13627), .ZN(n11736) );
  AOI21_X1 U8130 ( .B1(n7274), .B2(n11597), .A(n6587), .ZN(n7272) );
  NAND2_X1 U8131 ( .A1(n11583), .A2(n6613), .ZN(n6615) );
  AND2_X1 U8132 ( .A1(n10138), .A2(n6558), .ZN(n7190) );
  NAND2_X1 U8133 ( .A1(n6453), .A2(n6460), .ZN(n6921) );
  NAND2_X1 U8134 ( .A1(n6602), .A2(n11680), .ZN(n6922) );
  INV_X1 U8135 ( .A(n14149), .ZN(n13852) );
  AND4_X1 U8136 ( .A1(n11362), .A2(n11361), .A3(n11360), .A4(n11359), .ZN(
        n14052) );
  NAND4_X1 U8137 ( .A1(n11771), .A2(n11770), .A3(n11769), .A4(n11768), .ZN(
        n13933) );
  NAND2_X1 U8138 ( .A1(n14615), .A2(n14616), .ZN(n14614) );
  INV_X1 U8139 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n13799) );
  NAND2_X1 U8140 ( .A1(n6718), .A2(n6717), .ZN(n6716) );
  AOI21_X1 U8141 ( .B1(n6886), .B2(n14636), .A(n13796), .ZN(n6717) );
  INV_X1 U8142 ( .A(n13794), .ZN(n6886) );
  NAND2_X1 U8143 ( .A1(n13797), .A2(n13796), .ZN(n6719) );
  NAND2_X1 U8144 ( .A1(n11866), .A2(n11865), .ZN(n14098) );
  NAND2_X1 U8145 ( .A1(n13893), .A2(n7180), .ZN(n13880) );
  NAND2_X1 U8146 ( .A1(n7314), .A2(n7313), .ZN(n7312) );
  NAND2_X1 U8147 ( .A1(n13879), .A2(n14702), .ZN(n7313) );
  NAND2_X1 U8148 ( .A1(n7170), .A2(n7171), .ZN(n14011) );
  NAND2_X1 U8149 ( .A1(n14119), .A2(n14749), .ZN(n6805) );
  INV_X1 U8150 ( .A(n12058), .ZN(n13796) );
  NAND2_X1 U8151 ( .A1(n14579), .A2(n14578), .ZN(n14577) );
  NAND2_X1 U8152 ( .A1(n7122), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n7121) );
  XNOR2_X1 U8153 ( .A(n8301), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n8302) );
  OAI22_X1 U8154 ( .A1(n11898), .A2(n6946), .B1(n11897), .B2(n6945), .ZN(
        n11902) );
  INV_X1 U8155 ( .A(n11896), .ZN(n6945) );
  INV_X1 U8156 ( .A(n8347), .ZN(n7366) );
  INV_X1 U8157 ( .A(n8337), .ZN(n6688) );
  NAND2_X1 U8158 ( .A1(n6950), .A2(n11913), .ZN(n6949) );
  INV_X1 U8159 ( .A(n11924), .ZN(n6932) );
  NOR2_X1 U8160 ( .A1(n6934), .A2(n11924), .ZN(n6933) );
  NAND2_X1 U8161 ( .A1(n7398), .A2(n7397), .ZN(n7396) );
  INV_X1 U8162 ( .A(n8375), .ZN(n7397) );
  OR2_X1 U8163 ( .A1(n8362), .A2(n8361), .ZN(n8363) );
  AND2_X1 U8164 ( .A1(n8362), .A2(n8361), .ZN(n8364) );
  NAND2_X1 U8165 ( .A1(n7396), .A2(n7395), .ZN(n7394) );
  INV_X1 U8166 ( .A(n8369), .ZN(n7395) );
  NAND2_X1 U8167 ( .A1(n11937), .A2(n6937), .ZN(n6936) );
  NAND2_X1 U8168 ( .A1(n6943), .A2(n6523), .ZN(n6941) );
  NAND2_X1 U8169 ( .A1(n8385), .A2(n6515), .ZN(n6817) );
  NOR2_X1 U8170 ( .A1(n8385), .A2(n6515), .ZN(n6818) );
  NOR2_X1 U8171 ( .A1(n8418), .A2(n8420), .ZN(n7383) );
  AOI21_X1 U8172 ( .B1(n8425), .B2(n6834), .A(n6832), .ZN(n6831) );
  NAND2_X1 U8173 ( .A1(n8432), .A2(n6833), .ZN(n6832) );
  NAND2_X1 U8174 ( .A1(n6837), .A2(n6834), .ZN(n6833) );
  NAND2_X1 U8175 ( .A1(n11996), .A2(n11998), .ZN(n7258) );
  INV_X1 U8176 ( .A(n8445), .ZN(n7364) );
  NAND2_X1 U8177 ( .A1(n11858), .A2(n11844), .ZN(n11856) );
  INV_X1 U8178 ( .A(n15089), .ZN(n6756) );
  INV_X1 U8179 ( .A(n15099), .ZN(n6713) );
  AOI21_X1 U8180 ( .B1(n8451), .B2(n8450), .A(n8449), .ZN(n8452) );
  NAND2_X1 U8181 ( .A1(n13451), .A2(n11558), .ZN(n7328) );
  INV_X1 U8182 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n7463) );
  INV_X1 U8183 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7462) );
  INV_X1 U8184 ( .A(n12010), .ZN(n6919) );
  NOR2_X1 U8185 ( .A1(n12013), .A2(n12010), .ZN(n6920) );
  INV_X1 U8186 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9214) );
  AOI21_X1 U8187 ( .B1(n7239), .B2(n7241), .A(n7238), .ZN(n7237) );
  INV_X1 U8188 ( .A(n7852), .ZN(n7238) );
  OAI21_X1 U8189 ( .B1(n6450), .B2(n6703), .A(n6702), .ZN(n7759) );
  NAND2_X1 U8190 ( .A1(n6436), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n6702) );
  OAI21_X1 U8191 ( .B1(n6450), .B2(n10137), .A(n6708), .ZN(n7581) );
  NAND2_X1 U8192 ( .A1(n6436), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6708) );
  NAND2_X1 U8193 ( .A1(n12130), .A2(n7072), .ZN(n7071) );
  NAND2_X1 U8194 ( .A1(n10042), .A2(n10041), .ZN(n7090) );
  NAND2_X1 U8195 ( .A1(n7069), .A2(n7073), .ZN(n7066) );
  NOR2_X1 U8196 ( .A1(n12458), .A2(n7070), .ZN(n7068) );
  OR2_X1 U8197 ( .A1(n10544), .A2(n6735), .ZN(n10547) );
  NOR2_X1 U8198 ( .A1(n10521), .A2(n15161), .ZN(n6735) );
  NAND2_X1 U8199 ( .A1(n12584), .A2(n12585), .ZN(n12586) );
  NAND2_X1 U8200 ( .A1(n15028), .A2(n12588), .ZN(n12589) );
  AND2_X1 U8201 ( .A1(n12638), .A2(n12637), .ZN(n12640) );
  OAI21_X1 U8202 ( .B1(n14421), .B2(n12871), .A(n14427), .ZN(n12596) );
  NAND2_X1 U8203 ( .A1(n8707), .A2(n8706), .ZN(n9086) );
  NAND2_X1 U8204 ( .A1(n8705), .A2(n14320), .ZN(n9072) );
  INV_X1 U8205 ( .A(n9061), .ZN(n8705) );
  OR2_X1 U8206 ( .A1(n12698), .A2(n12677), .ZN(n12313) );
  INV_X1 U8207 ( .A(n6853), .ZN(n6851) );
  INV_X1 U8208 ( .A(n12310), .ZN(n6852) );
  OR2_X1 U8209 ( .A1(n9021), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n9032) );
  INV_X1 U8210 ( .A(n7051), .ZN(n7049) );
  AND2_X1 U8211 ( .A1(n8874), .A2(n6845), .ZN(n6844) );
  NAND2_X1 U8212 ( .A1(n6846), .A2(n12359), .ZN(n6845) );
  INV_X1 U8213 ( .A(n9103), .ZN(n7401) );
  AOI21_X1 U8214 ( .B1(n12222), .B2(n6848), .A(n6847), .ZN(n6846) );
  INV_X1 U8215 ( .A(n12225), .ZN(n6847) );
  INV_X1 U8216 ( .A(n12219), .ZN(n6848) );
  NOR2_X1 U8217 ( .A1(n9395), .A2(n9156), .ZN(n9170) );
  INV_X1 U8218 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8678) );
  INV_X1 U8219 ( .A(n7006), .ZN(n7005) );
  OAI21_X1 U8220 ( .B1(n8658), .B2(n7007), .A(n9027), .ZN(n7006) );
  INV_X1 U8221 ( .A(n8660), .ZN(n7007) );
  INV_X1 U8222 ( .A(n8654), .ZN(n7022) );
  OR2_X1 U8223 ( .A1(n12943), .A2(n7147), .ZN(n7146) );
  INV_X1 U8224 ( .A(n8099), .ZN(n7147) );
  NOR2_X1 U8225 ( .A1(n7155), .A2(n6667), .ZN(n6666) );
  INV_X1 U8226 ( .A(n7815), .ZN(n6667) );
  NAND2_X1 U8227 ( .A1(n7158), .A2(n7851), .ZN(n7155) );
  INV_X1 U8228 ( .A(n7156), .ZN(n7154) );
  NAND2_X1 U8229 ( .A1(n6666), .A2(n13029), .ZN(n6664) );
  XNOR2_X1 U8230 ( .A(n10274), .B(n8086), .ZN(n7644) );
  NOR2_X1 U8231 ( .A1(n8522), .A2(n8523), .ZN(n6771) );
  NAND2_X1 U8232 ( .A1(n8494), .A2(n8493), .ZN(n6773) );
  INV_X1 U8233 ( .A(n8537), .ZN(n7391) );
  INV_X1 U8234 ( .A(n8536), .ZN(n7390) );
  NOR2_X1 U8235 ( .A1(n6828), .A2(n6469), .ZN(n6827) );
  INV_X1 U8236 ( .A(n8459), .ZN(n6828) );
  NAND2_X1 U8237 ( .A1(n7377), .A2(n6474), .ZN(n7375) );
  NAND2_X1 U8238 ( .A1(n7140), .A2(n6467), .ZN(n7139) );
  OR2_X1 U8239 ( .A1(n8043), .A2(n8042), .ZN(n8067) );
  INV_X1 U8240 ( .A(n11530), .ZN(n7357) );
  OR2_X1 U8241 ( .A1(n7931), .A2(n7930), .ZN(n7952) );
  INV_X1 U8242 ( .A(n7211), .ZN(n7205) );
  INV_X1 U8243 ( .A(n10902), .ZN(n7359) );
  NOR2_X1 U8244 ( .A1(n7710), .A2(n7709), .ZN(n7731) );
  INV_X1 U8245 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7709) );
  NOR2_X1 U8246 ( .A1(n7638), .A2(n7637), .ZN(n7661) );
  AND2_X1 U8247 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7616) );
  NOR2_X1 U8248 ( .A1(n9727), .A2(n10073), .ZN(n9796) );
  NAND2_X1 U8249 ( .A1(n9786), .A2(n9791), .ZN(n9924) );
  INV_X1 U8250 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7500) );
  INV_X1 U8251 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7469) );
  NOR2_X1 U8252 ( .A1(n7743), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n7765) );
  OR2_X1 U8253 ( .A1(n7727), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n7743) );
  AND2_X1 U8254 ( .A1(n7545), .A2(n7141), .ZN(n7548) );
  INV_X1 U8255 ( .A(n11231), .ZN(n7281) );
  NAND2_X1 U8256 ( .A1(n11134), .A2(n6607), .ZN(n6606) );
  INV_X1 U8257 ( .A(n11130), .ZN(n6607) );
  INV_X1 U8258 ( .A(n10182), .ZN(n9300) );
  NAND2_X1 U8259 ( .A1(n11763), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n11798) );
  INV_X1 U8260 ( .A(n11765), .ZN(n11763) );
  NAND2_X1 U8261 ( .A1(n11720), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n11744) );
  INV_X1 U8262 ( .A(n11722), .ZN(n11720) );
  INV_X1 U8263 ( .A(n13849), .ZN(n6811) );
  NOR2_X1 U8264 ( .A1(n14001), .A2(n14149), .ZN(n6960) );
  NAND2_X1 U8265 ( .A1(n7296), .A2(n7295), .ZN(n7294) );
  INV_X1 U8266 ( .A(n7299), .ZN(n7295) );
  NOR2_X1 U8267 ( .A1(n11356), .A2(n11355), .ZN(n11614) );
  OR2_X1 U8268 ( .A1(n11309), .A2(n11308), .ZN(n11356) );
  AND2_X1 U8269 ( .A1(n11038), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n11288) );
  NAND2_X1 U8270 ( .A1(n10852), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10877) );
  NAND2_X1 U8271 ( .A1(n14815), .A2(n11139), .ZN(n6787) );
  AOI21_X1 U8272 ( .B1(n14724), .B2(n14719), .A(n10747), .ZN(n10790) );
  NAND2_X1 U8273 ( .A1(n6648), .A2(n7316), .ZN(n13921) );
  AOI21_X1 U8274 ( .B1(n7317), .B2(n13958), .A(n6578), .ZN(n7316) );
  NAND2_X1 U8275 ( .A1(n13959), .A2(n7317), .ZN(n6648) );
  NAND2_X1 U8276 ( .A1(n6640), .A2(n6499), .ZN(n14013) );
  NOR2_X1 U8277 ( .A1(n6962), .A2(n13686), .ZN(n6961) );
  INV_X1 U8278 ( .A(n6963), .ZN(n6962) );
  NAND2_X1 U8279 ( .A1(n8172), .A2(n8171), .ZN(n8177) );
  NAND2_X1 U8280 ( .A1(n8037), .A2(n8036), .ZN(n8057) );
  NAND2_X1 U8281 ( .A1(n6763), .A2(n7965), .ZN(n6759) );
  INV_X1 U8282 ( .A(n7252), .ZN(n7249) );
  NAND2_X1 U8283 ( .A1(n7874), .A2(n7873), .ZN(n6625) );
  INV_X1 U8284 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9210) );
  XNOR2_X1 U8285 ( .A(n7854), .B(n9568), .ZN(n7852) );
  NAND2_X1 U8286 ( .A1(n7242), .A2(n7816), .ZN(n7241) );
  INV_X1 U8287 ( .A(n7835), .ZN(n7242) );
  XNOR2_X1 U8288 ( .A(n7759), .B(SI_11_), .ZN(n7762) );
  AOI21_X1 U8289 ( .B1(n7676), .B2(n6770), .A(n6769), .ZN(n6768) );
  INV_X1 U8290 ( .A(n7672), .ZN(n6770) );
  INV_X1 U8291 ( .A(n7699), .ZN(n6769) );
  OAI21_X1 U8292 ( .B1(n6450), .B2(n9367), .A(n6697), .ZN(n7631) );
  NAND2_X1 U8293 ( .A1(n6436), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6697) );
  NAND2_X1 U8294 ( .A1(n6449), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6699) );
  INV_X1 U8295 ( .A(P1_RD_REG_SCAN_IN), .ZN(n6621) );
  INV_X1 U8296 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n6620) );
  INV_X1 U8297 ( .A(P2_RD_REG_SCAN_IN), .ZN(n6619) );
  AND2_X1 U8298 ( .A1(n8205), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7124) );
  INV_X1 U8299 ( .A(n8257), .ZN(n7125) );
  XNOR2_X1 U8300 ( .A(n8209), .B(n7117), .ZN(n8254) );
  AOI21_X1 U8301 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n8220), .A(n8219), .ZN(
        n8221) );
  NOR2_X1 U8302 ( .A1(n8252), .A2(n8251), .ZN(n8219) );
  OAI21_X1 U8303 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n14627), .A(n8230), .ZN(
        n8240) );
  INV_X1 U8304 ( .A(n12151), .ZN(n7098) );
  INV_X1 U8305 ( .A(n12130), .ZN(n7073) );
  NOR2_X1 U8306 ( .A1(n12154), .A2(n12156), .ZN(n12157) );
  INV_X1 U8307 ( .A(n12155), .ZN(n12156) );
  AND2_X1 U8308 ( .A1(n8699), .A2(n12469), .ZN(n8983) );
  NAND2_X1 U8309 ( .A1(n6556), .A2(n6859), .ZN(n6858) );
  NAND2_X1 U8310 ( .A1(n6860), .A2(n12397), .ZN(n6859) );
  OR2_X1 U8311 ( .A1(n8729), .A2(n6874), .ZN(n7045) );
  NAND2_X1 U8312 ( .A1(n6739), .A2(n6738), .ZN(n9864) );
  OR2_X1 U8313 ( .A1(n12646), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n6739) );
  NAND2_X1 U8314 ( .A1(n12646), .A2(n9828), .ZN(n6738) );
  NAND2_X1 U8315 ( .A1(n10545), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n6988) );
  OR2_X1 U8316 ( .A1(n14935), .A2(n10597), .ZN(n6873) );
  NOR2_X1 U8317 ( .A1(n14961), .A2(n10527), .ZN(n14976) );
  INV_X1 U8318 ( .A(n6884), .ZN(n10950) );
  XNOR2_X1 U8319 ( .A(n12586), .B(n12563), .ZN(n15019) );
  XNOR2_X1 U8320 ( .A(n12589), .B(n12605), .ZN(n15046) );
  NAND2_X1 U8321 ( .A1(n15079), .A2(n12592), .ZN(n15098) );
  INV_X1 U8322 ( .A(n15110), .ZN(n6757) );
  NAND2_X1 U8323 ( .A1(n6883), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n6882) );
  NAND2_X1 U8324 ( .A1(n12575), .A2(n6883), .ZN(n6881) );
  INV_X1 U8325 ( .A(n14432), .ZN(n6883) );
  XNOR2_X1 U8326 ( .A(n12596), .B(n14438), .ZN(n14440) );
  NAND2_X1 U8327 ( .A1(n14440), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n14439) );
  INV_X1 U8328 ( .A(n7405), .ZN(n7404) );
  OAI21_X1 U8329 ( .B1(n7409), .B2(n7406), .A(n6496), .ZN(n7405) );
  NAND2_X1 U8330 ( .A1(n12312), .A2(n12304), .ZN(n12724) );
  NAND2_X1 U8331 ( .A1(n9026), .A2(n12295), .ZN(n12734) );
  NAND2_X1 U8332 ( .A1(n6870), .A2(n6868), .ZN(n12759) );
  AOI21_X1 U8333 ( .B1(n12789), .B2(n6871), .A(n6869), .ZN(n6868) );
  NOR2_X1 U8334 ( .A1(n9002), .A2(n6872), .ZN(n6871) );
  OR2_X1 U8335 ( .A1(n8996), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9007) );
  OR2_X1 U8336 ( .A1(n12788), .A2(n12789), .ZN(n12786) );
  AND4_X1 U8337 ( .A1(n8989), .A2(n8988), .A3(n8987), .A4(n8986), .ZN(n12800)
         );
  NAND2_X1 U8338 ( .A1(n12813), .A2(n12271), .ZN(n12802) );
  AND2_X1 U8339 ( .A1(n12275), .A2(n12276), .ZN(n12801) );
  AOI21_X1 U8340 ( .B1(n7058), .B2(n7056), .A(n7055), .ZN(n7054) );
  INV_X1 U8341 ( .A(n12262), .ZN(n7056) );
  NAND2_X1 U8342 ( .A1(n8696), .A2(n8695), .ZN(n8946) );
  OR2_X1 U8343 ( .A1(n8896), .A2(n8692), .ZN(n8917) );
  AND2_X1 U8344 ( .A1(n7416), .A2(n7415), .ZN(n7414) );
  NAND2_X1 U8345 ( .A1(n7419), .A2(n7421), .ZN(n7415) );
  OR2_X1 U8346 ( .A1(n8822), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8853) );
  INV_X1 U8347 ( .A(n9104), .ZN(n7402) );
  AND2_X1 U8348 ( .A1(n7400), .A2(n9108), .ZN(n7399) );
  NAND2_X1 U8349 ( .A1(n9104), .A2(n7401), .ZN(n7400) );
  NAND2_X1 U8350 ( .A1(n11093), .A2(n12360), .ZN(n11092) );
  OAI21_X1 U8351 ( .B1(n10829), .B2(n12359), .A(n6846), .ZN(n11074) );
  NAND2_X1 U8352 ( .A1(n10831), .A2(n9103), .ZN(n10933) );
  NAND2_X1 U8353 ( .A1(n8690), .A2(n8689), .ZN(n8822) );
  INV_X1 U8354 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n8689) );
  INV_X1 U8355 ( .A(n8808), .ZN(n8690) );
  OR2_X1 U8356 ( .A1(n8794), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8808) );
  NAND2_X1 U8357 ( .A1(n10441), .A2(n9101), .ZN(n10620) );
  INV_X1 U8358 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n8687) );
  INV_X1 U8359 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10594) );
  INV_X1 U8360 ( .A(n7043), .ZN(n7042) );
  OAI22_X1 U8361 ( .A1(n8888), .A2(n9335), .B1(n9834), .B2(n10521), .ZN(n7043)
         );
  AND2_X1 U8362 ( .A1(n10049), .A2(n12327), .ZN(n12769) );
  NOR2_X1 U8363 ( .A1(n9880), .A2(n15144), .ZN(n10589) );
  NAND2_X1 U8364 ( .A1(n9186), .A2(n9185), .ZN(n9201) );
  OR2_X1 U8365 ( .A1(n9886), .A2(n9386), .ZN(n9880) );
  NAND2_X1 U8366 ( .A1(n8674), .A2(n8673), .ZN(n9181) );
  OAI21_X1 U8367 ( .B1(n9046), .B2(P1_DATAO_REG_24__SCAN_IN), .A(n8665), .ZN(
        n9056) );
  OR2_X1 U8368 ( .A1(n9056), .A2(n9055), .ZN(n9058) );
  INV_X1 U8369 ( .A(n7448), .ZN(n7443) );
  OR2_X1 U8370 ( .A1(n8599), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n9160) );
  NAND2_X1 U8371 ( .A1(n8649), .A2(n8648), .ZN(n8979) );
  NAND2_X1 U8372 ( .A1(n8966), .A2(n8647), .ZN(n8649) );
  NAND2_X1 U8373 ( .A1(n8680), .A2(n7108), .ZN(n8941) );
  NAND2_X1 U8374 ( .A1(n8911), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8640) );
  NAND2_X1 U8375 ( .A1(n7009), .A2(n7008), .ZN(n8908) );
  AOI21_X1 U8376 ( .B1(n7010), .B2(n7012), .A(n6589), .ZN(n7008) );
  INV_X1 U8377 ( .A(n7029), .ZN(n7028) );
  AOI21_X1 U8378 ( .B1(n7029), .B2(n7027), .A(n6553), .ZN(n7026) );
  AOI21_X1 U8379 ( .B1(n8622), .B2(n8623), .A(n6554), .ZN(n7029) );
  OR2_X1 U8380 ( .A1(n8828), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8829) );
  NOR2_X1 U8381 ( .A1(n8829), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8861) );
  AND2_X1 U8382 ( .A1(n8623), .A2(n8621), .ZN(n8802) );
  INV_X1 U8383 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7429) );
  INV_X1 U8384 ( .A(n7016), .ZN(n7015) );
  AOI21_X1 U8385 ( .B1(n7016), .B2(n7014), .A(n6552), .ZN(n7013) );
  XNOR2_X1 U8386 ( .A(n10137), .B(P1_DATAO_REG_4__SCAN_IN), .ZN(n8770) );
  AND2_X1 U8387 ( .A1(n9369), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8615) );
  NAND2_X1 U8388 ( .A1(n8002), .A2(n8001), .ZN(n8018) );
  INV_X1 U8389 ( .A(n6659), .ZN(n6654) );
  INV_X1 U8390 ( .A(n13013), .ZN(n6674) );
  NOR2_X1 U8391 ( .A1(n6674), .A2(n6675), .ZN(n6672) );
  INV_X1 U8392 ( .A(n12948), .ZN(n6675) );
  AND2_X1 U8393 ( .A1(n12121), .A2(n7755), .ZN(n6680) );
  NAND2_X1 U8394 ( .A1(n7160), .A2(n10208), .ZN(n12119) );
  XNOR2_X1 U8395 ( .A(n12126), .B(n8086), .ZN(n12094) );
  NAND2_X1 U8396 ( .A1(n7748), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7776) );
  XNOR2_X1 U8397 ( .A(n8312), .B(n7590), .ZN(n9943) );
  NAND2_X1 U8398 ( .A1(n7912), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7931) );
  INV_X1 U8399 ( .A(n7913), .ZN(n7912) );
  NAND2_X1 U8400 ( .A1(n8080), .A2(n7148), .ZN(n13062) );
  NAND2_X1 U8401 ( .A1(n7841), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7886) );
  INV_X1 U8402 ( .A(n6704), .ZN(n8480) );
  BUF_X1 U8404 ( .A(n7591), .Z(n8186) );
  NOR2_X1 U8405 ( .A1(n10372), .A2(n6973), .ZN(n10376) );
  AND2_X1 U8406 ( .A1(n10373), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6973) );
  NOR2_X1 U8407 ( .A1(n10375), .A2(n10376), .ZN(n10497) );
  NOR2_X1 U8408 ( .A1(n6974), .A2(n10497), .ZN(n10500) );
  AND2_X1 U8409 ( .A1(n10501), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6974) );
  NAND2_X1 U8410 ( .A1(n10500), .A2(n10499), .ZN(n11111) );
  OR2_X1 U8411 ( .A1(n7818), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n7837) );
  NOR2_X1 U8412 ( .A1(n14855), .A2(n6976), .ZN(n11115) );
  AND2_X1 U8413 ( .A1(n14861), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6976) );
  NOR2_X1 U8414 ( .A1(n11115), .A2(n11114), .ZN(n13147) );
  NOR2_X1 U8415 ( .A1(n13147), .A2(n6975), .ZN(n13162) );
  AND2_X1 U8416 ( .A1(n13148), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6975) );
  INV_X1 U8417 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n7485) );
  NAND2_X1 U8418 ( .A1(n13442), .A2(n11561), .ZN(n13250) );
  NAND2_X1 U8419 ( .A1(n13444), .A2(n13075), .ZN(n11561) );
  OAI21_X1 U8420 ( .B1(n13292), .B2(n7319), .A(n7318), .ZN(n13244) );
  INV_X1 U8421 ( .A(n7320), .ZN(n7319) );
  AOI21_X1 U8422 ( .B1(n7320), .B2(n7323), .A(n6472), .ZN(n7318) );
  NOR2_X1 U8423 ( .A1(n7325), .A2(n13270), .ZN(n7320) );
  AND2_X1 U8424 ( .A1(n8121), .A2(n8111), .ZN(n13266) );
  NAND2_X1 U8425 ( .A1(n6629), .A2(n11556), .ZN(n13275) );
  INV_X1 U8426 ( .A(n7218), .ZN(n7217) );
  NOR3_X1 U8427 ( .A1(n13340), .A2(n13465), .A3(n13462), .ZN(n13315) );
  NOR2_X1 U8428 ( .A1(n13340), .A2(n7139), .ZN(n13296) );
  AND2_X1 U8429 ( .A1(n13354), .A2(n11530), .ZN(n13335) );
  AOI21_X1 U8430 ( .B1(n6459), .B2(n7223), .A(n6507), .ZN(n7221) );
  INV_X1 U8431 ( .A(n7349), .ZN(n7348) );
  AOI21_X1 U8432 ( .B1(n7349), .B2(n7347), .A(n7346), .ZN(n7345) );
  INV_X1 U8433 ( .A(n11386), .ZN(n7347) );
  NAND2_X1 U8434 ( .A1(n7134), .A2(n7133), .ZN(n13410) );
  INV_X1 U8435 ( .A(n7134), .ZN(n11384) );
  INV_X1 U8436 ( .A(n14508), .ZN(n7135) );
  INV_X1 U8437 ( .A(n11149), .ZN(n6727) );
  NAND2_X1 U8438 ( .A1(n7138), .A2(n7137), .ZN(n10909) );
  INV_X1 U8439 ( .A(n7136), .ZN(n11151) );
  INV_X1 U8440 ( .A(n7341), .ZN(n7340) );
  NAND2_X1 U8441 ( .A1(n10428), .A2(n10427), .ZN(n10472) );
  NAND2_X1 U8442 ( .A1(n7131), .A2(n7130), .ZN(n10402) );
  NAND2_X1 U8443 ( .A1(n10395), .A2(n7343), .ZN(n10428) );
  NAND2_X1 U8444 ( .A1(n10395), .A2(n10394), .ZN(n10397) );
  INV_X1 U8445 ( .A(n10391), .ZN(n10284) );
  INV_X1 U8446 ( .A(n13051), .ZN(n13370) );
  AND2_X1 U8447 ( .A1(n9431), .A2(n8192), .ZN(n13372) );
  NAND2_X1 U8448 ( .A1(n9728), .A2(n9729), .ZN(n9727) );
  INV_X1 U8449 ( .A(n9582), .ZN(n7198) );
  NOR2_X1 U8450 ( .A1(n9462), .A2(n9998), .ZN(n7165) );
  INV_X1 U8451 ( .A(n7879), .ZN(n7499) );
  NAND2_X1 U8452 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n7475) );
  OR2_X1 U8453 ( .A1(n7612), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n7657) );
  OR2_X1 U8454 ( .A1(n7566), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n7584) );
  NAND2_X1 U8455 ( .A1(n13562), .A2(n7278), .ZN(n7276) );
  INV_X1 U8456 ( .A(n7277), .ZN(n7275) );
  OR2_X1 U8457 ( .A1(n10877), .A2(n10876), .ZN(n11007) );
  INV_X1 U8458 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n11006) );
  NOR2_X1 U8459 ( .A1(n11007), .A2(n11006), .ZN(n11038) );
  NOR2_X1 U8460 ( .A1(n11682), .A2(n13647), .ZN(n11702) );
  NAND2_X1 U8461 ( .A1(n11663), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11682) );
  OR2_X1 U8462 ( .A1(n11230), .A2(n11229), .ZN(n11231) );
  AND2_X1 U8463 ( .A1(n10187), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13664) );
  NAND2_X1 U8464 ( .A1(n12027), .A2(n12029), .ZN(n7254) );
  INV_X1 U8465 ( .A(n6909), .ZN(n6908) );
  NAND2_X1 U8466 ( .A1(n13722), .A2(n6714), .ZN(n9303) );
  NAND2_X1 U8467 ( .A1(n6715), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6714) );
  NAND2_X1 U8468 ( .A1(n6892), .A2(n6891), .ZN(n6890) );
  NAND2_X1 U8469 ( .A1(n6715), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6891) );
  NOR2_X1 U8470 ( .A1(n9741), .A2(n6900), .ZN(n13743) );
  AND2_X1 U8471 ( .A1(n10321), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6900) );
  NOR2_X1 U8472 ( .A1(n13743), .A2(n13742), .ZN(n13741) );
  NAND2_X1 U8473 ( .A1(n10351), .A2(n10350), .ZN(n13756) );
  NAND2_X1 U8474 ( .A1(n13756), .A2(n6894), .ZN(n13757) );
  OR2_X1 U8475 ( .A1(n13762), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6894) );
  NAND2_X1 U8476 ( .A1(n13757), .A2(n13758), .ZN(n13781) );
  NOR2_X1 U8477 ( .A1(n7179), .A2(n7178), .ZN(n7177) );
  INV_X1 U8478 ( .A(n7180), .ZN(n7178) );
  NAND2_X1 U8479 ( .A1(n13925), .A2(n14705), .ZN(n7314) );
  NAND2_X1 U8480 ( .A1(n6960), .A2(n6959), .ZN(n13969) );
  INV_X1 U8481 ( .A(n6960), .ZN(n13986) );
  OAI21_X1 U8482 ( .B1(n14161), .B2(n14040), .A(n14159), .ZN(n13998) );
  NAND2_X1 U8483 ( .A1(n6792), .A2(n6791), .ZN(n14044) );
  AOI21_X1 U8484 ( .B1(n6793), .B2(n6797), .A(n6579), .ZN(n6791) );
  NAND2_X1 U8485 ( .A1(n6644), .A2(n11950), .ZN(n11306) );
  NOR2_X1 U8486 ( .A1(n11304), .A2(n6646), .ZN(n6645) );
  INV_X1 U8487 ( .A(n11302), .ZN(n6646) );
  NAND2_X1 U8488 ( .A1(n11029), .A2(n6963), .ZN(n14092) );
  NAND2_X1 U8489 ( .A1(n11029), .A2(n14544), .ZN(n14091) );
  INV_X1 U8490 ( .A(n7309), .ZN(n7308) );
  AOI21_X1 U8491 ( .B1(n12043), .B2(n10886), .A(n6516), .ZN(n7309) );
  OR2_X1 U8492 ( .A1(n10732), .A2(n10731), .ZN(n10758) );
  OR2_X1 U8493 ( .A1(n10333), .A2(n10332), .ZN(n10732) );
  NOR2_X1 U8494 ( .A1(n6956), .A2(n14712), .ZN(n6954) );
  NAND2_X1 U8495 ( .A1(n14736), .A2(n14785), .ZN(n14735) );
  NAND2_X1 U8496 ( .A1(n14736), .A2(n6955), .ZN(n14713) );
  OAI211_X1 U8497 ( .C1(n10766), .C2(n7304), .A(n7301), .B(n12038), .ZN(n10797) );
  NOR2_X1 U8498 ( .A1(n7304), .A2(n7305), .ZN(n7302) );
  NOR2_X1 U8499 ( .A1(n10172), .A2(n10171), .ZN(n10233) );
  NAND2_X1 U8500 ( .A1(n6638), .A2(n12035), .ZN(n14746) );
  NAND2_X1 U8501 ( .A1(n14743), .A2(n14741), .ZN(n6638) );
  AND4_X2 U8502 ( .A1(n9611), .A2(n9610), .A3(n9609), .A4(n9608), .ZN(n13581)
         );
  OR2_X1 U8503 ( .A1(n10225), .A2(n9517), .ZN(n10791) );
  NAND2_X1 U8504 ( .A1(n9601), .A2(n11853), .ZN(n11867) );
  AND2_X1 U8505 ( .A1(n11852), .A2(n11851), .ZN(n14103) );
  OR2_X1 U8506 ( .A1(n13917), .A2(n13916), .ZN(n14127) );
  NAND2_X1 U8507 ( .A1(n11303), .A2(n11302), .ZN(n14083) );
  NAND2_X1 U8508 ( .A1(n11284), .A2(n7185), .ZN(n14077) );
  INV_X1 U8509 ( .A(n11895), .ZN(n14781) );
  OAI211_X1 U8510 ( .C1(n6953), .C2(n6952), .A(n6951), .B(n14756), .ZN(n14767)
         );
  INV_X1 U8511 ( .A(n14757), .ZN(n6951) );
  INV_X1 U8512 ( .A(n11090), .ZN(n9406) );
  NOR2_X1 U8513 ( .A1(n8500), .A2(n8499), .ZN(n6775) );
  INV_X1 U8514 ( .A(n8504), .ZN(n6776) );
  INV_X1 U8515 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7176) );
  INV_X1 U8516 ( .A(n8169), .ZN(n8106) );
  XNOR2_X1 U8517 ( .A(n9222), .B(n9221), .ZN(n10181) );
  OR2_X1 U8518 ( .A1(n9591), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n10083) );
  NAND2_X1 U8519 ( .A1(n7817), .A2(n7816), .ZN(n7836) );
  NAND2_X1 U8520 ( .A1(n6914), .A2(n6913), .ZN(n7790) );
  AND2_X1 U8521 ( .A1(n6626), .A2(n7243), .ZN(n6913) );
  OAI21_X1 U8522 ( .B1(n7725), .B2(n7247), .A(n7245), .ZN(n7787) );
  OAI21_X1 U8523 ( .B1(n6630), .B2(SI_10_), .A(n7741), .ZN(n7723) );
  NAND2_X1 U8524 ( .A1(n7725), .A2(n7724), .ZN(n7742) );
  NAND2_X1 U8525 ( .A1(n6450), .A2(n8608), .ZN(n6726) );
  INV_X1 U8526 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n8261) );
  NOR2_X1 U8527 ( .A1(n8212), .A2(n8211), .ZN(n8272) );
  NOR2_X1 U8528 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n8253), .ZN(n8211) );
  OAI21_X1 U8529 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n8225), .A(n8224), .ZN(
        n8247) );
  INV_X1 U8530 ( .A(n12551), .ZN(n11184) );
  NAND2_X1 U8531 ( .A1(n6721), .A2(n11472), .ZN(n12131) );
  NAND2_X1 U8532 ( .A1(n9039), .A2(n9038), .ZN(n12725) );
  NAND2_X1 U8533 ( .A1(n7105), .A2(n7106), .ZN(n11413) );
  INV_X1 U8534 ( .A(n7104), .ZN(n7106) );
  NAND2_X1 U8535 ( .A1(n7084), .A2(n7089), .ZN(n10452) );
  NAND2_X1 U8536 ( .A1(n7086), .A2(n7085), .ZN(n7084) );
  NAND2_X1 U8537 ( .A1(n8995), .A2(n8994), .ZN(n12439) );
  AND4_X1 U8538 ( .A1(n8860), .A2(n8859), .A3(n8858), .A4(n8857), .ZN(n11257)
         );
  OR2_X1 U8539 ( .A1(n11050), .A2(n11081), .ZN(n11051) );
  INV_X1 U8540 ( .A(n12505), .ZN(n12525) );
  NAND2_X1 U8541 ( .A1(n12557), .A2(n7094), .ZN(n7093) );
  NAND2_X1 U8542 ( .A1(n9018), .A2(n9017), .ZN(n12750) );
  NAND2_X1 U8543 ( .A1(n7076), .A2(n12164), .ZN(n12449) );
  NAND2_X1 U8544 ( .A1(n12475), .A2(n12476), .ZN(n7076) );
  NAND2_X1 U8545 ( .A1(n7085), .A2(n7088), .ZN(n7081) );
  OR2_X1 U8546 ( .A1(n8888), .A2(n9332), .ZN(n8727) );
  NAND2_X1 U8547 ( .A1(n7100), .A2(n7099), .ZN(n12485) );
  INV_X1 U8548 ( .A(n12484), .ZN(n7100) );
  NAND2_X1 U8549 ( .A1(n7103), .A2(n7102), .ZN(n7101) );
  INV_X1 U8550 ( .A(n11417), .ZN(n7103) );
  OR2_X1 U8551 ( .A1(n10050), .A2(n10049), .ZN(n12505) );
  NOR2_X1 U8552 ( .A1(n12143), .A2(n6522), .ZN(n12500) );
  NOR2_X1 U8553 ( .A1(n12467), .A2(n12140), .ZN(n12143) );
  AND2_X1 U8554 ( .A1(n9898), .A2(n9897), .ZN(n12461) );
  INV_X1 U8555 ( .A(n12534), .ZN(n12499) );
  AND2_X1 U8556 ( .A1(n9094), .A2(n9093), .ZN(n12676) );
  AOI21_X1 U8557 ( .B1(n7077), .B2(n7079), .A(n6513), .ZN(n7074) );
  INV_X1 U8558 ( .A(n12528), .ZN(n12515) );
  INV_X1 U8559 ( .A(n12461), .ZN(n12531) );
  AND2_X1 U8560 ( .A1(n12353), .A2(n9129), .ZN(n12185) );
  INV_X1 U8561 ( .A(n12453), .ZN(n12691) );
  INV_X1 U8562 ( .A(n12677), .ZN(n12707) );
  INV_X1 U8563 ( .A(n12694), .ZN(n12720) );
  INV_X1 U8564 ( .A(n12746), .ZN(n12770) );
  INV_X1 U8565 ( .A(n11423), .ZN(n12548) );
  INV_X1 U8566 ( .A(n11257), .ZN(n12234) );
  INV_X1 U8567 ( .A(n10921), .ZN(n12553) );
  INV_X1 U8568 ( .A(P3_U3897), .ZN(n12558) );
  NAND2_X1 U8569 ( .A1(n8753), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8722) );
  NOR2_X1 U8570 ( .A1(n9903), .A2(n9902), .ZN(n9905) );
  INV_X1 U8571 ( .A(n6989), .ZN(n10531) );
  OAI21_X1 U8572 ( .B1(n6987), .B2(n14939), .A(n6986), .ZN(n14935) );
  INV_X1 U8573 ( .A(n6873), .ZN(n14934) );
  INV_X1 U8574 ( .A(n6993), .ZN(n14993) );
  NAND2_X1 U8575 ( .A1(n14987), .A2(n6577), .ZN(n10962) );
  AND2_X1 U8576 ( .A1(n9850), .A2(n9842), .ZN(n14960) );
  NAND2_X1 U8577 ( .A1(n6877), .A2(n6876), .ZN(n15024) );
  NAND2_X1 U8578 ( .A1(n6747), .A2(n6748), .ZN(n15034) );
  AOI21_X1 U8579 ( .B1(n15013), .B2(n15011), .A(n6752), .ZN(n15036) );
  NAND2_X1 U8580 ( .A1(n6477), .A2(n6996), .ZN(n6995) );
  AND2_X1 U8581 ( .A1(n15052), .A2(n12619), .ZN(n15073) );
  INV_X1 U8582 ( .A(n6985), .ZN(n12571) );
  NAND2_X1 U8583 ( .A1(n15087), .A2(n12631), .ZN(n15111) );
  NAND2_X1 U8584 ( .A1(n15087), .A2(n6478), .ZN(n15112) );
  NOR2_X1 U8585 ( .A1(n14404), .A2(n14405), .ZN(n14403) );
  NAND2_X1 U8586 ( .A1(n6878), .A2(n14960), .ZN(n14467) );
  NAND2_X1 U8587 ( .A1(n6880), .A2(n14464), .ZN(n6878) );
  NAND2_X1 U8588 ( .A1(n14466), .A2(n14465), .ZN(n6880) );
  INV_X1 U8589 ( .A(n6991), .ZN(n14466) );
  NAND2_X1 U8590 ( .A1(n14464), .A2(n12580), .ZN(n12582) );
  NOR2_X1 U8591 ( .A1(n14457), .A2(n6742), .ZN(n12650) );
  AND2_X1 U8592 ( .A1(n9850), .A2(n12646), .ZN(n15107) );
  NAND2_X1 U8593 ( .A1(n12335), .A2(n12334), .ZN(n14475) );
  NAND2_X1 U8594 ( .A1(n6857), .A2(n6861), .ZN(n12398) );
  NAND2_X1 U8595 ( .A1(n7431), .A2(n7430), .ZN(n9187) );
  AND2_X1 U8596 ( .A1(n11509), .A2(n11508), .ZN(n12086) );
  NAND2_X1 U8597 ( .A1(n9085), .A2(n9084), .ZN(n12170) );
  OR2_X1 U8598 ( .A1(n12333), .A2(n11332), .ZN(n9084) );
  NAND2_X1 U8599 ( .A1(n12710), .A2(n12310), .ZN(n12697) );
  NAND2_X1 U8600 ( .A1(n7403), .A2(n7409), .ZN(n12731) );
  OR2_X1 U8601 ( .A1(n12756), .A2(n7411), .ZN(n7403) );
  NAND2_X1 U8602 ( .A1(n7413), .A2(n7412), .ZN(n12742) );
  NAND2_X1 U8603 ( .A1(n7432), .A2(n7435), .ZN(n12809) );
  NAND2_X1 U8604 ( .A1(n11439), .A2(n7437), .ZN(n7432) );
  AOI21_X1 U8605 ( .B1(n11439), .B2(n12376), .A(n7438), .ZN(n11462) );
  NAND2_X1 U8606 ( .A1(n7057), .A2(n12262), .ZN(n11465) );
  OR2_X1 U8607 ( .A1(n11438), .A2(n8936), .ZN(n7057) );
  NAND2_X1 U8608 ( .A1(n7050), .A2(n7051), .ZN(n11375) );
  NAND2_X1 U8609 ( .A1(n11247), .A2(n12247), .ZN(n11223) );
  NAND2_X1 U8610 ( .A1(n11064), .A2(n9110), .ZN(n11243) );
  NAND2_X1 U8611 ( .A1(n10932), .A2(n12222), .ZN(n10931) );
  NAND2_X1 U8612 ( .A1(n10829), .A2(n12219), .ZN(n10932) );
  AND2_X1 U8613 ( .A1(n12818), .A2(n10590), .ZN(n12821) );
  NAND2_X1 U8614 ( .A1(n10593), .A2(n10592), .ZN(n12815) );
  INV_X2 U8615 ( .A(n12818), .ZN(n15136) );
  NOR2_X1 U8616 ( .A1(n12660), .A2(n12659), .ZN(n14474) );
  INV_X1 U8617 ( .A(n9201), .ZN(n12422) );
  AND2_X1 U8618 ( .A1(n9071), .A2(n9070), .ZN(n12884) );
  NAND2_X1 U8619 ( .A1(n8971), .A2(n8970), .ZN(n12918) );
  AND2_X1 U8620 ( .A1(n8958), .A2(n8957), .ZN(n12922) );
  INV_X2 U8621 ( .A(n15157), .ZN(n15158) );
  OR2_X1 U8622 ( .A1(n15157), .A2(n15144), .ZN(n12926) );
  OAI21_X1 U8623 ( .B1(n9395), .B2(P3_D_REG_1__SCAN_IN), .A(n9144), .ZN(n10584) );
  INV_X1 U8624 ( .A(n9386), .ZN(n9423) );
  INV_X1 U8625 ( .A(n8715), .ZN(n12935) );
  NAND2_X1 U8626 ( .A1(n7004), .A2(n8660), .ZN(n9028) );
  NAND2_X1 U8627 ( .A1(n8659), .A2(n8658), .ZN(n7004) );
  NAND2_X1 U8628 ( .A1(n7023), .A2(n8654), .ZN(n9004) );
  NAND2_X1 U8629 ( .A1(n7025), .A2(n7024), .ZN(n7023) );
  NAND2_X1 U8630 ( .A1(n8597), .A2(n8599), .ZN(n10196) );
  INV_X1 U8631 ( .A(SI_19_), .ZN(n10012) );
  INV_X1 U8632 ( .A(SI_17_), .ZN(n9757) );
  INV_X1 U8633 ( .A(SI_16_), .ZN(n9647) );
  INV_X1 U8634 ( .A(SI_15_), .ZN(n9568) );
  NAND2_X1 U8635 ( .A1(n7035), .A2(n7033), .ZN(n8940) );
  NAND2_X1 U8636 ( .A1(n7035), .A2(n8642), .ZN(n8938) );
  INV_X1 U8637 ( .A(SI_14_), .ZN(n14351) );
  INV_X1 U8638 ( .A(SI_12_), .ZN(n14350) );
  OR2_X1 U8639 ( .A1(n8906), .A2(n8905), .ZN(n15068) );
  INV_X1 U8640 ( .A(SI_11_), .ZN(n9384) );
  NAND2_X1 U8641 ( .A1(n8846), .A2(n8632), .ZN(n8887) );
  INV_X1 U8642 ( .A(n10542), .ZN(n14967) );
  AND2_X1 U8643 ( .A1(n9430), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14905) );
  NAND2_X1 U8644 ( .A1(n13062), .A2(n8099), .ZN(n12942) );
  XNOR2_X1 U8645 ( .A(n8018), .B(n8016), .ZN(n12949) );
  OR2_X1 U8646 ( .A1(n12120), .A2(n7739), .ZN(n7740) );
  NAND2_X1 U8647 ( .A1(n10208), .A2(n7720), .ZN(n12963) );
  NAND2_X1 U8648 ( .A1(n8080), .A2(n6659), .ZN(n6651) );
  INV_X1 U8649 ( .A(n13066), .ZN(n13054) );
  INV_X1 U8650 ( .A(n13021), .ZN(n6676) );
  NAND2_X1 U8651 ( .A1(n6671), .A2(n6669), .ZN(n12995) );
  INV_X1 U8652 ( .A(n6670), .ZN(n6669) );
  NAND2_X1 U8653 ( .A1(n12949), .A2(n6672), .ZN(n6671) );
  OAI21_X1 U8654 ( .B1(n8019), .B2(n6674), .A(n8054), .ZN(n6670) );
  NAND2_X1 U8655 ( .A1(n7624), .A2(n9970), .ZN(n9979) );
  NAND2_X1 U8656 ( .A1(n9988), .A2(n7600), .ZN(n7624) );
  NAND2_X1 U8657 ( .A1(n7893), .A2(n13006), .ZN(n13012) );
  NAND2_X1 U8658 ( .A1(n6673), .A2(n8019), .ZN(n13014) );
  NAND2_X1 U8659 ( .A1(n12949), .A2(n12948), .ZN(n6673) );
  XNOR2_X1 U8660 ( .A(n8053), .B(n8051), .ZN(n13013) );
  XNOR2_X1 U8661 ( .A(n9969), .B(n7598), .ZN(n9989) );
  NAND2_X1 U8662 ( .A1(n9990), .A2(n7597), .ZN(n9988) );
  AND2_X1 U8663 ( .A1(n9989), .A2(n7596), .ZN(n7597) );
  AND2_X1 U8664 ( .A1(n8181), .A2(n8166), .ZN(n14523) );
  NAND2_X1 U8665 ( .A1(n10031), .A2(n7695), .ZN(n12968) );
  NAND2_X1 U8666 ( .A1(n6701), .A2(n8050), .ZN(n9859) );
  INV_X1 U8667 ( .A(n6677), .ZN(n13022) );
  NAND2_X1 U8668 ( .A1(n6668), .A2(n7814), .ZN(n13031) );
  NAND2_X1 U8669 ( .A1(n13012), .A2(n7897), .ZN(n13057) );
  NAND2_X1 U8670 ( .A1(n9979), .A2(n7628), .ZN(n10092) );
  NAND2_X1 U8671 ( .A1(n8080), .A2(n8079), .ZN(n13064) );
  NAND2_X1 U8672 ( .A1(n14504), .A2(n7831), .ZN(n9233) );
  NOR2_X1 U8673 ( .A1(n8539), .A2(n7459), .ZN(n8546) );
  NAND2_X1 U8674 ( .A1(n7571), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7353) );
  NAND2_X1 U8675 ( .A1(n8069), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7352) );
  AND2_X1 U8676 ( .A1(n7525), .A2(n7524), .ZN(n6693) );
  AND2_X1 U8677 ( .A1(n9427), .A2(n6565), .ZN(n9527) );
  NOR2_X1 U8678 ( .A1(n6978), .A2(n9527), .ZN(n9530) );
  NOR2_X1 U8679 ( .A1(n9526), .A2(n6979), .ZN(n6978) );
  INV_X1 U8680 ( .A(n6972), .ZN(n13115) );
  INV_X1 U8681 ( .A(n6970), .ZN(n13130) );
  NAND2_X1 U8682 ( .A1(n13142), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6969) );
  NOR2_X1 U8683 ( .A1(n9802), .A2(n6584), .ZN(n9805) );
  NAND2_X1 U8684 ( .A1(n9805), .A2(n9804), .ZN(n10116) );
  XNOR2_X1 U8685 ( .A(n13162), .B(n13168), .ZN(n13149) );
  INV_X1 U8686 ( .A(n7128), .ZN(n13236) );
  NAND2_X1 U8687 ( .A1(n8180), .A2(n8179), .ZN(n13438) );
  NAND2_X1 U8688 ( .A1(n7321), .A2(n7324), .ZN(n13260) );
  OAI21_X1 U8689 ( .B1(n13292), .B2(n13289), .A(n6480), .ZN(n13277) );
  NAND2_X1 U8690 ( .A1(n13309), .A2(n11554), .ZN(n13290) );
  NAND2_X1 U8691 ( .A1(n7232), .A2(n7231), .ZN(n13349) );
  AND2_X1 U8692 ( .A1(n7232), .A2(n6504), .ZN(n13346) );
  AND2_X1 U8693 ( .A1(n11548), .A2(n11547), .ZN(n13353) );
  NAND2_X1 U8694 ( .A1(n7351), .A2(n7349), .ZN(n11524) );
  NAND2_X1 U8695 ( .A1(n7351), .A2(n11388), .ZN(n11390) );
  NAND2_X1 U8696 ( .A1(n13503), .A2(n11382), .ZN(n11543) );
  NAND2_X1 U8697 ( .A1(n11211), .A2(n11201), .ZN(n13503) );
  INV_X1 U8698 ( .A(n11211), .ZN(n11213) );
  NAND2_X1 U8699 ( .A1(n7202), .A2(n7207), .ZN(n11268) );
  NAND2_X1 U8700 ( .A1(n11144), .A2(n7211), .ZN(n7202) );
  NAND2_X1 U8701 ( .A1(n7206), .A2(n7213), .ZN(n11210) );
  OR2_X1 U8702 ( .A1(n11144), .A2(n11143), .ZN(n7206) );
  NAND2_X1 U8703 ( .A1(n10903), .A2(n10902), .ZN(n11145) );
  NAND2_X1 U8704 ( .A1(n7224), .A2(n7225), .ZN(n10905) );
  NAND2_X1 U8705 ( .A1(n7226), .A2(n7229), .ZN(n10668) );
  NAND2_X1 U8706 ( .A1(n7228), .A2(n7227), .ZN(n7226) );
  NAND2_X1 U8707 ( .A1(n10015), .A2(n10014), .ZN(n10016) );
  INV_X1 U8708 ( .A(n9728), .ZN(n9627) );
  INV_X1 U8709 ( .A(n13424), .ZN(n13325) );
  INV_X1 U8710 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n7337) );
  OR2_X1 U8711 ( .A1(n13470), .A2(n13469), .ZN(n13529) );
  NAND3_X1 U8712 ( .A1(n9996), .A2(n9642), .A3(n9641), .ZN(n14928) );
  NOR2_X1 U8713 ( .A1(n7497), .A2(n6840), .ZN(n6838) );
  NAND2_X1 U8714 ( .A1(n7518), .A2(n7521), .ZN(n6840) );
  CLKBUF_X1 U8715 ( .A(n13548), .Z(n6698) );
  NAND2_X1 U8716 ( .A1(n8145), .A2(n8144), .ZN(n11338) );
  OR2_X1 U8717 ( .A1(n8148), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n8144) );
  XNOR2_X1 U8718 ( .A(n8151), .B(n8150), .ZN(n11087) );
  OAI21_X1 U8719 ( .B1(n8157), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8151) );
  INV_X1 U8720 ( .A(n7517), .ZN(n11099) );
  AOI21_X1 U8721 ( .B1(n7482), .B2(n7481), .A(n7480), .ZN(n6650) );
  INV_X1 U8722 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10944) );
  INV_X1 U8723 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10217) );
  INV_X1 U8724 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9454) );
  INV_X1 U8725 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9404) );
  INV_X1 U8726 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9387) );
  INV_X1 U8727 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9378) );
  INV_X1 U8728 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9373) );
  INV_X1 U8729 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9370) );
  INV_X1 U8730 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9355) );
  AND4_X1 U8731 ( .A1(n11294), .A2(n11293), .A3(n11292), .A4(n11291), .ZN(
        n14085) );
  NOR2_X1 U8732 ( .A1(n13562), .A2(n13563), .ZN(n13671) );
  NAND2_X1 U8733 ( .A1(n13642), .A2(n11696), .ZN(n13569) );
  NAND2_X1 U8734 ( .A1(n11135), .A2(n11134), .ZN(n11232) );
  NAND2_X1 U8735 ( .A1(n10157), .A2(n10156), .ZN(n13579) );
  INV_X1 U8736 ( .A(n13577), .ZN(n10156) );
  INV_X1 U8737 ( .A(n14683), .ZN(n11139) );
  AND2_X1 U8738 ( .A1(n9693), .A2(n9694), .ZN(n9704) );
  INV_X1 U8739 ( .A(n9691), .ZN(n9692) );
  NAND2_X1 U8740 ( .A1(n13634), .A2(n11658), .ZN(n13595) );
  NAND2_X1 U8741 ( .A1(n11662), .A2(n11661), .ZN(n14154) );
  NAND2_X1 U8742 ( .A1(n7276), .A2(n7277), .ZN(n13611) );
  OAI21_X1 U8743 ( .B1(n13642), .B2(n6612), .A(n6609), .ZN(n13626) );
  INV_X1 U8744 ( .A(n13570), .ZN(n6612) );
  INV_X1 U8745 ( .A(n7270), .ZN(n7269) );
  NAND2_X1 U8746 ( .A1(n10219), .A2(n10166), .ZN(n10167) );
  AND2_X1 U8747 ( .A1(n10982), .A2(n7289), .ZN(n7285) );
  AND2_X1 U8748 ( .A1(n7286), .A2(n7289), .ZN(n10983) );
  NAND2_X1 U8749 ( .A1(n11456), .A2(n11455), .ZN(n11583) );
  NAND2_X1 U8750 ( .A1(n13593), .A2(n11677), .ZN(n13643) );
  INV_X1 U8751 ( .A(n7279), .ZN(n11396) );
  NAND2_X1 U8752 ( .A1(n11232), .A2(n11231), .ZN(n11233) );
  OAI22_X1 U8753 ( .A1(n6487), .A2(n13619), .B1(n11609), .B2(n11608), .ZN(
        n13653) );
  NAND2_X1 U8754 ( .A1(n11758), .A2(n11757), .ZN(n13660) );
  AND2_X1 U8755 ( .A1(n10826), .A2(n14792), .ZN(n13685) );
  NAND2_X1 U8756 ( .A1(n9684), .A2(n9682), .ZN(n13688) );
  AND2_X1 U8757 ( .A1(n9707), .A2(n9678), .ZN(n14705) );
  NOR2_X1 U8758 ( .A1(n9681), .A2(n10184), .ZN(n12081) );
  OR2_X1 U8759 ( .A1(n11618), .A2(n11617), .ZN(n14065) );
  INV_X1 U8760 ( .A(n14052), .ZN(n13844) );
  NAND2_X1 U8761 ( .A1(n11814), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9524) );
  NAND2_X1 U8762 ( .A1(n6470), .A2(n14367), .ZN(n6926) );
  AND2_X1 U8763 ( .A1(n6925), .A2(n6924), .ZN(n6923) );
  INV_X1 U8764 ( .A(n6892), .ZN(n13718) );
  AND2_X1 U8765 ( .A1(n6890), .A2(n6889), .ZN(n9482) );
  INV_X1 U8766 ( .A(n9308), .ZN(n6889) );
  INV_X1 U8767 ( .A(n6890), .ZN(n9309) );
  NAND2_X1 U8768 ( .A1(n13735), .A2(n6533), .ZN(n9491) );
  NAND2_X1 U8769 ( .A1(n9491), .A2(n9492), .ZN(n9745) );
  NOR2_X1 U8770 ( .A1(n13741), .A2(n6899), .ZN(n9744) );
  AND2_X1 U8771 ( .A1(n13748), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6899) );
  NAND2_X1 U8772 ( .A1(n9744), .A2(n9743), .ZN(n9957) );
  AND2_X1 U8773 ( .A1(n9817), .A2(n9653), .ZN(n14610) );
  NOR2_X1 U8774 ( .A1(n14605), .A2(n6888), .ZN(n14615) );
  AND2_X1 U8775 ( .A1(n14610), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6888) );
  INV_X1 U8776 ( .A(n13784), .ZN(n13785) );
  INV_X1 U8777 ( .A(n14665), .ZN(n14636) );
  INV_X1 U8778 ( .A(n13808), .ZN(n13807) );
  NAND2_X1 U8779 ( .A1(n6807), .A2(n6809), .ZN(n13937) );
  NAND2_X1 U8780 ( .A1(n13963), .A2(n7317), .ZN(n13932) );
  NAND2_X1 U8781 ( .A1(n13854), .A2(n7188), .ZN(n13951) );
  NAND2_X1 U8782 ( .A1(n13854), .A2(n13853), .ZN(n13968) );
  NAND2_X1 U8783 ( .A1(n7292), .A2(n7296), .ZN(n14051) );
  NAND2_X1 U8784 ( .A1(n11353), .A2(n7299), .ZN(n7292) );
  NAND2_X1 U8785 ( .A1(n13815), .A2(n13814), .ZN(n14062) );
  NAND2_X1 U8786 ( .A1(n6794), .A2(n6795), .ZN(n14060) );
  OR2_X1 U8787 ( .A1(n11341), .A2(n6797), .ZN(n6794) );
  NAND2_X1 U8788 ( .A1(n11341), .A2(n11340), .ZN(n13842) );
  NAND2_X1 U8789 ( .A1(n11344), .A2(n11343), .ZN(n13843) );
  AND2_X1 U8790 ( .A1(n7184), .A2(n7183), .ZN(n11295) );
  AND2_X1 U8791 ( .A1(n6789), .A2(n6790), .ZN(n11002) );
  NAND2_X1 U8792 ( .A1(n10887), .A2(n10886), .ZN(n11003) );
  NAND2_X1 U8793 ( .A1(n7168), .A2(n7167), .ZN(n10998) );
  NAND2_X1 U8794 ( .A1(n6786), .A2(n10755), .ZN(n10756) );
  NAND2_X1 U8795 ( .A1(n14687), .A2(n10754), .ZN(n6786) );
  OR2_X1 U8796 ( .A1(n6442), .A2(n10662), .ZN(n14047) );
  OR2_X1 U8797 ( .A1(n6442), .A2(n12058), .ZN(n14695) );
  INV_X1 U8798 ( .A(n14047), .ZN(n14754) );
  NAND2_X2 U8799 ( .A1(n9686), .A2(n9685), .ZN(n14751) );
  AND2_X1 U8800 ( .A1(n14110), .A2(n14111), .ZN(n6725) );
  NAND2_X1 U8801 ( .A1(n14117), .A2(n6694), .ZN(n14202) );
  NAND2_X1 U8802 ( .A1(n6696), .A2(n14824), .ZN(n6695) );
  OAI21_X1 U8803 ( .B1(n6493), .B2(n14826), .A(n6803), .ZN(n6800) );
  NAND2_X1 U8804 ( .A1(n6488), .A2(n13893), .ZN(n14119) );
  AND2_X1 U8805 ( .A1(n14827), .A2(n14749), .ZN(n6798) );
  OR4_X1 U8806 ( .A1(n14165), .A2(n14164), .A3(n14163), .A4(n14162), .ZN(
        n14210) );
  NAND2_X1 U8807 ( .A1(n10181), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9407) );
  OAI21_X1 U8808 ( .B1(n10312), .B2(n9268), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9270) );
  NAND2_X1 U8809 ( .A1(n9245), .A2(n7453), .ZN(n9268) );
  XNOR2_X1 U8810 ( .A(n6618), .B(P1_IR_REG_26__SCAN_IN), .ZN(n11334) );
  OAI21_X1 U8811 ( .B1(n9230), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6618) );
  OR2_X1 U8812 ( .A1(n9255), .A2(n9220), .ZN(n9259) );
  NOR2_X1 U8813 ( .A1(n9257), .A2(n9256), .ZN(n9258) );
  INV_X1 U8814 ( .A(n9602), .ZN(n11853) );
  INV_X1 U8815 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10942) );
  INV_X1 U8816 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10513) );
  NAND2_X1 U8817 ( .A1(n7925), .A2(n7262), .ZN(n7906) );
  INV_X1 U8818 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10086) );
  INV_X1 U8819 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9419) );
  NOR2_X1 U8820 ( .A1(n9418), .A2(n9417), .ZN(n14597) );
  INV_X1 U8821 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9403) );
  INV_X1 U8822 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9381) );
  NAND2_X1 U8823 ( .A1(n7630), .A2(n6682), .ZN(n6681) );
  NOR2_X1 U8824 ( .A1(n7633), .A2(n6901), .ZN(n6682) );
  INV_X1 U8825 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9364) );
  INV_X1 U8826 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10147) );
  MUX2_X1 U8827 ( .A(n14216), .B(n9294), .S(P1_IR_REG_2__SCAN_IN), .Z(n9295)
         );
  NAND2_X1 U8828 ( .A1(n6896), .A2(n9297), .ZN(n9599) );
  OAI21_X1 U8829 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(P1_IR_REG_1__SCAN_IN), .A(
        n6898), .ZN(n6897) );
  CLKBUF_X1 U8830 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n14377) );
  NOR2_X1 U8831 ( .A1(n8264), .A2(n15183), .ZN(n14383) );
  INV_X1 U8832 ( .A(n7126), .ZN(n8258) );
  OAI21_X1 U8833 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n8266), .A(n15179), .ZN(
        n15168) );
  INV_X1 U8834 ( .A(n8281), .ZN(n7113) );
  XNOR2_X1 U8835 ( .A(n8285), .B(n8284), .ZN(n14394) );
  INV_X1 U8836 ( .A(n8283), .ZN(n8284) );
  NAND2_X1 U8837 ( .A1(n14394), .A2(n14393), .ZN(n14392) );
  OAI21_X1 U8838 ( .B1(n14558), .B2(n14557), .A(n6732), .ZN(n6731) );
  INV_X1 U8839 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n6732) );
  NAND2_X1 U8840 ( .A1(n14566), .A2(n14564), .ZN(n14569) );
  INV_X1 U8841 ( .A(n8295), .ZN(n7111) );
  AOI211_X1 U8842 ( .C1(n12411), .C2(n12410), .A(n12409), .B(n12408), .ZN(
        n12418) );
  OAI211_X1 U8843 ( .C1(n12658), .C2(n15116), .A(n6711), .B(n6710), .ZN(
        P3_U3201) );
  NAND2_X1 U8844 ( .A1(n12657), .A2(n15107), .ZN(n6710) );
  NOR2_X1 U8845 ( .A1(n12656), .A2(n12655), .ZN(n6711) );
  XNOR2_X1 U8846 ( .A(n12582), .B(n12581), .ZN(n12658) );
  AOI21_X1 U8847 ( .B1(P3_REG1_REG_28__SCAN_IN), .B2(n15164), .A(n6586), .ZN(
        n6706) );
  INV_X1 U8848 ( .A(n9990), .ZN(n7575) );
  OAI21_X1 U8849 ( .B1(n13227), .B2(n9998), .A(n6980), .ZN(P2_U3233) );
  AOI21_X1 U8850 ( .B1(n6982), .B2(n9998), .A(n6981), .ZN(n6980) );
  OAI21_X1 U8851 ( .B1(n14871), .B2(n6622), .A(n13228), .ZN(n6981) );
  NAND2_X1 U8852 ( .A1(n7339), .A2(n7333), .ZN(n7329) );
  OR2_X1 U8853 ( .A1(n6443), .A2(n7193), .ZN(n7192) );
  NAND2_X1 U8854 ( .A1(n6635), .A2(n6443), .ZN(n7194) );
  INV_X1 U8855 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n7193) );
  INV_X1 U8856 ( .A(n6684), .ZN(n6683) );
  NAND2_X1 U8857 ( .A1(n6716), .A2(n6719), .ZN(n6685) );
  OAI211_X1 U8858 ( .C1(n14123), .C2(n6802), .A(n6801), .B(n6799), .ZN(
        P1_U3523) );
  NAND2_X1 U8859 ( .A1(n14827), .A2(n14805), .ZN(n6802) );
  NAND2_X1 U8860 ( .A1(n14119), .A2(n6798), .ZN(n6801) );
  INV_X1 U8861 ( .A(n6800), .ZN(n6799) );
  XNOR2_X1 U8862 ( .A(n6733), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  NAND2_X1 U8863 ( .A1(n7120), .A2(n6734), .ZN(n6733) );
  XNOR2_X1 U8864 ( .A(n8302), .B(n6604), .ZN(n7118) );
  CLKBUF_X3 U8865 ( .A(n8344), .Z(n8514) );
  NAND2_X2 U8866 ( .A1(n9514), .A2(n10182), .ZN(n10161) );
  AND2_X1 U8867 ( .A1(n10135), .A2(n14090), .ZN(n10328) );
  NAND2_X2 U8868 ( .A1(n8303), .A2(n9998), .ZN(n8344) );
  NOR2_X1 U8869 ( .A1(n12443), .A2(n7098), .ZN(n6455) );
  AND2_X1 U8870 ( .A1(n6520), .A2(n7229), .ZN(n6456) );
  NOR2_X1 U8871 ( .A1(n9514), .A2(n9300), .ZN(n10135) );
  INV_X1 U8872 ( .A(n10161), .ZN(n9765) );
  INV_X1 U8873 ( .A(n10151), .ZN(n6715) );
  AND2_X1 U8874 ( .A1(n9197), .A2(n9095), .ZN(n12320) );
  INV_X2 U8875 ( .A(n10225), .ZN(n10326) );
  OR2_X1 U8876 ( .A1(n8451), .A2(n8450), .ZN(n6457) );
  NAND2_X1 U8877 ( .A1(n13950), .A2(n13958), .ZN(n6458) );
  NAND2_X1 U8878 ( .A1(n11781), .A2(n11780), .ZN(n14121) );
  NAND2_X1 U8879 ( .A1(n7801), .A2(n7800), .ZN(n11146) );
  INV_X1 U8880 ( .A(n6877), .ZN(n15027) );
  OR2_X1 U8881 ( .A1(n15008), .A2(n12565), .ZN(n6877) );
  INV_X1 U8882 ( .A(n12061), .ZN(n6906) );
  AND2_X1 U8883 ( .A1(n7222), .A2(n11542), .ZN(n6459) );
  INV_X1 U8884 ( .A(n12808), .ZN(n7434) );
  AND2_X1 U8885 ( .A1(n11492), .A2(n14377), .ZN(n6460) );
  INV_X1 U8886 ( .A(n12483), .ZN(n7099) );
  AND2_X1 U8887 ( .A1(n11401), .A2(n7283), .ZN(n6461) );
  AND2_X1 U8888 ( .A1(n12126), .A2(n13086), .ZN(n6462) );
  INV_X1 U8889 ( .A(n11597), .ZN(n7278) );
  AND3_X1 U8890 ( .A1(n7363), .A2(n7362), .A3(n7585), .ZN(n6463) );
  AND2_X1 U8891 ( .A1(n7171), .A2(n7169), .ZN(n6464) );
  NOR2_X1 U8892 ( .A1(n9605), .A2(n10717), .ZN(n6465) );
  NOR2_X1 U8893 ( .A1(n7572), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6466) );
  INV_X1 U8894 ( .A(n7240), .ZN(n7239) );
  OAI21_X1 U8895 ( .B1(n7794), .B2(n7241), .A(n7834), .ZN(n7240) );
  NOR2_X1 U8896 ( .A1(n13456), .A2(n13462), .ZN(n6467) );
  INV_X1 U8897 ( .A(n7208), .ZN(n7207) );
  NAND2_X1 U8898 ( .A1(n7209), .A2(n11208), .ZN(n7208) );
  INV_X1 U8899 ( .A(n7420), .ZN(n7419) );
  OAI21_X1 U8900 ( .B1(n12243), .B2(n7421), .A(n12549), .ZN(n7420) );
  AND2_X1 U8901 ( .A1(n13472), .A2(n13357), .ZN(n6468) );
  NOR2_X1 U8902 ( .A1(n6458), .A2(n6813), .ZN(n6812) );
  NAND2_X1 U8903 ( .A1(n8108), .A2(n8107), .ZN(n13444) );
  INV_X1 U8904 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7164) );
  NOR2_X1 U8905 ( .A1(n7375), .A2(n7374), .ZN(n6469) );
  INV_X1 U8906 ( .A(n12287), .ZN(n6869) );
  AND2_X1 U8907 ( .A1(n14370), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6470) );
  AND2_X1 U8908 ( .A1(n9519), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6471) );
  AND2_X1 U8909 ( .A1(n13444), .A2(n11560), .ZN(n6472) );
  OR2_X1 U8910 ( .A1(n12069), .A2(n12075), .ZN(n6473) );
  AND2_X1 U8911 ( .A1(n8454), .A2(n8453), .ZN(n6474) );
  AND2_X1 U8912 ( .A1(n11552), .A2(n11551), .ZN(n6475) );
  AND2_X1 U8913 ( .A1(n12567), .A2(n12605), .ZN(n6476) );
  AND2_X1 U8914 ( .A1(n6999), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n6477) );
  AND2_X1 U8915 ( .A1(n12631), .A2(n6757), .ZN(n6478) );
  NAND2_X1 U8916 ( .A1(n8183), .A2(n13377), .ZN(n14507) );
  INV_X1 U8917 ( .A(n12975), .ZN(n7130) );
  INV_X1 U8918 ( .A(n9459), .ZN(n6701) );
  INV_X2 U8919 ( .A(n9766), .ZN(n11807) );
  NAND2_X2 U8920 ( .A1(n9521), .A2(n9519), .ZN(n9605) );
  NAND2_X2 U8921 ( .A1(n7551), .A2(n7550), .ZN(n8319) );
  OR2_X1 U8922 ( .A1(n8967), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n6479) );
  INV_X1 U8923 ( .A(n7571), .ZN(n7686) );
  NAND2_X1 U8924 ( .A1(n7044), .A2(n8743), .ZN(n10051) );
  OR2_X1 U8925 ( .A1(n13300), .A2(n13077), .ZN(n6480) );
  NAND2_X2 U8926 ( .A1(n11501), .A2(n12935), .ZN(n8731) );
  INV_X1 U8927 ( .A(n9521), .ZN(n14367) );
  NAND2_X1 U8928 ( .A1(n13636), .A2(n13635), .ZN(n13634) );
  AND2_X1 U8929 ( .A1(n7144), .A2(n7143), .ZN(n6481) );
  NAND4_X1 U8930 ( .A1(n8885), .A2(n8884), .A3(n8883), .A4(n8882), .ZN(n12549)
         );
  OAI211_X1 U8931 ( .C1(n6444), .C2(n10151), .A(n10150), .B(n10149), .ZN(
        n14753) );
  INV_X1 U8932 ( .A(n11267), .ZN(n7204) );
  NAND2_X1 U8933 ( .A1(n9458), .A2(n7490), .ZN(n7590) );
  NAND2_X1 U8934 ( .A1(n7248), .A2(n7741), .ZN(n7247) );
  NAND4_X1 U8935 ( .A1(n8902), .A2(n7448), .A3(n7442), .A4(n7061), .ZN(n6482)
         );
  OR2_X1 U8936 ( .A1(n7610), .A2(n9596), .ZN(n6483) );
  XNOR2_X1 U8937 ( .A(n14121), .B(n13832), .ZN(n13896) );
  AND2_X1 U8938 ( .A1(n11551), .A2(n11553), .ZN(n6484) );
  NAND2_X1 U8939 ( .A1(n11975), .A2(n13821), .ZN(n14039) );
  OR2_X1 U8940 ( .A1(n14070), .A2(n13844), .ZN(n6485) );
  INV_X1 U8941 ( .A(n13877), .ZN(n7179) );
  NOR2_X1 U8942 ( .A1(n10051), .A2(n10101), .ZN(n6486) );
  AND2_X1 U8943 ( .A1(n6615), .A2(n7272), .ZN(n6487) );
  OR2_X1 U8944 ( .A1(n13894), .A2(n13896), .ZN(n6488) );
  AND3_X1 U8945 ( .A1(n8752), .A2(n8751), .A3(n8750), .ZN(n6489) );
  INV_X1 U8946 ( .A(n14742), .ZN(n12035) );
  NAND2_X1 U8947 ( .A1(n11892), .A2(n11891), .ZN(n14742) );
  AND2_X1 U8948 ( .A1(n11264), .A2(n9999), .ZN(n8303) );
  INV_X1 U8949 ( .A(n13850), .ZN(n6813) );
  AND2_X1 U8950 ( .A1(n7136), .A2(n7135), .ZN(n6490) );
  AND2_X1 U8951 ( .A1(n8588), .A2(n8912), .ZN(n6491) );
  OR2_X1 U8952 ( .A1(n7377), .A2(n6474), .ZN(n6492) );
  AND2_X1 U8953 ( .A1(n6804), .A2(n14122), .ZN(n6493) );
  AND2_X1 U8954 ( .A1(n8349), .A2(n8348), .ZN(n6494) );
  AND2_X1 U8955 ( .A1(n6863), .A2(n6867), .ZN(n6495) );
  OR2_X1 U8956 ( .A1(n12736), .A2(n12540), .ZN(n6496) );
  INV_X1 U8957 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8684) );
  OR2_X1 U8958 ( .A1(n13335), .A2(n13347), .ZN(n6497) );
  INV_X1 U8959 ( .A(n14703), .ZN(n10752) );
  OR2_X1 U8960 ( .A1(n13481), .A2(n13358), .ZN(n6498) );
  AOI21_X1 U8961 ( .B1(n9195), .B2(n12766), .A(n9194), .ZN(n12419) );
  AND2_X1 U8962 ( .A1(n14010), .A2(n13821), .ZN(n6499) );
  OR3_X1 U8963 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        P3_IR_REG_1__SCAN_IN), .ZN(n6500) );
  XNOR2_X1 U8964 ( .A(n13868), .B(n13812), .ZN(n6501) );
  NAND2_X1 U8965 ( .A1(n8737), .A2(n8584), .ZN(n8772) );
  OR2_X1 U8966 ( .A1(n13340), .A2(n13465), .ZN(n6502) );
  INV_X1 U8967 ( .A(n11938), .ZN(n6937) );
  AND2_X1 U8968 ( .A1(n12808), .A2(n7437), .ZN(n6503) );
  INV_X1 U8969 ( .A(n12546), .ZN(n12811) );
  OR2_X1 U8970 ( .A1(n13477), .A2(n13373), .ZN(n6504) );
  NAND2_X1 U8971 ( .A1(n12482), .A2(n12770), .ZN(n6505) );
  AND2_X1 U8972 ( .A1(n6970), .A2(n6969), .ZN(n6506) );
  XNOR2_X1 U8973 ( .A(n14133), .B(n13924), .ZN(n13938) );
  INV_X1 U8974 ( .A(n13938), .ZN(n6814) );
  AND2_X1 U8975 ( .A1(n13498), .A2(n13080), .ZN(n6507) );
  AND2_X1 U8976 ( .A1(n12049), .A2(n7183), .ZN(n6508) );
  OR2_X1 U8977 ( .A1(n8380), .A2(n8379), .ZN(n6509) );
  AND2_X1 U8978 ( .A1(n9045), .A2(n12312), .ZN(n6510) );
  OR2_X1 U8979 ( .A1(n8391), .A2(n8390), .ZN(n6511) );
  OR2_X1 U8980 ( .A1(n8355), .A2(n8354), .ZN(n6512) );
  AND2_X1 U8981 ( .A1(n12165), .A2(n12677), .ZN(n6513) );
  AND2_X1 U8982 ( .A1(n12152), .A2(n12758), .ZN(n6514) );
  AND2_X1 U8983 ( .A1(n8383), .A2(n8382), .ZN(n6515) );
  AND2_X1 U8984 ( .A1(n11936), .A2(n11405), .ZN(n6516) );
  OR2_X1 U8985 ( .A1(n13702), .A2(n6617), .ZN(n6517) );
  NOR2_X1 U8986 ( .A1(n7460), .A2(n7357), .ZN(n6518) );
  OR2_X1 U8987 ( .A1(n14438), .A2(n12577), .ZN(n6519) );
  OR2_X1 U8988 ( .A1(n12126), .A2(n13086), .ZN(n6520) );
  NOR2_X1 U8989 ( .A1(n9521), .A2(n9520), .ZN(n6521) );
  NOR2_X1 U8990 ( .A1(n12142), .A2(n12497), .ZN(n6522) );
  AND2_X1 U8991 ( .A1(n11948), .A2(n11949), .ZN(n6523) );
  OR2_X1 U8992 ( .A1(n8445), .A2(n7365), .ZN(n6524) );
  AND2_X1 U8993 ( .A1(n14113), .A2(n6725), .ZN(n6525) );
  AND2_X1 U8994 ( .A1(n13963), .A2(n13830), .ZN(n6526) );
  AND2_X1 U8995 ( .A1(n11146), .A2(n14499), .ZN(n6527) );
  NAND2_X1 U8996 ( .A1(n11287), .A2(n11286), .ZN(n13686) );
  INV_X1 U8997 ( .A(n10482), .ZN(n7227) );
  NAND2_X1 U8998 ( .A1(n12100), .A2(n13085), .ZN(n6528) );
  INV_X1 U8999 ( .A(n11914), .ZN(n6950) );
  NAND2_X1 U9000 ( .A1(n6778), .A2(SI_5_), .ZN(n7629) );
  INV_X1 U9001 ( .A(n7629), .ZN(n6901) );
  INV_X1 U9002 ( .A(n7323), .ZN(n7322) );
  NAND2_X1 U9003 ( .A1(n7328), .A2(n6480), .ZN(n7323) );
  AND2_X1 U9004 ( .A1(n6787), .A2(n10754), .ZN(n6529) );
  INV_X1 U9005 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7123) );
  NOR2_X1 U9006 ( .A1(n14403), .A2(n12575), .ZN(n6530) );
  OR2_X1 U9007 ( .A1(n11998), .A2(n11996), .ZN(n6531) );
  AND2_X1 U9008 ( .A1(n11535), .A2(n7327), .ZN(n6532) );
  OR2_X1 U9009 ( .A1(n9490), .A2(n10170), .ZN(n6533) );
  INV_X1 U9010 ( .A(n7325), .ZN(n7324) );
  NOR2_X1 U9011 ( .A1(n6532), .A2(n7326), .ZN(n7325) );
  AND2_X1 U9012 ( .A1(n13848), .A2(n14054), .ZN(n6534) );
  AND2_X1 U9013 ( .A1(n8085), .A2(n8084), .ZN(n13282) );
  NAND2_X1 U9014 ( .A1(n14549), .A2(n11405), .ZN(n6535) );
  AND2_X1 U9015 ( .A1(n11792), .A2(n11791), .ZN(n6536) );
  AND2_X1 U9016 ( .A1(n11624), .A2(n11623), .ZN(n6537) );
  AND2_X1 U9017 ( .A1(n7570), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6538) );
  INV_X1 U9018 ( .A(n7283), .ZN(n7282) );
  NOR2_X1 U9019 ( .A1(n13843), .A2(n14064), .ZN(n6539) );
  NOR2_X1 U9020 ( .A1(n11273), .A2(n13082), .ZN(n6540) );
  NOR2_X1 U9021 ( .A1(n11936), .A2(n11405), .ZN(n6541) );
  NOR2_X1 U9022 ( .A1(n11146), .A2(n14499), .ZN(n6542) );
  NAND2_X1 U9023 ( .A1(n6987), .A2(n14939), .ZN(n6986) );
  OR2_X1 U9024 ( .A1(n12925), .A2(n12546), .ZN(n12264) );
  INV_X1 U9025 ( .A(n12264), .ZN(n7055) );
  INV_X1 U9026 ( .A(n7088), .ZN(n7087) );
  NAND2_X1 U9027 ( .A1(n10488), .A2(n12556), .ZN(n7088) );
  INV_X1 U9028 ( .A(n6956), .ZN(n6955) );
  NAND2_X1 U9029 ( .A1(n14785), .A2(n6957), .ZN(n6956) );
  INV_X1 U9030 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n12929) );
  AND2_X1 U9031 ( .A1(n12878), .A2(n12660), .ZN(n12399) );
  OR2_X1 U9032 ( .A1(n13998), .A2(n13999), .ZN(n13997) );
  INV_X1 U9033 ( .A(n13997), .ZN(n6808) );
  OR2_X1 U9034 ( .A1(n10182), .A2(n9277), .ZN(n6543) );
  INV_X1 U9035 ( .A(n12370), .ZN(n11222) );
  NAND2_X1 U9036 ( .A1(n12463), .A2(n12545), .ZN(n6544) );
  NOR2_X1 U9037 ( .A1(n12750), .A2(n12541), .ZN(n6545) );
  NOR2_X1 U9038 ( .A1(n9177), .A2(n11510), .ZN(n6546) );
  INV_X1 U9039 ( .A(n7070), .ZN(n7069) );
  NAND2_X1 U9040 ( .A1(n12137), .A2(n7071), .ZN(n7070) );
  OAI211_X1 U9041 ( .C1(n8080), .C2(n6661), .A(n6651), .B(n6656), .ZN(n8184)
         );
  OR2_X1 U9042 ( .A1(n7444), .A2(n7443), .ZN(n6547) );
  INV_X1 U9043 ( .A(n7441), .ZN(n7438) );
  NAND2_X1 U9044 ( .A1(n11444), .A2(n12547), .ZN(n7441) );
  OR2_X1 U9045 ( .A1(n7366), .A2(n8343), .ZN(n6548) );
  INV_X1 U9046 ( .A(n7423), .ZN(n7422) );
  INV_X1 U9047 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9367) );
  AND2_X1 U9048 ( .A1(n6664), .A2(n7153), .ZN(n6549) );
  AND2_X1 U9049 ( .A1(n7855), .A2(n9568), .ZN(n6550) );
  NAND2_X1 U9050 ( .A1(n8204), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n6551) );
  AND2_X1 U9051 ( .A1(n10137), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6552) );
  AND2_X1 U9052 ( .A1(n9378), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n6553) );
  AND2_X1 U9053 ( .A1(n9381), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n6554) );
  INV_X1 U9054 ( .A(n7234), .ZN(n7233) );
  NAND2_X1 U9055 ( .A1(n11549), .A2(n11547), .ZN(n7234) );
  INV_X1 U9056 ( .A(n6968), .ZN(n13863) );
  AND2_X1 U9057 ( .A1(n13675), .A2(n13674), .ZN(n6555) );
  INV_X1 U9058 ( .A(n7412), .ZN(n7411) );
  AND2_X1 U9059 ( .A1(n12748), .A2(n6505), .ZN(n7412) );
  AND2_X1 U9060 ( .A1(n6866), .A2(n6865), .ZN(n6556) );
  INV_X1 U9061 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7518) );
  INV_X1 U9062 ( .A(n7461), .ZN(n7398) );
  INV_X1 U9063 ( .A(n7149), .ZN(n7148) );
  NAND2_X1 U9064 ( .A1(n7150), .A2(n8079), .ZN(n7149) );
  INV_X1 U9065 ( .A(n11994), .ZN(n6931) );
  NAND2_X1 U9066 ( .A1(n7485), .A2(n7469), .ZN(n7491) );
  OR2_X1 U9067 ( .A1(n11417), .A2(n7104), .ZN(n6557) );
  NAND2_X1 U9068 ( .A1(n8064), .A2(n8063), .ZN(n13456) );
  OR2_X1 U9069 ( .A1(n11680), .A2(n10140), .ZN(n6558) );
  OR2_X1 U9070 ( .A1(n8209), .A2(n7117), .ZN(n6559) );
  OR2_X1 U9071 ( .A1(n12073), .A2(n12072), .ZN(n6560) );
  AND2_X1 U9072 ( .A1(n6943), .A2(n11940), .ZN(n6561) );
  AND2_X1 U9073 ( .A1(n6943), .A2(n11944), .ZN(n6562) );
  AND2_X1 U9074 ( .A1(n7225), .A2(n6528), .ZN(n6563) );
  AND2_X1 U9075 ( .A1(n8460), .A2(n6492), .ZN(n6564) );
  NAND2_X1 U9076 ( .A1(n7042), .A2(n8747), .ZN(n15129) );
  AND2_X1 U9077 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(
        n6565) );
  INV_X1 U9078 ( .A(n7297), .ZN(n7296) );
  OAI21_X1 U9079 ( .B1(n13818), .B2(n7298), .A(n13817), .ZN(n7297) );
  OR2_X1 U9080 ( .A1(n12029), .A2(n12027), .ZN(n6566) );
  OR2_X1 U9081 ( .A1(n7364), .A2(n8446), .ZN(n6567) );
  AND2_X1 U9082 ( .A1(n12696), .A2(n6850), .ZN(n6568) );
  AND2_X1 U9083 ( .A1(n6495), .A2(n12397), .ZN(n6569) );
  OR2_X1 U9084 ( .A1(n6950), .A2(n11913), .ZN(n6570) );
  AND2_X1 U9085 ( .A1(n6805), .A2(n6804), .ZN(n6571) );
  OR2_X1 U9086 ( .A1(n6937), .A2(n11937), .ZN(n6572) );
  OR2_X1 U9087 ( .A1(n11987), .A2(n11985), .ZN(n6573) );
  OR2_X1 U9088 ( .A1(n12009), .A2(n12007), .ZN(n6574) );
  AND2_X1 U9089 ( .A1(n6930), .A2(n6531), .ZN(n6575) );
  NAND2_X1 U9090 ( .A1(n10252), .A2(n9465), .ZN(n9459) );
  INV_X1 U9091 ( .A(n7758), .ZN(n6679) );
  OR2_X1 U9092 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n6576) );
  INV_X1 U9093 ( .A(n7059), .ZN(n7058) );
  NAND2_X1 U9094 ( .A1(n12373), .A2(n7060), .ZN(n7059) );
  INV_X1 U9095 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9413) );
  INV_X1 U9096 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9759) );
  INV_X1 U9097 ( .A(n12783), .ZN(n12789) );
  AND2_X1 U9098 ( .A1(n12279), .A2(n12283), .ZN(n12783) );
  INV_X1 U9099 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n6874) );
  NAND2_X1 U9100 ( .A1(n11583), .A2(n11582), .ZN(n13562) );
  XNOR2_X1 U9101 ( .A(n14012), .B(n13996), .ZN(n14010) );
  INV_X1 U9102 ( .A(n14010), .ZN(n7169) );
  INV_X1 U9103 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7117) );
  INV_X1 U9104 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6703) );
  NAND2_X1 U9105 ( .A1(n11027), .A2(n11026), .ZN(n11946) );
  INV_X1 U9106 ( .A(n11946), .ZN(n14544) );
  OR2_X1 U9107 ( .A1(n10530), .A2(n14994), .ZN(n6577) );
  INV_X1 U9108 ( .A(n13465), .ZN(n7140) );
  OAI21_X1 U9109 ( .B1(n6721), .B2(n7073), .A(n7069), .ZN(n12457) );
  NAND2_X1 U9110 ( .A1(n12786), .A2(n12279), .ZN(n12773) );
  INV_X1 U9111 ( .A(n14144), .ZN(n6959) );
  INV_X1 U9112 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7108) );
  INV_X1 U9113 ( .A(n15026), .ZN(n6876) );
  NAND2_X1 U9114 ( .A1(n11718), .A2(n11717), .ZN(n14139) );
  INV_X1 U9115 ( .A(n8460), .ZN(n7374) );
  AND2_X1 U9116 ( .A1(n14133), .A2(n13960), .ZN(n6578) );
  AND2_X1 U9117 ( .A1(n14070), .A2(n13844), .ZN(n6579) );
  AND2_X1 U9118 ( .A1(n14504), .A2(n7156), .ZN(n6580) );
  INV_X1 U9119 ( .A(n7132), .ZN(n13408) );
  NOR2_X1 U9120 ( .A1(n13410), .A2(n13493), .ZN(n7132) );
  INV_X1 U9121 ( .A(n8641), .ZN(n7036) );
  AND2_X1 U9122 ( .A1(n7276), .A2(n7274), .ZN(n6581) );
  AND2_X1 U9123 ( .A1(n14126), .A2(n13933), .ZN(n6582) );
  AND2_X1 U9124 ( .A1(n6876), .A2(n15049), .ZN(n6583) );
  AND2_X1 U9125 ( .A1(n9808), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6584) );
  AND2_X1 U9126 ( .A1(n12485), .A2(n6455), .ZN(n6585) );
  NOR2_X1 U9127 ( .A1(n9177), .A2(n12876), .ZN(n6586) );
  AND2_X1 U9128 ( .A1(n11600), .A2(n11599), .ZN(n6587) );
  OR2_X1 U9129 ( .A1(n12616), .A2(n15033), .ZN(n6588) );
  AND2_X1 U9130 ( .A1(n6703), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n6589) );
  INV_X1 U9131 ( .A(n11541), .ZN(n7338) );
  NAND2_X1 U9132 ( .A1(n11540), .A2(n11539), .ZN(n11541) );
  OR2_X1 U9133 ( .A1(n7964), .A2(n10012), .ZN(n6590) );
  NOR2_X1 U9134 ( .A1(n8937), .A2(n7034), .ZN(n7033) );
  INV_X1 U9135 ( .A(n7968), .ZN(n6762) );
  AND2_X1 U9136 ( .A1(n6748), .A2(n6588), .ZN(n6591) );
  OR2_X1 U9137 ( .A1(n8406), .A2(n8407), .ZN(n6592) );
  OR2_X1 U9138 ( .A1(n7382), .A2(n8419), .ZN(n6593) );
  OR2_X1 U9139 ( .A1(n7372), .A2(n7371), .ZN(n6594) );
  INV_X1 U9140 ( .A(n9260), .ZN(n11843) );
  NAND2_X1 U9141 ( .A1(n9259), .A2(n9258), .ZN(n9260) );
  INV_X1 U9142 ( .A(n15049), .ZN(n12605) );
  NAND2_X1 U9143 ( .A1(n6649), .A2(n10028), .ZN(n10031) );
  INV_X2 U9144 ( .A(n15164), .ZN(n15166) );
  NAND2_X1 U9145 ( .A1(n11099), .A2(n11264), .ZN(n9571) );
  INV_X1 U9146 ( .A(n9571), .ZN(n7166) );
  OAI211_X1 U9147 ( .C1(n6639), .C2(n6637), .A(n10650), .B(n6636), .ZN(n14726)
         );
  NAND2_X1 U9148 ( .A1(n7882), .A2(n7881), .ZN(n13498) );
  INV_X1 U9149 ( .A(n13498), .ZN(n7133) );
  AND2_X1 U9150 ( .A1(n10745), .A2(n10744), .ZN(n14719) );
  AND2_X1 U9151 ( .A1(n6780), .A2(n6779), .ZN(n14740) );
  INV_X1 U9152 ( .A(n8653), .ZN(n7024) );
  INV_X1 U9153 ( .A(n7138), .ZN(n10676) );
  NOR2_X1 U9154 ( .A1(n10478), .A2(n12126), .ZN(n7138) );
  NAND2_X1 U9155 ( .A1(n10017), .A2(n10018), .ZN(n10295) );
  INV_X1 U9156 ( .A(n10295), .ZN(n7131) );
  AND2_X1 U9157 ( .A1(n6786), .A2(n6784), .ZN(n6595) );
  AND2_X1 U9158 ( .A1(n7269), .A2(n10219), .ZN(n6596) );
  AND2_X1 U9159 ( .A1(n11266), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6597) );
  NOR2_X1 U9160 ( .A1(n8656), .A2(n7022), .ZN(n7021) );
  AND2_X1 U9161 ( .A1(n7084), .A2(n7082), .ZN(n6598) );
  INV_X1 U9162 ( .A(n14454), .ZN(n6743) );
  INV_X1 U9163 ( .A(n14933), .ZN(n14931) );
  INV_X1 U9164 ( .A(n14793), .ZN(n6957) );
  INV_X1 U9165 ( .A(n10692), .ZN(n6953) );
  AND2_X1 U9166 ( .A1(n14933), .A2(n14533), .ZN(n6599) );
  NAND2_X1 U9167 ( .A1(n7774), .A2(n7773), .ZN(n12100) );
  INV_X1 U9168 ( .A(n12100), .ZN(n7137) );
  OR2_X1 U9169 ( .A1(n12593), .A2(n14481), .ZN(n6600) );
  NAND2_X1 U9170 ( .A1(n12615), .A2(n12614), .ZN(n6601) );
  INV_X1 U9171 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7110) );
  INV_X1 U9172 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7521) );
  AND2_X1 U9173 ( .A1(n7488), .A2(n7487), .ZN(n9998) );
  XOR2_X1 U9174 ( .A(n9267), .B(P2_DATAO_REG_0__SCAN_IN), .Z(n6602) );
  OR2_X1 U9175 ( .A1(n11867), .A2(n13796), .ZN(n14797) );
  AND2_X1 U9176 ( .A1(n8548), .A2(n9998), .ZN(n6603) );
  XOR2_X1 U9177 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n6604) );
  INV_X1 U9178 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6979) );
  INV_X1 U9179 ( .A(n9278), .ZN(n6617) );
  NAND2_X1 U9180 ( .A1(n9272), .A2(n9243), .ZN(n9230) );
  NOR2_X2 U9181 ( .A1(n10209), .A2(n9217), .ZN(n7290) );
  NAND4_X1 U9182 ( .A1(n9213), .A2(n9212), .A3(n9211), .A4(n9210), .ZN(n10209)
         );
  NAND4_X1 U9183 ( .A1(n6620), .A2(n6619), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7259) );
  NAND4_X1 U9184 ( .A1(n13799), .A2(n6622), .A3(P3_ADDR_REG_19__SCAN_IN), .A4(
        n6621), .ZN(n7260) );
  NAND2_X1 U9185 ( .A1(n6915), .A2(n6917), .ZN(n6626) );
  NAND2_X1 U9186 ( .A1(n7926), .A2(n6764), .ZN(n6763) );
  INV_X1 U9187 ( .A(n7904), .ZN(n6627) );
  OAI21_X1 U9188 ( .B1(n9354), .B2(n9413), .A(n6631), .ZN(n6630) );
  NAND2_X1 U9189 ( .A1(n9354), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n6631) );
  INV_X1 U9190 ( .A(n13375), .ZN(n6633) );
  NAND2_X1 U9191 ( .A1(n13390), .A2(n11545), .ZN(n6634) );
  AND2_X1 U9192 ( .A1(n10649), .A2(n6643), .ZN(n10686) );
  NAND2_X1 U9193 ( .A1(n11303), .A2(n6645), .ZN(n6644) );
  NAND2_X2 U9194 ( .A1(n11351), .A2(n11954), .ZN(n11353) );
  OR2_X2 U9195 ( .A1(n11306), .A2(n12049), .ZN(n11351) );
  NAND2_X1 U9196 ( .A1(n9246), .A2(n9247), .ZN(n6647) );
  NAND2_X2 U9197 ( .A1(n13921), .A2(n13922), .ZN(n13920) );
  NAND2_X2 U9198 ( .A1(n10848), .A2(n10847), .ZN(n10849) );
  OR2_X2 U9199 ( .A1(n10774), .A2(n12042), .ZN(n10848) );
  OAI21_X2 U9200 ( .B1(n14681), .B2(n10771), .A(n10772), .ZN(n10774) );
  AND2_X2 U9201 ( .A1(n14370), .A2(n9521), .ZN(n11814) );
  NAND2_X1 U9202 ( .A1(n10089), .A2(n7649), .ZN(n6649) );
  AND2_X2 U9203 ( .A1(n7517), .A2(n11102), .ZN(n9999) );
  NAND3_X1 U9204 ( .A1(n7468), .A2(n7679), .A3(n7164), .ZN(n7482) );
  INV_X1 U9205 ( .A(n13030), .ZN(n6668) );
  OAI211_X1 U9206 ( .C1(n6680), .C2(n6679), .A(n12095), .B(n6678), .ZN(n12102)
         );
  NAND3_X1 U9207 ( .A1(n7758), .A2(n7160), .A3(n10208), .ZN(n6678) );
  NAND2_X1 U9208 ( .A1(n12119), .A2(n6680), .ZN(n12128) );
  XNOR2_X1 U9209 ( .A(n8000), .B(n7998), .ZN(n13042) );
  NAND2_X1 U9210 ( .A1(n7982), .A2(n7981), .ZN(n8000) );
  OR2_X1 U9211 ( .A1(n7669), .A2(n7670), .ZN(n7671) );
  NAND2_X1 U9212 ( .A1(n9303), .A2(n9304), .ZN(n9489) );
  NAND2_X1 U9213 ( .A1(n7651), .A2(n6681), .ZN(n10320) );
  INV_X1 U9214 ( .A(n6897), .ZN(n6896) );
  NAND2_X1 U9215 ( .A1(n6685), .A2(n6683), .ZN(P1_U3262) );
  OAI21_X1 U9216 ( .B1(n14679), .B2(n13799), .A(n13798), .ZN(n6684) );
  NAND2_X1 U9217 ( .A1(n9322), .A2(n9323), .ZN(n9321) );
  OR2_X1 U9218 ( .A1(n9599), .A2(n10718), .ZN(n6686) );
  AOI21_X1 U9219 ( .B1(n10726), .B2(P1_REG2_REG_9__SCAN_IN), .A(n10352), .ZN(
        n14591) );
  AOI21_X1 U9220 ( .B1(n13783), .B2(P1_REG2_REG_14__SCAN_IN), .A(n14619), .ZN(
        n13774) );
  AOI21_X1 U9221 ( .B1(n13762), .B2(P1_REG2_REG_11__SCAN_IN), .A(n13761), .ZN(
        n13765) );
  AOI21_X1 U9222 ( .B1(n14649), .B2(P1_REG2_REG_16__SCAN_IN), .A(n14644), .ZN(
        n14655) );
  OAI21_X1 U9223 ( .B1(n13795), .B2(n14669), .A(n14618), .ZN(n6885) );
  INV_X1 U9224 ( .A(n6885), .ZN(n6718) );
  AOI21_X1 U9225 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n14661), .A(n14653), .ZN(
        n13776) );
  AOI21_X1 U9226 ( .B1(n14610), .B2(P1_REG2_REG_13__SCAN_IN), .A(n14602), .ZN(
        n14621) );
  NAND2_X1 U9227 ( .A1(n6457), .A2(n6564), .ZN(n6829) );
  OAI21_X1 U9228 ( .B1(n8364), .B2(n7456), .A(n8363), .ZN(n8370) );
  OAI21_X1 U9229 ( .B1(n6822), .B2(n6820), .A(n6819), .ZN(n8355) );
  OAI21_X1 U9230 ( .B1(n8386), .B2(n6818), .A(n6817), .ZN(n8391) );
  AOI21_X1 U9231 ( .B1(n8441), .B2(n8440), .A(n8439), .ZN(n6815) );
  OAI21_X1 U9232 ( .B1(n8425), .B2(n6837), .A(n6834), .ZN(n8431) );
  OAI21_X1 U9233 ( .B1(n8339), .B2(n8338), .A(n6687), .ZN(n7369) );
  NAND2_X1 U9234 ( .A1(n6689), .A2(n6688), .ZN(n6687) );
  NAND2_X1 U9235 ( .A1(n8339), .A2(n8338), .ZN(n6689) );
  OAI21_X2 U9236 ( .B1(n7879), .B2(n7497), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n7498) );
  AOI21_X1 U9237 ( .B1(n8368), .B2(n7396), .A(n7392), .ZN(n8380) );
  OAI21_X1 U9238 ( .B1(n8452), .B2(n6829), .A(n6827), .ZN(n6826) );
  NOR2_X1 U9239 ( .A1(n6494), .A2(n6821), .ZN(n6820) );
  INV_X1 U9240 ( .A(n8381), .ZN(n6690) );
  NAND2_X1 U9241 ( .A1(n6690), .A2(n6509), .ZN(n8386) );
  INV_X1 U9242 ( .A(n8392), .ZN(n6691) );
  NAND2_X1 U9243 ( .A1(n6691), .A2(n6511), .ZN(n8398) );
  INV_X1 U9244 ( .A(n8356), .ZN(n6692) );
  NAND2_X1 U9245 ( .A1(n6692), .A2(n6512), .ZN(n8362) );
  OAI21_X1 U9246 ( .B1(n6816), .B2(n6815), .A(n6567), .ZN(n8451) );
  NAND2_X1 U9247 ( .A1(n9736), .A2(n9735), .ZN(n9944) );
  NAND2_X2 U9248 ( .A1(n7199), .A2(n6693), .ZN(n13097) );
  NAND2_X1 U9249 ( .A1(n9951), .A2(n7560), .ZN(n9822) );
  INV_X1 U9250 ( .A(n9822), .ZN(n6709) );
  OAI21_X1 U9251 ( .B1(n11353), .B2(n7297), .A(n7293), .ZN(n13820) );
  XNOR2_X1 U9252 ( .A(n9943), .B(n7534), .ZN(n9735) );
  NAND2_X1 U9253 ( .A1(n9944), .A2(n7536), .ZN(n7556) );
  OR2_X1 U9254 ( .A1(n7677), .A2(n7676), .ZN(n7678) );
  OAI21_X1 U9255 ( .B1(n6450), .B2(n9759), .A(n6699), .ZN(n7538) );
  NAND2_X1 U9256 ( .A1(n12102), .A2(n7785), .ZN(n13030) );
  NAND2_X1 U9257 ( .A1(n12968), .A2(n7698), .ZN(n7716) );
  NAND4_X2 U9258 ( .A1(n7595), .A2(n7594), .A3(n7593), .A4(n7592), .ZN(n13093)
         );
  NAND2_X2 U9259 ( .A1(n6700), .A2(n6483), .ZN(n8312) );
  INV_X1 U9260 ( .A(n7516), .ZN(n6700) );
  NAND2_X1 U9261 ( .A1(n11211), .A2(n6459), .ZN(n7220) );
  NAND2_X1 U9262 ( .A1(n10285), .A2(n10284), .ZN(n10390) );
  NAND2_X1 U9263 ( .A1(n14514), .A2(n14513), .ZN(n14512) );
  NAND2_X1 U9264 ( .A1(n14512), .A2(n7872), .ZN(n7893) );
  NAND2_X1 U9265 ( .A1(n10146), .A2(n10145), .ZN(n13578) );
  NAND2_X1 U9266 ( .A1(n9770), .A2(n9771), .ZN(n10146) );
  AND2_X1 U9267 ( .A1(n7526), .A2(n7527), .ZN(n7199) );
  NAND2_X1 U9268 ( .A1(n6723), .A2(n9702), .ZN(n9769) );
  NAND2_X1 U9269 ( .A1(n13248), .A2(n11562), .ZN(n7197) );
  INV_X1 U9270 ( .A(n10286), .ZN(n10285) );
  NAND2_X1 U9271 ( .A1(n9459), .A2(n7198), .ZN(n9575) );
  NAND2_X1 U9272 ( .A1(n13831), .A2(n13859), .ZN(n13898) );
  NAND2_X1 U9273 ( .A1(n14726), .A2(n7302), .ZN(n7301) );
  OAI211_X1 U9274 ( .C1(n14123), .C2(n14797), .A(n6805), .B(n6493), .ZN(n14203) );
  NAND2_X2 U9275 ( .A1(n10672), .A2(n10671), .ZN(n10674) );
  NAND2_X1 U9276 ( .A1(n6728), .A2(n6727), .ZN(n11199) );
  NAND2_X1 U9277 ( .A1(n6729), .A2(n9925), .ZN(n10020) );
  NAND2_X1 U9278 ( .A1(n13882), .A2(n13860), .ZN(n13862) );
  NAND2_X1 U9279 ( .A1(n6812), .A2(n6811), .ZN(n6810) );
  NAND2_X1 U9280 ( .A1(n7704), .A2(n7703), .ZN(n7722) );
  OAI21_X1 U9281 ( .B1(n7510), .B2(SI_1_), .A(n7236), .ZN(n7514) );
  AND2_X2 U9282 ( .A1(n6705), .A2(n9132), .ZN(n12672) );
  NAND3_X1 U9283 ( .A1(n9123), .A2(n9178), .A3(n12766), .ZN(n6705) );
  OR2_X2 U9284 ( .A1(n9118), .A2(n12320), .ZN(n11504) );
  NAND2_X1 U9285 ( .A1(n6707), .A2(n6706), .ZN(P3_U3487) );
  NAND2_X1 U9286 ( .A1(n9174), .A2(n15166), .ZN(n6707) );
  NAND4_X2 U9287 ( .A1(n7062), .A2(n8902), .A3(n8684), .A4(n7448), .ZN(n8712)
         );
  NOR2_X4 U9288 ( .A1(n8676), .A2(n6842), .ZN(n7448) );
  INV_X1 U9289 ( .A(n10091), .ZN(n7648) );
  NAND2_X1 U9290 ( .A1(n7647), .A2(n7649), .ZN(n10091) );
  INV_X1 U9291 ( .A(n9823), .ZN(n6722) );
  NAND2_X2 U9292 ( .A1(n7569), .A2(n7568), .ZN(n10006) );
  NOR2_X1 U9293 ( .A1(n14670), .A2(n13777), .ZN(n13778) );
  NAND2_X1 U9294 ( .A1(n14562), .A2(n14561), .ZN(n14560) );
  XNOR2_X1 U9295 ( .A(n8280), .B(n7113), .ZN(n14391) );
  XNOR2_X1 U9296 ( .A(n8296), .B(n7111), .ZN(n14402) );
  NAND2_X1 U9297 ( .A1(n15175), .A2(n15176), .ZN(n15174) );
  NAND2_X1 U9298 ( .A1(n14378), .A2(n14379), .ZN(n7122) );
  INV_X1 U9299 ( .A(n8292), .ZN(n8294) );
  NAND2_X1 U9300 ( .A1(n7120), .A2(n7121), .ZN(n7119) );
  XNOR2_X1 U9301 ( .A(n7119), .B(n7118), .ZN(SUB_1596_U4) );
  INV_X1 U9302 ( .A(n7291), .ZN(n9388) );
  NAND2_X1 U9303 ( .A1(n15172), .A2(n15171), .ZN(n15170) );
  NAND2_X1 U9304 ( .A1(n15174), .A2(n7114), .ZN(n8280) );
  NAND2_X1 U9305 ( .A1(n6730), .A2(n14577), .ZN(n8296) );
  NAND2_X1 U9306 ( .A1(n14556), .A2(n6731), .ZN(n14562) );
  NAND2_X1 U9307 ( .A1(n10489), .A2(n10490), .ZN(n10706) );
  NAND2_X4 U9308 ( .A1(n14367), .A2(n14370), .ZN(n11816) );
  XNOR2_X1 U9309 ( .A(n13878), .B(n7179), .ZN(n7315) );
  INV_X1 U9310 ( .A(n7231), .ZN(n7230) );
  INV_X1 U9311 ( .A(n7762), .ZN(n7248) );
  OR2_X1 U9312 ( .A1(n10748), .A2(n7908), .ZN(n7685) );
  NAND2_X2 U9313 ( .A1(n7655), .A2(n7654), .ZN(n7673) );
  NAND2_X2 U9314 ( .A1(n7771), .A2(n9354), .ZN(n8487) );
  INV_X1 U9315 ( .A(n9701), .ZN(n6723) );
  NAND2_X1 U9316 ( .A1(n10162), .A2(n10163), .ZN(n10219) );
  NAND2_X1 U9317 ( .A1(n7286), .A2(n7285), .ZN(n11131) );
  OAI21_X2 U9318 ( .B1(n7608), .B2(n6901), .A(n6724), .ZN(n7651) );
  NAND2_X1 U9319 ( .A1(n7605), .A2(n7604), .ZN(n7608) );
  NAND2_X1 U9320 ( .A1(n13898), .A2(n13833), .ZN(n13878) );
  NAND2_X1 U9321 ( .A1(n14112), .A2(n6525), .ZN(n14201) );
  OAI21_X2 U9322 ( .B1(n10849), .B2(n7308), .A(n7306), .ZN(n11033) );
  NAND2_X1 U9323 ( .A1(n7608), .A2(n7607), .ZN(n7630) );
  OAI21_X1 U9324 ( .B1(n6449), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n6726), .ZN(
        n6918) );
  NAND3_X2 U9325 ( .A1(n7353), .A2(n6825), .A3(n7352), .ZN(n13094) );
  AOI22_X4 U9326 ( .A1(n13304), .A2(n13308), .B1(n11534), .B2(n13462), .ZN(
        n13292) );
  INV_X1 U9327 ( .A(n9931), .ZN(n6729) );
  INV_X1 U9328 ( .A(n11148), .ZN(n6728) );
  NAND2_X1 U9329 ( .A1(n7677), .A2(n7676), .ZN(n7700) );
  OAI21_X2 U9330 ( .B1(n13329), .B2(n11533), .A(n11532), .ZN(n13304) );
  NAND2_X1 U9331 ( .A1(n7651), .A2(n7650), .ZN(n7655) );
  AOI21_X2 U9332 ( .B1(n13404), .B2(n11527), .A(n11526), .ZN(n13391) );
  NAND2_X1 U9333 ( .A1(n7194), .A2(n7192), .ZN(P2_U3496) );
  OAI21_X1 U9334 ( .B1(n10395), .B2(n7342), .A(n7340), .ZN(n10474) );
  XNOR2_X1 U9335 ( .A(n11537), .B(n11563), .ZN(n7339) );
  NOR2_X1 U9336 ( .A1(n8256), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n8207) );
  NOR2_X2 U9337 ( .A1(n8294), .A2(n8293), .ZN(n14573) );
  NAND2_X1 U9338 ( .A1(n14378), .A2(n14379), .ZN(n6734) );
  XNOR2_X2 U9339 ( .A(n6740), .B(P3_IR_REG_27__SCAN_IN), .ZN(n10514) );
  NAND3_X1 U9340 ( .A1(n7448), .A2(n8902), .A3(n7062), .ZN(n6741) );
  NAND2_X1 U9341 ( .A1(n6747), .A2(n6591), .ZN(n15053) );
  INV_X1 U9342 ( .A(n15088), .ZN(n6753) );
  AOI21_X1 U9343 ( .B1(n6753), .B2(n6478), .A(n6754), .ZN(n12638) );
  NAND2_X1 U9344 ( .A1(n6758), .A2(n6760), .ZN(n8037) );
  NAND3_X1 U9345 ( .A1(n6764), .A2(n7968), .A3(n7926), .ZN(n6758) );
  NAND2_X1 U9346 ( .A1(n7926), .A2(n7925), .ZN(n7966) );
  NAND2_X1 U9347 ( .A1(n7673), .A2(n6768), .ZN(n6765) );
  NAND2_X1 U9348 ( .A1(n6766), .A2(n6765), .ZN(n6914) );
  NAND2_X1 U9349 ( .A1(n7673), .A2(n7672), .ZN(n7677) );
  OAI21_X1 U9350 ( .B1(SI_5_), .B2(n6778), .A(n7629), .ZN(n7606) );
  MUX2_X1 U9351 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n9354), .Z(n6778) );
  NAND3_X1 U9352 ( .A1(n11887), .A2(n14741), .A3(n10658), .ZN(n6779) );
  NAND3_X1 U9353 ( .A1(n6781), .A2(n10658), .A3(n10657), .ZN(n6780) );
  NAND2_X1 U9354 ( .A1(n6781), .A2(n10657), .ZN(n10685) );
  OAI21_X1 U9355 ( .B1(n6784), .B2(n6783), .A(n6782), .ZN(n10891) );
  NAND2_X1 U9356 ( .A1(n11341), .A2(n6793), .ZN(n6792) );
  OR2_X1 U9357 ( .A1(n14827), .A2(n11782), .ZN(n6803) );
  NAND2_X1 U9358 ( .A1(n6494), .A2(n6821), .ZN(n6819) );
  INV_X1 U9359 ( .A(n8350), .ZN(n6821) );
  OAI21_X1 U9360 ( .B1(n7369), .B2(n7367), .A(n6548), .ZN(n6822) );
  NOR2_X1 U9361 ( .A1(n6466), .A2(n6538), .ZN(n6825) );
  NAND3_X1 U9362 ( .A1(n6830), .A2(n7387), .A3(n6826), .ZN(n7384) );
  NAND3_X1 U9363 ( .A1(n7373), .A2(n7375), .A3(n7374), .ZN(n6830) );
  INV_X1 U9364 ( .A(n6831), .ZN(n8430) );
  NAND2_X1 U9365 ( .A1(n6841), .A2(n6838), .ZN(n13539) );
  NAND2_X1 U9366 ( .A1(n6841), .A2(n6839), .ZN(n7520) );
  NAND3_X1 U9367 ( .A1(n8679), .A2(n8677), .A3(n8678), .ZN(n6842) );
  NAND2_X1 U9368 ( .A1(n10829), .A2(n6846), .ZN(n6843) );
  NAND2_X1 U9369 ( .A1(n6843), .A2(n6844), .ZN(n8880) );
  OR2_X1 U9370 ( .A1(n9045), .A2(n6852), .ZN(n6849) );
  NAND2_X1 U9371 ( .A1(n6849), .A2(n6568), .ZN(n12695) );
  NAND2_X1 U9372 ( .A1(n11246), .A2(n6855), .ZN(n7050) );
  NAND2_X1 U9373 ( .A1(n7050), .A2(n7048), .ZN(n8924) );
  NAND2_X1 U9374 ( .A1(n12678), .A2(n6495), .ZN(n6857) );
  AOI21_X1 U9375 ( .B1(n12678), .B2(n6569), .A(n6858), .ZN(n12403) );
  NAND2_X1 U9376 ( .A1(n12678), .A2(n6863), .ZN(n11509) );
  NAND2_X1 U9377 ( .A1(n12678), .A2(n12318), .ZN(n11507) );
  INV_X1 U9378 ( .A(n12396), .ZN(n6866) );
  NAND2_X1 U9379 ( .A1(n12788), .A2(n6871), .ZN(n6870) );
  XNOR2_X2 U9380 ( .A(n8744), .B(P3_IR_REG_2__SCAN_IN), .ZN(n10521) );
  OAI21_X2 U9381 ( .B1(n14404), .B2(n6882), .A(n6881), .ZN(n14433) );
  XNOR2_X2 U9382 ( .A(n12574), .B(n14408), .ZN(n14404) );
  NAND3_X1 U9383 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .A3(
        n14377), .ZN(n6898) );
  NAND3_X1 U9384 ( .A1(n6501), .A2(n6907), .A3(n6906), .ZN(n6905) );
  MUX2_X1 U9385 ( .A(n12065), .B(n12066), .S(n12068), .Z(n6909) );
  NOR2_X1 U9386 ( .A1(n6918), .A2(n14225), .ZN(n7512) );
  XNOR2_X2 U9387 ( .A(n8004), .B(SI_22_), .ZN(n11678) );
  OAI21_X2 U9388 ( .B1(n7984), .B2(n7983), .A(n7985), .ZN(n8004) );
  XNOR2_X2 U9389 ( .A(n8025), .B(SI_21_), .ZN(n7984) );
  AND2_X2 U9390 ( .A1(n14376), .A2(n6444), .ZN(n14149) );
  XNOR2_X2 U9391 ( .A(n11679), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14376) );
  OAI22_X2 U9392 ( .A1(n12011), .A2(n6920), .B1(n12012), .B2(n6919), .ZN(
        n12016) );
  NAND2_X1 U9393 ( .A1(n12016), .A2(n12017), .ZN(n12015) );
  NAND2_X1 U9394 ( .A1(n6922), .A2(n6921), .ZN(n9278) );
  NAND3_X2 U9395 ( .A1(n9253), .A2(n6926), .A3(n6923), .ZN(n13702) );
  NAND2_X1 U9396 ( .A1(n13702), .A2(n9278), .ZN(n10655) );
  NAND2_X1 U9397 ( .A1(n6928), .A2(n6575), .ZN(n7257) );
  NAND3_X1 U9398 ( .A1(n11993), .A2(n6929), .A3(n11992), .ZN(n6928) );
  OR2_X1 U9399 ( .A1(n6931), .A2(n11995), .ZN(n6930) );
  OAI22_X2 U9400 ( .A1(n11926), .A2(n6933), .B1(n11925), .B2(n6932), .ZN(
        n11930) );
  NAND2_X1 U9401 ( .A1(n6935), .A2(n6936), .ZN(n11942) );
  NAND3_X1 U9402 ( .A1(n11935), .A2(n6572), .A3(n11934), .ZN(n6935) );
  NAND2_X1 U9403 ( .A1(n6938), .A2(n6939), .ZN(n11991) );
  NAND3_X1 U9404 ( .A1(n11984), .A2(n6573), .A3(n11983), .ZN(n6938) );
  NAND2_X1 U9405 ( .A1(n11941), .A2(n6561), .ZN(n6942) );
  NAND2_X1 U9406 ( .A1(n11945), .A2(n6562), .ZN(n6940) );
  NAND3_X1 U9407 ( .A1(n6942), .A2(n6941), .A3(n6940), .ZN(n11958) );
  NAND2_X1 U9408 ( .A1(n11902), .A2(n11901), .ZN(n11900) );
  NOR2_X1 U9409 ( .A1(n6947), .A2(n11896), .ZN(n6946) );
  NAND2_X1 U9410 ( .A1(n6948), .A2(n6949), .ZN(n11917) );
  NAND3_X1 U9411 ( .A1(n11912), .A2(n6570), .A3(n11911), .ZN(n6948) );
  NAND2_X2 U9412 ( .A1(n14757), .A2(n14773), .ZN(n14755) );
  AND2_X2 U9413 ( .A1(n6953), .A2(n6952), .ZN(n14757) );
  INV_X1 U9414 ( .A(n10695), .ZN(n6952) );
  INV_X1 U9415 ( .A(n6958), .ZN(n14714) );
  NOR2_X2 U9416 ( .A1(n13953), .A2(n14133), .ZN(n13939) );
  NAND2_X2 U9417 ( .A1(n11029), .A2(n6961), .ZN(n11346) );
  XNOR2_X1 U9418 ( .A(n7506), .B(n7507), .ZN(n9526) );
  INV_X1 U9419 ( .A(n15095), .ZN(n6984) );
  NOR2_X2 U9420 ( .A1(n14447), .A2(n14448), .ZN(n14449) );
  AOI21_X1 U9421 ( .B1(n15027), .B2(n6476), .A(n6995), .ZN(n6994) );
  NAND2_X1 U9422 ( .A1(n15024), .A2(n6476), .ZN(n6998) );
  NAND2_X1 U9423 ( .A1(n15026), .A2(n6476), .ZN(n6996) );
  NAND3_X1 U9424 ( .A1(n6998), .A2(n6999), .A3(n6997), .ZN(n15044) );
  NAND2_X1 U9425 ( .A1(n9083), .A2(n8672), .ZN(n8674) );
  NAND2_X1 U9426 ( .A1(n9069), .A2(n8669), .ZN(n7001) );
  NAND2_X1 U9427 ( .A1(n8631), .A2(n7010), .ZN(n7009) );
  XNOR2_X2 U9428 ( .A(n8664), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n9046) );
  OAI21_X1 U9429 ( .B1(n8758), .B2(n8615), .A(n8616), .ZN(n8771) );
  NAND2_X1 U9430 ( .A1(n8991), .A2(n7021), .ZN(n7018) );
  OAI21_X1 U9431 ( .B1(n8803), .B2(n8622), .A(n8623), .ZN(n8815) );
  NAND2_X1 U9432 ( .A1(n8926), .A2(n7033), .ZN(n7030) );
  NAND2_X1 U9433 ( .A1(n12723), .A2(n12382), .ZN(n9045) );
  NAND2_X1 U9434 ( .A1(n12734), .A2(n12306), .ZN(n7038) );
  NOR2_X2 U9435 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n8737) );
  NAND3_X1 U9436 ( .A1(n10101), .A2(n7044), .A3(n8743), .ZN(n12203) );
  OR2_X1 U9437 ( .A1(n8731), .A2(n7047), .ZN(n7046) );
  AND3_X1 U9438 ( .A1(n8742), .A2(n7046), .A3(n7045), .ZN(n7044) );
  INV_X1 U9439 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n7047) );
  OAI21_X1 U9440 ( .B1(n11438), .B2(n7059), .A(n7054), .ZN(n12814) );
  NAND3_X1 U9441 ( .A1(n8902), .A2(n7448), .A3(n7442), .ZN(n9137) );
  NAND2_X1 U9442 ( .A1(n8902), .A2(n8588), .ZN(n8904) );
  AND2_X4 U9443 ( .A1(n8786), .A2(n8587), .ZN(n8902) );
  NAND2_X1 U9444 ( .A1(n12475), .A2(n7077), .ZN(n7075) );
  OAI21_X1 U9445 ( .B1(n10451), .B2(n7081), .A(n7080), .ZN(n10489) );
  OR2_X1 U9446 ( .A1(n7082), .A2(n7087), .ZN(n7080) );
  OR2_X1 U9447 ( .A1(n10449), .A2(n10051), .ZN(n7089) );
  NAND2_X1 U9448 ( .A1(n10448), .A2(n10602), .ZN(n7092) );
  NAND2_X2 U9449 ( .A1(n10042), .A2(n10041), .ZN(n10448) );
  NAND3_X1 U9450 ( .A1(n10042), .A2(n10041), .A3(n10052), .ZN(n7091) );
  INV_X1 U9451 ( .A(n10448), .ZN(n12153) );
  NAND2_X1 U9452 ( .A1(n10098), .A2(n7093), .ZN(n10047) );
  NOR2_X1 U9453 ( .A1(n7090), .A2(n10052), .ZN(n7094) );
  NAND2_X1 U9454 ( .A1(n12484), .A2(n6455), .ZN(n7096) );
  OAI21_X1 U9455 ( .B1(n11254), .B2(n6557), .A(n7101), .ZN(n11420) );
  INV_X1 U9456 ( .A(n11254), .ZN(n7105) );
  NOR2_X1 U9457 ( .A1(n11254), .A2(n11253), .ZN(n11256) );
  OAI21_X2 U9458 ( .B1(n10707), .B2(n12555), .A(n10706), .ZN(n10782) );
  NOR2_X4 U9459 ( .A1(n14755), .A2(n11895), .ZN(n14736) );
  NOR2_X4 U9460 ( .A1(n11017), .A2(n11939), .ZN(n11029) );
  NOR2_X2 U9461 ( .A1(n11346), .A2(n13843), .ZN(n14067) );
  NOR2_X2 U9462 ( .A1(n8288), .A2(n8287), .ZN(n14396) );
  INV_X1 U9463 ( .A(n15177), .ZN(n7115) );
  NOR2_X2 U9464 ( .A1(n14386), .A2(n8276), .ZN(n15175) );
  AOI21_X2 U9465 ( .B1(n7126), .B2(n7125), .A(n7124), .ZN(n8206) );
  NAND2_X2 U9466 ( .A1(n7468), .A2(n7679), .ZN(n7879) );
  NOR2_X1 U9467 ( .A1(n8319), .A2(n9578), .ZN(n9728) );
  NAND2_X1 U9468 ( .A1(n11570), .A2(n11569), .ZN(n13235) );
  NAND2_X1 U9469 ( .A1(n11570), .A2(n7127), .ZN(n7128) );
  OR2_X1 U9470 ( .A1(n13237), .A2(n13432), .ZN(n7129) );
  NAND3_X1 U9471 ( .A1(n7129), .A2(n13505), .A3(n7128), .ZN(n13431) );
  NOR2_X2 U9472 ( .A1(n10402), .A2(n10424), .ZN(n10433) );
  NOR2_X2 U9473 ( .A1(n9936), .A2(n10274), .ZN(n10017) );
  NOR2_X2 U9474 ( .A1(n13408), .A2(n13488), .ZN(n13396) );
  NOR2_X2 U9475 ( .A1(n11269), .A2(n13504), .ZN(n7134) );
  NOR2_X2 U9476 ( .A1(n10909), .A2(n11146), .ZN(n7136) );
  NOR3_X4 U9477 ( .A1(n13340), .A2(n7139), .A3(n13451), .ZN(n13280) );
  INV_X1 U9478 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7141) );
  NAND2_X1 U9479 ( .A1(n7556), .A2(n7142), .ZN(n9951) );
  NOR3_X1 U9480 ( .A1(n9946), .A2(n9945), .A3(n7142), .ZN(n9947) );
  XNOR2_X1 U9481 ( .A(n7558), .B(n7557), .ZN(n7142) );
  INV_X1 U9482 ( .A(n14501), .ZN(n7159) );
  NOR2_X2 U9483 ( .A1(n9571), .A2(n9462), .ZN(n13505) );
  OR2_X1 U9484 ( .A1(n10891), .A2(n13694), .ZN(n7167) );
  OAI21_X1 U9485 ( .B1(n14044), .B2(n13847), .A(n13846), .ZN(n14026) );
  NAND3_X1 U9486 ( .A1(n9247), .A2(n7176), .A3(n9246), .ZN(n14217) );
  NAND2_X1 U9487 ( .A1(n13893), .A2(n7177), .ZN(n13882) );
  NAND2_X1 U9488 ( .A1(n11284), .A2(n7181), .ZN(n7184) );
  INV_X1 U9489 ( .A(n7184), .ZN(n14076) );
  NAND2_X1 U9490 ( .A1(n14723), .A2(n11895), .ZN(n14725) );
  AND3_X2 U9491 ( .A1(n10132), .A2(n10134), .A3(n7191), .ZN(n14723) );
  AND2_X1 U9492 ( .A1(n10131), .A2(n10133), .ZN(n7191) );
  XNOR2_X2 U9493 ( .A(n13097), .B(n8312), .ZN(n9582) );
  NAND2_X1 U9494 ( .A1(n11144), .A2(n7203), .ZN(n7201) );
  OAI21_X1 U9495 ( .B1(n7216), .B2(n9930), .A(n10021), .ZN(n7215) );
  NAND2_X1 U9496 ( .A1(n7220), .A2(n7221), .ZN(n13419) );
  NAND2_X1 U9497 ( .A1(n10483), .A2(n6456), .ZN(n7224) );
  NAND2_X1 U9498 ( .A1(n7224), .A2(n6563), .ZN(n10907) );
  NAND2_X1 U9499 ( .A1(n7537), .A2(n7236), .ZN(n7542) );
  NAND2_X1 U9500 ( .A1(n7510), .A2(SI_1_), .ZN(n7236) );
  NAND2_X1 U9501 ( .A1(n7249), .A2(n7964), .ZN(n7250) );
  NAND3_X1 U9502 ( .A1(n7250), .A2(n12022), .A3(n7946), .ZN(n11629) );
  AND2_X1 U9503 ( .A1(n7250), .A2(n7946), .ZN(n11625) );
  INV_X1 U9504 ( .A(n7964), .ZN(n7251) );
  NAND3_X1 U9505 ( .A1(n12021), .A2(n12020), .A3(n6566), .ZN(n7253) );
  NAND2_X1 U9506 ( .A1(n7253), .A2(n7254), .ZN(n12077) );
  NAND2_X1 U9507 ( .A1(n7255), .A2(n7256), .ZN(n12011) );
  NAND3_X1 U9508 ( .A1(n12006), .A2(n6574), .A3(n12005), .ZN(n7255) );
  NAND2_X1 U9509 ( .A1(n7257), .A2(n7258), .ZN(n12001) );
  NAND3_X1 U9510 ( .A1(n7260), .A2(n7259), .A3(P1_DATAO_REG_1__SCAN_IN), .ZN(
        n7508) );
  NAND2_X1 U9511 ( .A1(n7904), .A2(n9968), .ZN(n7262) );
  INV_X1 U9512 ( .A(n9275), .ZN(n7263) );
  OAI21_X2 U9513 ( .B1(n13634), .B2(n7266), .A(n7264), .ZN(n13642) );
  NAND2_X1 U9514 ( .A1(n10219), .A2(n7270), .ZN(n10319) );
  NOR2_X1 U9515 ( .A1(n11396), .A2(n7282), .ZN(n11402) );
  NAND2_X1 U9516 ( .A1(n11397), .A2(n11398), .ZN(n7283) );
  NAND2_X1 U9517 ( .A1(n9261), .A2(n9219), .ZN(n9254) );
  NAND2_X1 U9518 ( .A1(n10819), .A2(n7287), .ZN(n7286) );
  NAND2_X1 U9519 ( .A1(n10819), .A2(n10818), .ZN(n10820) );
  INV_X1 U9520 ( .A(n7286), .ZN(n10975) );
  NOR2_X1 U9521 ( .A1(n10821), .A2(n7288), .ZN(n7287) );
  INV_X1 U9522 ( .A(n10818), .ZN(n7288) );
  NAND2_X1 U9523 ( .A1(n10976), .A2(n10977), .ZN(n7289) );
  NAND3_X1 U9524 ( .A1(n7291), .A2(n7290), .A3(n9218), .ZN(n9495) );
  NOR2_X2 U9525 ( .A1(n9260), .A2(n9602), .ZN(n9514) );
  NAND2_X1 U9526 ( .A1(n7303), .A2(n10766), .ZN(n14728) );
  NAND2_X1 U9527 ( .A1(n14726), .A2(n14725), .ZN(n7303) );
  INV_X1 U9528 ( .A(n10794), .ZN(n7304) );
  INV_X1 U9529 ( .A(n14725), .ZN(n7305) );
  NOR2_X1 U9530 ( .A1(n13244), .A2(n13249), .ZN(n13243) );
  NAND4_X1 U9531 ( .A1(n7332), .A2(n7330), .A3(n7336), .A4(n7329), .ZN(
        P2_U3528) );
  NAND2_X1 U9532 ( .A1(n7331), .A2(n6599), .ZN(n7330) );
  INV_X1 U9533 ( .A(n13436), .ZN(n7331) );
  OR2_X1 U9534 ( .A1(n14933), .A2(n7337), .ZN(n7336) );
  OAI21_X1 U9535 ( .B1(n7343), .B2(n7342), .A(n10471), .ZN(n7341) );
  NOR2_X1 U9536 ( .A1(n10422), .A2(n7344), .ZN(n7343) );
  OAI21_X2 U9537 ( .B1(n11387), .B2(n7348), .A(n7345), .ZN(n13404) );
  NAND2_X1 U9538 ( .A1(n7355), .A2(n13347), .ZN(n7354) );
  OAI21_X1 U9539 ( .B1(n10674), .B2(n7360), .A(n7358), .ZN(n11148) );
  INV_X1 U9540 ( .A(n8446), .ZN(n7365) );
  NOR2_X1 U9541 ( .A1(n8347), .A2(n7368), .ZN(n7367) );
  INV_X1 U9542 ( .A(n8343), .ZN(n7368) );
  NAND3_X1 U9543 ( .A1(n8403), .A2(n8402), .A3(n6594), .ZN(n7370) );
  NAND2_X1 U9544 ( .A1(n7370), .A2(n6592), .ZN(n8413) );
  INV_X1 U9545 ( .A(n8407), .ZN(n7371) );
  INV_X1 U9546 ( .A(n8406), .ZN(n7372) );
  NAND3_X1 U9547 ( .A1(n7376), .A2(n6457), .A3(n6492), .ZN(n7373) );
  INV_X1 U9548 ( .A(n8452), .ZN(n7376) );
  INV_X1 U9549 ( .A(n8455), .ZN(n7377) );
  NAND2_X1 U9550 ( .A1(n7379), .A2(n7378), .ZN(n8339) );
  OR2_X1 U9551 ( .A1(n8333), .A2(n8334), .ZN(n7378) );
  NAND3_X1 U9552 ( .A1(n7380), .A2(n8329), .A3(n8330), .ZN(n7379) );
  NAND2_X1 U9553 ( .A1(n7381), .A2(n6593), .ZN(n8425) );
  NAND2_X1 U9554 ( .A1(n7384), .A2(n7385), .ZN(n8547) );
  OAI21_X1 U9555 ( .B1(n8370), .B2(n7394), .A(n7393), .ZN(n7392) );
  AND2_X2 U9556 ( .A1(n7407), .A2(n7404), .ZN(n12719) );
  OR2_X2 U9557 ( .A1(n12756), .A2(n7408), .ZN(n7407) );
  NAND2_X1 U9558 ( .A1(n11065), .A2(n7418), .ZN(n7417) );
  NAND2_X2 U9559 ( .A1(n7417), .A2(n7414), .ZN(n11217) );
  OAI21_X1 U9560 ( .B1(n12243), .B2(n7424), .A(n12246), .ZN(n7423) );
  NAND2_X1 U9561 ( .A1(n9110), .A2(n7425), .ZN(n7424) );
  INV_X1 U9562 ( .A(n12549), .ZN(n7425) );
  OR2_X1 U9563 ( .A1(n8756), .A2(n9346), .ZN(n7427) );
  NAND3_X1 U9564 ( .A1(n7429), .A2(n8584), .A3(n8737), .ZN(n8787) );
  NAND3_X1 U9565 ( .A1(n10441), .A2(n9101), .A3(n12361), .ZN(n10622) );
  NAND2_X1 U9566 ( .A1(n9118), .A2(n9122), .ZN(n7431) );
  NAND2_X1 U9567 ( .A1(n11504), .A2(n9122), .ZN(n9178) );
  INV_X1 U9568 ( .A(n9118), .ZN(n11505) );
  INV_X1 U9569 ( .A(n7444), .ZN(n8680) );
  NAND2_X1 U9570 ( .A1(n10572), .A2(n10571), .ZN(n10819) );
  OAI21_X2 U9571 ( .B1(n8303), .B2(n7489), .A(n13226), .ZN(n9458) );
  INV_X1 U9572 ( .A(n14027), .ZN(n13848) );
  INV_X1 U9573 ( .A(n10165), .ZN(n10162) );
  OR2_X1 U9574 ( .A1(n9406), .A2(n11334), .ZN(n9512) );
  OAI211_X1 U9575 ( .C1(n11168), .C2(n9397), .A(n11334), .B(n9396), .ZN(n9675)
         );
  NAND2_X1 U9576 ( .A1(n8006), .A2(n8005), .ZN(n8008) );
  NAND2_X1 U9577 ( .A1(n11842), .A2(n11844), .ZN(n14685) );
  AND2_X1 U9578 ( .A1(n9264), .A2(n9254), .ZN(n9602) );
  AND2_X2 U9579 ( .A1(n10020), .A2(n10019), .ZN(n10023) );
  NAND2_X1 U9580 ( .A1(n10920), .A2(n11050), .ZN(n11052) );
  NAND2_X1 U9581 ( .A1(n10919), .A2(n10918), .ZN(n10920) );
  NAND2_X1 U9582 ( .A1(n12087), .A2(n7451), .ZN(n12827) );
  OAI21_X2 U9583 ( .B1(n12148), .B2(n12542), .A(n12432), .ZN(n12484) );
  NAND2_X1 U9584 ( .A1(n11506), .A2(n12766), .ZN(n11516) );
  MUX2_X2 U9585 ( .A(P3_REG0_REG_28__SCAN_IN), .B(n9174), .S(n15158), .Z(n9175) );
  NAND2_X2 U9586 ( .A1(n10686), .A2(n12034), .ZN(n14743) );
  NAND2_X1 U9587 ( .A1(n11879), .A2(n10649), .ZN(n10656) );
  OR2_X1 U9588 ( .A1(n7478), .A2(n7475), .ZN(n7477) );
  NAND2_X1 U9589 ( .A1(n9465), .A2(n9857), .ZN(n8557) );
  AOI22_X1 U9590 ( .A1(n10782), .A2(n10781), .B1(n10780), .B2(n10834), .ZN(
        n10784) );
  INV_X1 U9591 ( .A(n9882), .ZN(n11836) );
  NOR2_X2 U9592 ( .A1(n10312), .A2(n9240), .ZN(n9272) );
  INV_X1 U9593 ( .A(n7522), .ZN(n13546) );
  NAND2_X1 U9594 ( .A1(n13700), .A2(n9765), .ZN(n9695) );
  NAND2_X1 U9595 ( .A1(n8714), .A2(n12935), .ZN(n8729) );
  OR2_X1 U9596 ( .A1(n12422), .A2(n12926), .ZN(n7445) );
  OR2_X1 U9597 ( .A1(n9177), .A2(n12926), .ZN(n7446) );
  AND3_X1 U9598 ( .A1(n11638), .A2(n11637), .A3(n11636), .ZN(n14054) );
  INV_X1 U9599 ( .A(n11201), .ZN(n11212) );
  OR2_X1 U9600 ( .A1(n12422), .A2(n12876), .ZN(n7447) );
  OR2_X1 U9601 ( .A1(n13841), .A2(n13840), .ZN(n7450) );
  OR2_X1 U9602 ( .A1(n12086), .A2(n15146), .ZN(n7451) );
  INV_X1 U9603 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9220) );
  INV_X1 U9604 ( .A(n13444), .ZN(n13265) );
  AND2_X1 U9605 ( .A1(n9244), .A2(n9271), .ZN(n7453) );
  OR2_X1 U9606 ( .A1(n11871), .A2(n12072), .ZN(n7454) );
  INV_X1 U9607 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7509) );
  INV_X1 U9608 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9269) );
  CLKBUF_X2 U9609 ( .A(P1_U4016), .Z(n13701) );
  INV_X1 U9610 ( .A(n14105), .ZN(n13899) );
  AND2_X1 U9611 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n7455) );
  NAND2_X2 U9612 ( .A1(n13869), .A2(n14751), .ZN(n14691) );
  INV_X1 U9613 ( .A(n9421), .ZN(n9410) );
  AND2_X1 U9614 ( .A1(n8360), .A2(n8359), .ZN(n7456) );
  XNOR2_X1 U9615 ( .A(n13226), .B(n8573), .ZN(n7457) );
  AND3_X1 U9616 ( .A1(n8538), .A2(n8537), .A3(n8536), .ZN(n7459) );
  AND2_X1 U9617 ( .A1(n13472), .A2(n12987), .ZN(n7460) );
  AND2_X1 U9618 ( .A1(n8374), .A2(n8373), .ZN(n7461) );
  INV_X1 U9619 ( .A(n14693), .ZN(n10753) );
  INV_X1 U9620 ( .A(n8308), .ZN(n8307) );
  AOI21_X1 U9621 ( .B1(n8370), .B2(n8369), .A(n8367), .ZN(n8368) );
  INV_X1 U9622 ( .A(n8419), .ZN(n8420) );
  OR2_X1 U9623 ( .A1(n11991), .A2(n11990), .ZN(n11992) );
  INV_X1 U9624 ( .A(n8432), .ZN(n8433) );
  NAND2_X1 U9625 ( .A1(n8436), .A2(n8435), .ZN(n8441) );
  INV_X1 U9626 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8677) );
  INV_X1 U9627 ( .A(n8021), .ZN(n8027) );
  INV_X1 U9628 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9244) );
  NAND2_X1 U9629 ( .A1(n12400), .A2(n12878), .ZN(n12401) );
  INV_X1 U9630 ( .A(n8972), .ZN(n8699) );
  OR2_X1 U9631 ( .A1(n8103), .A2(n11195), .ZN(n8104) );
  NAND2_X1 U9632 ( .A1(n12386), .A2(n12401), .ZN(n12402) );
  INV_X1 U9633 ( .A(n9032), .ZN(n8704) );
  INV_X1 U9634 ( .A(n14952), .ZN(n10534) );
  INV_X1 U9635 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n14291) );
  INV_X1 U9636 ( .A(n12320), .ZN(n9119) );
  OR2_X1 U9637 ( .A1(n9040), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9049) );
  INV_X1 U9638 ( .A(n8959), .ZN(n8698) );
  INV_X1 U9639 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8681) );
  INV_X1 U9640 ( .A(n7952), .ZN(n7951) );
  AND2_X1 U9641 ( .A1(n7731), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7748) );
  NAND2_X1 U9642 ( .A1(n11199), .A2(n11198), .ZN(n11276) );
  INV_X1 U9643 ( .A(n11744), .ZN(n11742) );
  INV_X1 U9644 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10876) );
  INV_X1 U9645 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10171) );
  OR2_X1 U9646 ( .A1(n10743), .A2(n12036), .ZN(n10744) );
  INV_X1 U9647 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9223) );
  INV_X1 U9648 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9219) );
  INV_X1 U9649 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9206) );
  INV_X1 U9650 ( .A(n9007), .ZN(n8702) );
  OR2_X1 U9651 ( .A1(n9049), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9061) );
  NAND2_X1 U9652 ( .A1(n8704), .A2(n8703), .ZN(n9040) );
  INV_X1 U9653 ( .A(n12564), .ZN(n12562) );
  INV_X1 U9654 ( .A(n12537), .ZN(n11510) );
  NAND2_X1 U9655 ( .A1(n8983), .A2(n8700), .ZN(n8996) );
  NAND2_X1 U9656 ( .A1(n8694), .A2(n8693), .ZN(n8930) );
  INV_X1 U9657 ( .A(n7990), .ZN(n7988) );
  INV_X1 U9658 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7637) );
  OR2_X1 U9659 ( .A1(n8110), .A2(n8109), .ZN(n8121) );
  OR2_X1 U9660 ( .A1(n7971), .A2(n12986), .ZN(n7990) );
  NAND2_X1 U9661 ( .A1(n7951), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n7971) );
  OR2_X1 U9662 ( .A1(n7776), .A2(n7775), .ZN(n7802) );
  AND2_X1 U9663 ( .A1(n10367), .A2(n10366), .ZN(n10504) );
  AND2_X1 U9664 ( .A1(n9435), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9438) );
  OR2_X1 U9665 ( .A1(n8087), .A2(n13067), .ZN(n8110) );
  INV_X1 U9666 ( .A(n13308), .ZN(n11553) );
  OR2_X1 U9667 ( .A1(n7688), .A2(n7687), .ZN(n7710) );
  INV_X1 U9668 ( .A(n11579), .ZN(n11580) );
  INV_X1 U9669 ( .A(n10815), .ZN(n10816) );
  INV_X1 U9670 ( .A(n11447), .ZN(n11450) );
  NAND2_X1 U9671 ( .A1(n11742), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n11765) );
  OR2_X1 U9672 ( .A1(n11631), .A2(n11630), .ZN(n11651) );
  NAND2_X1 U9673 ( .A1(n14115), .A2(n14105), .ZN(n13860) );
  INV_X1 U9674 ( .A(n13896), .ZN(n13859) );
  NAND2_X1 U9675 ( .A1(n11288), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n11309) );
  INV_X1 U9676 ( .A(n11840), .ZN(n9601) );
  OR2_X1 U9677 ( .A1(n11939), .A2(n13692), .ZN(n11023) );
  NAND2_X1 U9678 ( .A1(n7791), .A2(SI_13_), .ZN(n7816) );
  INV_X1 U9679 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9361) );
  NOR2_X1 U9680 ( .A1(n8247), .A2(n8246), .ZN(n8227) );
  OR2_X1 U9681 ( .A1(n10917), .A2(n10921), .ZN(n10918) );
  NAND2_X1 U9682 ( .A1(n8702), .A2(n8701), .ZN(n9021) );
  OR2_X1 U9683 ( .A1(n10050), .A2(n9879), .ZN(n12527) );
  XNOR2_X1 U9684 ( .A(n12405), .B(n12404), .ZN(n12407) );
  INV_X1 U9685 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n10709) );
  INV_X1 U9686 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n11183) );
  AND2_X1 U9687 ( .A1(n9839), .A2(n9838), .ZN(n9850) );
  AND2_X1 U9688 ( .A1(n12264), .A2(n12269), .ZN(n12373) );
  INV_X1 U9689 ( .A(n15134), .ZN(n12816) );
  OR2_X1 U9690 ( .A1(n10584), .A2(n10040), .ZN(n9168) );
  INV_X1 U9691 ( .A(n12670), .ZN(n9177) );
  OR2_X1 U9692 ( .A1(n10049), .A2(n12317), .ZN(n12799) );
  INV_X1 U9693 ( .A(n10442), .ZN(n12363) );
  INV_X1 U9694 ( .A(n10303), .ZN(n12367) );
  NOR2_X1 U9695 ( .A1(n9171), .A2(n9170), .ZN(n9896) );
  OAI21_X1 U9696 ( .B1(n9160), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9162) );
  AND2_X1 U9697 ( .A1(n8657), .A2(n8655), .ZN(n9003) );
  XNOR2_X1 U9698 ( .A(n9364), .B(P1_DATAO_REG_5__SCAN_IN), .ZN(n8784) );
  NAND2_X1 U9699 ( .A1(n7988), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8043) );
  INV_X1 U9700 ( .A(n7842), .ZN(n7841) );
  INV_X1 U9701 ( .A(n8050), .ZN(n9856) );
  INV_X1 U9702 ( .A(n13029), .ZN(n7814) );
  OR2_X1 U9703 ( .A1(n8193), .A2(n8577), .ZN(n13066) );
  NOR2_X1 U9704 ( .A1(n8121), .A2(n8120), .ZN(n11565) );
  INV_X1 U9705 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n14854) );
  NAND2_X1 U9706 ( .A1(n13074), .A2(n13370), .ZN(n11540) );
  INV_X1 U9707 ( .A(n13084), .ZN(n14499) );
  INV_X1 U9708 ( .A(n13381), .ZN(n13415) );
  OAI21_X1 U9709 ( .B1(P2_D_REG_1__SCAN_IN), .B2(n8163), .A(n14908), .ZN(n9995) );
  AND2_X1 U9710 ( .A1(n7765), .A2(n7764), .ZN(n7769) );
  NAND2_X1 U9711 ( .A1(n11581), .A2(n11580), .ZN(n11582) );
  NAND2_X1 U9712 ( .A1(n11127), .A2(n11129), .ZN(n11130) );
  INV_X1 U9713 ( .A(n13925), .ZN(n13832) );
  NAND2_X1 U9714 ( .A1(n10817), .A2(n10816), .ZN(n10818) );
  INV_X1 U9715 ( .A(n13924), .ZN(n13960) );
  OR2_X1 U9716 ( .A1(n12077), .A2(n12076), .ZN(n12078) );
  NOR2_X1 U9717 ( .A1(n11651), .A2(n13637), .ZN(n11663) );
  INV_X1 U9718 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n11136) );
  OR2_X1 U9719 ( .A1(n14587), .A2(n9302), .ZN(n14669) );
  INV_X1 U9720 ( .A(n13858), .ZN(n13922) );
  INV_X1 U9721 ( .A(n12050), .ZN(n14061) );
  INV_X1 U9722 ( .A(n13693), .ZN(n11405) );
  NAND2_X1 U9723 ( .A1(n14693), .A2(n14703), .ZN(n10755) );
  NAND2_X1 U9724 ( .A1(n13699), .A2(n6952), .ZN(n11887) );
  INV_X1 U9725 ( .A(n13992), .ZN(n13999) );
  NAND2_X1 U9726 ( .A1(n9603), .A2(n10662), .ZN(n14792) );
  INV_X1 U9727 ( .A(n13692), .ZN(n11239) );
  INV_X1 U9728 ( .A(n12039), .ZN(n14700) );
  OR2_X1 U9729 ( .A1(n9675), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9513) );
  XNOR2_X1 U9730 ( .A(n7900), .B(n9757), .ZN(n7898) );
  XNOR2_X1 U9731 ( .A(n7832), .B(SI_14_), .ZN(n7835) );
  NAND2_X1 U9732 ( .A1(n7580), .A2(n7579), .ZN(n7603) );
  AOI22_X1 U9733 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14613), .B1(n8245), .B2(
        n8229), .ZN(n8242) );
  NAND2_X1 U9734 ( .A1(n11052), .A2(n11051), .ZN(n11054) );
  AND2_X1 U9735 ( .A1(n12353), .A2(n12352), .ZN(n12660) );
  AND2_X1 U9736 ( .A1(n9079), .A2(n9078), .ZN(n12453) );
  INV_X1 U9737 ( .A(n15109), .ZN(n15090) );
  INV_X1 U9738 ( .A(n15101), .ZN(n15000) );
  INV_X1 U9739 ( .A(n12815), .ZN(n14471) );
  AND2_X1 U9740 ( .A1(n12255), .A2(n12256), .ZN(n12372) );
  AND2_X1 U9741 ( .A1(n9109), .A2(n12237), .ZN(n12360) );
  AND2_X1 U9742 ( .A1(n10589), .A2(n10603), .ZN(n15134) );
  AND3_X1 U9743 ( .A1(n9168), .A2(n9163), .A3(n9171), .ZN(n10587) );
  AND3_X1 U9744 ( .A1(n8894), .A2(n8893), .A3(n8892), .ZN(n12246) );
  AND2_X1 U9745 ( .A1(n10603), .A2(n9134), .ZN(n15143) );
  OR2_X1 U9746 ( .A1(n15125), .A2(n15143), .ZN(n15150) );
  NAND2_X1 U9747 ( .A1(n8952), .A2(n8646), .ZN(n8966) );
  INV_X1 U9748 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8817) );
  INV_X1 U9749 ( .A(n13081), .ZN(n11391) );
  NOR2_X1 U9750 ( .A1(n7457), .A2(n8574), .ZN(n8575) );
  OR2_X1 U9751 ( .A1(n13252), .A2(n8124), .ZN(n8129) );
  NAND2_X1 U9752 ( .A1(n7591), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n7524) );
  INV_X1 U9753 ( .A(n14862), .ZN(n13184) );
  OR2_X1 U9754 ( .A1(n9441), .A2(n11538), .ZN(n14856) );
  NOR2_X1 U9755 ( .A1(n9440), .A2(n9439), .ZN(n14862) );
  AND2_X1 U9756 ( .A1(n9442), .A2(n11538), .ZN(n13224) );
  OR2_X1 U9757 ( .A1(n9464), .A2(n9463), .ZN(n13406) );
  OR2_X1 U9758 ( .A1(n14872), .A2(n9457), .ZN(n13377) );
  AND2_X1 U9759 ( .A1(n13394), .A2(n13226), .ZN(n13424) );
  AND2_X1 U9760 ( .A1(n13394), .A2(n10002), .ZN(n13381) );
  AND2_X1 U9761 ( .A1(n9458), .A2(n10420), .ZN(n13516) );
  INV_X1 U9762 ( .A(n13516), .ZN(n14533) );
  INV_X1 U9763 ( .A(n10420), .ZN(n14927) );
  NAND2_X1 U9764 ( .A1(n9432), .A2(n14905), .ZN(n14872) );
  AND2_X1 U9765 ( .A1(n7613), .A2(n7657), .ZN(n13125) );
  INV_X1 U9766 ( .A(n13688), .ZN(n13645) );
  OAI211_X1 U9767 ( .C1(n7454), .C2(n12079), .A(n7458), .B(n12078), .ZN(n12080) );
  OR2_X1 U9768 ( .A1(n9605), .A2(n13906), .ZN(n11784) );
  OR2_X1 U9769 ( .A1(n9605), .A2(n13628), .ZN(n11726) );
  OR2_X1 U9770 ( .A1(n14587), .A2(n9707), .ZN(n14618) );
  OR2_X1 U9771 ( .A1(n14587), .A2(n14582), .ZN(n14665) );
  INV_X1 U9772 ( .A(n14669), .ZN(n14633) );
  INV_X1 U9773 ( .A(n14618), .ZN(n14676) );
  INV_X1 U9774 ( .A(n13829), .ZN(n13958) );
  INV_X1 U9775 ( .A(n14161), .ZN(n14012) );
  INV_X1 U9776 ( .A(n14695), .ZN(n14759) );
  INV_X1 U9777 ( .A(n9680), .ZN(n10639) );
  INV_X1 U9778 ( .A(n14824), .ZN(n14197) );
  NAND2_X1 U9779 ( .A1(n10791), .A2(n14797), .ZN(n14824) );
  NAND2_X1 U9780 ( .A1(n9513), .A2(n9512), .ZN(n9680) );
  AND2_X1 U9781 ( .A1(n9363), .A2(n9379), .ZN(n13734) );
  AND3_X1 U9782 ( .A1(n9159), .A2(n9158), .A3(n9157), .ZN(n9886) );
  NAND2_X1 U9783 ( .A1(n9881), .A2(n10589), .ZN(n12528) );
  NAND2_X1 U9784 ( .A1(n9878), .A2(n9877), .ZN(n12534) );
  INV_X1 U9785 ( .A(n12676), .ZN(n12538) );
  INV_X1 U9786 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n15007) );
  INV_X1 U9787 ( .A(n14960), .ZN(n15116) );
  AND2_X1 U9788 ( .A1(n11221), .A2(n11220), .ZN(n14490) );
  INV_X1 U9789 ( .A(n12821), .ZN(n12666) );
  NAND2_X1 U9790 ( .A1(n15166), .A2(n15152), .ZN(n12876) );
  NAND2_X1 U9791 ( .A1(n9164), .A2(n10587), .ZN(n15164) );
  INV_X1 U9792 ( .A(n12439), .ZN(n12910) );
  AND2_X1 U9793 ( .A1(n14490), .A2(n14489), .ZN(n14498) );
  AND2_X1 U9794 ( .A1(n9173), .A2(n9172), .ZN(n15157) );
  AND2_X1 U9795 ( .A1(n9423), .A2(n9395), .ZN(n9421) );
  NAND2_X1 U9796 ( .A1(n9885), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9386) );
  INV_X1 U9797 ( .A(SI_18_), .ZN(n9968) );
  INV_X1 U9798 ( .A(SI_13_), .ZN(n9412) );
  NAND2_X1 U9799 ( .A1(n8833), .A2(n8832), .ZN(n12609) );
  INV_X1 U9800 ( .A(n10521), .ZN(n10545) );
  INV_X1 U9801 ( .A(n8200), .ZN(n8201) );
  INV_X1 U9802 ( .A(n14507), .ZN(n14515) );
  NAND2_X1 U9803 ( .A1(n8576), .A2(n8575), .ZN(n8582) );
  NAND2_X1 U9804 ( .A1(n8117), .A2(n8116), .ZN(n13075) );
  OR2_X1 U9805 ( .A1(n7808), .A2(n7807), .ZN(n13084) );
  INV_X1 U9806 ( .A(n13224), .ZN(n14864) );
  NAND2_X1 U9807 ( .A1(n13394), .A2(n10058), .ZN(n13421) );
  AND3_X2 U9808 ( .A1(n9996), .A2(n9642), .A3(n9994), .ZN(n14933) );
  OR2_X1 U9809 ( .A1(n13510), .A2(n13509), .ZN(n13536) );
  NOR2_X1 U9810 ( .A1(n14873), .A2(n14872), .ZN(n14888) );
  CLKBUF_X1 U9811 ( .A(n14888), .Z(n14910) );
  INV_X1 U9812 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9594) );
  INV_X1 U9813 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9369) );
  INV_X1 U9814 ( .A(n11923), .ZN(n14815) );
  NAND4_X1 U9815 ( .A1(n11786), .A2(n11785), .A3(n11784), .A4(n11783), .ZN(
        n13925) );
  NAND2_X1 U9816 ( .A1(n11670), .A2(n11669), .ZN(n14017) );
  NOR2_X1 U9817 ( .A1(n9407), .A2(n10182), .ZN(P1_U4016) );
  INV_X1 U9818 ( .A(n13581), .ZN(n13699) );
  INV_X1 U9819 ( .A(n14585), .ZN(n14679) );
  INV_X1 U9820 ( .A(n14697), .ZN(n14059) );
  INV_X1 U9821 ( .A(n14839), .ZN(n14837) );
  INV_X1 U9822 ( .A(n14827), .ZN(n14826) );
  NAND2_X1 U9823 ( .A1(n9685), .A2(n9675), .ZN(n14765) );
  INV_X1 U9824 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10215) );
  AND2_X2 U9825 ( .A1(n9423), .A2(n9886), .ZN(P3_U3897) );
  AND2_X1 U9826 ( .A1(n14905), .A2(n9232), .ZN(P2_U3947) );
  NOR2_X1 U9827 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7465) );
  NAND4_X1 U9828 ( .A1(n7465), .A2(n7464), .A3(n7463), .A4(n7462), .ZN(n7858)
         );
  NOR2_X1 U9829 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n7466) );
  NAND2_X1 U9830 ( .A1(n7856), .A2(n7466), .ZN(n7467) );
  NOR2_X2 U9831 ( .A1(n7858), .A2(n7467), .ZN(n7468) );
  AND2_X2 U9832 ( .A1(n6463), .A2(n7548), .ZN(n7679) );
  NAND2_X1 U9833 ( .A1(n7476), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7473) );
  INV_X1 U9834 ( .A(n7478), .ZN(n7483) );
  AND2_X1 U9835 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n7481) );
  INV_X1 U9836 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n13538) );
  NAND2_X1 U9837 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .ZN(n7479) );
  AOI22_X1 U9838 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(n13538), .B1(n7479), .B2(
        P2_IR_REG_31__SCAN_IN), .ZN(n7480) );
  NAND2_X1 U9839 ( .A1(n7482), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7486) );
  INV_X1 U9840 ( .A(n7486), .ZN(n7484) );
  NAND2_X1 U9841 ( .A1(n7484), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n7488) );
  NAND2_X1 U9842 ( .A1(n7486), .A2(n7485), .ZN(n7487) );
  INV_X1 U9843 ( .A(n9999), .ZN(n7490) );
  INV_X1 U9844 ( .A(n7491), .ZN(n7494) );
  NOR2_X1 U9845 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n7493) );
  NOR2_X1 U9846 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n7492) );
  INV_X1 U9847 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7495) );
  NAND3_X1 U9848 ( .A1(n8141), .A2(n7500), .A3(n7495), .ZN(n7505) );
  INV_X1 U9849 ( .A(n7505), .ZN(n7496) );
  NAND2_X1 U9850 ( .A1(n7452), .A2(n7496), .ZN(n7497) );
  NAND3_X1 U9851 ( .A1(n8141), .A2(n7500), .A3(P2_IR_REG_27__SCAN_IN), .ZN(
        n7502) );
  XNOR2_X1 U9852 ( .A(P2_IR_REG_31__SCAN_IN), .B(P2_IR_REG_27__SCAN_IN), .ZN(
        n7501) );
  NAND2_X1 U9853 ( .A1(n7502), .A2(n7501), .ZN(n7503) );
  INV_X1 U9854 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n7507) );
  NAND2_X1 U9855 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7506) );
  OAI22_X1 U9856 ( .A1(n8487), .A2(n9355), .B1(n7771), .B2(n9526), .ZN(n7516)
         );
  OAI21_X2 U9857 ( .B1(n6448), .B2(n7509), .A(n7508), .ZN(n7510) );
  INV_X1 U9858 ( .A(n7514), .ZN(n7511) );
  INV_X1 U9859 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8725) );
  NAND2_X1 U9860 ( .A1(n7511), .A2(n7512), .ZN(n7537) );
  INV_X1 U9861 ( .A(n7512), .ZN(n7513) );
  NAND2_X1 U9862 ( .A1(n7514), .A2(n7513), .ZN(n7515) );
  NAND2_X1 U9863 ( .A1(n7537), .A2(n7515), .ZN(n9596) );
  NAND2_X1 U9864 ( .A1(n7571), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7527) );
  AND2_X4 U9865 ( .A1(n11576), .A2(n7522), .ZN(n8069) );
  NAND2_X1 U9866 ( .A1(n6447), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7526) );
  NAND2_X1 U9867 ( .A1(n8050), .A2(n13097), .ZN(n7534) );
  INV_X1 U9868 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9475) );
  NAND2_X1 U9869 ( .A1(n6436), .A2(SI_0_), .ZN(n7528) );
  XNOR2_X1 U9870 ( .A(n7528), .B(n8608), .ZN(n13552) );
  MUX2_X1 U9871 ( .A(n9475), .B(n13552), .S(n7771), .Z(n9857) );
  INV_X1 U9872 ( .A(n9857), .ZN(n10252) );
  OR2_X1 U9873 ( .A1(n7590), .A2(n10252), .ZN(n7533) );
  NAND2_X1 U9874 ( .A1(n6446), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7532) );
  NAND2_X1 U9875 ( .A1(n7571), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7529) );
  AND2_X1 U9876 ( .A1(n9859), .A2(n7533), .ZN(n9736) );
  INV_X1 U9877 ( .A(n9943), .ZN(n7535) );
  NAND2_X1 U9878 ( .A1(n7535), .A2(n7534), .ZN(n7536) );
  INV_X1 U9879 ( .A(n7542), .ZN(n7539) );
  NAND2_X1 U9880 ( .A1(n7538), .A2(SI_2_), .ZN(n7561) );
  OAI21_X1 U9881 ( .B1(n7538), .B2(SI_2_), .A(n7561), .ZN(n7540) );
  NAND2_X1 U9882 ( .A1(n7539), .A2(n7540), .ZN(n7543) );
  INV_X1 U9883 ( .A(n7540), .ZN(n7541) );
  NAND2_X1 U9884 ( .A1(n7542), .A2(n7541), .ZN(n7562) );
  NAND2_X1 U9885 ( .A1(n7543), .A2(n7562), .ZN(n9758) );
  NAND2_X1 U9886 ( .A1(n7544), .A2(n8509), .ZN(n7551) );
  INV_X1 U9887 ( .A(n7545), .ZN(n7546) );
  NAND2_X1 U9888 ( .A1(n7546), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7547) );
  MUX2_X1 U9889 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7547), .S(
        P2_IR_REG_2__SCAN_IN), .Z(n7549) );
  INV_X1 U9890 ( .A(n7548), .ZN(n7566) );
  NAND2_X1 U9891 ( .A1(n7549), .A2(n7566), .ZN(n9534) );
  INV_X1 U9892 ( .A(n9534), .ZN(n9551) );
  AOI22_X1 U9893 ( .A1(n7582), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n9428), .B2(
        n9551), .ZN(n7550) );
  XNOR2_X1 U9894 ( .A(n7590), .B(n8319), .ZN(n7557) );
  NAND2_X1 U9895 ( .A1(n8186), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7555) );
  NAND2_X1 U9896 ( .A1(n8069), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7554) );
  NAND2_X1 U9897 ( .A1(n7570), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7553) );
  NAND2_X1 U9898 ( .A1(n7571), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n7552) );
  NAND2_X1 U9899 ( .A1(n8050), .A2(n13095), .ZN(n7558) );
  INV_X1 U9900 ( .A(n7557), .ZN(n7559) );
  NAND2_X1 U9901 ( .A1(n7559), .A2(n7558), .ZN(n7560) );
  NAND2_X1 U9902 ( .A1(n7562), .A2(n7561), .ZN(n7578) );
  MUX2_X1 U9903 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n6450), .Z(n7564) );
  NAND2_X1 U9904 ( .A1(n7564), .A2(SI_3_), .ZN(n7579) );
  OAI21_X1 U9905 ( .B1(n7564), .B2(SI_3_), .A(n7579), .ZN(n7576) );
  XNOR2_X1 U9906 ( .A(n7578), .B(n7576), .ZN(n9365) );
  NAND2_X1 U9907 ( .A1(n9365), .A2(n8509), .ZN(n7569) );
  NAND2_X1 U9908 ( .A1(n7566), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7565) );
  MUX2_X1 U9909 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7565), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n7567) );
  AOI22_X1 U9910 ( .A1(n7582), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n9428), .B2(
        n13110), .ZN(n7568) );
  XNOR2_X1 U9911 ( .A(n7590), .B(n10006), .ZN(n9981) );
  INV_X1 U9912 ( .A(n7591), .ZN(n7572) );
  AND2_X1 U9913 ( .A1(n8050), .A2(n13094), .ZN(n7573) );
  NAND2_X1 U9914 ( .A1(n9981), .A2(n7573), .ZN(n7596) );
  OR2_X1 U9915 ( .A1(n9981), .A2(n7573), .ZN(n7574) );
  NAND2_X1 U9916 ( .A1(n7596), .A2(n7574), .ZN(n9823) );
  INV_X1 U9917 ( .A(n7576), .ZN(n7577) );
  NAND2_X1 U9918 ( .A1(n7578), .A2(n7577), .ZN(n7580) );
  NAND2_X1 U9919 ( .A1(n7581), .A2(SI_4_), .ZN(n7604) );
  OAI21_X1 U9920 ( .B1(n7581), .B2(SI_4_), .A(n7604), .ZN(n7601) );
  XNOR2_X1 U9921 ( .A(n7603), .B(n7601), .ZN(n10136) );
  NAND2_X1 U9922 ( .A1(n10136), .A2(n8509), .ZN(n7589) );
  NAND2_X1 U9923 ( .A1(n7584), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7583) );
  MUX2_X1 U9924 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7583), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n7587) );
  INV_X1 U9925 ( .A(n7584), .ZN(n7586) );
  INV_X1 U9926 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7585) );
  NAND2_X1 U9927 ( .A1(n7586), .A2(n7585), .ZN(n7612) );
  NAND2_X1 U9928 ( .A1(n7587), .A2(n7612), .ZN(n9554) );
  INV_X1 U9929 ( .A(n9554), .ZN(n14846) );
  AOI22_X1 U9930 ( .A1(n7582), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n9428), .B2(
        n14846), .ZN(n7588) );
  NAND2_X1 U9931 ( .A1(n8477), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n7595) );
  NAND2_X1 U9932 ( .A1(n8069), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7594) );
  NAND2_X1 U9933 ( .A1(n7570), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7593) );
  INV_X1 U9934 ( .A(n7616), .ZN(n7618) );
  OAI21_X1 U9935 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n7618), .ZN(n10069) );
  OR2_X1 U9936 ( .A1(n8124), .A2(n10069), .ZN(n7592) );
  NAND2_X1 U9937 ( .A1(n8050), .A2(n13093), .ZN(n7598) );
  INV_X1 U9938 ( .A(n9969), .ZN(n7599) );
  NAND2_X1 U9939 ( .A1(n7599), .A2(n7598), .ZN(n7600) );
  INV_X1 U9940 ( .A(n7601), .ZN(n7602) );
  NAND2_X1 U9941 ( .A1(n7603), .A2(n7602), .ZN(n7605) );
  INV_X1 U9942 ( .A(n7606), .ZN(n7607) );
  OR2_X1 U9943 ( .A1(n7608), .A2(n7607), .ZN(n7609) );
  NAND2_X1 U9944 ( .A1(n7630), .A2(n7609), .ZN(n10220) );
  OR2_X1 U9945 ( .A1(n10220), .A2(n7908), .ZN(n7615) );
  NAND2_X1 U9946 ( .A1(n7612), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7611) );
  MUX2_X1 U9947 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7611), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n7613) );
  AOI22_X1 U9948 ( .A1(n7582), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9428), .B2(
        n13125), .ZN(n7614) );
  NAND2_X1 U9949 ( .A1(n7615), .A2(n7614), .ZN(n9973) );
  XNOR2_X1 U9950 ( .A(n9973), .B(n8086), .ZN(n7625) );
  NAND2_X1 U9951 ( .A1(n8477), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7623) );
  NAND2_X1 U9952 ( .A1(n8069), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7622) );
  NAND2_X1 U9953 ( .A1(n6704), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7621) );
  NAND2_X1 U9954 ( .A1(n7616), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7638) );
  INV_X1 U9955 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7617) );
  NAND2_X1 U9956 ( .A1(n7618), .A2(n7617), .ZN(n7619) );
  NAND2_X1 U9957 ( .A1(n7638), .A2(n7619), .ZN(n10266) );
  OR2_X1 U9958 ( .A1(n7572), .A2(n10266), .ZN(n7620) );
  NAND4_X1 U9959 ( .A1(n7623), .A2(n7622), .A3(n7621), .A4(n7620), .ZN(n13092)
         );
  NAND2_X1 U9960 ( .A1(n8050), .A2(n13092), .ZN(n7626) );
  XNOR2_X1 U9961 ( .A(n7625), .B(n7626), .ZN(n9970) );
  INV_X1 U9962 ( .A(n7625), .ZN(n7627) );
  NAND2_X1 U9963 ( .A1(n7627), .A2(n7626), .ZN(n7628) );
  NAND2_X1 U9964 ( .A1(n7631), .A2(SI_6_), .ZN(n7650) );
  OAI21_X1 U9965 ( .B1(SI_6_), .B2(n7631), .A(n7650), .ZN(n7632) );
  NAND2_X1 U9966 ( .A1(n7657), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7634) );
  XNOR2_X1 U9967 ( .A(n7634), .B(P2_IR_REG_6__SCAN_IN), .ZN(n13142) );
  AOI22_X1 U9968 ( .A1(n7582), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9428), .B2(
        n13142), .ZN(n7635) );
  NAND2_X1 U9969 ( .A1(n8477), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n7643) );
  NAND2_X1 U9970 ( .A1(n8069), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7642) );
  NAND2_X1 U9971 ( .A1(n6704), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7641) );
  INV_X1 U9972 ( .A(n7661), .ZN(n7663) );
  NAND2_X1 U9973 ( .A1(n7638), .A2(n7637), .ZN(n7639) );
  NAND2_X1 U9974 ( .A1(n7663), .A2(n7639), .ZN(n10275) );
  OR2_X1 U9975 ( .A1(n8124), .A2(n10275), .ZN(n7640) );
  NAND4_X1 U9976 ( .A1(n7643), .A2(n7642), .A3(n7641), .A4(n7640), .ZN(n13091)
         );
  AND2_X1 U9977 ( .A1(n8050), .A2(n13091), .ZN(n7645) );
  NAND2_X1 U9978 ( .A1(n7644), .A2(n7645), .ZN(n7649) );
  INV_X1 U9979 ( .A(n7644), .ZN(n10030) );
  INV_X1 U9980 ( .A(n7645), .ZN(n7646) );
  NAND2_X1 U9981 ( .A1(n10030), .A2(n7646), .ZN(n7647) );
  MUX2_X1 U9982 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6450), .Z(n7652) );
  NAND2_X1 U9983 ( .A1(n7652), .A2(SI_7_), .ZN(n7672) );
  OAI21_X1 U9984 ( .B1(n7652), .B2(SI_7_), .A(n7672), .ZN(n7653) );
  INV_X1 U9985 ( .A(n7653), .ZN(n7654) );
  OR2_X1 U9986 ( .A1(n7655), .A2(n7654), .ZN(n7656) );
  NAND2_X1 U9987 ( .A1(n7673), .A2(n7656), .ZN(n10561) );
  OR2_X1 U9988 ( .A1(n10561), .A2(n7908), .ZN(n7660) );
  OAI21_X1 U9989 ( .B1(n7657), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7658) );
  XNOR2_X1 U9990 ( .A(n7658), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9660) );
  AOI22_X1 U9991 ( .A1(n8510), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n9428), .B2(
        n9660), .ZN(n7659) );
  XNOR2_X1 U9992 ( .A(n10289), .B(n8086), .ZN(n7669) );
  NAND2_X1 U9993 ( .A1(n8069), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7668) );
  NAND2_X1 U9994 ( .A1(n6704), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7667) );
  NAND2_X1 U9995 ( .A1(n8477), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7666) );
  NAND2_X1 U9996 ( .A1(n7661), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7688) );
  INV_X1 U9997 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7662) );
  NAND2_X1 U9998 ( .A1(n7663), .A2(n7662), .ZN(n7664) );
  NAND2_X1 U9999 ( .A1(n7688), .A2(n7664), .ZN(n10255) );
  OR2_X1 U10000 ( .A1(n8124), .A2(n10255), .ZN(n7665) );
  NAND4_X1 U10001 ( .A1(n7668), .A2(n7667), .A3(n7666), .A4(n7665), .ZN(n13090) );
  AND2_X1 U10002 ( .A1(n8050), .A2(n13090), .ZN(n7670) );
  NAND2_X1 U10003 ( .A1(n7669), .A2(n7670), .ZN(n7694) );
  INV_X1 U10004 ( .A(n7669), .ZN(n12976) );
  AND2_X1 U10005 ( .A1(n7694), .A2(n7671), .ZN(n10028) );
  MUX2_X1 U10006 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n6436), .Z(n7674) );
  NAND2_X1 U10007 ( .A1(n7674), .A2(SI_8_), .ZN(n7699) );
  OAI21_X1 U10008 ( .B1(SI_8_), .B2(n7674), .A(n7699), .ZN(n7675) );
  INV_X1 U10009 ( .A(n7675), .ZN(n7676) );
  NAND2_X1 U10010 ( .A1(n7700), .A2(n7678), .ZN(n10748) );
  INV_X1 U10011 ( .A(n7679), .ZN(n7680) );
  NAND2_X1 U10012 ( .A1(n7680), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7681) );
  MUX2_X1 U10013 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7681), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n7683) );
  INV_X1 U10014 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7682) );
  NAND2_X1 U10015 ( .A1(n7679), .A2(n7682), .ZN(n7727) );
  NAND2_X1 U10016 ( .A1(n7683), .A2(n7727), .ZN(n9667) );
  INV_X1 U10017 ( .A(n9667), .ZN(n9808) );
  AOI22_X1 U10018 ( .A1(n8510), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n9428), .B2(
        n9808), .ZN(n7684) );
  INV_X2 U10019 ( .A(n7686), .ZN(n8477) );
  NAND2_X1 U10020 ( .A1(n8477), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7693) );
  NAND2_X1 U10021 ( .A1(n8069), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7692) );
  NAND2_X1 U10022 ( .A1(n6704), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7691) );
  INV_X1 U10023 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7687) );
  NAND2_X1 U10024 ( .A1(n7688), .A2(n7687), .ZN(n7689) );
  NAND2_X1 U10025 ( .A1(n7710), .A2(n7689), .ZN(n12970) );
  OR2_X1 U10026 ( .A1(n8124), .A2(n12970), .ZN(n7690) );
  NAND4_X1 U10027 ( .A1(n7693), .A2(n7692), .A3(n7691), .A4(n7690), .ZN(n13089) );
  NAND2_X1 U10028 ( .A1(n8050), .A2(n13089), .ZN(n7697) );
  AND2_X1 U10029 ( .A1(n12978), .A2(n7694), .ZN(n7695) );
  INV_X1 U10030 ( .A(n7696), .ZN(n10203) );
  NAND2_X1 U10031 ( .A1(n10203), .A2(n7697), .ZN(n7698) );
  MUX2_X1 U10032 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n6436), .Z(n7701) );
  NAND2_X1 U10033 ( .A1(n7701), .A2(SI_9_), .ZN(n7721) );
  OAI21_X1 U10034 ( .B1(n7701), .B2(SI_9_), .A(n7721), .ZN(n7702) );
  INV_X1 U10035 ( .A(n7702), .ZN(n7703) );
  OR2_X1 U10036 ( .A1(n7704), .A2(n7703), .ZN(n7705) );
  NAND2_X1 U10037 ( .A1(n7722), .A2(n7705), .ZN(n10725) );
  OR2_X1 U10038 ( .A1(n10725), .A2(n7908), .ZN(n7708) );
  NAND2_X1 U10039 ( .A1(n7727), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7706) );
  XNOR2_X1 U10040 ( .A(n7706), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10120) );
  AOI22_X1 U10041 ( .A1(n7582), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n9428), .B2(
        n10120), .ZN(n7707) );
  NAND2_X2 U10042 ( .A1(n7708), .A2(n7707), .ZN(n10424) );
  XNOR2_X1 U10043 ( .A(n10424), .B(n8086), .ZN(n7717) );
  NAND2_X1 U10044 ( .A1(n8069), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7715) );
  NAND2_X1 U10045 ( .A1(n6704), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7714) );
  NAND2_X1 U10046 ( .A1(n8477), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7713) );
  INV_X1 U10047 ( .A(n7731), .ZN(n7733) );
  NAND2_X1 U10048 ( .A1(n7710), .A2(n7709), .ZN(n7711) );
  NAND2_X1 U10049 ( .A1(n7733), .A2(n7711), .ZN(n10404) );
  OR2_X1 U10050 ( .A1(n8124), .A2(n10404), .ZN(n7712) );
  NAND4_X1 U10051 ( .A1(n7715), .A2(n7714), .A3(n7713), .A4(n7712), .ZN(n13088) );
  NAND2_X1 U10052 ( .A1(n8050), .A2(n13088), .ZN(n7718) );
  XNOR2_X1 U10053 ( .A(n7717), .B(n7718), .ZN(n10202) );
  INV_X1 U10054 ( .A(n7717), .ZN(n7719) );
  NAND2_X1 U10055 ( .A1(n7719), .A2(n7718), .ZN(n7720) );
  INV_X1 U10056 ( .A(n7723), .ZN(n7724) );
  OR2_X1 U10057 ( .A1(n7725), .A2(n7724), .ZN(n7726) );
  NAND2_X1 U10058 ( .A1(n7742), .A2(n7726), .ZN(n10843) );
  NAND2_X1 U10059 ( .A1(n7743), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7728) );
  XNOR2_X1 U10060 ( .A(n7728), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10373) );
  AOI22_X1 U10061 ( .A1(n7582), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n9428), 
        .B2(n10373), .ZN(n7729) );
  NAND2_X2 U10062 ( .A1(n7730), .A2(n7729), .ZN(n12966) );
  NAND2_X1 U10063 ( .A1(n8477), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7738) );
  NAND2_X1 U10064 ( .A1(n8069), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7737) );
  NAND2_X1 U10065 ( .A1(n6704), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7736) );
  INV_X1 U10066 ( .A(n7748), .ZN(n7749) );
  INV_X1 U10067 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7732) );
  NAND2_X1 U10068 ( .A1(n7733), .A2(n7732), .ZN(n7734) );
  NAND2_X1 U10069 ( .A1(n7749), .A2(n7734), .ZN(n12956) );
  OR2_X1 U10070 ( .A1(n8124), .A2(n12956), .ZN(n7735) );
  NAND4_X1 U10071 ( .A1(n7738), .A2(n7737), .A3(n7736), .A4(n7735), .ZN(n13087) );
  AND2_X1 U10072 ( .A1(n8050), .A2(n13087), .ZN(n7739) );
  NAND2_X1 U10073 ( .A1(n12120), .A2(n7739), .ZN(n7755) );
  NAND2_X1 U10074 ( .A1(n7755), .A2(n7740), .ZN(n12962) );
  NAND2_X1 U10075 ( .A1(n10883), .A2(n8509), .ZN(n7747) );
  INV_X1 U10076 ( .A(n7765), .ZN(n7744) );
  NAND2_X1 U10077 ( .A1(n7744), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7745) );
  XNOR2_X1 U10078 ( .A(n7745), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10501) );
  AOI22_X1 U10079 ( .A1(n7582), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n9428), 
        .B2(n10501), .ZN(n7746) );
  NAND2_X1 U10080 ( .A1(n8069), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7754) );
  NAND2_X1 U10081 ( .A1(n6704), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7753) );
  NAND2_X1 U10082 ( .A1(n8477), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7752) );
  INV_X1 U10083 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10368) );
  NAND2_X1 U10084 ( .A1(n7749), .A2(n10368), .ZN(n7750) );
  NAND2_X1 U10085 ( .A1(n7776), .A2(n7750), .ZN(n12118) );
  OR2_X1 U10086 ( .A1(n8124), .A2(n12118), .ZN(n7751) );
  NAND4_X1 U10087 ( .A1(n7754), .A2(n7753), .A3(n7752), .A4(n7751), .ZN(n13086) );
  NAND2_X1 U10088 ( .A1(n8050), .A2(n13086), .ZN(n7756) );
  XNOR2_X1 U10089 ( .A(n12094), .B(n7756), .ZN(n12121) );
  INV_X1 U10090 ( .A(n12094), .ZN(n7757) );
  NAND2_X1 U10091 ( .A1(n7757), .A2(n7756), .ZN(n7758) );
  INV_X1 U10092 ( .A(n7759), .ZN(n7760) );
  NAND2_X1 U10093 ( .A1(n7760), .A2(n9384), .ZN(n7761) );
  MUX2_X1 U10094 ( .A(n8635), .B(n9594), .S(n6436), .Z(n7788) );
  XNOR2_X1 U10095 ( .A(n7787), .B(n7786), .ZN(n10999) );
  NAND2_X1 U10096 ( .A1(n10999), .A2(n8509), .ZN(n7774) );
  INV_X1 U10097 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n7764) );
  INV_X1 U10098 ( .A(n7769), .ZN(n7766) );
  NAND2_X1 U10099 ( .A1(n7766), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7767) );
  MUX2_X1 U10100 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7767), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n7770) );
  INV_X1 U10101 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7768) );
  NAND2_X1 U10102 ( .A1(n7769), .A2(n7768), .ZN(n7818) );
  NAND2_X1 U10103 ( .A1(n7770), .A2(n7818), .ZN(n11105) );
  OAI22_X1 U10104 ( .A1(n11105), .A2(n7771), .B1(n8487), .B2(n9594), .ZN(n7772) );
  INV_X1 U10105 ( .A(n7772), .ZN(n7773) );
  XNOR2_X1 U10106 ( .A(n12100), .B(n8086), .ZN(n7782) );
  NAND2_X1 U10107 ( .A1(n8069), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7781) );
  NAND2_X1 U10108 ( .A1(n8477), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7780) );
  INV_X1 U10109 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7775) );
  NAND2_X1 U10110 ( .A1(n7776), .A2(n7775), .ZN(n7777) );
  NAND2_X1 U10111 ( .A1(n7802), .A2(n7777), .ZN(n12093) );
  OR2_X1 U10112 ( .A1(n7572), .A2(n12093), .ZN(n7779) );
  INV_X1 U10113 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10678) );
  OR2_X1 U10114 ( .A1(n8480), .A2(n10678), .ZN(n7778) );
  NAND4_X1 U10115 ( .A1(n7781), .A2(n7780), .A3(n7779), .A4(n7778), .ZN(n13085) );
  NAND2_X1 U10116 ( .A1(n8050), .A2(n13085), .ZN(n7783) );
  XNOR2_X1 U10117 ( .A(n7782), .B(n7783), .ZN(n12095) );
  INV_X1 U10118 ( .A(n7782), .ZN(n7784) );
  NAND2_X1 U10119 ( .A1(n7784), .A2(n7783), .ZN(n7785) );
  NAND2_X1 U10120 ( .A1(n7788), .A2(n14350), .ZN(n7789) );
  MUX2_X1 U10121 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n6436), .Z(n7791) );
  INV_X1 U10122 ( .A(n7791), .ZN(n7792) );
  NAND2_X1 U10123 ( .A1(n7792), .A2(n9412), .ZN(n7793) );
  NAND2_X1 U10124 ( .A1(n7816), .A2(n7793), .ZN(n7796) );
  NAND2_X1 U10125 ( .A1(n7797), .A2(n7796), .ZN(n7798) );
  NAND2_X1 U10126 ( .A1(n7817), .A2(n7798), .ZN(n11025) );
  OR2_X1 U10127 ( .A1(n11025), .A2(n7908), .ZN(n7801) );
  NAND2_X1 U10128 ( .A1(n7818), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7799) );
  XNOR2_X1 U10129 ( .A(n7799), .B(P2_IR_REG_13__SCAN_IN), .ZN(n14861) );
  AOI22_X1 U10130 ( .A1(n14861), .A2(n9428), .B1(n7582), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n7800) );
  XNOR2_X1 U10131 ( .A(n11146), .B(n8086), .ZN(n7809) );
  INV_X1 U10132 ( .A(n7822), .ZN(n7824) );
  NAND2_X1 U10133 ( .A1(n7802), .A2(n14854), .ZN(n7803) );
  NAND2_X1 U10134 ( .A1(n7824), .A2(n7803), .ZN(n13033) );
  NAND2_X1 U10135 ( .A1(n8069), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7804) );
  OAI21_X1 U10136 ( .B1(n13033), .B2(n7572), .A(n7804), .ZN(n7808) );
  INV_X1 U10137 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7806) );
  NAND2_X1 U10138 ( .A1(n6704), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7805) );
  OAI21_X1 U10139 ( .B1(n7686), .B2(n7806), .A(n7805), .ZN(n7807) );
  AND2_X1 U10140 ( .A1(n8050), .A2(n13084), .ZN(n7810) );
  NAND2_X1 U10141 ( .A1(n7809), .A2(n7810), .ZN(n7815) );
  INV_X1 U10142 ( .A(n7809), .ZN(n7812) );
  INV_X1 U10143 ( .A(n7810), .ZN(n7811) );
  NAND2_X1 U10144 ( .A1(n7812), .A2(n7811), .ZN(n7813) );
  NAND2_X1 U10145 ( .A1(n7815), .A2(n7813), .ZN(n13029) );
  MUX2_X1 U10146 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n6450), .Z(n7832) );
  XNOR2_X1 U10147 ( .A(n7836), .B(n7835), .ZN(n11281) );
  NAND2_X1 U10148 ( .A1(n11281), .A2(n8509), .ZN(n7821) );
  NAND2_X1 U10149 ( .A1(n7837), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7819) );
  XNOR2_X1 U10150 ( .A(n7819), .B(P2_IR_REG_14__SCAN_IN), .ZN(n13148) );
  AOI22_X1 U10151 ( .A1(n13148), .A2(n9428), .B1(n7582), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n7820) );
  XNOR2_X1 U10152 ( .A(n14508), .B(n8130), .ZN(n7830) );
  INV_X1 U10153 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7828) );
  INV_X1 U10154 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7823) );
  NAND2_X1 U10155 ( .A1(n7824), .A2(n7823), .ZN(n7825) );
  NAND2_X1 U10156 ( .A1(n7842), .A2(n7825), .ZN(n14511) );
  OR2_X1 U10157 ( .A1(n14511), .A2(n8124), .ZN(n7827) );
  AOI22_X1 U10158 ( .A1(n6704), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8069), .B2(
        P2_REG1_REG_14__SCAN_IN), .ZN(n7826) );
  OAI211_X1 U10159 ( .C1(n7686), .C2(n7828), .A(n7827), .B(n7826), .ZN(n13083)
         );
  NAND2_X1 U10160 ( .A1(n13083), .A2(n8050), .ZN(n7829) );
  XNOR2_X1 U10161 ( .A(n7830), .B(n7829), .ZN(n14500) );
  NAND2_X1 U10162 ( .A1(n7830), .A2(n7829), .ZN(n7831) );
  INV_X1 U10163 ( .A(n7832), .ZN(n7833) );
  NAND2_X1 U10164 ( .A1(n7833), .A2(n14351), .ZN(n7834) );
  MUX2_X1 U10165 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n6436), .Z(n7854) );
  XNOR2_X1 U10166 ( .A(n7853), .B(n7852), .ZN(n11285) );
  NAND2_X1 U10167 ( .A1(n11285), .A2(n8509), .ZN(n7840) );
  OAI21_X1 U10168 ( .B1(n7837), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7838) );
  XNOR2_X1 U10169 ( .A(n7838), .B(P2_IR_REG_15__SCAN_IN), .ZN(n13168) );
  AOI22_X1 U10170 ( .A1(n13168), .A2(n9428), .B1(n7582), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n7839) );
  XNOR2_X1 U10171 ( .A(n11273), .B(n8086), .ZN(n7846) );
  INV_X1 U10172 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n11271) );
  INV_X1 U10173 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n13150) );
  NAND2_X1 U10174 ( .A1(n7842), .A2(n13150), .ZN(n7843) );
  NAND2_X1 U10175 ( .A1(n7886), .A2(n7843), .ZN(n11270) );
  OR2_X1 U10176 ( .A1(n11270), .A2(n8124), .ZN(n7845) );
  AOI22_X1 U10177 ( .A1(n8477), .A2(P2_REG0_REG_15__SCAN_IN), .B1(n8069), .B2(
        P2_REG1_REG_15__SCAN_IN), .ZN(n7844) );
  OAI211_X1 U10178 ( .C1(n8480), .C2(n11271), .A(n7845), .B(n7844), .ZN(n13082) );
  AND2_X1 U10179 ( .A1(n13082), .A2(n8050), .ZN(n7847) );
  NAND2_X1 U10180 ( .A1(n7846), .A2(n7847), .ZN(n7851) );
  INV_X1 U10181 ( .A(n7846), .ZN(n7849) );
  INV_X1 U10182 ( .A(n7847), .ZN(n7848) );
  NAND2_X1 U10183 ( .A1(n7849), .A2(n7848), .ZN(n7850) );
  NAND2_X1 U10184 ( .A1(n7851), .A2(n7850), .ZN(n9234) );
  INV_X1 U10185 ( .A(n7854), .ZN(n7855) );
  MUX2_X1 U10186 ( .A(n10215), .B(n10217), .S(n6450), .Z(n7875) );
  XNOR2_X1 U10187 ( .A(n7874), .B(n7873), .ZN(n11342) );
  NAND2_X1 U10188 ( .A1(n11342), .A2(n8509), .ZN(n7864) );
  INV_X1 U10189 ( .A(n7856), .ZN(n7857) );
  NOR2_X1 U10190 ( .A1(n7858), .A2(n7857), .ZN(n7859) );
  NAND2_X1 U10191 ( .A1(n7679), .A2(n7859), .ZN(n7861) );
  NAND2_X1 U10192 ( .A1(n7861), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7860) );
  MUX2_X1 U10193 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7860), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n7862) );
  OR2_X1 U10194 ( .A1(n7861), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n7877) );
  AND2_X1 U10195 ( .A1(n7862), .A2(n7877), .ZN(n13172) );
  AOI22_X1 U10196 ( .A1(n8510), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n9428), 
        .B2(n13172), .ZN(n7863) );
  XNOR2_X1 U10197 ( .A(n13504), .B(n8086), .ZN(n13005) );
  INV_X1 U10198 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7884) );
  XNOR2_X1 U10199 ( .A(n7886), .B(n7884), .ZN(n14527) );
  OR2_X1 U10200 ( .A1(n14527), .A2(n8124), .ZN(n7869) );
  INV_X1 U10201 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13188) );
  NAND2_X1 U10202 ( .A1(n8069), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7866) );
  NAND2_X1 U10203 ( .A1(n8477), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7865) );
  OAI211_X1 U10204 ( .C1(n8480), .C2(n13188), .A(n7866), .B(n7865), .ZN(n7867)
         );
  INV_X1 U10205 ( .A(n7867), .ZN(n7868) );
  NAND2_X1 U10206 ( .A1(n7869), .A2(n7868), .ZN(n13081) );
  NAND2_X1 U10207 ( .A1(n13081), .A2(n8050), .ZN(n7870) );
  XNOR2_X1 U10208 ( .A(n13005), .B(n7870), .ZN(n14513) );
  INV_X1 U10209 ( .A(n13005), .ZN(n7871) );
  NAND2_X1 U10210 ( .A1(n7871), .A2(n7870), .ZN(n7872) );
  NAND2_X1 U10211 ( .A1(n7875), .A2(n9647), .ZN(n7876) );
  MUX2_X1 U10212 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n6450), .Z(n7900) );
  XNOR2_X1 U10213 ( .A(n7899), .B(n7898), .ZN(n11601) );
  NAND2_X1 U10214 ( .A1(n11601), .A2(n8509), .ZN(n7882) );
  NAND2_X1 U10215 ( .A1(n7877), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7878) );
  MUX2_X1 U10216 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7878), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n7880) );
  NAND2_X1 U10217 ( .A1(n7880), .A2(n7879), .ZN(n13198) );
  INV_X1 U10218 ( .A(n13198), .ZN(n13203) );
  AOI22_X1 U10219 ( .A1(n8510), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n9428), 
        .B2(n13203), .ZN(n7881) );
  XNOR2_X1 U10220 ( .A(n13498), .B(n8086), .ZN(n7894) );
  INV_X1 U10221 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7883) );
  OAI21_X1 U10222 ( .B1(n7886), .B2(n7884), .A(n7883), .ZN(n7887) );
  NAND2_X1 U10223 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_REG3_REG_17__SCAN_IN), 
        .ZN(n7885) );
  AND2_X1 U10224 ( .A1(n7887), .A2(n7913), .ZN(n13001) );
  NAND2_X1 U10225 ( .A1(n13001), .A2(n8186), .ZN(n7892) );
  INV_X1 U10226 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n14345) );
  NAND2_X1 U10227 ( .A1(n8477), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n7889) );
  NAND2_X1 U10228 ( .A1(n8069), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7888) );
  OAI211_X1 U10229 ( .C1(n14345), .C2(n8480), .A(n7889), .B(n7888), .ZN(n7890)
         );
  INV_X1 U10230 ( .A(n7890), .ZN(n7891) );
  NAND2_X1 U10231 ( .A1(n7892), .A2(n7891), .ZN(n13080) );
  NAND2_X1 U10232 ( .A1(n13080), .A2(n8050), .ZN(n7895) );
  XNOR2_X1 U10233 ( .A(n7894), .B(n7895), .ZN(n13006) );
  INV_X1 U10234 ( .A(n7894), .ZN(n7896) );
  NAND2_X1 U10235 ( .A1(n7896), .A2(n7895), .ZN(n7897) );
  NAND2_X1 U10236 ( .A1(n7899), .A2(n7898), .ZN(n7903) );
  INV_X1 U10237 ( .A(n7900), .ZN(n7901) );
  NAND2_X1 U10238 ( .A1(n7901), .A2(n9757), .ZN(n7902) );
  NAND2_X1 U10239 ( .A1(n7903), .A2(n7902), .ZN(n7904) );
  INV_X1 U10240 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10511) );
  MUX2_X1 U10241 ( .A(n10513), .B(n10511), .S(n6436), .Z(n7905) );
  NAND2_X1 U10242 ( .A1(n7906), .A2(n7905), .ZN(n7907) );
  NAND2_X1 U10243 ( .A1(n7926), .A2(n7907), .ZN(n11611) );
  OR2_X1 U10244 ( .A1(n11611), .A2(n7908), .ZN(n7911) );
  NAND2_X1 U10245 ( .A1(n7879), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7909) );
  XNOR2_X1 U10246 ( .A(n7909), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13211) );
  AOI22_X1 U10247 ( .A1(n8510), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n9428), 
        .B2(n13211), .ZN(n7910) );
  XNOR2_X1 U10248 ( .A(n13493), .B(n8086), .ZN(n12108) );
  INV_X1 U10249 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n14308) );
  NAND2_X1 U10250 ( .A1(n7913), .A2(n14308), .ZN(n7914) );
  NAND2_X1 U10251 ( .A1(n7931), .A2(n7914), .ZN(n13411) );
  OR2_X1 U10252 ( .A1(n13411), .A2(n8124), .ZN(n7920) );
  INV_X1 U10253 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n7917) );
  NAND2_X1 U10254 ( .A1(n8477), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7916) );
  NAND2_X1 U10255 ( .A1(n8069), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n7915) );
  OAI211_X1 U10256 ( .C1(n7917), .C2(n8480), .A(n7916), .B(n7915), .ZN(n7918)
         );
  INV_X1 U10257 ( .A(n7918), .ZN(n7919) );
  NAND2_X1 U10258 ( .A1(n7920), .A2(n7919), .ZN(n13079) );
  AND2_X1 U10259 ( .A1(n13079), .A2(n8050), .ZN(n7921) );
  NAND2_X1 U10260 ( .A1(n12108), .A2(n7921), .ZN(n7939) );
  INV_X1 U10261 ( .A(n12108), .ZN(n7923) );
  INV_X1 U10262 ( .A(n7921), .ZN(n7922) );
  NAND2_X1 U10263 ( .A1(n7923), .A2(n7922), .ZN(n7924) );
  NAND2_X1 U10264 ( .A1(n7939), .A2(n7924), .ZN(n13058) );
  NAND2_X1 U10265 ( .A1(n7966), .A2(SI_19_), .ZN(n7945) );
  OR2_X1 U10266 ( .A1(n7966), .A2(SI_19_), .ZN(n7927) );
  MUX2_X1 U10267 ( .A(n10942), .B(n10944), .S(n6450), .Z(n7964) );
  NAND2_X1 U10268 ( .A1(n11625), .A2(n8509), .ZN(n7929) );
  AOI22_X1 U10269 ( .A1(n8510), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9428), 
        .B2(n9998), .ZN(n7928) );
  NAND2_X2 U10270 ( .A1(n7929), .A2(n7928), .ZN(n13488) );
  XNOR2_X1 U10271 ( .A(n13488), .B(n8086), .ZN(n7941) );
  INV_X1 U10272 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7930) );
  NAND2_X1 U10273 ( .A1(n7931), .A2(n7930), .ZN(n7932) );
  AND2_X1 U10274 ( .A1(n7952), .A2(n7932), .ZN(n13397) );
  NAND2_X1 U10275 ( .A1(n13397), .A2(n8186), .ZN(n7938) );
  INV_X1 U10276 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n7935) );
  NAND2_X1 U10277 ( .A1(n8069), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n7934) );
  NAND2_X1 U10278 ( .A1(n8477), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n7933) );
  OAI211_X1 U10279 ( .C1(n8480), .C2(n7935), .A(n7934), .B(n7933), .ZN(n7936)
         );
  INV_X1 U10280 ( .A(n7936), .ZN(n7937) );
  NAND2_X1 U10281 ( .A1(n7938), .A2(n7937), .ZN(n13371) );
  NAND2_X1 U10282 ( .A1(n13371), .A2(n8050), .ZN(n7942) );
  XNOR2_X1 U10283 ( .A(n7941), .B(n7942), .ZN(n12109) );
  INV_X1 U10284 ( .A(n7941), .ZN(n7943) );
  NAND2_X1 U10285 ( .A1(n7943), .A2(n7942), .ZN(n7944) );
  NAND2_X1 U10286 ( .A1(n7946), .A2(n7945), .ZN(n7948) );
  MUX2_X1 U10287 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n6436), .Z(n7967) );
  XNOR2_X1 U10288 ( .A(n7967), .B(SI_20_), .ZN(n7947) );
  NAND2_X1 U10289 ( .A1(n11647), .A2(n8509), .ZN(n7950) );
  NAND2_X1 U10290 ( .A1(n8510), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7949) );
  XNOR2_X1 U10291 ( .A(n13481), .B(n8130), .ZN(n7959) );
  INV_X1 U10292 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13024) );
  NAND2_X1 U10293 ( .A1(n7952), .A2(n13024), .ZN(n7953) );
  NAND2_X1 U10294 ( .A1(n7971), .A2(n7953), .ZN(n13378) );
  OR2_X1 U10295 ( .A1(n13378), .A2(n7572), .ZN(n7958) );
  INV_X1 U10296 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n13379) );
  NAND2_X1 U10297 ( .A1(n8477), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n7955) );
  NAND2_X1 U10298 ( .A1(n8069), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n7954) );
  OAI211_X1 U10299 ( .C1(n13379), .C2(n8480), .A(n7955), .B(n7954), .ZN(n7956)
         );
  INV_X1 U10300 ( .A(n7956), .ZN(n7957) );
  NAND2_X1 U10301 ( .A1(n7958), .A2(n7957), .ZN(n13358) );
  NAND2_X1 U10302 ( .A1(n13358), .A2(n8050), .ZN(n7960) );
  NAND2_X1 U10303 ( .A1(n7959), .A2(n7960), .ZN(n13021) );
  INV_X1 U10304 ( .A(n7959), .ZN(n7962) );
  INV_X1 U10305 ( .A(n7960), .ZN(n7961) );
  NAND2_X1 U10306 ( .A1(n7962), .A2(n7961), .ZN(n13020) );
  INV_X1 U10307 ( .A(n7967), .ZN(n7963) );
  INV_X1 U10308 ( .A(SI_20_), .ZN(n10197) );
  AOI22_X1 U10309 ( .A1(n10012), .A2(n7964), .B1(n7963), .B2(n10197), .ZN(
        n7965) );
  NAND2_X1 U10310 ( .A1(n7967), .A2(SI_20_), .ZN(n7968) );
  MUX2_X1 U10311 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n6450), .Z(n8026) );
  XNOR2_X1 U10312 ( .A(n7984), .B(n8026), .ZN(n11659) );
  NAND2_X1 U10313 ( .A1(n11659), .A2(n8509), .ZN(n7970) );
  NAND2_X1 U10314 ( .A1(n8510), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7969) );
  XNOR2_X1 U10315 ( .A(n13477), .B(n8086), .ZN(n7980) );
  INV_X1 U10316 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12986) );
  NAND2_X1 U10317 ( .A1(n7971), .A2(n12986), .ZN(n7972) );
  AND2_X1 U10318 ( .A1(n7990), .A2(n7972), .ZN(n12988) );
  NAND2_X1 U10319 ( .A1(n12988), .A2(n8186), .ZN(n7977) );
  INV_X1 U10320 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n13361) );
  NAND2_X1 U10321 ( .A1(n8069), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n7974) );
  NAND2_X1 U10322 ( .A1(n8477), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n7973) );
  OAI211_X1 U10323 ( .C1(n13361), .C2(n8480), .A(n7974), .B(n7973), .ZN(n7975)
         );
  INV_X1 U10324 ( .A(n7975), .ZN(n7976) );
  NAND2_X1 U10325 ( .A1(n7977), .A2(n7976), .ZN(n13373) );
  NAND2_X1 U10326 ( .A1(n13373), .A2(n8050), .ZN(n7978) );
  XNOR2_X1 U10327 ( .A(n7980), .B(n7978), .ZN(n12984) );
  INV_X1 U10328 ( .A(n7978), .ZN(n7979) );
  NAND2_X1 U10329 ( .A1(n7980), .A2(n7979), .ZN(n7981) );
  INV_X1 U10330 ( .A(n8026), .ZN(n7983) );
  NAND2_X1 U10331 ( .A1(n8025), .A2(SI_21_), .ZN(n7985) );
  MUX2_X1 U10332 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n6436), .Z(n8021) );
  XNOR2_X1 U10333 ( .A(n11678), .B(n8021), .ZN(n11263) );
  NAND2_X1 U10334 ( .A1(n11263), .A2(n8509), .ZN(n7987) );
  NAND2_X1 U10335 ( .A1(n8510), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n7986) );
  NAND2_X2 U10336 ( .A1(n7987), .A2(n7986), .ZN(n13472) );
  XNOR2_X1 U10337 ( .A(n13472), .B(n8130), .ZN(n7998) );
  INV_X1 U10338 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n7989) );
  NAND2_X1 U10339 ( .A1(n7990), .A2(n7989), .ZN(n7991) );
  NAND2_X1 U10340 ( .A1(n8043), .A2(n7991), .ZN(n13342) );
  OR2_X1 U10341 ( .A1(n13342), .A2(n7572), .ZN(n7997) );
  INV_X1 U10342 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n7994) );
  NAND2_X1 U10343 ( .A1(n8477), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n7993) );
  NAND2_X1 U10344 ( .A1(n8069), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n7992) );
  OAI211_X1 U10345 ( .C1(n7994), .C2(n8480), .A(n7993), .B(n7992), .ZN(n7995)
         );
  INV_X1 U10346 ( .A(n7995), .ZN(n7996) );
  NAND2_X1 U10347 ( .A1(n7997), .A2(n7996), .ZN(n13357) );
  AND2_X1 U10348 ( .A1(n13357), .A2(n8050), .ZN(n13041) );
  NAND2_X1 U10349 ( .A1(n13042), .A2(n13041), .ZN(n8002) );
  INV_X1 U10350 ( .A(n7998), .ZN(n7999) );
  NAND2_X1 U10351 ( .A1(n8000), .A2(n7999), .ZN(n8001) );
  INV_X1 U10352 ( .A(n11678), .ZN(n8003) );
  NAND2_X1 U10353 ( .A1(n8003), .A2(n8021), .ZN(n8006) );
  NAND2_X1 U10354 ( .A1(n8004), .A2(SI_22_), .ZN(n8005) );
  MUX2_X1 U10355 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n6436), .Z(n8030) );
  XNOR2_X1 U10356 ( .A(n8030), .B(SI_23_), .ZN(n8007) );
  NAND2_X1 U10357 ( .A1(n11697), .A2(n8509), .ZN(n8010) );
  NAND2_X1 U10358 ( .A1(n8510), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8009) );
  XNOR2_X1 U10359 ( .A(n13465), .B(n8130), .ZN(n8016) );
  XNOR2_X1 U10360 ( .A(n8043), .B(P2_REG3_REG_23__SCAN_IN), .ZN(n13321) );
  NAND2_X1 U10361 ( .A1(n13321), .A2(n8186), .ZN(n8015) );
  INV_X1 U10362 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13322) );
  NAND2_X1 U10363 ( .A1(n8477), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8012) );
  NAND2_X1 U10364 ( .A1(n8069), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8011) );
  OAI211_X1 U10365 ( .C1(n13322), .C2(n8480), .A(n8012), .B(n8011), .ZN(n8013)
         );
  INV_X1 U10366 ( .A(n8013), .ZN(n8014) );
  NAND2_X1 U10367 ( .A1(n8015), .A2(n8014), .ZN(n13338) );
  AND2_X1 U10368 ( .A1(n13338), .A2(n8050), .ZN(n12948) );
  INV_X1 U10369 ( .A(n8016), .ZN(n8017) );
  NAND2_X1 U10370 ( .A1(n8018), .A2(n8017), .ZN(n8019) );
  INV_X1 U10371 ( .A(n8030), .ZN(n8020) );
  INV_X1 U10372 ( .A(SI_23_), .ZN(n10631) );
  NAND2_X1 U10373 ( .A1(n8020), .A2(n10631), .ZN(n8029) );
  INV_X1 U10374 ( .A(SI_22_), .ZN(n9029) );
  NAND2_X1 U10375 ( .A1(n8027), .A2(n9029), .ZN(n8022) );
  NAND2_X1 U10376 ( .A1(n8029), .A2(n8022), .ZN(n8034) );
  NOR2_X1 U10377 ( .A1(n8026), .A2(SI_21_), .ZN(n8023) );
  NOR2_X1 U10378 ( .A1(n8034), .A2(n8023), .ZN(n8024) );
  NAND2_X1 U10379 ( .A1(n8026), .A2(SI_21_), .ZN(n8033) );
  NOR2_X1 U10380 ( .A1(n8027), .A2(n9029), .ZN(n8028) );
  NAND2_X1 U10381 ( .A1(n8029), .A2(n8028), .ZN(n8032) );
  NAND2_X1 U10382 ( .A1(n8030), .A2(SI_23_), .ZN(n8031) );
  OAI211_X1 U10383 ( .C1(n8034), .C2(n8033), .A(n8032), .B(n8031), .ZN(n8035)
         );
  INV_X1 U10384 ( .A(n8035), .ZN(n8036) );
  MUX2_X1 U10385 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n6450), .Z(n8058) );
  XNOR2_X1 U10386 ( .A(n8058), .B(SI_24_), .ZN(n8038) );
  XNOR2_X1 U10387 ( .A(n8057), .B(n8038), .ZN(n11715) );
  NAND2_X1 U10388 ( .A1(n11715), .A2(n8509), .ZN(n8040) );
  NAND2_X1 U10389 ( .A1(n8510), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8039) );
  XNOR2_X1 U10390 ( .A(n13462), .B(n8086), .ZN(n8053) );
  INV_X1 U10391 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n12952) );
  INV_X1 U10392 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8041) );
  OAI21_X1 U10393 ( .B1(n8043), .B2(n12952), .A(n8041), .ZN(n8044) );
  NAND2_X1 U10394 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(P2_REG3_REG_23__SCAN_IN), 
        .ZN(n8042) );
  NAND2_X1 U10395 ( .A1(n8044), .A2(n8067), .ZN(n13311) );
  OR2_X1 U10396 ( .A1(n13311), .A2(n8124), .ZN(n8049) );
  INV_X1 U10397 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13310) );
  NAND2_X1 U10398 ( .A1(n8477), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8046) );
  NAND2_X1 U10399 ( .A1(n8069), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8045) );
  OAI211_X1 U10400 ( .C1(n13310), .C2(n8480), .A(n8046), .B(n8045), .ZN(n8047)
         );
  INV_X1 U10401 ( .A(n8047), .ZN(n8048) );
  NAND2_X1 U10402 ( .A1(n8049), .A2(n8048), .ZN(n13078) );
  NAND2_X1 U10403 ( .A1(n13078), .A2(n8050), .ZN(n8051) );
  INV_X1 U10404 ( .A(n8051), .ZN(n8052) );
  NAND2_X1 U10405 ( .A1(n8053), .A2(n8052), .ZN(n8054) );
  INV_X1 U10406 ( .A(n8058), .ZN(n8055) );
  INV_X1 U10407 ( .A(SI_24_), .ZN(n10928) );
  NAND2_X1 U10408 ( .A1(n8055), .A2(n10928), .ZN(n8056) );
  NAND2_X1 U10409 ( .A1(n8058), .A2(SI_24_), .ZN(n8059) );
  INV_X1 U10410 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11738) );
  INV_X1 U10411 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11172) );
  MUX2_X1 U10412 ( .A(n11738), .B(n11172), .S(n6436), .Z(n8060) );
  INV_X1 U10413 ( .A(SI_25_), .ZN(n11830) );
  NAND2_X1 U10414 ( .A1(n8060), .A2(n11830), .ZN(n8083) );
  INV_X1 U10415 ( .A(n8060), .ZN(n8061) );
  NAND2_X1 U10416 ( .A1(n8061), .A2(SI_25_), .ZN(n8062) );
  NAND2_X1 U10417 ( .A1(n8083), .A2(n8062), .ZN(n8081) );
  XNOR2_X1 U10418 ( .A(n8082), .B(n8081), .ZN(n11737) );
  NAND2_X1 U10419 ( .A1(n11737), .A2(n8509), .ZN(n8064) );
  NAND2_X1 U10420 ( .A1(n8510), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8063) );
  XNOR2_X1 U10421 ( .A(n13456), .B(n8086), .ZN(n8078) );
  INV_X1 U10422 ( .A(n8067), .ZN(n8065) );
  NAND2_X1 U10423 ( .A1(n8065), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n8087) );
  INV_X1 U10424 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8066) );
  NAND2_X1 U10425 ( .A1(n8067), .A2(n8066), .ZN(n8068) );
  NAND2_X1 U10426 ( .A1(n8087), .A2(n8068), .ZN(n12996) );
  OR2_X1 U10427 ( .A1(n12996), .A2(n7572), .ZN(n8075) );
  INV_X1 U10428 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8072) );
  NAND2_X1 U10429 ( .A1(n8477), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8071) );
  NAND2_X1 U10430 ( .A1(n8069), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8070) );
  OAI211_X1 U10431 ( .C1(n8072), .C2(n8480), .A(n8071), .B(n8070), .ZN(n8073)
         );
  INV_X1 U10432 ( .A(n8073), .ZN(n8074) );
  NAND2_X1 U10433 ( .A1(n13077), .A2(n8050), .ZN(n8076) );
  XNOR2_X1 U10434 ( .A(n8078), .B(n8076), .ZN(n12994) );
  INV_X1 U10435 ( .A(n8076), .ZN(n8077) );
  NAND2_X1 U10436 ( .A1(n8078), .A2(n8077), .ZN(n8079) );
  INV_X1 U10437 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n11760) );
  INV_X1 U10438 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n11336) );
  MUX2_X1 U10439 ( .A(n11760), .B(n11336), .S(n6450), .Z(n8100) );
  NAND2_X1 U10440 ( .A1(n11759), .A2(n8509), .ZN(n8085) );
  NAND2_X1 U10441 ( .A1(n8510), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8084) );
  XNOR2_X1 U10442 ( .A(n13282), .B(n8086), .ZN(n8094) );
  INV_X1 U10443 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n13067) );
  NAND2_X1 U10444 ( .A1(n8087), .A2(n13067), .ZN(n8088) );
  NAND2_X1 U10445 ( .A1(n8110), .A2(n8088), .ZN(n13284) );
  OR2_X1 U10446 ( .A1(n13284), .A2(n8124), .ZN(n8093) );
  INV_X1 U10447 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n13283) );
  NAND2_X1 U10448 ( .A1(n8069), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8090) );
  NAND2_X1 U10449 ( .A1(n8477), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8089) );
  OAI211_X1 U10450 ( .C1(n13283), .C2(n8480), .A(n8090), .B(n8089), .ZN(n8091)
         );
  INV_X1 U10451 ( .A(n8091), .ZN(n8092) );
  NAND2_X1 U10452 ( .A1(n13076), .A2(n8050), .ZN(n8095) );
  NAND2_X1 U10453 ( .A1(n8094), .A2(n8095), .ZN(n8099) );
  INV_X1 U10454 ( .A(n8094), .ZN(n8097) );
  INV_X1 U10455 ( .A(n8095), .ZN(n8096) );
  NAND2_X1 U10456 ( .A1(n8097), .A2(n8096), .ZN(n8098) );
  NAND2_X1 U10457 ( .A1(n8099), .A2(n8098), .ZN(n13065) );
  INV_X1 U10458 ( .A(n8100), .ZN(n8101) );
  INV_X1 U10459 ( .A(SI_26_), .ZN(n11195) );
  INV_X1 U10460 ( .A(SI_27_), .ZN(n11332) );
  MUX2_X1 U10461 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n6436), .Z(n8168) );
  NAND2_X1 U10462 ( .A1(n13547), .A2(n8509), .ZN(n8108) );
  NAND2_X1 U10463 ( .A1(n8510), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8107) );
  XNOR2_X1 U10464 ( .A(n13444), .B(n8130), .ZN(n8119) );
  INV_X1 U10465 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8109) );
  NAND2_X1 U10466 ( .A1(n8110), .A2(n8109), .ZN(n8111) );
  NAND2_X1 U10467 ( .A1(n13266), .A2(n8186), .ZN(n8117) );
  INV_X1 U10468 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8114) );
  NAND2_X1 U10469 ( .A1(n8477), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8113) );
  NAND2_X1 U10470 ( .A1(n8069), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8112) );
  OAI211_X1 U10471 ( .C1(n8114), .C2(n8480), .A(n8113), .B(n8112), .ZN(n8115)
         );
  INV_X1 U10472 ( .A(n8115), .ZN(n8116) );
  NAND2_X1 U10473 ( .A1(n13075), .A2(n8050), .ZN(n8118) );
  XNOR2_X1 U10474 ( .A(n8119), .B(n8118), .ZN(n12943) );
  INV_X1 U10475 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8120) );
  INV_X1 U10476 ( .A(n11565), .ZN(n8123) );
  NAND2_X1 U10477 ( .A1(n8121), .A2(n8120), .ZN(n8122) );
  NAND2_X1 U10478 ( .A1(n8123), .A2(n8122), .ZN(n13252) );
  INV_X1 U10479 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13251) );
  NAND2_X1 U10480 ( .A1(n8477), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8126) );
  NAND2_X1 U10481 ( .A1(n8069), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8125) );
  OAI211_X1 U10482 ( .C1(n13251), .C2(n8480), .A(n8126), .B(n8125), .ZN(n8127)
         );
  INV_X1 U10483 ( .A(n8127), .ZN(n8128) );
  NAND2_X1 U10484 ( .A1(n13074), .A2(n8050), .ZN(n8131) );
  XNOR2_X1 U10485 ( .A(n8131), .B(n8130), .ZN(n8132) );
  INV_X1 U10486 ( .A(n8184), .ZN(n8167) );
  NOR4_X1 U10487 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n8136) );
  NOR4_X1 U10488 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n8135) );
  NOR4_X1 U10489 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8134) );
  NOR4_X1 U10490 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n8133) );
  NAND4_X1 U10491 ( .A1(n8136), .A2(n8135), .A3(n8134), .A4(n8133), .ZN(n8156)
         );
  NOR2_X1 U10492 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .ZN(
        n8140) );
  NOR4_X1 U10493 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n8139) );
  NOR4_X1 U10494 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n8138) );
  NOR4_X1 U10495 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n8137) );
  NAND4_X1 U10496 ( .A1(n8140), .A2(n8139), .A3(n8138), .A4(n8137), .ZN(n8155)
         );
  NAND2_X1 U10497 ( .A1(n8148), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8143) );
  MUX2_X1 U10498 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8143), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8145) );
  NAND2_X1 U10499 ( .A1(n8146), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8147) );
  MUX2_X1 U10500 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8147), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8149) );
  NAND2_X1 U10501 ( .A1(n8149), .A2(n8148), .ZN(n11170) );
  INV_X1 U10502 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8150) );
  INV_X1 U10503 ( .A(P2_B_REG_SCAN_IN), .ZN(n8152) );
  XOR2_X1 U10504 ( .A(n11087), .B(n8152), .Z(n8153) );
  OAI21_X1 U10505 ( .B1(n8156), .B2(n8155), .A(n14873), .ZN(n8194) );
  NAND2_X1 U10506 ( .A1(n8157), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8159) );
  XNOR2_X1 U10507 ( .A(n8159), .B(n8158), .ZN(n9430) );
  INV_X1 U10508 ( .A(n14872), .ZN(n8160) );
  AND2_X1 U10509 ( .A1(n8194), .A2(n8160), .ZN(n9456) );
  NAND2_X1 U10510 ( .A1(n11087), .A2(n11338), .ZN(n14906) );
  INV_X1 U10511 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n8161) );
  NAND2_X1 U10512 ( .A1(n14873), .A2(n8161), .ZN(n8162) );
  NAND2_X1 U10513 ( .A1(n9456), .A2(n9994), .ZN(n8164) );
  INV_X1 U10514 ( .A(n14873), .ZN(n8163) );
  NAND2_X1 U10515 ( .A1(n11338), .A2(n11170), .ZN(n14908) );
  NOR2_X1 U10516 ( .A1(n8164), .A2(n9995), .ZN(n8181) );
  INV_X1 U10517 ( .A(n9431), .ZN(n8165) );
  NAND2_X1 U10518 ( .A1(n13226), .A2(n11102), .ZN(n8577) );
  NAND2_X1 U10519 ( .A1(n7166), .A2(n8577), .ZN(n14922) );
  AND2_X1 U10520 ( .A1(n8165), .A2(n14922), .ZN(n8166) );
  NAND2_X1 U10521 ( .A1(n8167), .A2(n14523), .ZN(n8203) );
  NAND2_X1 U10522 ( .A1(n8169), .A2(n8168), .ZN(n8172) );
  NAND2_X1 U10523 ( .A1(n8170), .A2(SI_27_), .ZN(n8171) );
  INV_X1 U10524 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14257) );
  INV_X1 U10525 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n11503) );
  MUX2_X1 U10526 ( .A(n14257), .B(n11503), .S(n6450), .Z(n8173) );
  INV_X1 U10527 ( .A(SI_28_), .ZN(n12940) );
  NAND2_X1 U10528 ( .A1(n8173), .A2(n12940), .ZN(n8465) );
  INV_X1 U10529 ( .A(n8173), .ZN(n8174) );
  NAND2_X1 U10530 ( .A1(n8174), .A2(SI_28_), .ZN(n8175) );
  NAND2_X1 U10531 ( .A1(n8465), .A2(n8175), .ZN(n8176) );
  NAND2_X1 U10532 ( .A1(n8177), .A2(n8176), .ZN(n8178) );
  NAND2_X1 U10533 ( .A1(n8466), .A2(n8178), .ZN(n11793) );
  NAND2_X1 U10534 ( .A1(n11793), .A2(n8509), .ZN(n8180) );
  NAND2_X1 U10535 ( .A1(n8510), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8179) );
  INV_X1 U10536 ( .A(n8181), .ZN(n8193) );
  NAND2_X1 U10537 ( .A1(n7166), .A2(n9462), .ZN(n10001) );
  OR2_X1 U10538 ( .A1(n8193), .A2(n10001), .ZN(n8183) );
  NOR2_X1 U10539 ( .A1(n9462), .A2(n13226), .ZN(n8182) );
  NAND2_X1 U10540 ( .A1(n14927), .A2(n11099), .ZN(n9457) );
  NAND2_X1 U10541 ( .A1(n13438), .A2(n8185), .ZN(n8202) );
  NAND2_X1 U10542 ( .A1(n11565), .A2(n8186), .ZN(n8191) );
  INV_X1 U10543 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n11567) );
  NAND2_X1 U10544 ( .A1(n8477), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8188) );
  NAND2_X1 U10545 ( .A1(n8069), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8187) );
  OAI211_X1 U10546 ( .C1(n11567), .C2(n8480), .A(n8188), .B(n8187), .ZN(n8189)
         );
  INV_X1 U10547 ( .A(n8189), .ZN(n8190) );
  NAND2_X1 U10548 ( .A1(n8191), .A2(n8190), .ZN(n13073) );
  INV_X1 U10549 ( .A(n8192), .ZN(n9439) );
  NAND2_X1 U10550 ( .A1(n9431), .A2(n9439), .ZN(n13051) );
  AOI22_X1 U10551 ( .A1(n13073), .A2(n13372), .B1(n13075), .B2(n13370), .ZN(
        n13245) );
  INV_X1 U10552 ( .A(n13252), .ZN(n8198) );
  NAND2_X1 U10553 ( .A1(n8194), .A2(n9994), .ZN(n8195) );
  OAI21_X1 U10554 ( .B1(n9995), .B2(n8195), .A(n9457), .ZN(n8197) );
  NAND2_X1 U10555 ( .A1(n9431), .A2(n8577), .ZN(n9455) );
  AND3_X1 U10556 ( .A1(n9432), .A2(n9430), .A3(n9455), .ZN(n8196) );
  NAND2_X1 U10557 ( .A1(n8197), .A2(n8196), .ZN(n9733) );
  INV_X1 U10558 ( .A(n14528), .ZN(n13036) );
  AOI22_X1 U10559 ( .A1(n8198), .A2(n13036), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n8199) );
  OAI21_X1 U10560 ( .B1(n13245), .B2(n13066), .A(n8199), .ZN(n8200) );
  OAI211_X1 U10561 ( .C1(n8203), .C2(n13438), .A(n8202), .B(n8201), .ZN(
        P2_U3192) );
  XNOR2_X1 U10562 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n8299) );
  INV_X1 U10563 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n14652) );
  AND2_X1 U10564 ( .A1(n14652), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n8232) );
  INV_X1 U10565 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14410) );
  INV_X1 U10566 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14627) );
  XNOR2_X1 U10567 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n8243) );
  INV_X1 U10568 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14613) );
  INV_X1 U10569 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14311) );
  INV_X1 U10570 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n8225) );
  XNOR2_X1 U10571 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n8248) );
  INV_X1 U10572 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n8220) );
  INV_X1 U10573 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n8218) );
  XNOR2_X1 U10574 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n8278) );
  NAND2_X1 U10575 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(n8261), .ZN(n8260) );
  XNOR2_X1 U10576 ( .A(n8205), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n8257) );
  NOR2_X1 U10577 ( .A1(n8206), .A2(n7123), .ZN(n8208) );
  INV_X1 U10578 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n14264) );
  NOR2_X1 U10579 ( .A1(n8210), .A2(n14264), .ZN(n8212) );
  INV_X1 U10580 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9480) );
  NAND2_X1 U10581 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n9480), .ZN(n8213) );
  NAND2_X1 U10582 ( .A1(n8214), .A2(P3_ADDR_REG_7__SCAN_IN), .ZN(n8216) );
  XNOR2_X1 U10583 ( .A(n8214), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n8277) );
  NAND2_X1 U10584 ( .A1(n8278), .A2(n8279), .ZN(n8217) );
  XOR2_X1 U10585 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), .Z(
        n8251) );
  INV_X1 U10586 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14601) );
  NAND2_X1 U10587 ( .A1(n8221), .A2(n14601), .ZN(n8223) );
  XNOR2_X1 U10588 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(n8221), .ZN(n8250) );
  NAND2_X1 U10589 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(n8250), .ZN(n8222) );
  NAND2_X1 U10590 ( .A1(n8248), .A2(n8249), .ZN(n8224) );
  NAND2_X1 U10591 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(n14311), .ZN(n8226) );
  OAI21_X1 U10592 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n14311), .A(n8226), .ZN(
        n8246) );
  INV_X1 U10593 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n8228) );
  NAND2_X1 U10594 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n8228), .ZN(n8229) );
  NAND2_X1 U10595 ( .A1(n8243), .A2(n8242), .ZN(n8230) );
  INV_X1 U10596 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14640) );
  NAND2_X1 U10597 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14640), .ZN(n8231) );
  AOI22_X1 U10598 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14410), .B1(n8240), 
        .B2(n8231), .ZN(n8239) );
  OAI22_X1 U10599 ( .A1(n8232), .A2(n8239), .B1(P3_ADDR_REG_16__SCAN_IN), .B2(
        n14652), .ZN(n8233) );
  NOR2_X1 U10600 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n8233), .ZN(n8236) );
  INV_X1 U10601 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n8234) );
  XNOR2_X1 U10602 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n8233), .ZN(n8237) );
  NOR2_X1 U10603 ( .A1(n8234), .A2(n8237), .ZN(n8235) );
  NOR2_X1 U10604 ( .A1(n8236), .A2(n8235), .ZN(n8298) );
  XNOR2_X1 U10605 ( .A(n8299), .B(n8298), .ZN(n14379) );
  XNOR2_X1 U10606 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n8237), .ZN(n8295) );
  XOR2_X1 U10607 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .Z(n8238) );
  XNOR2_X1 U10608 ( .A(n8239), .B(n8238), .ZN(n14578) );
  XNOR2_X1 U10609 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .ZN(n8241) );
  XOR2_X1 U10610 ( .A(n8241), .B(n8240), .Z(n8293) );
  XNOR2_X1 U10611 ( .A(n8243), .B(n8242), .ZN(n14570) );
  XOR2_X1 U10612 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .Z(n8244) );
  XOR2_X1 U10613 ( .A(n8245), .B(n8244), .Z(n8289) );
  XNOR2_X1 U10614 ( .A(n8247), .B(n8246), .ZN(n14561) );
  XOR2_X1 U10615 ( .A(n8249), .B(n8248), .Z(n14557) );
  XNOR2_X1 U10616 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n8250), .ZN(n8287) );
  XNOR2_X1 U10617 ( .A(n8252), .B(n8251), .ZN(n8283) );
  INV_X1 U10618 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14349) );
  XNOR2_X1 U10619 ( .A(n14349), .B(n8253), .ZN(n8268) );
  INV_X1 U10620 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14853) );
  NAND2_X1 U10621 ( .A1(n8255), .A2(n14853), .ZN(n8267) );
  XNOR2_X1 U10622 ( .A(P2_ADDR_REG_4__SCAN_IN), .B(n8255), .ZN(n15169) );
  INV_X1 U10623 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n13716) );
  XNOR2_X1 U10624 ( .A(n8256), .B(n13716), .ZN(n15180) );
  XOR2_X1 U10625 ( .A(n8258), .B(n8257), .Z(n14384) );
  INV_X1 U10626 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n8263) );
  NOR2_X1 U10627 ( .A1(n8262), .A2(n8263), .ZN(n8264) );
  OAI21_X1 U10628 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n8261), .A(n8260), .ZN(
        n15173) );
  NAND2_X1 U10629 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15173), .ZN(n15185) );
  XNOR2_X1 U10630 ( .A(n8263), .B(n8262), .ZN(n15184) );
  NOR2_X1 U10631 ( .A1(n15185), .A2(n15184), .ZN(n15183) );
  NOR2_X1 U10632 ( .A1(n14384), .A2(n14383), .ZN(n8265) );
  NAND2_X1 U10633 ( .A1(n14384), .A2(n14383), .ZN(n14382) );
  NOR2_X1 U10634 ( .A1(n15180), .A2(n15181), .ZN(n8266) );
  NAND2_X1 U10635 ( .A1(n15180), .A2(n15181), .ZN(n15179) );
  NAND2_X1 U10636 ( .A1(n15169), .A2(n15168), .ZN(n15167) );
  NAND2_X1 U10637 ( .A1(n8267), .A2(n15167), .ZN(n8269) );
  NAND2_X1 U10638 ( .A1(n8268), .A2(n8269), .ZN(n8270) );
  INV_X1 U10639 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15171) );
  INV_X1 U10640 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n8274) );
  NOR2_X1 U10641 ( .A1(n8275), .A2(n8274), .ZN(n8276) );
  NAND2_X1 U10642 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n15007), .ZN(n8271) );
  OAI21_X1 U10643 ( .B1(n15007), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n8271), .ZN(
        n8273) );
  XOR2_X1 U10644 ( .A(n8273), .B(n8272), .Z(n14388) );
  XNOR2_X1 U10645 ( .A(n8275), .B(n8274), .ZN(n14387) );
  NOR2_X1 U10646 ( .A1(n14388), .A2(n14387), .ZN(n14386) );
  INV_X1 U10647 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n15176) );
  XNOR2_X1 U10648 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n8277), .ZN(n15177) );
  XOR2_X1 U10649 ( .A(n8279), .B(n8278), .Z(n8281) );
  INV_X1 U10650 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14390) );
  NAND2_X1 U10651 ( .A1(n14391), .A2(n14390), .ZN(n14389) );
  NAND2_X1 U10652 ( .A1(n8281), .A2(n8280), .ZN(n8282) );
  NAND2_X1 U10653 ( .A1(n8283), .A2(n8285), .ZN(n8286) );
  INV_X1 U10654 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14393) );
  INV_X1 U10655 ( .A(n14396), .ZN(n14397) );
  INV_X1 U10656 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14399) );
  NAND2_X1 U10657 ( .A1(n8288), .A2(n8287), .ZN(n14398) );
  NAND2_X1 U10658 ( .A1(n14399), .A2(n14398), .ZN(n14395) );
  NAND2_X1 U10659 ( .A1(n14557), .A2(n14558), .ZN(n14556) );
  INV_X1 U10660 ( .A(n14565), .ZN(n14566) );
  INV_X1 U10661 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14870) );
  NAND2_X1 U10662 ( .A1(n8290), .A2(n8289), .ZN(n14567) );
  NAND2_X1 U10663 ( .A1(n14870), .A2(n14567), .ZN(n14564) );
  NOR2_X1 U10664 ( .A1(n14570), .A2(n14569), .ZN(n8291) );
  NAND2_X1 U10665 ( .A1(n14570), .A2(n14569), .ZN(n14568) );
  OAI21_X1 U10666 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(n8291), .A(n14568), .ZN(
        n8292) );
  INV_X1 U10667 ( .A(n14573), .ZN(n14574) );
  INV_X1 U10668 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n14576) );
  NAND2_X1 U10669 ( .A1(n8294), .A2(n8293), .ZN(n14575) );
  NAND2_X1 U10670 ( .A1(n14576), .A2(n14575), .ZN(n14572) );
  NAND2_X1 U10671 ( .A1(n8295), .A2(n8296), .ZN(n8297) );
  INV_X1 U10672 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14401) );
  NAND2_X1 U10673 ( .A1(n14402), .A2(n14401), .ZN(n14400) );
  NAND2_X1 U10674 ( .A1(n8297), .A2(n14400), .ZN(n14378) );
  INV_X1 U10675 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14680) );
  NAND2_X1 U10676 ( .A1(n8299), .A2(n8298), .ZN(n8300) );
  OAI21_X1 U10677 ( .B1(n14680), .B2(P3_ADDR_REG_18__SCAN_IN), .A(n8300), .ZN(
        n8301) );
  NAND2_X1 U10678 ( .A1(n8340), .A2(n13097), .ZN(n8305) );
  NAND2_X1 U10679 ( .A1(n8344), .A2(n8312), .ZN(n8304) );
  AND2_X1 U10680 ( .A1(n8305), .A2(n8304), .ZN(n8316) );
  NAND2_X1 U10681 ( .A1(n8344), .A2(n10252), .ZN(n8306) );
  NAND3_X1 U10682 ( .A1(n8557), .A2(n8307), .A3(n8306), .ZN(n8311) );
  NAND2_X1 U10683 ( .A1(n8308), .A2(n10252), .ZN(n8309) );
  NAND3_X1 U10684 ( .A1(n9465), .A2(n8309), .A3(n8344), .ZN(n8310) );
  NAND2_X1 U10685 ( .A1(n8311), .A2(n8310), .ZN(n8315) );
  INV_X1 U10686 ( .A(n8312), .ZN(n10384) );
  NAND2_X1 U10687 ( .A1(n13097), .A2(n8344), .ZN(n8313) );
  OAI21_X1 U10688 ( .B1(n10384), .B2(n8344), .A(n8313), .ZN(n8314) );
  OAI21_X1 U10689 ( .B1(n8316), .B2(n8315), .A(n8314), .ZN(n8324) );
  NAND2_X1 U10690 ( .A1(n8316), .A2(n8315), .ZN(n8323) );
  NAND2_X1 U10691 ( .A1(n8319), .A2(n8344), .ZN(n8318) );
  NAND2_X1 U10692 ( .A1(n8340), .A2(n13095), .ZN(n8317) );
  AND2_X1 U10693 ( .A1(n8318), .A2(n8317), .ZN(n8326) );
  NAND2_X1 U10694 ( .A1(n8340), .A2(n8319), .ZN(n8321) );
  NAND2_X1 U10695 ( .A1(n13095), .A2(n8344), .ZN(n8320) );
  NAND2_X1 U10696 ( .A1(n8321), .A2(n8320), .ZN(n8325) );
  NAND2_X1 U10697 ( .A1(n8326), .A2(n8325), .ZN(n8322) );
  NAND3_X1 U10698 ( .A1(n8324), .A2(n8323), .A3(n8322), .ZN(n8330) );
  INV_X1 U10699 ( .A(n8325), .ZN(n8328) );
  INV_X1 U10700 ( .A(n8326), .ZN(n8327) );
  NAND2_X1 U10701 ( .A1(n8328), .A2(n8327), .ZN(n8329) );
  NAND2_X1 U10702 ( .A1(n10006), .A2(n8344), .ZN(n8332) );
  NAND2_X1 U10703 ( .A1(n8340), .A2(n13094), .ZN(n8331) );
  NAND2_X1 U10704 ( .A1(n8332), .A2(n8331), .ZN(n8334) );
  NAND2_X1 U10705 ( .A1(n10073), .A2(n8541), .ZN(n8336) );
  NAND2_X1 U10706 ( .A1(n13093), .A2(n8514), .ZN(n8335) );
  NAND2_X1 U10707 ( .A1(n8336), .A2(n8335), .ZN(n8338) );
  AOI22_X1 U10708 ( .A1(n10073), .A2(n8514), .B1(n8340), .B2(n13093), .ZN(
        n8337) );
  NAND2_X1 U10709 ( .A1(n9973), .A2(n8344), .ZN(n8342) );
  NAND2_X1 U10710 ( .A1(n8340), .A2(n13092), .ZN(n8341) );
  NAND2_X1 U10711 ( .A1(n8342), .A2(n8341), .ZN(n8343) );
  NAND2_X1 U10712 ( .A1(n9973), .A2(n8340), .ZN(n8346) );
  NAND2_X1 U10713 ( .A1(n13092), .A2(n8514), .ZN(n8345) );
  NAND2_X1 U10714 ( .A1(n8346), .A2(n8345), .ZN(n8347) );
  NAND2_X1 U10715 ( .A1(n10274), .A2(n8541), .ZN(n8349) );
  NAND2_X1 U10716 ( .A1(n13091), .A2(n8344), .ZN(n8348) );
  AOI22_X1 U10717 ( .A1(n10274), .A2(n8344), .B1(n8541), .B2(n13091), .ZN(
        n8350) );
  NAND2_X1 U10718 ( .A1(n10289), .A2(n8514), .ZN(n8352) );
  NAND2_X1 U10719 ( .A1(n8541), .A2(n13090), .ZN(n8351) );
  NAND2_X1 U10720 ( .A1(n8352), .A2(n8351), .ZN(n8354) );
  AOI22_X1 U10721 ( .A1(n10289), .A2(n8541), .B1(n13090), .B2(n8514), .ZN(
        n8353) );
  AOI21_X1 U10722 ( .B1(n8355), .B2(n8354), .A(n8353), .ZN(n8356) );
  NAND2_X1 U10723 ( .A1(n12975), .A2(n8541), .ZN(n8358) );
  NAND2_X1 U10724 ( .A1(n13089), .A2(n8514), .ZN(n8357) );
  NAND2_X1 U10725 ( .A1(n8358), .A2(n8357), .ZN(n8361) );
  NAND2_X1 U10726 ( .A1(n12975), .A2(n8514), .ZN(n8360) );
  NAND2_X1 U10727 ( .A1(n8541), .A2(n13089), .ZN(n8359) );
  NAND2_X1 U10728 ( .A1(n10424), .A2(n8514), .ZN(n8366) );
  NAND2_X1 U10729 ( .A1(n8541), .A2(n13088), .ZN(n8365) );
  NAND2_X1 U10730 ( .A1(n8366), .A2(n8365), .ZN(n8369) );
  AOI22_X1 U10731 ( .A1(n10424), .A2(n8541), .B1(n13088), .B2(n8514), .ZN(
        n8367) );
  NAND2_X1 U10732 ( .A1(n12966), .A2(n8340), .ZN(n8372) );
  NAND2_X1 U10733 ( .A1(n13087), .A2(n8514), .ZN(n8371) );
  NAND2_X1 U10734 ( .A1(n8372), .A2(n8371), .ZN(n8375) );
  NAND2_X1 U10735 ( .A1(n12966), .A2(n8514), .ZN(n8374) );
  NAND2_X1 U10736 ( .A1(n8541), .A2(n13087), .ZN(n8373) );
  NAND2_X1 U10737 ( .A1(n12126), .A2(n8514), .ZN(n8377) );
  NAND2_X1 U10738 ( .A1(n8541), .A2(n13086), .ZN(n8376) );
  NAND2_X1 U10739 ( .A1(n8377), .A2(n8376), .ZN(n8379) );
  AOI22_X1 U10740 ( .A1(n12126), .A2(n8541), .B1(n13086), .B2(n8514), .ZN(
        n8378) );
  AOI21_X1 U10741 ( .B1(n8380), .B2(n8379), .A(n8378), .ZN(n8381) );
  NAND2_X1 U10742 ( .A1(n12100), .A2(n8340), .ZN(n8383) );
  NAND2_X1 U10743 ( .A1(n13085), .A2(n8514), .ZN(n8382) );
  INV_X1 U10744 ( .A(n13085), .ZN(n10901) );
  NAND2_X1 U10745 ( .A1(n12100), .A2(n8514), .ZN(n8384) );
  OAI21_X1 U10746 ( .B1(n10901), .B2(n8514), .A(n8384), .ZN(n8385) );
  NAND2_X1 U10747 ( .A1(n11146), .A2(n8514), .ZN(n8388) );
  NAND2_X1 U10748 ( .A1(n8541), .A2(n13084), .ZN(n8387) );
  NAND2_X1 U10749 ( .A1(n8388), .A2(n8387), .ZN(n8390) );
  AOI22_X1 U10750 ( .A1(n11146), .A2(n8541), .B1(n13084), .B2(n8514), .ZN(
        n8389) );
  AOI21_X1 U10751 ( .B1(n8391), .B2(n8390), .A(n8389), .ZN(n8392) );
  NAND2_X1 U10752 ( .A1(n14508), .A2(n8340), .ZN(n8394) );
  NAND2_X1 U10753 ( .A1(n13083), .A2(n8514), .ZN(n8393) );
  NAND2_X1 U10754 ( .A1(n8394), .A2(n8393), .ZN(n8399) );
  NAND2_X1 U10755 ( .A1(n8398), .A2(n8399), .ZN(n8397) );
  INV_X1 U10756 ( .A(n13083), .ZN(n9235) );
  NAND2_X1 U10757 ( .A1(n14508), .A2(n8514), .ZN(n8395) );
  OAI21_X1 U10758 ( .B1(n9235), .B2(n8514), .A(n8395), .ZN(n8396) );
  NAND2_X1 U10759 ( .A1(n8397), .A2(n8396), .ZN(n8403) );
  INV_X1 U10760 ( .A(n8398), .ZN(n8401) );
  INV_X1 U10761 ( .A(n8399), .ZN(n8400) );
  NAND2_X1 U10762 ( .A1(n8401), .A2(n8400), .ZN(n8402) );
  NAND2_X1 U10763 ( .A1(n11273), .A2(n8514), .ZN(n8405) );
  NAND2_X1 U10764 ( .A1(n13082), .A2(n8541), .ZN(n8404) );
  NAND2_X1 U10765 ( .A1(n8405), .A2(n8404), .ZN(n8407) );
  AOI22_X1 U10766 ( .A1(n11273), .A2(n8541), .B1(n13082), .B2(n8514), .ZN(
        n8406) );
  NAND2_X1 U10767 ( .A1(n13504), .A2(n8541), .ZN(n8409) );
  NAND2_X1 U10768 ( .A1(n13081), .A2(n8514), .ZN(n8408) );
  NAND2_X1 U10769 ( .A1(n8409), .A2(n8408), .ZN(n8412) );
  AOI22_X1 U10770 ( .A1(n13504), .A2(n8514), .B1(n8541), .B2(n13081), .ZN(
        n8410) );
  AOI21_X1 U10771 ( .B1(n8413), .B2(n8412), .A(n8410), .ZN(n8411) );
  NOR2_X1 U10772 ( .A1(n8413), .A2(n8412), .ZN(n8414) );
  NAND2_X1 U10773 ( .A1(n13498), .A2(n8514), .ZN(n8416) );
  NAND2_X1 U10774 ( .A1(n13080), .A2(n8340), .ZN(n8415) );
  NAND2_X1 U10775 ( .A1(n8416), .A2(n8415), .ZN(n8419) );
  INV_X1 U10776 ( .A(n13080), .ZN(n14517) );
  NAND2_X1 U10777 ( .A1(n13498), .A2(n8541), .ZN(n8417) );
  OAI21_X1 U10778 ( .B1(n14517), .B2(n8541), .A(n8417), .ZN(n8418) );
  NAND2_X1 U10779 ( .A1(n13493), .A2(n8541), .ZN(n8422) );
  NAND2_X1 U10780 ( .A1(n13079), .A2(n8514), .ZN(n8421) );
  NAND2_X1 U10781 ( .A1(n8422), .A2(n8421), .ZN(n8424) );
  AOI22_X1 U10782 ( .A1(n13493), .A2(n8514), .B1(n8541), .B2(n13079), .ZN(
        n8423) );
  NAND2_X1 U10783 ( .A1(n13488), .A2(n8514), .ZN(n8427) );
  NAND2_X1 U10784 ( .A1(n13371), .A2(n8340), .ZN(n8426) );
  NAND2_X1 U10785 ( .A1(n8427), .A2(n8426), .ZN(n8432) );
  INV_X1 U10786 ( .A(n13371), .ZN(n13053) );
  NAND2_X1 U10787 ( .A1(n13488), .A2(n8541), .ZN(n8428) );
  OAI21_X1 U10788 ( .B1(n13053), .B2(n8541), .A(n8428), .ZN(n8429) );
  NAND2_X1 U10789 ( .A1(n8430), .A2(n8429), .ZN(n8436) );
  INV_X1 U10790 ( .A(n8431), .ZN(n8434) );
  NAND2_X1 U10791 ( .A1(n8434), .A2(n8433), .ZN(n8435) );
  NAND2_X1 U10792 ( .A1(n13481), .A2(n8541), .ZN(n8438) );
  NAND2_X1 U10793 ( .A1(n13358), .A2(n8514), .ZN(n8437) );
  NAND2_X1 U10794 ( .A1(n8438), .A2(n8437), .ZN(n8440) );
  AOI22_X1 U10795 ( .A1(n13481), .A2(n8514), .B1(n8541), .B2(n13358), .ZN(
        n8439) );
  NAND2_X1 U10796 ( .A1(n13477), .A2(n8514), .ZN(n8443) );
  NAND2_X1 U10797 ( .A1(n13373), .A2(n8541), .ZN(n8442) );
  NAND2_X1 U10798 ( .A1(n8443), .A2(n8442), .ZN(n8446) );
  INV_X1 U10799 ( .A(n13373), .ZN(n13045) );
  NAND2_X1 U10800 ( .A1(n13477), .A2(n8541), .ZN(n8444) );
  OAI21_X1 U10801 ( .B1(n13045), .B2(n8541), .A(n8444), .ZN(n8445) );
  NAND2_X1 U10802 ( .A1(n13472), .A2(n8541), .ZN(n8448) );
  NAND2_X1 U10803 ( .A1(n13357), .A2(n8344), .ZN(n8447) );
  NAND2_X1 U10804 ( .A1(n8448), .A2(n8447), .ZN(n8450) );
  AOI22_X1 U10805 ( .A1(n13472), .A2(n8514), .B1(n8541), .B2(n13357), .ZN(
        n8449) );
  NAND2_X1 U10806 ( .A1(n13465), .A2(n8514), .ZN(n8454) );
  NAND2_X1 U10807 ( .A1(n13338), .A2(n8340), .ZN(n8453) );
  AOI22_X1 U10808 ( .A1(n13465), .A2(n8541), .B1(n13338), .B2(n8514), .ZN(
        n8455) );
  NAND2_X1 U10809 ( .A1(n13462), .A2(n8340), .ZN(n8457) );
  NAND2_X1 U10810 ( .A1(n13078), .A2(n8514), .ZN(n8456) );
  NAND2_X1 U10811 ( .A1(n8457), .A2(n8456), .ZN(n8460) );
  INV_X1 U10812 ( .A(n13078), .ZN(n11534) );
  NAND2_X1 U10813 ( .A1(n13462), .A2(n8514), .ZN(n8458) );
  OAI21_X1 U10814 ( .B1(n11534), .B2(n8514), .A(n8458), .ZN(n8459) );
  NAND2_X1 U10815 ( .A1(n13456), .A2(n8514), .ZN(n8462) );
  NAND2_X1 U10816 ( .A1(n13077), .A2(n8340), .ZN(n8461) );
  NAND2_X1 U10817 ( .A1(n8462), .A2(n8461), .ZN(n8464) );
  AOI22_X1 U10818 ( .A1(n13451), .A2(n8541), .B1(n13076), .B2(n8514), .ZN(
        n8537) );
  OAI22_X1 U10819 ( .A1(n13282), .A2(n8340), .B1(n11558), .B2(n8514), .ZN(
        n8536) );
  AOI22_X1 U10820 ( .A1(n13456), .A2(n8541), .B1(n13077), .B2(n8514), .ZN(
        n8463) );
  INV_X1 U10821 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14369) );
  INV_X1 U10822 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13545) );
  MUX2_X1 U10823 ( .A(n14369), .B(n13545), .S(n6450), .Z(n8467) );
  XNOR2_X1 U10824 ( .A(n8467), .B(SI_29_), .ZN(n8485) );
  INV_X1 U10825 ( .A(SI_29_), .ZN(n12937) );
  NAND2_X1 U10826 ( .A1(n8467), .A2(n12937), .ZN(n8495) );
  NAND2_X1 U10827 ( .A1(n8504), .A2(n8495), .ZN(n8471) );
  MUX2_X1 U10828 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6450), .Z(n8468) );
  NAND2_X1 U10829 ( .A1(n8468), .A2(SI_30_), .ZN(n8498) );
  INV_X1 U10830 ( .A(n8468), .ZN(n8469) );
  INV_X1 U10831 ( .A(SI_30_), .ZN(n12332) );
  NAND2_X1 U10832 ( .A1(n8469), .A2(n12332), .ZN(n8496) );
  AND2_X1 U10833 ( .A1(n8498), .A2(n8496), .ZN(n8470) );
  NAND2_X1 U10834 ( .A1(n11850), .A2(n8509), .ZN(n8473) );
  INV_X1 U10835 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12338) );
  OR2_X1 U10836 ( .A1(n8487), .A2(n12338), .ZN(n8472) );
  NAND2_X2 U10837 ( .A1(n8473), .A2(n8472), .ZN(n13241) );
  INV_X1 U10838 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n13238) );
  NAND2_X1 U10839 ( .A1(n8069), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8475) );
  NAND2_X1 U10840 ( .A1(n8477), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8474) );
  OAI211_X1 U10841 ( .C1(n8480), .C2(n13238), .A(n8475), .B(n8474), .ZN(n13072) );
  AND2_X1 U10842 ( .A1(n8541), .A2(n13072), .ZN(n8476) );
  AOI21_X1 U10843 ( .B1(n13241), .B2(n8514), .A(n8476), .ZN(n8535) );
  NAND2_X1 U10844 ( .A1(n13241), .A2(n8340), .ZN(n8484) );
  INV_X1 U10845 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n13230) );
  NAND2_X1 U10846 ( .A1(n8069), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8479) );
  NAND2_X1 U10847 ( .A1(n8477), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8478) );
  OAI211_X1 U10848 ( .C1(n8480), .C2(n13230), .A(n8479), .B(n8478), .ZN(n13231) );
  NAND2_X1 U10849 ( .A1(n13231), .A2(n8514), .ZN(n8540) );
  NOR2_X1 U10850 ( .A1(n11264), .A2(n13226), .ZN(n9464) );
  NAND2_X1 U10851 ( .A1(n9464), .A2(n11102), .ZN(n8481) );
  NAND4_X1 U10852 ( .A1(n8540), .A2(n7517), .A3(n8577), .A4(n8481), .ZN(n8482)
         );
  NAND2_X1 U10853 ( .A1(n8482), .A2(n13072), .ZN(n8483) );
  NAND2_X1 U10854 ( .A1(n8484), .A2(n8483), .ZN(n8534) );
  NAND2_X1 U10855 ( .A1(n8535), .A2(n8534), .ZN(n8494) );
  NAND2_X1 U10856 ( .A1(n13544), .A2(n8509), .ZN(n8489) );
  OR2_X1 U10857 ( .A1(n8487), .A2(n13545), .ZN(n8488) );
  AND2_X1 U10858 ( .A1(n13073), .A2(n8541), .ZN(n8490) );
  AOI21_X1 U10859 ( .B1(n13434), .B2(n8514), .A(n8490), .ZN(n8529) );
  NAND2_X1 U10860 ( .A1(n13434), .A2(n8340), .ZN(n8492) );
  NAND2_X1 U10861 ( .A1(n13073), .A2(n8514), .ZN(n8491) );
  NAND2_X1 U10862 ( .A1(n8492), .A2(n8491), .ZN(n8528) );
  NAND2_X1 U10863 ( .A1(n8529), .A2(n8528), .ZN(n8493) );
  NAND2_X1 U10864 ( .A1(n8496), .A2(n8495), .ZN(n8502) );
  MUX2_X1 U10865 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6449), .Z(n8497) );
  XNOR2_X1 U10866 ( .A(n8497), .B(SI_31_), .ZN(n8500) );
  NOR2_X1 U10867 ( .A1(n8502), .A2(n8500), .ZN(n8508) );
  XNOR2_X1 U10868 ( .A(n8500), .B(n8498), .ZN(n8507) );
  INV_X1 U10869 ( .A(n8498), .ZN(n8499) );
  INV_X1 U10870 ( .A(n8500), .ZN(n8501) );
  NOR2_X1 U10871 ( .A1(n8502), .A2(n8501), .ZN(n8503) );
  NAND2_X1 U10872 ( .A1(n8504), .A2(n8503), .ZN(n8505) );
  NAND2_X1 U10873 ( .A1(n14222), .A2(n8509), .ZN(n8512) );
  NAND2_X1 U10874 ( .A1(n8510), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8511) );
  AND2_X1 U10875 ( .A1(n13074), .A2(n8541), .ZN(n8513) );
  AOI21_X1 U10876 ( .B1(n13438), .B2(n8514), .A(n8513), .ZN(n8527) );
  NAND2_X1 U10877 ( .A1(n13438), .A2(n8340), .ZN(n8516) );
  NAND2_X1 U10878 ( .A1(n13074), .A2(n8514), .ZN(n8515) );
  NAND2_X1 U10879 ( .A1(n8516), .A2(n8515), .ZN(n8526) );
  NAND2_X1 U10880 ( .A1(n8527), .A2(n8526), .ZN(n8517) );
  AND2_X1 U10881 ( .A1(n13075), .A2(n8541), .ZN(n8518) );
  AOI21_X1 U10882 ( .B1(n13444), .B2(n8344), .A(n8518), .ZN(n8523) );
  NAND2_X1 U10883 ( .A1(n13444), .A2(n8340), .ZN(n8520) );
  NAND2_X1 U10884 ( .A1(n13075), .A2(n8514), .ZN(n8519) );
  NAND2_X1 U10885 ( .A1(n8520), .A2(n8519), .ZN(n8522) );
  AND2_X1 U10886 ( .A1(n8523), .A2(n8522), .ZN(n8521) );
  NOR2_X1 U10887 ( .A1(n8524), .A2(n8521), .ZN(n8538) );
  INV_X1 U10888 ( .A(n8525), .ZN(n8570) );
  OAI22_X1 U10889 ( .A1(n8529), .A2(n8528), .B1(n8527), .B2(n8526), .ZN(n8531)
         );
  OAI21_X1 U10890 ( .B1(n8570), .B2(n8531), .A(n8530), .ZN(n8532) );
  OAI211_X1 U10891 ( .C1(n8535), .C2(n8534), .A(n8533), .B(n8532), .ZN(n8539)
         );
  AND2_X1 U10892 ( .A1(n8541), .A2(n13231), .ZN(n8544) );
  INV_X1 U10893 ( .A(n8540), .ZN(n8542) );
  NOR2_X1 U10894 ( .A1(n8542), .A2(n8541), .ZN(n8543) );
  MUX2_X1 U10895 ( .A(n8544), .B(n8543), .S(n13427), .Z(n8545) );
  INV_X1 U10896 ( .A(n11264), .ZN(n8580) );
  MUX2_X1 U10897 ( .A(n7517), .B(n8580), .S(n11102), .Z(n8548) );
  INV_X1 U10898 ( .A(n8577), .ZN(n8549) );
  AOI211_X1 U10899 ( .C1(n7517), .C2(n13226), .A(n8549), .B(n8303), .ZN(n8550)
         );
  NAND2_X1 U10900 ( .A1(n8552), .A2(n8550), .ZN(n8551) );
  INV_X1 U10901 ( .A(n9430), .ZN(n9429) );
  AND2_X1 U10902 ( .A1(n9429), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11328) );
  INV_X1 U10903 ( .A(n11328), .ZN(n8579) );
  OAI211_X1 U10904 ( .C1(n8552), .C2(n6603), .A(n8551), .B(n11328), .ZN(n8583)
         );
  NAND2_X1 U10905 ( .A1(n8552), .A2(n11102), .ZN(n8576) );
  NAND2_X1 U10906 ( .A1(n13438), .A2(n13074), .ZN(n11562) );
  OR2_X1 U10907 ( .A1(n13438), .A2(n13074), .ZN(n8553) );
  INV_X1 U10908 ( .A(n13075), .ZN(n11560) );
  XNOR2_X1 U10909 ( .A(n13444), .B(n11560), .ZN(n13270) );
  XNOR2_X1 U10910 ( .A(n13451), .B(n11558), .ZN(n13276) );
  INV_X1 U10911 ( .A(n13357), .ZN(n12987) );
  INV_X1 U10912 ( .A(n13338), .ZN(n13046) );
  OR2_X1 U10913 ( .A1(n13465), .A2(n13046), .ZN(n11531) );
  NAND2_X1 U10914 ( .A1(n13465), .A2(n13046), .ZN(n11532) );
  NAND2_X1 U10915 ( .A1(n11531), .A2(n11532), .ZN(n13328) );
  XNOR2_X1 U10916 ( .A(n13456), .B(n13077), .ZN(n13291) );
  XNOR2_X1 U10917 ( .A(n13481), .B(n13358), .ZN(n13376) );
  XNOR2_X1 U10918 ( .A(n13488), .B(n13053), .ZN(n13392) );
  INV_X1 U10919 ( .A(n13079), .ZN(n11525) );
  XNOR2_X1 U10920 ( .A(n13493), .B(n11525), .ZN(n13403) );
  XNOR2_X1 U10921 ( .A(n13504), .B(n11391), .ZN(n11201) );
  NAND2_X1 U10922 ( .A1(n13498), .A2(n14517), .ZN(n8554) );
  NAND2_X1 U10923 ( .A1(n11523), .A2(n8554), .ZN(n11389) );
  INV_X1 U10924 ( .A(n13082), .ZN(n14520) );
  XNOR2_X1 U10925 ( .A(n11273), .B(n14520), .ZN(n11267) );
  NAND2_X1 U10926 ( .A1(n14508), .A2(n9235), .ZN(n11198) );
  OR2_X1 U10927 ( .A1(n14508), .A2(n9235), .ZN(n8555) );
  NAND2_X1 U10928 ( .A1(n11198), .A2(n8555), .ZN(n11149) );
  XNOR2_X1 U10929 ( .A(n11146), .B(n14499), .ZN(n10908) );
  XNOR2_X1 U10930 ( .A(n12100), .B(n10901), .ZN(n10673) );
  INV_X1 U10931 ( .A(n13086), .ZN(n12960) );
  XNOR2_X1 U10932 ( .A(n12126), .B(n12960), .ZN(n10475) );
  INV_X1 U10933 ( .A(n13088), .ZN(n12972) );
  NAND2_X1 U10934 ( .A1(n10424), .A2(n12972), .ZN(n10427) );
  OR2_X1 U10935 ( .A1(n10424), .A2(n12972), .ZN(n8556) );
  INV_X1 U10936 ( .A(n13090), .ZN(n10288) );
  XNOR2_X1 U10937 ( .A(n10289), .B(n10288), .ZN(n10021) );
  XNOR2_X1 U10938 ( .A(n10274), .B(n13091), .ZN(n9925) );
  OR2_X1 U10939 ( .A1(n9465), .A2(n9857), .ZN(n9461) );
  AND2_X1 U10940 ( .A1(n9461), .A2(n8557), .ZN(n10249) );
  NAND4_X1 U10941 ( .A1(n10249), .A2(n9462), .A3(n9582), .A4(n9630), .ZN(n8558) );
  NOR2_X1 U10942 ( .A1(n9721), .A2(n8558), .ZN(n8559) );
  XNOR2_X1 U10943 ( .A(n9973), .B(n13092), .ZN(n9785) );
  XNOR2_X1 U10944 ( .A(n10073), .B(n13093), .ZN(n9787) );
  NAND4_X1 U10945 ( .A1(n9925), .A2(n8559), .A3(n9785), .A4(n9787), .ZN(n8560)
         );
  NOR2_X1 U10946 ( .A1(n10021), .A2(n8560), .ZN(n8561) );
  XNOR2_X1 U10947 ( .A(n12975), .B(n13089), .ZN(n10391) );
  NAND4_X1 U10948 ( .A1(n10429), .A2(n10396), .A3(n8561), .A4(n10391), .ZN(
        n8562) );
  OR4_X1 U10949 ( .A1(n10908), .A2(n10673), .A3(n10475), .A4(n8562), .ZN(n8563) );
  OR4_X1 U10950 ( .A1(n11389), .A2(n11267), .A3(n11149), .A4(n8563), .ZN(n8564) );
  OR3_X1 U10951 ( .A1(n13403), .A2(n11201), .A3(n8564), .ZN(n8565) );
  NOR2_X1 U10952 ( .A1(n13392), .A2(n8565), .ZN(n8566) );
  AND2_X1 U10953 ( .A1(n13376), .A2(n8566), .ZN(n8567) );
  XNOR2_X1 U10954 ( .A(n13462), .B(n13078), .ZN(n13308) );
  XNOR2_X1 U10955 ( .A(n13477), .B(n13373), .ZN(n13355) );
  NAND4_X1 U10956 ( .A1(n13291), .A2(n8567), .A3(n13308), .A4(n13355), .ZN(
        n8568) );
  NOR4_X1 U10957 ( .A1(n8570), .A2(n13249), .A3(n13270), .A4(n8569), .ZN(n8572) );
  XNOR2_X1 U10958 ( .A(n13241), .B(n13072), .ZN(n8571) );
  NAND3_X1 U10959 ( .A1(n8572), .A2(n11563), .A3(n8571), .ZN(n8573) );
  NAND2_X1 U10960 ( .A1(n11328), .A2(n11099), .ZN(n8574) );
  OR4_X1 U10961 ( .A1(n14872), .A2(n6698), .A3(n13051), .A4(n8577), .ZN(n8578)
         );
  OAI211_X1 U10962 ( .C1(n8580), .C2(n8579), .A(n8578), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8581) );
  NAND3_X1 U10963 ( .A1(n8583), .A2(n8582), .A3(n8581), .ZN(P2_U3328) );
  NOR2_X1 U10964 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n8586) );
  NAND2_X1 U10965 ( .A1(n8955), .A2(n8591), .ZN(n8967) );
  INV_X1 U10966 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8589) );
  XNOR2_X2 U10967 ( .A(n8590), .B(n8589), .ZN(n12654) );
  NAND2_X1 U10968 ( .A1(n9160), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8594) );
  NAND2_X1 U10969 ( .A1(n8595), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8596) );
  MUX2_X1 U10970 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8596), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8597) );
  NAND2_X1 U10971 ( .A1(n12415), .A2(n10196), .ZN(n8598) );
  NAND2_X1 U10972 ( .A1(n12404), .A2(n8598), .ZN(n8602) );
  NAND2_X1 U10973 ( .A1(n8599), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8600) );
  MUX2_X1 U10974 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8600), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n8601) );
  INV_X2 U10975 ( .A(n12195), .ZN(n10414) );
  NAND2_X1 U10976 ( .A1(n8602), .A2(n10414), .ZN(n8605) );
  INV_X1 U10977 ( .A(n12415), .ZN(n9134) );
  NAND2_X1 U10978 ( .A1(n10414), .A2(n10196), .ZN(n8603) );
  NAND2_X1 U10979 ( .A1(n9134), .A2(n8603), .ZN(n8604) );
  NAND2_X1 U10980 ( .A1(n8605), .A2(n8604), .ZN(n9883) );
  NAND2_X1 U10981 ( .A1(n12654), .A2(n10196), .ZN(n9167) );
  INV_X1 U10982 ( .A(n9167), .ZN(n12411) );
  NAND2_X1 U10983 ( .A1(n9134), .A2(n10414), .ZN(n15144) );
  NAND3_X1 U10984 ( .A1(n9883), .A2(n12411), .A3(n15144), .ZN(n8607) );
  AND2_X1 U10985 ( .A1(n12415), .A2(n9165), .ZN(n8606) );
  NAND2_X1 U10986 ( .A1(n12654), .A2(n8606), .ZN(n9133) );
  NAND2_X1 U10987 ( .A1(n8607), .A2(n9133), .ZN(n15125) );
  AND2_X1 U10988 ( .A1(n12404), .A2(n10196), .ZN(n10603) );
  INV_X1 U10989 ( .A(n15150), .ZN(n14483) );
  XNOR2_X1 U10990 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8741) );
  NAND2_X1 U10991 ( .A1(n8608), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8740) );
  INV_X1 U10992 ( .A(n8740), .ZN(n8609) );
  NAND2_X1 U10993 ( .A1(n8741), .A2(n8609), .ZN(n8611) );
  NAND2_X1 U10994 ( .A1(n9355), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8610) );
  NAND2_X1 U10995 ( .A1(n8611), .A2(n8610), .ZN(n8746) );
  NAND2_X1 U10996 ( .A1(n9759), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8612) );
  NAND2_X1 U10997 ( .A1(n8746), .A2(n8612), .ZN(n8614) );
  NAND2_X1 U10998 ( .A1(n9370), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8613) );
  NAND2_X1 U10999 ( .A1(n8614), .A2(n8613), .ZN(n8758) );
  NAND2_X1 U11000 ( .A1(n10147), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8616) );
  INV_X1 U11001 ( .A(n8770), .ZN(n8617) );
  INV_X1 U11002 ( .A(n8784), .ZN(n8618) );
  NAND2_X1 U11003 ( .A1(n8785), .A2(n8618), .ZN(n8620) );
  NAND2_X1 U11004 ( .A1(n9364), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8619) );
  NAND2_X1 U11005 ( .A1(n9367), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8621) );
  INV_X1 U11006 ( .A(n8802), .ZN(n8622) );
  XNOR2_X1 U11007 ( .A(n9387), .B(P2_DATAO_REG_8__SCAN_IN), .ZN(n8834) );
  INV_X1 U11008 ( .A(n8834), .ZN(n8624) );
  NAND2_X1 U11009 ( .A1(n9387), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8625) );
  NAND2_X1 U11010 ( .A1(n9403), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8628) );
  NAND2_X1 U11011 ( .A1(n9404), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8627) );
  NAND2_X1 U11012 ( .A1(n8628), .A2(n8627), .ZN(n8864) );
  NAND2_X1 U11013 ( .A1(n9419), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8632) );
  NAND2_X1 U11014 ( .A1(n9413), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8629) );
  NAND2_X1 U11015 ( .A1(n8632), .A2(n8629), .ZN(n8844) );
  INV_X1 U11016 ( .A(n8844), .ZN(n8630) );
  NAND2_X1 U11017 ( .A1(n9454), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8633) );
  XNOR2_X1 U11018 ( .A(n8635), .B(P1_DATAO_REG_12__SCAN_IN), .ZN(n8907) );
  INV_X1 U11019 ( .A(n8907), .ZN(n8634) );
  NAND2_X1 U11020 ( .A1(n8635), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8636) );
  INV_X1 U11021 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9654) );
  NAND2_X1 U11022 ( .A1(n8638), .A2(n9654), .ZN(n8639) );
  INV_X1 U11023 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9819) );
  AND2_X1 U11024 ( .A1(n9819), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8641) );
  INV_X1 U11025 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9821) );
  NAND2_X1 U11026 ( .A1(n9821), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8642) );
  NAND2_X1 U11027 ( .A1(n10086), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8644) );
  INV_X1 U11028 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10087) );
  NAND2_X1 U11029 ( .A1(n10087), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8643) );
  NAND2_X1 U11030 ( .A1(n8644), .A2(n8643), .ZN(n8937) );
  NAND2_X1 U11031 ( .A1(n10215), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8646) );
  NAND2_X1 U11032 ( .A1(n10217), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8645) );
  INV_X1 U11033 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10315) );
  NAND2_X1 U11034 ( .A1(n10315), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8647) );
  INV_X1 U11035 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10314) );
  NAND2_X1 U11036 ( .A1(n10314), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8648) );
  XNOR2_X1 U11037 ( .A(n10513), .B(P1_DATAO_REG_18__SCAN_IN), .ZN(n8978) );
  INV_X1 U11038 ( .A(n8978), .ZN(n8650) );
  NAND2_X1 U11039 ( .A1(n10513), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8651) );
  NOR2_X1 U11040 ( .A1(n10944), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8653) );
  NAND2_X1 U11041 ( .A1(n10944), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8654) );
  INV_X1 U11042 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11648) );
  NAND2_X1 U11043 ( .A1(n11648), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8657) );
  INV_X1 U11044 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11104) );
  NAND2_X1 U11045 ( .A1(n11104), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8655) );
  INV_X1 U11046 ( .A(n9003), .ZN(n8656) );
  INV_X1 U11047 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11101) );
  XNOR2_X1 U11048 ( .A(n11101), .B(P2_DATAO_REG_21__SCAN_IN), .ZN(n9015) );
  INV_X1 U11049 ( .A(n9015), .ZN(n8658) );
  NAND2_X1 U11050 ( .A1(n11101), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8660) );
  XNOR2_X1 U11051 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .ZN(n9027) );
  INV_X1 U11052 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11266) );
  XNOR2_X1 U11053 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n9036) );
  INV_X1 U11054 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8661) );
  NAND2_X1 U11055 ( .A1(n8661), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8662) );
  INV_X1 U11056 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11088) );
  NAND2_X1 U11057 ( .A1(n8664), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8665) );
  NAND2_X1 U11058 ( .A1(n11738), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8667) );
  NAND2_X1 U11059 ( .A1(n11172), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8666) );
  NAND2_X1 U11060 ( .A1(n8667), .A2(n8666), .ZN(n9055) );
  NAND2_X1 U11061 ( .A1(n11760), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8670) );
  NAND2_X1 U11062 ( .A1(n11336), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8668) );
  NAND2_X1 U11063 ( .A1(n8670), .A2(n8668), .ZN(n9068) );
  INV_X1 U11064 ( .A(n9068), .ZN(n8669) );
  INV_X1 U11065 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14373) );
  NAND2_X1 U11066 ( .A1(n14373), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8673) );
  INV_X1 U11067 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13550) );
  NAND2_X1 U11068 ( .A1(n13550), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8671) );
  NAND2_X1 U11069 ( .A1(n8673), .A2(n8671), .ZN(n9082) );
  INV_X1 U11070 ( .A(n9082), .ZN(n8672) );
  NAND2_X1 U11071 ( .A1(n14257), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9182) );
  NAND2_X1 U11072 ( .A1(n11503), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8675) );
  NAND2_X1 U11073 ( .A1(n9182), .A2(n8675), .ZN(n9179) );
  XNOR2_X1 U11074 ( .A(n9181), .B(n9179), .ZN(n12938) );
  NOR2_X1 U11075 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), 
        .ZN(n8679) );
  XNOR2_X2 U11076 ( .A(n8683), .B(n8682), .ZN(n9130) );
  NAND2_X1 U11077 ( .A1(n12938), .A2(n12343), .ZN(n8686) );
  OR2_X1 U11078 ( .A1(n12333), .A2(n12940), .ZN(n8685) );
  NAND2_X1 U11079 ( .A1(n8687), .A2(n10594), .ZN(n8778) );
  INV_X1 U11080 ( .A(n8778), .ZN(n8688) );
  NAND2_X1 U11081 ( .A1(n8688), .A2(n10709), .ZN(n8794) );
  NAND2_X1 U11082 ( .A1(n11430), .A2(n14291), .ZN(n8692) );
  INV_X1 U11083 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8693) );
  INV_X1 U11084 ( .A(n8930), .ZN(n8696) );
  INV_X1 U11085 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n8695) );
  INV_X1 U11086 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n8697) );
  INV_X1 U11087 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n12469) );
  INV_X1 U11088 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n8700) );
  INV_X1 U11089 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n8701) );
  INV_X1 U11090 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n8703) );
  INV_X1 U11091 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n14320) );
  INV_X1 U11092 ( .A(n9072), .ZN(n8707) );
  INV_X1 U11093 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n8706) );
  INV_X1 U11094 ( .A(n9088), .ZN(n8708) );
  INV_X1 U11095 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n12184) );
  NAND2_X1 U11096 ( .A1(n8708), .A2(n12184), .ZN(n12420) );
  NAND2_X1 U11097 ( .A1(n9088), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8709) );
  NAND2_X1 U11098 ( .A1(n12420), .A2(n8709), .ZN(n12183) );
  OR2_X1 U11099 ( .A1(P3_IR_REG_28__SCAN_IN), .A2(P3_IR_REG_29__SCAN_IN), .ZN(
        n8710) );
  OR2_X2 U11100 ( .A1(n8712), .A2(n8710), .ZN(n12930) );
  NAND2_X2 U11101 ( .A1(n12930), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8711) );
  XNOR2_X2 U11102 ( .A(n8711), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8714) );
  NAND2_X1 U11104 ( .A1(n12183), .A2(n9089), .ZN(n8720) );
  INV_X1 U11105 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12664) );
  INV_X1 U11106 ( .A(n8714), .ZN(n11501) );
  NAND2_X1 U11107 ( .A1(n12346), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8717) );
  NAND2_X1 U11108 ( .A1(n6445), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8716) );
  OAI211_X1 U11109 ( .C1(n12350), .C2(n12664), .A(n8717), .B(n8716), .ZN(n8718) );
  INV_X1 U11110 ( .A(n8718), .ZN(n8719) );
  XNOR2_X2 U11111 ( .A(n12670), .B(n12537), .ZN(n12321) );
  NAND2_X1 U11112 ( .A1(n9188), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8724) );
  NAND2_X1 U11113 ( .A1(n9089), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8723) );
  OR2_X1 U11114 ( .A1(n8756), .A2(n14225), .ZN(n8728) );
  NAND2_X1 U11115 ( .A1(n8725), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8726) );
  AND2_X1 U11116 ( .A1(n8740), .A2(n8726), .ZN(n9332) );
  OAI211_X1 U11117 ( .C1(n14322), .C2(n9834), .A(n8728), .B(n8727), .ZN(n9882)
         );
  NAND2_X1 U11118 ( .A1(n8753), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8735) );
  INV_X1 U11119 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n9829) );
  OR2_X1 U11120 ( .A1(n8729), .A2(n9829), .ZN(n8734) );
  INV_X1 U11121 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10608) );
  OR2_X1 U11122 ( .A1(n8748), .A2(n10608), .ZN(n8733) );
  INV_X1 U11123 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n8730) );
  NAND2_X1 U11124 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n8736) );
  INV_X1 U11125 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n9909) );
  MUX2_X1 U11126 ( .A(n8736), .B(P3_IR_REG_31__SCAN_IN), .S(n9909), .Z(n8739)
         );
  INV_X1 U11127 ( .A(n8737), .ZN(n8738) );
  INV_X1 U11128 ( .A(SI_1_), .ZN(n9346) );
  XNOR2_X1 U11129 ( .A(n8741), .B(n8740), .ZN(n9347) );
  NAND2_X1 U11130 ( .A1(n12193), .A2(n12196), .ZN(n10045) );
  NAND2_X1 U11131 ( .A1(n9097), .A2(n10602), .ZN(n12191) );
  NAND2_X1 U11132 ( .A1(n10045), .A2(n12191), .ZN(n15121) );
  NAND2_X1 U11133 ( .A1(n9089), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8743) );
  NAND2_X1 U11134 ( .A1(n8753), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8742) );
  OR2_X1 U11135 ( .A1(n8737), .A2(n12929), .ZN(n8744) );
  XNOR2_X1 U11136 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8745) );
  XNOR2_X1 U11137 ( .A(n8746), .B(n8745), .ZN(n9335) );
  OR2_X1 U11138 ( .A1(n8756), .A2(SI_2_), .ZN(n8747) );
  NAND2_X1 U11139 ( .A1(n10051), .A2(n15129), .ZN(n12190) );
  NAND2_X1 U11140 ( .A1(n12203), .A2(n12190), .ZN(n12200) );
  INV_X1 U11141 ( .A(n12200), .ZN(n15120) );
  NAND2_X1 U11142 ( .A1(n15121), .A2(n15120), .ZN(n15119) );
  NAND2_X1 U11143 ( .A1(n15119), .A2(n12203), .ZN(n10301) );
  INV_X1 U11144 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10597) );
  OR2_X1 U11145 ( .A1(n8729), .A2(n10597), .ZN(n8752) );
  OR2_X1 U11146 ( .A1(n8748), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8751) );
  NAND2_X1 U11147 ( .A1(n8749), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8750) );
  INV_X1 U11148 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n8754) );
  OR2_X1 U11149 ( .A1(n9127), .A2(n8754), .ZN(n8755) );
  INV_X1 U11150 ( .A(n12556), .ZN(n15123) );
  OR2_X1 U11151 ( .A1(n12333), .A2(SI_3_), .ZN(n8763) );
  XNOR2_X1 U11152 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8757) );
  XNOR2_X1 U11153 ( .A(n8758), .B(n8757), .ZN(n9338) );
  OR2_X1 U11154 ( .A1(n8888), .A2(n9338), .ZN(n8762) );
  INV_X1 U11155 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8760) );
  NAND2_X1 U11156 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n6500), .ZN(n8759) );
  XNOR2_X1 U11157 ( .A(n8760), .B(n8759), .ZN(n14939) );
  INV_X1 U11158 ( .A(n14939), .ZN(n10546) );
  OR2_X1 U11159 ( .A1(n9834), .A2(n10546), .ZN(n8761) );
  NAND2_X1 U11160 ( .A1(n15123), .A2(n10595), .ZN(n12210) );
  INV_X1 U11161 ( .A(n10595), .ZN(n10462) );
  NAND2_X1 U11162 ( .A1(n12556), .A2(n10462), .ZN(n12204) );
  NAND2_X1 U11163 ( .A1(n12210), .A2(n12204), .ZN(n10303) );
  NAND2_X1 U11164 ( .A1(n10301), .A2(n12367), .ZN(n10300) );
  NAND2_X1 U11165 ( .A1(n10300), .A2(n12210), .ZN(n10440) );
  NAND2_X1 U11166 ( .A1(n9188), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8769) );
  INV_X1 U11167 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10543) );
  OR2_X1 U11168 ( .A1(n9127), .A2(n10543), .ZN(n8768) );
  NAND2_X1 U11169 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8764) );
  AND2_X1 U11170 ( .A1(n8778), .A2(n8764), .ZN(n10698) );
  OR2_X1 U11171 ( .A1(n6452), .A2(n10698), .ZN(n8767) );
  INV_X1 U11172 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n8765) );
  OR2_X1 U11173 ( .A1(n8731), .A2(n8765), .ZN(n8766) );
  OR2_X1 U11174 ( .A1(n12333), .A2(SI_4_), .ZN(n8777) );
  XNOR2_X1 U11175 ( .A(n8771), .B(n8770), .ZN(n9351) );
  OR2_X1 U11176 ( .A1(n8888), .A2(n9351), .ZN(n8776) );
  NAND2_X1 U11177 ( .A1(n8772), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8773) );
  MUX2_X1 U11178 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8773), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n8774) );
  AND2_X1 U11179 ( .A1(n8787), .A2(n8774), .ZN(n10542) );
  OR2_X1 U11180 ( .A1(n9834), .A2(n10542), .ZN(n8775) );
  NAND2_X1 U11181 ( .A1(n10710), .A2(n10494), .ZN(n12211) );
  INV_X1 U11182 ( .A(n10710), .ZN(n12555) );
  INV_X1 U11183 ( .A(n10494), .ZN(n10699) );
  NAND2_X1 U11184 ( .A1(n12555), .A2(n10699), .ZN(n12212) );
  NAND2_X1 U11185 ( .A1(n12211), .A2(n12212), .ZN(n10442) );
  NAND2_X1 U11186 ( .A1(n10440), .A2(n12363), .ZN(n10439) );
  NAND2_X1 U11187 ( .A1(n10439), .A2(n12211), .ZN(n10619) );
  NAND2_X1 U11188 ( .A1(n6445), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8783) );
  INV_X1 U11189 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10633) );
  OR2_X1 U11190 ( .A1(n12350), .A2(n10633), .ZN(n8782) );
  INV_X1 U11191 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10515) );
  OR2_X1 U11192 ( .A1(n9127), .A2(n10515), .ZN(n8781) );
  NAND2_X1 U11193 ( .A1(n8778), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8779) );
  AND2_X1 U11194 ( .A1(n8794), .A2(n8779), .ZN(n10715) );
  OR2_X1 U11195 ( .A1(n6452), .A2(n10715), .ZN(n8780) );
  OR2_X1 U11196 ( .A1(n12333), .A2(SI_5_), .ZN(n8793) );
  XNOR2_X1 U11197 ( .A(n8785), .B(n8784), .ZN(n9348) );
  OR2_X1 U11198 ( .A1(n8888), .A2(n9348), .ZN(n8792) );
  INV_X1 U11199 ( .A(n8786), .ZN(n8790) );
  NAND2_X1 U11200 ( .A1(n8787), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8788) );
  MUX2_X1 U11201 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8788), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n8789) );
  NAND2_X1 U11202 ( .A1(n8790), .A2(n8789), .ZN(n14977) );
  INV_X1 U11203 ( .A(n14977), .ZN(n10550) );
  OR2_X1 U11204 ( .A1(n6439), .A2(n10550), .ZN(n8791) );
  NAND2_X1 U11205 ( .A1(n10834), .A2(n10712), .ZN(n12216) );
  INV_X1 U11206 ( .A(n10834), .ZN(n12554) );
  INV_X1 U11207 ( .A(n10712), .ZN(n10809) );
  NAND2_X1 U11208 ( .A1(n12554), .A2(n10809), .ZN(n12215) );
  NAND2_X1 U11209 ( .A1(n10619), .A2(n12358), .ZN(n10618) );
  NAND2_X1 U11210 ( .A1(n10618), .A2(n12216), .ZN(n10830) );
  NAND2_X1 U11211 ( .A1(n9188), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8800) );
  INV_X1 U11212 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10541) );
  OR2_X1 U11213 ( .A1(n9127), .A2(n10541), .ZN(n8799) );
  NAND2_X1 U11214 ( .A1(n8794), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8795) );
  AND2_X1 U11215 ( .A1(n8808), .A2(n8795), .ZN(n10991) );
  OR2_X1 U11216 ( .A1(n6452), .A2(n10991), .ZN(n8798) );
  INV_X1 U11217 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n8796) );
  OR2_X1 U11218 ( .A1(n8731), .A2(n8796), .ZN(n8797) );
  OR2_X1 U11219 ( .A1(n8786), .A2(n12929), .ZN(n8801) );
  XNOR2_X1 U11220 ( .A(n8801), .B(n8816), .ZN(n14994) );
  INV_X1 U11221 ( .A(SI_6_), .ZN(n9333) );
  OR2_X1 U11222 ( .A1(n12333), .A2(n9333), .ZN(n8805) );
  XNOR2_X1 U11223 ( .A(n8803), .B(n8802), .ZN(n9334) );
  OR2_X1 U11224 ( .A1(n8888), .A2(n9334), .ZN(n8804) );
  OAI211_X1 U11225 ( .C1(n9834), .C2(n14994), .A(n8805), .B(n8804), .ZN(n10787) );
  NAND2_X1 U11226 ( .A1(n10921), .A2(n10787), .ZN(n12219) );
  INV_X1 U11227 ( .A(n10787), .ZN(n10992) );
  NAND2_X1 U11228 ( .A1(n12553), .A2(n10992), .ZN(n12220) );
  NAND2_X1 U11229 ( .A1(n12219), .A2(n12220), .ZN(n10832) );
  INV_X1 U11230 ( .A(n10832), .ZN(n12362) );
  NAND2_X1 U11231 ( .A1(n6445), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8813) );
  INV_X1 U11232 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n8806) );
  OR2_X1 U11233 ( .A1(n12350), .A2(n8806), .ZN(n8812) );
  INV_X1 U11234 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n8807) );
  OR2_X1 U11235 ( .A1(n9127), .A2(n8807), .ZN(n8811) );
  NAND2_X1 U11236 ( .A1(n8808), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8809) );
  AND2_X1 U11237 ( .A1(n8822), .A2(n8809), .ZN(n11120) );
  OR2_X1 U11238 ( .A1(n6452), .A2(n11120), .ZN(n8810) );
  OR2_X1 U11239 ( .A1(n12333), .A2(SI_7_), .ZN(n8821) );
  XNOR2_X1 U11240 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n8814) );
  XNOR2_X1 U11241 ( .A(n8815), .B(n8814), .ZN(n9343) );
  OR2_X1 U11242 ( .A1(n8888), .A2(n9343), .ZN(n8820) );
  NAND2_X1 U11243 ( .A1(n8786), .A2(n8816), .ZN(n8828) );
  NAND2_X1 U11244 ( .A1(n8828), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8818) );
  XNOR2_X1 U11245 ( .A(n8818), .B(n8817), .ZN(n10963) );
  INV_X1 U11246 ( .A(n10963), .ZN(n10951) );
  OR2_X1 U11247 ( .A1(n9834), .A2(n10951), .ZN(n8819) );
  NAND2_X1 U11248 ( .A1(n11081), .A2(n10924), .ZN(n12225) );
  INV_X1 U11249 ( .A(n11081), .ZN(n12552) );
  INV_X1 U11250 ( .A(n10924), .ZN(n11121) );
  NAND2_X1 U11251 ( .A1(n12552), .A2(n11121), .ZN(n12226) );
  NAND2_X1 U11252 ( .A1(n12225), .A2(n12226), .ZN(n12359) );
  INV_X1 U11253 ( .A(n12359), .ZN(n12222) );
  NAND2_X1 U11254 ( .A1(n9188), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8827) );
  NAND2_X1 U11255 ( .A1(n12346), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8826) );
  NAND2_X1 U11256 ( .A1(n6445), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8825) );
  NAND2_X1 U11257 ( .A1(n8822), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8823) );
  AND2_X1 U11258 ( .A1(n8853), .A2(n8823), .ZN(n11082) );
  OR2_X1 U11259 ( .A1(n6452), .A2(n11082), .ZN(n8824) );
  NAND4_X1 U11260 ( .A1(n8827), .A2(n8826), .A3(n8825), .A4(n8824), .ZN(n12551) );
  INV_X1 U11261 ( .A(n8861), .ZN(n8833) );
  NAND2_X1 U11262 ( .A1(n8829), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8831) );
  MUX2_X1 U11263 ( .A(n8831), .B(P3_IR_REG_31__SCAN_IN), .S(n8830), .Z(n8832)
         );
  XNOR2_X1 U11264 ( .A(n8835), .B(n8834), .ZN(n9342) );
  OR2_X1 U11265 ( .A1(n8888), .A2(n9342), .ZN(n8837) );
  INV_X1 U11266 ( .A(SI_8_), .ZN(n9341) );
  OR2_X1 U11267 ( .A1(n12333), .A2(n9341), .ZN(n8836) );
  OAI211_X1 U11268 ( .C1(n6439), .C2(n12609), .A(n8837), .B(n8836), .ZN(n12230) );
  XNOR2_X1 U11269 ( .A(n12551), .B(n12230), .ZN(n12365) );
  NAND2_X1 U11270 ( .A1(n9188), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8843) );
  INV_X1 U11271 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n12583) );
  OR2_X1 U11272 ( .A1(n9127), .A2(n12583), .ZN(n8842) );
  NAND2_X1 U11273 ( .A1(n8855), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8838) );
  AND2_X1 U11274 ( .A1(n8896), .A2(n8838), .ZN(n11262) );
  OR2_X1 U11275 ( .A1(n6452), .A2(n11262), .ZN(n8841) );
  INV_X1 U11276 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n8839) );
  OR2_X1 U11277 ( .A1(n8731), .A2(n8839), .ZN(n8840) );
  NAND2_X1 U11278 ( .A1(n8845), .A2(n8844), .ZN(n8847) );
  AND2_X1 U11279 ( .A1(n8847), .A2(n8846), .ZN(n9376) );
  OR2_X1 U11280 ( .A1(n8888), .A2(n9376), .ZN(n8851) );
  OR2_X1 U11281 ( .A1(n12333), .A2(SI_10_), .ZN(n8850) );
  INV_X1 U11282 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8862) );
  NAND2_X1 U11283 ( .A1(n8861), .A2(n8862), .ZN(n8889) );
  NAND2_X1 U11284 ( .A1(n8889), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8848) );
  XNOR2_X1 U11285 ( .A(n8848), .B(P3_IR_REG_10__SCAN_IN), .ZN(n12617) );
  OR2_X1 U11286 ( .A1(n6439), .A2(n12617), .ZN(n8849) );
  INV_X1 U11287 ( .A(n15153), .ZN(n11068) );
  NAND2_X1 U11288 ( .A1(n12550), .A2(n11068), .ZN(n12241) );
  INV_X1 U11289 ( .A(n12241), .ZN(n8871) );
  NAND2_X1 U11290 ( .A1(n9188), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8860) );
  INV_X1 U11291 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n8852) );
  OR2_X1 U11292 ( .A1(n9127), .A2(n8852), .ZN(n8859) );
  NAND2_X1 U11293 ( .A1(n8853), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n8854) );
  AND2_X1 U11294 ( .A1(n8855), .A2(n8854), .ZN(n11186) );
  OR2_X1 U11295 ( .A1(n6452), .A2(n11186), .ZN(n8858) );
  INV_X1 U11296 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n8856) );
  OR2_X1 U11297 ( .A1(n8731), .A2(n8856), .ZN(n8857) );
  OR2_X1 U11298 ( .A1(n8861), .A2(n12929), .ZN(n8863) );
  XNOR2_X1 U11299 ( .A(n8863), .B(n8862), .ZN(n15014) );
  INV_X1 U11300 ( .A(n15014), .ZN(n12563) );
  OR2_X1 U11301 ( .A1(n12333), .A2(SI_9_), .ZN(n8869) );
  NAND2_X1 U11302 ( .A1(n8865), .A2(n8864), .ZN(n8866) );
  AND2_X1 U11303 ( .A1(n8867), .A2(n8866), .ZN(n9356) );
  OR2_X1 U11304 ( .A1(n8888), .A2(n9356), .ZN(n8868) );
  OAI211_X1 U11305 ( .C1(n12563), .C2(n6439), .A(n8869), .B(n8868), .ZN(n15145) );
  INV_X1 U11306 ( .A(n15145), .ZN(n12235) );
  NAND2_X1 U11307 ( .A1(n11257), .A2(n12235), .ZN(n11061) );
  NAND2_X1 U11308 ( .A1(n11245), .A2(n15153), .ZN(n12240) );
  AND2_X1 U11309 ( .A1(n11061), .A2(n12240), .ZN(n8870) );
  OR2_X1 U11310 ( .A1(n8871), .A2(n8870), .ZN(n8876) );
  INV_X1 U11311 ( .A(n8876), .ZN(n8873) );
  NAND2_X1 U11312 ( .A1(n12234), .A2(n15145), .ZN(n11060) );
  AND2_X1 U11313 ( .A1(n11060), .A2(n12241), .ZN(n8872) );
  AND2_X1 U11314 ( .A1(n12365), .A2(n8875), .ZN(n8874) );
  INV_X1 U11315 ( .A(n8875), .ZN(n8878) );
  NAND2_X1 U11316 ( .A1(n11184), .A2(n12230), .ZN(n11059) );
  AND2_X1 U11317 ( .A1(n11059), .A2(n8876), .ZN(n8877) );
  OR2_X1 U11318 ( .A1(n8878), .A2(n8877), .ZN(n8879) );
  NAND2_X1 U11319 ( .A1(n8880), .A2(n8879), .ZN(n11246) );
  INV_X1 U11320 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n8881) );
  OR2_X1 U11321 ( .A1(n9127), .A2(n8881), .ZN(n8885) );
  NAND2_X1 U11322 ( .A1(n6445), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8884) );
  XNOR2_X1 U11323 ( .A(n8896), .B(n11430), .ZN(n11433) );
  OR2_X1 U11324 ( .A1(n6452), .A2(n11433), .ZN(n8883) );
  INV_X1 U11325 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n12602) );
  OR2_X1 U11326 ( .A1(n12350), .A2(n12602), .ZN(n8882) );
  XNOR2_X1 U11327 ( .A(n9454), .B(P2_DATAO_REG_11__SCAN_IN), .ZN(n8886) );
  XNOR2_X1 U11328 ( .A(n8887), .B(n8886), .ZN(n9382) );
  OR2_X1 U11329 ( .A1(n9382), .A2(n8888), .ZN(n8894) );
  OR2_X1 U11330 ( .A1(n12333), .A2(SI_11_), .ZN(n8893) );
  OAI21_X1 U11331 ( .B1(n8889), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8891) );
  INV_X1 U11332 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8890) );
  XNOR2_X1 U11333 ( .A(n8891), .B(n8890), .ZN(n15049) );
  OR2_X1 U11334 ( .A1(n9834), .A2(n12605), .ZN(n8892) );
  XNOR2_X1 U11335 ( .A(n12549), .B(n12246), .ZN(n12374) );
  NAND2_X1 U11336 ( .A1(n7425), .A2(n12246), .ZN(n12247) );
  NAND2_X1 U11337 ( .A1(n12346), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8901) );
  INV_X1 U11338 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n8895) );
  OR2_X1 U11339 ( .A1(n8731), .A2(n8895), .ZN(n8900) );
  OAI21_X1 U11340 ( .B1(n8896), .B2(P3_REG3_REG_11__SCAN_IN), .A(
        P3_REG3_REG_12__SCAN_IN), .ZN(n8897) );
  AND2_X1 U11341 ( .A1(n8917), .A2(n8897), .ZN(n11488) );
  OR2_X1 U11342 ( .A1(n6452), .A2(n11488), .ZN(n8899) );
  INV_X1 U11343 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12620) );
  OR2_X1 U11344 ( .A1(n12350), .A2(n12620), .ZN(n8898) );
  INV_X1 U11345 ( .A(n9834), .ZN(n8992) );
  NOR2_X1 U11346 ( .A1(n8902), .A2(n12929), .ZN(n8903) );
  MUX2_X1 U11347 ( .A(n12929), .B(n8903), .S(P3_IR_REG_12__SCAN_IN), .Z(n8906)
         );
  INV_X1 U11348 ( .A(n8904), .ZN(n8905) );
  INV_X1 U11349 ( .A(n15068), .ZN(n12623) );
  AOI22_X1 U11350 ( .A1(n8993), .A2(SI_12_), .B1(n8992), .B2(n12623), .ZN(
        n8910) );
  XNOR2_X1 U11351 ( .A(n8908), .B(n8907), .ZN(n9393) );
  NAND2_X1 U11352 ( .A1(n9393), .A2(n12343), .ZN(n8909) );
  NAND2_X1 U11353 ( .A1(n8910), .A2(n8909), .ZN(n14487) );
  NAND2_X1 U11354 ( .A1(n11423), .A2(n14487), .ZN(n12250) );
  INV_X1 U11355 ( .A(n14487), .ZN(n11224) );
  NAND2_X1 U11356 ( .A1(n12548), .A2(n11224), .ZN(n12251) );
  NAND2_X1 U11357 ( .A1(n12250), .A2(n12251), .ZN(n12370) );
  XNOR2_X1 U11358 ( .A(n8911), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n9411) );
  NAND2_X1 U11359 ( .A1(n9411), .A2(n12343), .ZN(n8915) );
  NAND2_X1 U11360 ( .A1(n8904), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8913) );
  INV_X1 U11361 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8912) );
  XNOR2_X1 U11362 ( .A(n8913), .B(n8912), .ZN(n15084) );
  AOI22_X1 U11363 ( .A1(n8993), .A2(n9412), .B1(n8992), .B2(n15084), .ZN(n8914) );
  NAND2_X1 U11364 ( .A1(n8915), .A2(n8914), .ZN(n14482) );
  INV_X1 U11365 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n8916) );
  OR2_X1 U11366 ( .A1(n9127), .A2(n8916), .ZN(n8922) );
  NAND2_X1 U11367 ( .A1(n6445), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8921) );
  NAND2_X1 U11368 ( .A1(n8917), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8918) );
  AND2_X1 U11369 ( .A1(n8930), .A2(n8918), .ZN(n11421) );
  OR2_X1 U11370 ( .A1(n6452), .A2(n11421), .ZN(n8920) );
  INV_X1 U11371 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12626) );
  OR2_X1 U11372 ( .A1(n12350), .A2(n12626), .ZN(n8919) );
  NAND4_X1 U11373 ( .A1(n8922), .A2(n8921), .A3(n8920), .A4(n8919), .ZN(n11485) );
  OR2_X1 U11374 ( .A1(n14482), .A2(n11485), .ZN(n12255) );
  INV_X1 U11375 ( .A(n12255), .ZN(n8923) );
  NAND2_X1 U11376 ( .A1(n14482), .A2(n11485), .ZN(n12256) );
  NAND2_X1 U11377 ( .A1(n8924), .A2(n12256), .ZN(n11438) );
  XNOR2_X1 U11378 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8925) );
  XNOR2_X1 U11379 ( .A(n8926), .B(n8925), .ZN(n9426) );
  NAND2_X1 U11380 ( .A1(n9426), .A2(n12343), .ZN(n8929) );
  NAND2_X1 U11381 ( .A1(n7444), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8927) );
  XNOR2_X1 U11382 ( .A(n8927), .B(n7108), .ZN(n15100) );
  AOI22_X1 U11383 ( .A1(n8993), .A2(n14351), .B1(n8992), .B2(n15100), .ZN(
        n8928) );
  NAND2_X1 U11384 ( .A1(n8929), .A2(n8928), .ZN(n14477) );
  NAND2_X1 U11385 ( .A1(n12346), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8935) );
  NAND2_X1 U11386 ( .A1(n9188), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8934) );
  NAND2_X1 U11387 ( .A1(n6445), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8933) );
  NAND2_X1 U11388 ( .A1(n8930), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8931) );
  AND2_X1 U11389 ( .A1(n8946), .A2(n8931), .ZN(n11474) );
  OR2_X1 U11390 ( .A1(n6452), .A2(n11474), .ZN(n8932) );
  NAND4_X1 U11391 ( .A1(n8935), .A2(n8934), .A3(n8933), .A4(n8932), .ZN(n12547) );
  NAND2_X1 U11392 ( .A1(n14477), .A2(n12547), .ZN(n12260) );
  INV_X1 U11393 ( .A(n12260), .ZN(n8936) );
  OR2_X1 U11394 ( .A1(n14477), .A2(n12547), .ZN(n12262) );
  NAND2_X1 U11395 ( .A1(n8938), .A2(n8937), .ZN(n8939) );
  NAND2_X1 U11396 ( .A1(n8940), .A2(n8939), .ZN(n9567) );
  NAND2_X1 U11397 ( .A1(n9567), .A2(n12343), .ZN(n8945) );
  NAND2_X1 U11398 ( .A1(n8941), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8943) );
  XNOR2_X1 U11399 ( .A(n8943), .B(n8942), .ZN(n14408) );
  AOI22_X1 U11400 ( .A1(n8993), .A2(n9568), .B1(n8992), .B2(n14408), .ZN(n8944) );
  INV_X1 U11401 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n14335) );
  OR2_X1 U11402 ( .A1(n9127), .A2(n14335), .ZN(n8951) );
  INV_X1 U11403 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n14244) );
  OR2_X1 U11404 ( .A1(n6440), .A2(n14244), .ZN(n8950) );
  NAND2_X1 U11405 ( .A1(n8946), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8947) );
  AND2_X1 U11406 ( .A1(n8959), .A2(n8947), .ZN(n11466) );
  OR2_X1 U11407 ( .A1(n6452), .A2(n11466), .ZN(n8949) );
  INV_X1 U11408 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14405) );
  OR2_X1 U11409 ( .A1(n12350), .A2(n14405), .ZN(n8948) );
  NAND4_X1 U11410 ( .A1(n8951), .A2(n8950), .A3(n8949), .A4(n8948), .ZN(n12546) );
  NAND2_X1 U11411 ( .A1(n12925), .A2(n12546), .ZN(n12269) );
  OAI21_X1 U11412 ( .B1(n8954), .B2(n8953), .A(n8952), .ZN(n9646) );
  OR2_X1 U11413 ( .A1(n9646), .A2(n8888), .ZN(n8958) );
  OR2_X1 U11414 ( .A1(n8955), .A2(n12929), .ZN(n8956) );
  XNOR2_X1 U11415 ( .A(n8956), .B(P3_IR_REG_16__SCAN_IN), .ZN(n14421) );
  AOI22_X1 U11416 ( .A1(n8993), .A2(SI_16_), .B1(n8992), .B2(n14421), .ZN(
        n8957) );
  NAND2_X1 U11417 ( .A1(n9188), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8964) );
  INV_X1 U11418 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12871) );
  OR2_X1 U11419 ( .A1(n9127), .A2(n12871), .ZN(n8963) );
  NAND2_X1 U11420 ( .A1(n6445), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8962) );
  NAND2_X1 U11421 ( .A1(n8959), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8960) );
  AND2_X1 U11422 ( .A1(n8972), .A2(n8960), .ZN(n12817) );
  OR2_X1 U11423 ( .A1(n6452), .A2(n12817), .ZN(n8961) );
  NAND4_X1 U11424 ( .A1(n8964), .A2(n8963), .A3(n8962), .A4(n8961), .ZN(n12545) );
  NAND2_X1 U11425 ( .A1(n12922), .A2(n12545), .ZN(n12270) );
  NAND2_X1 U11426 ( .A1(n12463), .A2(n12798), .ZN(n12271) );
  NAND2_X1 U11427 ( .A1(n12270), .A2(n12271), .ZN(n12808) );
  NAND2_X1 U11428 ( .A1(n12814), .A2(n7434), .ZN(n12813) );
  XNOR2_X1 U11429 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .ZN(n8965) );
  XNOR2_X1 U11430 ( .A(n8966), .B(n8965), .ZN(n9756) );
  NAND2_X1 U11431 ( .A1(n9756), .A2(n12343), .ZN(n8971) );
  NAND2_X1 U11432 ( .A1(n8967), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8969) );
  INV_X1 U11433 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8968) );
  XNOR2_X1 U11434 ( .A(n8969), .B(n8968), .ZN(n12643) );
  AOI22_X1 U11435 ( .A1(n8993), .A2(n9757), .B1(n8992), .B2(n12643), .ZN(n8970) );
  INV_X1 U11436 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12867) );
  OR2_X1 U11437 ( .A1(n9127), .A2(n12867), .ZN(n8976) );
  NAND2_X1 U11438 ( .A1(n6445), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8975) );
  XNOR2_X1 U11439 ( .A(n8972), .B(n12469), .ZN(n12803) );
  OR2_X1 U11440 ( .A1(n6452), .A2(n12803), .ZN(n8974) );
  INV_X1 U11441 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14448) );
  OR2_X1 U11442 ( .A1(n12350), .A2(n14448), .ZN(n8973) );
  NAND4_X1 U11443 ( .A1(n8976), .A2(n8975), .A3(n8974), .A4(n8973), .ZN(n12544) );
  NAND2_X1 U11444 ( .A1(n12918), .A2(n12544), .ZN(n12276) );
  NAND2_X1 U11445 ( .A1(n12802), .A2(n12801), .ZN(n8977) );
  NAND2_X1 U11446 ( .A1(n8977), .A2(n12275), .ZN(n12788) );
  XNOR2_X1 U11447 ( .A(n8979), .B(n8978), .ZN(n9966) );
  NAND2_X1 U11448 ( .A1(n9966), .A2(n12343), .ZN(n8982) );
  NAND2_X1 U11449 ( .A1(n6479), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8980) );
  XNOR2_X1 U11450 ( .A(n8980), .B(P3_IR_REG_18__SCAN_IN), .ZN(n14454) );
  AOI22_X1 U11451 ( .A1(n8993), .A2(SI_18_), .B1(n8992), .B2(n14454), .ZN(
        n8981) );
  NAND2_X1 U11452 ( .A1(n8982), .A2(n8981), .ZN(n12139) );
  NAND2_X1 U11453 ( .A1(n12346), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8989) );
  INV_X1 U11454 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12791) );
  OR2_X1 U11455 ( .A1(n12350), .A2(n12791), .ZN(n8988) );
  INV_X1 U11456 ( .A(n8983), .ZN(n8984) );
  NAND2_X1 U11457 ( .A1(n8984), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8985) );
  AND2_X1 U11458 ( .A1(n8996), .A2(n8985), .ZN(n12790) );
  OR2_X1 U11459 ( .A1(n6452), .A2(n12790), .ZN(n8987) );
  INV_X1 U11460 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12912) );
  OR2_X1 U11461 ( .A1(n8731), .A2(n12912), .ZN(n8986) );
  OR2_X1 U11462 ( .A1(n12139), .A2(n12800), .ZN(n12279) );
  NAND2_X1 U11463 ( .A1(n12139), .A2(n12800), .ZN(n12283) );
  AOI22_X1 U11464 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(
        P1_DATAO_REG_19__SCAN_IN), .B1(n10944), .B2(n10942), .ZN(n8990) );
  XNOR2_X1 U11465 ( .A(n8991), .B(n8990), .ZN(n10011) );
  NAND2_X1 U11466 ( .A1(n10011), .A2(n12343), .ZN(n8995) );
  AOI22_X1 U11467 ( .A1(n8993), .A2(SI_19_), .B1(n8992), .B2(n12404), .ZN(
        n8994) );
  NAND2_X1 U11468 ( .A1(n6445), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9001) );
  INV_X1 U11469 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12859) );
  OR2_X1 U11470 ( .A1(n9127), .A2(n12859), .ZN(n9000) );
  NAND2_X1 U11471 ( .A1(n8996), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8997) );
  AND2_X1 U11472 ( .A1(n9007), .A2(n8997), .ZN(n12775) );
  OR2_X1 U11473 ( .A1(n12775), .A2(n6452), .ZN(n8999) );
  INV_X1 U11474 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12776) );
  OR2_X1 U11475 ( .A1(n12350), .A2(n12776), .ZN(n8998) );
  INV_X1 U11476 ( .A(n12288), .ZN(n9002) );
  NAND2_X1 U11477 ( .A1(n12439), .A2(n12785), .ZN(n12287) );
  XNOR2_X1 U11478 ( .A(n9004), .B(n9003), .ZN(n10195) );
  NAND2_X1 U11479 ( .A1(n10195), .A2(n12343), .ZN(n9006) );
  OR2_X1 U11480 ( .A1(n12333), .A2(n10197), .ZN(n9005) );
  NAND2_X1 U11481 ( .A1(n9007), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9008) );
  NAND2_X1 U11482 ( .A1(n9021), .A2(n9008), .ZN(n12761) );
  NAND2_X1 U11483 ( .A1(n9089), .A2(n12761), .ZN(n9013) );
  INV_X1 U11484 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12855) );
  OR2_X1 U11485 ( .A1(n9127), .A2(n12855), .ZN(n9012) );
  INV_X1 U11486 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12904) );
  OR2_X1 U11487 ( .A1(n6440), .A2(n12904), .ZN(n9011) );
  INV_X1 U11488 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n9009) );
  OR2_X1 U11489 ( .A1(n12350), .A2(n9009), .ZN(n9010) );
  NAND2_X1 U11490 ( .A1(n12482), .A2(n12746), .ZN(n12293) );
  NAND2_X1 U11491 ( .A1(n12292), .A2(n12293), .ZN(n12760) );
  XNOR2_X1 U11492 ( .A(n9016), .B(n9015), .ZN(n10411) );
  NAND2_X1 U11493 ( .A1(n10411), .A2(n12343), .ZN(n9018) );
  INV_X1 U11494 ( .A(SI_21_), .ZN(n10413) );
  OR2_X1 U11495 ( .A1(n12333), .A2(n10413), .ZN(n9017) );
  NAND2_X1 U11496 ( .A1(n9188), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n9020) );
  INV_X1 U11497 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n14237) );
  OR2_X1 U11498 ( .A1(n9127), .A2(n14237), .ZN(n9019) );
  AND2_X1 U11499 ( .A1(n9020), .A2(n9019), .ZN(n9025) );
  NAND2_X1 U11500 ( .A1(n9021), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n9022) );
  NAND2_X1 U11501 ( .A1(n9032), .A2(n9022), .ZN(n12751) );
  NAND2_X1 U11502 ( .A1(n12751), .A2(n9089), .ZN(n9024) );
  NAND2_X1 U11503 ( .A1(n6445), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n9023) );
  NAND2_X1 U11504 ( .A1(n12750), .A2(n12758), .ZN(n12294) );
  NAND2_X1 U11505 ( .A1(n12749), .A2(n12294), .ZN(n9026) );
  XNOR2_X1 U11506 ( .A(n9028), .B(n9027), .ZN(n10459) );
  NAND2_X1 U11507 ( .A1(n10459), .A2(n12343), .ZN(n9031) );
  OR2_X1 U11508 ( .A1(n12333), .A2(n9029), .ZN(n9030) );
  INV_X1 U11509 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n14334) );
  NAND2_X1 U11510 ( .A1(n9032), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9033) );
  NAND2_X1 U11511 ( .A1(n9040), .A2(n9033), .ZN(n12737) );
  NAND2_X1 U11512 ( .A1(n12737), .A2(n9089), .ZN(n9035) );
  AOI22_X1 U11513 ( .A1(n9188), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n12346), 
        .B2(P3_REG1_REG_22__SCAN_IN), .ZN(n9034) );
  OAI211_X1 U11514 ( .C1(n8731), .C2(n14334), .A(n9035), .B(n9034), .ZN(n12540) );
  NAND2_X1 U11515 ( .A1(n12736), .A2(n12747), .ZN(n12306) );
  XNOR2_X1 U11516 ( .A(n9037), .B(n9036), .ZN(n10629) );
  NAND2_X1 U11517 ( .A1(n10629), .A2(n12343), .ZN(n9039) );
  OR2_X1 U11518 ( .A1(n12333), .A2(n10631), .ZN(n9038) );
  NAND2_X1 U11519 ( .A1(n9040), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9041) );
  NAND2_X1 U11520 ( .A1(n9049), .A2(n9041), .ZN(n12726) );
  NAND2_X1 U11521 ( .A1(n12726), .A2(n9089), .ZN(n9044) );
  AOI22_X1 U11522 ( .A1(n9188), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n12346), 
        .B2(P3_REG1_REG_23__SCAN_IN), .ZN(n9043) );
  INV_X1 U11523 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n14266) );
  OR2_X1 U11524 ( .A1(n8731), .A2(n14266), .ZN(n9042) );
  NAND2_X1 U11525 ( .A1(n12725), .A2(n12733), .ZN(n12304) );
  INV_X1 U11526 ( .A(n12724), .ZN(n12382) );
  XNOR2_X1 U11527 ( .A(n9046), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n10927) );
  NAND2_X1 U11528 ( .A1(n10927), .A2(n12343), .ZN(n9048) );
  NAND2_X1 U11529 ( .A1(n9049), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9050) );
  NAND2_X1 U11530 ( .A1(n9061), .A2(n9050), .ZN(n12713) );
  INV_X1 U11531 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n9053) );
  NAND2_X1 U11532 ( .A1(n12346), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9052) );
  NAND2_X1 U11533 ( .A1(n6445), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n9051) );
  OAI211_X1 U11534 ( .C1(n9053), .C2(n12350), .A(n9052), .B(n9051), .ZN(n9054)
         );
  AOI21_X1 U11535 ( .B1(n12713), .B2(n9089), .A(n9054), .ZN(n12694) );
  XNOR2_X1 U11536 ( .A(n12712), .B(n12694), .ZN(n12705) );
  NAND2_X1 U11537 ( .A1(n12712), .A2(n12694), .ZN(n12310) );
  NAND2_X1 U11538 ( .A1(n9056), .A2(n9055), .ZN(n9057) );
  NAND2_X1 U11539 ( .A1(n9058), .A2(n9057), .ZN(n11831) );
  NAND2_X1 U11540 ( .A1(n9061), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9062) );
  NAND2_X1 U11541 ( .A1(n9072), .A2(n9062), .ZN(n12699) );
  NAND2_X1 U11542 ( .A1(n12699), .A2(n9089), .ZN(n9067) );
  INV_X1 U11543 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n14293) );
  NAND2_X1 U11544 ( .A1(n9188), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9064) );
  NAND2_X1 U11545 ( .A1(n6445), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n9063) );
  OAI211_X1 U11546 ( .C1(n9127), .C2(n14293), .A(n9064), .B(n9063), .ZN(n9065)
         );
  INV_X1 U11547 ( .A(n9065), .ZN(n9066) );
  NAND2_X1 U11548 ( .A1(n12698), .A2(n12677), .ZN(n12680) );
  XNOR2_X1 U11549 ( .A(n9069), .B(n9068), .ZN(n11194) );
  NAND2_X1 U11550 ( .A1(n11194), .A2(n12343), .ZN(n9071) );
  OR2_X1 U11551 ( .A1(n12333), .A2(n11195), .ZN(n9070) );
  NAND2_X1 U11552 ( .A1(n9072), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9073) );
  NAND2_X1 U11553 ( .A1(n9086), .A2(n9073), .ZN(n12683) );
  NAND2_X1 U11554 ( .A1(n12683), .A2(n9089), .ZN(n9079) );
  INV_X1 U11555 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n9076) );
  NAND2_X1 U11556 ( .A1(n6445), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n9075) );
  NAND2_X1 U11557 ( .A1(n12346), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9074) );
  OAI211_X1 U11558 ( .C1(n12350), .C2(n9076), .A(n9075), .B(n9074), .ZN(n9077)
         );
  INV_X1 U11559 ( .A(n9077), .ZN(n9078) );
  NAND2_X1 U11560 ( .A1(n12516), .A2(n12453), .ZN(n12319) );
  NAND2_X1 U11561 ( .A1(n12318), .A2(n12319), .ZN(n12673) );
  INV_X1 U11562 ( .A(n12680), .ZN(n9080) );
  NOR2_X1 U11563 ( .A1(n12673), .A2(n9080), .ZN(n9081) );
  NAND2_X1 U11564 ( .A1(n12695), .A2(n9081), .ZN(n12678) );
  XNOR2_X1 U11565 ( .A(n9083), .B(n9082), .ZN(n11331) );
  NAND2_X1 U11566 ( .A1(n11331), .A2(n12343), .ZN(n9085) );
  NAND2_X1 U11567 ( .A1(n9086), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9087) );
  NAND2_X1 U11568 ( .A1(n9088), .A2(n9087), .ZN(n11517) );
  NAND2_X1 U11569 ( .A1(n11517), .A2(n9089), .ZN(n9094) );
  INV_X1 U11570 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n11518) );
  NAND2_X1 U11571 ( .A1(n12346), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n9091) );
  NAND2_X1 U11572 ( .A1(n6445), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n9090) );
  OAI211_X1 U11573 ( .C1(n12350), .C2(n11518), .A(n9091), .B(n9090), .ZN(n9092) );
  INV_X1 U11574 ( .A(n9092), .ZN(n9093) );
  NAND2_X1 U11575 ( .A1(n12170), .A2(n12676), .ZN(n9197) );
  NAND2_X1 U11576 ( .A1(n11509), .A2(n9197), .ZN(n9096) );
  XOR2_X1 U11577 ( .A(n12321), .B(n9096), .Z(n12667) );
  INV_X1 U11578 ( .A(n12758), .ZN(n12541) );
  INV_X1 U11579 ( .A(n12139), .ZN(n12914) );
  NAND2_X1 U11580 ( .A1(n12559), .A2(n9882), .ZN(n10604) );
  NAND2_X1 U11581 ( .A1(n10043), .A2(n10604), .ZN(n9099) );
  NAND2_X1 U11582 ( .A1(n9097), .A2(n10052), .ZN(n9098) );
  NAND2_X1 U11583 ( .A1(n9099), .A2(n9098), .ZN(n15118) );
  INV_X1 U11584 ( .A(n15129), .ZN(n10101) );
  NAND2_X1 U11585 ( .A1(n10304), .A2(n10303), .ZN(n10302) );
  NAND2_X1 U11586 ( .A1(n12556), .A2(n10595), .ZN(n9100) );
  NAND2_X1 U11587 ( .A1(n12555), .A2(n10494), .ZN(n9101) );
  NAND2_X1 U11588 ( .A1(n10834), .A2(n10809), .ZN(n9102) );
  AND2_X2 U11589 ( .A1(n10622), .A2(n9102), .ZN(n10833) );
  NAND2_X1 U11590 ( .A1(n12553), .A2(n10787), .ZN(n9103) );
  INV_X1 U11591 ( .A(n12230), .ZN(n12229) );
  NAND2_X1 U11592 ( .A1(n11184), .A2(n12229), .ZN(n9105) );
  AND2_X1 U11593 ( .A1(n12359), .A2(n9105), .ZN(n9104) );
  INV_X1 U11594 ( .A(n9105), .ZN(n9107) );
  INV_X1 U11595 ( .A(n12365), .ZN(n9106) );
  NAND2_X1 U11596 ( .A1(n12552), .A2(n10924), .ZN(n11075) );
  AND2_X1 U11597 ( .A1(n9106), .A2(n11075), .ZN(n11076) );
  OR2_X1 U11598 ( .A1(n9107), .A2(n11076), .ZN(n9108) );
  NAND2_X1 U11599 ( .A1(n11257), .A2(n15145), .ZN(n9109) );
  NAND2_X1 U11600 ( .A1(n12234), .A2(n12235), .ZN(n12237) );
  NAND2_X1 U11601 ( .A1(n12240), .A2(n12241), .ZN(n12243) );
  NAND2_X1 U11602 ( .A1(n12550), .A2(n15153), .ZN(n9110) );
  INV_X1 U11603 ( .A(n11485), .ZN(n11441) );
  NAND2_X1 U11604 ( .A1(n12262), .A2(n12260), .ZN(n12376) );
  INV_X1 U11605 ( .A(n14477), .ZN(n11444) );
  INV_X1 U11606 ( .A(n12544), .ZN(n12812) );
  NAND2_X1 U11607 ( .A1(n12288), .A2(n12287), .ZN(n12774) );
  OAI21_X2 U11608 ( .B1(n12785), .B2(n12910), .A(n12767), .ZN(n12756) );
  NAND2_X1 U11609 ( .A1(n12295), .A2(n12294), .ZN(n12748) );
  NAND2_X1 U11610 ( .A1(n12736), .A2(n12540), .ZN(n9111) );
  NAND2_X1 U11611 ( .A1(n12719), .A2(n12724), .ZN(n12718) );
  INV_X1 U11612 ( .A(n12733), .ZN(n12539) );
  NAND2_X1 U11613 ( .A1(n12725), .A2(n12539), .ZN(n9112) );
  NAND2_X1 U11614 ( .A1(n12718), .A2(n9112), .ZN(n12706) );
  NAND2_X1 U11615 ( .A1(n12706), .A2(n12705), .ZN(n12704) );
  NAND2_X1 U11616 ( .A1(n12712), .A2(n12720), .ZN(n9113) );
  NAND2_X1 U11617 ( .A1(n12704), .A2(n9113), .ZN(n12690) );
  NAND2_X1 U11618 ( .A1(n12690), .A2(n12689), .ZN(n12688) );
  NAND2_X1 U11619 ( .A1(n12698), .A2(n12707), .ZN(n9114) );
  NAND2_X1 U11620 ( .A1(n12688), .A2(n9114), .ZN(n12674) );
  NAND2_X1 U11621 ( .A1(n12884), .A2(n12453), .ZN(n9115) );
  NAND2_X1 U11622 ( .A1(n12674), .A2(n9115), .ZN(n9117) );
  NAND2_X1 U11623 ( .A1(n12516), .A2(n12691), .ZN(n9116) );
  NAND2_X1 U11624 ( .A1(n9117), .A2(n9116), .ZN(n9118) );
  INV_X1 U11625 ( .A(n11504), .ZN(n9120) );
  NOR2_X1 U11626 ( .A1(n12170), .A2(n12538), .ZN(n9121) );
  OAI21_X1 U11627 ( .B1(n9120), .B2(n9121), .A(n12321), .ZN(n9123) );
  NAND2_X1 U11628 ( .A1(n12404), .A2(n12415), .ZN(n9166) );
  NAND2_X1 U11629 ( .A1(n12195), .A2(n9165), .ZN(n12406) );
  NOR2_X1 U11630 ( .A1(n12321), .A2(n9121), .ZN(n9122) );
  OR2_X1 U11631 ( .A1(n12420), .A2(n6452), .ZN(n12353) );
  INV_X1 U11632 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9126) );
  NAND2_X1 U11633 ( .A1(n9188), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9125) );
  NAND2_X1 U11634 ( .A1(n6445), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9124) );
  OAI211_X1 U11635 ( .C1(n9127), .C2(n9126), .A(n9125), .B(n9124), .ZN(n9128)
         );
  INV_X1 U11636 ( .A(n9128), .ZN(n9129) );
  INV_X1 U11637 ( .A(n9130), .ZN(n12412) );
  NAND2_X1 U11638 ( .A1(n12412), .A2(n10514), .ZN(n9841) );
  NAND2_X1 U11639 ( .A1(n9834), .A2(n9841), .ZN(n10049) );
  OAI22_X1 U11640 ( .A1(n12185), .A2(n15122), .B1(n12676), .B2(n12799), .ZN(
        n9131) );
  INV_X1 U11641 ( .A(n9131), .ZN(n9132) );
  OAI21_X1 U11642 ( .B1(n14483), .B2(n12667), .A(n12672), .ZN(n9174) );
  NAND2_X1 U11643 ( .A1(n9167), .A2(n12327), .ZN(n9889) );
  NAND2_X1 U11644 ( .A1(n9133), .A2(n12317), .ZN(n10583) );
  AND2_X1 U11645 ( .A1(n9889), .A2(n10583), .ZN(n10585) );
  OAI22_X1 U11646 ( .A1(n12404), .A2(n9134), .B1(n9165), .B2(n15144), .ZN(
        n9135) );
  AOI21_X1 U11647 ( .B1(n9135), .B2(n9167), .A(n12327), .ZN(n9145) );
  NAND2_X1 U11648 ( .A1(n6547), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9136) );
  MUX2_X1 U11649 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9136), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n9138) );
  NAND2_X1 U11650 ( .A1(n9138), .A2(n9137), .ZN(n10930) );
  XNOR2_X1 U11651 ( .A(n10930), .B(P3_B_REG_SCAN_IN), .ZN(n9141) );
  NAND2_X1 U11652 ( .A1(n9137), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9139) );
  MUX2_X1 U11653 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9139), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n9140) );
  NAND2_X1 U11654 ( .A1(n9140), .A2(n6482), .ZN(n11829) );
  NAND2_X1 U11655 ( .A1(n9141), .A2(n11829), .ZN(n9143) );
  NAND2_X1 U11656 ( .A1(n6482), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9142) );
  INV_X1 U11657 ( .A(n9159), .ZN(n11197) );
  NAND2_X1 U11658 ( .A1(n11197), .A2(n11829), .ZN(n9144) );
  MUX2_X1 U11659 ( .A(n10585), .B(n9145), .S(n10584), .Z(n9164) );
  NAND2_X1 U11660 ( .A1(n11197), .A2(n10930), .ZN(n9422) );
  NOR2_X1 U11661 ( .A1(P3_D_REG_22__SCAN_IN), .A2(P3_D_REG_7__SCAN_IN), .ZN(
        n9149) );
  NOR4_X1 U11662 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_2__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_17__SCAN_IN), .ZN(n9148) );
  NOR4_X1 U11663 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_10__SCAN_IN), .ZN(n9147) );
  NOR4_X1 U11664 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n9146) );
  NAND4_X1 U11665 ( .A1(n9149), .A2(n9148), .A3(n9147), .A4(n9146), .ZN(n9155)
         );
  NOR4_X1 U11666 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n9153) );
  NOR4_X1 U11667 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_11__SCAN_IN), .ZN(n9152) );
  NOR4_X1 U11668 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_8__SCAN_IN), .ZN(n9151) );
  NOR4_X1 U11669 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n9150) );
  NAND4_X1 U11670 ( .A1(n9153), .A2(n9152), .A3(n9151), .A4(n9150), .ZN(n9154)
         );
  NOR2_X1 U11671 ( .A1(n9155), .A2(n9154), .ZN(n9156) );
  INV_X1 U11672 ( .A(n10930), .ZN(n9158) );
  INV_X1 U11673 ( .A(n11829), .ZN(n9157) );
  INV_X1 U11674 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9161) );
  NOR2_X1 U11675 ( .A1(n9170), .A2(n9880), .ZN(n9163) );
  NAND2_X1 U11676 ( .A1(n10584), .A2(n10040), .ZN(n9171) );
  INV_X1 U11677 ( .A(n15144), .ZN(n15152) );
  NAND2_X1 U11678 ( .A1(n10414), .A2(n9165), .ZN(n12392) );
  OR2_X1 U11679 ( .A1(n9166), .A2(n12392), .ZN(n9884) );
  NOR2_X1 U11680 ( .A1(n9167), .A2(n12317), .ZN(n10107) );
  INV_X1 U11681 ( .A(n9880), .ZN(n9877) );
  NAND2_X1 U11682 ( .A1(n10107), .A2(n9877), .ZN(n9895) );
  OAI21_X1 U11683 ( .B1(n9884), .B2(n9880), .A(n9895), .ZN(n9169) );
  NOR2_X1 U11684 ( .A1(n9168), .A2(n9170), .ZN(n9893) );
  NAND2_X1 U11685 ( .A1(n9169), .A2(n9893), .ZN(n9173) );
  NAND3_X1 U11686 ( .A1(n9896), .A2(n9877), .A3(n9883), .ZN(n9172) );
  INV_X1 U11687 ( .A(n9175), .ZN(n9176) );
  NAND2_X1 U11688 ( .A1(n9176), .A2(n7446), .ZN(P3_U3455) );
  INV_X1 U11689 ( .A(n9179), .ZN(n9180) );
  NAND2_X1 U11690 ( .A1(n9181), .A2(n9180), .ZN(n9183) );
  AOI22_X1 U11691 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n13545), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n14369), .ZN(n9184) );
  XNOR2_X1 U11692 ( .A(n11494), .B(n9184), .ZN(n12936) );
  OR2_X1 U11693 ( .A1(n12936), .A2(n8888), .ZN(n9186) );
  OR2_X1 U11694 ( .A1(n12333), .A2(n12937), .ZN(n9185) );
  NAND2_X1 U11695 ( .A1(n9201), .A2(n12185), .ZN(n12393) );
  XNOR2_X1 U11696 ( .A(n9187), .B(n9196), .ZN(n9195) );
  INV_X1 U11697 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14492) );
  NAND2_X1 U11698 ( .A1(n9188), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9190) );
  NAND2_X1 U11699 ( .A1(n12346), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9189) );
  OAI211_X1 U11700 ( .C1(n14492), .C2(n8731), .A(n9190), .B(n9189), .ZN(n9191)
         );
  INV_X1 U11701 ( .A(n9191), .ZN(n9192) );
  INV_X1 U11702 ( .A(P3_B_REG_SCAN_IN), .ZN(n9193) );
  OAI21_X1 U11703 ( .B1(n9130), .B2(n9193), .A(n12769), .ZN(n12659) );
  OAI22_X1 U11704 ( .A1(n11510), .A2(n12799), .B1(n12354), .B2(n12659), .ZN(
        n9194) );
  INV_X1 U11705 ( .A(n9197), .ZN(n9198) );
  AOI21_X1 U11706 ( .B1(n11510), .B2(n12670), .A(n9198), .ZN(n12325) );
  NOR2_X1 U11707 ( .A1(n12670), .A2(n11510), .ZN(n12324) );
  XOR2_X1 U11708 ( .A(n12384), .B(n12398), .Z(n12424) );
  NAND2_X1 U11709 ( .A1(n12424), .A2(n15150), .ZN(n9199) );
  NAND2_X1 U11710 ( .A1(n12419), .A2(n9199), .ZN(n9203) );
  INV_X1 U11711 ( .A(n9200), .ZN(n9202) );
  NAND2_X1 U11712 ( .A1(n9202), .A2(n7445), .ZN(P3_U3456) );
  INV_X1 U11713 ( .A(n9204), .ZN(n9205) );
  NAND2_X1 U11714 ( .A1(n9205), .A2(n7447), .ZN(P3_U3488) );
  NAND4_X1 U11715 ( .A1(n9208), .A2(n9207), .A3(n9361), .A4(n9291), .ZN(n9209)
         );
  NOR2_X1 U11716 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), 
        .ZN(n9213) );
  NAND3_X1 U11717 ( .A1(n9216), .A2(n9215), .A3(n9214), .ZN(n9217) );
  OAI21_X1 U11718 ( .B1(n9265), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9222) );
  INV_X1 U11719 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9221) );
  NOR2_X1 U11720 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), 
        .ZN(n9225) );
  NAND4_X1 U11721 ( .A1(n9225), .A2(n9224), .A3(n9218), .A4(n9223), .ZN(n9240)
         );
  INV_X1 U11722 ( .A(n9272), .ZN(n9226) );
  NAND2_X1 U11723 ( .A1(n9226), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9227) );
  MUX2_X1 U11724 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9227), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n9228) );
  NAND2_X1 U11725 ( .A1(n9228), .A2(n9230), .ZN(n11090) );
  NAND2_X1 U11726 ( .A1(n9230), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9229) );
  XNOR2_X1 U11727 ( .A(n9229), .B(P1_IR_REG_25__SCAN_IN), .ZN(n11168) );
  AND2_X1 U11728 ( .A1(n9406), .A2(n11168), .ZN(n9231) );
  INV_X1 U11729 ( .A(n9432), .ZN(n9232) );
  INV_X2 U11730 ( .A(n14523), .ZN(n14502) );
  AOI211_X1 U11731 ( .C1(n9233), .C2(n9234), .A(n14502), .B(n6580), .ZN(n9239)
         );
  INV_X1 U11732 ( .A(n11273), .ZN(n11322) );
  NOR2_X1 U11733 ( .A1(n11322), .A2(n14515), .ZN(n9238) );
  NAND2_X1 U11734 ( .A1(n13054), .A2(n13372), .ZN(n14518) );
  OAI22_X1 U11735 ( .A1(n14518), .A2(n11391), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13150), .ZN(n9237) );
  NAND2_X1 U11736 ( .A1(n13054), .A2(n13370), .ZN(n14519) );
  OAI22_X1 U11737 ( .A1(n14519), .A2(n9235), .B1(n11270), .B2(n14528), .ZN(
        n9236) );
  OR4_X1 U11738 ( .A1(n9239), .A2(n9238), .A3(n9237), .A4(n9236), .ZN(P2_U3213) );
  AND2_X1 U11739 ( .A1(n14377), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n13709) );
  INV_X1 U11740 ( .A(n9240), .ZN(n9245) );
  XNOR2_X2 U11741 ( .A(n9248), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9521) );
  XNOR2_X2 U11742 ( .A(n9249), .B(P1_IR_REG_29__SCAN_IN), .ZN(n9519) );
  INV_X1 U11743 ( .A(n9605), .ZN(n9250) );
  NAND2_X1 U11744 ( .A1(n9250), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9253) );
  INV_X1 U11745 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9251) );
  INV_X1 U11746 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9252) );
  INV_X1 U11747 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9277) );
  NAND2_X1 U11748 ( .A1(n9254), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9255) );
  INV_X1 U11749 ( .A(n9261), .ZN(n9262) );
  NAND2_X1 U11750 ( .A1(n9262), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9263) );
  MUX2_X1 U11751 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9263), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n9264) );
  XNOR2_X2 U11752 ( .A(n9266), .B(P1_IR_REG_22__SCAN_IN), .ZN(n11840) );
  NAND2_X1 U11753 ( .A1(n13702), .A2(n10328), .ZN(n9276) );
  INV_X1 U11754 ( .A(n14377), .ZN(n14583) );
  NOR2_X1 U11755 ( .A1(n6450), .A2(n14225), .ZN(n9267) );
  XNOR2_X2 U11756 ( .A(n9270), .B(n9269), .ZN(n11492) );
  NAND2_X1 U11757 ( .A1(n9272), .A2(n9271), .ZN(n9273) );
  OAI22_X1 U11758 ( .A1(n6617), .A2(n10161), .B1(n10182), .B2(n14583), .ZN(
        n9275) );
  NAND2_X1 U11759 ( .A1(n13702), .A2(n9765), .ZN(n9279) );
  INV_X1 U11760 ( .A(n10135), .ZN(n9766) );
  OAI21_X1 U11761 ( .B1(n9280), .B2(n9691), .A(n9693), .ZN(n9683) );
  INV_X1 U11762 ( .A(n9683), .ZN(n9282) );
  MUX2_X1 U11763 ( .A(n13709), .B(n9282), .S(n6453), .Z(n9284) );
  INV_X1 U11764 ( .A(n11492), .ZN(n9707) );
  INV_X1 U11765 ( .A(n6453), .ZN(n14582) );
  AOI21_X1 U11766 ( .B1(n14582), .B2(n9251), .A(n11492), .ZN(n14581) );
  OAI21_X1 U11767 ( .B1(n14581), .B2(n14377), .A(n13701), .ZN(n9283) );
  AOI21_X1 U11768 ( .B1(n9284), .B2(n9707), .A(n9283), .ZN(n9330) );
  INV_X1 U11769 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n14326) );
  OR2_X1 U11770 ( .A1(n9285), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n9287) );
  NAND2_X1 U11771 ( .A1(n9287), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9286) );
  MUX2_X1 U11772 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9286), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n9290) );
  INV_X1 U11773 ( .A(n9287), .ZN(n9289) );
  INV_X1 U11774 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9288) );
  NAND2_X1 U11775 ( .A1(n9289), .A2(n9288), .ZN(n9360) );
  NAND2_X1 U11776 ( .A1(n9290), .A2(n9360), .ZN(n10140) );
  MUX2_X1 U11777 ( .A(n14326), .B(P1_REG2_REG_4__SCAN_IN), .S(n10140), .Z(
        n9304) );
  INV_X1 U11778 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9774) );
  NAND2_X1 U11779 ( .A1(n9285), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9292) );
  XNOR2_X1 U11780 ( .A(n9291), .B(n9292), .ZN(n10151) );
  INV_X1 U11781 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9298) );
  NOR2_X1 U11782 ( .A1(n9293), .A2(n14216), .ZN(n9294) );
  INV_X1 U11783 ( .A(n9295), .ZN(n9296) );
  NAND2_X1 U11784 ( .A1(n9296), .A2(n9285), .ZN(n9762) );
  MUX2_X1 U11785 ( .A(n9298), .B(P1_REG2_REG_2__SCAN_IN), .S(n9762), .Z(n9323)
         );
  INV_X1 U11786 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10718) );
  INV_X1 U11787 ( .A(n9293), .ZN(n9297) );
  XNOR2_X1 U11788 ( .A(n9599), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n13710) );
  NAND2_X1 U11789 ( .A1(n13710), .A2(n13709), .ZN(n13708) );
  OAI21_X1 U11790 ( .B1(n9298), .B2(n9762), .A(n9321), .ZN(n13723) );
  XNOR2_X1 U11791 ( .A(n10151), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n13724) );
  NAND2_X1 U11792 ( .A1(n13723), .A2(n13724), .ZN(n13722) );
  NAND2_X1 U11793 ( .A1(n11840), .A2(n11843), .ZN(n11868) );
  INV_X1 U11794 ( .A(n11868), .ZN(n9678) );
  NAND2_X1 U11795 ( .A1(n9678), .A2(n10181), .ZN(n9299) );
  AND2_X1 U11796 ( .A1(n11680), .A2(n9299), .ZN(n9310) );
  OR2_X1 U11797 ( .A1(n9300), .A2(n9407), .ZN(n9681) );
  INV_X1 U11798 ( .A(n10181), .ZN(n9301) );
  NAND2_X1 U11799 ( .A1(n9301), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12084) );
  NAND2_X1 U11800 ( .A1(n9681), .A2(n12084), .ZN(n9311) );
  NAND2_X1 U11801 ( .A1(n9310), .A2(n9311), .ZN(n14587) );
  OR2_X1 U11802 ( .A1(n11492), .A2(n6453), .ZN(n9302) );
  OAI211_X1 U11803 ( .C1(n9304), .C2(n9303), .A(n14633), .B(n9489), .ZN(n9305)
         );
  INV_X1 U11804 ( .A(n9305), .ZN(n9317) );
  INV_X1 U11805 ( .A(n9762), .ZN(n9307) );
  INV_X1 U11806 ( .A(n9599), .ZN(n13707) );
  INV_X1 U11807 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9306) );
  XNOR2_X1 U11808 ( .A(n9599), .B(n9306), .ZN(n13704) );
  NOR3_X1 U11809 ( .A1(n13704), .A2(n9277), .A3(n14583), .ZN(n13703) );
  AOI21_X1 U11810 ( .B1(P1_REG1_REG_1__SCAN_IN), .B2(n13707), .A(n13703), .ZN(
        n9320) );
  INV_X1 U11811 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9607) );
  MUX2_X1 U11812 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9607), .S(n9762), .Z(n9319)
         );
  NOR2_X1 U11813 ( .A1(n9320), .A2(n9319), .ZN(n9318) );
  XOR2_X1 U11814 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10151), .Z(n13719) );
  XOR2_X1 U11815 ( .A(n10140), .B(P1_REG1_REG_4__SCAN_IN), .Z(n9308) );
  AOI211_X1 U11816 ( .C1(n9309), .C2(n9308), .A(n14665), .B(n9482), .ZN(n9316)
         );
  INV_X1 U11817 ( .A(n9310), .ZN(n9312) );
  AND2_X1 U11818 ( .A1(n9312), .A2(n9311), .ZN(n14585) );
  NAND2_X1 U11819 ( .A1(n14585), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n9314) );
  AND2_X1 U11820 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10189) );
  INV_X1 U11821 ( .A(n10189), .ZN(n9313) );
  OAI211_X1 U11822 ( .C1(n14618), .C2(n10140), .A(n9314), .B(n9313), .ZN(n9315) );
  OR4_X1 U11823 ( .A1(n9330), .A2(n9317), .A3(n9316), .A4(n9315), .ZN(P1_U3247) );
  AOI211_X1 U11824 ( .C1(n9320), .C2(n9319), .A(n9318), .B(n14665), .ZN(n9329)
         );
  OAI211_X1 U11825 ( .C1(n9323), .C2(n9322), .A(n14633), .B(n9321), .ZN(n9324)
         );
  INV_X1 U11826 ( .A(n9324), .ZN(n9328) );
  NAND2_X1 U11827 ( .A1(n14585), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n9326) );
  NAND2_X1 U11828 ( .A1(P1_U3086), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9325) );
  OAI211_X1 U11829 ( .C1(n14618), .C2(n9762), .A(n9326), .B(n9325), .ZN(n9327)
         );
  OR4_X1 U11830 ( .A1(n9330), .A2(n9329), .A3(n9328), .A4(n9327), .ZN(P1_U3245) );
  INV_X1 U11831 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n14322) );
  NOR2_X1 U11832 ( .A1(n6450), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12927) );
  INV_X2 U11833 ( .A(n12927), .ZN(n11500) );
  NAND2_X1 U11834 ( .A1(n6436), .A2(P3_U3151), .ZN(n12939) );
  INV_X1 U11835 ( .A(SI_0_), .ZN(n14225) );
  OAI222_X1 U11836 ( .A1(P3_U3151), .A2(n14322), .B1(n11500), .B2(n9332), .C1(
        n12939), .C2(n14225), .ZN(P3_U3295) );
  OAI222_X1 U11837 ( .A1(P3_U3151), .A2(n14994), .B1(n11500), .B2(n9334), .C1(
        n9333), .C2(n12939), .ZN(P3_U3289) );
  INV_X1 U11838 ( .A(n9335), .ZN(n9337) );
  INV_X1 U11839 ( .A(SI_2_), .ZN(n9336) );
  OAI222_X1 U11840 ( .A1(n10545), .A2(P3_U3151), .B1(n11500), .B2(n9337), .C1(
        n9336), .C2(n12939), .ZN(P3_U3293) );
  INV_X1 U11841 ( .A(n9338), .ZN(n9340) );
  INV_X1 U11842 ( .A(SI_3_), .ZN(n9339) );
  OAI222_X1 U11843 ( .A1(n14939), .A2(P3_U3151), .B1(n11500), .B2(n9340), .C1(
        n9339), .C2(n12939), .ZN(P3_U3292) );
  CLKBUF_X1 U11844 ( .A(n12939), .Z(n12933) );
  OAI222_X1 U11845 ( .A1(n12609), .A2(P3_U3151), .B1(n11500), .B2(n9342), .C1(
        n9341), .C2(n12933), .ZN(P3_U3287) );
  INV_X1 U11846 ( .A(n9343), .ZN(n9345) );
  INV_X1 U11847 ( .A(SI_7_), .ZN(n9344) );
  OAI222_X1 U11848 ( .A1(n10963), .A2(P3_U3151), .B1(n11500), .B2(n9345), .C1(
        n9344), .C2(n12933), .ZN(P3_U3288) );
  OAI222_X1 U11849 ( .A1(n11500), .A2(n9347), .B1(n12933), .B2(n9346), .C1(
        P3_U3151), .C2(n9844), .ZN(P3_U3294) );
  INV_X1 U11850 ( .A(SI_5_), .ZN(n9350) );
  INV_X1 U11851 ( .A(n9348), .ZN(n9349) );
  OAI222_X1 U11852 ( .A1(P3_U3151), .A2(n14977), .B1(n12933), .B2(n9350), .C1(
        n11500), .C2(n9349), .ZN(P3_U3290) );
  INV_X1 U11853 ( .A(SI_4_), .ZN(n9353) );
  INV_X1 U11854 ( .A(n9351), .ZN(n9352) );
  OAI222_X1 U11855 ( .A1(P3_U3151), .A2(n14967), .B1(n12933), .B2(n9353), .C1(
        n11500), .C2(n9352), .ZN(P3_U3291) );
  AND2_X1 U11856 ( .A1(n9354), .A2(P2_U3088), .ZN(n13541) );
  INV_X2 U11857 ( .A(n13541), .ZN(n13551) );
  OAI222_X1 U11858 ( .A1(P2_U3088), .A2(n9526), .B1(n13549), .B2(n9596), .C1(
        n9355), .C2(n13551), .ZN(P2_U3326) );
  INV_X1 U11859 ( .A(SI_9_), .ZN(n9358) );
  INV_X1 U11860 ( .A(n9356), .ZN(n9357) );
  OAI222_X1 U11861 ( .A1(P3_U3151), .A2(n15014), .B1(n12933), .B2(n9358), .C1(
        n11500), .C2(n9357), .ZN(P3_U3286) );
  NAND2_X1 U11862 ( .A1(n9360), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9359) );
  MUX2_X1 U11863 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9359), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n9363) );
  INV_X1 U11864 ( .A(n9360), .ZN(n9362) );
  NAND2_X1 U11865 ( .A1(n9362), .A2(n9361), .ZN(n9379) );
  INV_X1 U11866 ( .A(n13734), .ZN(n9490) );
  NOR2_X1 U11867 ( .A1(n6449), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14221) );
  INV_X2 U11868 ( .A(n14221), .ZN(n14375) );
  AND2_X1 U11869 ( .A1(n6436), .A2(P1_U3086), .ZN(n9592) );
  INV_X2 U11870 ( .A(n9592), .ZN(n14372) );
  OAI222_X1 U11871 ( .A1(P1_U3086), .A2(n9490), .B1(n14375), .B2(n10220), .C1(
        n9364), .C2(n14372), .ZN(P1_U3350) );
  INV_X1 U11872 ( .A(n9365), .ZN(n10148) );
  OAI222_X1 U11873 ( .A1(n14372), .A2(n10147), .B1(n14375), .B2(n10148), .C1(
        n10151), .C2(P1_U3086), .ZN(P1_U3352) );
  OAI222_X1 U11874 ( .A1(P1_U3086), .A2(n9599), .B1(n14375), .B2(n9596), .C1(
        n7509), .C2(n14372), .ZN(P1_U3354) );
  OAI222_X1 U11875 ( .A1(P1_U3086), .A2(n9762), .B1(n14375), .B2(n9758), .C1(
        n9759), .C2(n14372), .ZN(P1_U3353) );
  INV_X1 U11876 ( .A(n10136), .ZN(n9371) );
  OAI222_X1 U11877 ( .A1(n14372), .A2(n10137), .B1(n14375), .B2(n9371), .C1(
        n10140), .C2(P1_U3086), .ZN(P1_U3351) );
  NAND2_X1 U11878 ( .A1(n9379), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9366) );
  XNOR2_X1 U11879 ( .A(n9366), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10321) );
  INV_X1 U11880 ( .A(n10321), .ZN(n9746) );
  OAI222_X1 U11881 ( .A1(P1_U3086), .A2(n9746), .B1(n14375), .B2(n10320), .C1(
        n9367), .C2(n14372), .ZN(P1_U3349) );
  INV_X1 U11882 ( .A(n13110), .ZN(n9368) );
  OAI222_X1 U11883 ( .A1(n13551), .A2(n9369), .B1(n13549), .B2(n10148), .C1(
        P2_U3088), .C2(n9368), .ZN(P2_U3324) );
  OAI222_X1 U11884 ( .A1(P2_U3088), .A2(n9534), .B1(n13549), .B2(n9758), .C1(
        n9370), .C2(n13551), .ZN(P2_U3325) );
  INV_X1 U11885 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9372) );
  OAI222_X1 U11886 ( .A1(n13551), .A2(n9372), .B1(n13549), .B2(n9371), .C1(
        P2_U3088), .C2(n9554), .ZN(P2_U3323) );
  INV_X1 U11887 ( .A(n13142), .ZN(n9556) );
  OAI222_X1 U11888 ( .A1(P2_U3088), .A2(n9556), .B1(n13549), .B2(n10320), .C1(
        n9373), .C2(n13551), .ZN(P2_U3321) );
  INV_X1 U11889 ( .A(n13125), .ZN(n9375) );
  INV_X1 U11890 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9374) );
  OAI222_X1 U11891 ( .A1(P2_U3088), .A2(n9375), .B1(n13549), .B2(n10220), .C1(
        n9374), .C2(n13551), .ZN(P2_U3322) );
  INV_X1 U11892 ( .A(n12617), .ZN(n15033) );
  INV_X1 U11893 ( .A(SI_10_), .ZN(n14254) );
  INV_X1 U11894 ( .A(n9376), .ZN(n9377) );
  OAI222_X1 U11895 ( .A1(P3_U3151), .A2(n15033), .B1(n12933), .B2(n14254), 
        .C1(n11500), .C2(n9377), .ZN(P3_U3285) );
  INV_X1 U11896 ( .A(n9660), .ZN(n9563) );
  OAI222_X1 U11897 ( .A1(P2_U3088), .A2(n9563), .B1(n13549), .B2(n10561), .C1(
        n9378), .C2(n13551), .ZN(P2_U3320) );
  OAI21_X1 U11898 ( .B1(n9379), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9380) );
  XNOR2_X1 U11899 ( .A(n9380), .B(P1_IR_REG_7__SCAN_IN), .ZN(n13748) );
  INV_X1 U11900 ( .A(n13748), .ZN(n9747) );
  OAI222_X1 U11901 ( .A1(P1_U3086), .A2(n9747), .B1(n14375), .B2(n10561), .C1(
        n9381), .C2(n14372), .ZN(P1_U3348) );
  INV_X1 U11902 ( .A(n9382), .ZN(n9383) );
  OAI222_X1 U11903 ( .A1(P3_U3151), .A2(n15049), .B1(n12933), .B2(n9384), .C1(
        n11500), .C2(n9383), .ZN(P3_U3284) );
  NAND2_X1 U11904 ( .A1(n9386), .A2(P3_D_REG_1__SCAN_IN), .ZN(n9385) );
  OAI21_X1 U11905 ( .B1(n10584), .B2(n9386), .A(n9385), .ZN(P3_U3377) );
  OAI222_X1 U11906 ( .A1(P2_U3088), .A2(n9667), .B1(n13549), .B2(n10748), .C1(
        n9387), .C2(n13551), .ZN(P2_U3319) );
  NAND2_X1 U11907 ( .A1(n9388), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9389) );
  MUX2_X1 U11908 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9389), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n9390) );
  INV_X1 U11909 ( .A(n9390), .ZN(n9391) );
  NOR2_X1 U11910 ( .A1(n9391), .A2(n10211), .ZN(n10749) );
  INV_X1 U11911 ( .A(n10749), .ZN(n9953) );
  INV_X1 U11912 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9392) );
  OAI222_X1 U11913 ( .A1(P1_U3086), .A2(n9953), .B1(n14375), .B2(n10748), .C1(
        n9392), .C2(n14372), .ZN(P1_U3347) );
  INV_X1 U11914 ( .A(n9393), .ZN(n9394) );
  OAI222_X1 U11915 ( .A1(n12933), .A2(n14350), .B1(n11500), .B2(n9394), .C1(
        n15068), .C2(P3_U3151), .ZN(P3_U3283) );
  INV_X1 U11916 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n14241) );
  NOR2_X1 U11917 ( .A1(n9421), .A2(n14241), .ZN(P3_U3243) );
  INV_X1 U11918 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n14314) );
  NOR2_X1 U11919 ( .A1(n9421), .A2(n14314), .ZN(P3_U3258) );
  INV_X1 U11920 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n14277) );
  NOR2_X1 U11921 ( .A1(n9421), .A2(n14277), .ZN(P3_U3234) );
  INV_X1 U11922 ( .A(n9681), .ZN(n9685) );
  NAND2_X1 U11923 ( .A1(n11090), .A2(P1_B_REG_SCAN_IN), .ZN(n9397) );
  INV_X1 U11924 ( .A(P1_B_REG_SCAN_IN), .ZN(n13802) );
  NAND2_X1 U11925 ( .A1(n9406), .A2(n13802), .ZN(n9396) );
  INV_X1 U11926 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9672) );
  INV_X1 U11927 ( .A(n9407), .ZN(n9399) );
  OR2_X1 U11928 ( .A1(n11334), .A2(n11168), .ZN(n9676) );
  INV_X1 U11929 ( .A(n9676), .ZN(n9398) );
  AOI22_X1 U11930 ( .A1(n14765), .A2(n9672), .B1(n9399), .B2(n9398), .ZN(
        P1_U3446) );
  NOR2_X1 U11931 ( .A1(n10211), .A2(n14216), .ZN(n9400) );
  MUX2_X1 U11932 ( .A(n14216), .B(n9400), .S(P1_IR_REG_9__SCAN_IN), .Z(n9402)
         );
  INV_X1 U11933 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9401) );
  NOR2_X1 U11934 ( .A1(n9402), .A2(n9416), .ZN(n10726) );
  INV_X1 U11935 ( .A(n10726), .ZN(n9961) );
  OAI222_X1 U11936 ( .A1(P1_U3086), .A2(n9961), .B1(n14375), .B2(n10725), .C1(
        n9403), .C2(n14372), .ZN(P1_U3346) );
  INV_X1 U11937 ( .A(n10120), .ZN(n9405) );
  OAI222_X1 U11938 ( .A1(P2_U3088), .A2(n9405), .B1(n13549), .B2(n10725), .C1(
        n9404), .C2(n13551), .ZN(P2_U3318) );
  INV_X1 U11939 ( .A(n14765), .ZN(n14764) );
  OAI22_X1 U11940 ( .A1(n14764), .A2(P1_D_REG_0__SCAN_IN), .B1(n9407), .B2(
        n9512), .ZN(n9408) );
  INV_X1 U11941 ( .A(n9408), .ZN(P1_U3445) );
  INV_X1 U11942 ( .A(n9465), .ZN(n9858) );
  INV_X2 U11943 ( .A(P2_U3947), .ZN(n13096) );
  MUX2_X1 U11944 ( .A(n9858), .B(n8725), .S(n13096), .Z(n9409) );
  INV_X1 U11945 ( .A(n9409), .ZN(P2_U3531) );
  AND2_X1 U11946 ( .A1(n9410), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U11947 ( .A1(n9410), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U11948 ( .A1(n9410), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U11949 ( .A1(n9410), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U11950 ( .A1(n9410), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U11951 ( .A1(n9410), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U11952 ( .A1(n9410), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U11953 ( .A1(n9410), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U11954 ( .A1(n9410), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U11955 ( .A1(n9410), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  OAI222_X1 U11956 ( .A1(P3_U3151), .A2(n15084), .B1(n12939), .B2(n9412), .C1(
        n11500), .C2(n9411), .ZN(P3_U3282) );
  INV_X1 U11957 ( .A(n10373), .ZN(n10126) );
  OAI222_X1 U11958 ( .A1(P2_U3088), .A2(n10126), .B1(n13549), .B2(n10843), 
        .C1(n9413), .C2(n13551), .ZN(P2_U3317) );
  NOR2_X1 U11959 ( .A1(n9416), .A2(n14216), .ZN(n9414) );
  MUX2_X1 U11960 ( .A(n14216), .B(n9414), .S(P1_IR_REG_10__SCAN_IN), .Z(n9418)
         );
  INV_X1 U11961 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9415) );
  NAND2_X1 U11962 ( .A1(n9416), .A2(n9415), .ZN(n9591) );
  INV_X1 U11963 ( .A(n9591), .ZN(n9417) );
  INV_X1 U11964 ( .A(n14597), .ZN(n9420) );
  OAI222_X1 U11965 ( .A1(P1_U3086), .A2(n9420), .B1(n14375), .B2(n10843), .C1(
        n9419), .C2(n14372), .ZN(P1_U3345) );
  INV_X1 U11966 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n9425) );
  INV_X1 U11967 ( .A(n9422), .ZN(n9424) );
  AOI22_X1 U11968 ( .A1(n9410), .A2(n9425), .B1(n9424), .B2(n9423), .ZN(
        P3_U3376) );
  AND2_X1 U11969 ( .A1(n9410), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U11970 ( .A1(n9410), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U11971 ( .A1(n9410), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U11972 ( .A1(n9410), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U11973 ( .A1(n9410), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U11974 ( .A1(n9410), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U11975 ( .A1(n9410), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U11976 ( .A1(n9410), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U11977 ( .A1(n9410), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U11978 ( .A1(n9410), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U11979 ( .A1(n9410), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U11980 ( .A1(n9410), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U11981 ( .A1(n9410), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U11982 ( .A1(n9410), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U11983 ( .A1(n9410), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U11984 ( .A1(n9410), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U11985 ( .A1(n9410), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  OAI222_X1 U11986 ( .A1(n15100), .A2(P3_U3151), .B1(n11500), .B2(n9426), .C1(
        n12933), .C2(n14351), .ZN(P3_U3281) );
  NAND2_X1 U11987 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9437) );
  INV_X1 U11988 ( .A(n9427), .ZN(n9436) );
  OAI21_X1 U11989 ( .B1(n9432), .B2(n9429), .A(n9428), .ZN(n9434) );
  NAND3_X1 U11990 ( .A1(n9432), .A2(n9431), .A3(n9430), .ZN(n9433) );
  NAND2_X1 U11991 ( .A1(n9434), .A2(n9433), .ZN(n9448) );
  INV_X1 U11992 ( .A(n9448), .ZN(n9435) );
  NAND2_X1 U11993 ( .A1(n9438), .A2(n9439), .ZN(n9441) );
  INV_X1 U11994 ( .A(n6698), .ZN(n11538) );
  AOI211_X1 U11995 ( .C1(n9437), .C2(n9436), .A(n9527), .B(n14856), .ZN(n9447)
         );
  INV_X1 U11996 ( .A(n9438), .ZN(n9440) );
  XNOR2_X1 U11997 ( .A(n9526), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n9444) );
  AND2_X1 U11998 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9443) );
  INV_X1 U11999 ( .A(n9441), .ZN(n9442) );
  NAND2_X1 U12000 ( .A1(n9444), .A2(n9443), .ZN(n9533) );
  OAI211_X1 U12001 ( .C1(n9444), .C2(n9443), .A(n13224), .B(n9533), .ZN(n9445)
         );
  OAI21_X1 U12002 ( .B1(n13184), .B2(n9526), .A(n9445), .ZN(n9446) );
  NOR2_X1 U12003 ( .A1(n9447), .A2(n9446), .ZN(n9450) );
  AND2_X1 U12004 ( .A1(n9448), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14840) );
  AOI22_X1 U12005 ( .A1(n14840), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n9449) );
  NAND2_X1 U12006 ( .A1(n9450), .A2(n9449), .ZN(P2_U3215) );
  NOR2_X1 U12007 ( .A1(n14585), .A2(n13701), .ZN(P1_U3085) );
  NAND2_X1 U12008 ( .A1(n9591), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9451) );
  XNOR2_X1 U12009 ( .A(n9451), .B(P1_IR_REG_11__SCAN_IN), .ZN(n13762) );
  INV_X1 U12010 ( .A(n13762), .ZN(n9452) );
  INV_X1 U12011 ( .A(n10883), .ZN(n9453) );
  OAI222_X1 U12012 ( .A1(n9452), .A2(P1_U3086), .B1(n14375), .B2(n9453), .C1(
        n6703), .C2(n14372), .ZN(P1_U3344) );
  INV_X1 U12013 ( .A(n10501), .ZN(n10371) );
  OAI222_X1 U12014 ( .A1(n13551), .A2(n9454), .B1(n13549), .B2(n9453), .C1(
        P2_U3088), .C2(n10371), .ZN(P2_U3316) );
  AND2_X1 U12015 ( .A1(n9995), .A2(n9457), .ZN(n9642) );
  NAND2_X1 U12016 ( .A1(n9582), .A2(n6701), .ZN(n9460) );
  AND2_X1 U12017 ( .A1(n9575), .A2(n9460), .ZN(n10388) );
  INV_X1 U12018 ( .A(n9461), .ZN(n9581) );
  XNOR2_X1 U12019 ( .A(n9582), .B(n9581), .ZN(n9468) );
  AND2_X1 U12020 ( .A1(n7517), .A2(n9462), .ZN(n9463) );
  NAND2_X1 U12021 ( .A1(n13370), .A2(n9465), .ZN(n9467) );
  NAND2_X1 U12022 ( .A1(n13095), .A2(n13372), .ZN(n9466) );
  NAND2_X1 U12023 ( .A1(n9467), .A2(n9466), .ZN(n9734) );
  AOI21_X1 U12024 ( .B1(n9468), .B2(n13406), .A(n9734), .ZN(n10382) );
  NAND2_X1 U12025 ( .A1(n10384), .A2(n9857), .ZN(n9578) );
  OAI211_X1 U12026 ( .C1(n10384), .C2(n9857), .A(n13505), .B(n9578), .ZN(
        n10383) );
  INV_X1 U12027 ( .A(n10383), .ZN(n9469) );
  AOI21_X1 U12028 ( .B1(n13513), .B2(n8312), .A(n9469), .ZN(n9470) );
  OAI211_X1 U12029 ( .C1(n13516), .C2(n10388), .A(n10382), .B(n9470), .ZN(
        n9711) );
  NAND2_X1 U12030 ( .A1(n14933), .A2(n9711), .ZN(n9471) );
  OAI21_X1 U12031 ( .B1(n14933), .B2(n6979), .A(n9471), .ZN(P2_U3500) );
  INV_X1 U12032 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9472) );
  NAND2_X1 U12033 ( .A1(n13224), .A2(n9472), .ZN(n9473) );
  OAI211_X1 U12034 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n14856), .A(n9473), .B(
        n13184), .ZN(n9474) );
  INV_X1 U12035 ( .A(n9474), .ZN(n9477) );
  INV_X1 U12036 ( .A(n14856), .ZN(n13223) );
  AOI22_X1 U12037 ( .A1(n13223), .A2(P2_REG1_REG_0__SCAN_IN), .B1(n13224), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n9476) );
  MUX2_X1 U12038 ( .A(n9477), .B(n9476), .S(n9475), .Z(n9479) );
  AOI22_X1 U12039 ( .A1(n14840), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n9478) );
  NAND2_X1 U12040 ( .A1(n9479), .A2(n9478), .ZN(P2_U3214) );
  NAND2_X1 U12041 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n10340) );
  OAI21_X1 U12042 ( .B1(n14679), .B2(n9480), .A(n10340), .ZN(n9487) );
  INV_X1 U12043 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9481) );
  MUX2_X1 U12044 ( .A(n9481), .B(P1_REG1_REG_6__SCAN_IN), .S(n10321), .Z(n9485) );
  INV_X1 U12045 ( .A(n10140), .ZN(n9483) );
  AOI21_X1 U12046 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9483), .A(n9482), .ZN(
        n13730) );
  INV_X1 U12047 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10169) );
  MUX2_X1 U12048 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10169), .S(n13734), .Z(
        n13729) );
  NAND2_X1 U12049 ( .A1(n13730), .A2(n13729), .ZN(n13728) );
  OAI21_X1 U12050 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n13734), .A(n13728), .ZN(
        n9484) );
  NOR2_X1 U12051 ( .A1(n9484), .A2(n9485), .ZN(n9741) );
  AOI211_X1 U12052 ( .C1(n9485), .C2(n9484), .A(n14665), .B(n9741), .ZN(n9486)
         );
  AOI211_X1 U12053 ( .C1(n14676), .C2(n10321), .A(n9487), .B(n9486), .ZN(n9494) );
  INV_X1 U12054 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9488) );
  MUX2_X1 U12055 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n9488), .S(n10321), .Z(n9492) );
  INV_X1 U12056 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10170) );
  OAI21_X1 U12057 ( .B1(n14326), .B2(n10140), .A(n9489), .ZN(n13736) );
  MUX2_X1 U12058 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10170), .S(n13734), .Z(
        n13737) );
  NAND2_X1 U12059 ( .A1(n13736), .A2(n13737), .ZN(n13735) );
  OAI211_X1 U12060 ( .C1(n9492), .C2(n9491), .A(n14633), .B(n9745), .ZN(n9493)
         );
  NAND2_X1 U12061 ( .A1(n9494), .A2(n9493), .ZN(P1_U3249) );
  NAND2_X1 U12062 ( .A1(n9495), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9496) );
  INV_X1 U12063 ( .A(n14797), .ZN(n14805) );
  NAND2_X1 U12064 ( .A1(n14805), .A2(n9260), .ZN(n10180) );
  INV_X1 U12065 ( .A(n9675), .ZN(n9507) );
  NOR4_X1 U12066 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9500) );
  NOR4_X1 U12067 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n9499) );
  NOR4_X1 U12068 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9498) );
  NOR4_X1 U12069 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9497) );
  AND4_X1 U12070 ( .A1(n9500), .A2(n9499), .A3(n9498), .A4(n9497), .ZN(n9506)
         );
  NOR2_X1 U12071 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .ZN(
        n9504) );
  NOR4_X1 U12072 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n9503) );
  NOR4_X1 U12073 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n9502) );
  NOR4_X1 U12074 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n9501) );
  AND4_X1 U12075 ( .A1(n9504), .A2(n9503), .A3(n9502), .A4(n9501), .ZN(n9505)
         );
  NAND2_X1 U12076 ( .A1(n9506), .A2(n9505), .ZN(n9673) );
  NAND2_X1 U12077 ( .A1(n9507), .A2(n9673), .ZN(n9509) );
  OAI21_X1 U12078 ( .B1(n9675), .B2(P1_D_REG_1__SCAN_IN), .A(n9676), .ZN(n9508) );
  AND2_X1 U12079 ( .A1(n9509), .A2(n9508), .ZN(n9510) );
  AND2_X1 U12080 ( .A1(n10180), .A2(n9510), .ZN(n9620) );
  NAND2_X1 U12081 ( .A1(n11853), .A2(n13796), .ZN(n9511) );
  AND2_X1 U12082 ( .A1(n9678), .A2(n9511), .ZN(n10184) );
  AND3_X2 U12083 ( .A1(n9620), .A2(n12081), .A3(n10639), .ZN(n14839) );
  AND2_X1 U12084 ( .A1(n11840), .A2(n13796), .ZN(n9515) );
  NAND2_X1 U12085 ( .A1(n9514), .A2(n11840), .ZN(n9516) );
  NAND2_X1 U12086 ( .A1(n9516), .A2(n13796), .ZN(n9517) );
  OAI21_X1 U12087 ( .B1(n13702), .B2(n9278), .A(n10655), .ZN(n12032) );
  INV_X1 U12088 ( .A(n12032), .ZN(n10646) );
  NAND2_X1 U12089 ( .A1(n11840), .A2(n12058), .ZN(n11842) );
  NAND2_X1 U12090 ( .A1(n11843), .A2(n9602), .ZN(n11844) );
  NAND2_X1 U12091 ( .A1(n9678), .A2(n11492), .ZN(n14720) );
  INV_X1 U12092 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9518) );
  OR2_X2 U12093 ( .A1(n11816), .A2(n9518), .ZN(n9523) );
  INV_X1 U12094 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10717) );
  NAND2_X1 U12095 ( .A1(n9519), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9520) );
  NOR2_X1 U12096 ( .A1(n6465), .A2(n6521), .ZN(n9522) );
  NAND3_X2 U12097 ( .A1(n9522), .A2(n9523), .A3(n9524), .ZN(n13700) );
  AOI22_X1 U12098 ( .A1(n10646), .A2(n14685), .B1(n14702), .B2(n13700), .ZN(
        n10638) );
  OR3_X1 U12099 ( .A1(n6617), .A2(n11843), .A3(n11840), .ZN(n10644) );
  OAI211_X1 U12100 ( .C1(n14197), .C2(n12032), .A(n10638), .B(n10644), .ZN(
        n9621) );
  NAND2_X1 U12101 ( .A1(n9621), .A2(n14839), .ZN(n9525) );
  OAI21_X1 U12102 ( .B1(n14839), .B2(n9277), .A(n9525), .ZN(P1_U3528) );
  INV_X1 U12103 ( .A(n9526), .ZN(n9531) );
  INV_X1 U12104 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9528) );
  MUX2_X1 U12105 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n9528), .S(n9534), .Z(n9529)
         );
  NOR2_X1 U12106 ( .A1(n9530), .A2(n9529), .ZN(n9544) );
  AOI211_X1 U12107 ( .C1(n9530), .C2(n9529), .A(n9544), .B(n14856), .ZN(n9541)
         );
  NAND2_X1 U12108 ( .A1(n9531), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9532) );
  NAND2_X1 U12109 ( .A1(n9533), .A2(n9532), .ZN(n9535) );
  INV_X1 U12110 ( .A(n9535), .ZN(n9539) );
  INV_X1 U12111 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10061) );
  MUX2_X1 U12112 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10061), .S(n9534), .Z(n9538) );
  MUX2_X1 U12113 ( .A(n10061), .B(P2_REG2_REG_2__SCAN_IN), .S(n9534), .Z(n9536) );
  NAND2_X1 U12114 ( .A1(n9536), .A2(n9535), .ZN(n13106) );
  INV_X1 U12115 ( .A(n13106), .ZN(n9537) );
  AOI211_X1 U12116 ( .C1(n9539), .C2(n9538), .A(n9537), .B(n14864), .ZN(n9540)
         );
  AOI211_X1 U12117 ( .C1(n14862), .C2(n9551), .A(n9541), .B(n9540), .ZN(n9543)
         );
  AOI22_X1 U12118 ( .A1(n14840), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n9542) );
  NAND2_X1 U12119 ( .A1(n9543), .A2(n9542), .ZN(P2_U3216) );
  AOI21_X1 U12120 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n9551), .A(n9544), .ZN(
        n13100) );
  INV_X1 U12121 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9545) );
  MUX2_X1 U12122 ( .A(n9545), .B(P2_REG1_REG_3__SCAN_IN), .S(n13110), .Z(
        n13099) );
  NOR2_X1 U12123 ( .A1(n13100), .A2(n13099), .ZN(n13098) );
  AOI21_X1 U12124 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n13110), .A(n13098), .ZN(
        n14843) );
  INV_X1 U12125 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9546) );
  MUX2_X1 U12126 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9546), .S(n9554), .Z(n14842) );
  NOR2_X1 U12127 ( .A1(n14843), .A2(n14842), .ZN(n14841) );
  AOI21_X1 U12128 ( .B1(n14846), .B2(P2_REG1_REG_4__SCAN_IN), .A(n14841), .ZN(
        n13117) );
  INV_X1 U12129 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9547) );
  MUX2_X1 U12130 ( .A(n9547), .B(P2_REG1_REG_5__SCAN_IN), .S(n13125), .Z(
        n13116) );
  INV_X1 U12131 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9548) );
  MUX2_X1 U12132 ( .A(n9548), .B(P2_REG1_REG_6__SCAN_IN), .S(n13142), .Z(
        n13131) );
  INV_X1 U12133 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9549) );
  MUX2_X1 U12134 ( .A(n9549), .B(P2_REG1_REG_7__SCAN_IN), .S(n9660), .Z(n9550)
         );
  NOR2_X1 U12135 ( .A1(n6506), .A2(n9550), .ZN(n9656) );
  AOI211_X1 U12136 ( .C1(n6506), .C2(n9550), .A(n14856), .B(n9656), .ZN(n9566)
         );
  NAND2_X1 U12137 ( .A1(n9551), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n13105) );
  INV_X1 U12138 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9552) );
  MUX2_X1 U12139 ( .A(n9552), .B(P2_REG2_REG_3__SCAN_IN), .S(n13110), .Z(
        n13107) );
  AOI21_X1 U12140 ( .B1(n13106), .B2(n13105), .A(n13107), .ZN(n13104) );
  AOI21_X1 U12141 ( .B1(n13110), .B2(P2_REG2_REG_3__SCAN_IN), .A(n13104), .ZN(
        n14849) );
  INV_X1 U12142 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9553) );
  MUX2_X1 U12143 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n9553), .S(n9554), .Z(n14848) );
  NOR2_X1 U12144 ( .A1(n14849), .A2(n14848), .ZN(n14847) );
  NOR2_X1 U12145 ( .A1(n9554), .A2(n9553), .ZN(n13121) );
  INV_X1 U12146 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10265) );
  MUX2_X1 U12147 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10265), .S(n13125), .Z(
        n9555) );
  OAI21_X1 U12148 ( .B1(n14847), .B2(n13121), .A(n9555), .ZN(n13139) );
  NAND2_X1 U12149 ( .A1(n13125), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n13138) );
  INV_X1 U12150 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n14230) );
  MUX2_X1 U12151 ( .A(n14230), .B(P2_REG2_REG_6__SCAN_IN), .S(n13142), .Z(
        n13137) );
  AOI21_X1 U12152 ( .B1(n13139), .B2(n13138), .A(n13137), .ZN(n13136) );
  NOR2_X1 U12153 ( .A1(n9556), .A2(n14230), .ZN(n9559) );
  INV_X1 U12154 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9557) );
  MUX2_X1 U12155 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9557), .S(n9660), .Z(n9558)
         );
  OAI21_X1 U12156 ( .B1(n13136), .B2(n9559), .A(n9558), .ZN(n9663) );
  INV_X1 U12157 ( .A(n9663), .ZN(n9561) );
  NOR3_X1 U12158 ( .A1(n13136), .A2(n9559), .A3(n9558), .ZN(n9560) );
  NOR3_X1 U12159 ( .A1(n9561), .A2(n14864), .A3(n9560), .ZN(n9565) );
  NAND2_X1 U12160 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10034) );
  NAND2_X1 U12161 ( .A1(n14840), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n9562) );
  OAI211_X1 U12162 ( .C1(n13184), .C2(n9563), .A(n10034), .B(n9562), .ZN(n9564) );
  OR3_X1 U12163 ( .A1(n9566), .A2(n9565), .A3(n9564), .ZN(P2_U3221) );
  OAI222_X1 U12164 ( .A1(P3_U3151), .A2(n14408), .B1(n12933), .B2(n9568), .C1(
        n11500), .C2(n9567), .ZN(P3_U3280) );
  AND2_X1 U12165 ( .A1(n9458), .A2(n13294), .ZN(n9570) );
  INV_X1 U12166 ( .A(n13097), .ZN(n9569) );
  INV_X1 U12167 ( .A(n13372), .ZN(n13052) );
  OAI22_X1 U12168 ( .A1(n10249), .A2(n9570), .B1(n9569), .B2(n13052), .ZN(
        n10246) );
  OAI22_X1 U12169 ( .A1(n10249), .A2(n10420), .B1(n9571), .B2(n9857), .ZN(
        n9572) );
  NOR2_X1 U12170 ( .A1(n10246), .A2(n9572), .ZN(n14913) );
  NAND2_X1 U12171 ( .A1(n14931), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9573) );
  OAI21_X1 U12172 ( .B1(n14931), .B2(n14913), .A(n9573), .ZN(P2_U3499) );
  OR2_X1 U12173 ( .A1(n13097), .A2(n8312), .ZN(n9574) );
  INV_X1 U12174 ( .A(n9630), .ZN(n9576) );
  NAND2_X1 U12175 ( .A1(n9577), .A2(n9576), .ZN(n9624) );
  OAI21_X1 U12176 ( .B1(n9577), .B2(n9576), .A(n9624), .ZN(n10059) );
  INV_X1 U12177 ( .A(n8319), .ZN(n9942) );
  NAND2_X1 U12178 ( .A1(n9578), .A2(n8319), .ZN(n9579) );
  AND3_X1 U12179 ( .A1(n9627), .A2(n13505), .A3(n9579), .ZN(n10064) );
  INV_X1 U12180 ( .A(n10064), .ZN(n9580) );
  OAI21_X1 U12181 ( .B1(n9942), .B2(n14922), .A(n9580), .ZN(n9589) );
  NAND2_X1 U12182 ( .A1(n9582), .A2(n9581), .ZN(n9584) );
  OR2_X1 U12183 ( .A1(n13097), .A2(n10384), .ZN(n9583) );
  NAND2_X1 U12184 ( .A1(n9584), .A2(n9583), .ZN(n9631) );
  XNOR2_X1 U12185 ( .A(n9631), .B(n9630), .ZN(n9585) );
  NAND2_X1 U12186 ( .A1(n9585), .A2(n13406), .ZN(n9588) );
  NAND2_X1 U12187 ( .A1(n13370), .A2(n13097), .ZN(n9587) );
  NAND2_X1 U12188 ( .A1(n13094), .A2(n13372), .ZN(n9586) );
  AND2_X1 U12189 ( .A1(n9587), .A2(n9586), .ZN(n9941) );
  NAND2_X1 U12190 ( .A1(n9588), .A2(n9941), .ZN(n10063) );
  AOI211_X1 U12191 ( .C1(n14533), .C2(n10059), .A(n9589), .B(n10063), .ZN(
        n9643) );
  NAND2_X1 U12192 ( .A1(n14931), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9590) );
  OAI21_X1 U12193 ( .B1(n9643), .B2(n14931), .A(n9590), .ZN(P2_U3501) );
  INV_X1 U12194 ( .A(n10999), .ZN(n9595) );
  NAND2_X1 U12195 ( .A1(n10083), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9650) );
  XNOR2_X1 U12196 ( .A(n9650), .B(P1_IR_REG_12__SCAN_IN), .ZN(n13782) );
  AOI22_X1 U12197 ( .A1(n13782), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9592), .ZN(n9593) );
  OAI21_X1 U12198 ( .B1(n9595), .B2(n14375), .A(n9593), .ZN(P1_U3343) );
  OAI222_X1 U12199 ( .A1(P2_U3088), .A2(n11105), .B1(n13549), .B2(n9595), .C1(
        n9594), .C2(n13551), .ZN(P2_U3315) );
  OR2_X1 U12200 ( .A1(n11610), .A2(n9596), .ZN(n9598) );
  NAND2_X4 U12201 ( .A1(n6444), .A2(n6450), .ZN(n12023) );
  OAI211_X2 U12202 ( .C1(n11680), .C2(n9599), .A(n9598), .B(n9597), .ZN(n11876) );
  NAND2_X1 U12203 ( .A1(n13700), .A2(n9600), .ZN(n10649) );
  INV_X1 U12204 ( .A(n10656), .ZN(n12033) );
  XNOR2_X1 U12205 ( .A(n12033), .B(n10655), .ZN(n10724) );
  INV_X1 U12206 ( .A(n10724), .ZN(n9618) );
  NAND3_X1 U12207 ( .A1(n9601), .A2(n12058), .A3(n9260), .ZN(n9603) );
  NAND2_X1 U12208 ( .A1(n9260), .A2(n9602), .ZN(n12059) );
  OR2_X1 U12209 ( .A1(n12059), .A2(n11840), .ZN(n10662) );
  NAND2_X1 U12210 ( .A1(n11872), .A2(n6617), .ZN(n10692) );
  OAI21_X1 U12211 ( .B1(n11872), .B2(n6617), .A(n10692), .ZN(n9612) );
  INV_X1 U12212 ( .A(n9612), .ZN(n9604) );
  NAND2_X1 U12213 ( .A1(n9604), .A2(n14756), .ZN(n10719) );
  OAI21_X1 U12214 ( .B1(n11872), .B2(n14821), .A(n10719), .ZN(n9617) );
  NAND2_X1 U12215 ( .A1(n11814), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9611) );
  INV_X1 U12216 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10691) );
  OR2_X1 U12217 ( .A1(n9605), .A2(n10691), .ZN(n9610) );
  INV_X1 U12218 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9606) );
  OR2_X1 U12219 ( .A1(n11816), .A2(n9606), .ZN(n9609) );
  OR2_X1 U12220 ( .A1(n11818), .A2(n9607), .ZN(n9608) );
  XNOR2_X1 U12221 ( .A(n9612), .B(n13700), .ZN(n9613) );
  AOI21_X1 U12222 ( .B1(n9613), .B2(n14685), .A(n13702), .ZN(n9616) );
  AOI21_X1 U12223 ( .B1(n12033), .B2(n13702), .A(n14744), .ZN(n9614) );
  NOR2_X1 U12224 ( .A1(n9614), .A2(n14705), .ZN(n9615) );
  OAI222_X1 U12225 ( .A1(n14720), .A2(n13581), .B1(n10791), .B2(n10724), .C1(
        n9616), .C2(n9615), .ZN(n10716) );
  AOI211_X1 U12226 ( .C1(n14805), .C2(n9618), .A(n9617), .B(n10716), .ZN(
        n14766) );
  NAND2_X1 U12227 ( .A1(n14837), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9619) );
  OAI21_X1 U12228 ( .B1(n14766), .B2(n14837), .A(n9619), .ZN(P1_U3529) );
  AND3_X2 U12229 ( .A1(n9620), .A2(n12081), .A3(n9680), .ZN(n14827) );
  NAND2_X1 U12230 ( .A1(n9621), .A2(n14827), .ZN(n9622) );
  OAI21_X1 U12231 ( .B1(n14827), .B2(n9252), .A(n9622), .ZN(P1_U3459) );
  OR2_X1 U12232 ( .A1(n13095), .A2(n8319), .ZN(n9623) );
  NAND2_X1 U12233 ( .A1(n9624), .A2(n9623), .ZN(n9717) );
  NAND2_X1 U12234 ( .A1(n9717), .A2(n9721), .ZN(n9719) );
  OR2_X1 U12235 ( .A1(n13094), .A2(n10006), .ZN(n9625) );
  NAND2_X1 U12236 ( .A1(n9719), .A2(n9625), .ZN(n9626) );
  INV_X1 U12237 ( .A(n9787), .ZN(n9637) );
  NAND2_X1 U12238 ( .A1(n9626), .A2(n9637), .ZN(n9784) );
  OAI21_X1 U12239 ( .B1(n9626), .B2(n9637), .A(n9784), .ZN(n10068) );
  INV_X1 U12240 ( .A(n10073), .ZN(n9629) );
  INV_X1 U12241 ( .A(n10006), .ZN(n9729) );
  INV_X1 U12242 ( .A(n9727), .ZN(n9628) );
  INV_X1 U12243 ( .A(n9796), .ZN(n9798) );
  OAI21_X1 U12244 ( .B1(n9629), .B2(n9628), .A(n9798), .ZN(n10070) );
  INV_X1 U12245 ( .A(n13505), .ZN(n13409) );
  OAI22_X1 U12246 ( .A1(n10070), .A2(n13409), .B1(n9629), .B2(n14922), .ZN(
        n9639) );
  INV_X1 U12247 ( .A(n13092), .ZN(n10093) );
  NAND2_X1 U12248 ( .A1(n9631), .A2(n9630), .ZN(n9633) );
  INV_X1 U12249 ( .A(n13095), .ZN(n9720) );
  NAND2_X1 U12250 ( .A1(n9720), .A2(n8319), .ZN(n9632) );
  NAND2_X1 U12251 ( .A1(n9633), .A2(n9632), .ZN(n9722) );
  INV_X1 U12252 ( .A(n9721), .ZN(n9634) );
  NAND2_X1 U12253 ( .A1(n9722), .A2(n9634), .ZN(n9636) );
  NAND2_X1 U12254 ( .A1(n10006), .A2(n9983), .ZN(n9635) );
  NAND2_X1 U12255 ( .A1(n9636), .A2(n9635), .ZN(n9788) );
  XNOR2_X1 U12256 ( .A(n9788), .B(n9637), .ZN(n9638) );
  OAI222_X1 U12257 ( .A1(n13052), .A2(n10093), .B1(n13051), .B2(n9983), .C1(
        n13294), .C2(n9638), .ZN(n10074) );
  AOI211_X1 U12258 ( .C1(n14533), .C2(n10068), .A(n9639), .B(n10074), .ZN(
        n9714) );
  NAND2_X1 U12259 ( .A1(n14931), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9640) );
  OAI21_X1 U12260 ( .B1(n9714), .B2(n14931), .A(n9640), .ZN(P2_U3503) );
  INV_X1 U12261 ( .A(n9994), .ZN(n9641) );
  INV_X1 U12262 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9645) );
  OR2_X1 U12263 ( .A1(n9643), .A2(n14928), .ZN(n9644) );
  OAI21_X1 U12264 ( .B1(n6443), .B2(n9645), .A(n9644), .ZN(P2_U3436) );
  INV_X1 U12265 ( .A(n14421), .ZN(n12641) );
  OAI222_X1 U12266 ( .A1(n12939), .A2(n9647), .B1(n11500), .B2(n9646), .C1(
        n12641), .C2(P3_U3151), .ZN(P3_U3279) );
  INV_X1 U12267 ( .A(n14861), .ZN(n9649) );
  INV_X1 U12268 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9648) );
  OAI222_X1 U12269 ( .A1(P2_U3088), .A2(n9649), .B1(n13549), .B2(n11025), .C1(
        n9648), .C2(n13551), .ZN(P2_U3314) );
  INV_X1 U12270 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10080) );
  NAND2_X1 U12271 ( .A1(n9650), .A2(n10080), .ZN(n9651) );
  NAND2_X1 U12272 ( .A1(n9651), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9652) );
  INV_X1 U12273 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n10081) );
  NAND2_X1 U12274 ( .A1(n9652), .A2(n10081), .ZN(n9817) );
  OR2_X1 U12275 ( .A1(n9652), .A2(n10081), .ZN(n9653) );
  INV_X1 U12276 ( .A(n14610), .ZN(n13771) );
  OAI222_X1 U12277 ( .A1(P1_U3086), .A2(n13771), .B1(n14375), .B2(n11025), 
        .C1(n9654), .C2(n14372), .ZN(P1_U3342) );
  INV_X1 U12278 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n14271) );
  NAND2_X1 U12279 ( .A1(n12234), .A2(P3_U3897), .ZN(n9655) );
  OAI21_X1 U12280 ( .B1(P3_U3897), .B2(n14271), .A(n9655), .ZN(P3_U3500) );
  INV_X1 U12281 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9657) );
  MUX2_X1 U12282 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9657), .S(n9667), .Z(n9658)
         );
  AOI211_X1 U12283 ( .C1(n9659), .C2(n9658), .A(n14856), .B(n9802), .ZN(n9670)
         );
  NAND2_X1 U12284 ( .A1(n9660), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9662) );
  INV_X1 U12285 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n14242) );
  MUX2_X1 U12286 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n14242), .S(n9667), .Z(n9661) );
  AOI21_X1 U12287 ( .B1(n9663), .B2(n9662), .A(n9661), .ZN(n9807) );
  AND3_X1 U12288 ( .A1(n9663), .A2(n9662), .A3(n9661), .ZN(n9664) );
  NOR3_X1 U12289 ( .A1(n9807), .A2(n9664), .A3(n14864), .ZN(n9669) );
  NAND2_X1 U12290 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n12971) );
  INV_X1 U12291 ( .A(n12971), .ZN(n9665) );
  AOI21_X1 U12292 ( .B1(n14840), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n9665), .ZN(
        n9666) );
  OAI21_X1 U12293 ( .B1(n13184), .B2(n9667), .A(n9666), .ZN(n9668) );
  OR3_X1 U12294 ( .A1(n9670), .A2(n9669), .A3(n9668), .ZN(P2_U3222) );
  NOR2_X1 U12295 ( .A1(n9673), .A2(n9672), .ZN(n9674) );
  OR2_X1 U12296 ( .A1(n9675), .A2(n9674), .ZN(n9677) );
  AND2_X1 U12297 ( .A1(n9677), .A2(n9676), .ZN(n10178) );
  NAND2_X1 U12298 ( .A1(n12081), .A2(n10178), .ZN(n10640) );
  NAND2_X1 U12299 ( .A1(n10639), .A2(n9678), .ZN(n9679) );
  OR2_X1 U12300 ( .A1(n10640), .A2(n9679), .ZN(n9706) );
  INV_X1 U12301 ( .A(n6433), .ZN(n13683) );
  NOR2_X1 U12302 ( .A1(n9681), .A2(n9680), .ZN(n9684) );
  AND3_X1 U12303 ( .A1(n14821), .A2(n10178), .A3(n11868), .ZN(n9682) );
  NAND2_X1 U12304 ( .A1(n9683), .A2(n13645), .ZN(n9689) );
  NAND2_X1 U12305 ( .A1(n9684), .A2(n10178), .ZN(n9687) );
  INV_X1 U12306 ( .A(n10180), .ZN(n9686) );
  NAND2_X1 U12307 ( .A1(n9687), .A2(n14751), .ZN(n10826) );
  INV_X1 U12308 ( .A(n10826), .ZN(n13621) );
  NOR2_X1 U12309 ( .A1(n13621), .A2(n10184), .ZN(n9772) );
  INV_X1 U12310 ( .A(n9772), .ZN(n9705) );
  AOI22_X1 U12311 ( .A1(n9705), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n9278), .B2(
        n13685), .ZN(n9688) );
  OAI211_X1 U12312 ( .C1(n9671), .C2(n13683), .A(n9689), .B(n9688), .ZN(
        P1_U3232) );
  INV_X1 U12313 ( .A(P3_DATAO_REG_20__SCAN_IN), .ZN(n14309) );
  NAND2_X1 U12314 ( .A1(n12770), .A2(P3_U3897), .ZN(n9690) );
  OAI21_X1 U12315 ( .B1(P3_U3897), .B2(n14309), .A(n9690), .ZN(P3_U3511) );
  NAND2_X1 U12316 ( .A1(n9692), .A2(n10326), .ZN(n9694) );
  NAND2_X1 U12317 ( .A1(n11876), .A2(n10135), .ZN(n9696) );
  NAND2_X1 U12318 ( .A1(n9696), .A2(n9695), .ZN(n9697) );
  XNOR2_X1 U12319 ( .A(n9697), .B(n10225), .ZN(n9699) );
  AOI22_X1 U12320 ( .A1(n13700), .A2(n10328), .B1(n9765), .B2(n11876), .ZN(
        n9698) );
  NAND2_X1 U12321 ( .A1(n9699), .A2(n9698), .ZN(n9768) );
  INV_X1 U12322 ( .A(n9704), .ZN(n9702) );
  INV_X1 U12323 ( .A(n9769), .ZN(n9703) );
  AOI21_X1 U12324 ( .B1(n9704), .B2(n9701), .A(n9703), .ZN(n9710) );
  AOI22_X1 U12325 ( .A1(n9705), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n13685), .B2(
        n11876), .ZN(n9709) );
  INV_X1 U12326 ( .A(n9706), .ZN(n13582) );
  NAND2_X1 U12327 ( .A1(n13582), .A2(n9707), .ZN(n13667) );
  INV_X1 U12328 ( .A(n13667), .ZN(n13681) );
  AOI22_X1 U12329 ( .A1(n13681), .A2(n13702), .B1(n13699), .B2(n6433), .ZN(
        n9708) );
  OAI211_X1 U12330 ( .C1(n9710), .C2(n13688), .A(n9709), .B(n9708), .ZN(
        P1_U3222) );
  INV_X1 U12331 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9713) );
  NAND2_X1 U12332 ( .A1(n6443), .A2(n9711), .ZN(n9712) );
  OAI21_X1 U12333 ( .B1(n6443), .B2(n9713), .A(n9712), .ZN(P2_U3433) );
  INV_X1 U12334 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9716) );
  OR2_X1 U12335 ( .A1(n9714), .A2(n14928), .ZN(n9715) );
  OAI21_X1 U12336 ( .B1(n6443), .B2(n9716), .A(n9715), .ZN(P2_U3442) );
  INV_X1 U12337 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n14272) );
  OR2_X1 U12338 ( .A1(n9717), .A2(n9721), .ZN(n9718) );
  NAND2_X1 U12339 ( .A1(n9719), .A2(n9718), .ZN(n9726) );
  INV_X1 U12340 ( .A(n9726), .ZN(n10010) );
  INV_X1 U12341 ( .A(n9458), .ZN(n10401) );
  INV_X1 U12342 ( .A(n13093), .ZN(n9972) );
  OAI22_X1 U12343 ( .A1(n9972), .A2(n13052), .B1(n9720), .B2(n13051), .ZN(
        n9725) );
  XNOR2_X1 U12344 ( .A(n9721), .B(n9722), .ZN(n9723) );
  NOR2_X1 U12345 ( .A1(n9723), .A2(n13294), .ZN(n9724) );
  AOI211_X1 U12346 ( .C1(n10401), .C2(n9726), .A(n9725), .B(n9724), .ZN(n10007) );
  OAI21_X1 U12347 ( .B1(n9729), .B2(n9728), .A(n9727), .ZN(n10004) );
  INV_X1 U12348 ( .A(n10004), .ZN(n9730) );
  AOI22_X1 U12349 ( .A1(n9730), .A2(n13505), .B1(n13513), .B2(n10006), .ZN(
        n9731) );
  OAI211_X1 U12350 ( .C1(n10010), .C2(n10420), .A(n10007), .B(n9731), .ZN(
        n13521) );
  NAND2_X1 U12351 ( .A1(n13521), .A2(n6443), .ZN(n9732) );
  OAI21_X1 U12352 ( .B1(n6443), .B2(n14272), .A(n9732), .ZN(P2_U3439) );
  NOR2_X1 U12353 ( .A1(n9733), .A2(P2_U3088), .ZN(n9940) );
  INV_X1 U12354 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10381) );
  AOI22_X1 U12355 ( .A1(n13054), .A2(n9734), .B1(n14507), .B2(n8312), .ZN(
        n9739) );
  OAI21_X1 U12356 ( .B1(n9736), .B2(n9735), .A(n9944), .ZN(n9737) );
  NAND2_X1 U12357 ( .A1(n14523), .A2(n9737), .ZN(n9738) );
  OAI211_X1 U12358 ( .C1(n9940), .C2(n10381), .A(n9739), .B(n9738), .ZN(
        P2_U3194) );
  INV_X1 U12359 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n14258) );
  NAND2_X1 U12360 ( .A1(n11485), .A2(P3_U3897), .ZN(n9740) );
  OAI21_X1 U12361 ( .B1(P3_U3897), .B2(n14258), .A(n9740), .ZN(P3_U3504) );
  INV_X1 U12362 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9742) );
  MUX2_X1 U12363 ( .A(n9742), .B(P1_REG1_REG_7__SCAN_IN), .S(n13748), .Z(
        n13742) );
  INV_X1 U12364 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10573) );
  MUX2_X1 U12365 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10573), .S(n10749), .Z(
        n9743) );
  OAI21_X1 U12366 ( .B1(n9744), .B2(n9743), .A(n9957), .ZN(n9754) );
  INV_X1 U12367 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10331) );
  OAI21_X1 U12368 ( .B1(n9488), .B2(n9746), .A(n9745), .ZN(n13750) );
  MUX2_X1 U12369 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10331), .S(n13748), .Z(
        n13751) );
  NAND2_X1 U12370 ( .A1(n13750), .A2(n13751), .ZN(n13749) );
  OAI21_X1 U12371 ( .B1(n9747), .B2(n10331), .A(n13749), .ZN(n9750) );
  INV_X1 U12372 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9748) );
  MUX2_X1 U12373 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n9748), .S(n10749), .Z(n9749) );
  NAND2_X1 U12374 ( .A1(n9750), .A2(n9749), .ZN(n9952) );
  OAI211_X1 U12375 ( .C1(n9750), .C2(n9749), .A(n9952), .B(n14633), .ZN(n9752)
         );
  INV_X1 U12376 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n14306) );
  NOR2_X1 U12377 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14306), .ZN(n10823) );
  AOI21_X1 U12378 ( .B1(n14585), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n10823), .ZN(
        n9751) );
  OAI211_X1 U12379 ( .C1(n14618), .C2(n9953), .A(n9752), .B(n9751), .ZN(n9753)
         );
  AOI21_X1 U12380 ( .B1(n9754), .B2(n14636), .A(n9753), .ZN(n9755) );
  INV_X1 U12381 ( .A(n9755), .ZN(P1_U3251) );
  OAI222_X1 U12382 ( .A1(P3_U3151), .A2(n12643), .B1(n12939), .B2(n9757), .C1(
        n11500), .C2(n9756), .ZN(P3_U3278) );
  INV_X1 U12383 ( .A(n10328), .ZN(n10153) );
  OR2_X1 U12384 ( .A1(n13581), .A2(n10153), .ZN(n9764) );
  OR2_X1 U12385 ( .A1(n11610), .A2(n9758), .ZN(n9761) );
  OR2_X1 U12386 ( .A1(n12023), .A2(n9759), .ZN(n9760) );
  NAND2_X1 U12387 ( .A1(n10695), .A2(n11775), .ZN(n9763) );
  NAND2_X1 U12388 ( .A1(n9764), .A2(n9763), .ZN(n10142) );
  OAI22_X1 U12389 ( .A1(n13581), .A2(n10161), .B1(n6952), .B2(n9766), .ZN(
        n9767) );
  XNOR2_X1 U12390 ( .A(n9767), .B(n10225), .ZN(n10144) );
  XNOR2_X1 U12391 ( .A(n10142), .B(n10144), .ZN(n9771) );
  NAND2_X1 U12392 ( .A1(n9769), .A2(n9768), .ZN(n9770) );
  OAI21_X1 U12393 ( .B1(n9771), .B2(n9770), .A(n10146), .ZN(n9781) );
  NAND2_X1 U12394 ( .A1(n10695), .A2(n14792), .ZN(n14768) );
  OAI22_X1 U12395 ( .A1(n9772), .A2(n10691), .B1(n13621), .B2(n14768), .ZN(
        n9780) );
  NAND2_X1 U12396 ( .A1(n11846), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9778) );
  OR2_X1 U12397 ( .A1(n9605), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9777) );
  INV_X1 U12398 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9773) );
  OR2_X1 U12399 ( .A1(n11818), .A2(n9773), .ZN(n9776) );
  OR2_X1 U12400 ( .A1(n11839), .A2(n9774), .ZN(n9775) );
  AND4_X2 U12401 ( .A1(n9778), .A2(n9777), .A3(n9776), .A4(n9775), .ZN(n10687)
         );
  OAI22_X1 U12402 ( .A1(n13683), .A2(n10687), .B1(n9671), .B2(n13667), .ZN(
        n9779) );
  AOI211_X1 U12403 ( .C1(n9781), .C2(n13645), .A(n9780), .B(n9779), .ZN(n9782)
         );
  INV_X1 U12404 ( .A(n9782), .ZN(P1_U3237) );
  INV_X1 U12405 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9801) );
  OR2_X1 U12406 ( .A1(n10073), .A2(n13093), .ZN(n9783) );
  NAND2_X1 U12407 ( .A1(n9784), .A2(n9783), .ZN(n9786) );
  INV_X1 U12408 ( .A(n9785), .ZN(n9791) );
  OAI21_X1 U12409 ( .B1(n9786), .B2(n9791), .A(n9924), .ZN(n9795) );
  INV_X1 U12410 ( .A(n9795), .ZN(n10272) );
  INV_X1 U12411 ( .A(n13091), .ZN(n10035) );
  OAI22_X1 U12412 ( .A1(n9972), .A2(n13051), .B1(n10035), .B2(n13052), .ZN(
        n9794) );
  NAND2_X1 U12413 ( .A1(n9788), .A2(n9787), .ZN(n9790) );
  NAND2_X1 U12414 ( .A1(n10073), .A2(n9972), .ZN(n9789) );
  XNOR2_X1 U12415 ( .A(n9928), .B(n9791), .ZN(n9792) );
  NOR2_X1 U12416 ( .A1(n9792), .A2(n13294), .ZN(n9793) );
  AOI211_X1 U12417 ( .C1(n10401), .C2(n9795), .A(n9794), .B(n9793), .ZN(n10264) );
  INV_X1 U12418 ( .A(n9973), .ZN(n10267) );
  NAND2_X1 U12419 ( .A1(n9796), .A2(n10267), .ZN(n9936) );
  INV_X1 U12420 ( .A(n9936), .ZN(n9797) );
  AOI211_X1 U12421 ( .C1(n9973), .C2(n9798), .A(n13409), .B(n9797), .ZN(n10269) );
  AOI21_X1 U12422 ( .B1(n13513), .B2(n9973), .A(n10269), .ZN(n9799) );
  OAI211_X1 U12423 ( .C1(n10272), .C2(n10420), .A(n10264), .B(n9799), .ZN(
        n13520) );
  NAND2_X1 U12424 ( .A1(n13520), .A2(n6443), .ZN(n9800) );
  OAI21_X1 U12425 ( .B1(n6443), .B2(n9801), .A(n9800), .ZN(P2_U3445) );
  INV_X1 U12426 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9803) );
  MUX2_X1 U12427 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n9803), .S(n10120), .Z(n9804) );
  OAI21_X1 U12428 ( .B1(n9805), .B2(n9804), .A(n10116), .ZN(n9806) );
  NAND2_X1 U12429 ( .A1(n9806), .A2(n13223), .ZN(n9816) );
  AOI21_X1 U12430 ( .B1(n9808), .B2(P2_REG2_REG_8__SCAN_IN), .A(n9807), .ZN(
        n9811) );
  INV_X1 U12431 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9809) );
  MUX2_X1 U12432 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n9809), .S(n10120), .Z(n9810) );
  NAND2_X1 U12433 ( .A1(n9811), .A2(n9810), .ZN(n10119) );
  OAI21_X1 U12434 ( .B1(n9811), .B2(n9810), .A(n10119), .ZN(n9814) );
  INV_X1 U12435 ( .A(n14840), .ZN(n14871) );
  NAND2_X1 U12436 ( .A1(n14862), .A2(n10120), .ZN(n9812) );
  NAND2_X1 U12437 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n10199) );
  OAI211_X1 U12438 ( .C1(n14393), .C2(n14871), .A(n9812), .B(n10199), .ZN(
        n9813) );
  AOI21_X1 U12439 ( .B1(n9814), .B2(n13224), .A(n9813), .ZN(n9815) );
  NAND2_X1 U12440 ( .A1(n9816), .A2(n9815), .ZN(P2_U3223) );
  INV_X1 U12441 ( .A(n11281), .ZN(n9820) );
  NAND2_X1 U12442 ( .A1(n9817), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9818) );
  XNOR2_X1 U12443 ( .A(n9818), .B(P1_IR_REG_14__SCAN_IN), .ZN(n13783) );
  INV_X1 U12444 ( .A(n13783), .ZN(n14617) );
  OAI222_X1 U12445 ( .A1(n14372), .A2(n9819), .B1(n14375), .B2(n9820), .C1(
        n14617), .C2(P1_U3086), .ZN(P1_U3341) );
  INV_X1 U12446 ( .A(n13148), .ZN(n11107) );
  OAI222_X1 U12447 ( .A1(n13551), .A2(n9821), .B1(n13549), .B2(n9820), .C1(
        P2_U3088), .C2(n11107), .ZN(P2_U3313) );
  AOI211_X1 U12448 ( .C1(n9823), .C2(n9822), .A(n14502), .B(n7575), .ZN(n9827)
         );
  INV_X1 U12449 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n13102) );
  INV_X1 U12450 ( .A(n14519), .ZN(n12979) );
  INV_X1 U12451 ( .A(n14518), .ZN(n9861) );
  AOI22_X1 U12452 ( .A1(n12979), .A2(n13095), .B1(n9861), .B2(n13093), .ZN(
        n9825) );
  AOI22_X1 U12453 ( .A1(n14507), .A2(n10006), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n9824) );
  OAI211_X1 U12454 ( .C1(n14528), .C2(P2_REG3_REG_3__SCAN_IN), .A(n9825), .B(
        n9824), .ZN(n9826) );
  OR2_X1 U12455 ( .A1(n9827), .A2(n9826), .ZN(P2_U3190) );
  INV_X1 U12456 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11833) );
  INV_X1 U12457 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n9828) );
  NOR2_X1 U12458 ( .A1(n10517), .A2(n9829), .ZN(n9830) );
  AOI21_X1 U12459 ( .B1(P3_REG1_REG_1__SCAN_IN), .B2(n12646), .A(n9830), .ZN(
        n9831) );
  INV_X1 U12460 ( .A(n9844), .ZN(n9852) );
  NAND2_X1 U12461 ( .A1(n9831), .A2(n9852), .ZN(n9901) );
  OAI21_X1 U12462 ( .B1(n9831), .B2(n9852), .A(n9901), .ZN(n9832) );
  AOI21_X1 U12463 ( .B1(n9872), .B2(n9832), .A(n9903), .ZN(n9855) );
  NAND2_X1 U12464 ( .A1(P3_U3897), .A2(n9130), .ZN(n15109) );
  NAND2_X1 U12465 ( .A1(n12327), .A2(n9885), .ZN(n9833) );
  AND2_X1 U12466 ( .A1(n6439), .A2(n9833), .ZN(n9839) );
  OR2_X1 U12467 ( .A1(n9885), .A2(P3_U3151), .ZN(n12417) );
  NAND2_X1 U12468 ( .A1(n9880), .A2(n12417), .ZN(n9838) );
  NAND2_X1 U12469 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n14322), .ZN(n9906) );
  NOR2_X1 U12470 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n9906), .ZN(n9835) );
  AOI21_X1 U12471 ( .B1(n9852), .B2(n9906), .A(n9835), .ZN(n9837) );
  AND2_X1 U12472 ( .A1(n9837), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9907) );
  INV_X1 U12473 ( .A(n9907), .ZN(n9836) );
  OAI21_X1 U12474 ( .B1(P3_REG1_REG_1__SCAN_IN), .B2(n9837), .A(n9836), .ZN(
        n9849) );
  INV_X1 U12475 ( .A(n9838), .ZN(n9840) );
  OR2_X1 U12476 ( .A1(n9840), .A2(n9839), .ZN(n15104) );
  OAI22_X1 U12477 ( .A1(n15104), .A2(n6720), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10608), .ZN(n9848) );
  INV_X1 U12478 ( .A(n9841), .ZN(n9842) );
  AND2_X1 U12479 ( .A1(n14322), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9866) );
  NAND2_X1 U12480 ( .A1(n8737), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9843) );
  OAI21_X1 U12481 ( .B1(n9844), .B2(n9866), .A(n9843), .ZN(n9845) );
  AOI21_X1 U12482 ( .B1(n9829), .B2(n9845), .A(n9915), .ZN(n9846) );
  NOR2_X1 U12483 ( .A1(n15116), .A2(n9846), .ZN(n9847) );
  AOI211_X1 U12484 ( .C1(n15107), .C2(n9849), .A(n9848), .B(n9847), .ZN(n9854)
         );
  INV_X1 U12485 ( .A(n9850), .ZN(n9851) );
  MUX2_X1 U12486 ( .A(n12558), .B(n9851), .S(n9130), .Z(n15101) );
  NAND2_X1 U12487 ( .A1(n15000), .A2(n9852), .ZN(n9853) );
  OAI211_X1 U12488 ( .C1(n9855), .C2(n15109), .A(n9854), .B(n9853), .ZN(
        P3_U3183) );
  INV_X1 U12489 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10248) );
  NOR2_X1 U12490 ( .A1(n14502), .A2(n9856), .ZN(n13040) );
  INV_X1 U12491 ( .A(n13040), .ZN(n12977) );
  OAI22_X1 U12492 ( .A1(n12977), .A2(n9858), .B1(n9857), .B2(n14502), .ZN(
        n9860) );
  NAND2_X1 U12493 ( .A1(n9860), .A2(n9859), .ZN(n9863) );
  AOI22_X1 U12494 ( .A1(n9861), .A2(n13097), .B1(n10252), .B2(n14507), .ZN(
        n9862) );
  OAI211_X1 U12495 ( .C1(n9940), .C2(n10248), .A(n9863), .B(n9862), .ZN(
        P2_U3204) );
  NOR3_X1 U12496 ( .A1(n14960), .A2(n15107), .A3(n15090), .ZN(n9873) );
  INV_X1 U12497 ( .A(n15104), .ZN(n15082) );
  OR2_X1 U12498 ( .A1(n15109), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9865) );
  INV_X1 U12499 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n14239) );
  OAI22_X1 U12500 ( .A1(n9865), .A2(n9864), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14239), .ZN(n9869) );
  INV_X1 U12501 ( .A(n9866), .ZN(n9867) );
  INV_X1 U12502 ( .A(n15107), .ZN(n9914) );
  OAI22_X1 U12503 ( .A1(n15116), .A2(n9867), .B1(n9914), .B2(n9906), .ZN(n9868) );
  AOI211_X1 U12504 ( .C1(n15082), .C2(P3_ADDR_REG_0__SCAN_IN), .A(n9869), .B(
        n9868), .ZN(n9871) );
  NAND2_X1 U12505 ( .A1(n15000), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9870) );
  OAI211_X1 U12506 ( .C1(n9873), .C2(n9872), .A(n9871), .B(n9870), .ZN(
        P3_U3182) );
  NAND2_X1 U12507 ( .A1(n12559), .A2(n11836), .ZN(n12194) );
  INV_X1 U12508 ( .A(n12194), .ZN(n12198) );
  NOR2_X1 U12509 ( .A1(n12193), .A2(n12198), .ZN(n12368) );
  NAND3_X1 U12510 ( .A1(n9893), .A2(n15144), .A3(n9883), .ZN(n9876) );
  INV_X1 U12511 ( .A(n9884), .ZN(n9874) );
  NAND2_X1 U12512 ( .A1(n9896), .A2(n9874), .ZN(n9875) );
  NAND2_X1 U12513 ( .A1(n9876), .A2(n9875), .ZN(n9878) );
  INV_X1 U12514 ( .A(n9895), .ZN(n12413) );
  NAND2_X1 U12515 ( .A1(n12413), .A2(n9896), .ZN(n10050) );
  INV_X1 U12516 ( .A(n10049), .ZN(n9879) );
  INV_X1 U12517 ( .A(n12527), .ZN(n12503) );
  OR2_X1 U12518 ( .A1(n9893), .A2(n10603), .ZN(n9881) );
  AOI22_X1 U12519 ( .A1(n12557), .A2(n12503), .B1(n12515), .B2(n9882), .ZN(
        n9900) );
  INV_X1 U12520 ( .A(n9883), .ZN(n9892) );
  OR2_X1 U12521 ( .A1(n9896), .A2(n9884), .ZN(n9891) );
  INV_X1 U12522 ( .A(n9885), .ZN(n9887) );
  NOR2_X1 U12523 ( .A1(n9887), .A2(n9886), .ZN(n9888) );
  AND2_X1 U12524 ( .A1(n9889), .A2(n9888), .ZN(n9890) );
  OAI211_X1 U12525 ( .C1(n9893), .C2(n9892), .A(n9891), .B(n9890), .ZN(n9894)
         );
  NAND2_X1 U12526 ( .A1(n9894), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9898) );
  OR2_X1 U12527 ( .A1(n9896), .A2(n9895), .ZN(n9897) );
  NAND2_X1 U12528 ( .A1(n12461), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10104) );
  NAND2_X1 U12529 ( .A1(n10104), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9899) );
  OAI211_X1 U12530 ( .C1(n12368), .C2(n12534), .A(n9900), .B(n9899), .ZN(
        P3_U3172) );
  INV_X1 U12531 ( .A(n9901), .ZN(n9902) );
  MUX2_X1 U12532 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12646), .Z(n10518) );
  XOR2_X1 U12533 ( .A(n10521), .B(n10518), .Z(n9904) );
  NOR2_X1 U12534 ( .A1(n9905), .A2(n9904), .ZN(n10519) );
  AOI21_X1 U12535 ( .B1(n9905), .B2(n9904), .A(n10519), .ZN(n9922) );
  INV_X1 U12536 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n15161) );
  MUX2_X1 U12537 ( .A(P3_REG1_REG_2__SCAN_IN), .B(n15161), .S(n10521), .Z(
        n9911) );
  INV_X1 U12538 ( .A(n9906), .ZN(n9908) );
  AOI21_X1 U12539 ( .B1(n9909), .B2(n9908), .A(n9907), .ZN(n9910) );
  NOR2_X1 U12540 ( .A1(n9910), .A2(n9911), .ZN(n10544) );
  AOI21_X1 U12541 ( .B1(n9911), .B2(n9910), .A(n10544), .ZN(n9913) );
  AOI22_X1 U12542 ( .A1(n15082), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n9912) );
  OAI21_X1 U12543 ( .B1(n9914), .B2(n9913), .A(n9912), .ZN(n9920) );
  AOI21_X1 U12544 ( .B1(n9917), .B2(n9916), .A(n10531), .ZN(n9918) );
  NOR2_X1 U12545 ( .A1(n15116), .A2(n9918), .ZN(n9919) );
  AOI211_X1 U12546 ( .C1(n15000), .C2(n10521), .A(n9920), .B(n9919), .ZN(n9921) );
  OAI21_X1 U12547 ( .B1(n9922), .B2(n15109), .A(n9921), .ZN(P3_U3184) );
  INV_X1 U12548 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9939) );
  NAND2_X1 U12549 ( .A1(n10267), .A2(n10093), .ZN(n9923) );
  INV_X1 U12550 ( .A(n9925), .ZN(n9930) );
  OAI21_X1 U12551 ( .B1(n9926), .B2(n9930), .A(n10015), .ZN(n9935) );
  INV_X1 U12552 ( .A(n9935), .ZN(n10281) );
  OAI22_X1 U12553 ( .A1(n10288), .A2(n13052), .B1(n10093), .B2(n13051), .ZN(
        n9934) );
  AND2_X1 U12554 ( .A1(n9973), .A2(n10093), .ZN(n9927) );
  NAND2_X1 U12555 ( .A1(n10267), .A2(n13092), .ZN(n9929) );
  NAND2_X1 U12556 ( .A1(n9931), .A2(n9930), .ZN(n9932) );
  AOI21_X1 U12557 ( .B1(n10020), .B2(n9932), .A(n13294), .ZN(n9933) );
  AOI211_X1 U12558 ( .C1(n10401), .C2(n9935), .A(n9934), .B(n9933), .ZN(n10273) );
  AOI21_X1 U12559 ( .B1(n10274), .B2(n9936), .A(n10017), .ZN(n10278) );
  AOI22_X1 U12560 ( .A1(n10278), .A2(n13505), .B1(n13513), .B2(n10274), .ZN(
        n9937) );
  OAI211_X1 U12561 ( .C1(n10281), .C2(n10420), .A(n10273), .B(n9937), .ZN(
        n13519) );
  NAND2_X1 U12562 ( .A1(n13519), .A2(n6443), .ZN(n9938) );
  OAI21_X1 U12563 ( .B1(n6443), .B2(n9939), .A(n9938), .ZN(P2_U3448) );
  INV_X1 U12564 ( .A(n9940), .ZN(n9949) );
  OAI22_X1 U12565 ( .A1(n14515), .A2(n9942), .B1(n9941), .B2(n13066), .ZN(
        n9948) );
  AOI22_X1 U12566 ( .A1(n13040), .A2(n13097), .B1(n14523), .B2(n9943), .ZN(
        n9946) );
  INV_X1 U12567 ( .A(n9944), .ZN(n9945) );
  AOI211_X1 U12568 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(n9949), .A(n9948), .B(
        n9947), .ZN(n9950) );
  OAI21_X1 U12569 ( .B1(n9951), .B2(n14502), .A(n9950), .ZN(P2_U3209) );
  OAI21_X1 U12570 ( .B1(n9748), .B2(n9953), .A(n9952), .ZN(n9956) );
  INV_X1 U12571 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9954) );
  MUX2_X1 U12572 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n9954), .S(n10726), .Z(n9955) );
  AND2_X1 U12573 ( .A1(n9956), .A2(n9955), .ZN(n10352) );
  OAI21_X1 U12574 ( .B1(n9956), .B2(n9955), .A(n14633), .ZN(n9965) );
  INV_X1 U12575 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10729) );
  MUX2_X1 U12576 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10729), .S(n10726), .Z(
        n9959) );
  OAI21_X1 U12577 ( .B1(n10749), .B2(P1_REG1_REG_8__SCAN_IN), .A(n9957), .ZN(
        n9958) );
  NAND2_X1 U12578 ( .A1(n9958), .A2(n9959), .ZN(n10348) );
  OAI21_X1 U12579 ( .B1(n9959), .B2(n9958), .A(n10348), .ZN(n9960) );
  NAND2_X1 U12580 ( .A1(n9960), .A2(n14636), .ZN(n9964) );
  AND2_X1 U12581 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n10985) );
  NOR2_X1 U12582 ( .A1(n14618), .A2(n9961), .ZN(n9962) );
  AOI211_X1 U12583 ( .C1(n14585), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n10985), .B(
        n9962), .ZN(n9963) );
  OAI211_X1 U12584 ( .C1(n10352), .C2(n9965), .A(n9964), .B(n9963), .ZN(
        P1_U3252) );
  INV_X1 U12585 ( .A(n9966), .ZN(n9967) );
  OAI222_X1 U12586 ( .A1(P3_U3151), .A2(n6743), .B1(n12933), .B2(n9968), .C1(
        n11500), .C2(n9967), .ZN(P3_U3277) );
  AOI22_X1 U12587 ( .A1(n13040), .A2(n13093), .B1(n14523), .B2(n9969), .ZN(
        n9971) );
  NOR2_X1 U12588 ( .A1(n9971), .A2(n9970), .ZN(n9977) );
  OAI22_X1 U12589 ( .A1(n9972), .A2(n14519), .B1(n14518), .B2(n10035), .ZN(
        n9976) );
  NAND2_X1 U12590 ( .A1(n14507), .A2(n9973), .ZN(n9974) );
  NAND2_X1 U12591 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n13119) );
  OAI211_X1 U12592 ( .C1(n14528), .C2(n10266), .A(n9974), .B(n13119), .ZN(
        n9975) );
  AOI211_X1 U12593 ( .C1(n9977), .C2(n9988), .A(n9976), .B(n9975), .ZN(n9978)
         );
  OAI21_X1 U12594 ( .B1(n9979), .B2(n14502), .A(n9978), .ZN(P2_U3199) );
  INV_X1 U12595 ( .A(n10069), .ZN(n9987) );
  AND2_X1 U12596 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n14845) );
  AOI21_X1 U12597 ( .B1(n14507), .B2(n10073), .A(n14845), .ZN(n9980) );
  OAI21_X1 U12598 ( .B1(n14518), .B2(n10093), .A(n9980), .ZN(n9986) );
  INV_X1 U12599 ( .A(n9989), .ZN(n9982) );
  NAND3_X1 U12600 ( .A1(n13040), .A2(n9982), .A3(n9981), .ZN(n9984) );
  AOI21_X1 U12601 ( .B1(n9984), .B2(n14519), .A(n9983), .ZN(n9985) );
  AOI211_X1 U12602 ( .C1(n13036), .C2(n9987), .A(n9986), .B(n9985), .ZN(n9993)
         );
  OAI21_X1 U12603 ( .B1(n9990), .B2(n9989), .A(n9988), .ZN(n9991) );
  NAND2_X1 U12604 ( .A1(n9991), .A2(n14523), .ZN(n9992) );
  NAND2_X1 U12605 ( .A1(n9993), .A2(n9992), .ZN(P2_U3202) );
  NOR2_X1 U12606 ( .A1(n9995), .A2(n9994), .ZN(n9997) );
  NAND2_X1 U12607 ( .A1(n9997), .A2(n9996), .ZN(n10003) );
  INV_X2 U12608 ( .A(n13426), .ZN(n13394) );
  AND2_X1 U12609 ( .A1(n9999), .A2(n9998), .ZN(n10000) );
  NAND2_X1 U12610 ( .A1(n13394), .A2(n10000), .ZN(n10438) );
  INV_X1 U12611 ( .A(n10001), .ZN(n10002) );
  NOR2_X1 U12612 ( .A1(n10003), .A2(n8050), .ZN(n13385) );
  INV_X1 U12613 ( .A(n13385), .ZN(n10071) );
  OAI22_X1 U12614 ( .A1(n10071), .A2(n10004), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n13377), .ZN(n10005) );
  AOI21_X1 U12615 ( .B1(n13381), .B2(n10006), .A(n10005), .ZN(n10009) );
  MUX2_X1 U12616 ( .A(n9552), .B(n10007), .S(n13394), .Z(n10008) );
  OAI211_X1 U12617 ( .C1(n10010), .C2(n10438), .A(n10009), .B(n10008), .ZN(
        P2_U3262) );
  INV_X1 U12618 ( .A(n10011), .ZN(n10013) );
  OAI222_X1 U12619 ( .A1(n11500), .A2(n10013), .B1(n12933), .B2(n10012), .C1(
        P3_U3151), .C2(n12654), .ZN(P3_U3276) );
  OR2_X1 U12620 ( .A1(n10274), .A2(n13091), .ZN(n10014) );
  OAI21_X1 U12621 ( .B1(n10016), .B2(n10021), .A(n10283), .ZN(n10262) );
  INV_X1 U12622 ( .A(n10289), .ZN(n10018) );
  OAI211_X1 U12623 ( .C1(n10018), .C2(n10017), .A(n13505), .B(n10295), .ZN(
        n10258) );
  OAI21_X1 U12624 ( .B1(n10018), .B2(n14922), .A(n10258), .ZN(n10026) );
  NAND2_X1 U12625 ( .A1(n10274), .A2(n10035), .ZN(n10019) );
  INV_X1 U12626 ( .A(n10021), .ZN(n10022) );
  OAI211_X1 U12627 ( .C1(n10023), .C2(n10022), .A(n10291), .B(n13406), .ZN(
        n10025) );
  AOI22_X1 U12628 ( .A1(n13370), .A2(n13091), .B1(n13089), .B2(n13372), .ZN(
        n10024) );
  NAND2_X1 U12629 ( .A1(n10025), .A2(n10024), .ZN(n10259) );
  AOI211_X1 U12630 ( .C1(n14533), .C2(n10262), .A(n10026), .B(n10259), .ZN(
        n10112) );
  NAND2_X1 U12631 ( .A1(n14931), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10027) );
  OAI21_X1 U12632 ( .B1(n10112), .B2(n14931), .A(n10027), .ZN(P2_U3506) );
  INV_X1 U12633 ( .A(n10028), .ZN(n10029) );
  AOI21_X1 U12634 ( .B1(n10089), .B2(n10029), .A(n14502), .ZN(n10033) );
  NOR3_X1 U12635 ( .A1(n12977), .A2(n10030), .A3(n10035), .ZN(n10032) );
  OAI21_X1 U12636 ( .B1(n10033), .B2(n10032), .A(n10031), .ZN(n10039) );
  INV_X1 U12637 ( .A(n13089), .ZN(n10393) );
  OAI21_X1 U12638 ( .B1(n14518), .B2(n10393), .A(n10034), .ZN(n10037) );
  OAI22_X1 U12639 ( .A1(n14519), .A2(n10035), .B1(n14528), .B2(n10255), .ZN(
        n10036) );
  AOI211_X1 U12640 ( .C1(n10289), .C2(n14507), .A(n10037), .B(n10036), .ZN(
        n10038) );
  NAND2_X1 U12641 ( .A1(n10039), .A2(n10038), .ZN(P2_U3185) );
  INV_X1 U12642 ( .A(n10604), .ZN(n10048) );
  INV_X1 U12643 ( .A(n10043), .ZN(n12199) );
  NOR3_X1 U12644 ( .A1(n12199), .A2(n12153), .A3(n12193), .ZN(n10046) );
  NAND2_X1 U12645 ( .A1(n10604), .A2(n12153), .ZN(n10044) );
  AOI21_X1 U12646 ( .B1(n10045), .B2(n10044), .A(n10047), .ZN(n10100) );
  AOI211_X1 U12647 ( .C1(n10048), .C2(n10047), .A(n10046), .B(n10100), .ZN(
        n10056) );
  INV_X1 U12648 ( .A(n10051), .ZN(n10455) );
  OAI22_X1 U12649 ( .A1(n10455), .A2(n12527), .B1(n10052), .B2(n12528), .ZN(
        n10053) );
  AOI21_X1 U12650 ( .B1(n12525), .B2(n12559), .A(n10053), .ZN(n10055) );
  NAND2_X1 U12651 ( .A1(n10104), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n10054) );
  OAI211_X1 U12652 ( .C1(n10056), .C2(n12534), .A(n10055), .B(n10054), .ZN(
        P3_U3162) );
  NAND2_X1 U12653 ( .A1(n9458), .A2(n13226), .ZN(n10057) );
  AND2_X1 U12654 ( .A1(n8086), .A2(n10057), .ZN(n10058) );
  INV_X1 U12655 ( .A(n10059), .ZN(n10067) );
  INV_X1 U12656 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10060) );
  OAI22_X1 U12657 ( .A1(n13394), .A2(n10061), .B1(n10060), .B2(n13377), .ZN(
        n10062) );
  AOI21_X1 U12658 ( .B1(n13381), .B2(n8319), .A(n10062), .ZN(n10066) );
  AOI22_X1 U12659 ( .A1(n13424), .A2(n10064), .B1(n13394), .B2(n10063), .ZN(
        n10065) );
  OAI211_X1 U12660 ( .C1(n13421), .C2(n10067), .A(n10066), .B(n10065), .ZN(
        P2_U3263) );
  INV_X1 U12661 ( .A(n10068), .ZN(n10078) );
  OAI22_X1 U12662 ( .A1(n10071), .A2(n10070), .B1(n10069), .B2(n13377), .ZN(
        n10072) );
  AOI21_X1 U12663 ( .B1(n13381), .B2(n10073), .A(n10072), .ZN(n10077) );
  INV_X1 U12664 ( .A(n10074), .ZN(n10075) );
  MUX2_X1 U12665 ( .A(n9553), .B(n10075), .S(n13394), .Z(n10076) );
  OAI211_X1 U12666 ( .C1(n10078), .C2(n13421), .A(n10077), .B(n10076), .ZN(
        P2_U3261) );
  INV_X1 U12667 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n10079) );
  NAND3_X1 U12668 ( .A1(n10081), .A2(n10080), .A3(n10079), .ZN(n10082) );
  OAI21_X1 U12669 ( .B1(n10083), .B2(n10082), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n10085) );
  INV_X1 U12670 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n10084) );
  XNOR2_X1 U12671 ( .A(n10085), .B(n10084), .ZN(n13786) );
  INV_X1 U12672 ( .A(n11285), .ZN(n10088) );
  OAI222_X1 U12673 ( .A1(P1_U3086), .A2(n13786), .B1(n14375), .B2(n10088), 
        .C1(n10086), .C2(n14372), .ZN(P1_U3340) );
  INV_X1 U12674 ( .A(n13168), .ZN(n13161) );
  OAI222_X1 U12675 ( .A1(P2_U3088), .A2(n13161), .B1(n13549), .B2(n10088), 
        .C1(n10087), .C2(n13551), .ZN(P2_U3312) );
  INV_X1 U12676 ( .A(n10089), .ZN(n10090) );
  AOI211_X1 U12677 ( .C1(n10092), .C2(n10091), .A(n14502), .B(n10090), .ZN(
        n10097) );
  OAI22_X1 U12678 ( .A1(n10288), .A2(n14518), .B1(n14519), .B2(n10093), .ZN(
        n10096) );
  NAND2_X1 U12679 ( .A1(n14507), .A2(n10274), .ZN(n10094) );
  NAND2_X1 U12680 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n13134) );
  OAI211_X1 U12681 ( .C1(n14528), .C2(n10275), .A(n10094), .B(n13134), .ZN(
        n10095) );
  OR3_X1 U12682 ( .A1(n10097), .A2(n10096), .A3(n10095), .ZN(P2_U3211) );
  XNOR2_X1 U12683 ( .A(n15129), .B(n10448), .ZN(n10449) );
  XNOR2_X1 U12684 ( .A(n10449), .B(n10051), .ZN(n10450) );
  INV_X1 U12685 ( .A(n10098), .ZN(n10099) );
  NOR2_X1 U12686 ( .A1(n10100), .A2(n10099), .ZN(n10451) );
  XOR2_X1 U12687 ( .A(n10450), .B(n10451), .Z(n10106) );
  AOI22_X1 U12688 ( .A1(n12556), .A2(n12503), .B1(n12515), .B2(n10101), .ZN(
        n10102) );
  OAI21_X1 U12689 ( .B1(n9097), .B2(n12505), .A(n10102), .ZN(n10103) );
  AOI21_X1 U12690 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n10104), .A(n10103), .ZN(
        n10105) );
  OAI21_X1 U12691 ( .B1(n10106), .B2(n12534), .A(n10105), .ZN(P3_U3177) );
  OR3_X1 U12692 ( .A1(n12368), .A2(n15152), .A3(n10107), .ZN(n10108) );
  OAI21_X1 U12693 ( .B1(n9097), .B2(n15122), .A(n10108), .ZN(n11832) );
  INV_X1 U12694 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10109) );
  OAI22_X1 U12695 ( .A1(n11836), .A2(n12926), .B1(n15158), .B2(n10109), .ZN(
        n10110) );
  AOI21_X1 U12696 ( .B1(n11832), .B2(n15158), .A(n10110), .ZN(n10111) );
  INV_X1 U12697 ( .A(n10111), .ZN(P3_U3390) );
  INV_X1 U12698 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10114) );
  OR2_X1 U12699 ( .A1(n10112), .A2(n14928), .ZN(n10113) );
  OAI21_X1 U12700 ( .B1(n6443), .B2(n10114), .A(n10113), .ZN(P2_U3451) );
  INV_X1 U12701 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10115) );
  MUX2_X1 U12702 ( .A(n10115), .B(P2_REG1_REG_10__SCAN_IN), .S(n10373), .Z(
        n10118) );
  OAI21_X1 U12703 ( .B1(n10120), .B2(P2_REG1_REG_9__SCAN_IN), .A(n10116), .ZN(
        n10117) );
  NOR2_X1 U12704 ( .A1(n10117), .A2(n10118), .ZN(n10372) );
  AOI211_X1 U12705 ( .C1(n10118), .C2(n10117), .A(n14856), .B(n10372), .ZN(
        n10129) );
  OAI21_X1 U12706 ( .B1(n10120), .B2(P2_REG2_REG_9__SCAN_IN), .A(n10119), .ZN(
        n10123) );
  INV_X1 U12707 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10121) );
  MUX2_X1 U12708 ( .A(n10121), .B(P2_REG2_REG_10__SCAN_IN), .S(n10373), .Z(
        n10122) );
  NOR2_X1 U12709 ( .A1(n10123), .A2(n10122), .ZN(n10363) );
  AOI211_X1 U12710 ( .C1(n10123), .C2(n10122), .A(n14864), .B(n10363), .ZN(
        n10128) );
  NAND2_X1 U12711 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n12958)
         );
  INV_X1 U12712 ( .A(n12958), .ZN(n10124) );
  AOI21_X1 U12713 ( .B1(n14840), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n10124), 
        .ZN(n10125) );
  OAI21_X1 U12714 ( .B1(n13184), .B2(n10126), .A(n10125), .ZN(n10127) );
  OR3_X1 U12715 ( .A1(n10129), .A2(n10128), .A3(n10127), .ZN(P2_U3224) );
  NAND2_X1 U12716 ( .A1(n11845), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10134) );
  OR2_X1 U12717 ( .A1(n11839), .A2(n14326), .ZN(n10133) );
  NAND2_X1 U12718 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n10172) );
  OAI21_X1 U12719 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n10172), .ZN(n10188) );
  OR2_X1 U12720 ( .A1(n9605), .A2(n10188), .ZN(n10132) );
  INV_X1 U12721 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10130) );
  OR2_X1 U12722 ( .A1(n11816), .A2(n10130), .ZN(n10131) );
  NAND2_X1 U12723 ( .A1(n12022), .A2(n10136), .ZN(n10139) );
  OR2_X1 U12724 ( .A1(n12023), .A2(n10137), .ZN(n10138) );
  AOI22_X1 U12725 ( .A1(n13697), .A2(n11775), .B1(n11807), .B2(n11895), .ZN(
        n10141) );
  XOR2_X1 U12726 ( .A(n10326), .B(n10141), .Z(n10168) );
  INV_X1 U12727 ( .A(n10142), .ZN(n10143) );
  NAND2_X1 U12728 ( .A1(n10144), .A2(n10143), .ZN(n10145) );
  INV_X1 U12729 ( .A(n13578), .ZN(n10157) );
  OR2_X1 U12730 ( .A1(n12023), .A2(n10147), .ZN(n10150) );
  OR2_X1 U12731 ( .A1(n11610), .A2(n10148), .ZN(n10149) );
  OAI22_X1 U12732 ( .A1(n10687), .A2(n10161), .B1(n14773), .B2(n9766), .ZN(
        n10152) );
  XNOR2_X1 U12733 ( .A(n10152), .B(n10326), .ZN(n10159) );
  OR2_X1 U12734 ( .A1(n10687), .A2(n10153), .ZN(n10155) );
  NAND2_X1 U12735 ( .A1(n14753), .A2(n11775), .ZN(n10154) );
  NAND2_X1 U12736 ( .A1(n10155), .A2(n10154), .ZN(n10158) );
  XNOR2_X1 U12737 ( .A(n10159), .B(n10158), .ZN(n13577) );
  NAND2_X1 U12738 ( .A1(n10159), .A2(n10158), .ZN(n10160) );
  AOI22_X1 U12739 ( .A1(n13697), .A2(n11808), .B1(n11775), .B2(n11895), .ZN(
        n10163) );
  INV_X1 U12740 ( .A(n10163), .ZN(n10164) );
  AOI21_X1 U12741 ( .B1(n10168), .B2(n10167), .A(n6596), .ZN(n10194) );
  NAND2_X1 U12742 ( .A1(n11846), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n10177) );
  OR2_X1 U12743 ( .A1(n11818), .A2(n10169), .ZN(n10176) );
  OR2_X1 U12744 ( .A1(n11839), .A2(n10170), .ZN(n10175) );
  AND2_X1 U12745 ( .A1(n10172), .A2(n10171), .ZN(n10173) );
  OR2_X1 U12746 ( .A1(n10173), .A2(n10233), .ZN(n14732) );
  OR2_X1 U12747 ( .A1(n9605), .A2(n14732), .ZN(n10174) );
  NAND4_X1 U12748 ( .A1(n10177), .A2(n10176), .A3(n10175), .A4(n10174), .ZN(
        n13696) );
  NAND2_X1 U12749 ( .A1(n6433), .A2(n13696), .ZN(n10191) );
  NAND2_X1 U12750 ( .A1(n10639), .A2(n10178), .ZN(n10179) );
  NAND2_X1 U12751 ( .A1(n10180), .A2(n10179), .ZN(n10186) );
  NAND2_X1 U12752 ( .A1(n10182), .A2(n10181), .ZN(n10183) );
  NOR2_X1 U12753 ( .A1(n10184), .A2(n10183), .ZN(n10185) );
  NAND2_X1 U12754 ( .A1(n10186), .A2(n10185), .ZN(n10187) );
  INV_X1 U12755 ( .A(n10188), .ZN(n10663) );
  AOI21_X1 U12756 ( .B1(n13664), .B2(n10663), .A(n10189), .ZN(n10190) );
  OAI211_X1 U12757 ( .C1(n10687), .C2(n13667), .A(n10191), .B(n10190), .ZN(
        n10192) );
  AOI21_X1 U12758 ( .B1(n13685), .B2(n11895), .A(n10192), .ZN(n10193) );
  OAI21_X1 U12759 ( .B1(n10194), .B2(n13688), .A(n10193), .ZN(P1_U3230) );
  INV_X1 U12760 ( .A(n10195), .ZN(n10198) );
  OAI222_X1 U12761 ( .A1(n11500), .A2(n10198), .B1(n12933), .B2(n10197), .C1(
        P3_U3151), .C2(n10196), .ZN(P3_U3275) );
  OAI21_X1 U12762 ( .B1(n14519), .B2(n10393), .A(n10199), .ZN(n10201) );
  INV_X1 U12763 ( .A(n13087), .ZN(n10476) );
  OAI22_X1 U12764 ( .A1(n14518), .A2(n10476), .B1(n14528), .B2(n10404), .ZN(
        n10200) );
  AOI211_X1 U12765 ( .C1(n10424), .C2(n14507), .A(n10201), .B(n10200), .ZN(
        n10207) );
  INV_X1 U12766 ( .A(n10202), .ZN(n10205) );
  OAI22_X1 U12767 ( .A1(n12977), .A2(n10393), .B1(n10203), .B2(n14502), .ZN(
        n10204) );
  NAND3_X1 U12768 ( .A1(n12968), .A2(n10205), .A3(n10204), .ZN(n10206) );
  OAI211_X1 U12769 ( .C1(n10208), .C2(n14502), .A(n10207), .B(n10206), .ZN(
        P2_U3203) );
  INV_X1 U12770 ( .A(n10209), .ZN(n10210) );
  NAND2_X1 U12771 ( .A1(n10211), .A2(n10210), .ZN(n10213) );
  NAND2_X1 U12772 ( .A1(n10213), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10212) );
  MUX2_X1 U12773 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10212), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n10214) );
  OR2_X1 U12774 ( .A1(n10213), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n10310) );
  AND2_X1 U12775 ( .A1(n10214), .A2(n10310), .ZN(n14649) );
  INV_X1 U12776 ( .A(n14649), .ZN(n10216) );
  INV_X1 U12777 ( .A(n11342), .ZN(n10218) );
  OAI222_X1 U12778 ( .A1(P1_U3086), .A2(n10216), .B1(n14375), .B2(n10218), 
        .C1(n10215), .C2(n14372), .ZN(P1_U3339) );
  INV_X1 U12779 ( .A(n13172), .ZN(n13189) );
  OAI222_X1 U12780 ( .A1(P2_U3088), .A2(n13189), .B1(n13549), .B2(n10218), 
        .C1(n10217), .C2(n13551), .ZN(P2_U3311) );
  NAND2_X1 U12781 ( .A1(n13696), .A2(n11775), .ZN(n10224) );
  AOI22_X1 U12782 ( .A1(n11627), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n11626), 
        .B2(n13734), .ZN(n10222) );
  OR2_X1 U12783 ( .A1(n10220), .A2(n11610), .ZN(n10221) );
  NAND2_X1 U12784 ( .A1(n10222), .A2(n10221), .ZN(n14734) );
  NAND2_X1 U12785 ( .A1(n14734), .A2(n11807), .ZN(n10223) );
  NAND2_X1 U12786 ( .A1(n10224), .A2(n10223), .ZN(n10226) );
  XNOR2_X1 U12787 ( .A(n10226), .B(n10225), .ZN(n10227) );
  AOI22_X1 U12788 ( .A1(n13696), .A2(n11808), .B1(n14734), .B2(n11775), .ZN(
        n10228) );
  AND2_X1 U12789 ( .A1(n10227), .A2(n10228), .ZN(n10318) );
  INV_X1 U12790 ( .A(n10318), .ZN(n10231) );
  INV_X1 U12791 ( .A(n10227), .ZN(n10230) );
  INV_X1 U12792 ( .A(n10228), .ZN(n10229) );
  NAND2_X1 U12793 ( .A1(n10230), .A2(n10229), .ZN(n10317) );
  NAND2_X1 U12794 ( .A1(n10231), .A2(n10317), .ZN(n10232) );
  XNOR2_X1 U12795 ( .A(n10319), .B(n10232), .ZN(n10245) );
  NAND2_X1 U12796 ( .A1(n11845), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10239) );
  OR2_X1 U12797 ( .A1(n11839), .A2(n9488), .ZN(n10238) );
  NAND2_X1 U12798 ( .A1(n10233), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10333) );
  OR2_X1 U12799 ( .A1(n10233), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10234) );
  NAND2_X1 U12800 ( .A1(n10333), .A2(n10234), .ZN(n10802) );
  OR2_X1 U12801 ( .A1(n9605), .A2(n10802), .ZN(n10237) );
  INV_X1 U12802 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10235) );
  OR2_X1 U12803 ( .A1(n11816), .A2(n10235), .ZN(n10236) );
  NAND4_X1 U12804 ( .A1(n10239), .A2(n10238), .A3(n10237), .A4(n10236), .ZN(
        n14704) );
  NAND2_X1 U12805 ( .A1(n6433), .A2(n14704), .ZN(n10242) );
  INV_X1 U12806 ( .A(n14732), .ZN(n10240) );
  AND2_X1 U12807 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n13733) );
  AOI21_X1 U12808 ( .B1(n13664), .B2(n10240), .A(n13733), .ZN(n10241) );
  OAI211_X1 U12809 ( .C1(n14723), .C2(n13667), .A(n10242), .B(n10241), .ZN(
        n10243) );
  AOI21_X1 U12810 ( .B1(n13685), .B2(n14734), .A(n10243), .ZN(n10244) );
  OAI21_X1 U12811 ( .B1(n10245), .B2(n13688), .A(n10244), .ZN(P1_U3227) );
  NAND2_X1 U12812 ( .A1(n13394), .A2(n10246), .ZN(n10247) );
  OAI21_X1 U12813 ( .B1(n13377), .B2(n10248), .A(n10247), .ZN(n10251) );
  NOR2_X1 U12814 ( .A1(n10438), .A2(n10249), .ZN(n10250) );
  AOI211_X1 U12815 ( .C1(n13426), .C2(P2_REG2_REG_0__SCAN_IN), .A(n10251), .B(
        n10250), .ZN(n10254) );
  OAI21_X1 U12816 ( .B1(n13381), .B2(n13385), .A(n10252), .ZN(n10253) );
  NAND2_X1 U12817 ( .A1(n10254), .A2(n10253), .ZN(P2_U3265) );
  INV_X1 U12818 ( .A(n13421), .ZN(n13272) );
  INV_X1 U12819 ( .A(n13377), .ZN(n13412) );
  INV_X1 U12820 ( .A(n10255), .ZN(n10256) );
  AOI22_X1 U12821 ( .A1(n13381), .A2(n10289), .B1(n13412), .B2(n10256), .ZN(
        n10257) );
  OAI21_X1 U12822 ( .B1(n13325), .B2(n10258), .A(n10257), .ZN(n10261) );
  MUX2_X1 U12823 ( .A(n10259), .B(P2_REG2_REG_7__SCAN_IN), .S(n13426), .Z(
        n10260) );
  AOI211_X1 U12824 ( .C1(n13272), .C2(n10262), .A(n10261), .B(n10260), .ZN(
        n10263) );
  INV_X1 U12825 ( .A(n10263), .ZN(P2_U3258) );
  MUX2_X1 U12826 ( .A(n10265), .B(n10264), .S(n13394), .Z(n10271) );
  OAI22_X1 U12827 ( .A1(n13415), .A2(n10267), .B1(n13377), .B2(n10266), .ZN(
        n10268) );
  AOI21_X1 U12828 ( .B1(n13424), .B2(n10269), .A(n10268), .ZN(n10270) );
  OAI211_X1 U12829 ( .C1(n10272), .C2(n10438), .A(n10271), .B(n10270), .ZN(
        P2_U3260) );
  MUX2_X1 U12830 ( .A(n14230), .B(n10273), .S(n13394), .Z(n10280) );
  INV_X1 U12831 ( .A(n10274), .ZN(n10276) );
  OAI22_X1 U12832 ( .A1(n13415), .A2(n10276), .B1(n13377), .B2(n10275), .ZN(
        n10277) );
  AOI21_X1 U12833 ( .B1(n13385), .B2(n10278), .A(n10277), .ZN(n10279) );
  OAI211_X1 U12834 ( .C1(n10281), .C2(n10438), .A(n10280), .B(n10279), .ZN(
        P2_U3259) );
  OR2_X1 U12835 ( .A1(n10289), .A2(n13090), .ZN(n10282) );
  NAND2_X1 U12836 ( .A1(n10286), .A2(n10391), .ZN(n10287) );
  NAND2_X1 U12837 ( .A1(n10390), .A2(n10287), .ZN(n14914) );
  AOI22_X1 U12838 ( .A1(n13370), .A2(n13090), .B1(n13088), .B2(n13372), .ZN(
        n10294) );
  OR2_X1 U12839 ( .A1(n10289), .A2(n10288), .ZN(n10290) );
  NAND2_X1 U12840 ( .A1(n10291), .A2(n10290), .ZN(n10392) );
  XOR2_X1 U12841 ( .A(n10392), .B(n10391), .Z(n10292) );
  NAND2_X1 U12842 ( .A1(n10292), .A2(n13406), .ZN(n10293) );
  OAI211_X1 U12843 ( .C1(n14914), .C2(n9458), .A(n10294), .B(n10293), .ZN(
        n14916) );
  NAND2_X1 U12844 ( .A1(n14916), .A2(n13394), .ZN(n10299) );
  OAI22_X1 U12845 ( .A1(n13394), .A2(n14242), .B1(n12970), .B2(n13377), .ZN(
        n10297) );
  OAI211_X1 U12846 ( .C1(n7130), .C2(n7131), .A(n13505), .B(n10402), .ZN(
        n14915) );
  NOR2_X1 U12847 ( .A1(n14915), .A2(n13325), .ZN(n10296) );
  AOI211_X1 U12848 ( .C1(n13381), .C2(n12975), .A(n10297), .B(n10296), .ZN(
        n10298) );
  OAI211_X1 U12849 ( .C1(n14914), .C2(n10438), .A(n10299), .B(n10298), .ZN(
        P2_U3257) );
  OAI21_X1 U12850 ( .B1(n10301), .B2(n12367), .A(n10300), .ZN(n10599) );
  OAI211_X1 U12851 ( .C1(n10304), .C2(n10303), .A(n12766), .B(n10302), .ZN(
        n10306) );
  INV_X1 U12852 ( .A(n12799), .ZN(n11219) );
  AOI22_X1 U12853 ( .A1(n12555), .A2(n12769), .B1(n11219), .B2(n10051), .ZN(
        n10305) );
  NAND2_X1 U12854 ( .A1(n10306), .A2(n10305), .ZN(n10582) );
  AOI21_X1 U12855 ( .B1(n15150), .B2(n10599), .A(n10582), .ZN(n10465) );
  INV_X1 U12856 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n10307) );
  OAI22_X1 U12857 ( .A1(n10462), .A2(n12926), .B1(n15158), .B2(n10307), .ZN(
        n10308) );
  INV_X1 U12858 ( .A(n10308), .ZN(n10309) );
  OAI21_X1 U12859 ( .B1(n10465), .B2(n15157), .A(n10309), .ZN(P3_U3399) );
  NAND2_X1 U12860 ( .A1(n10310), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10311) );
  MUX2_X1 U12861 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10311), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n10313) );
  NAND2_X1 U12862 ( .A1(n10313), .A2(n10312), .ZN(n13789) );
  INV_X1 U12863 ( .A(n11601), .ZN(n10316) );
  OAI222_X1 U12864 ( .A1(P1_U3086), .A2(n13789), .B1(n14375), .B2(n10316), 
        .C1(n10314), .C2(n14372), .ZN(P1_U3338) );
  OAI222_X1 U12865 ( .A1(P2_U3088), .A2(n13198), .B1(n13549), .B2(n10316), 
        .C1(n10315), .C2(n13551), .ZN(P2_U3310) );
  OR2_X1 U12866 ( .A1(n10320), .A2(n11610), .ZN(n10323) );
  AOI22_X1 U12867 ( .A1(n11627), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n11626), 
        .B2(n10321), .ZN(n10322) );
  NAND2_X1 U12868 ( .A1(n10323), .A2(n10322), .ZN(n14793) );
  NAND2_X1 U12869 ( .A1(n14793), .A2(n11807), .ZN(n10325) );
  NAND2_X1 U12870 ( .A1(n14704), .A2(n11775), .ZN(n10324) );
  NAND2_X1 U12871 ( .A1(n10325), .A2(n10324), .ZN(n10327) );
  XNOR2_X1 U12872 ( .A(n10327), .B(n10326), .ZN(n10564) );
  AOI22_X1 U12873 ( .A1(n14793), .A2(n11775), .B1(n11808), .B2(n14704), .ZN(
        n10565) );
  XNOR2_X1 U12874 ( .A(n10564), .B(n10565), .ZN(n10329) );
  NAND2_X1 U12875 ( .A1(n10330), .A2(n10329), .ZN(n10568) );
  OAI211_X1 U12876 ( .C1(n10330), .C2(n10329), .A(n10568), .B(n13645), .ZN(
        n10347) );
  NAND2_X1 U12877 ( .A1(n11845), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10339) );
  OR2_X1 U12878 ( .A1(n11839), .A2(n10331), .ZN(n10338) );
  INV_X1 U12879 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10332) );
  NAND2_X1 U12880 ( .A1(n10333), .A2(n10332), .ZN(n10334) );
  NAND2_X1 U12881 ( .A1(n10732), .A2(n10334), .ZN(n14709) );
  OR2_X1 U12882 ( .A1(n9605), .A2(n14709), .ZN(n10337) );
  INV_X1 U12883 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10335) );
  OR2_X1 U12884 ( .A1(n11816), .A2(n10335), .ZN(n10336) );
  NAND4_X1 U12885 ( .A1(n10339), .A2(n10338), .A3(n10337), .A4(n10336), .ZN(
        n14682) );
  NAND2_X1 U12886 ( .A1(n6433), .A2(n14682), .ZN(n10344) );
  INV_X1 U12887 ( .A(n10802), .ZN(n10342) );
  INV_X1 U12888 ( .A(n10340), .ZN(n10341) );
  AOI21_X1 U12889 ( .B1(n13664), .B2(n10342), .A(n10341), .ZN(n10343) );
  OAI211_X1 U12890 ( .C1(n10793), .C2(n13667), .A(n10344), .B(n10343), .ZN(
        n10345) );
  AOI21_X1 U12891 ( .B1(n13685), .B2(n14793), .A(n10345), .ZN(n10346) );
  NAND2_X1 U12892 ( .A1(n10347), .A2(n10346), .ZN(P1_U3239) );
  OAI21_X1 U12893 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n10726), .A(n10348), .ZN(
        n14593) );
  INV_X1 U12894 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10349) );
  MUX2_X1 U12895 ( .A(n10349), .B(P1_REG1_REG_10__SCAN_IN), .S(n14597), .Z(
        n14594) );
  NOR2_X1 U12896 ( .A1(n14593), .A2(n14594), .ZN(n14592) );
  INV_X1 U12897 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10851) );
  MUX2_X1 U12898 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10851), .S(n13762), .Z(
        n10350) );
  OAI21_X1 U12899 ( .B1(n10351), .B2(n10350), .A(n13756), .ZN(n10361) );
  INV_X1 U12900 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10353) );
  MUX2_X1 U12901 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10353), .S(n14597), .Z(
        n10354) );
  INV_X1 U12902 ( .A(n10354), .ZN(n14590) );
  NOR2_X1 U12903 ( .A1(n14591), .A2(n14590), .ZN(n14589) );
  AOI21_X1 U12904 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n14597), .A(n14589), 
        .ZN(n10356) );
  XNOR2_X1 U12905 ( .A(n13762), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n10355) );
  NOR2_X1 U12906 ( .A1(n10356), .A2(n10355), .ZN(n13761) );
  AOI211_X1 U12907 ( .C1(n10356), .C2(n10355), .A(n14669), .B(n13761), .ZN(
        n10360) );
  INV_X1 U12908 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10358) );
  NAND2_X1 U12909 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n11235)
         );
  NAND2_X1 U12910 ( .A1(n14676), .A2(n13762), .ZN(n10357) );
  OAI211_X1 U12911 ( .C1(n14679), .C2(n10358), .A(n11235), .B(n10357), .ZN(
        n10359) );
  AOI211_X1 U12912 ( .C1(n10361), .C2(n14636), .A(n10360), .B(n10359), .ZN(
        n10362) );
  INV_X1 U12913 ( .A(n10362), .ZN(P1_U3254) );
  AOI21_X1 U12914 ( .B1(n10373), .B2(P2_REG2_REG_10__SCAN_IN), .A(n10363), 
        .ZN(n10367) );
  INV_X1 U12915 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10364) );
  MUX2_X1 U12916 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n10364), .S(n10501), .Z(
        n10366) );
  INV_X1 U12917 ( .A(n10504), .ZN(n10365) );
  OAI21_X1 U12918 ( .B1(n10367), .B2(n10366), .A(n10365), .ZN(n10379) );
  NOR2_X1 U12919 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10368), .ZN(n10369) );
  AOI21_X1 U12920 ( .B1(n14840), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n10369), 
        .ZN(n10370) );
  OAI21_X1 U12921 ( .B1(n13184), .B2(n10371), .A(n10370), .ZN(n10378) );
  INV_X1 U12922 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10374) );
  MUX2_X1 U12923 ( .A(n10374), .B(P2_REG1_REG_11__SCAN_IN), .S(n10501), .Z(
        n10375) );
  AOI211_X1 U12924 ( .C1(n10376), .C2(n10375), .A(n14856), .B(n10497), .ZN(
        n10377) );
  AOI211_X1 U12925 ( .C1(n13224), .C2(n10379), .A(n10378), .B(n10377), .ZN(
        n10380) );
  INV_X1 U12926 ( .A(n10380), .ZN(P2_U3225) );
  OAI22_X1 U12927 ( .A1(n13426), .A2(n10382), .B1(n10381), .B2(n13377), .ZN(
        n10386) );
  OAI22_X1 U12928 ( .A1(n10384), .A2(n13415), .B1(n13325), .B2(n10383), .ZN(
        n10385) );
  AOI211_X1 U12929 ( .C1(P2_REG2_REG_1__SCAN_IN), .C2(n13426), .A(n10386), .B(
        n10385), .ZN(n10387) );
  OAI21_X1 U12930 ( .B1(n13421), .B2(n10388), .A(n10387), .ZN(P2_U3264) );
  NAND2_X1 U12931 ( .A1(n12975), .A2(n13089), .ZN(n10389) );
  NAND2_X1 U12932 ( .A1(n10390), .A2(n10389), .ZN(n10423) );
  XNOR2_X1 U12933 ( .A(n10423), .B(n10396), .ZN(n10415) );
  OAI22_X1 U12934 ( .A1(n10476), .A2(n13052), .B1(n10393), .B2(n13051), .ZN(
        n10400) );
  OR2_X1 U12935 ( .A1(n12975), .A2(n10393), .ZN(n10394) );
  INV_X1 U12936 ( .A(n10396), .ZN(n10422) );
  NAND2_X1 U12937 ( .A1(n10397), .A2(n10422), .ZN(n10398) );
  AOI21_X1 U12938 ( .B1(n10428), .B2(n10398), .A(n13294), .ZN(n10399) );
  AOI211_X1 U12939 ( .C1(n10415), .C2(n10401), .A(n10400), .B(n10399), .ZN(
        n10418) );
  AOI21_X1 U12940 ( .B1(n10424), .B2(n10402), .A(n10433), .ZN(n10416) );
  INV_X1 U12941 ( .A(n10424), .ZN(n10403) );
  NOR2_X1 U12942 ( .A1(n10403), .A2(n13415), .ZN(n10406) );
  OAI22_X1 U12943 ( .A1(n13394), .A2(n9809), .B1(n10404), .B2(n13377), .ZN(
        n10405) );
  AOI211_X1 U12944 ( .C1(n10416), .C2(n13385), .A(n10406), .B(n10405), .ZN(
        n10409) );
  INV_X1 U12945 ( .A(n10438), .ZN(n10407) );
  NAND2_X1 U12946 ( .A1(n10415), .A2(n10407), .ZN(n10408) );
  OAI211_X1 U12947 ( .C1(n10418), .C2(n13426), .A(n10409), .B(n10408), .ZN(
        P2_U3256) );
  NAND2_X1 U12948 ( .A1(n12558), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n10410) );
  OAI21_X1 U12949 ( .B1(n12185), .B2(n12558), .A(n10410), .ZN(P3_U3520) );
  INV_X1 U12950 ( .A(n10411), .ZN(n10412) );
  OAI222_X1 U12951 ( .A1(P3_U3151), .A2(n10414), .B1(n12933), .B2(n10413), 
        .C1(n11500), .C2(n10412), .ZN(P3_U3274) );
  INV_X1 U12952 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n14226) );
  INV_X1 U12953 ( .A(n10415), .ZN(n10419) );
  AOI22_X1 U12954 ( .A1(n10416), .A2(n13505), .B1(n13513), .B2(n10424), .ZN(
        n10417) );
  OAI211_X1 U12955 ( .C1(n10420), .C2(n10419), .A(n10418), .B(n10417), .ZN(
        n13518) );
  NAND2_X1 U12956 ( .A1(n13518), .A2(n6443), .ZN(n10421) );
  OAI21_X1 U12957 ( .B1(n6443), .B2(n14226), .A(n10421), .ZN(P2_U3457) );
  NAND2_X1 U12958 ( .A1(n10423), .A2(n10422), .ZN(n10426) );
  NAND2_X1 U12959 ( .A1(n10424), .A2(n13088), .ZN(n10425) );
  XOR2_X1 U12960 ( .A(n10483), .B(n10429), .Z(n14920) );
  XNOR2_X1 U12961 ( .A(n10472), .B(n10429), .ZN(n10431) );
  OAI22_X1 U12962 ( .A1(n12960), .A2(n13052), .B1(n12972), .B2(n13051), .ZN(
        n10430) );
  AOI21_X1 U12963 ( .B1(n10431), .B2(n13406), .A(n10430), .ZN(n10432) );
  OAI21_X1 U12964 ( .B1(n14920), .B2(n9458), .A(n10432), .ZN(n14924) );
  NAND2_X1 U12965 ( .A1(n14924), .A2(n13394), .ZN(n10437) );
  OAI22_X1 U12966 ( .A1(n13394), .A2(n10121), .B1(n12956), .B2(n13377), .ZN(
        n10435) );
  INV_X1 U12967 ( .A(n12966), .ZN(n14923) );
  NAND2_X1 U12968 ( .A1(n14923), .A2(n10433), .ZN(n10478) );
  OAI211_X1 U12969 ( .C1(n14923), .C2(n10433), .A(n13505), .B(n10478), .ZN(
        n14921) );
  NOR2_X1 U12970 ( .A1(n14921), .A2(n13325), .ZN(n10434) );
  AOI211_X1 U12971 ( .C1(n13381), .C2(n12966), .A(n10435), .B(n10434), .ZN(
        n10436) );
  OAI211_X1 U12972 ( .C1(n14920), .C2(n10438), .A(n10437), .B(n10436), .ZN(
        P2_U3255) );
  OAI21_X1 U12973 ( .B1(n10440), .B2(n12363), .A(n10439), .ZN(n10703) );
  OAI211_X1 U12974 ( .C1(n10443), .C2(n10442), .A(n10441), .B(n12766), .ZN(
        n10445) );
  AOI22_X1 U12975 ( .A1(n12769), .A2(n12554), .B1(n12556), .B2(n11219), .ZN(
        n10444) );
  NAND2_X1 U12976 ( .A1(n10445), .A2(n10444), .ZN(n10700) );
  AOI21_X1 U12977 ( .B1(n15150), .B2(n10703), .A(n10700), .ZN(n10468) );
  OAI22_X1 U12978 ( .A1(n10699), .A2(n12926), .B1(n15158), .B2(n8765), .ZN(
        n10446) );
  INV_X1 U12979 ( .A(n10446), .ZN(n10447) );
  OAI21_X1 U12980 ( .B1(n10468), .B2(n15157), .A(n10447), .ZN(P3_U3402) );
  XNOR2_X1 U12981 ( .A(n10595), .B(n10448), .ZN(n10487) );
  XNOR2_X1 U12982 ( .A(n10487), .B(n15123), .ZN(n10453) );
  AOI211_X1 U12983 ( .C1(n10453), .C2(n10452), .A(n12534), .B(n6598), .ZN(
        n10454) );
  INV_X1 U12984 ( .A(n10454), .ZN(n10458) );
  AND2_X1 U12985 ( .A1(P3_U3151), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n14942) );
  OAI22_X1 U12986 ( .A1(n10455), .A2(n12505), .B1(n10710), .B2(n12527), .ZN(
        n10456) );
  AOI211_X1 U12987 ( .C1(n12515), .C2(n10595), .A(n14942), .B(n10456), .ZN(
        n10457) );
  OAI211_X1 U12988 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12461), .A(n10458), .B(
        n10457), .ZN(P3_U3158) );
  INV_X1 U12989 ( .A(n10459), .ZN(n10461) );
  OAI22_X1 U12990 ( .A1(n12415), .A2(P3_U3151), .B1(SI_22_), .B2(n12933), .ZN(
        n10460) );
  AOI21_X1 U12991 ( .B1(n10461), .B2(n12927), .A(n10460), .ZN(P3_U3273) );
  OAI22_X1 U12992 ( .A1(n12876), .A2(n10462), .B1(n15166), .B2(n8754), .ZN(
        n10463) );
  INV_X1 U12993 ( .A(n10463), .ZN(n10464) );
  OAI21_X1 U12994 ( .B1(n10465), .B2(n15164), .A(n10464), .ZN(P3_U3462) );
  OAI22_X1 U12995 ( .A1(n12876), .A2(n10699), .B1(n15166), .B2(n10543), .ZN(
        n10466) );
  INV_X1 U12996 ( .A(n10466), .ZN(n10467) );
  OAI21_X1 U12997 ( .B1(n10468), .B2(n15164), .A(n10467), .ZN(P3_U3463) );
  INV_X1 U12998 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n14252) );
  INV_X1 U12999 ( .A(n12354), .ZN(n10469) );
  NAND2_X1 U13000 ( .A1(n10469), .A2(P3_U3897), .ZN(n10470) );
  OAI21_X1 U13001 ( .B1(P3_U3897), .B2(n14252), .A(n10470), .ZN(P3_U3521) );
  OR2_X1 U13002 ( .A1(n12966), .A2(n10476), .ZN(n10471) );
  NAND2_X1 U13003 ( .A1(n12966), .A2(n10476), .ZN(n10473) );
  NAND2_X1 U13004 ( .A1(n10474), .A2(n10473), .ZN(n10670) );
  XNOR2_X1 U13005 ( .A(n10670), .B(n10669), .ZN(n10477) );
  OAI22_X1 U13006 ( .A1(n10901), .A2(n13052), .B1(n10476), .B2(n13051), .ZN(
        n12116) );
  AOI21_X1 U13007 ( .B1(n10477), .B2(n13406), .A(n12116), .ZN(n10613) );
  AOI211_X1 U13008 ( .C1(n12126), .C2(n10478), .A(n13409), .B(n7138), .ZN(
        n10612) );
  INV_X1 U13009 ( .A(n12126), .ZN(n10481) );
  INV_X1 U13010 ( .A(n12118), .ZN(n10479) );
  AOI22_X1 U13011 ( .A1(n13426), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n10479), 
        .B2(n13412), .ZN(n10480) );
  OAI21_X1 U13012 ( .B1(n10481), .B2(n13415), .A(n10480), .ZN(n10485) );
  AND2_X1 U13013 ( .A1(n12966), .A2(n13087), .ZN(n10482) );
  XNOR2_X1 U13014 ( .A(n10668), .B(n10669), .ZN(n10615) );
  NOR2_X1 U13015 ( .A1(n10615), .A2(n13421), .ZN(n10484) );
  AOI211_X1 U13016 ( .C1(n10612), .C2(n13424), .A(n10485), .B(n10484), .ZN(
        n10486) );
  OAI21_X1 U13017 ( .B1(n13426), .B2(n10613), .A(n10486), .ZN(P2_U3254) );
  XNOR2_X1 U13018 ( .A(n10494), .B(n7090), .ZN(n10705) );
  XNOR2_X1 U13019 ( .A(n12555), .B(n10705), .ZN(n10490) );
  INV_X1 U13020 ( .A(n10487), .ZN(n10488) );
  OAI21_X1 U13021 ( .B1(n10490), .B2(n10489), .A(n10706), .ZN(n10491) );
  NAND2_X1 U13022 ( .A1(n10491), .A2(n12499), .ZN(n10496) );
  NAND2_X1 U13023 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_U3151), .ZN(n14969) );
  INV_X1 U13024 ( .A(n14969), .ZN(n10493) );
  OAI22_X1 U13025 ( .A1(n10834), .A2(n12527), .B1(n15123), .B2(n12505), .ZN(
        n10492) );
  AOI211_X1 U13026 ( .C1(n10494), .C2(n12515), .A(n10493), .B(n10492), .ZN(
        n10495) );
  OAI211_X1 U13027 ( .C1(n10698), .C2(n12461), .A(n10496), .B(n10495), .ZN(
        P3_U3170) );
  INV_X1 U13028 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10498) );
  MUX2_X1 U13029 ( .A(n10498), .B(P2_REG1_REG_12__SCAN_IN), .S(n11105), .Z(
        n10499) );
  OAI21_X1 U13030 ( .B1(n10500), .B2(n10499), .A(n11111), .ZN(n10509) );
  NOR2_X1 U13031 ( .A1(n10501), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10502) );
  MUX2_X1 U13032 ( .A(n10678), .B(P2_REG2_REG_12__SCAN_IN), .S(n11105), .Z(
        n10503) );
  OAI21_X1 U13033 ( .B1(n10504), .B2(n10502), .A(n10503), .ZN(n11106) );
  OR3_X1 U13034 ( .A1(n10504), .A2(n10503), .A3(n10502), .ZN(n10505) );
  AOI21_X1 U13035 ( .B1(n11106), .B2(n10505), .A(n14864), .ZN(n10508) );
  NAND2_X1 U13036 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n12091)
         );
  NAND2_X1 U13037 ( .A1(n14840), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n10506) );
  OAI211_X1 U13038 ( .C1(n13184), .C2(n11105), .A(n12091), .B(n10506), .ZN(
        n10507) );
  AOI211_X1 U13039 ( .C1(n10509), .C2(n13223), .A(n10508), .B(n10507), .ZN(
        n10510) );
  INV_X1 U13040 ( .A(n10510), .ZN(P2_U3226) );
  INV_X1 U13041 ( .A(n13211), .ZN(n13204) );
  OAI222_X1 U13042 ( .A1(P2_U3088), .A2(n13204), .B1(n13549), .B2(n11611), 
        .C1(n10511), .C2(n13551), .ZN(P2_U3309) );
  NAND2_X1 U13043 ( .A1(n10312), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10512) );
  XNOR2_X1 U13044 ( .A(n10512), .B(n9218), .ZN(n13790) );
  OAI222_X1 U13045 ( .A1(P1_U3086), .A2(n13790), .B1(n14375), .B2(n11611), 
        .C1(n10513), .C2(n14372), .ZN(P1_U3337) );
  INV_X2 U13046 ( .A(n10514), .ZN(n12646) );
  MUX2_X1 U13047 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12646), .Z(n10964) );
  XNOR2_X1 U13048 ( .A(n10964), .B(n10963), .ZN(n10965) );
  MUX2_X1 U13049 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12646), .Z(n10530) );
  XOR2_X1 U13050 ( .A(n14994), .B(n10530), .Z(n14988) );
  MUX2_X1 U13051 ( .A(n10633), .B(n10515), .S(n12646), .Z(n10528) );
  NOR2_X1 U13052 ( .A1(n10528), .A2(n10550), .ZN(n14973) );
  INV_X1 U13053 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10532) );
  MUX2_X1 U13054 ( .A(n10532), .B(n10543), .S(n12646), .Z(n10526) );
  AND2_X1 U13055 ( .A1(n10526), .A2(n10542), .ZN(n10527) );
  NOR2_X1 U13056 ( .A1(n12646), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n10516) );
  AOI21_X1 U13057 ( .B1(n8754), .B2(n10517), .A(n10516), .ZN(n10522) );
  NOR2_X1 U13058 ( .A1(n10522), .A2(n14939), .ZN(n10524) );
  INV_X1 U13059 ( .A(n10518), .ZN(n10520) );
  AOI21_X1 U13060 ( .B1(n10521), .B2(n10520), .A(n10519), .ZN(n14938) );
  AOI21_X1 U13061 ( .B1(n10522), .B2(n14939), .A(n10524), .ZN(n10523) );
  INV_X1 U13062 ( .A(n10523), .ZN(n14937) );
  NOR2_X1 U13063 ( .A1(n14938), .A2(n14937), .ZN(n14936) );
  NOR2_X1 U13064 ( .A1(n10524), .A2(n14936), .ZN(n14962) );
  INV_X1 U13065 ( .A(n10527), .ZN(n10525) );
  OAI21_X1 U13066 ( .B1(n10542), .B2(n10526), .A(n10525), .ZN(n14963) );
  NOR2_X1 U13067 ( .A1(n14962), .A2(n14963), .ZN(n14961) );
  AND2_X1 U13068 ( .A1(n10528), .A2(n10550), .ZN(n14974) );
  INV_X1 U13069 ( .A(n14974), .ZN(n10529) );
  XNOR2_X1 U13070 ( .A(n10965), .B(n10962), .ZN(n10560) );
  NAND2_X1 U13071 ( .A1(n14967), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n10535) );
  NAND2_X1 U13072 ( .A1(n10542), .A2(n10532), .ZN(n10533) );
  NAND2_X1 U13073 ( .A1(n10535), .A2(n10533), .ZN(n14952) );
  NAND2_X1 U13074 ( .A1(n14949), .A2(n10534), .ZN(n14950) );
  NOR2_X1 U13075 ( .A1(n10550), .A2(n10536), .ZN(n10537) );
  NAND2_X1 U13076 ( .A1(n14994), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n10539) );
  OR2_X1 U13077 ( .A1(n14994), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n10538) );
  NAND2_X1 U13078 ( .A1(n10539), .A2(n10538), .ZN(n14992) );
  XNOR2_X1 U13079 ( .A(n8806), .B(n10952), .ZN(n10540) );
  NAND2_X1 U13080 ( .A1(n10540), .A2(n14960), .ZN(n10559) );
  NAND2_X1 U13081 ( .A1(n14994), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n10553) );
  MUX2_X1 U13082 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n10541), .S(n14994), .Z(
        n14996) );
  NAND2_X1 U13083 ( .A1(n14967), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n10549) );
  MUX2_X1 U13084 ( .A(n10543), .B(P3_REG1_REG_4__SCAN_IN), .S(n10542), .Z(
        n14956) );
  NAND2_X1 U13085 ( .A1(n14939), .A2(n10547), .ZN(n10548) );
  XNOR2_X1 U13086 ( .A(n10547), .B(n10546), .ZN(n14944) );
  NAND2_X1 U13087 ( .A1(P3_REG1_REG_3__SCAN_IN), .A2(n14944), .ZN(n14943) );
  NAND2_X1 U13088 ( .A1(n10548), .A2(n14943), .ZN(n14957) );
  NAND2_X1 U13089 ( .A1(n14956), .A2(n14957), .ZN(n14955) );
  NAND2_X1 U13090 ( .A1(n10549), .A2(n14955), .ZN(n10551) );
  NAND2_X1 U13091 ( .A1(n14977), .A2(n10551), .ZN(n10552) );
  XNOR2_X1 U13092 ( .A(n10551), .B(n10550), .ZN(n14982) );
  NAND2_X1 U13093 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n14982), .ZN(n14981) );
  NAND2_X1 U13094 ( .A1(n10552), .A2(n14981), .ZN(n14997) );
  NAND2_X1 U13095 ( .A1(n14996), .A2(n14997), .ZN(n14995) );
  NAND2_X1 U13096 ( .A1(n10553), .A2(n14995), .ZN(n10945) );
  XNOR2_X1 U13097 ( .A(n10945), .B(n10951), .ZN(n10554) );
  NAND2_X1 U13098 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n10554), .ZN(n10946) );
  OAI21_X1 U13099 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n10554), .A(n10946), .ZN(
        n10557) );
  AND2_X1 U13100 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n10923) );
  AOI21_X1 U13101 ( .B1(n15082), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n10923), .ZN(
        n10555) );
  OAI21_X1 U13102 ( .B1(n15101), .B2(n10963), .A(n10555), .ZN(n10556) );
  AOI21_X1 U13103 ( .B1(n15107), .B2(n10557), .A(n10556), .ZN(n10558) );
  OAI211_X1 U13104 ( .C1(n10560), .C2(n15109), .A(n10559), .B(n10558), .ZN(
        P3_U3189) );
  OR2_X1 U13105 ( .A1(n10561), .A2(n11610), .ZN(n10563) );
  AOI22_X1 U13106 ( .A1(n11627), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n11626), 
        .B2(n13748), .ZN(n10562) );
  NAND2_X1 U13107 ( .A1(n10563), .A2(n10562), .ZN(n14712) );
  INV_X1 U13108 ( .A(n14712), .ZN(n14800) );
  INV_X1 U13109 ( .A(n13685), .ZN(n13652) );
  INV_X1 U13110 ( .A(n10565), .ZN(n10566) );
  NAND2_X1 U13111 ( .A1(n10564), .A2(n10566), .ZN(n10567) );
  NAND2_X1 U13112 ( .A1(n10568), .A2(n10567), .ZN(n10572) );
  AND2_X1 U13113 ( .A1(n14682), .A2(n11808), .ZN(n10569) );
  AOI21_X1 U13114 ( .B1(n14712), .B2(n11775), .A(n10569), .ZN(n10815) );
  AOI22_X1 U13115 ( .A1(n14712), .A2(n11807), .B1(n11775), .B2(n14682), .ZN(
        n10570) );
  XNOR2_X1 U13116 ( .A(n10570), .B(n10326), .ZN(n10814) );
  XOR2_X1 U13117 ( .A(n10815), .B(n10814), .Z(n10571) );
  OAI211_X1 U13118 ( .C1(n10572), .C2(n10571), .A(n10819), .B(n13645), .ZN(
        n10581) );
  NAND2_X1 U13119 ( .A1(n11846), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10577) );
  OR2_X1 U13120 ( .A1(n11818), .A2(n10573), .ZN(n10576) );
  OR2_X1 U13121 ( .A1(n11839), .A2(n9748), .ZN(n10575) );
  XNOR2_X1 U13122 ( .A(n10732), .B(n14306), .ZN(n14690) );
  OR2_X1 U13123 ( .A1(n9605), .A2(n14690), .ZN(n10574) );
  NAND4_X1 U13124 ( .A1(n10577), .A2(n10576), .A3(n10575), .A4(n10574), .ZN(
        n14703) );
  INV_X1 U13125 ( .A(n13664), .ZN(n13679) );
  NAND2_X1 U13126 ( .A1(n13681), .A2(n14704), .ZN(n10578) );
  NAND2_X1 U13127 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n13745) );
  OAI211_X1 U13128 ( .C1(n13679), .C2(n14709), .A(n10578), .B(n13745), .ZN(
        n10579) );
  AOI21_X1 U13129 ( .B1(n6433), .B2(n14703), .A(n10579), .ZN(n10580) );
  OAI211_X1 U13130 ( .C1(n14800), .C2(n13652), .A(n10581), .B(n10580), .ZN(
        P1_U3213) );
  INV_X1 U13131 ( .A(n10582), .ZN(n10601) );
  INV_X1 U13132 ( .A(n10583), .ZN(n10586) );
  MUX2_X1 U13133 ( .A(n10586), .B(n10585), .S(n10584), .Z(n10588) );
  NAND2_X1 U13134 ( .A1(n10588), .A2(n10587), .ZN(n10591) );
  AND2_X1 U13135 ( .A1(n10603), .A2(n12195), .ZN(n15131) );
  OR2_X1 U13136 ( .A1(n15125), .A2(n15131), .ZN(n10590) );
  INV_X1 U13137 ( .A(n10591), .ZN(n10593) );
  NOR2_X1 U13138 ( .A1(n10603), .A2(n15144), .ZN(n10592) );
  AOI22_X1 U13139 ( .A1(n14471), .A2(n10595), .B1(n15134), .B2(n10594), .ZN(
        n10596) );
  OAI21_X1 U13140 ( .B1(n10597), .B2(n12818), .A(n10596), .ZN(n10598) );
  AOI21_X1 U13141 ( .B1(n10599), .B2(n12821), .A(n10598), .ZN(n10600) );
  OAI21_X1 U13142 ( .B1(n10601), .B2(n15136), .A(n10600), .ZN(P3_U3230) );
  AND2_X1 U13143 ( .A1(n10602), .A2(n15152), .ZN(n15138) );
  INV_X1 U13144 ( .A(n10603), .ZN(n15130) );
  XNOR2_X1 U13145 ( .A(n10043), .B(n10604), .ZN(n10605) );
  NAND2_X1 U13146 ( .A1(n10605), .A2(n12766), .ZN(n10607) );
  AOI22_X1 U13147 ( .A1(n12769), .A2(n10051), .B1(n12559), .B2(n11219), .ZN(
        n10606) );
  NAND2_X1 U13148 ( .A1(n10607), .A2(n10606), .ZN(n15137) );
  AOI21_X1 U13149 ( .B1(n15138), .B2(n15130), .A(n15137), .ZN(n10611) );
  XNOR2_X1 U13150 ( .A(n12199), .B(n12193), .ZN(n15139) );
  OAI22_X1 U13151 ( .A1(n12818), .A2(n9829), .B1(n10608), .B2(n12816), .ZN(
        n10609) );
  AOI21_X1 U13152 ( .B1(n15139), .B2(n12821), .A(n10609), .ZN(n10610) );
  OAI21_X1 U13153 ( .B1(n10611), .B2(n15136), .A(n10610), .ZN(P3_U3232) );
  INV_X1 U13154 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10617) );
  AOI21_X1 U13155 ( .B1(n13513), .B2(n12126), .A(n10612), .ZN(n10614) );
  OAI211_X1 U13156 ( .C1(n10615), .C2(n13516), .A(n10614), .B(n10613), .ZN(
        n13517) );
  NAND2_X1 U13157 ( .A1(n13517), .A2(n6443), .ZN(n10616) );
  OAI21_X1 U13158 ( .B1(n6443), .B2(n10617), .A(n10616), .ZN(P2_U3463) );
  OAI21_X1 U13159 ( .B1(n10619), .B2(n12358), .A(n10618), .ZN(n10635) );
  INV_X1 U13160 ( .A(n10635), .ZN(n10625) );
  NAND2_X1 U13161 ( .A1(n10620), .A2(n12358), .ZN(n10621) );
  NAND2_X1 U13162 ( .A1(n10622), .A2(n10621), .ZN(n10624) );
  OAI22_X1 U13163 ( .A1(n10710), .A2(n12799), .B1(n10921), .B2(n15122), .ZN(
        n10623) );
  AOI21_X1 U13164 ( .B1(n10624), .B2(n12766), .A(n10623), .ZN(n10632) );
  OAI21_X1 U13165 ( .B1(n10625), .B2(n14483), .A(n10632), .ZN(n10811) );
  INV_X1 U13166 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n10626) );
  OAI22_X1 U13167 ( .A1(n10809), .A2(n12926), .B1(n15158), .B2(n10626), .ZN(
        n10627) );
  AOI21_X1 U13168 ( .B1(n10811), .B2(n15158), .A(n10627), .ZN(n10628) );
  INV_X1 U13169 ( .A(n10628), .ZN(P3_U3405) );
  NAND2_X1 U13170 ( .A1(n10629), .A2(n12927), .ZN(n10630) );
  OAI211_X1 U13171 ( .C1(n10631), .C2(n12933), .A(n10630), .B(n12417), .ZN(
        P3_U3272) );
  MUX2_X1 U13172 ( .A(n10633), .B(n10632), .S(n12818), .Z(n10637) );
  OAI22_X1 U13173 ( .A1(n12815), .A2(n10809), .B1(n10715), .B2(n12816), .ZN(
        n10634) );
  AOI21_X1 U13174 ( .B1(n10635), .B2(n12821), .A(n10634), .ZN(n10636) );
  NAND2_X1 U13175 ( .A1(n10637), .A2(n10636), .ZN(P3_U3228) );
  INV_X1 U13176 ( .A(n10638), .ZN(n10642) );
  INV_X1 U13177 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n14325) );
  OAI22_X1 U13178 ( .A1(n10644), .A2(n11853), .B1(n14325), .B2(n14751), .ZN(
        n10641) );
  OR2_X1 U13179 ( .A1(n10640), .A2(n10639), .ZN(n13869) );
  OAI21_X1 U13180 ( .B1(n10642), .B2(n10641), .A(n14691), .ZN(n10648) );
  NAND2_X1 U13181 ( .A1(n9514), .A2(n12058), .ZN(n11870) );
  AND2_X1 U13182 ( .A1(n10791), .A2(n11870), .ZN(n10643) );
  OAI22_X1 U13183 ( .A1(n14695), .A2(n10644), .B1(n14691), .B2(n9251), .ZN(
        n10645) );
  AOI21_X1 U13184 ( .B1(n10646), .B2(n14697), .A(n10645), .ZN(n10647) );
  NAND2_X1 U13185 ( .A1(n10648), .A2(n10647), .ZN(P1_U3293) );
  NAND2_X1 U13186 ( .A1(n13581), .A2(n10695), .ZN(n14741) );
  INV_X1 U13187 ( .A(n10687), .ZN(n13698) );
  NAND2_X1 U13188 ( .A1(n13698), .A2(n14773), .ZN(n11892) );
  INV_X1 U13189 ( .A(n12036), .ZN(n10650) );
  NAND3_X1 U13190 ( .A1(n14746), .A2(n11891), .A3(n12036), .ZN(n10651) );
  NAND2_X1 U13191 ( .A1(n14726), .A2(n10651), .ZN(n10654) );
  INV_X1 U13192 ( .A(n14705), .ZN(n14722) );
  NAND2_X1 U13193 ( .A1(n13696), .A2(n14702), .ZN(n10652) );
  OAI21_X1 U13194 ( .B1(n10687), .B2(n14722), .A(n10652), .ZN(n10653) );
  AOI21_X1 U13195 ( .B1(n10654), .B2(n14685), .A(n10653), .ZN(n14780) );
  MUX2_X1 U13196 ( .A(n14326), .B(n14780), .S(n14691), .Z(n10667) );
  NAND2_X1 U13197 ( .A1(n9671), .A2(n11872), .ZN(n10657) );
  NAND2_X1 U13198 ( .A1(n13581), .A2(n6952), .ZN(n10658) );
  NAND2_X1 U13199 ( .A1(n14740), .A2(n14742), .ZN(n10741) );
  NAND2_X1 U13200 ( .A1(n10687), .A2(n14773), .ZN(n10739) );
  NAND2_X1 U13201 ( .A1(n10741), .A2(n10739), .ZN(n10659) );
  XNOR2_X1 U13202 ( .A(n10659), .B(n12036), .ZN(n14783) );
  INV_X1 U13203 ( .A(n14755), .ZN(n10661) );
  INV_X1 U13204 ( .A(n14736), .ZN(n10660) );
  OAI211_X1 U13205 ( .C1(n14781), .C2(n10661), .A(n10660), .B(n14756), .ZN(
        n14779) );
  INV_X1 U13206 ( .A(n14751), .ZN(n14710) );
  AOI22_X1 U13207 ( .A1(n14754), .A2(n11895), .B1(n14710), .B2(n10663), .ZN(
        n10664) );
  OAI21_X1 U13208 ( .B1(n14779), .B2(n14695), .A(n10664), .ZN(n10665) );
  AOI21_X1 U13209 ( .B1(n14783), .B2(n14697), .A(n10665), .ZN(n10666) );
  NAND2_X1 U13210 ( .A1(n10667), .A2(n10666), .ZN(P1_U3289) );
  XOR2_X1 U13211 ( .A(n10673), .B(n10905), .Z(n10870) );
  INV_X1 U13212 ( .A(n10870), .ZN(n10684) );
  NAND2_X1 U13213 ( .A1(n10670), .A2(n10669), .ZN(n10672) );
  NAND2_X1 U13214 ( .A1(n12126), .A2(n12960), .ZN(n10671) );
  AOI21_X1 U13215 ( .B1(n10674), .B2(n10673), .A(n13294), .ZN(n10675) );
  OAI22_X1 U13216 ( .A1(n14499), .A2(n13052), .B1(n12960), .B2(n13051), .ZN(
        n12090) );
  AOI21_X1 U13217 ( .B1(n10675), .B2(n10903), .A(n12090), .ZN(n10868) );
  INV_X1 U13218 ( .A(n10868), .ZN(n10682) );
  AOI21_X1 U13219 ( .B1(n12100), .B2(n10676), .A(n13409), .ZN(n10677) );
  NAND2_X1 U13220 ( .A1(n10677), .A2(n10909), .ZN(n10867) );
  OAI22_X1 U13221 ( .A1(n13394), .A2(n10678), .B1(n12093), .B2(n13377), .ZN(
        n10679) );
  AOI21_X1 U13222 ( .B1(n12100), .B2(n13381), .A(n10679), .ZN(n10680) );
  OAI21_X1 U13223 ( .B1(n10867), .B2(n13325), .A(n10680), .ZN(n10681) );
  AOI21_X1 U13224 ( .B1(n10682), .B2(n13394), .A(n10681), .ZN(n10683) );
  OAI21_X1 U13225 ( .B1(n10684), .B2(n13421), .A(n10683), .ZN(P2_U3253) );
  XNOR2_X1 U13226 ( .A(n10685), .B(n12034), .ZN(n14769) );
  NOR2_X1 U13227 ( .A1(n6442), .A2(n11870), .ZN(n14760) );
  INV_X1 U13228 ( .A(n14760), .ZN(n10806) );
  OAI21_X1 U13229 ( .B1(n12034), .B2(n10686), .A(n14743), .ZN(n10689) );
  OAI22_X1 U13230 ( .A1(n9671), .A2(n14722), .B1(n10687), .B2(n14720), .ZN(
        n10688) );
  AOI21_X1 U13231 ( .B1(n10689), .B2(n14685), .A(n10688), .ZN(n10690) );
  OAI21_X1 U13232 ( .B1(n14769), .B2(n10791), .A(n10690), .ZN(n14771) );
  NAND2_X1 U13233 ( .A1(n14771), .A2(n14691), .ZN(n10697) );
  OAI22_X1 U13234 ( .A1(n14691), .A2(n9298), .B1(n10691), .B2(n14751), .ZN(
        n10694) );
  NOR2_X1 U13235 ( .A1(n14767), .A2(n14695), .ZN(n10693) );
  AOI211_X1 U13236 ( .C1(n14754), .C2(n10695), .A(n10694), .B(n10693), .ZN(
        n10696) );
  OAI211_X1 U13237 ( .C1(n14769), .C2(n10806), .A(n10697), .B(n10696), .ZN(
        P1_U3291) );
  OAI22_X1 U13238 ( .A1(n12815), .A2(n10699), .B1(n10698), .B2(n12816), .ZN(
        n10702) );
  MUX2_X1 U13239 ( .A(n10700), .B(P3_REG2_REG_4__SCAN_IN), .S(n15136), .Z(
        n10701) );
  AOI211_X1 U13240 ( .C1(n12821), .C2(n10703), .A(n10702), .B(n10701), .ZN(
        n10704) );
  INV_X1 U13241 ( .A(n10704), .ZN(P3_U3229) );
  INV_X1 U13242 ( .A(n10705), .ZN(n10707) );
  XNOR2_X1 U13243 ( .A(n10712), .B(n12180), .ZN(n10780) );
  XNOR2_X1 U13244 ( .A(n12554), .B(n10780), .ZN(n10781) );
  XNOR2_X1 U13245 ( .A(n10782), .B(n10781), .ZN(n10708) );
  NAND2_X1 U13246 ( .A1(n10708), .A2(n12499), .ZN(n10714) );
  NOR2_X1 U13247 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10709), .ZN(n14980) );
  OAI22_X1 U13248 ( .A1(n10710), .A2(n12505), .B1(n10921), .B2(n12527), .ZN(
        n10711) );
  AOI211_X1 U13249 ( .C1(n12515), .C2(n10712), .A(n14980), .B(n10711), .ZN(
        n10713) );
  OAI211_X1 U13250 ( .C1(n10715), .C2(n12461), .A(n10714), .B(n10713), .ZN(
        P3_U3167) );
  NAND2_X1 U13251 ( .A1(n10716), .A2(n14691), .ZN(n10723) );
  OAI22_X1 U13252 ( .A1(n14691), .A2(n10718), .B1(n10717), .B2(n14751), .ZN(
        n10721) );
  NOR2_X1 U13253 ( .A1(n10719), .A2(n14695), .ZN(n10720) );
  AOI211_X1 U13254 ( .C1(n14754), .C2(n11876), .A(n10721), .B(n10720), .ZN(
        n10722) );
  OAI211_X1 U13255 ( .C1(n10724), .C2(n10806), .A(n10723), .B(n10722), .ZN(
        P1_U3292) );
  OR2_X1 U13256 ( .A1(n10725), .A2(n11610), .ZN(n10728) );
  AOI22_X1 U13257 ( .A1(n11627), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n11626), 
        .B2(n10726), .ZN(n10727) );
  NAND2_X1 U13258 ( .A1(n11814), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10738) );
  OR2_X1 U13259 ( .A1(n11818), .A2(n10729), .ZN(n10737) );
  INV_X1 U13260 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10730) );
  OAI21_X1 U13261 ( .B1(n10732), .B2(n14306), .A(n10730), .ZN(n10733) );
  NAND2_X1 U13262 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n10731) );
  NAND2_X1 U13263 ( .A1(n10733), .A2(n10758), .ZN(n10984) );
  OR2_X1 U13264 ( .A1(n9605), .A2(n10984), .ZN(n10736) );
  INV_X1 U13265 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10734) );
  OR2_X1 U13266 ( .A1(n11816), .A2(n10734), .ZN(n10735) );
  NAND4_X1 U13267 ( .A1(n10738), .A2(n10737), .A3(n10736), .A4(n10735), .ZN(
        n14683) );
  XNOR2_X1 U13268 ( .A(n11923), .B(n11139), .ZN(n12042) );
  INV_X1 U13269 ( .A(n12042), .ZN(n10757) );
  NAND2_X1 U13270 ( .A1(n14723), .A2(n14781), .ZN(n10742) );
  AND2_X1 U13271 ( .A1(n10739), .A2(n10742), .ZN(n10740) );
  NAND2_X1 U13272 ( .A1(n10741), .A2(n10740), .ZN(n10745) );
  INV_X1 U13273 ( .A(n10742), .ZN(n10743) );
  NAND2_X1 U13274 ( .A1(n10793), .A2(n14734), .ZN(n10794) );
  NAND2_X1 U13275 ( .A1(n13696), .A2(n14785), .ZN(n10746) );
  NAND2_X1 U13276 ( .A1(n10794), .A2(n10746), .ZN(n14724) );
  NOR2_X1 U13277 ( .A1(n13696), .A2(n14734), .ZN(n10747) );
  XNOR2_X1 U13278 ( .A(n14793), .B(n14704), .ZN(n12038) );
  OAI22_X1 U13279 ( .A1(n10790), .A2(n12038), .B1(n14793), .B2(n14704), .ZN(
        n14699) );
  XNOR2_X1 U13280 ( .A(n14712), .B(n14682), .ZN(n12039) );
  INV_X1 U13281 ( .A(n14682), .ZN(n10792) );
  AOI22_X1 U13282 ( .A1(n14699), .A2(n14700), .B1(n10792), .B2(n14800), .ZN(
        n14687) );
  OR2_X1 U13283 ( .A1(n10748), .A2(n11610), .ZN(n10751) );
  AOI22_X1 U13284 ( .A1(n11627), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n11626), 
        .B2(n10749), .ZN(n10750) );
  NAND2_X1 U13285 ( .A1(n10751), .A2(n10750), .ZN(n14693) );
  NAND2_X1 U13286 ( .A1(n10753), .A2(n10752), .ZN(n10754) );
  AOI21_X1 U13287 ( .B1(n10757), .B2(n10756), .A(n6595), .ZN(n14813) );
  NAND2_X1 U13288 ( .A1(n11845), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10765) );
  OR2_X1 U13289 ( .A1(n11839), .A2(n10353), .ZN(n10764) );
  INV_X1 U13290 ( .A(n10852), .ZN(n10760) );
  NAND2_X1 U13291 ( .A1(n10758), .A2(n11136), .ZN(n10759) );
  NAND2_X1 U13292 ( .A1(n10760), .A2(n10759), .ZN(n10861) );
  OR2_X1 U13293 ( .A1(n9605), .A2(n10861), .ZN(n10763) );
  INV_X1 U13294 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10761) );
  OR2_X1 U13295 ( .A1(n11816), .A2(n10761), .ZN(n10762) );
  NAND4_X1 U13296 ( .A1(n10765), .A2(n10764), .A3(n10763), .A4(n10762), .ZN(
        n13694) );
  INV_X1 U13297 ( .A(n14724), .ZN(n10766) );
  INV_X1 U13298 ( .A(n14704), .ZN(n14721) );
  NAND2_X1 U13299 ( .A1(n14793), .A2(n14721), .ZN(n10767) );
  NAND2_X1 U13300 ( .A1(n10797), .A2(n10767), .ZN(n14701) );
  OR2_X1 U13301 ( .A1(n14712), .A2(n10792), .ZN(n10768) );
  NAND2_X1 U13302 ( .A1(n14701), .A2(n10768), .ZN(n10770) );
  NAND2_X1 U13303 ( .A1(n14712), .A2(n10792), .ZN(n10769) );
  INV_X1 U13304 ( .A(n14686), .ZN(n10771) );
  OR2_X1 U13305 ( .A1(n14693), .A2(n10752), .ZN(n10772) );
  INV_X1 U13306 ( .A(n10848), .ZN(n10773) );
  AOI21_X1 U13307 ( .B1(n12042), .B2(n10774), .A(n10773), .ZN(n10775) );
  OAI222_X1 U13308 ( .A1(n14720), .A2(n10888), .B1(n14722), .B2(n10752), .C1(
        n14744), .C2(n10775), .ZN(n14816) );
  NAND2_X1 U13309 ( .A1(n14816), .A2(n14691), .ZN(n10779) );
  OAI22_X1 U13310 ( .A1(n14691), .A2(n9954), .B1(n10984), .B2(n14751), .ZN(
        n10777) );
  NAND2_X1 U13311 ( .A1(n14688), .A2(n14815), .ZN(n10892) );
  OAI211_X1 U13312 ( .C1(n14688), .C2(n14815), .A(n14756), .B(n10892), .ZN(
        n14814) );
  NOR2_X1 U13313 ( .A1(n14814), .A2(n14695), .ZN(n10776) );
  AOI211_X1 U13314 ( .C1(n14754), .C2(n11923), .A(n10777), .B(n10776), .ZN(
        n10778) );
  OAI211_X1 U13315 ( .C1(n14813), .C2(n14059), .A(n10779), .B(n10778), .ZN(
        P1_U3284) );
  XNOR2_X1 U13316 ( .A(n10787), .B(n12180), .ZN(n10917) );
  XNOR2_X1 U13317 ( .A(n12553), .B(n10917), .ZN(n10783) );
  NAND2_X1 U13318 ( .A1(n10784), .A2(n10783), .ZN(n10919) );
  OAI211_X1 U13319 ( .C1(n10784), .C2(n10783), .A(n10919), .B(n12499), .ZN(
        n10789) );
  NAND2_X1 U13320 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n15005) );
  INV_X1 U13321 ( .A(n15005), .ZN(n10786) );
  OAI22_X1 U13322 ( .A1(n10834), .A2(n12505), .B1(n11081), .B2(n12527), .ZN(
        n10785) );
  AOI211_X1 U13323 ( .C1(n12515), .C2(n10787), .A(n10786), .B(n10785), .ZN(
        n10788) );
  OAI211_X1 U13324 ( .C1(n10991), .C2(n12461), .A(n10789), .B(n10788), .ZN(
        P3_U3179) );
  XNOR2_X1 U13325 ( .A(n10790), .B(n12038), .ZN(n10800) );
  INV_X1 U13326 ( .A(n10800), .ZN(n14796) );
  INV_X1 U13327 ( .A(n10791), .ZN(n14749) );
  OAI22_X1 U13328 ( .A1(n10793), .A2(n14722), .B1(n10792), .B2(n14720), .ZN(
        n10799) );
  INV_X1 U13329 ( .A(n12038), .ZN(n10795) );
  NAND3_X1 U13330 ( .A1(n14728), .A2(n10795), .A3(n10794), .ZN(n10796) );
  AOI21_X1 U13331 ( .B1(n10797), .B2(n10796), .A(n14744), .ZN(n10798) );
  AOI211_X1 U13332 ( .C1(n10800), .C2(n14749), .A(n10799), .B(n10798), .ZN(
        n14795) );
  MUX2_X1 U13333 ( .A(n9488), .B(n14795), .S(n14691), .Z(n10805) );
  AOI21_X1 U13334 ( .B1(n14735), .B2(n14793), .A(n14090), .ZN(n10801) );
  AND2_X1 U13335 ( .A1(n10801), .A2(n14713), .ZN(n14791) );
  OAI22_X1 U13336 ( .A1(n14047), .A2(n6957), .B1(n14751), .B2(n10802), .ZN(
        n10803) );
  AOI21_X1 U13337 ( .B1(n14791), .B2(n14759), .A(n10803), .ZN(n10804) );
  OAI211_X1 U13338 ( .C1(n14796), .C2(n10806), .A(n10805), .B(n10804), .ZN(
        P1_U3287) );
  OAI22_X1 U13339 ( .A1(n12876), .A2(n11836), .B1(n15166), .B2(n9828), .ZN(
        n10807) );
  AOI21_X1 U13340 ( .B1(n11832), .B2(n15166), .A(n10807), .ZN(n10808) );
  INV_X1 U13341 ( .A(n10808), .ZN(P3_U3459) );
  OAI22_X1 U13342 ( .A1(n12876), .A2(n10809), .B1(n15166), .B2(n10515), .ZN(
        n10810) );
  AOI21_X1 U13343 ( .B1(n10811), .B2(n15166), .A(n10810), .ZN(n10812) );
  INV_X1 U13344 ( .A(n10812), .ZN(P3_U3464) );
  AOI22_X1 U13345 ( .A1(n14693), .A2(n11807), .B1(n11775), .B2(n14703), .ZN(
        n10813) );
  XNOR2_X1 U13346 ( .A(n10813), .B(n10326), .ZN(n10976) );
  AOI22_X1 U13347 ( .A1(n14693), .A2(n11775), .B1(n11808), .B2(n14703), .ZN(
        n10977) );
  XNOR2_X1 U13348 ( .A(n10976), .B(n10977), .ZN(n10821) );
  INV_X1 U13349 ( .A(n10814), .ZN(n10817) );
  AOI21_X1 U13350 ( .B1(n10821), .B2(n10820), .A(n10975), .ZN(n10828) );
  AND2_X1 U13351 ( .A1(n14693), .A2(n14792), .ZN(n14806) );
  NOR2_X1 U13352 ( .A1(n13679), .A2(n14690), .ZN(n10822) );
  AOI211_X1 U13353 ( .C1(n13681), .C2(n14682), .A(n10823), .B(n10822), .ZN(
        n10824) );
  OAI21_X1 U13354 ( .B1(n11139), .B2(n13683), .A(n10824), .ZN(n10825) );
  AOI21_X1 U13355 ( .B1(n14806), .B2(n10826), .A(n10825), .ZN(n10827) );
  OAI21_X1 U13356 ( .B1(n10828), .B2(n13688), .A(n10827), .ZN(P1_U3221) );
  OAI21_X1 U13357 ( .B1(n10830), .B2(n12362), .A(n10829), .ZN(n10996) );
  OAI211_X1 U13358 ( .C1(n10833), .C2(n10832), .A(n10831), .B(n12766), .ZN(
        n10837) );
  OAI22_X1 U13359 ( .A1(n10834), .A2(n12799), .B1(n11081), .B2(n15122), .ZN(
        n10835) );
  INV_X1 U13360 ( .A(n10835), .ZN(n10836) );
  NAND2_X1 U13361 ( .A1(n10837), .A2(n10836), .ZN(n10993) );
  AOI21_X1 U13362 ( .B1(n15150), .B2(n10996), .A(n10993), .ZN(n10842) );
  OAI22_X1 U13363 ( .A1(n10992), .A2(n12926), .B1(n15158), .B2(n8796), .ZN(
        n10838) );
  INV_X1 U13364 ( .A(n10838), .ZN(n10839) );
  OAI21_X1 U13365 ( .B1(n10842), .B2(n15157), .A(n10839), .ZN(P3_U3408) );
  OAI22_X1 U13366 ( .A1(n12876), .A2(n10992), .B1(n15166), .B2(n10541), .ZN(
        n10840) );
  INV_X1 U13367 ( .A(n10840), .ZN(n10841) );
  OAI21_X1 U13368 ( .B1(n10842), .B2(n15164), .A(n10841), .ZN(P3_U3465) );
  INV_X1 U13369 ( .A(n10891), .ZN(n10846) );
  OR2_X1 U13370 ( .A1(n10843), .A2(n11610), .ZN(n10845) );
  AOI22_X1 U13371 ( .A1(n11627), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n11626), 
        .B2(n14597), .ZN(n10844) );
  XNOR2_X1 U13372 ( .A(n11927), .B(n10888), .ZN(n12043) );
  XNOR2_X1 U13373 ( .A(n10846), .B(n12043), .ZN(n14825) );
  NAND2_X1 U13374 ( .A1(n11923), .A2(n11139), .ZN(n10847) );
  AOI21_X1 U13375 ( .B1(n10849), .B2(n12043), .A(n14744), .ZN(n10850) );
  AOI22_X1 U13376 ( .A1(n10850), .A2(n10887), .B1(n14705), .B2(n14683), .ZN(
        n14820) );
  NOR2_X1 U13377 ( .A1(n14820), .A2(n6442), .ZN(n10865) );
  INV_X1 U13378 ( .A(n11927), .ZN(n14822) );
  XNOR2_X1 U13379 ( .A(n10892), .B(n14822), .ZN(n10860) );
  NAND2_X1 U13380 ( .A1(n11814), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10858) );
  OR2_X1 U13381 ( .A1(n11818), .A2(n10851), .ZN(n10857) );
  OR2_X1 U13382 ( .A1(n10852), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10853) );
  NAND2_X1 U13383 ( .A1(n10877), .A2(n10853), .ZN(n11236) );
  OR2_X1 U13384 ( .A1(n9605), .A2(n11236), .ZN(n10856) );
  INV_X1 U13385 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10854) );
  OR2_X1 U13386 ( .A1(n11816), .A2(n10854), .ZN(n10855) );
  NAND4_X1 U13387 ( .A1(n10858), .A2(n10857), .A3(n10856), .A4(n10855), .ZN(
        n13693) );
  AND2_X1 U13388 ( .A1(n13693), .A2(n14702), .ZN(n10859) );
  AOI21_X1 U13389 ( .B1(n10860), .B2(n14756), .A(n10859), .ZN(n14819) );
  INV_X1 U13390 ( .A(n10861), .ZN(n11137) );
  AOI22_X1 U13391 ( .A1(n6442), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n11137), 
        .B2(n14710), .ZN(n10863) );
  NAND2_X1 U13392 ( .A1(n11927), .A2(n14754), .ZN(n10862) );
  OAI211_X1 U13393 ( .C1(n14819), .C2(n14695), .A(n10863), .B(n10862), .ZN(
        n10864) );
  AOI211_X1 U13394 ( .C1(n14825), .C2(n14697), .A(n10865), .B(n10864), .ZN(
        n10866) );
  INV_X1 U13395 ( .A(n10866), .ZN(P1_U3283) );
  OAI211_X1 U13396 ( .C1(n7137), .C2(n14922), .A(n10868), .B(n10867), .ZN(
        n10869) );
  AOI21_X1 U13397 ( .B1(n10870), .B2(n14533), .A(n10869), .ZN(n10874) );
  INV_X1 U13398 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10871) );
  OR2_X1 U13399 ( .A1(n6443), .A2(n10871), .ZN(n10872) );
  OAI21_X1 U13400 ( .B1(n10874), .B2(n14928), .A(n10872), .ZN(P2_U3466) );
  NAND2_X1 U13401 ( .A1(n14931), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n10873) );
  OAI21_X1 U13402 ( .B1(n10874), .B2(n14931), .A(n10873), .ZN(P2_U3511) );
  NAND2_X1 U13403 ( .A1(n11846), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n10882) );
  INV_X1 U13404 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n13755) );
  OR2_X1 U13405 ( .A1(n11818), .A2(n13755), .ZN(n10881) );
  INV_X1 U13406 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10875) );
  OR2_X1 U13407 ( .A1(n11839), .A2(n10875), .ZN(n10880) );
  NAND2_X1 U13408 ( .A1(n10877), .A2(n10876), .ZN(n10878) );
  NAND2_X1 U13409 ( .A1(n11007), .A2(n10878), .ZN(n11018) );
  OR2_X1 U13410 ( .A1(n9605), .A2(n11018), .ZN(n10879) );
  NAND4_X1 U13411 ( .A1(n10882), .A2(n10881), .A3(n10880), .A4(n10879), .ZN(
        n13692) );
  NAND2_X1 U13412 ( .A1(n10883), .A2(n12022), .ZN(n10885) );
  AOI22_X1 U13413 ( .A1(n11627), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n11626), 
        .B2(n13762), .ZN(n10884) );
  XNOR2_X1 U13414 ( .A(n11936), .B(n11405), .ZN(n12044) );
  OR2_X1 U13415 ( .A1(n11927), .A2(n10888), .ZN(n10886) );
  XOR2_X1 U13416 ( .A(n12044), .B(n11003), .Z(n10889) );
  OAI222_X1 U13417 ( .A1(n14720), .A2(n11239), .B1(n10889), .B2(n14744), .C1(
        n14722), .C2(n10888), .ZN(n14551) );
  INV_X1 U13418 ( .A(n14551), .ZN(n10900) );
  AOI21_X1 U13419 ( .B1(n10891), .B2(n13694), .A(n11927), .ZN(n10890) );
  XNOR2_X1 U13420 ( .A(n10998), .B(n12044), .ZN(n14552) );
  OR2_X2 U13421 ( .A1(n10892), .A2(n11927), .ZN(n10893) );
  INV_X1 U13422 ( .A(n10893), .ZN(n10894) );
  INV_X1 U13423 ( .A(n11936), .ZN(n14549) );
  OR2_X2 U13424 ( .A1(n10893), .A2(n11936), .ZN(n11017) );
  OAI211_X1 U13425 ( .C1(n10894), .C2(n14549), .A(n14756), .B(n11017), .ZN(
        n14548) );
  INV_X1 U13426 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10895) );
  OAI22_X1 U13427 ( .A1(n14691), .A2(n10895), .B1(n11236), .B2(n14751), .ZN(
        n10896) );
  AOI21_X1 U13428 ( .B1(n11936), .B2(n14754), .A(n10896), .ZN(n10897) );
  OAI21_X1 U13429 ( .B1(n14548), .B2(n14695), .A(n10897), .ZN(n10898) );
  AOI21_X1 U13430 ( .B1(n14552), .B2(n14697), .A(n10898), .ZN(n10899) );
  OAI21_X1 U13431 ( .B1(n6442), .B2(n10900), .A(n10899), .ZN(P1_U3282) );
  OR2_X1 U13432 ( .A1(n12100), .A2(n10901), .ZN(n10902) );
  XOR2_X1 U13433 ( .A(n11145), .B(n10908), .Z(n10904) );
  AOI22_X1 U13434 ( .A1(n13083), .A2(n13372), .B1(n13370), .B2(n13085), .ZN(
        n13034) );
  OAI21_X1 U13435 ( .B1(n10904), .B2(n13294), .A(n13034), .ZN(n14531) );
  INV_X1 U13436 ( .A(n14531), .ZN(n10916) );
  OR2_X1 U13437 ( .A1(n12100), .A2(n13085), .ZN(n10906) );
  NAND2_X1 U13438 ( .A1(n10907), .A2(n10906), .ZN(n11144) );
  XNOR2_X1 U13439 ( .A(n11144), .B(n10908), .ZN(n14534) );
  INV_X1 U13440 ( .A(n11146), .ZN(n14530) );
  INV_X1 U13441 ( .A(n10909), .ZN(n10910) );
  OAI211_X1 U13442 ( .C1(n14530), .C2(n10910), .A(n13505), .B(n11151), .ZN(
        n14529) );
  INV_X1 U13443 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10911) );
  OAI22_X1 U13444 ( .A1(n13394), .A2(n10911), .B1(n13033), .B2(n13377), .ZN(
        n10912) );
  AOI21_X1 U13445 ( .B1(n11146), .B2(n13381), .A(n10912), .ZN(n10913) );
  OAI21_X1 U13446 ( .B1(n14529), .B2(n13325), .A(n10913), .ZN(n10914) );
  AOI21_X1 U13447 ( .B1(n14534), .B2(n13272), .A(n10914), .ZN(n10915) );
  OAI21_X1 U13448 ( .B1(n10916), .B2(n13426), .A(n10915), .ZN(P2_U3252) );
  XNOR2_X1 U13449 ( .A(n12359), .B(n12153), .ZN(n11050) );
  OAI211_X1 U13450 ( .C1(n10920), .C2(n11050), .A(n11052), .B(n12499), .ZN(
        n10926) );
  OAI22_X1 U13451 ( .A1(n11184), .A2(n12527), .B1(n10921), .B2(n12505), .ZN(
        n10922) );
  AOI211_X1 U13452 ( .C1(n12515), .C2(n10924), .A(n10923), .B(n10922), .ZN(
        n10925) );
  OAI211_X1 U13453 ( .C1(n11120), .C2(n12461), .A(n10926), .B(n10925), .ZN(
        P3_U3153) );
  INV_X1 U13454 ( .A(n10927), .ZN(n10929) );
  OAI222_X1 U13455 ( .A1(P3_U3151), .A2(n10930), .B1(n11500), .B2(n10929), 
        .C1(n10928), .C2(n12933), .ZN(P3_U3271) );
  OAI21_X1 U13456 ( .B1(n10932), .B2(n12222), .A(n10931), .ZN(n11125) );
  NAND2_X1 U13457 ( .A1(n10933), .A2(n12359), .ZN(n11077) );
  OAI211_X1 U13458 ( .C1(n10933), .C2(n12359), .A(n11077), .B(n12766), .ZN(
        n10935) );
  AOI22_X1 U13459 ( .A1(n12553), .A2(n11219), .B1(n12769), .B2(n12551), .ZN(
        n10934) );
  NAND2_X1 U13460 ( .A1(n10935), .A2(n10934), .ZN(n11122) );
  AOI21_X1 U13461 ( .B1(n15150), .B2(n11125), .A(n11122), .ZN(n10941) );
  OAI22_X1 U13462 ( .A1(n12876), .A2(n11121), .B1(n15166), .B2(n8807), .ZN(
        n10936) );
  INV_X1 U13463 ( .A(n10936), .ZN(n10937) );
  OAI21_X1 U13464 ( .B1(n10941), .B2(n15164), .A(n10937), .ZN(P3_U3466) );
  INV_X1 U13465 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n10938) );
  OAI22_X1 U13466 ( .A1(n11121), .A2(n12926), .B1(n15158), .B2(n10938), .ZN(
        n10939) );
  INV_X1 U13467 ( .A(n10939), .ZN(n10940) );
  OAI21_X1 U13468 ( .B1(n10941), .B2(n15157), .A(n10940), .ZN(P3_U3411) );
  INV_X1 U13469 ( .A(n11625), .ZN(n10943) );
  OAI222_X1 U13470 ( .A1(n13796), .A2(P1_U3086), .B1(n14375), .B2(n10943), 
        .C1(n10942), .C2(n14372), .ZN(P1_U3336) );
  OAI222_X1 U13471 ( .A1(n13551), .A2(n10944), .B1(P2_U3088), .B2(n13226), 
        .C1(n13549), .C2(n10943), .ZN(P2_U3308) );
  NAND2_X1 U13472 ( .A1(n10963), .A2(n10945), .ZN(n10947) );
  NAND2_X1 U13473 ( .A1(n10947), .A2(n10946), .ZN(n10949) );
  INV_X1 U13474 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n10960) );
  MUX2_X1 U13475 ( .A(P3_REG1_REG_8__SCAN_IN), .B(n10960), .S(n12609), .Z(
        n10948) );
  NAND2_X1 U13476 ( .A1(n10948), .A2(n10949), .ZN(n12584) );
  OAI21_X1 U13477 ( .B1(n10949), .B2(n10948), .A(n12584), .ZN(n10973) );
  AND2_X1 U13478 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n11056) );
  NOR2_X1 U13479 ( .A1(n10951), .A2(n10950), .ZN(n10954) );
  NOR2_X1 U13480 ( .A1(n10954), .A2(n10953), .ZN(n10957) );
  NAND2_X1 U13481 ( .A1(n12609), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n12560) );
  OAI21_X1 U13482 ( .B1(n12609), .B2(P3_REG2_REG_8__SCAN_IN), .A(n12560), .ZN(
        n10956) );
  INV_X1 U13483 ( .A(n12561), .ZN(n10955) );
  AOI21_X1 U13484 ( .B1(n10957), .B2(n10956), .A(n10955), .ZN(n10958) );
  NOR2_X1 U13485 ( .A1(n15116), .A2(n10958), .ZN(n10959) );
  AOI211_X1 U13486 ( .C1(n15082), .C2(P3_ADDR_REG_8__SCAN_IN), .A(n11056), .B(
        n10959), .ZN(n10971) );
  INV_X1 U13487 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10961) );
  MUX2_X1 U13488 ( .A(n10961), .B(n10960), .S(n12646), .Z(n12611) );
  XNOR2_X1 U13489 ( .A(n12611), .B(n12609), .ZN(n10968) );
  INV_X1 U13490 ( .A(n10962), .ZN(n10966) );
  OAI22_X1 U13491 ( .A1(n10966), .A2(n10965), .B1(n10964), .B2(n10963), .ZN(
        n10967) );
  NAND2_X1 U13492 ( .A1(n10967), .A2(n10968), .ZN(n12612) );
  OAI21_X1 U13493 ( .B1(n10968), .B2(n10967), .A(n12612), .ZN(n10969) );
  NAND2_X1 U13494 ( .A1(n10969), .A2(n15090), .ZN(n10970) );
  OAI211_X1 U13495 ( .C1(n15101), .C2(n12609), .A(n10971), .B(n10970), .ZN(
        n10972) );
  AOI21_X1 U13496 ( .B1(n15107), .B2(n10973), .A(n10972), .ZN(n10974) );
  INV_X1 U13497 ( .A(n10974), .ZN(P3_U3190) );
  NAND2_X1 U13498 ( .A1(n11923), .A2(n11807), .ZN(n10979) );
  NAND2_X1 U13499 ( .A1(n14683), .A2(n11775), .ZN(n10978) );
  NAND2_X1 U13500 ( .A1(n10979), .A2(n10978), .ZN(n10980) );
  XNOR2_X1 U13501 ( .A(n10980), .B(n10326), .ZN(n11127) );
  AND2_X1 U13502 ( .A1(n14683), .A2(n11808), .ZN(n10981) );
  AOI21_X1 U13503 ( .B1(n11923), .B2(n11775), .A(n10981), .ZN(n11128) );
  XNOR2_X1 U13504 ( .A(n11127), .B(n11128), .ZN(n10982) );
  OAI211_X1 U13505 ( .C1(n10983), .C2(n10982), .A(n11131), .B(n13645), .ZN(
        n10990) );
  INV_X1 U13506 ( .A(n10984), .ZN(n10986) );
  AOI21_X1 U13507 ( .B1(n13664), .B2(n10986), .A(n10985), .ZN(n10987) );
  OAI21_X1 U13508 ( .B1(n13667), .B2(n10752), .A(n10987), .ZN(n10988) );
  AOI21_X1 U13509 ( .B1(n6433), .B2(n13694), .A(n10988), .ZN(n10989) );
  OAI211_X1 U13510 ( .C1(n14815), .C2(n13652), .A(n10990), .B(n10989), .ZN(
        P1_U3231) );
  OAI22_X1 U13511 ( .A1(n12815), .A2(n10992), .B1(n10991), .B2(n12816), .ZN(
        n10995) );
  MUX2_X1 U13512 ( .A(n10993), .B(P3_REG2_REG_6__SCAN_IN), .S(n15136), .Z(
        n10994) );
  AOI211_X1 U13513 ( .C1(n12821), .C2(n10996), .A(n10995), .B(n10994), .ZN(
        n10997) );
  INV_X1 U13514 ( .A(n10997), .ZN(P3_U3227) );
  NAND2_X1 U13515 ( .A1(n10999), .A2(n12022), .ZN(n11001) );
  AOI22_X1 U13516 ( .A1(n11627), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n11626), 
        .B2(n13782), .ZN(n11000) );
  XNOR2_X1 U13517 ( .A(n11939), .B(n11239), .ZN(n12045) );
  OAI21_X1 U13518 ( .B1(n11002), .B2(n12045), .A(n11024), .ZN(n11173) );
  INV_X1 U13519 ( .A(n12045), .ZN(n11032) );
  XNOR2_X1 U13520 ( .A(n11033), .B(n11032), .ZN(n11004) );
  NOR2_X1 U13521 ( .A1(n11004), .A2(n14744), .ZN(n11016) );
  NAND2_X1 U13522 ( .A1(n11845), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11014) );
  INV_X1 U13523 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11005) );
  OR2_X1 U13524 ( .A1(n11839), .A2(n11005), .ZN(n11013) );
  INV_X1 U13525 ( .A(n11038), .ZN(n11009) );
  NAND2_X1 U13526 ( .A1(n11007), .A2(n11006), .ZN(n11008) );
  NAND2_X1 U13527 ( .A1(n11009), .A2(n11008), .ZN(n11458) );
  OR2_X1 U13528 ( .A1(n9605), .A2(n11458), .ZN(n11012) );
  INV_X1 U13529 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11010) );
  OR2_X1 U13530 ( .A1(n11816), .A2(n11010), .ZN(n11011) );
  NAND4_X1 U13531 ( .A1(n11014), .A2(n11013), .A3(n11012), .A4(n11011), .ZN(
        n14086) );
  INV_X1 U13532 ( .A(n14086), .ZN(n11947) );
  OAI22_X1 U13533 ( .A1(n11947), .A2(n14720), .B1(n11405), .B2(n14722), .ZN(
        n11015) );
  AOI211_X1 U13534 ( .C1(n11173), .C2(n14749), .A(n11016), .B(n11015), .ZN(
        n11176) );
  INV_X1 U13535 ( .A(n11939), .ZN(n11409) );
  AOI211_X1 U13536 ( .C1(n11939), .C2(n11017), .A(n14090), .B(n11029), .ZN(
        n11174) );
  NAND2_X1 U13537 ( .A1(n11174), .A2(n14759), .ZN(n11020) );
  INV_X1 U13538 ( .A(n11018), .ZN(n11403) );
  AOI22_X1 U13539 ( .A1(n6442), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n11403), 
        .B2(n14710), .ZN(n11019) );
  OAI211_X1 U13540 ( .C1(n11409), .C2(n14047), .A(n11020), .B(n11019), .ZN(
        n11021) );
  AOI21_X1 U13541 ( .B1(n11173), .B2(n14760), .A(n11021), .ZN(n11022) );
  OAI21_X1 U13542 ( .B1(n11176), .B2(n6442), .A(n11022), .ZN(P1_U3281) );
  NAND2_X1 U13543 ( .A1(n11024), .A2(n11023), .ZN(n11028) );
  OR2_X1 U13544 ( .A1(n11025), .A2(n11610), .ZN(n11027) );
  AOI22_X1 U13545 ( .A1(n11627), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n11626), 
        .B2(n14610), .ZN(n11026) );
  XNOR2_X1 U13546 ( .A(n11946), .B(n11947), .ZN(n12047) );
  NAND2_X1 U13547 ( .A1(n11028), .A2(n12047), .ZN(n11284) );
  OAI21_X1 U13548 ( .B1(n11028), .B2(n12047), .A(n11284), .ZN(n14547) );
  INV_X1 U13549 ( .A(n14547), .ZN(n11049) );
  OAI22_X1 U13550 ( .A1(n14691), .A2(n11005), .B1(n11458), .B2(n14751), .ZN(
        n11031) );
  OAI211_X1 U13551 ( .C1(n11029), .C2(n14544), .A(n14091), .B(n14756), .ZN(
        n14543) );
  NOR2_X1 U13552 ( .A1(n14543), .A2(n14695), .ZN(n11030) );
  AOI211_X1 U13553 ( .C1(n14754), .C2(n11946), .A(n11031), .B(n11030), .ZN(
        n11048) );
  NAND2_X1 U13554 ( .A1(n11033), .A2(n11032), .ZN(n11035) );
  OR2_X1 U13555 ( .A1(n11939), .A2(n11239), .ZN(n11034) );
  INV_X1 U13556 ( .A(n12047), .ZN(n11300) );
  XNOR2_X1 U13557 ( .A(n11301), .B(n11300), .ZN(n11036) );
  NOR2_X1 U13558 ( .A1(n11036), .A2(n14744), .ZN(n14546) );
  NAND2_X1 U13559 ( .A1(n11846), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n11043) );
  INV_X1 U13560 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11037) );
  OR2_X1 U13561 ( .A1(n11839), .A2(n11037), .ZN(n11042) );
  NOR2_X1 U13562 ( .A1(n11038), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n11039) );
  OR2_X1 U13563 ( .A1(n11288), .A2(n11039), .ZN(n14080) );
  OR2_X1 U13564 ( .A1(n9605), .A2(n14080), .ZN(n11041) );
  INV_X1 U13565 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n13779) );
  OR2_X1 U13566 ( .A1(n11818), .A2(n13779), .ZN(n11040) );
  OR2_X1 U13567 ( .A1(n11585), .A2(n14720), .ZN(n11045) );
  NAND2_X1 U13568 ( .A1(n13692), .A2(n14705), .ZN(n11044) );
  AND2_X1 U13569 ( .A1(n11045), .A2(n11044), .ZN(n14542) );
  INV_X1 U13570 ( .A(n14542), .ZN(n11046) );
  OAI21_X1 U13571 ( .B1(n14546), .B2(n11046), .A(n14691), .ZN(n11047) );
  OAI211_X1 U13572 ( .C1(n11049), .C2(n14059), .A(n11048), .B(n11047), .ZN(
        P1_U3280) );
  XNOR2_X1 U13573 ( .A(n12230), .B(n12180), .ZN(n11180) );
  XNOR2_X1 U13574 ( .A(n11180), .B(n12551), .ZN(n11053) );
  OAI211_X1 U13575 ( .C1(n11054), .C2(n11053), .A(n11179), .B(n12499), .ZN(
        n11058) );
  OAI22_X1 U13576 ( .A1(n11081), .A2(n12505), .B1(n11257), .B2(n12527), .ZN(
        n11055) );
  AOI211_X1 U13577 ( .C1(n12515), .C2(n12230), .A(n11056), .B(n11055), .ZN(
        n11057) );
  OAI211_X1 U13578 ( .C1(n11082), .C2(n12461), .A(n11058), .B(n11057), .ZN(
        P3_U3161) );
  NAND2_X1 U13579 ( .A1(n11074), .A2(n12365), .ZN(n11073) );
  NAND2_X1 U13580 ( .A1(n11073), .A2(n11059), .ZN(n11091) );
  NAND2_X1 U13581 ( .A1(n11091), .A2(n11060), .ZN(n11062) );
  NAND2_X1 U13582 ( .A1(n11062), .A2(n11061), .ZN(n11063) );
  INV_X1 U13583 ( .A(n12243), .ZN(n12366) );
  XNOR2_X1 U13584 ( .A(n11063), .B(n12366), .ZN(n15151) );
  INV_X1 U13585 ( .A(n15151), .ZN(n11072) );
  OAI211_X1 U13586 ( .C1(n11065), .C2(n12243), .A(n11064), .B(n12766), .ZN(
        n11067) );
  AOI22_X1 U13587 ( .A1(n12234), .A2(n11219), .B1(n12769), .B2(n12549), .ZN(
        n11066) );
  NAND2_X1 U13588 ( .A1(n11067), .A2(n11066), .ZN(n15156) );
  NAND2_X1 U13589 ( .A1(n15156), .A2(n12818), .ZN(n11071) );
  OAI22_X1 U13590 ( .A1(n12815), .A2(n11068), .B1(n11262), .B2(n12816), .ZN(
        n11069) );
  AOI21_X1 U13591 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n15136), .A(n11069), 
        .ZN(n11070) );
  OAI211_X1 U13592 ( .C1(n12666), .C2(n11072), .A(n11071), .B(n11070), .ZN(
        P3_U3223) );
  OAI21_X1 U13593 ( .B1(n11074), .B2(n12365), .A(n11073), .ZN(n11161) );
  INV_X1 U13594 ( .A(n11161), .ZN(n11086) );
  NAND2_X1 U13595 ( .A1(n11077), .A2(n11075), .ZN(n11079) );
  AND2_X1 U13596 ( .A1(n11077), .A2(n11076), .ZN(n11078) );
  AOI21_X1 U13597 ( .B1(n12365), .B2(n11079), .A(n11078), .ZN(n11080) );
  OAI222_X1 U13598 ( .A1(n15122), .A2(n11257), .B1(n12799), .B2(n11081), .C1(
        n15128), .C2(n11080), .ZN(n11160) );
  NAND2_X1 U13599 ( .A1(n11160), .A2(n12818), .ZN(n11085) );
  OAI22_X1 U13600 ( .A1(n12815), .A2(n12229), .B1(n11082), .B2(n12816), .ZN(
        n11083) );
  AOI21_X1 U13601 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n15136), .A(n11083), .ZN(
        n11084) );
  OAI211_X1 U13602 ( .C1(n11086), .C2(n12666), .A(n11085), .B(n11084), .ZN(
        P3_U3225) );
  INV_X1 U13603 ( .A(n11715), .ZN(n11089) );
  OAI222_X1 U13604 ( .A1(n13551), .A2(n11088), .B1(n13549), .B2(n11089), .C1(
        n11087), .C2(P2_U3088), .ZN(P2_U3303) );
  INV_X1 U13605 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11716) );
  OAI222_X1 U13606 ( .A1(P1_U3086), .A2(n11090), .B1(n14375), .B2(n11089), 
        .C1(n11716), .C2(n14372), .ZN(P1_U3331) );
  XNOR2_X1 U13607 ( .A(n11091), .B(n12360), .ZN(n15147) );
  NAND2_X1 U13608 ( .A1(n12818), .A2(n15131), .ZN(n11519) );
  INV_X1 U13609 ( .A(n15125), .ZN(n11513) );
  OAI211_X1 U13610 ( .C1(n11093), .C2(n12360), .A(n11092), .B(n12766), .ZN(
        n11095) );
  AOI22_X1 U13611 ( .A1(n12550), .A2(n12769), .B1(n11219), .B2(n12551), .ZN(
        n11094) );
  OAI211_X1 U13612 ( .C1(n15147), .C2(n11513), .A(n11095), .B(n11094), .ZN(
        n15149) );
  NAND2_X1 U13613 ( .A1(n15149), .A2(n12818), .ZN(n11098) );
  OAI22_X1 U13614 ( .A1(n12815), .A2(n15145), .B1(n11186), .B2(n12816), .ZN(
        n11096) );
  AOI21_X1 U13615 ( .B1(n15136), .B2(P3_REG2_REG_9__SCAN_IN), .A(n11096), .ZN(
        n11097) );
  OAI211_X1 U13616 ( .C1(n15147), .C2(n11519), .A(n11098), .B(n11097), .ZN(
        P3_U3224) );
  INV_X1 U13617 ( .A(n11659), .ZN(n11100) );
  INV_X1 U13618 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11660) );
  OAI222_X1 U13619 ( .A1(P1_U3086), .A2(n9260), .B1(n14375), .B2(n11100), .C1(
        n11660), .C2(n14372), .ZN(P1_U3334) );
  OAI222_X1 U13620 ( .A1(n13551), .A2(n11101), .B1(n13549), .B2(n11100), .C1(
        n11099), .C2(P2_U3088), .ZN(P2_U3306) );
  INV_X1 U13621 ( .A(n11647), .ZN(n11103) );
  OAI222_X1 U13622 ( .A1(P1_U3086), .A2(n11853), .B1(n14375), .B2(n11103), 
        .C1(n11648), .C2(n14372), .ZN(P1_U3335) );
  OAI222_X1 U13623 ( .A1(n13551), .A2(n11104), .B1(n13549), .B2(n11103), .C1(
        n11102), .C2(P2_U3088), .ZN(P2_U3307) );
  INV_X1 U13624 ( .A(n11105), .ZN(n11112) );
  OAI21_X1 U13625 ( .B1(n11112), .B2(P2_REG2_REG_12__SCAN_IN), .A(n11106), 
        .ZN(n14865) );
  MUX2_X1 U13626 ( .A(n10911), .B(P2_REG2_REG_13__SCAN_IN), .S(n14861), .Z(
        n14866) );
  NOR2_X1 U13627 ( .A1(n14865), .A2(n14866), .ZN(n14863) );
  AOI21_X1 U13628 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n14861), .A(n14863), 
        .ZN(n11108) );
  NAND2_X1 U13629 ( .A1(n11108), .A2(n11107), .ZN(n13153) );
  OAI21_X1 U13630 ( .B1(n11108), .B2(n11107), .A(n13153), .ZN(n11109) );
  NOR2_X1 U13631 ( .A1(n11109), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n13155) );
  AOI21_X1 U13632 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n11109), .A(n13155), 
        .ZN(n11119) );
  INV_X1 U13633 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n11110) );
  NAND2_X1 U13634 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14509)
         );
  OAI21_X1 U13635 ( .B1(n14871), .B2(n11110), .A(n14509), .ZN(n11117) );
  OAI21_X1 U13636 ( .B1(n11112), .B2(P2_REG1_REG_12__SCAN_IN), .A(n11111), 
        .ZN(n14857) );
  INV_X1 U13637 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11113) );
  MUX2_X1 U13638 ( .A(n11113), .B(P2_REG1_REG_13__SCAN_IN), .S(n14861), .Z(
        n14858) );
  NOR2_X1 U13639 ( .A1(n14857), .A2(n14858), .ZN(n14855) );
  XNOR2_X1 U13640 ( .A(n13148), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n11114) );
  AOI211_X1 U13641 ( .C1(n11115), .C2(n11114), .A(n14856), .B(n13147), .ZN(
        n11116) );
  AOI211_X1 U13642 ( .C1(n14862), .C2(n13148), .A(n11117), .B(n11116), .ZN(
        n11118) );
  OAI21_X1 U13643 ( .B1(n11119), .B2(n14864), .A(n11118), .ZN(P2_U3228) );
  OAI22_X1 U13644 ( .A1(n12815), .A2(n11121), .B1(n11120), .B2(n12816), .ZN(
        n11124) );
  MUX2_X1 U13645 ( .A(n11122), .B(P3_REG2_REG_7__SCAN_IN), .S(n15136), .Z(
        n11123) );
  AOI211_X1 U13646 ( .C1(n12821), .C2(n11125), .A(n11124), .B(n11123), .ZN(
        n11126) );
  INV_X1 U13647 ( .A(n11126), .ZN(P3_U3226) );
  INV_X1 U13648 ( .A(n11128), .ZN(n11129) );
  AND2_X1 U13649 ( .A1(n13694), .A2(n11808), .ZN(n11132) );
  AOI21_X1 U13650 ( .B1(n11927), .B2(n11775), .A(n11132), .ZN(n11229) );
  AOI22_X1 U13651 ( .A1(n11927), .A2(n11807), .B1(n11775), .B2(n13694), .ZN(
        n11133) );
  XNOR2_X1 U13652 ( .A(n11133), .B(n10326), .ZN(n11230) );
  XOR2_X1 U13653 ( .A(n11229), .B(n11230), .Z(n11134) );
  OAI211_X1 U13654 ( .C1(n11135), .C2(n11134), .A(n11232), .B(n13645), .ZN(
        n11142) );
  NOR2_X1 U13655 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11136), .ZN(n14598) );
  AOI21_X1 U13656 ( .B1(n13664), .B2(n11137), .A(n14598), .ZN(n11138) );
  OAI21_X1 U13657 ( .B1(n13667), .B2(n11139), .A(n11138), .ZN(n11140) );
  AOI21_X1 U13658 ( .B1(n6433), .B2(n13693), .A(n11140), .ZN(n11141) );
  OAI211_X1 U13659 ( .C1(n14822), .C2(n13652), .A(n11142), .B(n11141), .ZN(
        P1_U3217) );
  NOR2_X1 U13660 ( .A1(n11146), .A2(n13084), .ZN(n11143) );
  XNOR2_X1 U13661 ( .A(n11210), .B(n11149), .ZN(n13515) );
  INV_X1 U13662 ( .A(n11199), .ZN(n11147) );
  AOI21_X1 U13663 ( .B1(n11149), .B2(n11148), .A(n11147), .ZN(n11150) );
  OAI222_X1 U13664 ( .A1(n13052), .A2(n14520), .B1(n13051), .B2(n14499), .C1(
        n13294), .C2(n11150), .ZN(n13511) );
  NAND2_X1 U13665 ( .A1(n14508), .A2(n11151), .ZN(n11152) );
  NAND2_X1 U13666 ( .A1(n11152), .A2(n13505), .ZN(n11153) );
  NOR2_X1 U13667 ( .A1(n6490), .A2(n11153), .ZN(n13512) );
  NAND2_X1 U13668 ( .A1(n13512), .A2(n13424), .ZN(n11157) );
  INV_X1 U13669 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n11154) );
  OAI22_X1 U13670 ( .A1(n13394), .A2(n11154), .B1(n14511), .B2(n13377), .ZN(
        n11155) );
  AOI21_X1 U13671 ( .B1(n14508), .B2(n13381), .A(n11155), .ZN(n11156) );
  NAND2_X1 U13672 ( .A1(n11157), .A2(n11156), .ZN(n11158) );
  AOI21_X1 U13673 ( .B1(n13511), .B2(n13394), .A(n11158), .ZN(n11159) );
  OAI21_X1 U13674 ( .B1(n13421), .B2(n13515), .A(n11159), .ZN(P2_U3251) );
  AOI21_X1 U13675 ( .B1(n15150), .B2(n11161), .A(n11160), .ZN(n11167) );
  OAI22_X1 U13676 ( .A1(n12876), .A2(n12229), .B1(n15166), .B2(n10960), .ZN(
        n11162) );
  INV_X1 U13677 ( .A(n11162), .ZN(n11163) );
  OAI21_X1 U13678 ( .B1(n11167), .B2(n15164), .A(n11163), .ZN(P3_U3467) );
  INV_X1 U13679 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n11164) );
  OAI22_X1 U13680 ( .A1(n12229), .A2(n12926), .B1(n15158), .B2(n11164), .ZN(
        n11165) );
  INV_X1 U13681 ( .A(n11165), .ZN(n11166) );
  OAI21_X1 U13682 ( .B1(n11167), .B2(n15157), .A(n11166), .ZN(P3_U3414) );
  INV_X1 U13683 ( .A(n11168), .ZN(n11169) );
  INV_X1 U13684 ( .A(n11737), .ZN(n11171) );
  OAI222_X1 U13685 ( .A1(P1_U3086), .A2(n11169), .B1(n14375), .B2(n11171), 
        .C1(n11738), .C2(n14372), .ZN(P1_U3330) );
  OAI222_X1 U13686 ( .A1(n13551), .A2(n11172), .B1(n13549), .B2(n11171), .C1(
        n11170), .C2(P2_U3088), .ZN(P2_U3302) );
  INV_X1 U13687 ( .A(n11173), .ZN(n11177) );
  AOI21_X1 U13688 ( .B1(n11939), .B2(n14792), .A(n11174), .ZN(n11175) );
  OAI211_X1 U13689 ( .C1(n11177), .C2(n14797), .A(n11176), .B(n11175), .ZN(
        n11191) );
  NAND2_X1 U13690 ( .A1(n11191), .A2(n14839), .ZN(n11178) );
  OAI21_X1 U13691 ( .B1(n14839), .B2(n13755), .A(n11178), .ZN(P1_U3540) );
  XNOR2_X1 U13692 ( .A(n15145), .B(n12180), .ZN(n11252) );
  XNOR2_X1 U13693 ( .A(n12234), .B(n11252), .ZN(n11182) );
  OAI21_X1 U13694 ( .B1(n11184), .B2(n11180), .A(n11179), .ZN(n11181) );
  NOR2_X2 U13695 ( .A1(n11181), .A2(n11182), .ZN(n11254) );
  AOI21_X1 U13696 ( .B1(n11182), .B2(n11181), .A(n11254), .ZN(n11190) );
  NOR2_X1 U13697 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11183), .ZN(n15017) );
  OAI22_X1 U13698 ( .A1(n11184), .A2(n12505), .B1(n11245), .B2(n12527), .ZN(
        n11185) );
  AOI211_X1 U13699 ( .C1(n12515), .C2(n12235), .A(n15017), .B(n11185), .ZN(
        n11189) );
  INV_X1 U13700 ( .A(n11186), .ZN(n11187) );
  NAND2_X1 U13701 ( .A1(n12531), .A2(n11187), .ZN(n11188) );
  OAI211_X1 U13702 ( .C1(n11190), .C2(n12534), .A(n11189), .B(n11188), .ZN(
        P3_U3171) );
  INV_X1 U13703 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11193) );
  NAND2_X1 U13704 ( .A1(n11191), .A2(n14827), .ZN(n11192) );
  OAI21_X1 U13705 ( .B1(n14827), .B2(n11193), .A(n11192), .ZN(P1_U3495) );
  INV_X1 U13706 ( .A(n11194), .ZN(n11196) );
  OAI222_X1 U13707 ( .A1(P3_U3151), .A2(n11197), .B1(n11500), .B2(n11196), 
        .C1(n11195), .C2(n12933), .ZN(P3_U3269) );
  NAND2_X1 U13708 ( .A1(n11276), .A2(n7204), .ZN(n11275) );
  NAND2_X1 U13709 ( .A1(n11273), .A2(n14520), .ZN(n11200) );
  XNOR2_X1 U13710 ( .A(n11387), .B(n11212), .ZN(n11202) );
  NAND2_X1 U13711 ( .A1(n11202), .A2(n13406), .ZN(n11204) );
  AOI22_X1 U13712 ( .A1(n13080), .A2(n13372), .B1(n13370), .B2(n13082), .ZN(
        n11203) );
  NAND2_X1 U13713 ( .A1(n11204), .A2(n11203), .ZN(n13510) );
  INV_X1 U13714 ( .A(n13510), .ZN(n11216) );
  NAND2_X1 U13715 ( .A1(n11322), .A2(n6490), .ZN(n11269) );
  NAND2_X1 U13716 ( .A1(n11269), .A2(n13504), .ZN(n11205) );
  AND2_X1 U13717 ( .A1(n11384), .A2(n11205), .ZN(n13506) );
  OAI22_X1 U13718 ( .A1(n13394), .A2(n13188), .B1(n14527), .B2(n13377), .ZN(
        n11207) );
  INV_X1 U13719 ( .A(n13504), .ZN(n14516) );
  NOR2_X1 U13720 ( .A1(n14516), .A2(n13415), .ZN(n11206) );
  AOI211_X1 U13721 ( .C1(n13506), .C2(n13385), .A(n11207), .B(n11206), .ZN(
        n11215) );
  AND2_X1 U13722 ( .A1(n14508), .A2(n13083), .ZN(n11209) );
  OR2_X1 U13723 ( .A1(n14508), .A2(n13083), .ZN(n11208) );
  NAND2_X1 U13724 ( .A1(n11213), .A2(n11212), .ZN(n13502) );
  NAND3_X1 U13725 ( .A1(n13503), .A2(n13502), .A3(n13272), .ZN(n11214) );
  OAI211_X1 U13726 ( .C1(n11216), .C2(n13426), .A(n11215), .B(n11214), .ZN(
        P2_U3249) );
  XNOR2_X1 U13727 ( .A(n11217), .B(n11222), .ZN(n11218) );
  NAND2_X1 U13728 ( .A1(n11218), .A2(n12766), .ZN(n11221) );
  AOI22_X1 U13729 ( .A1(n11219), .A2(n12549), .B1(n11485), .B2(n12769), .ZN(
        n11220) );
  XNOR2_X1 U13730 ( .A(n11223), .B(n11222), .ZN(n14488) );
  NOR2_X1 U13731 ( .A1(n12815), .A2(n11224), .ZN(n11226) );
  OAI22_X1 U13732 ( .A1(n12818), .A2(n12620), .B1(n11488), .B2(n12816), .ZN(
        n11225) );
  AOI211_X1 U13733 ( .C1(n14488), .C2(n12821), .A(n11226), .B(n11225), .ZN(
        n11227) );
  OAI21_X1 U13734 ( .B1(n14490), .B2(n15136), .A(n11227), .ZN(P3_U3221) );
  AOI22_X1 U13735 ( .A1(n11936), .A2(n11807), .B1(n11775), .B2(n13693), .ZN(
        n11228) );
  XNOR2_X1 U13736 ( .A(n11228), .B(n10326), .ZN(n11397) );
  AOI22_X1 U13737 ( .A1(n11936), .A2(n11775), .B1(n11808), .B2(n13693), .ZN(
        n11398) );
  XNOR2_X1 U13738 ( .A(n11397), .B(n11398), .ZN(n11234) );
  AOI21_X1 U13739 ( .B1(n11234), .B2(n11233), .A(n11396), .ZN(n11242) );
  OAI21_X1 U13740 ( .B1(n13679), .B2(n11236), .A(n11235), .ZN(n11237) );
  AOI21_X1 U13741 ( .B1(n13681), .B2(n13694), .A(n11237), .ZN(n11238) );
  OAI21_X1 U13742 ( .B1(n11239), .B2(n13683), .A(n11238), .ZN(n11240) );
  AOI21_X1 U13743 ( .B1(n11936), .B2(n13685), .A(n11240), .ZN(n11241) );
  OAI21_X1 U13744 ( .B1(n11242), .B2(n13688), .A(n11241), .ZN(P1_U3236) );
  XOR2_X1 U13745 ( .A(n12374), .B(n11243), .Z(n11244) );
  OAI222_X1 U13746 ( .A1(n12799), .A2(n11245), .B1(n15122), .B2(n11423), .C1(
        n11244), .C2(n15128), .ZN(n11369) );
  INV_X1 U13747 ( .A(n11369), .ZN(n11251) );
  OAI21_X1 U13748 ( .B1(n11246), .B2(n12374), .A(n11247), .ZN(n11370) );
  INV_X1 U13749 ( .A(n12246), .ZN(n11437) );
  NOR2_X1 U13750 ( .A1(n12815), .A2(n11437), .ZN(n11249) );
  OAI22_X1 U13751 ( .A1(n12818), .A2(n12602), .B1(n11433), .B2(n12816), .ZN(
        n11248) );
  AOI211_X1 U13752 ( .C1(n11370), .C2(n12821), .A(n11249), .B(n11248), .ZN(
        n11250) );
  OAI21_X1 U13753 ( .B1(n11251), .B2(n15136), .A(n11250), .ZN(P3_U3222) );
  NOR2_X1 U13754 ( .A1(n12234), .A2(n11252), .ZN(n11253) );
  XNOR2_X1 U13755 ( .A(n15153), .B(n12180), .ZN(n11410) );
  XNOR2_X1 U13756 ( .A(n12550), .B(n11410), .ZN(n11255) );
  OAI211_X1 U13757 ( .C1(n11256), .C2(n11255), .A(n11413), .B(n12499), .ZN(
        n11261) );
  NAND2_X1 U13758 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n15032)
         );
  INV_X1 U13759 ( .A(n15032), .ZN(n11259) );
  OAI22_X1 U13760 ( .A1(n7425), .A2(n12527), .B1(n11257), .B2(n12505), .ZN(
        n11258) );
  AOI211_X1 U13761 ( .C1(n15153), .C2(n12515), .A(n11259), .B(n11258), .ZN(
        n11260) );
  OAI211_X1 U13762 ( .C1(n11262), .C2(n12461), .A(n11261), .B(n11260), .ZN(
        P3_U3157) );
  INV_X1 U13763 ( .A(n11263), .ZN(n11265) );
  OAI222_X1 U13764 ( .A1(n13551), .A2(n11266), .B1(n13549), .B2(n11265), .C1(
        n11264), .C2(P2_U3088), .ZN(P2_U3305) );
  XNOR2_X1 U13765 ( .A(n11268), .B(n11267), .ZN(n11324) );
  OAI211_X1 U13766 ( .C1(n11322), .C2(n6490), .A(n13505), .B(n11269), .ZN(
        n11320) );
  OAI22_X1 U13767 ( .A1(n13394), .A2(n11271), .B1(n11270), .B2(n13377), .ZN(
        n11272) );
  AOI21_X1 U13768 ( .B1(n11273), .B2(n13381), .A(n11272), .ZN(n11274) );
  OAI21_X1 U13769 ( .B1(n11320), .B2(n13325), .A(n11274), .ZN(n11279) );
  OAI21_X1 U13770 ( .B1(n11276), .B2(n7204), .A(n11275), .ZN(n11277) );
  AOI222_X1 U13771 ( .A1(n13406), .A2(n11277), .B1(n13081), .B2(n13372), .C1(
        n13083), .C2(n13370), .ZN(n11321) );
  NOR2_X1 U13772 ( .A1(n11321), .A2(n13426), .ZN(n11278) );
  AOI211_X1 U13773 ( .C1(n11324), .C2(n13272), .A(n11279), .B(n11278), .ZN(
        n11280) );
  INV_X1 U13774 ( .A(n11280), .ZN(P2_U3250) );
  NAND2_X1 U13775 ( .A1(n11281), .A2(n12022), .ZN(n11283) );
  AOI22_X1 U13776 ( .A1(n11627), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n11626), 
        .B2(n13783), .ZN(n11282) );
  INV_X1 U13777 ( .A(n11585), .ZN(n13691) );
  NAND2_X1 U13778 ( .A1(n14194), .A2(n11585), .ZN(n11950) );
  NAND2_X1 U13779 ( .A1(n11951), .A2(n11950), .ZN(n14082) );
  INV_X1 U13780 ( .A(n14082), .ZN(n14078) );
  NAND2_X1 U13781 ( .A1(n11285), .A2(n12022), .ZN(n11287) );
  INV_X1 U13782 ( .A(n13786), .ZN(n14635) );
  AOI22_X1 U13783 ( .A1(n11627), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n11626), 
        .B2(n14635), .ZN(n11286) );
  NAND2_X1 U13784 ( .A1(n11845), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n11294) );
  INV_X1 U13785 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11296) );
  OR2_X1 U13786 ( .A1(n11839), .A2(n11296), .ZN(n11293) );
  OR2_X1 U13787 ( .A1(n11288), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n11289) );
  NAND2_X1 U13788 ( .A1(n11309), .A2(n11289), .ZN(n13678) );
  OR2_X1 U13789 ( .A1(n9605), .A2(n13678), .ZN(n11292) );
  INV_X1 U13790 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n11290) );
  OR2_X1 U13791 ( .A1(n11816), .A2(n11290), .ZN(n11291) );
  NAND2_X1 U13792 ( .A1(n13686), .A2(n14085), .ZN(n11955) );
  NAND2_X1 U13793 ( .A1(n11954), .A2(n11955), .ZN(n12049) );
  OAI21_X1 U13794 ( .B1(n11295), .B2(n12049), .A(n11341), .ZN(n14541) );
  INV_X1 U13795 ( .A(n14541), .ZN(n11319) );
  OAI22_X1 U13796 ( .A1(n14691), .A2(n11296), .B1(n13678), .B2(n14751), .ZN(
        n11299) );
  INV_X1 U13797 ( .A(n13686), .ZN(n14538) );
  AOI21_X1 U13798 ( .B1(n13686), .B2(n14092), .A(n14090), .ZN(n11297) );
  NAND2_X1 U13799 ( .A1(n11346), .A2(n11297), .ZN(n14537) );
  NOR2_X1 U13800 ( .A1(n14537), .A2(n14695), .ZN(n11298) );
  AOI211_X1 U13801 ( .C1(n14754), .C2(n13686), .A(n11299), .B(n11298), .ZN(
        n11318) );
  NAND2_X1 U13802 ( .A1(n11301), .A2(n11300), .ZN(n11303) );
  OR2_X1 U13803 ( .A1(n11946), .A2(n11947), .ZN(n11302) );
  INV_X1 U13804 ( .A(n11951), .ZN(n11304) );
  INV_X1 U13805 ( .A(n11351), .ZN(n11305) );
  AOI211_X1 U13806 ( .C1(n12049), .C2(n11306), .A(n14744), .B(n11305), .ZN(
        n14540) );
  NAND2_X1 U13807 ( .A1(n11814), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11315) );
  INV_X1 U13808 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n11307) );
  OR2_X1 U13809 ( .A1(n11818), .A2(n11307), .ZN(n11314) );
  INV_X1 U13810 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n11308) );
  NAND2_X1 U13811 ( .A1(n11309), .A2(n11308), .ZN(n11310) );
  NAND2_X1 U13812 ( .A1(n11356), .A2(n11310), .ZN(n13614) );
  OR2_X1 U13813 ( .A1(n9605), .A2(n13614), .ZN(n11313) );
  INV_X1 U13814 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n11311) );
  OR2_X1 U13815 ( .A1(n11816), .A2(n11311), .ZN(n11312) );
  NAND4_X1 U13816 ( .A1(n11315), .A2(n11314), .A3(n11313), .A4(n11312), .ZN(
        n14064) );
  AOI22_X1 U13817 ( .A1(n13691), .A2(n14705), .B1(n14702), .B2(n14064), .ZN(
        n14536) );
  INV_X1 U13818 ( .A(n14536), .ZN(n11316) );
  OAI21_X1 U13819 ( .B1(n14540), .B2(n11316), .A(n14691), .ZN(n11317) );
  OAI211_X1 U13820 ( .C1(n11319), .C2(n14059), .A(n11318), .B(n11317), .ZN(
        P1_U3278) );
  OAI211_X1 U13821 ( .C1(n11322), .C2(n14922), .A(n11321), .B(n11320), .ZN(
        n11323) );
  AOI21_X1 U13822 ( .B1(n11324), .B2(n14533), .A(n11323), .ZN(n11327) );
  NAND2_X1 U13823 ( .A1(n14931), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n11325) );
  OAI21_X1 U13824 ( .B1(n11327), .B2(n14931), .A(n11325), .ZN(P2_U3514) );
  NAND2_X1 U13825 ( .A1(n14928), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n11326) );
  OAI21_X1 U13826 ( .B1(n11327), .B2(n14928), .A(n11326), .ZN(P2_U3475) );
  INV_X1 U13827 ( .A(n11697), .ZN(n11330) );
  AOI21_X1 U13828 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n13541), .A(n11328), 
        .ZN(n11329) );
  OAI21_X1 U13829 ( .B1(n11330), .B2(n13549), .A(n11329), .ZN(P2_U3304) );
  INV_X1 U13830 ( .A(n11331), .ZN(n11333) );
  OAI222_X1 U13831 ( .A1(P3_U3151), .A2(n12646), .B1(n11500), .B2(n11333), 
        .C1(n11332), .C2(n12933), .ZN(P3_U3268) );
  INV_X1 U13832 ( .A(n11334), .ZN(n11335) );
  INV_X1 U13833 ( .A(n11759), .ZN(n11337) );
  OAI222_X1 U13834 ( .A1(n11335), .A2(P1_U3086), .B1(n14375), .B2(n11337), 
        .C1(n11760), .C2(n14372), .ZN(P1_U3329) );
  OAI222_X1 U13835 ( .A1(n11338), .A2(P2_U3088), .B1(n13549), .B2(n11337), 
        .C1(n11336), .C2(n13551), .ZN(P2_U3301) );
  INV_X1 U13836 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11698) );
  NAND2_X1 U13837 ( .A1(n11697), .A2(n14221), .ZN(n11339) );
  OAI211_X1 U13838 ( .C1(n11698), .C2(n14372), .A(n11339), .B(n12084), .ZN(
        P1_U3332) );
  INV_X1 U13839 ( .A(n14085), .ZN(n13690) );
  NAND2_X1 U13840 ( .A1(n11342), .A2(n12022), .ZN(n11344) );
  AOI22_X1 U13841 ( .A1(n11627), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n11626), 
        .B2(n14649), .ZN(n11343) );
  XNOR2_X1 U13842 ( .A(n13843), .B(n14064), .ZN(n12051) );
  XNOR2_X1 U13843 ( .A(n13842), .B(n11352), .ZN(n14189) );
  INV_X1 U13844 ( .A(n14189), .ZN(n11368) );
  INV_X1 U13845 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11345) );
  OAI22_X1 U13846 ( .A1(n14691), .A2(n11345), .B1(n13614), .B2(n14751), .ZN(
        n11350) );
  NAND2_X1 U13847 ( .A1(n11346), .A2(n13843), .ZN(n11347) );
  NAND2_X1 U13848 ( .A1(n11347), .A2(n14756), .ZN(n11348) );
  OR2_X1 U13849 ( .A1(n14067), .A2(n11348), .ZN(n14186) );
  NOR2_X1 U13850 ( .A1(n14186), .A2(n14695), .ZN(n11349) );
  AOI211_X1 U13851 ( .C1(n14754), .C2(n13843), .A(n11350), .B(n11349), .ZN(
        n11367) );
  NAND2_X1 U13852 ( .A1(n11353), .A2(n11352), .ZN(n11354) );
  AOI21_X1 U13853 ( .B1(n13815), .B2(n11354), .A(n14744), .ZN(n14188) );
  INV_X1 U13854 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n11355) );
  AND2_X1 U13855 ( .A1(n11356), .A2(n11355), .ZN(n11357) );
  NOR2_X1 U13856 ( .A1(n11614), .A2(n11357), .ZN(n14069) );
  NAND2_X1 U13857 ( .A1(n14069), .A2(n9250), .ZN(n11362) );
  INV_X1 U13858 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n13788) );
  OR2_X1 U13859 ( .A1(n11818), .A2(n13788), .ZN(n11361) );
  NAND2_X1 U13860 ( .A1(n11846), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n11360) );
  INV_X1 U13861 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n11358) );
  OR2_X1 U13862 ( .A1(n11839), .A2(n11358), .ZN(n11359) );
  OR2_X1 U13863 ( .A1(n14052), .A2(n14720), .ZN(n11364) );
  OR2_X1 U13864 ( .A1(n14085), .A2(n14722), .ZN(n11363) );
  AND2_X1 U13865 ( .A1(n11364), .A2(n11363), .ZN(n14185) );
  INV_X1 U13866 ( .A(n14185), .ZN(n11365) );
  OAI21_X1 U13867 ( .B1(n14188), .B2(n11365), .A(n14691), .ZN(n11366) );
  OAI211_X1 U13868 ( .C1(n11368), .C2(n14059), .A(n11367), .B(n11366), .ZN(
        P1_U3277) );
  INV_X1 U13869 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n11371) );
  AOI21_X1 U13870 ( .B1(n15150), .B2(n11370), .A(n11369), .ZN(n11373) );
  MUX2_X1 U13871 ( .A(n11371), .B(n11373), .S(n15158), .Z(n11372) );
  OAI21_X1 U13872 ( .B1(n12926), .B2(n11437), .A(n11372), .ZN(P3_U3423) );
  MUX2_X1 U13873 ( .A(n8881), .B(n11373), .S(n15166), .Z(n11374) );
  OAI21_X1 U13874 ( .B1(n12876), .B2(n11437), .A(n11374), .ZN(P3_U3470) );
  XOR2_X1 U13875 ( .A(n12372), .B(n11375), .Z(n14484) );
  INV_X1 U13876 ( .A(n12547), .ZN(n11464) );
  XNOR2_X1 U13877 ( .A(n11376), .B(n12372), .ZN(n11377) );
  OAI222_X1 U13878 ( .A1(n12799), .A2(n11423), .B1(n15122), .B2(n11464), .C1(
        n11377), .C2(n15128), .ZN(n14486) );
  NAND2_X1 U13879 ( .A1(n14486), .A2(n12818), .ZN(n11381) );
  INV_X1 U13880 ( .A(n14482), .ZN(n11379) );
  OAI22_X1 U13881 ( .A1(n12818), .A2(n12626), .B1(n11421), .B2(n12816), .ZN(
        n11378) );
  AOI21_X1 U13882 ( .B1(n11379), .B2(n14471), .A(n11378), .ZN(n11380) );
  OAI211_X1 U13883 ( .C1(n12666), .C2(n14484), .A(n11381), .B(n11380), .ZN(
        P3_U3220) );
  NAND2_X1 U13884 ( .A1(n13504), .A2(n13081), .ZN(n11382) );
  XNOR2_X1 U13885 ( .A(n11543), .B(n11389), .ZN(n13501) );
  INV_X1 U13886 ( .A(n13410), .ZN(n11383) );
  AOI211_X1 U13887 ( .C1(n13498), .C2(n11384), .A(n13409), .B(n11383), .ZN(
        n13497) );
  AOI22_X1 U13888 ( .A1(n13426), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13001), 
        .B2(n13412), .ZN(n11385) );
  OAI21_X1 U13889 ( .B1(n7133), .B2(n13415), .A(n11385), .ZN(n11394) );
  OR2_X1 U13890 ( .A1(n13504), .A2(n11391), .ZN(n11386) );
  NAND2_X1 U13891 ( .A1(n13504), .A2(n11391), .ZN(n11388) );
  AOI21_X1 U13892 ( .B1(n11390), .B2(n11389), .A(n13294), .ZN(n11392) );
  OAI22_X1 U13893 ( .A1(n11525), .A2(n13052), .B1(n11391), .B2(n13051), .ZN(
        n13002) );
  AOI21_X1 U13894 ( .B1(n11392), .B2(n11524), .A(n13002), .ZN(n13500) );
  NOR2_X1 U13895 ( .A1(n13500), .A2(n13426), .ZN(n11393) );
  AOI211_X1 U13896 ( .C1(n13497), .C2(n13424), .A(n11394), .B(n11393), .ZN(
        n11395) );
  OAI21_X1 U13897 ( .B1(n13421), .B2(n13501), .A(n11395), .ZN(P2_U3248) );
  AND2_X1 U13898 ( .A1(n13692), .A2(n11808), .ZN(n11399) );
  AOI21_X1 U13899 ( .B1(n11939), .B2(n11775), .A(n11399), .ZN(n11448) );
  AOI22_X1 U13900 ( .A1(n11939), .A2(n11807), .B1(n11775), .B2(n13692), .ZN(
        n11400) );
  XNOR2_X1 U13901 ( .A(n11400), .B(n10326), .ZN(n11447) );
  XOR2_X1 U13902 ( .A(n11448), .B(n11447), .Z(n11401) );
  OAI211_X1 U13903 ( .C1(n11402), .C2(n11401), .A(n11452), .B(n13645), .ZN(
        n11408) );
  AND2_X1 U13904 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n13760) );
  AOI21_X1 U13905 ( .B1(n13664), .B2(n11403), .A(n13760), .ZN(n11404) );
  OAI21_X1 U13906 ( .B1(n13667), .B2(n11405), .A(n11404), .ZN(n11406) );
  AOI21_X1 U13907 ( .B1(n6433), .B2(n14086), .A(n11406), .ZN(n11407) );
  OAI211_X1 U13908 ( .C1(n11409), .C2(n13652), .A(n11408), .B(n11407), .ZN(
        P1_U3224) );
  INV_X1 U13909 ( .A(n11410), .ZN(n11411) );
  NAND2_X1 U13910 ( .A1(n11411), .A2(n12550), .ZN(n11412) );
  XNOR2_X1 U13911 ( .A(n12246), .B(n12153), .ZN(n11428) );
  XNOR2_X1 U13912 ( .A(n14487), .B(n12180), .ZN(n11482) );
  NOR2_X1 U13913 ( .A1(n11482), .A2(n11423), .ZN(n11416) );
  AOI21_X1 U13914 ( .B1(n12549), .B2(n11428), .A(n11416), .ZN(n11418) );
  INV_X1 U13915 ( .A(n11428), .ZN(n11480) );
  NAND2_X1 U13916 ( .A1(n11480), .A2(n7425), .ZN(n11415) );
  INV_X1 U13917 ( .A(n11482), .ZN(n11414) );
  OAI22_X1 U13918 ( .A1(n11416), .A2(n11415), .B1(n11414), .B2(n12548), .ZN(
        n11417) );
  XNOR2_X1 U13919 ( .A(n14482), .B(n12180), .ZN(n11471) );
  XNOR2_X1 U13920 ( .A(n11471), .B(n11441), .ZN(n11419) );
  OAI211_X1 U13921 ( .C1(n11420), .C2(n11419), .A(n6721), .B(n12499), .ZN(
        n11427) );
  INV_X1 U13922 ( .A(n11421), .ZN(n11425) );
  AND2_X1 U13923 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n15081) );
  AOI21_X1 U13924 ( .B1(n12503), .B2(n12547), .A(n15081), .ZN(n11422) );
  OAI21_X1 U13925 ( .B1(n11423), .B2(n12505), .A(n11422), .ZN(n11424) );
  AOI21_X1 U13926 ( .B1(n11425), .B2(n12531), .A(n11424), .ZN(n11426) );
  OAI211_X1 U13927 ( .C1(n12528), .C2(n14482), .A(n11427), .B(n11426), .ZN(
        P3_U3174) );
  XNOR2_X1 U13928 ( .A(n11481), .B(n11428), .ZN(n11429) );
  NAND2_X1 U13929 ( .A1(n11429), .A2(n12549), .ZN(n11479) );
  OAI211_X1 U13930 ( .C1(n11429), .C2(n12549), .A(n11479), .B(n12499), .ZN(
        n11436) );
  NOR2_X1 U13931 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11430), .ZN(n15047) );
  AOI21_X1 U13932 ( .B1(n12548), .B2(n12503), .A(n15047), .ZN(n11432) );
  NAND2_X1 U13933 ( .A1(n12550), .A2(n12525), .ZN(n11431) );
  OAI211_X1 U13934 ( .C1(n12461), .C2(n11433), .A(n11432), .B(n11431), .ZN(
        n11434) );
  INV_X1 U13935 ( .A(n11434), .ZN(n11435) );
  OAI211_X1 U13936 ( .C1(n12528), .C2(n11437), .A(n11436), .B(n11435), .ZN(
        P3_U3176) );
  INV_X1 U13937 ( .A(n12376), .ZN(n12258) );
  XNOR2_X1 U13938 ( .A(n11438), .B(n12258), .ZN(n14478) );
  XNOR2_X1 U13939 ( .A(n11439), .B(n12376), .ZN(n11440) );
  OAI222_X1 U13940 ( .A1(n15122), .A2(n12811), .B1(n12799), .B2(n11441), .C1(
        n11440), .C2(n15128), .ZN(n14480) );
  NAND2_X1 U13941 ( .A1(n14480), .A2(n12818), .ZN(n11446) );
  INV_X1 U13942 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n11442) );
  OAI22_X1 U13943 ( .A1(n12818), .A2(n11442), .B1(n11474), .B2(n12816), .ZN(
        n11443) );
  AOI21_X1 U13944 ( .B1(n11444), .B2(n14471), .A(n11443), .ZN(n11445) );
  OAI211_X1 U13945 ( .C1(n14478), .C2(n12666), .A(n11446), .B(n11445), .ZN(
        P3_U3219) );
  INV_X1 U13946 ( .A(n11448), .ZN(n11449) );
  NAND2_X1 U13947 ( .A1(n11450), .A2(n11449), .ZN(n11451) );
  NAND2_X1 U13948 ( .A1(n11452), .A2(n11451), .ZN(n11456) );
  AND2_X1 U13949 ( .A1(n14086), .A2(n11808), .ZN(n11453) );
  AOI21_X1 U13950 ( .B1(n11946), .B2(n11775), .A(n11453), .ZN(n11579) );
  AOI22_X1 U13951 ( .A1(n11946), .A2(n11807), .B1(n11775), .B2(n14086), .ZN(
        n11454) );
  XNOR2_X1 U13952 ( .A(n11454), .B(n10326), .ZN(n11578) );
  XOR2_X1 U13953 ( .A(n11579), .B(n11578), .Z(n11455) );
  OAI211_X1 U13954 ( .C1(n11456), .C2(n11455), .A(n11583), .B(n13645), .ZN(
        n11461) );
  NAND2_X1 U13955 ( .A1(n13681), .A2(n13692), .ZN(n11457) );
  NAND2_X1 U13956 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14611)
         );
  OAI211_X1 U13957 ( .C1(n13679), .C2(n11458), .A(n11457), .B(n14611), .ZN(
        n11459) );
  AOI21_X1 U13958 ( .B1(n6433), .B2(n13691), .A(n11459), .ZN(n11460) );
  OAI211_X1 U13959 ( .C1(n14544), .C2(n13652), .A(n11461), .B(n11460), .ZN(
        P1_U3234) );
  XNOR2_X1 U13960 ( .A(n11462), .B(n12373), .ZN(n11463) );
  OAI222_X1 U13961 ( .A1(n15122), .A2(n12798), .B1(n12799), .B2(n11464), .C1(
        n11463), .C2(n15128), .ZN(n12873) );
  INV_X1 U13962 ( .A(n12873), .ZN(n11470) );
  XNOR2_X1 U13963 ( .A(n11465), .B(n12373), .ZN(n12874) );
  INV_X1 U13964 ( .A(n11466), .ZN(n12532) );
  AOI22_X1 U13965 ( .A1(n15136), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15134), 
        .B2(n12532), .ZN(n11467) );
  OAI21_X1 U13966 ( .B1(n12925), .B2(n12815), .A(n11467), .ZN(n11468) );
  AOI21_X1 U13967 ( .B1(n12874), .B2(n12821), .A(n11468), .ZN(n11469) );
  OAI21_X1 U13968 ( .B1(n11470), .B2(n15136), .A(n11469), .ZN(P3_U3218) );
  NAND2_X1 U13969 ( .A1(n11471), .A2(n11485), .ZN(n11472) );
  XNOR2_X1 U13970 ( .A(n14477), .B(n12180), .ZN(n12132) );
  XOR2_X1 U13971 ( .A(n12547), .B(n12132), .Z(n12129) );
  NAND2_X1 U13972 ( .A1(n12131), .A2(n12129), .ZN(n12522) );
  OAI211_X1 U13973 ( .C1(n12131), .C2(n12129), .A(n12522), .B(n12499), .ZN(
        n11478) );
  NAND2_X1 U13974 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n15102)
         );
  OAI21_X1 U13975 ( .B1(n12811), .B2(n12527), .A(n15102), .ZN(n11476) );
  NOR2_X1 U13976 ( .A1(n12461), .A2(n11474), .ZN(n11475) );
  AOI211_X1 U13977 ( .C1(n12525), .C2(n11485), .A(n11476), .B(n11475), .ZN(
        n11477) );
  OAI211_X1 U13978 ( .C1(n12528), .C2(n14477), .A(n11478), .B(n11477), .ZN(
        P3_U3155) );
  OAI21_X1 U13979 ( .B1(n11481), .B2(n11480), .A(n11479), .ZN(n11484) );
  XNOR2_X1 U13980 ( .A(n11482), .B(n12548), .ZN(n11483) );
  XNOR2_X1 U13981 ( .A(n11484), .B(n11483), .ZN(n11491) );
  NOR2_X1 U13982 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14291), .ZN(n15066) );
  AOI21_X1 U13983 ( .B1(n12503), .B2(n11485), .A(n15066), .ZN(n11487) );
  NAND2_X1 U13984 ( .A1(n12525), .A2(n12549), .ZN(n11486) );
  OAI211_X1 U13985 ( .C1(n12461), .C2(n11488), .A(n11487), .B(n11486), .ZN(
        n11489) );
  AOI21_X1 U13986 ( .B1(n12515), .B2(n14487), .A(n11489), .ZN(n11490) );
  OAI21_X1 U13987 ( .B1(n11491), .B2(n12534), .A(n11490), .ZN(P3_U3164) );
  INV_X1 U13988 ( .A(n11793), .ZN(n11502) );
  OAI222_X1 U13989 ( .A1(n11492), .A2(P1_U3086), .B1(n14375), .B2(n11502), 
        .C1(n14257), .C2(n14372), .ZN(P1_U3327) );
  NAND2_X1 U13990 ( .A1(n13545), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n11493) );
  NAND2_X1 U13991 ( .A1(n11494), .A2(n11493), .ZN(n11496) );
  NAND2_X1 U13992 ( .A1(n14369), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n11495) );
  NAND2_X1 U13993 ( .A1(n11496), .A2(n11495), .ZN(n12340) );
  INV_X1 U13994 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14366) );
  AOI22_X1 U13995 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n12338), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n14366), .ZN(n11497) );
  INV_X1 U13996 ( .A(n11497), .ZN(n11498) );
  XNOR2_X1 U13997 ( .A(n12340), .B(n11498), .ZN(n12331) );
  INV_X1 U13998 ( .A(n12331), .ZN(n11499) );
  OAI222_X1 U13999 ( .A1(n13551), .A2(n11503), .B1(n13549), .B2(n11502), .C1(
        n8192), .C2(P2_U3088), .ZN(P2_U3299) );
  OAI21_X1 U14000 ( .B1(n11505), .B2(n9119), .A(n11504), .ZN(n11506) );
  NAND2_X1 U14001 ( .A1(n11507), .A2(n9119), .ZN(n11508) );
  OAI22_X1 U14002 ( .A1(n11510), .A2(n15122), .B1(n12453), .B2(n12799), .ZN(
        n11511) );
  INV_X1 U14003 ( .A(n11511), .ZN(n11512) );
  INV_X1 U14004 ( .A(n11517), .ZN(n12173) );
  OAI22_X1 U14005 ( .A1(n12173), .A2(n12816), .B1(n12818), .B2(n11518), .ZN(
        n11521) );
  NOR2_X1 U14006 ( .A1(n12086), .A2(n11519), .ZN(n11520) );
  AOI211_X1 U14007 ( .C1(n14471), .C2(n12170), .A(n11521), .B(n11520), .ZN(
        n11522) );
  OAI21_X1 U14008 ( .B1(n12087), .B2(n15136), .A(n11522), .ZN(P3_U3206) );
  INV_X1 U14009 ( .A(n13438), .ZN(n11536) );
  NAND2_X1 U14010 ( .A1(n13493), .A2(n11525), .ZN(n11527) );
  NOR2_X1 U14011 ( .A1(n13493), .A2(n11525), .ZN(n11526) );
  OR2_X1 U14012 ( .A1(n13488), .A2(n13053), .ZN(n11528) );
  INV_X1 U14013 ( .A(n13358), .ZN(n12989) );
  NOR2_X1 U14014 ( .A1(n13481), .A2(n12989), .ZN(n11529) );
  NAND2_X1 U14015 ( .A1(n13477), .A2(n13045), .ZN(n11530) );
  INV_X1 U14016 ( .A(n11531), .ZN(n11533) );
  INV_X1 U14017 ( .A(n13291), .ZN(n13289) );
  INV_X1 U14018 ( .A(n13456), .ZN(n13300) );
  INV_X1 U14019 ( .A(n13276), .ZN(n11535) );
  AOI21_X1 U14020 ( .B1(n11536), .B2(n13074), .A(n13243), .ZN(n11537) );
  AOI21_X1 U14021 ( .B1(n11538), .B2(P2_B_REG_SCAN_IN), .A(n13052), .ZN(n13232) );
  NAND2_X1 U14022 ( .A1(n13232), .A2(n13072), .ZN(n11539) );
  INV_X1 U14023 ( .A(n13355), .ZN(n11549) );
  OR2_X1 U14024 ( .A1(n13498), .A2(n13080), .ZN(n11542) );
  INV_X1 U14025 ( .A(n13403), .ZN(n13420) );
  OR2_X1 U14026 ( .A1(n13493), .A2(n13079), .ZN(n11544) );
  NAND2_X1 U14027 ( .A1(n13417), .A2(n11544), .ZN(n13390) );
  NAND2_X1 U14028 ( .A1(n13488), .A2(n13371), .ZN(n11545) );
  OR2_X1 U14029 ( .A1(n13488), .A2(n13371), .ZN(n11546) );
  NAND2_X1 U14030 ( .A1(n13481), .A2(n13358), .ZN(n11547) );
  AND2_X1 U14031 ( .A1(n13465), .A2(n13338), .ZN(n11550) );
  OR2_X1 U14032 ( .A1(n13465), .A2(n13338), .ZN(n11551) );
  NAND2_X1 U14033 ( .A1(n13462), .A2(n13078), .ZN(n11554) );
  OR2_X1 U14034 ( .A1(n13456), .A2(n13077), .ZN(n11555) );
  NAND2_X1 U14035 ( .A1(n13456), .A2(n13077), .ZN(n11556) );
  NOR2_X1 U14036 ( .A1(n13282), .A2(n11558), .ZN(n11557) );
  NAND2_X1 U14037 ( .A1(n13282), .A2(n11558), .ZN(n11559) );
  NAND2_X1 U14038 ( .A1(n13250), .A2(n13249), .ZN(n13248) );
  NAND2_X1 U14039 ( .A1(n11565), .A2(n13412), .ZN(n11566) );
  OAI21_X1 U14040 ( .B1(n13394), .B2(n11567), .A(n11566), .ZN(n11568) );
  AOI21_X1 U14041 ( .B1(n13434), .B2(n13381), .A(n11568), .ZN(n11573) );
  INV_X1 U14042 ( .A(n13481), .ZN(n13382) );
  NAND2_X1 U14043 ( .A1(n13382), .A2(n13396), .ZN(n13384) );
  OR2_X2 U14044 ( .A1(n13384), .A2(n13477), .ZN(n13363) );
  OR2_X2 U14045 ( .A1(n13472), .A2(n13363), .ZN(n13340) );
  NAND2_X1 U14046 ( .A1(n13280), .A2(n13265), .ZN(n13264) );
  INV_X1 U14048 ( .A(n13254), .ZN(n11570) );
  INV_X1 U14049 ( .A(n13434), .ZN(n11569) );
  AOI21_X1 U14050 ( .B1(n13254), .B2(n13434), .A(n13409), .ZN(n11571) );
  NAND2_X1 U14051 ( .A1(n13433), .A2(n13424), .ZN(n11572) );
  OAI211_X1 U14052 ( .C1(n13436), .C2(n13421), .A(n11573), .B(n11572), .ZN(
        n11574) );
  INV_X1 U14053 ( .A(n11574), .ZN(n11575) );
  OAI21_X1 U14054 ( .B1(n13435), .B2(n13426), .A(n11575), .ZN(P2_U3236) );
  INV_X1 U14055 ( .A(n11850), .ZN(n14368) );
  OAI222_X1 U14056 ( .A1(n13549), .A2(n14368), .B1(P2_U3088), .B2(n11576), 
        .C1(n12338), .C2(n13551), .ZN(P2_U3297) );
  INV_X1 U14057 ( .A(n13843), .ZN(n13841) );
  INV_X1 U14058 ( .A(n14064), .ZN(n13840) );
  OAI22_X1 U14059 ( .A1(n13841), .A2(n10161), .B1(n13840), .B2(n10153), .ZN(
        n11598) );
  INV_X1 U14060 ( .A(n11598), .ZN(n11600) );
  AOI22_X1 U14061 ( .A1(n13843), .A2(n11807), .B1(n11775), .B2(n14064), .ZN(
        n11577) );
  XNOR2_X1 U14062 ( .A(n11577), .B(n10326), .ZN(n11599) );
  INV_X1 U14063 ( .A(n11578), .ZN(n11581) );
  NOR2_X1 U14064 ( .A1(n11585), .A2(n10153), .ZN(n11584) );
  AOI21_X1 U14065 ( .B1(n14194), .B2(n11775), .A(n11584), .ZN(n11595) );
  NAND2_X1 U14066 ( .A1(n14194), .A2(n11807), .ZN(n11587) );
  OR2_X1 U14067 ( .A1(n11585), .A2(n10161), .ZN(n11586) );
  NAND2_X1 U14068 ( .A1(n11587), .A2(n11586), .ZN(n11588) );
  XNOR2_X1 U14069 ( .A(n11588), .B(n10326), .ZN(n11594) );
  XOR2_X1 U14070 ( .A(n11595), .B(n11594), .Z(n13563) );
  NAND2_X1 U14071 ( .A1(n13686), .A2(n11807), .ZN(n11590) );
  OR2_X1 U14072 ( .A1(n14085), .A2(n10161), .ZN(n11589) );
  NAND2_X1 U14073 ( .A1(n11590), .A2(n11589), .ZN(n11591) );
  XNOR2_X1 U14074 ( .A(n11591), .B(n10326), .ZN(n13675) );
  NAND2_X1 U14075 ( .A1(n13686), .A2(n11775), .ZN(n11593) );
  OR2_X1 U14076 ( .A1(n14085), .A2(n10153), .ZN(n11592) );
  NAND2_X1 U14077 ( .A1(n11593), .A2(n11592), .ZN(n13674) );
  INV_X1 U14078 ( .A(n11594), .ZN(n11596) );
  NAND2_X1 U14079 ( .A1(n11596), .A2(n11595), .ZN(n13672) );
  OAI21_X1 U14080 ( .B1(n13675), .B2(n13674), .A(n13672), .ZN(n11597) );
  XOR2_X1 U14081 ( .A(n11598), .B(n11599), .Z(n13612) );
  NAND2_X1 U14082 ( .A1(n11601), .A2(n12022), .ZN(n11603) );
  INV_X1 U14083 ( .A(n13789), .ZN(n14661) );
  AOI22_X1 U14084 ( .A1(n11627), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n11626), 
        .B2(n14661), .ZN(n11602) );
  AOI22_X1 U14085 ( .A1(n14070), .A2(n11775), .B1(n11808), .B2(n13844), .ZN(
        n11607) );
  NAND2_X1 U14086 ( .A1(n14070), .A2(n11807), .ZN(n11605) );
  OR2_X1 U14087 ( .A1(n14052), .A2(n10161), .ZN(n11604) );
  NAND2_X1 U14088 ( .A1(n11605), .A2(n11604), .ZN(n11606) );
  XNOR2_X1 U14089 ( .A(n11606), .B(n10326), .ZN(n11609) );
  XOR2_X1 U14090 ( .A(n11607), .B(n11609), .Z(n13619) );
  INV_X1 U14091 ( .A(n11607), .ZN(n11608) );
  OR2_X1 U14092 ( .A1(n11611), .A2(n11610), .ZN(n11613) );
  INV_X1 U14093 ( .A(n13790), .ZN(n14675) );
  AOI22_X1 U14094 ( .A1(n11627), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n11626), 
        .B2(n14675), .ZN(n11612) );
  NAND2_X1 U14095 ( .A1(n14174), .A2(n11807), .ZN(n11620) );
  OR2_X1 U14096 ( .A1(n11614), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n11615) );
  NAND2_X1 U14097 ( .A1(n11631), .A2(n11615), .ZN(n14055) );
  INV_X1 U14098 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n11616) );
  OAI22_X1 U14099 ( .A1(n14055), .A2(n9605), .B1(n11816), .B2(n11616), .ZN(
        n11618) );
  INV_X1 U14100 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14671) );
  INV_X1 U14101 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14667) );
  OAI22_X1 U14102 ( .A1(n11839), .A2(n14671), .B1(n11818), .B2(n14667), .ZN(
        n11617) );
  NAND2_X1 U14103 ( .A1(n14065), .A2(n11775), .ZN(n11619) );
  NAND2_X1 U14104 ( .A1(n11620), .A2(n11619), .ZN(n11621) );
  XNOR2_X1 U14105 ( .A(n11621), .B(n10326), .ZN(n11622) );
  AOI22_X1 U14106 ( .A1(n14174), .A2(n11775), .B1(n11808), .B2(n14065), .ZN(
        n11623) );
  XNOR2_X1 U14107 ( .A(n11622), .B(n11623), .ZN(n13654) );
  INV_X1 U14108 ( .A(n11622), .ZN(n11624) );
  AOI22_X1 U14109 ( .A1(n11627), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n12058), 
        .B2(n11626), .ZN(n11628) );
  NAND2_X1 U14110 ( .A1(n14027), .A2(n11807), .ZN(n11640) );
  INV_X1 U14111 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n11630) );
  NAND2_X1 U14112 ( .A1(n11631), .A2(n11630), .ZN(n11632) );
  NAND2_X1 U14113 ( .A1(n11651), .A2(n11632), .ZN(n14032) );
  OR2_X1 U14114 ( .A1(n14032), .A2(n9605), .ZN(n11638) );
  INV_X1 U14115 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n11633) );
  OR2_X1 U14116 ( .A1(n11818), .A2(n11633), .ZN(n11635) );
  INV_X1 U14117 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14033) );
  OR2_X1 U14118 ( .A1(n11839), .A2(n14033), .ZN(n11634) );
  AND2_X1 U14119 ( .A1(n11635), .A2(n11634), .ZN(n11637) );
  NAND2_X1 U14120 ( .A1(n11846), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n11636) );
  INV_X1 U14121 ( .A(n14054), .ZN(n14016) );
  NAND2_X1 U14122 ( .A1(n14016), .A2(n11775), .ZN(n11639) );
  NAND2_X1 U14123 ( .A1(n11640), .A2(n11639), .ZN(n11641) );
  XNOR2_X1 U14124 ( .A(n11641), .B(n10326), .ZN(n11643) );
  NOR2_X1 U14125 ( .A1(n14054), .A2(n10153), .ZN(n11642) );
  AOI21_X1 U14126 ( .B1(n14027), .B2(n11775), .A(n11642), .ZN(n11644) );
  XNOR2_X1 U14127 ( .A(n11643), .B(n11644), .ZN(n13587) );
  INV_X1 U14128 ( .A(n11643), .ZN(n11645) );
  OR2_X1 U14129 ( .A1(n11645), .A2(n11644), .ZN(n11646) );
  NAND2_X1 U14130 ( .A1(n11647), .A2(n12022), .ZN(n11650) );
  OR2_X1 U14131 ( .A1(n12023), .A2(n11648), .ZN(n11649) );
  INV_X1 U14132 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13637) );
  AND2_X1 U14133 ( .A1(n11651), .A2(n13637), .ZN(n11652) );
  OR2_X1 U14134 ( .A1(n11663), .A2(n11652), .ZN(n14018) );
  AOI22_X1 U14135 ( .A1(n11814), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n11845), 
        .B2(P1_REG1_REG_20__SCAN_IN), .ZN(n11654) );
  NAND2_X1 U14136 ( .A1(n11846), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n11653) );
  OAI211_X1 U14137 ( .C1(n14018), .C2(n9605), .A(n11654), .B(n11653), .ZN(
        n13996) );
  INV_X1 U14138 ( .A(n13996), .ZN(n14040) );
  OAI22_X1 U14139 ( .A1(n14161), .A2(n10161), .B1(n14040), .B2(n10153), .ZN(
        n11657) );
  OAI22_X1 U14140 ( .A1(n14161), .A2(n9766), .B1(n14040), .B2(n10161), .ZN(
        n11655) );
  XNOR2_X1 U14141 ( .A(n11655), .B(n10326), .ZN(n11656) );
  XOR2_X1 U14142 ( .A(n11657), .B(n11656), .Z(n13635) );
  NAND2_X1 U14143 ( .A1(n11656), .A2(n11657), .ZN(n11658) );
  NAND2_X1 U14144 ( .A1(n11659), .A2(n12022), .ZN(n11662) );
  OR2_X1 U14145 ( .A1(n12023), .A2(n11660), .ZN(n11661) );
  OR2_X1 U14146 ( .A1(n11663), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11664) );
  NAND2_X1 U14147 ( .A1(n11664), .A2(n11682), .ZN(n14002) );
  OR2_X1 U14148 ( .A1(n14002), .A2(n9605), .ZN(n11670) );
  INV_X1 U14149 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n11667) );
  NAND2_X1 U14150 ( .A1(n11845), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n11666) );
  NAND2_X1 U14151 ( .A1(n11846), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n11665) );
  OAI211_X1 U14152 ( .C1(n11839), .C2(n11667), .A(n11666), .B(n11665), .ZN(
        n11668) );
  INV_X1 U14153 ( .A(n11668), .ZN(n11669) );
  AOI22_X1 U14154 ( .A1(n14154), .A2(n11775), .B1(n11808), .B2(n14017), .ZN(
        n11675) );
  NAND2_X1 U14155 ( .A1(n14154), .A2(n11807), .ZN(n11672) );
  NAND2_X1 U14156 ( .A1(n14017), .A2(n11775), .ZN(n11671) );
  NAND2_X1 U14157 ( .A1(n11672), .A2(n11671), .ZN(n11673) );
  XNOR2_X1 U14158 ( .A(n11673), .B(n10326), .ZN(n11674) );
  XOR2_X1 U14159 ( .A(n11675), .B(n11674), .Z(n13596) );
  INV_X1 U14160 ( .A(n11674), .ZN(n11676) );
  NAND2_X1 U14161 ( .A1(n11676), .A2(n11675), .ZN(n11677) );
  OR2_X2 U14162 ( .A1(n11678), .A2(n6449), .ZN(n11679) );
  NAND2_X1 U14163 ( .A1(n14149), .A2(n11807), .ZN(n11691) );
  NAND2_X1 U14164 ( .A1(n11814), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n11689) );
  INV_X1 U14165 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n11681) );
  OR2_X1 U14166 ( .A1(n11816), .A2(n11681), .ZN(n11688) );
  INV_X1 U14167 ( .A(n11682), .ZN(n11684) );
  INV_X1 U14168 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13647) );
  INV_X1 U14169 ( .A(n11702), .ZN(n11683) );
  OAI21_X1 U14170 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n11684), .A(n11683), 
        .ZN(n13984) );
  OR2_X1 U14171 ( .A1(n9605), .A2(n13984), .ZN(n11687) );
  INV_X1 U14172 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n11685) );
  OR2_X1 U14173 ( .A1(n11818), .A2(n11685), .ZN(n11686) );
  NAND4_X1 U14174 ( .A1(n11689), .A2(n11688), .A3(n11687), .A4(n11686), .ZN(
        n13995) );
  NAND2_X1 U14175 ( .A1(n13995), .A2(n11775), .ZN(n11690) );
  NAND2_X1 U14176 ( .A1(n11691), .A2(n11690), .ZN(n11692) );
  XNOR2_X1 U14177 ( .A(n11692), .B(n10326), .ZN(n11693) );
  AOI22_X1 U14178 ( .A1(n14149), .A2(n11775), .B1(n11808), .B2(n13995), .ZN(
        n11694) );
  XNOR2_X1 U14179 ( .A(n11693), .B(n11694), .ZN(n13644) );
  INV_X1 U14180 ( .A(n11693), .ZN(n11695) );
  NAND2_X1 U14181 ( .A1(n11695), .A2(n11694), .ZN(n11696) );
  NAND2_X1 U14182 ( .A1(n11697), .A2(n12022), .ZN(n11700) );
  OR2_X1 U14183 ( .A1(n12023), .A2(n11698), .ZN(n11699) );
  NAND2_X1 U14184 ( .A1(n14144), .A2(n11807), .ZN(n11709) );
  NAND2_X1 U14185 ( .A1(n11845), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n11707) );
  INV_X1 U14186 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n11701) );
  OR2_X1 U14187 ( .A1(n11839), .A2(n11701), .ZN(n11706) );
  NAND2_X1 U14188 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(n11702), .ZN(n11722) );
  OAI21_X1 U14189 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n11702), .A(n11722), 
        .ZN(n13571) );
  OR2_X1 U14190 ( .A1(n9605), .A2(n13571), .ZN(n11705) );
  INV_X1 U14191 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n11703) );
  OR2_X1 U14192 ( .A1(n11816), .A2(n11703), .ZN(n11704) );
  NAND4_X1 U14193 ( .A1(n11707), .A2(n11706), .A3(n11705), .A4(n11704), .ZN(
        n13980) );
  NAND2_X1 U14194 ( .A1(n13980), .A2(n11775), .ZN(n11708) );
  NAND2_X1 U14195 ( .A1(n11709), .A2(n11708), .ZN(n11710) );
  XNOR2_X1 U14196 ( .A(n11710), .B(n10326), .ZN(n11711) );
  AOI22_X1 U14197 ( .A1(n14144), .A2(n11775), .B1(n11808), .B2(n13980), .ZN(
        n11712) );
  XNOR2_X1 U14198 ( .A(n11711), .B(n11712), .ZN(n13570) );
  INV_X1 U14199 ( .A(n11711), .ZN(n11713) );
  NAND2_X1 U14200 ( .A1(n11713), .A2(n11712), .ZN(n11714) );
  NAND2_X1 U14201 ( .A1(n11715), .A2(n12022), .ZN(n11718) );
  OR2_X1 U14202 ( .A1(n12023), .A2(n11716), .ZN(n11717) );
  NAND2_X1 U14203 ( .A1(n14139), .A2(n11807), .ZN(n11730) );
  NAND2_X1 U14204 ( .A1(n11845), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n11728) );
  INV_X1 U14205 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n11719) );
  OR2_X1 U14206 ( .A1(n11839), .A2(n11719), .ZN(n11727) );
  INV_X1 U14207 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n11721) );
  NAND2_X1 U14208 ( .A1(n11722), .A2(n11721), .ZN(n11723) );
  NAND2_X1 U14209 ( .A1(n11744), .A2(n11723), .ZN(n13628) );
  INV_X1 U14210 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n11724) );
  OR2_X1 U14211 ( .A1(n11816), .A2(n11724), .ZN(n11725) );
  NAND4_X1 U14212 ( .A1(n11728), .A2(n11727), .A3(n11726), .A4(n11725), .ZN(
        n14132) );
  NAND2_X1 U14213 ( .A1(n14132), .A2(n11775), .ZN(n11729) );
  NAND2_X1 U14214 ( .A1(n11730), .A2(n11729), .ZN(n11731) );
  XNOR2_X1 U14215 ( .A(n11731), .B(n10326), .ZN(n11732) );
  AOI22_X1 U14216 ( .A1(n14139), .A2(n11775), .B1(n11808), .B2(n14132), .ZN(
        n11733) );
  XNOR2_X1 U14217 ( .A(n11732), .B(n11733), .ZN(n13627) );
  INV_X1 U14218 ( .A(n11732), .ZN(n11734) );
  NAND2_X1 U14219 ( .A1(n11734), .A2(n11733), .ZN(n11735) );
  NAND2_X1 U14220 ( .A1(n11736), .A2(n11735), .ZN(n13603) );
  NAND2_X1 U14221 ( .A1(n11737), .A2(n12022), .ZN(n11740) );
  OR2_X1 U14222 ( .A1(n12023), .A2(n11738), .ZN(n11739) );
  NAND2_X1 U14223 ( .A1(n14133), .A2(n11807), .ZN(n11752) );
  NAND2_X1 U14224 ( .A1(n11845), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n11750) );
  INV_X1 U14225 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n11741) );
  OR2_X1 U14226 ( .A1(n11839), .A2(n11741), .ZN(n11749) );
  INV_X1 U14227 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n11743) );
  NAND2_X1 U14228 ( .A1(n11744), .A2(n11743), .ZN(n11745) );
  NAND2_X1 U14229 ( .A1(n11765), .A2(n11745), .ZN(n13942) );
  OR2_X1 U14230 ( .A1(n9605), .A2(n13942), .ZN(n11748) );
  INV_X1 U14231 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n11746) );
  OR2_X1 U14232 ( .A1(n11816), .A2(n11746), .ZN(n11747) );
  NAND4_X2 U14233 ( .A1(n11750), .A2(n11749), .A3(n11748), .A4(n11747), .ZN(
        n13924) );
  NAND2_X1 U14234 ( .A1(n13924), .A2(n11775), .ZN(n11751) );
  NAND2_X1 U14235 ( .A1(n11752), .A2(n11751), .ZN(n11753) );
  XNOR2_X1 U14236 ( .A(n11753), .B(n10326), .ZN(n11754) );
  AOI22_X1 U14237 ( .A1(n14133), .A2(n11775), .B1(n11808), .B2(n13924), .ZN(
        n11755) );
  XNOR2_X1 U14238 ( .A(n11754), .B(n11755), .ZN(n13604) );
  NAND2_X1 U14239 ( .A1(n13603), .A2(n13604), .ZN(n11758) );
  INV_X1 U14240 ( .A(n11754), .ZN(n11756) );
  NAND2_X1 U14241 ( .A1(n11756), .A2(n11755), .ZN(n11757) );
  NAND2_X1 U14242 ( .A1(n11759), .A2(n12022), .ZN(n11762) );
  OR2_X1 U14243 ( .A1(n12023), .A2(n11760), .ZN(n11761) );
  NAND2_X1 U14244 ( .A1(n14126), .A2(n11807), .ZN(n11773) );
  NAND2_X1 U14245 ( .A1(n11845), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n11771) );
  INV_X1 U14246 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n13914) );
  OR2_X1 U14247 ( .A1(n11839), .A2(n13914), .ZN(n11770) );
  INV_X1 U14248 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n11764) );
  NAND2_X1 U14249 ( .A1(n11765), .A2(n11764), .ZN(n11766) );
  NAND2_X1 U14250 ( .A1(n11798), .A2(n11766), .ZN(n13913) );
  OR2_X1 U14251 ( .A1(n9605), .A2(n13913), .ZN(n11769) );
  INV_X1 U14252 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n11767) );
  OR2_X1 U14253 ( .A1(n11816), .A2(n11767), .ZN(n11768) );
  NAND2_X1 U14254 ( .A1(n13933), .A2(n11775), .ZN(n11772) );
  NAND2_X1 U14255 ( .A1(n11773), .A2(n11772), .ZN(n11774) );
  XNOR2_X1 U14256 ( .A(n11774), .B(n10326), .ZN(n11776) );
  AOI22_X1 U14257 ( .A1(n14126), .A2(n11775), .B1(n11808), .B2(n13933), .ZN(
        n11777) );
  XNOR2_X1 U14258 ( .A(n11776), .B(n11777), .ZN(n13661) );
  INV_X1 U14259 ( .A(n11776), .ZN(n11778) );
  NAND2_X1 U14260 ( .A1(n11778), .A2(n11777), .ZN(n11779) );
  NAND2_X1 U14261 ( .A1(n13547), .A2(n12022), .ZN(n11781) );
  OR2_X1 U14262 ( .A1(n12023), .A2(n14373), .ZN(n11780) );
  NAND2_X1 U14263 ( .A1(n14121), .A2(n11807), .ZN(n11788) );
  NAND2_X1 U14264 ( .A1(n11845), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n11786) );
  INV_X1 U14265 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n13907) );
  OR2_X1 U14266 ( .A1(n11839), .A2(n13907), .ZN(n11785) );
  INV_X1 U14267 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n13556) );
  XNOR2_X1 U14268 ( .A(n11798), .B(n13556), .ZN(n13906) );
  INV_X1 U14269 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n11782) );
  OR2_X1 U14270 ( .A1(n11816), .A2(n11782), .ZN(n11783) );
  NAND2_X1 U14271 ( .A1(n13925), .A2(n11775), .ZN(n11787) );
  NAND2_X1 U14272 ( .A1(n11788), .A2(n11787), .ZN(n11789) );
  XNOR2_X1 U14273 ( .A(n11789), .B(n10326), .ZN(n11790) );
  AOI22_X1 U14274 ( .A1(n14121), .A2(n11775), .B1(n11808), .B2(n13925), .ZN(
        n11791) );
  XNOR2_X1 U14275 ( .A(n11790), .B(n11791), .ZN(n13555) );
  INV_X1 U14276 ( .A(n11790), .ZN(n11792) );
  NAND2_X1 U14277 ( .A1(n11793), .A2(n12022), .ZN(n11795) );
  OR2_X1 U14278 ( .A1(n12023), .A2(n14257), .ZN(n11794) );
  NAND2_X1 U14279 ( .A1(n11845), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n11806) );
  INV_X1 U14280 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n11796) );
  OR2_X1 U14281 ( .A1(n11839), .A2(n11796), .ZN(n11805) );
  INV_X1 U14282 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n11797) );
  OAI21_X1 U14283 ( .B1(n11798), .B2(n13556), .A(n11797), .ZN(n11801) );
  INV_X1 U14284 ( .A(n11798), .ZN(n11800) );
  AND2_X1 U14285 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n11799) );
  NAND2_X1 U14286 ( .A1(n11800), .A2(n11799), .ZN(n13865) );
  NAND2_X1 U14287 ( .A1(n11801), .A2(n13865), .ZN(n13884) );
  OR2_X1 U14288 ( .A1(n9605), .A2(n13884), .ZN(n11804) );
  INV_X1 U14289 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n11802) );
  OR2_X1 U14290 ( .A1(n11816), .A2(n11802), .ZN(n11803) );
  NAND4_X1 U14291 ( .A1(n11806), .A2(n11805), .A3(n11804), .A4(n11803), .ZN(
        n14105) );
  AOI22_X1 U14292 ( .A1(n14115), .A2(n11807), .B1(n11775), .B2(n14105), .ZN(
        n11811) );
  AOI22_X1 U14293 ( .A1(n14115), .A2(n11775), .B1(n11808), .B2(n14105), .ZN(
        n11809) );
  XNOR2_X1 U14294 ( .A(n11809), .B(n10326), .ZN(n11810) );
  XOR2_X1 U14295 ( .A(n11811), .B(n11810), .Z(n11812) );
  XNOR2_X1 U14296 ( .A(n11813), .B(n11812), .ZN(n11828) );
  NAND2_X1 U14297 ( .A1(n11814), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n11822) );
  INV_X1 U14298 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n11815) );
  OR2_X1 U14299 ( .A1(n11816), .A2(n11815), .ZN(n11821) );
  OR2_X1 U14300 ( .A1(n9605), .A2(n13865), .ZN(n11820) );
  INV_X1 U14301 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n11817) );
  OR2_X1 U14302 ( .A1(n11818), .A2(n11817), .ZN(n11819) );
  NAND4_X1 U14303 ( .A1(n11822), .A2(n11821), .A3(n11820), .A4(n11819), .ZN(
        n13879) );
  NAND2_X1 U14304 ( .A1(n6433), .A2(n13879), .ZN(n11825) );
  INV_X1 U14305 ( .A(n13884), .ZN(n11823) );
  AOI22_X1 U14306 ( .A1(n13664), .A2(n11823), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11824) );
  OAI211_X1 U14307 ( .C1(n13832), .C2(n13667), .A(n11825), .B(n11824), .ZN(
        n11826) );
  AOI21_X1 U14308 ( .B1(n14115), .B2(n13685), .A(n11826), .ZN(n11827) );
  OAI21_X1 U14309 ( .B1(n11828), .B2(n13688), .A(n11827), .ZN(P1_U3220) );
  OAI222_X1 U14310 ( .A1(n11500), .A2(n11831), .B1(n12933), .B2(n11830), .C1(
        P3_U3151), .C2(n11829), .ZN(P3_U3270) );
  AOI21_X1 U14311 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n15134), .A(n11832), .ZN(
        n11834) );
  MUX2_X1 U14312 ( .A(n11834), .B(n11833), .S(n15136), .Z(n11835) );
  OAI21_X1 U14313 ( .B1(n11836), .B2(n12815), .A(n11835), .ZN(P3_U3233) );
  INV_X1 U14314 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n13801) );
  NAND2_X1 U14315 ( .A1(n11845), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n11838) );
  NAND2_X1 U14316 ( .A1(n11846), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n11837) );
  OAI211_X1 U14317 ( .C1(n11839), .C2(n13801), .A(n11838), .B(n11837), .ZN(
        n13804) );
  OR2_X1 U14318 ( .A1(n11840), .A2(n12058), .ZN(n11841) );
  NAND2_X1 U14319 ( .A1(n11842), .A2(n11841), .ZN(n11854) );
  OR2_X1 U14320 ( .A1(n11854), .A2(n11843), .ZN(n11858) );
  INV_X1 U14321 ( .A(n11856), .ZN(n11849) );
  INV_X1 U14322 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n13809) );
  NAND2_X1 U14323 ( .A1(n11845), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n11848) );
  NAND2_X1 U14324 ( .A1(n11846), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n11847) );
  OAI211_X1 U14325 ( .C1(n11839), .C2(n13809), .A(n11848), .B(n11847), .ZN(
        n13868) );
  OAI21_X1 U14326 ( .B1(n13804), .B2(n11849), .A(n13868), .ZN(n11857) );
  NAND2_X1 U14327 ( .A1(n11850), .A2(n12022), .ZN(n11852) );
  OR2_X1 U14328 ( .A1(n12023), .A2(n14366), .ZN(n11851) );
  OR2_X1 U14329 ( .A1(n11854), .A2(n11853), .ZN(n11855) );
  AND2_X4 U14330 ( .A1(n11856), .A2(n11855), .ZN(n12026) );
  MUX2_X1 U14331 ( .A(n11857), .B(n14103), .S(n12026), .Z(n12071) );
  INV_X1 U14332 ( .A(n12071), .ZN(n11864) );
  NAND2_X1 U14333 ( .A1(n13812), .A2(n11873), .ZN(n11862) );
  NAND2_X1 U14334 ( .A1(n13804), .A2(n12026), .ZN(n11859) );
  NAND2_X1 U14335 ( .A1(n11859), .A2(n11858), .ZN(n11860) );
  NAND2_X1 U14336 ( .A1(n11860), .A2(n13868), .ZN(n11861) );
  NAND2_X1 U14337 ( .A1(n11862), .A2(n11861), .ZN(n12070) );
  INV_X1 U14338 ( .A(n12070), .ZN(n11863) );
  NAND2_X1 U14339 ( .A1(n11864), .A2(n11863), .ZN(n12069) );
  INV_X1 U14340 ( .A(n12069), .ZN(n11871) );
  NAND2_X1 U14341 ( .A1(n14222), .A2(n12022), .ZN(n11866) );
  INV_X1 U14342 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14218) );
  OR2_X1 U14343 ( .A1(n12023), .A2(n14218), .ZN(n11865) );
  INV_X1 U14344 ( .A(n13804), .ZN(n12062) );
  XNOR2_X1 U14345 ( .A(n14098), .B(n12062), .ZN(n12061) );
  NAND2_X1 U14346 ( .A1(n11868), .A2(n11867), .ZN(n11869) );
  NAND2_X1 U14347 ( .A1(n11870), .A2(n11869), .ZN(n12060) );
  INV_X1 U14348 ( .A(n12060), .ZN(n12065) );
  NAND2_X1 U14349 ( .A1(n6906), .A2(n12065), .ZN(n12072) );
  AOI21_X1 U14350 ( .B1(n9671), .B2(n12026), .A(n11872), .ZN(n11886) );
  NAND2_X1 U14351 ( .A1(n13700), .A2(n12026), .ZN(n11877) );
  AOI21_X1 U14352 ( .B1(n11877), .B2(n13700), .A(n11876), .ZN(n11885) );
  INV_X1 U14353 ( .A(n13702), .ZN(n11874) );
  NAND3_X1 U14354 ( .A1(n11874), .A2(n9278), .A3(n6454), .ZN(n11883) );
  OAI21_X1 U14355 ( .B1(n13702), .B2(n6617), .A(n12026), .ZN(n11875) );
  OAI21_X1 U14356 ( .B1(n11877), .B2(n11876), .A(n11875), .ZN(n11878) );
  NAND2_X1 U14357 ( .A1(n12032), .A2(n9514), .ZN(n11880) );
  NAND2_X1 U14358 ( .A1(n11880), .A2(n11879), .ZN(n11881) );
  NOR2_X1 U14359 ( .A1(n11878), .A2(n11881), .ZN(n11882) );
  NAND2_X1 U14360 ( .A1(n11883), .A2(n11882), .ZN(n11884) );
  OAI211_X1 U14361 ( .C1(n11886), .C2(n11885), .A(n11884), .B(n12034), .ZN(
        n11889) );
  MUX2_X1 U14362 ( .A(n11887), .B(n14741), .S(n6454), .Z(n11888) );
  NAND2_X1 U14363 ( .A1(n11889), .A2(n11888), .ZN(n11890) );
  NAND2_X1 U14364 ( .A1(n11890), .A2(n12035), .ZN(n11894) );
  MUX2_X1 U14365 ( .A(n11892), .B(n11891), .S(n11873), .Z(n11893) );
  NAND2_X1 U14366 ( .A1(n11894), .A2(n11893), .ZN(n11898) );
  MUX2_X1 U14367 ( .A(n13697), .B(n11895), .S(n11873), .Z(n11897) );
  MUX2_X1 U14368 ( .A(n11895), .B(n13697), .S(n11873), .Z(n11896) );
  MUX2_X1 U14369 ( .A(n14734), .B(n13696), .S(n11873), .Z(n11901) );
  MUX2_X1 U14370 ( .A(n13696), .B(n14734), .S(n11873), .Z(n11899) );
  NAND2_X1 U14371 ( .A1(n11900), .A2(n11899), .ZN(n11904) );
  OR2_X1 U14372 ( .A1(n11902), .A2(n11901), .ZN(n11903) );
  NAND2_X1 U14373 ( .A1(n11904), .A2(n11903), .ZN(n11907) );
  MUX2_X1 U14374 ( .A(n14704), .B(n14793), .S(n6454), .Z(n11908) );
  NAND2_X1 U14375 ( .A1(n11907), .A2(n11908), .ZN(n11906) );
  MUX2_X1 U14376 ( .A(n14793), .B(n14704), .S(n11873), .Z(n11905) );
  NAND2_X1 U14377 ( .A1(n11906), .A2(n11905), .ZN(n11912) );
  INV_X1 U14378 ( .A(n11907), .ZN(n11910) );
  INV_X1 U14379 ( .A(n11908), .ZN(n11909) );
  NAND2_X1 U14380 ( .A1(n11910), .A2(n11909), .ZN(n11911) );
  MUX2_X1 U14381 ( .A(n14682), .B(n14712), .S(n6911), .Z(n11914) );
  MUX2_X1 U14382 ( .A(n14712), .B(n14682), .S(n6911), .Z(n11913) );
  MUX2_X1 U14383 ( .A(n14703), .B(n14693), .S(n6454), .Z(n11918) );
  NAND2_X1 U14384 ( .A1(n11917), .A2(n11918), .ZN(n11916) );
  MUX2_X1 U14385 ( .A(n14703), .B(n14693), .S(n6911), .Z(n11915) );
  NAND2_X1 U14386 ( .A1(n11916), .A2(n11915), .ZN(n11922) );
  INV_X1 U14387 ( .A(n11917), .ZN(n11920) );
  INV_X1 U14388 ( .A(n11918), .ZN(n11919) );
  NAND2_X1 U14389 ( .A1(n11920), .A2(n11919), .ZN(n11921) );
  NAND2_X1 U14390 ( .A1(n11922), .A2(n11921), .ZN(n11926) );
  MUX2_X1 U14391 ( .A(n14683), .B(n11923), .S(n6911), .Z(n11925) );
  MUX2_X1 U14392 ( .A(n14683), .B(n11923), .S(n11873), .Z(n11924) );
  MUX2_X1 U14393 ( .A(n13694), .B(n11927), .S(n11873), .Z(n11931) );
  MUX2_X1 U14394 ( .A(n13694), .B(n11927), .S(n6911), .Z(n11928) );
  NAND2_X1 U14395 ( .A1(n11929), .A2(n11928), .ZN(n11935) );
  INV_X1 U14396 ( .A(n11930), .ZN(n11933) );
  INV_X1 U14397 ( .A(n11931), .ZN(n11932) );
  NAND2_X1 U14398 ( .A1(n11933), .A2(n11932), .ZN(n11934) );
  MUX2_X1 U14399 ( .A(n13693), .B(n11936), .S(n6911), .Z(n11938) );
  MUX2_X1 U14400 ( .A(n13693), .B(n11936), .S(n6454), .Z(n11937) );
  MUX2_X1 U14401 ( .A(n13692), .B(n11939), .S(n11873), .Z(n11943) );
  NAND2_X1 U14402 ( .A1(n11942), .A2(n11943), .ZN(n11941) );
  MUX2_X1 U14403 ( .A(n13692), .B(n11939), .S(n6911), .Z(n11940) );
  INV_X1 U14404 ( .A(n11942), .ZN(n11945) );
  INV_X1 U14405 ( .A(n11943), .ZN(n11944) );
  MUX2_X1 U14406 ( .A(n14086), .B(n11946), .S(n6911), .Z(n11949) );
  MUX2_X1 U14407 ( .A(n11947), .B(n14544), .S(n11873), .Z(n11948) );
  NAND2_X1 U14408 ( .A1(n11955), .A2(n11950), .ZN(n11953) );
  NAND2_X1 U14409 ( .A1(n11954), .A2(n11951), .ZN(n11952) );
  MUX2_X1 U14410 ( .A(n11953), .B(n11952), .S(n11873), .Z(n11957) );
  MUX2_X1 U14411 ( .A(n11955), .B(n11954), .S(n6911), .Z(n11956) );
  OAI21_X1 U14412 ( .B1(n11958), .B2(n11957), .A(n11956), .ZN(n11962) );
  XNOR2_X1 U14413 ( .A(n14070), .B(n14052), .ZN(n12050) );
  MUX2_X1 U14414 ( .A(n13840), .B(n13841), .S(n6454), .Z(n11967) );
  OR2_X1 U14415 ( .A1(n14070), .A2(n14052), .ZN(n13817) );
  NAND2_X1 U14416 ( .A1(n14070), .A2(n14052), .ZN(n13816) );
  AND2_X1 U14417 ( .A1(n14064), .A2(n6454), .ZN(n11959) );
  AOI21_X1 U14418 ( .B1(n13843), .B2(n6911), .A(n11959), .ZN(n11960) );
  NAND3_X1 U14419 ( .A1(n13817), .A2(n13816), .A3(n11960), .ZN(n11966) );
  OAI21_X1 U14420 ( .B1(n12050), .B2(n11967), .A(n11966), .ZN(n11961) );
  NAND2_X1 U14421 ( .A1(n11962), .A2(n11961), .ZN(n11970) );
  NAND2_X1 U14422 ( .A1(n14174), .A2(n14065), .ZN(n13845) );
  NAND2_X1 U14423 ( .A1(n13846), .A2(n13845), .ZN(n14050) );
  AND2_X1 U14424 ( .A1(n13844), .A2(n6911), .ZN(n11964) );
  OAI21_X1 U14425 ( .B1(n6911), .B2(n13844), .A(n14070), .ZN(n11963) );
  OAI21_X1 U14426 ( .B1(n11964), .B2(n14070), .A(n11963), .ZN(n11965) );
  OAI211_X1 U14427 ( .C1(n11967), .C2(n11966), .A(n14050), .B(n11965), .ZN(
        n11968) );
  INV_X1 U14428 ( .A(n11968), .ZN(n11969) );
  NAND2_X1 U14429 ( .A1(n11970), .A2(n11969), .ZN(n11974) );
  NAND2_X1 U14430 ( .A1(n14065), .A2(n11873), .ZN(n11972) );
  INV_X1 U14431 ( .A(n14065), .ZN(n14166) );
  NAND2_X1 U14432 ( .A1(n14166), .A2(n6911), .ZN(n11971) );
  MUX2_X1 U14433 ( .A(n11972), .B(n11971), .S(n14174), .Z(n11973) );
  AOI21_X1 U14434 ( .B1(n11974), .B2(n11973), .A(n14039), .ZN(n11979) );
  INV_X1 U14435 ( .A(n13821), .ZN(n11977) );
  INV_X1 U14436 ( .A(n11975), .ZN(n11976) );
  MUX2_X1 U14437 ( .A(n11977), .B(n11976), .S(n6454), .Z(n11978) );
  OR2_X1 U14438 ( .A1(n11979), .A2(n11978), .ZN(n11982) );
  MUX2_X1 U14439 ( .A(n14040), .B(n14161), .S(n6454), .Z(n11981) );
  MUX2_X1 U14440 ( .A(n13996), .B(n14012), .S(n6911), .Z(n11980) );
  OAI21_X1 U14441 ( .B1(n11982), .B2(n11981), .A(n11980), .ZN(n11984) );
  NAND2_X1 U14442 ( .A1(n11982), .A2(n11981), .ZN(n11983) );
  MUX2_X1 U14443 ( .A(n14017), .B(n14154), .S(n6911), .Z(n11986) );
  MUX2_X1 U14444 ( .A(n14017), .B(n14154), .S(n11873), .Z(n11985) );
  INV_X1 U14445 ( .A(n11986), .ZN(n11987) );
  MUX2_X1 U14446 ( .A(n13995), .B(n14149), .S(n6454), .Z(n11990) );
  NAND2_X1 U14447 ( .A1(n11991), .A2(n11990), .ZN(n11989) );
  MUX2_X1 U14448 ( .A(n13995), .B(n14149), .S(n6911), .Z(n11988) );
  NAND2_X1 U14449 ( .A1(n11989), .A2(n11988), .ZN(n11993) );
  MUX2_X1 U14450 ( .A(n13980), .B(n14144), .S(n6911), .Z(n11995) );
  MUX2_X1 U14451 ( .A(n13980), .B(n14144), .S(n11873), .Z(n11994) );
  MUX2_X1 U14452 ( .A(n14132), .B(n14139), .S(n6454), .Z(n11997) );
  MUX2_X1 U14453 ( .A(n14132), .B(n14139), .S(n6911), .Z(n11996) );
  INV_X1 U14454 ( .A(n11997), .ZN(n11998) );
  MUX2_X1 U14455 ( .A(n13924), .B(n14133), .S(n12026), .Z(n12002) );
  NAND2_X1 U14456 ( .A1(n12001), .A2(n12002), .ZN(n12000) );
  MUX2_X1 U14457 ( .A(n13924), .B(n14133), .S(n6454), .Z(n11999) );
  NAND2_X1 U14458 ( .A1(n12000), .A2(n11999), .ZN(n12006) );
  INV_X1 U14459 ( .A(n12001), .ZN(n12004) );
  INV_X1 U14460 ( .A(n12002), .ZN(n12003) );
  NAND2_X1 U14461 ( .A1(n12004), .A2(n12003), .ZN(n12005) );
  MUX2_X1 U14462 ( .A(n13933), .B(n14126), .S(n11873), .Z(n12008) );
  MUX2_X1 U14463 ( .A(n13933), .B(n14126), .S(n6911), .Z(n12007) );
  INV_X1 U14464 ( .A(n12008), .ZN(n12009) );
  MUX2_X1 U14465 ( .A(n14121), .B(n13925), .S(n6454), .Z(n12012) );
  MUX2_X1 U14466 ( .A(n13925), .B(n14121), .S(n11873), .Z(n12010) );
  INV_X1 U14467 ( .A(n12012), .ZN(n12013) );
  MUX2_X1 U14468 ( .A(n14105), .B(n14115), .S(n6454), .Z(n12017) );
  MUX2_X1 U14469 ( .A(n14105), .B(n14115), .S(n12026), .Z(n12014) );
  NAND2_X1 U14470 ( .A1(n12015), .A2(n12014), .ZN(n12021) );
  INV_X1 U14471 ( .A(n12016), .ZN(n12019) );
  INV_X1 U14472 ( .A(n12017), .ZN(n12018) );
  NAND2_X1 U14473 ( .A1(n12019), .A2(n12018), .ZN(n12020) );
  NAND2_X1 U14474 ( .A1(n13544), .A2(n12022), .ZN(n12025) );
  OR2_X1 U14475 ( .A1(n12023), .A2(n14369), .ZN(n12024) );
  MUX2_X1 U14476 ( .A(n13879), .B(n14109), .S(n12026), .Z(n12028) );
  MUX2_X1 U14477 ( .A(n13879), .B(n14109), .S(n11873), .Z(n12027) );
  INV_X1 U14478 ( .A(n12028), .ZN(n12029) );
  INV_X1 U14479 ( .A(n12077), .ZN(n12079) );
  INV_X1 U14480 ( .A(n13879), .ZN(n12030) );
  XNOR2_X1 U14481 ( .A(n14109), .B(n12030), .ZN(n13837) );
  XNOR2_X1 U14482 ( .A(n14115), .B(n13899), .ZN(n13877) );
  NAND2_X1 U14483 ( .A1(n14126), .A2(n13900), .ZN(n13895) );
  OR2_X1 U14484 ( .A1(n14126), .A2(n13900), .ZN(n12031) );
  NAND2_X1 U14485 ( .A1(n13895), .A2(n12031), .ZN(n13858) );
  INV_X1 U14486 ( .A(n14017), .ZN(n13823) );
  XNOR2_X1 U14487 ( .A(n14154), .B(n13823), .ZN(n13992) );
  NAND4_X1 U14488 ( .A1(n12035), .A2(n12034), .A3(n12033), .A4(n12032), .ZN(
        n12037) );
  NOR3_X1 U14489 ( .A1(n12037), .A2(n12036), .A3(n14724), .ZN(n12040) );
  NAND4_X1 U14490 ( .A1(n14686), .A2(n12040), .A3(n12039), .A4(n12038), .ZN(
        n12041) );
  OR4_X1 U14491 ( .A1(n12044), .A2(n12043), .A3(n12042), .A4(n12041), .ZN(
        n12046) );
  OR4_X1 U14492 ( .A1(n14082), .A2(n12047), .A3(n12046), .A4(n12045), .ZN(
        n12048) );
  NOR2_X1 U14493 ( .A1(n12049), .A2(n12048), .ZN(n12052) );
  NAND4_X1 U14494 ( .A1(n14050), .A2(n12052), .A3(n12051), .A4(n14061), .ZN(
        n12053) );
  NOR2_X1 U14495 ( .A1(n14039), .A2(n12053), .ZN(n12054) );
  XNOR2_X1 U14496 ( .A(n14139), .B(n14132), .ZN(n13829) );
  NAND4_X1 U14497 ( .A1(n13938), .A2(n12054), .A3(n13829), .A4(n14010), .ZN(
        n12055) );
  INV_X1 U14498 ( .A(n13980), .ZN(n13961) );
  XNOR2_X1 U14499 ( .A(n14144), .B(n13961), .ZN(n13827) );
  OR4_X2 U14500 ( .A1(n13877), .A2(n12056), .A3(n13896), .A4(n13827), .ZN(
        n12057) );
  AND2_X1 U14501 ( .A1(n12060), .A2(n12059), .ZN(n12067) );
  AND2_X1 U14502 ( .A1(n12061), .A2(n12067), .ZN(n12066) );
  NAND2_X1 U14503 ( .A1(n14098), .A2(n12062), .ZN(n12064) );
  OR2_X1 U14504 ( .A1(n14098), .A2(n12062), .ZN(n12063) );
  NAND2_X1 U14505 ( .A1(n12068), .A2(n12067), .ZN(n12075) );
  AND2_X1 U14506 ( .A1(n12071), .A2(n12070), .ZN(n12074) );
  INV_X1 U14507 ( .A(n12074), .ZN(n12073) );
  OR2_X1 U14508 ( .A1(n12075), .A2(n12074), .ZN(n12076) );
  INV_X1 U14509 ( .A(n12080), .ZN(n12085) );
  NAND3_X1 U14510 ( .A1(n12081), .A2(n14582), .A3(n14705), .ZN(n12082) );
  OAI211_X1 U14511 ( .C1(n11840), .C2(n12084), .A(n12082), .B(P1_B_REG_SCAN_IN), .ZN(n12083) );
  OAI21_X1 U14512 ( .B1(n12085), .B2(n12084), .A(n12083), .ZN(P1_U3242) );
  INV_X1 U14513 ( .A(n12170), .ZN(n12830) );
  INV_X1 U14514 ( .A(n15143), .ZN(n15146) );
  INV_X1 U14515 ( .A(n12088), .ZN(n12089) );
  OAI21_X1 U14516 ( .B1(n12830), .B2(n12926), .A(n12089), .ZN(P3_U3454) );
  NAND2_X1 U14517 ( .A1(n13054), .A2(n12090), .ZN(n12092) );
  OAI211_X1 U14518 ( .C1(n14528), .C2(n12093), .A(n12092), .B(n12091), .ZN(
        n12099) );
  INV_X1 U14519 ( .A(n12128), .ZN(n12097) );
  AOI22_X1 U14520 ( .A1(n12094), .A2(n14523), .B1(n13040), .B2(n13086), .ZN(
        n12096) );
  NOR3_X1 U14521 ( .A1(n12097), .A2(n12096), .A3(n12095), .ZN(n12098) );
  AOI211_X1 U14522 ( .C1(n12100), .C2(n14507), .A(n12099), .B(n12098), .ZN(
        n12101) );
  OAI21_X1 U14523 ( .B1(n12102), .B2(n14502), .A(n12101), .ZN(P2_U3196) );
  INV_X1 U14524 ( .A(n13397), .ZN(n12106) );
  NAND2_X1 U14525 ( .A1(n13358), .A2(n13372), .ZN(n12104) );
  NAND2_X1 U14526 ( .A1(n13079), .A2(n13370), .ZN(n12103) );
  NAND2_X1 U14527 ( .A1(n12104), .A2(n12103), .ZN(n13487) );
  NAND2_X1 U14528 ( .A1(n13054), .A2(n13487), .ZN(n12105) );
  NAND2_X1 U14529 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13228)
         );
  OAI211_X1 U14530 ( .C1(n14528), .C2(n12106), .A(n12105), .B(n13228), .ZN(
        n12113) );
  INV_X1 U14531 ( .A(n12107), .ZN(n13056) );
  NAND2_X1 U14532 ( .A1(n13056), .A2(n14523), .ZN(n12111) );
  NAND3_X1 U14533 ( .A1(n12108), .A2(n13040), .A3(n13079), .ZN(n12110) );
  AOI21_X1 U14534 ( .B1(n12111), .B2(n12110), .A(n12109), .ZN(n12112) );
  AOI211_X1 U14535 ( .C1(n13488), .C2(n14507), .A(n12113), .B(n12112), .ZN(
        n12114) );
  OAI21_X1 U14536 ( .B1(n12115), .B2(n14502), .A(n12114), .ZN(P2_U3191) );
  AOI22_X1 U14537 ( .A1(n13054), .A2(n12116), .B1(P2_REG3_REG_11__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12117) );
  OAI21_X1 U14538 ( .B1(n12118), .B2(n14528), .A(n12117), .ZN(n12125) );
  INV_X1 U14539 ( .A(n12119), .ZN(n12961) );
  NAND2_X1 U14540 ( .A1(n12961), .A2(n14523), .ZN(n12123) );
  NAND3_X1 U14541 ( .A1(n12120), .A2(n13040), .A3(n13087), .ZN(n12122) );
  AOI21_X1 U14542 ( .B1(n12123), .B2(n12122), .A(n12121), .ZN(n12124) );
  AOI211_X1 U14543 ( .C1(n12126), .C2(n14507), .A(n12125), .B(n12124), .ZN(
        n12127) );
  OAI21_X1 U14544 ( .B1(n12128), .B2(n14502), .A(n12127), .ZN(P2_U3208) );
  XNOR2_X1 U14545 ( .A(n12439), .B(n12180), .ZN(n12147) );
  INV_X1 U14546 ( .A(n12147), .ZN(n12148) );
  INV_X1 U14547 ( .A(n12785), .ZN(n12542) );
  XNOR2_X1 U14548 ( .A(n12925), .B(n12153), .ZN(n12133) );
  NAND2_X1 U14549 ( .A1(n12133), .A2(n12811), .ZN(n12519) );
  AND2_X1 U14550 ( .A1(n12129), .A2(n12519), .ZN(n12130) );
  INV_X1 U14551 ( .A(n12519), .ZN(n12136) );
  NAND2_X1 U14552 ( .A1(n12132), .A2(n12547), .ZN(n12521) );
  INV_X1 U14553 ( .A(n12133), .ZN(n12134) );
  NAND2_X1 U14554 ( .A1(n12134), .A2(n12546), .ZN(n12520) );
  AND2_X1 U14555 ( .A1(n12521), .A2(n12520), .ZN(n12135) );
  OR2_X1 U14556 ( .A1(n12136), .A2(n12135), .ZN(n12137) );
  XNOR2_X1 U14557 ( .A(n12922), .B(n12180), .ZN(n12138) );
  XNOR2_X1 U14558 ( .A(n12138), .B(n12545), .ZN(n12458) );
  XNOR2_X1 U14559 ( .A(n12918), .B(n12180), .ZN(n12141) );
  XNOR2_X1 U14560 ( .A(n12141), .B(n12544), .ZN(n12466) );
  XNOR2_X1 U14561 ( .A(n12139), .B(n12180), .ZN(n12144) );
  XOR2_X1 U14562 ( .A(n12800), .B(n12144), .Z(n12501) );
  INV_X1 U14563 ( .A(n12501), .ZN(n12142) );
  OR2_X1 U14564 ( .A1(n12466), .A2(n12142), .ZN(n12140) );
  NAND2_X1 U14565 ( .A1(n12141), .A2(n12544), .ZN(n12497) );
  INV_X1 U14566 ( .A(n12144), .ZN(n12145) );
  INV_X1 U14567 ( .A(n12800), .ZN(n12543) );
  NAND2_X1 U14568 ( .A1(n12145), .A2(n12543), .ZN(n12146) );
  NAND2_X1 U14569 ( .A1(n12500), .A2(n12146), .ZN(n12434) );
  XNOR2_X1 U14570 ( .A(n12147), .B(n12785), .ZN(n12435) );
  OR2_X2 U14571 ( .A1(n12434), .A2(n12435), .ZN(n12432) );
  XNOR2_X1 U14572 ( .A(n12482), .B(n12180), .ZN(n12149) );
  XNOR2_X1 U14573 ( .A(n12149), .B(n12746), .ZN(n12483) );
  INV_X1 U14574 ( .A(n12149), .ZN(n12150) );
  NAND2_X1 U14575 ( .A1(n12150), .A2(n12770), .ZN(n12151) );
  XNOR2_X1 U14576 ( .A(n12750), .B(n12180), .ZN(n12152) );
  XNOR2_X1 U14577 ( .A(n12152), .B(n12758), .ZN(n12443) );
  XNOR2_X1 U14578 ( .A(n12736), .B(n12153), .ZN(n12154) );
  XNOR2_X1 U14579 ( .A(n12725), .B(n12180), .ZN(n12158) );
  XNOR2_X1 U14580 ( .A(n12160), .B(n12158), .ZN(n12426) );
  NAND2_X1 U14581 ( .A1(n12426), .A2(n12733), .ZN(n12162) );
  INV_X1 U14582 ( .A(n12158), .ZN(n12159) );
  OR2_X1 U14583 ( .A1(n12160), .A2(n12159), .ZN(n12161) );
  NAND2_X1 U14584 ( .A1(n12162), .A2(n12161), .ZN(n12475) );
  XNOR2_X1 U14585 ( .A(n12712), .B(n12180), .ZN(n12163) );
  XNOR2_X1 U14586 ( .A(n12163), .B(n12720), .ZN(n12476) );
  NAND2_X1 U14587 ( .A1(n12163), .A2(n12694), .ZN(n12164) );
  XNOR2_X1 U14588 ( .A(n12698), .B(n12180), .ZN(n12165) );
  XNOR2_X1 U14589 ( .A(n12165), .B(n12707), .ZN(n12450) );
  XNOR2_X1 U14590 ( .A(n12884), .B(n12180), .ZN(n12166) );
  XNOR2_X1 U14591 ( .A(n12166), .B(n12453), .ZN(n12511) );
  NAND2_X1 U14592 ( .A1(n12510), .A2(n12511), .ZN(n12169) );
  INV_X1 U14593 ( .A(n12166), .ZN(n12167) );
  NAND2_X1 U14594 ( .A1(n12167), .A2(n12453), .ZN(n12168) );
  XNOR2_X1 U14595 ( .A(n12170), .B(n12180), .ZN(n12177) );
  XNOR2_X1 U14596 ( .A(n12177), .B(n12538), .ZN(n12178) );
  XNOR2_X1 U14597 ( .A(n12179), .B(n12178), .ZN(n12171) );
  NAND2_X1 U14598 ( .A1(n12171), .A2(n12499), .ZN(n12176) );
  AOI22_X1 U14599 ( .A1(n12691), .A2(n12525), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12172) );
  OAI21_X1 U14600 ( .B1(n12173), .B2(n12461), .A(n12172), .ZN(n12174) );
  AOI21_X1 U14601 ( .B1(n12503), .B2(n12537), .A(n12174), .ZN(n12175) );
  OAI211_X1 U14602 ( .C1(n12830), .C2(n12528), .A(n12176), .B(n12175), .ZN(
        P3_U3154) );
  AOI22_X1 U14603 ( .A1(n12179), .A2(n12178), .B1(n12676), .B2(n12177), .ZN(
        n12182) );
  XNOR2_X1 U14604 ( .A(n12321), .B(n12180), .ZN(n12181) );
  XNOR2_X1 U14605 ( .A(n12182), .B(n12181), .ZN(n12189) );
  INV_X1 U14606 ( .A(n12183), .ZN(n12665) );
  OAI22_X1 U14607 ( .A1(n12665), .A2(n12461), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12184), .ZN(n12187) );
  OAI22_X1 U14608 ( .A1(n12185), .A2(n12527), .B1(n12676), .B2(n12505), .ZN(
        n12186) );
  AOI211_X1 U14609 ( .C1(n12670), .C2(n12515), .A(n12187), .B(n12186), .ZN(
        n12188) );
  OAI21_X1 U14610 ( .B1(n12189), .B2(n12534), .A(n12188), .ZN(P3_U3160) );
  AND2_X1 U14611 ( .A1(n12190), .A2(n12204), .ZN(n12208) );
  NAND2_X1 U14612 ( .A1(n12191), .A2(n12317), .ZN(n12192) );
  AOI211_X1 U14613 ( .C1(n12195), .C2(n12194), .A(n12193), .B(n12192), .ZN(
        n12202) );
  XNOR2_X1 U14614 ( .A(n12196), .B(n12317), .ZN(n12197) );
  AOI21_X1 U14615 ( .B1(n12199), .B2(n12198), .A(n12197), .ZN(n12201) );
  NOR3_X1 U14616 ( .A1(n12202), .A2(n12201), .A3(n12200), .ZN(n12206) );
  AOI21_X1 U14617 ( .B1(n12210), .B2(n12203), .A(n12327), .ZN(n12205) );
  OAI21_X1 U14618 ( .B1(n12206), .B2(n12205), .A(n12204), .ZN(n12207) );
  OAI21_X1 U14619 ( .B1(n12208), .B2(n12317), .A(n12207), .ZN(n12209) );
  OAI211_X1 U14620 ( .C1(n12210), .C2(n12317), .A(n12209), .B(n12363), .ZN(
        n12214) );
  MUX2_X1 U14621 ( .A(n12212), .B(n12211), .S(n12317), .Z(n12213) );
  AND3_X1 U14622 ( .A1(n12214), .A2(n12358), .A3(n12213), .ZN(n12224) );
  NAND2_X1 U14623 ( .A1(n12220), .A2(n12215), .ZN(n12218) );
  NAND2_X1 U14624 ( .A1(n12219), .A2(n12216), .ZN(n12217) );
  MUX2_X1 U14625 ( .A(n12218), .B(n12217), .S(n12327), .Z(n12223) );
  MUX2_X1 U14626 ( .A(n12220), .B(n12219), .S(n12317), .Z(n12221) );
  OAI211_X1 U14627 ( .C1(n12224), .C2(n12223), .A(n12222), .B(n12221), .ZN(
        n12228) );
  MUX2_X1 U14628 ( .A(n12226), .B(n12225), .S(n12327), .Z(n12227) );
  NAND3_X1 U14629 ( .A1(n12228), .A2(n12365), .A3(n12227), .ZN(n12239) );
  NOR2_X1 U14630 ( .A1(n12229), .A2(n12327), .ZN(n12232) );
  NOR2_X1 U14631 ( .A1(n12230), .A2(n12317), .ZN(n12231) );
  MUX2_X1 U14632 ( .A(n12232), .B(n12231), .S(n12551), .Z(n12233) );
  NOR2_X1 U14633 ( .A1(n12360), .A2(n12233), .ZN(n12238) );
  MUX2_X1 U14634 ( .A(n12235), .B(n12234), .S(n12317), .Z(n12236) );
  AOI22_X1 U14635 ( .A1(n12239), .A2(n12238), .B1(n12237), .B2(n12236), .ZN(
        n12244) );
  MUX2_X1 U14636 ( .A(n12241), .B(n12240), .S(n12327), .Z(n12242) );
  OAI211_X1 U14637 ( .C1(n12244), .C2(n12243), .A(n12374), .B(n12242), .ZN(
        n12245) );
  INV_X1 U14638 ( .A(n12245), .ZN(n12254) );
  OAI21_X1 U14639 ( .B1(n7425), .B2(n12246), .A(n12251), .ZN(n12249) );
  NAND2_X1 U14640 ( .A1(n12250), .A2(n12247), .ZN(n12248) );
  MUX2_X1 U14641 ( .A(n12249), .B(n12248), .S(n12317), .Z(n12253) );
  MUX2_X1 U14642 ( .A(n12251), .B(n12250), .S(n12327), .Z(n12252) );
  OAI211_X1 U14643 ( .C1(n12254), .C2(n12253), .A(n12372), .B(n12252), .ZN(
        n12259) );
  MUX2_X1 U14644 ( .A(n12256), .B(n12255), .S(n12317), .Z(n12257) );
  NAND3_X1 U14645 ( .A1(n12259), .A2(n12258), .A3(n12257), .ZN(n12263) );
  INV_X1 U14646 ( .A(n12263), .ZN(n12261) );
  OAI21_X1 U14647 ( .B1(n12261), .B2(n8936), .A(n12373), .ZN(n12268) );
  NAND3_X1 U14648 ( .A1(n12263), .A2(n12327), .A3(n12262), .ZN(n12266) );
  INV_X1 U14649 ( .A(n12271), .ZN(n12265) );
  AOI211_X1 U14650 ( .C1(n12266), .C2(n12373), .A(n12265), .B(n7055), .ZN(
        n12267) );
  AOI21_X1 U14651 ( .B1(n12317), .B2(n12268), .A(n12267), .ZN(n12274) );
  AOI21_X1 U14652 ( .B1(n12270), .B2(n12269), .A(n12327), .ZN(n12273) );
  MUX2_X1 U14653 ( .A(n12271), .B(n12270), .S(n12327), .Z(n12272) );
  OAI21_X1 U14654 ( .B1(n12274), .B2(n12273), .A(n12272), .ZN(n12281) );
  INV_X1 U14655 ( .A(n12275), .ZN(n12280) );
  INV_X1 U14656 ( .A(n12276), .ZN(n12277) );
  NAND2_X1 U14657 ( .A1(n12283), .A2(n12277), .ZN(n12278) );
  NAND4_X1 U14658 ( .A1(n12288), .A2(n12327), .A3(n12279), .A4(n12278), .ZN(
        n12282) );
  AOI22_X1 U14659 ( .A1(n12281), .A2(n12801), .B1(n12280), .B2(n12282), .ZN(
        n12286) );
  INV_X1 U14660 ( .A(n12282), .ZN(n12285) );
  AND3_X1 U14661 ( .A1(n12287), .A2(n12317), .A3(n12283), .ZN(n12284) );
  OAI22_X1 U14662 ( .A1(n12286), .A2(n12789), .B1(n12285), .B2(n12284), .ZN(
        n12291) );
  MUX2_X1 U14663 ( .A(n6869), .B(n9002), .S(n12317), .Z(n12289) );
  NOR2_X1 U14664 ( .A1(n12760), .A2(n12289), .ZN(n12290) );
  AOI21_X1 U14665 ( .B1(n12291), .B2(n12290), .A(n12748), .ZN(n12300) );
  MUX2_X1 U14666 ( .A(n12293), .B(n12292), .S(n12327), .Z(n12299) );
  INV_X1 U14667 ( .A(n12294), .ZN(n12297) );
  INV_X1 U14668 ( .A(n12295), .ZN(n12296) );
  MUX2_X1 U14669 ( .A(n12297), .B(n12296), .S(n12317), .Z(n12298) );
  NAND2_X1 U14670 ( .A1(n12302), .A2(n12306), .ZN(n12735) );
  AOI211_X1 U14671 ( .C1(n12300), .C2(n12299), .A(n12298), .B(n12735), .ZN(
        n12301) );
  OAI22_X1 U14672 ( .A1(n12301), .A2(n12724), .B1(n12317), .B2(n12304), .ZN(
        n12308) );
  INV_X1 U14673 ( .A(n12302), .ZN(n12303) );
  NAND2_X1 U14674 ( .A1(n12304), .A2(n12303), .ZN(n12305) );
  MUX2_X1 U14675 ( .A(n12306), .B(n12305), .S(n12327), .Z(n12307) );
  NAND2_X1 U14676 ( .A1(n12308), .A2(n12307), .ZN(n12309) );
  OAI21_X1 U14677 ( .B1(n12309), .B2(n12705), .A(n12696), .ZN(n12316) );
  INV_X1 U14678 ( .A(n12705), .ZN(n12711) );
  XNOR2_X1 U14679 ( .A(n12310), .B(n12327), .ZN(n12311) );
  AOI21_X1 U14680 ( .B1(n12711), .B2(n12312), .A(n12311), .ZN(n12315) );
  INV_X1 U14681 ( .A(n12673), .ZN(n12679) );
  MUX2_X1 U14682 ( .A(n12313), .B(n12680), .S(n12317), .Z(n12314) );
  OAI211_X1 U14683 ( .C1(n12316), .C2(n12315), .A(n12679), .B(n12314), .ZN(
        n12323) );
  MUX2_X1 U14684 ( .A(n12319), .B(n12318), .S(n12317), .Z(n12322) );
  NAND2_X1 U14685 ( .A1(n12321), .A2(n12320), .ZN(n12385) );
  AOI21_X1 U14686 ( .B1(n12323), .B2(n12322), .A(n12385), .ZN(n12330) );
  OAI22_X1 U14687 ( .A1(n12385), .A2(n12327), .B1(n12325), .B2(n12324), .ZN(
        n12326) );
  INV_X1 U14688 ( .A(n12326), .ZN(n12329) );
  NAND2_X1 U14689 ( .A1(n12330), .A2(n12327), .ZN(n12328) );
  OAI211_X1 U14690 ( .C1(n12330), .C2(n12329), .A(n12328), .B(n12393), .ZN(
        n12337) );
  NAND2_X1 U14691 ( .A1(n12331), .A2(n12343), .ZN(n12335) );
  OR2_X1 U14692 ( .A1(n12333), .A2(n12332), .ZN(n12334) );
  NOR2_X1 U14693 ( .A1(n14475), .A2(n12354), .ZN(n12400) );
  INV_X1 U14694 ( .A(n12400), .ZN(n12336) );
  NAND3_X1 U14695 ( .A1(n12337), .A2(n12397), .A3(n12336), .ZN(n12357) );
  NOR2_X1 U14696 ( .A1(n12338), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12339) );
  OAI22_X1 U14697 ( .A1(n12340), .A2(n12339), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n14366), .ZN(n12342) );
  XNOR2_X1 U14698 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12341) );
  XNOR2_X1 U14699 ( .A(n12342), .B(n12341), .ZN(n12928) );
  NAND2_X1 U14700 ( .A1(n12928), .A2(n12343), .ZN(n12345) );
  INV_X1 U14701 ( .A(SI_31_), .ZN(n12934) );
  OR2_X1 U14702 ( .A1(n12333), .A2(n12934), .ZN(n12344) );
  INV_X1 U14703 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12663) );
  NAND2_X1 U14704 ( .A1(n12346), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12349) );
  INV_X1 U14705 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12347) );
  OR2_X1 U14706 ( .A1(n6440), .A2(n12347), .ZN(n12348) );
  OAI211_X1 U14707 ( .C1(n12350), .C2(n12663), .A(n12349), .B(n12348), .ZN(
        n12351) );
  INV_X1 U14708 ( .A(n12351), .ZN(n12352) );
  OR2_X1 U14709 ( .A1(n12878), .A2(n12660), .ZN(n12356) );
  NAND2_X1 U14710 ( .A1(n14475), .A2(n12354), .ZN(n12355) );
  NAND2_X1 U14711 ( .A1(n12356), .A2(n12355), .ZN(n12396) );
  INV_X1 U14712 ( .A(n12396), .ZN(n12388) );
  AOI21_X1 U14713 ( .B1(n12357), .B2(n12388), .A(n12399), .ZN(n12410) );
  INV_X1 U14714 ( .A(n12774), .ZN(n12379) );
  INV_X1 U14715 ( .A(n12358), .ZN(n12361) );
  NOR4_X1 U14716 ( .A1(n12361), .A2(n12360), .A3(n12359), .A4(n10043), .ZN(
        n12364) );
  NAND4_X1 U14717 ( .A1(n12364), .A2(n15120), .A3(n12363), .A4(n12362), .ZN(
        n12371) );
  NAND4_X1 U14718 ( .A1(n12368), .A2(n12367), .A3(n12366), .A4(n12365), .ZN(
        n12369) );
  NOR3_X1 U14719 ( .A1(n12371), .A2(n12370), .A3(n12369), .ZN(n12375) );
  NAND4_X1 U14720 ( .A1(n12375), .A2(n12374), .A3(n12373), .A4(n12372), .ZN(
        n12377) );
  NOR3_X1 U14721 ( .A1(n12377), .A2(n12808), .A3(n12376), .ZN(n12378) );
  NAND4_X1 U14722 ( .A1(n12379), .A2(n12783), .A3(n12801), .A4(n12378), .ZN(
        n12380) );
  NOR4_X1 U14723 ( .A1(n12735), .A2(n12760), .A3(n12748), .A4(n12380), .ZN(
        n12381) );
  NAND4_X1 U14724 ( .A1(n12696), .A2(n12382), .A3(n12381), .A4(n12711), .ZN(
        n12383) );
  NOR4_X1 U14725 ( .A1(n12400), .A2(n12384), .A3(n12673), .A4(n12383), .ZN(
        n12389) );
  INV_X1 U14726 ( .A(n12385), .ZN(n12387) );
  INV_X1 U14727 ( .A(n12399), .ZN(n12386) );
  NAND4_X1 U14728 ( .A1(n12389), .A2(n12388), .A3(n12387), .A4(n12386), .ZN(
        n12390) );
  XNOR2_X1 U14729 ( .A(n12390), .B(n12654), .ZN(n12391) );
  OAI22_X1 U14730 ( .A1(n12410), .A2(n15130), .B1(n12392), .B2(n12391), .ZN(
        n12409) );
  INV_X1 U14731 ( .A(n14475), .ZN(n12394) );
  INV_X1 U14732 ( .A(n12660), .ZN(n12536) );
  OAI21_X1 U14733 ( .B1(n12394), .B2(n12536), .A(n12393), .ZN(n12395) );
  NOR2_X1 U14734 ( .A1(n12407), .A2(n12406), .ZN(n12408) );
  NAND3_X1 U14735 ( .A1(n12413), .A2(n12412), .A3(n12646), .ZN(n12414) );
  OAI211_X1 U14736 ( .C1(n12415), .C2(n12417), .A(n12414), .B(P3_B_REG_SCAN_IN), .ZN(n12416) );
  OAI21_X1 U14737 ( .B1(n12418), .B2(n12417), .A(n12416), .ZN(P3_U3296) );
  NOR2_X1 U14738 ( .A1(n12420), .A2(n12816), .ZN(n12661) );
  AOI21_X1 U14739 ( .B1(n15136), .B2(P3_REG2_REG_29__SCAN_IN), .A(n12661), 
        .ZN(n12421) );
  OAI21_X1 U14740 ( .B1(n12422), .B2(n12815), .A(n12421), .ZN(n12423) );
  AOI21_X1 U14741 ( .B1(n12424), .B2(n12821), .A(n12423), .ZN(n12425) );
  OAI21_X1 U14742 ( .B1(n12419), .B2(n15136), .A(n12425), .ZN(P3_U3204) );
  XNOR2_X1 U14743 ( .A(n12426), .B(n12539), .ZN(n12431) );
  AOI22_X1 U14744 ( .A1(n12720), .A2(n12503), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12428) );
  NAND2_X1 U14745 ( .A1(n12531), .A2(n12726), .ZN(n12427) );
  OAI211_X1 U14746 ( .C1(n12747), .C2(n12505), .A(n12428), .B(n12427), .ZN(
        n12429) );
  AOI21_X1 U14747 ( .B1(n12725), .B2(n12515), .A(n12429), .ZN(n12430) );
  OAI21_X1 U14748 ( .B1(n12431), .B2(n12534), .A(n12430), .ZN(P3_U3156) );
  INV_X1 U14749 ( .A(n12432), .ZN(n12433) );
  AOI21_X1 U14750 ( .B1(n12435), .B2(n12434), .A(n12433), .ZN(n12441) );
  AOI22_X1 U14751 ( .A1(n12770), .A2(n12503), .B1(P3_REG3_REG_19__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12437) );
  NAND2_X1 U14752 ( .A1(n12543), .A2(n12525), .ZN(n12436) );
  OAI211_X1 U14753 ( .C1(n12775), .C2(n12461), .A(n12437), .B(n12436), .ZN(
        n12438) );
  AOI21_X1 U14754 ( .B1(n12439), .B2(n12515), .A(n12438), .ZN(n12440) );
  OAI21_X1 U14755 ( .B1(n12441), .B2(n12534), .A(n12440), .ZN(P3_U3159) );
  AOI21_X1 U14756 ( .B1(n12443), .B2(n12442), .A(n6585), .ZN(n12448) );
  AOI22_X1 U14757 ( .A1(n12770), .A2(n12525), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12445) );
  NAND2_X1 U14758 ( .A1(n12531), .A2(n12751), .ZN(n12444) );
  OAI211_X1 U14759 ( .C1(n12747), .C2(n12527), .A(n12445), .B(n12444), .ZN(
        n12446) );
  AOI21_X1 U14760 ( .B1(n12750), .B2(n12515), .A(n12446), .ZN(n12447) );
  OAI21_X1 U14761 ( .B1(n12448), .B2(n12534), .A(n12447), .ZN(P3_U3163) );
  XOR2_X1 U14762 ( .A(n12450), .B(n12449), .Z(n12456) );
  AOI22_X1 U14763 ( .A1(n12720), .A2(n12525), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12452) );
  NAND2_X1 U14764 ( .A1(n12699), .A2(n12531), .ZN(n12451) );
  OAI211_X1 U14765 ( .C1(n12453), .C2(n12527), .A(n12452), .B(n12451), .ZN(
        n12454) );
  AOI21_X1 U14766 ( .B1(n12698), .B2(n12515), .A(n12454), .ZN(n12455) );
  OAI21_X1 U14767 ( .B1(n12456), .B2(n12534), .A(n12455), .ZN(P3_U3165) );
  XOR2_X1 U14768 ( .A(n12458), .B(n12457), .Z(n12465) );
  AOI22_X1 U14769 ( .A1(n12503), .A2(n12544), .B1(P3_REG3_REG_16__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12460) );
  NAND2_X1 U14770 ( .A1(n12525), .A2(n12546), .ZN(n12459) );
  OAI211_X1 U14771 ( .C1(n12817), .C2(n12461), .A(n12460), .B(n12459), .ZN(
        n12462) );
  AOI21_X1 U14772 ( .B1(n12463), .B2(n12515), .A(n12462), .ZN(n12464) );
  OAI21_X1 U14773 ( .B1(n12465), .B2(n12534), .A(n12464), .ZN(P3_U3166) );
  AOI21_X1 U14774 ( .B1(n12467), .B2(n12466), .A(n12534), .ZN(n12468) );
  OR2_X1 U14775 ( .A1(n12467), .A2(n12466), .ZN(n12498) );
  NAND2_X1 U14776 ( .A1(n12468), .A2(n12498), .ZN(n12474) );
  INV_X1 U14777 ( .A(n12803), .ZN(n12472) );
  NOR2_X1 U14778 ( .A1(n12469), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14446) );
  AOI21_X1 U14779 ( .B1(n12543), .B2(n12503), .A(n14446), .ZN(n12470) );
  OAI21_X1 U14780 ( .B1(n12798), .B2(n12505), .A(n12470), .ZN(n12471) );
  AOI21_X1 U14781 ( .B1(n12472), .B2(n12531), .A(n12471), .ZN(n12473) );
  OAI211_X1 U14782 ( .C1(n12528), .C2(n12918), .A(n12474), .B(n12473), .ZN(
        P3_U3168) );
  XOR2_X1 U14783 ( .A(n12476), .B(n12475), .Z(n12481) );
  AOI22_X1 U14784 ( .A1(n12539), .A2(n12525), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12478) );
  NAND2_X1 U14785 ( .A1(n12531), .A2(n12713), .ZN(n12477) );
  OAI211_X1 U14786 ( .C1(n12677), .C2(n12527), .A(n12478), .B(n12477), .ZN(
        n12479) );
  AOI21_X1 U14787 ( .B1(n12712), .B2(n12515), .A(n12479), .ZN(n12480) );
  OAI21_X1 U14788 ( .B1(n12481), .B2(n12534), .A(n12480), .ZN(P3_U3169) );
  INV_X1 U14789 ( .A(n12482), .ZN(n12906) );
  AOI21_X1 U14790 ( .B1(n12484), .B2(n12483), .A(n12534), .ZN(n12486) );
  NAND2_X1 U14791 ( .A1(n12486), .A2(n12485), .ZN(n12490) );
  AOI22_X1 U14792 ( .A1(n12541), .A2(n12503), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12487) );
  OAI21_X1 U14793 ( .B1(n12785), .B2(n12505), .A(n12487), .ZN(n12488) );
  AOI21_X1 U14794 ( .B1(n12761), .B2(n12531), .A(n12488), .ZN(n12489) );
  OAI211_X1 U14795 ( .C1(n12906), .C2(n12528), .A(n12490), .B(n12489), .ZN(
        P3_U3173) );
  XNOR2_X1 U14796 ( .A(n12491), .B(n12540), .ZN(n12496) );
  AOI22_X1 U14797 ( .A1(n12541), .A2(n12525), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12493) );
  NAND2_X1 U14798 ( .A1(n12531), .A2(n12737), .ZN(n12492) );
  OAI211_X1 U14799 ( .C1(n12733), .C2(n12527), .A(n12493), .B(n12492), .ZN(
        n12494) );
  AOI21_X1 U14800 ( .B1(n12736), .B2(n12515), .A(n12494), .ZN(n12495) );
  OAI21_X1 U14801 ( .B1(n12496), .B2(n12534), .A(n12495), .ZN(P3_U3175) );
  NAND2_X1 U14802 ( .A1(n12498), .A2(n12497), .ZN(n12502) );
  OAI211_X1 U14803 ( .C1(n12502), .C2(n12501), .A(n12500), .B(n12499), .ZN(
        n12509) );
  INV_X1 U14804 ( .A(n12790), .ZN(n12507) );
  AND2_X1 U14805 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n14463) );
  AOI21_X1 U14806 ( .B1(n12542), .B2(n12503), .A(n14463), .ZN(n12504) );
  OAI21_X1 U14807 ( .B1(n12812), .B2(n12505), .A(n12504), .ZN(n12506) );
  AOI21_X1 U14808 ( .B1(n12507), .B2(n12531), .A(n12506), .ZN(n12508) );
  OAI211_X1 U14809 ( .C1(n12914), .C2(n12528), .A(n12509), .B(n12508), .ZN(
        P3_U3178) );
  XOR2_X1 U14810 ( .A(n12511), .B(n12510), .Z(n12518) );
  AOI22_X1 U14811 ( .A1(n12707), .A2(n12525), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12513) );
  NAND2_X1 U14812 ( .A1(n12683), .A2(n12531), .ZN(n12512) );
  OAI211_X1 U14813 ( .C1(n12676), .C2(n12527), .A(n12513), .B(n12512), .ZN(
        n12514) );
  AOI21_X1 U14814 ( .B1(n12516), .B2(n12515), .A(n12514), .ZN(n12517) );
  OAI21_X1 U14815 ( .B1(n12518), .B2(n12534), .A(n12517), .ZN(P3_U3180) );
  NAND2_X1 U14816 ( .A1(n12520), .A2(n12519), .ZN(n12524) );
  NAND2_X1 U14817 ( .A1(n12522), .A2(n12521), .ZN(n12523) );
  XOR2_X1 U14818 ( .A(n12524), .B(n12523), .Z(n12535) );
  NAND2_X1 U14819 ( .A1(n12525), .A2(n12547), .ZN(n12526) );
  NAND2_X1 U14820 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n14409)
         );
  OAI211_X1 U14821 ( .C1(n12798), .C2(n12527), .A(n12526), .B(n14409), .ZN(
        n12530) );
  NOR2_X1 U14822 ( .A1(n12925), .A2(n12528), .ZN(n12529) );
  AOI211_X1 U14823 ( .C1(n12532), .C2(n12531), .A(n12530), .B(n12529), .ZN(
        n12533) );
  OAI21_X1 U14824 ( .B1(n12535), .B2(n12534), .A(n12533), .ZN(P3_U3181) );
  MUX2_X1 U14825 ( .A(n12536), .B(P3_DATAO_REG_31__SCAN_IN), .S(n12558), .Z(
        P3_U3522) );
  MUX2_X1 U14826 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12537), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14827 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12538), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14828 ( .A(n12691), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12558), .Z(
        P3_U3517) );
  MUX2_X1 U14829 ( .A(n12707), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12558), .Z(
        P3_U3516) );
  MUX2_X1 U14830 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12720), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14831 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n12539), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U14832 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12540), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14833 ( .A(n12541), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12558), .Z(
        P3_U3512) );
  MUX2_X1 U14834 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12542), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14835 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12543), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14836 ( .A(n12544), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12558), .Z(
        P3_U3508) );
  MUX2_X1 U14837 ( .A(n12545), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12558), .Z(
        P3_U3507) );
  MUX2_X1 U14838 ( .A(n12546), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12558), .Z(
        P3_U3506) );
  MUX2_X1 U14839 ( .A(n12547), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12558), .Z(
        P3_U3505) );
  MUX2_X1 U14840 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12548), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14841 ( .A(n12549), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12558), .Z(
        P3_U3502) );
  MUX2_X1 U14842 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12550), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14843 ( .A(n12551), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12558), .Z(
        P3_U3499) );
  MUX2_X1 U14844 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12552), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14845 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12553), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14846 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12554), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14847 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12555), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14848 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12556), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14849 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n10051), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14850 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12557), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14851 ( .A(n12559), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12558), .Z(
        P3_U3491) );
  INV_X1 U14852 ( .A(n12643), .ZN(n14438) );
  INV_X1 U14853 ( .A(n15084), .ZN(n12629) );
  NAND2_X2 U14854 ( .A1(n12561), .A2(n12560), .ZN(n12564) );
  NOR2_X1 U14855 ( .A1(n12563), .A2(n12562), .ZN(n12565) );
  INV_X1 U14856 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15010) );
  INV_X1 U14857 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n12607) );
  OR2_X1 U14858 ( .A1(n12617), .A2(n12607), .ZN(n12567) );
  NAND2_X1 U14859 ( .A1(n12617), .A2(n12607), .ZN(n12566) );
  NAND2_X1 U14860 ( .A1(n12567), .A2(n12566), .ZN(n15026) );
  NOR2_X1 U14861 ( .A1(n12605), .A2(n12568), .ZN(n12569) );
  NOR2_X1 U14862 ( .A1(n12569), .A2(n15043), .ZN(n15062) );
  MUX2_X1 U14863 ( .A(n12620), .B(P3_REG2_REG_12__SCAN_IN), .S(n15068), .Z(
        n15061) );
  NAND2_X1 U14864 ( .A1(n15068), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12570) );
  NOR2_X1 U14865 ( .A1(n12629), .A2(n12571), .ZN(n12572) );
  NOR2_X1 U14866 ( .A1(n12572), .A2(n15077), .ZN(n15097) );
  NAND2_X1 U14867 ( .A1(n15100), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12635) );
  OR2_X1 U14868 ( .A1(n15100), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12573) );
  NAND2_X1 U14869 ( .A1(n12635), .A2(n12573), .ZN(n15096) );
  NOR2_X1 U14870 ( .A1(n15097), .A2(n15096), .ZN(n15095) );
  AND2_X1 U14871 ( .A1(n14408), .A2(n12574), .ZN(n12575) );
  INV_X1 U14872 ( .A(n14408), .ZN(n12637) );
  INV_X1 U14873 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12576) );
  AOI22_X1 U14874 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n14421), .B1(n12641), 
        .B2(n12576), .ZN(n14432) );
  AOI21_X2 U14875 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n12641), .A(n14433), 
        .ZN(n12577) );
  XNOR2_X1 U14876 ( .A(n14438), .B(n12577), .ZN(n14447) );
  NAND2_X1 U14877 ( .A1(n6743), .A2(n12791), .ZN(n12579) );
  NAND2_X1 U14878 ( .A1(n14454), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12578) );
  AND2_X1 U14879 ( .A1(n12579), .A2(n12578), .ZN(n14465) );
  OR2_X1 U14880 ( .A1(n14454), .A2(n12791), .ZN(n12580) );
  MUX2_X1 U14881 ( .A(P3_REG2_REG_19__SCAN_IN), .B(n12776), .S(n12654), .Z(
        n12647) );
  INV_X1 U14882 ( .A(n12647), .ZN(n12581) );
  AOI22_X1 U14883 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12641), .B1(n14421), 
        .B2(n12871), .ZN(n14429) );
  INV_X1 U14884 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14491) );
  NAND2_X1 U14885 ( .A1(n15033), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n12588) );
  MUX2_X1 U14886 ( .A(n12583), .B(P3_REG1_REG_10__SCAN_IN), .S(n12617), .Z(
        n15029) );
  NAND2_X1 U14887 ( .A1(n12609), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n12585) );
  NAND2_X1 U14888 ( .A1(n15014), .A2(n12586), .ZN(n12587) );
  NAND2_X1 U14889 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n15019), .ZN(n15018) );
  NAND2_X1 U14890 ( .A1(n12587), .A2(n15018), .ZN(n15030) );
  NAND2_X1 U14891 ( .A1(n15029), .A2(n15030), .ZN(n15028) );
  NAND2_X1 U14892 ( .A1(n15049), .A2(n12589), .ZN(n12590) );
  NAND2_X1 U14893 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n15046), .ZN(n15045) );
  NAND2_X1 U14894 ( .A1(n12590), .A2(n15045), .ZN(n15065) );
  MUX2_X1 U14895 ( .A(P3_REG1_REG_12__SCAN_IN), .B(n14491), .S(n15068), .Z(
        n15064) );
  NAND2_X1 U14896 ( .A1(n15065), .A2(n15064), .ZN(n15063) );
  NAND2_X1 U14897 ( .A1(n15084), .A2(n12591), .ZN(n12592) );
  XNOR2_X1 U14898 ( .A(n15100), .B(P3_REG1_REG_14__SCAN_IN), .ZN(n15099) );
  INV_X1 U14899 ( .A(n15100), .ZN(n12593) );
  INV_X1 U14900 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n14481) );
  NAND2_X1 U14901 ( .A1(n14408), .A2(n12594), .ZN(n12595) );
  XNOR2_X1 U14902 ( .A(n12637), .B(n12594), .ZN(n14407) );
  NAND2_X1 U14903 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n14407), .ZN(n14406) );
  NAND2_X1 U14904 ( .A1(n12595), .A2(n14406), .ZN(n14428) );
  NAND2_X1 U14905 ( .A1(n14429), .A2(n14428), .ZN(n14427) );
  NAND2_X1 U14906 ( .A1(n12643), .A2(n12596), .ZN(n12597) );
  NAND2_X1 U14907 ( .A1(n12597), .A2(n14439), .ZN(n14456) );
  XNOR2_X1 U14908 ( .A(n14454), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n14455) );
  AOI22_X1 U14909 ( .A1(n14456), .A2(n14455), .B1(P3_REG1_REG_18__SCAN_IN), 
        .B2(n6743), .ZN(n12598) );
  XNOR2_X1 U14910 ( .A(n12654), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12645) );
  XNOR2_X1 U14911 ( .A(n12598), .B(n12645), .ZN(n12657) );
  NAND2_X1 U14912 ( .A1(n12646), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n12599) );
  OAI21_X1 U14913 ( .B1(n12646), .B2(n14448), .A(n12599), .ZN(n12644) );
  OR2_X1 U14914 ( .A1(n12646), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12601) );
  AOI21_X1 U14915 ( .B1(n12646), .B2(n12871), .A(n14421), .ZN(n12600) );
  AND2_X1 U14916 ( .A1(n12601), .A2(n12600), .ZN(n14422) );
  OR2_X1 U14917 ( .A1(n12646), .A2(n12602), .ZN(n12604) );
  NAND2_X1 U14918 ( .A1(n12646), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n12603) );
  NAND2_X1 U14919 ( .A1(n12604), .A2(n12603), .ZN(n12618) );
  XNOR2_X1 U14920 ( .A(n12618), .B(n12605), .ZN(n15054) );
  NAND2_X1 U14921 ( .A1(n12646), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n12606) );
  OAI21_X1 U14922 ( .B1(n12646), .B2(n12607), .A(n12606), .ZN(n12616) );
  NAND2_X1 U14923 ( .A1(n10514), .A2(n15010), .ZN(n12608) );
  OAI211_X1 U14924 ( .C1(n10514), .C2(P3_REG1_REG_9__SCAN_IN), .A(n12608), .B(
        n15014), .ZN(n15011) );
  INV_X1 U14925 ( .A(n12609), .ZN(n12610) );
  NAND2_X1 U14926 ( .A1(n12611), .A2(n12610), .ZN(n12613) );
  NAND2_X1 U14927 ( .A1(n12613), .A2(n12612), .ZN(n15013) );
  OR2_X1 U14928 ( .A1(n12646), .A2(n15010), .ZN(n12615) );
  AOI21_X1 U14929 ( .B1(n12646), .B2(P3_REG1_REG_9__SCAN_IN), .A(n15014), .ZN(
        n12614) );
  XOR2_X1 U14930 ( .A(n12617), .B(n12616), .Z(n15035) );
  NAND2_X1 U14931 ( .A1(n15054), .A2(n15053), .ZN(n15052) );
  OR2_X1 U14932 ( .A1(n12618), .A2(n15049), .ZN(n12619) );
  OR2_X1 U14933 ( .A1(n12646), .A2(n12620), .ZN(n12622) );
  NAND2_X1 U14934 ( .A1(n12646), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n12621) );
  NAND2_X1 U14935 ( .A1(n12622), .A2(n12621), .ZN(n12624) );
  XNOR2_X1 U14936 ( .A(n12624), .B(n12623), .ZN(n15072) );
  NAND2_X1 U14937 ( .A1(n15073), .A2(n15072), .ZN(n15071) );
  NAND2_X1 U14938 ( .A1(n12624), .A2(n15068), .ZN(n12625) );
  OR2_X1 U14939 ( .A1(n12646), .A2(n12626), .ZN(n12628) );
  NAND2_X1 U14940 ( .A1(n12646), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n12627) );
  NAND2_X1 U14941 ( .A1(n12628), .A2(n12627), .ZN(n12630) );
  XNOR2_X1 U14942 ( .A(n12630), .B(n12629), .ZN(n15089) );
  OR2_X1 U14943 ( .A1(n12630), .A2(n15084), .ZN(n12631) );
  INV_X1 U14944 ( .A(n15096), .ZN(n12633) );
  NAND2_X1 U14945 ( .A1(n12646), .A2(n15099), .ZN(n12632) );
  OAI21_X1 U14946 ( .B1(n12646), .B2(n12633), .A(n12632), .ZN(n15110) );
  NAND3_X1 U14947 ( .A1(n12646), .A2(P3_REG1_REG_14__SCAN_IN), .A3(n15100), 
        .ZN(n12634) );
  OAI21_X1 U14948 ( .B1(n12646), .B2(n12635), .A(n12634), .ZN(n12636) );
  NOR2_X1 U14949 ( .A1(n12638), .A2(n12637), .ZN(n12639) );
  NOR2_X1 U14950 ( .A1(n12640), .A2(n12639), .ZN(n14415) );
  MUX2_X1 U14951 ( .A(n14405), .B(n14335), .S(n12646), .Z(n14414) );
  AND2_X1 U14952 ( .A1(n14415), .A2(n14414), .ZN(n14417) );
  NOR2_X1 U14953 ( .A1(n12640), .A2(n14417), .ZN(n14426) );
  AOI21_X1 U14954 ( .B1(n12646), .B2(P3_REG1_REG_16__SCAN_IN), .A(n12641), 
        .ZN(n12642) );
  OAI21_X1 U14955 ( .B1(n12646), .B2(n12576), .A(n12642), .ZN(n14424) );
  OAI21_X1 U14956 ( .B1(n14422), .B2(n14426), .A(n14424), .ZN(n14443) );
  XNOR2_X1 U14957 ( .A(n12644), .B(n12643), .ZN(n14442) );
  NOR2_X1 U14958 ( .A1(n14443), .A2(n14442), .ZN(n14441) );
  MUX2_X1 U14959 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12646), .Z(n14459) );
  NOR2_X1 U14960 ( .A1(n14458), .A2(n14459), .ZN(n14457) );
  INV_X1 U14961 ( .A(n12645), .ZN(n12648) );
  MUX2_X1 U14962 ( .A(n12648), .B(n12647), .S(n10514), .Z(n12649) );
  XNOR2_X1 U14963 ( .A(n12650), .B(n12649), .ZN(n12651) );
  NOR2_X1 U14964 ( .A1(n12651), .A2(n15109), .ZN(n12656) );
  NAND2_X1 U14965 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(P3_U3151), .ZN(n12653)
         );
  NAND2_X1 U14966 ( .A1(n15082), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12652) );
  OAI211_X1 U14967 ( .C1(n15101), .C2(n12654), .A(n12653), .B(n12652), .ZN(
        n12655) );
  NAND2_X1 U14968 ( .A1(n12878), .A2(n14471), .ZN(n12662) );
  AOI21_X1 U14969 ( .B1(n14474), .B2(n12818), .A(n12661), .ZN(n14473) );
  OAI211_X1 U14970 ( .C1(n12663), .C2(n12818), .A(n12662), .B(n14473), .ZN(
        P3_U3202) );
  OAI22_X1 U14971 ( .A1(n12665), .A2(n12816), .B1(n12818), .B2(n12664), .ZN(
        n12669) );
  NOR2_X1 U14972 ( .A1(n12667), .A2(n12666), .ZN(n12668) );
  AOI211_X1 U14973 ( .C1(n14471), .C2(n12670), .A(n12669), .B(n12668), .ZN(
        n12671) );
  OAI21_X1 U14974 ( .B1(n12672), .B2(n15136), .A(n12671), .ZN(P3_U3205) );
  XNOR2_X1 U14975 ( .A(n12674), .B(n12673), .ZN(n12675) );
  OAI222_X1 U14976 ( .A1(n12799), .A2(n12677), .B1(n15122), .B2(n12676), .C1(
        n12675), .C2(n15128), .ZN(n12831) );
  INV_X1 U14977 ( .A(n12831), .ZN(n12687) );
  INV_X1 U14978 ( .A(n12678), .ZN(n12682) );
  AOI21_X1 U14979 ( .B1(n12695), .B2(n12680), .A(n12679), .ZN(n12681) );
  NOR2_X1 U14980 ( .A1(n12682), .A2(n12681), .ZN(n12832) );
  AOI22_X1 U14981 ( .A1(n12683), .A2(n15134), .B1(n15136), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12684) );
  OAI21_X1 U14982 ( .B1(n12884), .B2(n12815), .A(n12684), .ZN(n12685) );
  AOI21_X1 U14983 ( .B1(n12832), .B2(n12821), .A(n12685), .ZN(n12686) );
  OAI21_X1 U14984 ( .B1(n12687), .B2(n15136), .A(n12686), .ZN(P3_U3207) );
  OAI211_X1 U14985 ( .C1(n12690), .C2(n12689), .A(n12688), .B(n12766), .ZN(
        n12693) );
  NAND2_X1 U14986 ( .A1(n12691), .A2(n12769), .ZN(n12692) );
  OAI211_X1 U14987 ( .C1(n12694), .C2(n12799), .A(n12693), .B(n12692), .ZN(
        n12835) );
  INV_X1 U14988 ( .A(n12835), .ZN(n12703) );
  OAI21_X1 U14989 ( .B1(n12697), .B2(n12696), .A(n12695), .ZN(n12836) );
  INV_X1 U14990 ( .A(n12698), .ZN(n12888) );
  AOI22_X1 U14991 ( .A1(n12699), .A2(n15134), .B1(n15136), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12700) );
  OAI21_X1 U14992 ( .B1(n12888), .B2(n12815), .A(n12700), .ZN(n12701) );
  AOI21_X1 U14993 ( .B1(n12836), .B2(n12821), .A(n12701), .ZN(n12702) );
  OAI21_X1 U14994 ( .B1(n12703), .B2(n15136), .A(n12702), .ZN(P3_U3208) );
  OAI211_X1 U14995 ( .C1(n12706), .C2(n12705), .A(n12704), .B(n12766), .ZN(
        n12709) );
  NAND2_X1 U14996 ( .A1(n12707), .A2(n12769), .ZN(n12708) );
  OAI211_X1 U14997 ( .C1(n12733), .C2(n12799), .A(n12709), .B(n12708), .ZN(
        n12838) );
  INV_X1 U14998 ( .A(n12838), .ZN(n12717) );
  OAI21_X1 U14999 ( .B1(n6510), .B2(n12711), .A(n12710), .ZN(n12839) );
  INV_X1 U15000 ( .A(n12712), .ZN(n12892) );
  AOI22_X1 U15001 ( .A1(n12713), .A2(n15134), .B1(n15136), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n12714) );
  OAI21_X1 U15002 ( .B1(n12892), .B2(n12815), .A(n12714), .ZN(n12715) );
  AOI21_X1 U15003 ( .B1(n12839), .B2(n12821), .A(n12715), .ZN(n12716) );
  OAI21_X1 U15004 ( .B1(n12717), .B2(n15136), .A(n12716), .ZN(P3_U3209) );
  OAI211_X1 U15005 ( .C1(n12719), .C2(n12724), .A(n12718), .B(n12766), .ZN(
        n12722) );
  NAND2_X1 U15006 ( .A1(n12720), .A2(n12769), .ZN(n12721) );
  OAI211_X1 U15007 ( .C1(n12747), .C2(n12799), .A(n12722), .B(n12721), .ZN(
        n12842) );
  INV_X1 U15008 ( .A(n12842), .ZN(n12730) );
  XNOR2_X1 U15009 ( .A(n12723), .B(n12724), .ZN(n12843) );
  INV_X1 U15010 ( .A(n12725), .ZN(n12895) );
  AOI22_X1 U15011 ( .A1(P3_REG2_REG_23__SCAN_IN), .A2(n15136), .B1(n12726), 
        .B2(n15134), .ZN(n12727) );
  OAI21_X1 U15012 ( .B1(n12895), .B2(n12815), .A(n12727), .ZN(n12728) );
  AOI21_X1 U15013 ( .B1(n12843), .B2(n12821), .A(n12728), .ZN(n12729) );
  OAI21_X1 U15014 ( .B1(n12730), .B2(n15136), .A(n12729), .ZN(P3_U3210) );
  XOR2_X1 U15015 ( .A(n12735), .B(n12731), .Z(n12732) );
  OAI222_X1 U15016 ( .A1(n15122), .A2(n12733), .B1(n12799), .B2(n12758), .C1(
        n15128), .C2(n12732), .ZN(n12846) );
  INV_X1 U15017 ( .A(n12846), .ZN(n12741) );
  XNOR2_X1 U15018 ( .A(n12734), .B(n12735), .ZN(n12847) );
  INV_X1 U15019 ( .A(n12736), .ZN(n12898) );
  AOI22_X1 U15020 ( .A1(n15136), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15134), 
        .B2(n12737), .ZN(n12738) );
  OAI21_X1 U15021 ( .B1(n12898), .B2(n12815), .A(n12738), .ZN(n12739) );
  AOI21_X1 U15022 ( .B1(n12847), .B2(n12821), .A(n12739), .ZN(n12740) );
  OAI21_X1 U15023 ( .B1(n12741), .B2(n15136), .A(n12740), .ZN(P3_U3211) );
  OAI21_X1 U15024 ( .B1(n12743), .B2(n12748), .A(n12742), .ZN(n12744) );
  INV_X1 U15025 ( .A(n12744), .ZN(n12745) );
  OAI222_X1 U15026 ( .A1(n15122), .A2(n12747), .B1(n12799), .B2(n12746), .C1(
        n15128), .C2(n12745), .ZN(n12850) );
  INV_X1 U15027 ( .A(n12850), .ZN(n12755) );
  XNOR2_X1 U15028 ( .A(n12749), .B(n12748), .ZN(n12851) );
  INV_X1 U15029 ( .A(n12750), .ZN(n12902) );
  AOI22_X1 U15030 ( .A1(n15136), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15134), 
        .B2(n12751), .ZN(n12752) );
  OAI21_X1 U15031 ( .B1(n12902), .B2(n12815), .A(n12752), .ZN(n12753) );
  AOI21_X1 U15032 ( .B1(n12851), .B2(n12821), .A(n12753), .ZN(n12754) );
  OAI21_X1 U15033 ( .B1(n12755), .B2(n15136), .A(n12754), .ZN(P3_U3212) );
  XNOR2_X1 U15034 ( .A(n12756), .B(n12760), .ZN(n12757) );
  OAI222_X1 U15035 ( .A1(n15122), .A2(n12758), .B1(n12799), .B2(n12785), .C1(
        n12757), .C2(n15128), .ZN(n12853) );
  INV_X1 U15036 ( .A(n12853), .ZN(n12765) );
  XOR2_X1 U15037 ( .A(n12760), .B(n12759), .Z(n12854) );
  AOI22_X1 U15038 ( .A1(n15136), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15134), 
        .B2(n12761), .ZN(n12762) );
  OAI21_X1 U15039 ( .B1(n12906), .B2(n12815), .A(n12762), .ZN(n12763) );
  AOI21_X1 U15040 ( .B1(n12854), .B2(n12821), .A(n12763), .ZN(n12764) );
  OAI21_X1 U15041 ( .B1(n12765), .B2(n15136), .A(n12764), .ZN(P3_U3213) );
  OAI211_X1 U15042 ( .C1(n12768), .C2(n12774), .A(n12767), .B(n12766), .ZN(
        n12772) );
  NAND2_X1 U15043 ( .A1(n12770), .A2(n12769), .ZN(n12771) );
  OAI211_X1 U15044 ( .C1(n12800), .C2(n12799), .A(n12772), .B(n12771), .ZN(
        n12857) );
  INV_X1 U15045 ( .A(n12857), .ZN(n12780) );
  XNOR2_X1 U15046 ( .A(n12773), .B(n12774), .ZN(n12858) );
  NOR2_X1 U15047 ( .A1(n12910), .A2(n12815), .ZN(n12778) );
  OAI22_X1 U15048 ( .A1(n12818), .A2(n12776), .B1(n12775), .B2(n12816), .ZN(
        n12777) );
  AOI211_X1 U15049 ( .C1(n12858), .C2(n12821), .A(n12778), .B(n12777), .ZN(
        n12779) );
  OAI21_X1 U15050 ( .B1(n12780), .B2(n15136), .A(n12779), .ZN(P3_U3214) );
  AOI21_X1 U15051 ( .B1(n12783), .B2(n12782), .A(n12781), .ZN(n12784) );
  OAI222_X1 U15052 ( .A1(n15122), .A2(n12785), .B1(n12799), .B2(n12812), .C1(
        n15128), .C2(n12784), .ZN(n12861) );
  INV_X1 U15053 ( .A(n12861), .ZN(n12795) );
  INV_X1 U15054 ( .A(n12786), .ZN(n12787) );
  AOI21_X1 U15055 ( .B1(n12789), .B2(n12788), .A(n12787), .ZN(n12862) );
  NOR2_X1 U15056 ( .A1(n12914), .A2(n12815), .ZN(n12793) );
  OAI22_X1 U15057 ( .A1(n12818), .A2(n12791), .B1(n12790), .B2(n12816), .ZN(
        n12792) );
  AOI211_X1 U15058 ( .C1(n12862), .C2(n12821), .A(n12793), .B(n12792), .ZN(
        n12794) );
  OAI21_X1 U15059 ( .B1(n12795), .B2(n15136), .A(n12794), .ZN(P3_U3215) );
  XNOR2_X1 U15060 ( .A(n12796), .B(n12801), .ZN(n12797) );
  OAI222_X1 U15061 ( .A1(n15122), .A2(n12800), .B1(n12799), .B2(n12798), .C1(
        n12797), .C2(n15128), .ZN(n12865) );
  INV_X1 U15062 ( .A(n12865), .ZN(n12807) );
  XNOR2_X1 U15063 ( .A(n12802), .B(n12801), .ZN(n12866) );
  NOR2_X1 U15064 ( .A1(n12918), .A2(n12815), .ZN(n12805) );
  OAI22_X1 U15065 ( .A1(n12818), .A2(n14448), .B1(n12803), .B2(n12816), .ZN(
        n12804) );
  AOI211_X1 U15066 ( .C1(n12866), .C2(n12821), .A(n12805), .B(n12804), .ZN(
        n12806) );
  OAI21_X1 U15067 ( .B1(n12807), .B2(n15136), .A(n12806), .ZN(P3_U3216) );
  XNOR2_X1 U15068 ( .A(n12809), .B(n12808), .ZN(n12810) );
  OAI222_X1 U15069 ( .A1(n15122), .A2(n12812), .B1(n12799), .B2(n12811), .C1(
        n12810), .C2(n15128), .ZN(n12869) );
  INV_X1 U15070 ( .A(n12869), .ZN(n12823) );
  OAI21_X1 U15071 ( .B1(n12814), .B2(n7434), .A(n12813), .ZN(n12870) );
  NOR2_X1 U15072 ( .A1(n12922), .A2(n12815), .ZN(n12820) );
  OAI22_X1 U15073 ( .A1(n12818), .A2(n12576), .B1(n12817), .B2(n12816), .ZN(
        n12819) );
  AOI211_X1 U15074 ( .C1(n12870), .C2(n12821), .A(n12820), .B(n12819), .ZN(
        n12822) );
  OAI21_X1 U15075 ( .B1(n12823), .B2(n15136), .A(n12822), .ZN(P3_U3217) );
  INV_X1 U15076 ( .A(n12878), .ZN(n12826) );
  NAND2_X1 U15077 ( .A1(n15164), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12825) );
  NAND2_X1 U15078 ( .A1(n14474), .A2(n15166), .ZN(n12824) );
  OAI211_X1 U15079 ( .C1(n12826), .C2(n12876), .A(n12825), .B(n12824), .ZN(
        P3_U3490) );
  INV_X1 U15080 ( .A(n12828), .ZN(n12829) );
  OAI21_X1 U15081 ( .B1(n12830), .B2(n12876), .A(n12829), .ZN(P3_U3486) );
  INV_X1 U15082 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12833) );
  AOI21_X1 U15083 ( .B1(n12832), .B2(n15150), .A(n12831), .ZN(n12881) );
  MUX2_X1 U15084 ( .A(n12833), .B(n12881), .S(n15166), .Z(n12834) );
  OAI21_X1 U15085 ( .B1(n12884), .B2(n12876), .A(n12834), .ZN(P3_U3485) );
  AOI21_X1 U15086 ( .B1(n15150), .B2(n12836), .A(n12835), .ZN(n12885) );
  MUX2_X1 U15087 ( .A(n14293), .B(n12885), .S(n15166), .Z(n12837) );
  OAI21_X1 U15088 ( .B1(n12888), .B2(n12876), .A(n12837), .ZN(P3_U3484) );
  INV_X1 U15089 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12840) );
  AOI21_X1 U15090 ( .B1(n15150), .B2(n12839), .A(n12838), .ZN(n12889) );
  MUX2_X1 U15091 ( .A(n12840), .B(n12889), .S(n15166), .Z(n12841) );
  OAI21_X1 U15092 ( .B1(n12892), .B2(n12876), .A(n12841), .ZN(P3_U3483) );
  INV_X1 U15093 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12844) );
  AOI21_X1 U15094 ( .B1(n15150), .B2(n12843), .A(n12842), .ZN(n12893) );
  MUX2_X1 U15095 ( .A(n12844), .B(n12893), .S(n15166), .Z(n12845) );
  OAI21_X1 U15096 ( .B1(n12895), .B2(n12876), .A(n12845), .ZN(P3_U3482) );
  INV_X1 U15097 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12848) );
  AOI21_X1 U15098 ( .B1(n15150), .B2(n12847), .A(n12846), .ZN(n12896) );
  MUX2_X1 U15099 ( .A(n12848), .B(n12896), .S(n15166), .Z(n12849) );
  OAI21_X1 U15100 ( .B1(n12898), .B2(n12876), .A(n12849), .ZN(P3_U3481) );
  AOI21_X1 U15101 ( .B1(n15150), .B2(n12851), .A(n12850), .ZN(n12899) );
  MUX2_X1 U15102 ( .A(n14237), .B(n12899), .S(n15166), .Z(n12852) );
  OAI21_X1 U15103 ( .B1(n12902), .B2(n12876), .A(n12852), .ZN(P3_U3480) );
  AOI21_X1 U15104 ( .B1(n12854), .B2(n15150), .A(n12853), .ZN(n12903) );
  MUX2_X1 U15105 ( .A(n12855), .B(n12903), .S(n15166), .Z(n12856) );
  OAI21_X1 U15106 ( .B1(n12906), .B2(n12876), .A(n12856), .ZN(P3_U3479) );
  AOI21_X1 U15107 ( .B1(n15150), .B2(n12858), .A(n12857), .ZN(n12907) );
  MUX2_X1 U15108 ( .A(n12859), .B(n12907), .S(n15166), .Z(n12860) );
  OAI21_X1 U15109 ( .B1(n12910), .B2(n12876), .A(n12860), .ZN(P3_U3478) );
  INV_X1 U15110 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12863) );
  AOI21_X1 U15111 ( .B1(n12862), .B2(n15150), .A(n12861), .ZN(n12911) );
  MUX2_X1 U15112 ( .A(n12863), .B(n12911), .S(n15166), .Z(n12864) );
  OAI21_X1 U15113 ( .B1(n12914), .B2(n12876), .A(n12864), .ZN(P3_U3477) );
  AOI21_X1 U15114 ( .B1(n12866), .B2(n15150), .A(n12865), .ZN(n12915) );
  MUX2_X1 U15115 ( .A(n12867), .B(n12915), .S(n15166), .Z(n12868) );
  OAI21_X1 U15116 ( .B1(n12876), .B2(n12918), .A(n12868), .ZN(P3_U3476) );
  AOI21_X1 U15117 ( .B1(n15150), .B2(n12870), .A(n12869), .ZN(n12919) );
  MUX2_X1 U15118 ( .A(n12871), .B(n12919), .S(n15166), .Z(n12872) );
  OAI21_X1 U15119 ( .B1(n12922), .B2(n12876), .A(n12872), .ZN(P3_U3475) );
  AOI21_X1 U15120 ( .B1(n12874), .B2(n15150), .A(n12873), .ZN(n12923) );
  MUX2_X1 U15121 ( .A(n14335), .B(n12923), .S(n15166), .Z(n12875) );
  OAI21_X1 U15122 ( .B1(n12876), .B2(n12925), .A(n12875), .ZN(P3_U3474) );
  INV_X1 U15123 ( .A(n12926), .ZN(n12877) );
  NAND2_X1 U15124 ( .A1(n12878), .A2(n12877), .ZN(n12880) );
  NAND2_X1 U15125 ( .A1(n14474), .A2(n15158), .ZN(n12879) );
  OAI211_X1 U15126 ( .C1(n12347), .C2(n15158), .A(n12880), .B(n12879), .ZN(
        P3_U3458) );
  INV_X1 U15127 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12882) );
  MUX2_X1 U15128 ( .A(n12882), .B(n12881), .S(n15158), .Z(n12883) );
  OAI21_X1 U15129 ( .B1(n12884), .B2(n12926), .A(n12883), .ZN(P3_U3453) );
  INV_X1 U15130 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12886) );
  MUX2_X1 U15131 ( .A(n12886), .B(n12885), .S(n15158), .Z(n12887) );
  OAI21_X1 U15132 ( .B1(n12888), .B2(n12926), .A(n12887), .ZN(P3_U3452) );
  INV_X1 U15133 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12890) );
  MUX2_X1 U15134 ( .A(n12890), .B(n12889), .S(n15158), .Z(n12891) );
  OAI21_X1 U15135 ( .B1(n12892), .B2(n12926), .A(n12891), .ZN(P3_U3451) );
  MUX2_X1 U15136 ( .A(n14266), .B(n12893), .S(n15158), .Z(n12894) );
  OAI21_X1 U15137 ( .B1(n12895), .B2(n12926), .A(n12894), .ZN(P3_U3450) );
  MUX2_X1 U15138 ( .A(n14334), .B(n12896), .S(n15158), .Z(n12897) );
  OAI21_X1 U15139 ( .B1(n12898), .B2(n12926), .A(n12897), .ZN(P3_U3449) );
  INV_X1 U15140 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12900) );
  MUX2_X1 U15141 ( .A(n12900), .B(n12899), .S(n15158), .Z(n12901) );
  OAI21_X1 U15142 ( .B1(n12902), .B2(n12926), .A(n12901), .ZN(P3_U3448) );
  MUX2_X1 U15143 ( .A(n12904), .B(n12903), .S(n15158), .Z(n12905) );
  OAI21_X1 U15144 ( .B1(n12906), .B2(n12926), .A(n12905), .ZN(P3_U3447) );
  INV_X1 U15145 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12908) );
  MUX2_X1 U15146 ( .A(n12908), .B(n12907), .S(n15158), .Z(n12909) );
  OAI21_X1 U15147 ( .B1(n12910), .B2(n12926), .A(n12909), .ZN(P3_U3446) );
  MUX2_X1 U15148 ( .A(n12912), .B(n12911), .S(n15158), .Z(n12913) );
  OAI21_X1 U15149 ( .B1(n12914), .B2(n12926), .A(n12913), .ZN(P3_U3444) );
  INV_X1 U15150 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12916) );
  MUX2_X1 U15151 ( .A(n12916), .B(n12915), .S(n15158), .Z(n12917) );
  OAI21_X1 U15152 ( .B1(n12926), .B2(n12918), .A(n12917), .ZN(P3_U3441) );
  INV_X1 U15153 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12920) );
  MUX2_X1 U15154 ( .A(n12920), .B(n12919), .S(n15158), .Z(n12921) );
  OAI21_X1 U15155 ( .B1(n12922), .B2(n12926), .A(n12921), .ZN(P3_U3438) );
  MUX2_X1 U15156 ( .A(n14244), .B(n12923), .S(n15158), .Z(n12924) );
  OAI21_X1 U15157 ( .B1(n12926), .B2(n12925), .A(n12924), .ZN(P3_U3435) );
  NAND2_X1 U15158 ( .A1(n12928), .A2(n12927), .ZN(n12932) );
  OR4_X1 U15159 ( .A1(n12930), .A2(P3_IR_REG_30__SCAN_IN), .A3(n12929), .A4(
        P3_U3151), .ZN(n12931) );
  OAI211_X1 U15160 ( .C1(n12934), .C2(n12933), .A(n12932), .B(n12931), .ZN(
        P3_U3264) );
  OAI222_X1 U15161 ( .A1(n12939), .A2(n12937), .B1(n11500), .B2(n12936), .C1(
        n12935), .C2(P3_U3151), .ZN(P3_U3266) );
  INV_X1 U15162 ( .A(n12938), .ZN(n12941) );
  XNOR2_X1 U15163 ( .A(n12942), .B(n12943), .ZN(n12947) );
  AOI22_X1 U15164 ( .A1(n13074), .A2(n13372), .B1(n13370), .B2(n13076), .ZN(
        n13261) );
  AOI22_X1 U15165 ( .A1(n13266), .A2(n13036), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12944) );
  OAI21_X1 U15166 ( .B1(n13261), .B2(n13066), .A(n12944), .ZN(n12945) );
  AOI21_X1 U15167 ( .B1(n13444), .B2(n14507), .A(n12945), .ZN(n12946) );
  OAI21_X1 U15168 ( .B1(n12947), .B2(n14502), .A(n12946), .ZN(P2_U3186) );
  NAND2_X1 U15169 ( .A1(n13040), .A2(n13338), .ZN(n12951) );
  OR2_X1 U15170 ( .A1(n12948), .A2(n14502), .ZN(n12950) );
  MUX2_X1 U15171 ( .A(n12951), .B(n12950), .S(n12949), .Z(n12955) );
  AOI22_X1 U15172 ( .A1(n13078), .A2(n13372), .B1(n13370), .B2(n13357), .ZN(
        n13331) );
  OAI22_X1 U15173 ( .A1(n13331), .A2(n13066), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12952), .ZN(n12953) );
  AOI21_X1 U15174 ( .B1(n13321), .B2(n13036), .A(n12953), .ZN(n12954) );
  OAI211_X1 U15175 ( .C1(n7140), .C2(n14515), .A(n12955), .B(n12954), .ZN(
        P2_U3188) );
  INV_X1 U15176 ( .A(n12956), .ZN(n12957) );
  AOI22_X1 U15177 ( .A1(n12979), .A2(n13088), .B1(n12957), .B2(n13036), .ZN(
        n12959) );
  OAI211_X1 U15178 ( .C1(n12960), .C2(n14518), .A(n12959), .B(n12958), .ZN(
        n12965) );
  AOI211_X1 U15179 ( .C1(n12963), .C2(n12962), .A(n14502), .B(n12961), .ZN(
        n12964) );
  AOI211_X1 U15180 ( .C1(n12966), .C2(n14507), .A(n12965), .B(n12964), .ZN(
        n12967) );
  INV_X1 U15181 ( .A(n12967), .ZN(P2_U3189) );
  OAI21_X1 U15182 ( .B1(n12978), .B2(n10031), .A(n12968), .ZN(n12969) );
  NAND2_X1 U15183 ( .A1(n12969), .A2(n14523), .ZN(n12983) );
  NOR2_X1 U15184 ( .A1(n14528), .A2(n12970), .ZN(n12974) );
  OAI21_X1 U15185 ( .B1(n14518), .B2(n12972), .A(n12971), .ZN(n12973) );
  AOI211_X1 U15186 ( .C1(n12975), .C2(n14507), .A(n12974), .B(n12973), .ZN(
        n12982) );
  NOR3_X1 U15187 ( .A1(n12978), .A2(n12977), .A3(n12976), .ZN(n12980) );
  OAI21_X1 U15188 ( .B1(n12980), .B2(n12979), .A(n13090), .ZN(n12981) );
  NAND3_X1 U15189 ( .A1(n12983), .A2(n12982), .A3(n12981), .ZN(P2_U3193) );
  XNOR2_X1 U15190 ( .A(n12985), .B(n12984), .ZN(n12993) );
  OAI22_X1 U15191 ( .A1(n14518), .A2(n12987), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12986), .ZN(n12991) );
  INV_X1 U15192 ( .A(n12988), .ZN(n13360) );
  OAI22_X1 U15193 ( .A1(n14519), .A2(n12989), .B1(n13360), .B2(n14528), .ZN(
        n12990) );
  AOI211_X1 U15194 ( .C1(n13477), .C2(n14507), .A(n12991), .B(n12990), .ZN(
        n12992) );
  OAI21_X1 U15195 ( .B1(n12993), .B2(n14502), .A(n12992), .ZN(P2_U3195) );
  XNOR2_X1 U15196 ( .A(n12995), .B(n12994), .ZN(n13000) );
  AOI22_X1 U15197 ( .A1(n13076), .A2(n13372), .B1(n13370), .B2(n13078), .ZN(
        n13293) );
  INV_X1 U15198 ( .A(n12996), .ZN(n13298) );
  AOI22_X1 U15199 ( .A1(n13298), .A2(n13036), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12997) );
  OAI21_X1 U15200 ( .B1(n13293), .B2(n13066), .A(n12997), .ZN(n12998) );
  AOI21_X1 U15201 ( .B1(n13456), .B2(n14507), .A(n12998), .ZN(n12999) );
  OAI21_X1 U15202 ( .B1(n13000), .B2(n14502), .A(n12999), .ZN(P2_U3197) );
  INV_X1 U15203 ( .A(n13001), .ZN(n13004) );
  AOI22_X1 U15204 ( .A1(n13054), .A2(n13002), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13003) );
  OAI21_X1 U15205 ( .B1(n13004), .B2(n14528), .A(n13003), .ZN(n13010) );
  INV_X1 U15206 ( .A(n14512), .ZN(n13008) );
  AOI22_X1 U15207 ( .A1(n13005), .A2(n14523), .B1(n13040), .B2(n13081), .ZN(
        n13007) );
  NOR3_X1 U15208 ( .A1(n13008), .A2(n13007), .A3(n13006), .ZN(n13009) );
  AOI211_X1 U15209 ( .C1(n13498), .C2(n14507), .A(n13010), .B(n13009), .ZN(
        n13011) );
  OAI21_X1 U15210 ( .B1(n13012), .B2(n14502), .A(n13011), .ZN(P2_U3200) );
  XNOR2_X1 U15211 ( .A(n13014), .B(n13013), .ZN(n13019) );
  AOI22_X1 U15212 ( .A1(n13077), .A2(n13372), .B1(n13370), .B2(n13338), .ZN(
        n13305) );
  INV_X1 U15213 ( .A(n13311), .ZN(n13015) );
  AOI22_X1 U15214 ( .A1(n13036), .A2(n13015), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13016) );
  OAI21_X1 U15215 ( .B1(n13305), .B2(n13066), .A(n13016), .ZN(n13017) );
  AOI21_X1 U15216 ( .B1(n13462), .B2(n14507), .A(n13017), .ZN(n13018) );
  OAI21_X1 U15217 ( .B1(n13019), .B2(n14502), .A(n13018), .ZN(P2_U3201) );
  NAND2_X1 U15218 ( .A1(n13021), .A2(n13020), .ZN(n13023) );
  XOR2_X1 U15219 ( .A(n13023), .B(n13022), .Z(n13028) );
  OAI22_X1 U15220 ( .A1(n14519), .A2(n13053), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13024), .ZN(n13026) );
  OAI22_X1 U15221 ( .A1(n14518), .A2(n13045), .B1(n14528), .B2(n13378), .ZN(
        n13025) );
  AOI211_X1 U15222 ( .C1(n13481), .C2(n14507), .A(n13026), .B(n13025), .ZN(
        n13027) );
  OAI21_X1 U15223 ( .B1(n13028), .B2(n14502), .A(n13027), .ZN(P2_U3205) );
  AOI21_X1 U15224 ( .B1(n13030), .B2(n13029), .A(n14502), .ZN(n13032) );
  NAND2_X1 U15225 ( .A1(n13032), .A2(n13031), .ZN(n13039) );
  INV_X1 U15226 ( .A(n13033), .ZN(n13037) );
  OAI22_X1 U15227 ( .A1(n13066), .A2(n13034), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14854), .ZN(n13035) );
  AOI21_X1 U15228 ( .B1(n13037), .B2(n13036), .A(n13035), .ZN(n13038) );
  OAI211_X1 U15229 ( .C1(n14530), .C2(n14515), .A(n13039), .B(n13038), .ZN(
        P2_U3206) );
  INV_X1 U15230 ( .A(n13472), .ZN(n13345) );
  NAND2_X1 U15231 ( .A1(n13040), .A2(n13357), .ZN(n13044) );
  OR2_X1 U15232 ( .A1(n13041), .A2(n14502), .ZN(n13043) );
  MUX2_X1 U15233 ( .A(n13044), .B(n13043), .S(n13042), .Z(n13050) );
  NOR2_X1 U15234 ( .A1(n14519), .A2(n13045), .ZN(n13048) );
  OAI22_X1 U15235 ( .A1(n13046), .A2(n14518), .B1(n13342), .B2(n14528), .ZN(
        n13047) );
  AOI211_X1 U15236 ( .C1(P2_REG3_REG_22__SCAN_IN), .C2(P2_U3088), .A(n13048), 
        .B(n13047), .ZN(n13049) );
  OAI211_X1 U15237 ( .C1(n13345), .C2(n14515), .A(n13050), .B(n13049), .ZN(
        P2_U3207) );
  OAI22_X1 U15238 ( .A1(n13053), .A2(n13052), .B1(n14517), .B2(n13051), .ZN(
        n13405) );
  NAND2_X1 U15239 ( .A1(n13054), .A2(n13405), .ZN(n13055) );
  NAND2_X1 U15240 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13208)
         );
  OAI211_X1 U15241 ( .C1(n14528), .C2(n13411), .A(n13055), .B(n13208), .ZN(
        n13060) );
  AOI211_X1 U15242 ( .C1(n13058), .C2(n13057), .A(n14502), .B(n13056), .ZN(
        n13059) );
  AOI211_X1 U15243 ( .C1(n13493), .C2(n14507), .A(n13060), .B(n13059), .ZN(
        n13061) );
  INV_X1 U15244 ( .A(n13061), .ZN(P2_U3210) );
  INV_X1 U15245 ( .A(n13062), .ZN(n13063) );
  AOI21_X1 U15246 ( .B1(n13065), .B2(n13064), .A(n13063), .ZN(n13071) );
  AOI22_X1 U15247 ( .A1(n13075), .A2(n13372), .B1(n13370), .B2(n13077), .ZN(
        n13278) );
  NOR2_X1 U15248 ( .A1(n13278), .A2(n13066), .ZN(n13069) );
  OAI22_X1 U15249 ( .A1(n13284), .A2(n14528), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13067), .ZN(n13068) );
  AOI211_X1 U15250 ( .C1(n13451), .C2(n14507), .A(n13069), .B(n13068), .ZN(
        n13070) );
  OAI21_X1 U15251 ( .B1(n13071), .B2(n14502), .A(n13070), .ZN(P2_U3212) );
  MUX2_X1 U15252 ( .A(n13231), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13096), .Z(
        P2_U3562) );
  MUX2_X1 U15253 ( .A(n13072), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13096), .Z(
        P2_U3561) );
  MUX2_X1 U15254 ( .A(n13073), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13096), .Z(
        P2_U3560) );
  MUX2_X1 U15255 ( .A(n13074), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13096), .Z(
        P2_U3559) );
  MUX2_X1 U15256 ( .A(n13075), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13096), .Z(
        P2_U3558) );
  MUX2_X1 U15257 ( .A(n13076), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13096), .Z(
        P2_U3557) );
  MUX2_X1 U15258 ( .A(n13077), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13096), .Z(
        P2_U3556) );
  MUX2_X1 U15259 ( .A(n13078), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13096), .Z(
        P2_U3555) );
  MUX2_X1 U15260 ( .A(n13338), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13096), .Z(
        P2_U3554) );
  MUX2_X1 U15261 ( .A(n13357), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13096), .Z(
        P2_U3553) );
  MUX2_X1 U15262 ( .A(n13373), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13096), .Z(
        P2_U3552) );
  MUX2_X1 U15263 ( .A(n13358), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13096), .Z(
        P2_U3551) );
  MUX2_X1 U15264 ( .A(n13371), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13096), .Z(
        P2_U3550) );
  MUX2_X1 U15265 ( .A(n13079), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13096), .Z(
        P2_U3549) );
  MUX2_X1 U15266 ( .A(n13080), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13096), .Z(
        P2_U3548) );
  MUX2_X1 U15267 ( .A(n13081), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13096), .Z(
        P2_U3547) );
  MUX2_X1 U15268 ( .A(n13082), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13096), .Z(
        P2_U3546) );
  MUX2_X1 U15269 ( .A(n13083), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13096), .Z(
        P2_U3545) );
  MUX2_X1 U15270 ( .A(n13084), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13096), .Z(
        P2_U3544) );
  MUX2_X1 U15271 ( .A(n13085), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13096), .Z(
        P2_U3543) );
  MUX2_X1 U15272 ( .A(n13086), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13096), .Z(
        P2_U3542) );
  MUX2_X1 U15273 ( .A(n13087), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13096), .Z(
        P2_U3541) );
  MUX2_X1 U15274 ( .A(n13088), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13096), .Z(
        P2_U3540) );
  MUX2_X1 U15275 ( .A(n13089), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13096), .Z(
        P2_U3539) );
  MUX2_X1 U15276 ( .A(n13090), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13096), .Z(
        P2_U3538) );
  MUX2_X1 U15277 ( .A(n13091), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13096), .Z(
        P2_U3537) );
  MUX2_X1 U15278 ( .A(n13092), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13096), .Z(
        P2_U3536) );
  MUX2_X1 U15279 ( .A(n13093), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13096), .Z(
        P2_U3535) );
  MUX2_X1 U15280 ( .A(n13094), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13096), .Z(
        P2_U3534) );
  MUX2_X1 U15281 ( .A(n13095), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13096), .Z(
        P2_U3533) );
  MUX2_X1 U15282 ( .A(n13097), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13096), .Z(
        P2_U3532) );
  AOI211_X1 U15283 ( .C1(n13100), .C2(n13099), .A(n13098), .B(n14856), .ZN(
        n13101) );
  INV_X1 U15284 ( .A(n13101), .ZN(n13114) );
  NOR2_X1 U15285 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13102), .ZN(n13103) );
  AOI21_X1 U15286 ( .B1(n14840), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n13103), .ZN(
        n13113) );
  INV_X1 U15287 ( .A(n13104), .ZN(n13109) );
  NAND3_X1 U15288 ( .A1(n13107), .A2(n13106), .A3(n13105), .ZN(n13108) );
  NAND3_X1 U15289 ( .A1(n13224), .A2(n13109), .A3(n13108), .ZN(n13112) );
  NAND2_X1 U15290 ( .A1(n14862), .A2(n13110), .ZN(n13111) );
  NAND4_X1 U15291 ( .A1(n13114), .A2(n13113), .A3(n13112), .A4(n13111), .ZN(
        P2_U3217) );
  AOI211_X1 U15292 ( .C1(n13117), .C2(n13116), .A(n14856), .B(n13115), .ZN(
        n13118) );
  INV_X1 U15293 ( .A(n13118), .ZN(n13129) );
  INV_X1 U15294 ( .A(n13119), .ZN(n13120) );
  AOI21_X1 U15295 ( .B1(n14840), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n13120), .ZN(
        n13128) );
  MUX2_X1 U15296 ( .A(n10265), .B(P2_REG2_REG_5__SCAN_IN), .S(n13125), .Z(
        n13123) );
  INV_X1 U15297 ( .A(n13121), .ZN(n13122) );
  NAND2_X1 U15298 ( .A1(n13123), .A2(n13122), .ZN(n13124) );
  OAI211_X1 U15299 ( .C1(n14847), .C2(n13124), .A(n13224), .B(n13139), .ZN(
        n13127) );
  NAND2_X1 U15300 ( .A1(n14862), .A2(n13125), .ZN(n13126) );
  NAND4_X1 U15301 ( .A1(n13129), .A2(n13128), .A3(n13127), .A4(n13126), .ZN(
        P2_U3219) );
  AOI211_X1 U15302 ( .C1(n13132), .C2(n13131), .A(n14856), .B(n13130), .ZN(
        n13133) );
  INV_X1 U15303 ( .A(n13133), .ZN(n13146) );
  INV_X1 U15304 ( .A(n13134), .ZN(n13135) );
  AOI21_X1 U15305 ( .B1(n14840), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n13135), .ZN(
        n13145) );
  INV_X1 U15306 ( .A(n13136), .ZN(n13141) );
  NAND3_X1 U15307 ( .A1(n13139), .A2(n13138), .A3(n13137), .ZN(n13140) );
  NAND3_X1 U15308 ( .A1(n13224), .A2(n13141), .A3(n13140), .ZN(n13144) );
  NAND2_X1 U15309 ( .A1(n14862), .A2(n13142), .ZN(n13143) );
  NAND4_X1 U15310 ( .A1(n13146), .A2(n13145), .A3(n13144), .A4(n13143), .ZN(
        P2_U3220) );
  NAND2_X1 U15311 ( .A1(n13149), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n13160) );
  OAI211_X1 U15312 ( .C1(n13149), .C2(P2_REG1_REG_15__SCAN_IN), .A(n13160), 
        .B(n13223), .ZN(n13159) );
  NOR2_X1 U15313 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13150), .ZN(n13152) );
  NOR2_X1 U15314 ( .A1(n13184), .A2(n13161), .ZN(n13151) );
  AOI211_X1 U15315 ( .C1(n14840), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n13152), 
        .B(n13151), .ZN(n13158) );
  INV_X1 U15316 ( .A(n13153), .ZN(n13154) );
  NOR2_X1 U15317 ( .A1(n13155), .A2(n13154), .ZN(n13167) );
  XNOR2_X1 U15318 ( .A(n13167), .B(n13161), .ZN(n13156) );
  NAND2_X1 U15319 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n13156), .ZN(n13169) );
  OAI211_X1 U15320 ( .C1(n13156), .C2(P2_REG2_REG_15__SCAN_IN), .A(n13224), 
        .B(n13169), .ZN(n13157) );
  NAND3_X1 U15321 ( .A1(n13159), .A2(n13158), .A3(n13157), .ZN(P2_U3229) );
  OAI21_X1 U15322 ( .B1(n13162), .B2(n13161), .A(n13160), .ZN(n13164) );
  XOR2_X1 U15323 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13172), .Z(n13163) );
  NAND2_X1 U15324 ( .A1(n13164), .A2(n13163), .ZN(n13179) );
  OAI211_X1 U15325 ( .C1(n13164), .C2(n13163), .A(n13179), .B(n13223), .ZN(
        n13178) );
  NAND2_X1 U15326 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n14525)
         );
  INV_X1 U15327 ( .A(n14525), .ZN(n13166) );
  NOR2_X1 U15328 ( .A1(n13184), .A2(n13189), .ZN(n13165) );
  AOI211_X1 U15329 ( .C1(n14840), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n13166), 
        .B(n13165), .ZN(n13177) );
  NAND2_X1 U15330 ( .A1(n13168), .A2(n13167), .ZN(n13170) );
  NAND2_X1 U15331 ( .A1(n13170), .A2(n13169), .ZN(n13175) );
  NAND2_X1 U15332 ( .A1(n13172), .A2(n13188), .ZN(n13171) );
  OAI21_X1 U15333 ( .B1(n13172), .B2(n13188), .A(n13171), .ZN(n13174) );
  NAND2_X1 U15334 ( .A1(n13189), .A2(n13188), .ZN(n13173) );
  OAI211_X1 U15335 ( .C1(n13189), .C2(n13188), .A(n13175), .B(n13173), .ZN(
        n13187) );
  OAI211_X1 U15336 ( .C1(n13175), .C2(n13174), .A(n13187), .B(n13224), .ZN(
        n13176) );
  NAND3_X1 U15337 ( .A1(n13178), .A2(n13177), .A3(n13176), .ZN(P2_U3230) );
  INV_X1 U15338 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n13180) );
  OAI21_X1 U15339 ( .B1(n13189), .B2(n13180), .A(n13179), .ZN(n13182) );
  XNOR2_X1 U15340 ( .A(n13198), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n13181) );
  OAI21_X1 U15341 ( .B1(n13182), .B2(n13181), .A(n13223), .ZN(n13196) );
  AND2_X1 U15342 ( .A1(n13182), .A2(n13181), .ZN(n13202) );
  AND2_X1 U15343 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13186) );
  NOR2_X1 U15344 ( .A1(n13184), .A2(n13198), .ZN(n13185) );
  AOI211_X1 U15345 ( .C1(n14840), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n13186), 
        .B(n13185), .ZN(n13195) );
  OAI21_X1 U15346 ( .B1(n13189), .B2(n13188), .A(n13187), .ZN(n13193) );
  NAND2_X1 U15347 ( .A1(n13198), .A2(n14345), .ZN(n13190) );
  OAI21_X1 U15348 ( .B1(n13198), .B2(n14345), .A(n13190), .ZN(n13191) );
  INV_X1 U15349 ( .A(n13191), .ZN(n13192) );
  NAND2_X1 U15350 ( .A1(n13192), .A2(n13193), .ZN(n13197) );
  OAI211_X1 U15351 ( .C1(n13193), .C2(n13192), .A(n13197), .B(n13224), .ZN(
        n13194) );
  OAI211_X1 U15352 ( .C1(n13196), .C2(n13202), .A(n13195), .B(n13194), .ZN(
        P2_U3231) );
  OAI21_X1 U15353 ( .B1(n13198), .B2(n14345), .A(n13197), .ZN(n13199) );
  NOR2_X1 U15354 ( .A1(n13199), .A2(n13211), .ZN(n13215) );
  AOI21_X1 U15355 ( .B1(n13211), .B2(n13199), .A(n13215), .ZN(n13200) );
  INV_X1 U15356 ( .A(n13200), .ZN(n13201) );
  NOR2_X1 U15357 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n13201), .ZN(n13216) );
  AOI21_X1 U15358 ( .B1(n13201), .B2(P2_REG2_REG_18__SCAN_IN), .A(n13216), 
        .ZN(n13214) );
  AOI21_X1 U15359 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n13203), .A(n13202), 
        .ZN(n13205) );
  NOR2_X1 U15360 ( .A1(n13205), .A2(n13204), .ZN(n13218) );
  AOI21_X1 U15361 ( .B1(n13205), .B2(n13204), .A(n13218), .ZN(n13207) );
  AND2_X1 U15362 ( .A1(n13207), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n13219) );
  INV_X1 U15363 ( .A(n13219), .ZN(n13206) );
  OAI211_X1 U15364 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n13207), .A(n13206), 
        .B(n13223), .ZN(n13213) );
  INV_X1 U15365 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n13209) );
  OAI21_X1 U15366 ( .B1(n14871), .B2(n13209), .A(n13208), .ZN(n13210) );
  AOI21_X1 U15367 ( .B1(n13211), .B2(n14862), .A(n13210), .ZN(n13212) );
  OAI211_X1 U15368 ( .C1(n13214), .C2(n14864), .A(n13213), .B(n13212), .ZN(
        P2_U3232) );
  NOR2_X1 U15369 ( .A1(n13216), .A2(n13215), .ZN(n13217) );
  XOR2_X1 U15370 ( .A(n13217), .B(P2_REG2_REG_19__SCAN_IN), .Z(n13225) );
  INV_X1 U15371 ( .A(n13225), .ZN(n13221) );
  NOR2_X1 U15372 ( .A1(n13219), .A2(n13218), .ZN(n13220) );
  XNOR2_X1 U15373 ( .A(n13220), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n13222) );
  AOI22_X1 U15374 ( .A1(n13225), .A2(n13224), .B1(n13223), .B2(n13222), .ZN(
        n13227) );
  XNOR2_X1 U15375 ( .A(n13236), .B(n13427), .ZN(n13229) );
  NAND2_X1 U15376 ( .A1(n13229), .A2(n13505), .ZN(n13428) );
  NOR2_X1 U15377 ( .A1(n13394), .A2(n13230), .ZN(n13233) );
  NAND2_X1 U15378 ( .A1(n13232), .A2(n13231), .ZN(n13430) );
  NOR2_X1 U15379 ( .A1(n13426), .A2(n13430), .ZN(n13239) );
  AOI211_X1 U15380 ( .C1(n13427), .C2(n13381), .A(n13233), .B(n13239), .ZN(
        n13234) );
  OAI21_X1 U15381 ( .B1(n13428), .B2(n13325), .A(n13234), .ZN(P2_U3234) );
  INV_X1 U15382 ( .A(n13235), .ZN(n13237) );
  INV_X1 U15383 ( .A(n13241), .ZN(n13432) );
  NOR2_X1 U15384 ( .A1(n13394), .A2(n13238), .ZN(n13240) );
  AOI211_X1 U15385 ( .C1(n13241), .C2(n13381), .A(n13240), .B(n13239), .ZN(
        n13242) );
  OAI21_X1 U15386 ( .B1(n13431), .B2(n13325), .A(n13242), .ZN(P2_U3235) );
  AOI211_X1 U15387 ( .C1(n13249), .C2(n13244), .A(n13294), .B(n13243), .ZN(
        n13247) );
  INV_X1 U15388 ( .A(n13245), .ZN(n13246) );
  NOR2_X1 U15389 ( .A1(n13247), .A2(n13246), .ZN(n13440) );
  OAI21_X1 U15390 ( .B1(n13250), .B2(n13249), .A(n13248), .ZN(n13441) );
  OAI22_X1 U15391 ( .A1(n13252), .A2(n13377), .B1(n13251), .B2(n13394), .ZN(
        n13253) );
  AOI21_X1 U15392 ( .B1(n13438), .B2(n13381), .A(n13253), .ZN(n13257) );
  AOI21_X1 U15393 ( .B1(n13264), .B2(n13438), .A(n13409), .ZN(n13255) );
  AND2_X1 U15394 ( .A1(n13255), .A2(n13254), .ZN(n13437) );
  NAND2_X1 U15395 ( .A1(n13437), .A2(n13424), .ZN(n13256) );
  OAI211_X1 U15396 ( .C1(n13441), .C2(n13421), .A(n13257), .B(n13256), .ZN(
        n13258) );
  INV_X1 U15397 ( .A(n13258), .ZN(n13259) );
  OAI21_X1 U15398 ( .B1(n13440), .B2(n13426), .A(n13259), .ZN(P2_U3237) );
  XNOR2_X1 U15399 ( .A(n13260), .B(n13270), .ZN(n13263) );
  INV_X1 U15400 ( .A(n13261), .ZN(n13262) );
  AOI21_X1 U15401 ( .B1(n13263), .B2(n13406), .A(n13262), .ZN(n13448) );
  OAI211_X1 U15402 ( .C1(n13280), .C2(n13265), .A(n13505), .B(n13264), .ZN(
        n13447) );
  AOI22_X1 U15403 ( .A1(n13266), .A2(n13412), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n13426), .ZN(n13268) );
  NAND2_X1 U15404 ( .A1(n13444), .A2(n13381), .ZN(n13267) );
  OAI211_X1 U15405 ( .C1(n13447), .C2(n13325), .A(n13268), .B(n13267), .ZN(
        n13269) );
  INV_X1 U15406 ( .A(n13269), .ZN(n13274) );
  OR2_X1 U15407 ( .A1(n13271), .A2(n13270), .ZN(n13443) );
  NAND3_X1 U15408 ( .A1(n13443), .A2(n13272), .A3(n13442), .ZN(n13273) );
  OAI211_X1 U15409 ( .C1(n13448), .C2(n13426), .A(n13274), .B(n13273), .ZN(
        P2_U3238) );
  XNOR2_X1 U15410 ( .A(n13275), .B(n13276), .ZN(n13453) );
  XNOR2_X1 U15411 ( .A(n13277), .B(n13276), .ZN(n13279) );
  OAI21_X1 U15412 ( .B1(n13279), .B2(n13294), .A(n13278), .ZN(n13449) );
  NAND2_X1 U15413 ( .A1(n13449), .A2(n13394), .ZN(n13288) );
  INV_X1 U15414 ( .A(n13296), .ZN(n13281) );
  AOI211_X1 U15415 ( .C1(n13451), .C2(n13281), .A(n13409), .B(n13280), .ZN(
        n13450) );
  NOR2_X1 U15416 ( .A1(n13282), .A2(n13415), .ZN(n13286) );
  OAI22_X1 U15417 ( .A1(n13284), .A2(n13377), .B1(n13283), .B2(n13394), .ZN(
        n13285) );
  AOI211_X1 U15418 ( .C1(n13450), .C2(n13424), .A(n13286), .B(n13285), .ZN(
        n13287) );
  OAI211_X1 U15419 ( .C1(n13453), .C2(n13421), .A(n13288), .B(n13287), .ZN(
        P2_U3239) );
  XNOR2_X1 U15420 ( .A(n13290), .B(n13289), .ZN(n13458) );
  XNOR2_X1 U15421 ( .A(n13292), .B(n13291), .ZN(n13295) );
  OAI21_X1 U15422 ( .B1(n13295), .B2(n13294), .A(n13293), .ZN(n13454) );
  NAND2_X1 U15423 ( .A1(n13454), .A2(n13394), .ZN(n13303) );
  INV_X1 U15424 ( .A(n13315), .ZN(n13297) );
  AOI211_X1 U15425 ( .C1(n13456), .C2(n13297), .A(n13409), .B(n13296), .ZN(
        n13455) );
  AOI22_X1 U15426 ( .A1(n13298), .A2(n13412), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n13426), .ZN(n13299) );
  OAI21_X1 U15427 ( .B1(n13300), .B2(n13415), .A(n13299), .ZN(n13301) );
  AOI21_X1 U15428 ( .B1(n13455), .B2(n13424), .A(n13301), .ZN(n13302) );
  OAI211_X1 U15429 ( .C1(n13458), .C2(n13421), .A(n13303), .B(n13302), .ZN(
        P2_U3240) );
  XNOR2_X1 U15430 ( .A(n13304), .B(n13308), .ZN(n13307) );
  INV_X1 U15431 ( .A(n13305), .ZN(n13306) );
  AOI21_X1 U15432 ( .B1(n13307), .B2(n13406), .A(n13306), .ZN(n13463) );
  OAI21_X1 U15433 ( .B1(n6475), .B2(n11553), .A(n13309), .ZN(n13459) );
  OAI22_X1 U15434 ( .A1(n13311), .A2(n13377), .B1(n13394), .B2(n13310), .ZN(
        n13312) );
  AOI21_X1 U15435 ( .B1(n13462), .B2(n13381), .A(n13312), .ZN(n13317) );
  NAND2_X1 U15436 ( .A1(n6502), .A2(n13462), .ZN(n13313) );
  NAND2_X1 U15437 ( .A1(n13313), .A2(n13505), .ZN(n13314) );
  NOR2_X1 U15438 ( .A1(n13315), .A2(n13314), .ZN(n13461) );
  NAND2_X1 U15439 ( .A1(n13461), .A2(n13424), .ZN(n13316) );
  OAI211_X1 U15440 ( .C1(n13459), .C2(n13421), .A(n13317), .B(n13316), .ZN(
        n13318) );
  INV_X1 U15441 ( .A(n13318), .ZN(n13319) );
  OAI21_X1 U15442 ( .B1(n13463), .B2(n13426), .A(n13319), .ZN(P2_U3241) );
  XNOR2_X1 U15443 ( .A(n13320), .B(n13328), .ZN(n13468) );
  INV_X1 U15444 ( .A(n13321), .ZN(n13323) );
  OAI22_X1 U15445 ( .A1(n13323), .A2(n13377), .B1(n13322), .B2(n13394), .ZN(
        n13327) );
  AOI21_X1 U15446 ( .B1(n13465), .B2(n13340), .A(n13409), .ZN(n13324) );
  NAND2_X1 U15447 ( .A1(n13324), .A2(n6502), .ZN(n13466) );
  NOR2_X1 U15448 ( .A1(n13466), .A2(n13325), .ZN(n13326) );
  AOI211_X1 U15449 ( .C1(n13381), .C2(n13465), .A(n13327), .B(n13326), .ZN(
        n13334) );
  XNOR2_X1 U15450 ( .A(n13329), .B(n13328), .ZN(n13330) );
  NAND2_X1 U15451 ( .A1(n13330), .A2(n13406), .ZN(n13332) );
  NAND2_X1 U15452 ( .A1(n13332), .A2(n13331), .ZN(n13470) );
  NAND2_X1 U15453 ( .A1(n13470), .A2(n13394), .ZN(n13333) );
  OAI211_X1 U15454 ( .C1(n13421), .C2(n13468), .A(n13334), .B(n13333), .ZN(
        P2_U3242) );
  INV_X1 U15455 ( .A(n13335), .ZN(n13337) );
  INV_X1 U15456 ( .A(n13347), .ZN(n13336) );
  OAI21_X1 U15457 ( .B1(n13337), .B2(n13336), .A(n6497), .ZN(n13339) );
  AOI222_X1 U15458 ( .A1(n13406), .A2(n13339), .B1(n13373), .B2(n13370), .C1(
        n13338), .C2(n13372), .ZN(n13474) );
  INV_X1 U15459 ( .A(n13340), .ZN(n13341) );
  AOI211_X1 U15460 ( .C1(n13472), .C2(n13363), .A(n13409), .B(n13341), .ZN(
        n13471) );
  INV_X1 U15461 ( .A(n13342), .ZN(n13343) );
  AOI22_X1 U15462 ( .A1(n13426), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n13343), 
        .B2(n13412), .ZN(n13344) );
  OAI21_X1 U15463 ( .B1(n13345), .B2(n13415), .A(n13344), .ZN(n13351) );
  OR2_X1 U15464 ( .A1(n13347), .A2(n13346), .ZN(n13348) );
  NAND2_X1 U15465 ( .A1(n13349), .A2(n13348), .ZN(n13475) );
  NOR2_X1 U15466 ( .A1(n13475), .A2(n13421), .ZN(n13350) );
  AOI211_X1 U15467 ( .C1(n13471), .C2(n13424), .A(n13351), .B(n13350), .ZN(
        n13352) );
  OAI21_X1 U15468 ( .B1(n13474), .B2(n13426), .A(n13352), .ZN(P2_U3243) );
  XNOR2_X1 U15469 ( .A(n13353), .B(n13355), .ZN(n13480) );
  OAI21_X1 U15470 ( .B1(n13356), .B2(n13355), .A(n13354), .ZN(n13359) );
  AOI222_X1 U15471 ( .A1(n13406), .A2(n13359), .B1(n13358), .B2(n13370), .C1(
        n13357), .C2(n13372), .ZN(n13479) );
  OAI22_X1 U15472 ( .A1(n13394), .A2(n13361), .B1(n13360), .B2(n13377), .ZN(
        n13362) );
  AOI21_X1 U15473 ( .B1(n13477), .B2(n13381), .A(n13362), .ZN(n13366) );
  AOI21_X1 U15474 ( .B1(n13384), .B2(n13477), .A(n13409), .ZN(n13364) );
  AND2_X1 U15475 ( .A1(n13364), .A2(n13363), .ZN(n13476) );
  NAND2_X1 U15476 ( .A1(n13476), .A2(n13424), .ZN(n13365) );
  OAI211_X1 U15477 ( .C1(n13479), .C2(n13426), .A(n13366), .B(n13365), .ZN(
        n13367) );
  INV_X1 U15478 ( .A(n13367), .ZN(n13368) );
  OAI21_X1 U15479 ( .B1(n13480), .B2(n13421), .A(n13368), .ZN(P2_U3244) );
  XOR2_X1 U15480 ( .A(n13369), .B(n13376), .Z(n13374) );
  AOI222_X1 U15481 ( .A1(n13406), .A2(n13374), .B1(n13373), .B2(n13372), .C1(
        n13371), .C2(n13370), .ZN(n13484) );
  XNOR2_X1 U15482 ( .A(n13375), .B(n13376), .ZN(n13485) );
  OAI22_X1 U15483 ( .A1(n13394), .A2(n13379), .B1(n13378), .B2(n13377), .ZN(
        n13380) );
  AOI21_X1 U15484 ( .B1(n13481), .B2(n13381), .A(n13380), .ZN(n13387) );
  OR2_X1 U15485 ( .A1(n13382), .A2(n13396), .ZN(n13383) );
  AND2_X1 U15486 ( .A1(n13384), .A2(n13383), .ZN(n13482) );
  NAND2_X1 U15487 ( .A1(n13482), .A2(n13385), .ZN(n13386) );
  OAI211_X1 U15488 ( .C1(n13485), .C2(n13421), .A(n13387), .B(n13386), .ZN(
        n13388) );
  INV_X1 U15489 ( .A(n13388), .ZN(n13389) );
  OAI21_X1 U15490 ( .B1(n13484), .B2(n13426), .A(n13389), .ZN(P2_U3245) );
  XOR2_X1 U15491 ( .A(n13390), .B(n13392), .Z(n13491) );
  XOR2_X1 U15492 ( .A(n13392), .B(n13391), .Z(n13393) );
  NAND2_X1 U15493 ( .A1(n13393), .A2(n13406), .ZN(n13489) );
  INV_X1 U15494 ( .A(n13489), .ZN(n13395) );
  OAI21_X1 U15495 ( .B1(n13395), .B2(n13487), .A(n13394), .ZN(n13402) );
  AOI211_X1 U15496 ( .C1(n13488), .C2(n13408), .A(n13409), .B(n13396), .ZN(
        n13486) );
  INV_X1 U15497 ( .A(n13488), .ZN(n13399) );
  AOI22_X1 U15498 ( .A1(n13426), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13397), 
        .B2(n13412), .ZN(n13398) );
  OAI21_X1 U15499 ( .B1(n13399), .B2(n13415), .A(n13398), .ZN(n13400) );
  AOI21_X1 U15500 ( .B1(n13486), .B2(n13424), .A(n13400), .ZN(n13401) );
  OAI211_X1 U15501 ( .C1(n13491), .C2(n13421), .A(n13402), .B(n13401), .ZN(
        P2_U3246) );
  XNOR2_X1 U15502 ( .A(n13404), .B(n13403), .ZN(n13407) );
  AOI21_X1 U15503 ( .B1(n13407), .B2(n13406), .A(n13405), .ZN(n13495) );
  AOI211_X1 U15504 ( .C1(n13493), .C2(n13410), .A(n13409), .B(n7132), .ZN(
        n13492) );
  INV_X1 U15505 ( .A(n13493), .ZN(n13416) );
  INV_X1 U15506 ( .A(n13411), .ZN(n13413) );
  AOI22_X1 U15507 ( .A1(n13426), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13413), 
        .B2(n13412), .ZN(n13414) );
  OAI21_X1 U15508 ( .B1(n13416), .B2(n13415), .A(n13414), .ZN(n13423) );
  INV_X1 U15509 ( .A(n13417), .ZN(n13418) );
  AOI21_X1 U15510 ( .B1(n13420), .B2(n13419), .A(n13418), .ZN(n13496) );
  NOR2_X1 U15511 ( .A1(n13496), .A2(n13421), .ZN(n13422) );
  AOI211_X1 U15512 ( .C1(n13492), .C2(n13424), .A(n13423), .B(n13422), .ZN(
        n13425) );
  OAI21_X1 U15513 ( .B1(n13426), .B2(n13495), .A(n13425), .ZN(P2_U3247) );
  INV_X1 U15514 ( .A(n13427), .ZN(n13429) );
  OAI211_X1 U15515 ( .C1(n13429), .C2(n14922), .A(n13428), .B(n13430), .ZN(
        n13522) );
  MUX2_X1 U15516 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13522), .S(n14933), .Z(
        P2_U3530) );
  OAI211_X1 U15517 ( .C1(n13432), .C2(n14922), .A(n13431), .B(n13430), .ZN(
        n13523) );
  MUX2_X1 U15518 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13523), .S(n14933), .Z(
        P2_U3529) );
  AOI21_X1 U15519 ( .B1(n13513), .B2(n13438), .A(n13437), .ZN(n13439) );
  OAI211_X1 U15520 ( .C1(n13516), .C2(n13441), .A(n13440), .B(n13439), .ZN(
        n13524) );
  MUX2_X1 U15521 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13524), .S(n14933), .Z(
        P2_U3527) );
  NAND3_X1 U15522 ( .A1(n13443), .A2(n13442), .A3(n14533), .ZN(n13446) );
  NAND2_X1 U15523 ( .A1(n13444), .A2(n13513), .ZN(n13445) );
  NAND4_X1 U15524 ( .A1(n13448), .A2(n13447), .A3(n13446), .A4(n13445), .ZN(
        n13525) );
  MUX2_X1 U15525 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13525), .S(n14933), .Z(
        P2_U3526) );
  OAI21_X1 U15526 ( .B1(n13516), .B2(n13453), .A(n13452), .ZN(n13526) );
  MUX2_X1 U15527 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13526), .S(n14933), .Z(
        P2_U3525) );
  AOI211_X1 U15528 ( .C1(n13513), .C2(n13456), .A(n13455), .B(n13454), .ZN(
        n13457) );
  OAI21_X1 U15529 ( .B1(n13516), .B2(n13458), .A(n13457), .ZN(n13527) );
  MUX2_X1 U15530 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13527), .S(n14933), .Z(
        P2_U3524) );
  NOR2_X1 U15531 ( .A1(n13459), .A2(n13516), .ZN(n13460) );
  AOI211_X1 U15532 ( .C1(n13513), .C2(n13462), .A(n13461), .B(n13460), .ZN(
        n13464) );
  NAND2_X1 U15533 ( .A1(n13464), .A2(n13463), .ZN(n13528) );
  MUX2_X1 U15534 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13528), .S(n14933), .Z(
        P2_U3523) );
  NAND2_X1 U15535 ( .A1(n13465), .A2(n13513), .ZN(n13467) );
  OAI211_X1 U15536 ( .C1(n13468), .C2(n13516), .A(n13467), .B(n13466), .ZN(
        n13469) );
  MUX2_X1 U15537 ( .A(n13529), .B(P2_REG1_REG_23__SCAN_IN), .S(n14931), .Z(
        P2_U3522) );
  AOI21_X1 U15538 ( .B1(n13513), .B2(n13472), .A(n13471), .ZN(n13473) );
  OAI211_X1 U15539 ( .C1(n13516), .C2(n13475), .A(n13474), .B(n13473), .ZN(
        n13530) );
  MUX2_X1 U15540 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13530), .S(n14933), .Z(
        P2_U3521) );
  AOI21_X1 U15541 ( .B1(n13513), .B2(n13477), .A(n13476), .ZN(n13478) );
  OAI211_X1 U15542 ( .C1(n13516), .C2(n13480), .A(n13479), .B(n13478), .ZN(
        n13531) );
  MUX2_X1 U15543 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13531), .S(n14933), .Z(
        P2_U3520) );
  AOI22_X1 U15544 ( .A1(n13482), .A2(n13505), .B1(n13513), .B2(n13481), .ZN(
        n13483) );
  OAI211_X1 U15545 ( .C1(n13516), .C2(n13485), .A(n13484), .B(n13483), .ZN(
        n13532) );
  MUX2_X1 U15546 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13532), .S(n14933), .Z(
        P2_U3519) );
  AOI211_X1 U15547 ( .C1(n13513), .C2(n13488), .A(n13487), .B(n13486), .ZN(
        n13490) );
  OAI211_X1 U15548 ( .C1(n13516), .C2(n13491), .A(n13490), .B(n13489), .ZN(
        n13533) );
  MUX2_X1 U15549 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13533), .S(n14933), .Z(
        P2_U3518) );
  AOI21_X1 U15550 ( .B1(n13513), .B2(n13493), .A(n13492), .ZN(n13494) );
  OAI211_X1 U15551 ( .C1(n13496), .C2(n13516), .A(n13495), .B(n13494), .ZN(
        n13534) );
  MUX2_X1 U15552 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13534), .S(n14933), .Z(
        P2_U3517) );
  AOI21_X1 U15553 ( .B1(n13513), .B2(n13498), .A(n13497), .ZN(n13499) );
  OAI211_X1 U15554 ( .C1(n13501), .C2(n13516), .A(n13500), .B(n13499), .ZN(
        n13535) );
  MUX2_X1 U15555 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13535), .S(n14933), .Z(
        P2_U3516) );
  NAND3_X1 U15556 ( .A1(n13503), .A2(n13502), .A3(n14533), .ZN(n13508) );
  AOI22_X1 U15557 ( .A1(n13506), .A2(n13505), .B1(n13513), .B2(n13504), .ZN(
        n13507) );
  NAND2_X1 U15558 ( .A1(n13508), .A2(n13507), .ZN(n13509) );
  MUX2_X1 U15559 ( .A(n13536), .B(P2_REG1_REG_16__SCAN_IN), .S(n14931), .Z(
        P2_U3515) );
  AOI211_X1 U15560 ( .C1(n13513), .C2(n14508), .A(n13512), .B(n13511), .ZN(
        n13514) );
  OAI21_X1 U15561 ( .B1(n13516), .B2(n13515), .A(n13514), .ZN(n13537) );
  MUX2_X1 U15562 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13537), .S(n14933), .Z(
        P2_U3513) );
  MUX2_X1 U15563 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n13517), .S(n14933), .Z(
        P2_U3510) );
  MUX2_X1 U15564 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n13518), .S(n14933), .Z(
        P2_U3508) );
  MUX2_X1 U15565 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n13519), .S(n14933), .Z(
        P2_U3505) );
  MUX2_X1 U15566 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n13520), .S(n14933), .Z(
        P2_U3504) );
  MUX2_X1 U15567 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n13521), .S(n14933), .Z(
        P2_U3502) );
  MUX2_X1 U15568 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13522), .S(n6443), .Z(
        P2_U3498) );
  MUX2_X1 U15569 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13523), .S(n6443), .Z(
        P2_U3497) );
  MUX2_X1 U15570 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13524), .S(n6443), .Z(
        P2_U3495) );
  MUX2_X1 U15571 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13525), .S(n6443), .Z(
        P2_U3494) );
  MUX2_X1 U15572 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13526), .S(n6443), .Z(
        P2_U3493) );
  MUX2_X1 U15573 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13527), .S(n6443), .Z(
        P2_U3492) );
  MUX2_X1 U15574 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13528), .S(n6443), .Z(
        P2_U3491) );
  MUX2_X1 U15575 ( .A(n13529), .B(P2_REG0_REG_23__SCAN_IN), .S(n14928), .Z(
        P2_U3490) );
  MUX2_X1 U15576 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13530), .S(n6443), .Z(
        P2_U3489) );
  MUX2_X1 U15577 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13531), .S(n6443), .Z(
        P2_U3488) );
  MUX2_X1 U15578 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13532), .S(n6443), .Z(
        P2_U3487) );
  MUX2_X1 U15579 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13533), .S(n6443), .Z(
        P2_U3486) );
  MUX2_X1 U15580 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13534), .S(n6443), .Z(
        P2_U3484) );
  MUX2_X1 U15581 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13535), .S(n6443), .Z(
        P2_U3481) );
  MUX2_X1 U15582 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13536), .S(n6443), .Z(
        P2_U3478) );
  MUX2_X1 U15583 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n13537), .S(n6443), .Z(
        P2_U3472) );
  INV_X1 U15584 ( .A(n14222), .ZN(n13543) );
  NOR4_X1 U15585 ( .A1(n13539), .A2(P2_IR_REG_30__SCAN_IN), .A3(n13538), .A4(
        P2_U3088), .ZN(n13540) );
  AOI21_X1 U15586 ( .B1(n13541), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13540), 
        .ZN(n13542) );
  OAI21_X1 U15587 ( .B1(n13543), .B2(n13549), .A(n13542), .ZN(P2_U3296) );
  INV_X1 U15588 ( .A(n13544), .ZN(n14371) );
  OAI222_X1 U15589 ( .A1(n13549), .A2(n14371), .B1(P2_U3088), .B2(n13546), 
        .C1(n13545), .C2(n13551), .ZN(P2_U3298) );
  INV_X1 U15590 ( .A(n13547), .ZN(n14374) );
  OAI222_X1 U15591 ( .A1(n13551), .A2(n13550), .B1(n13549), .B2(n14374), .C1(
        P2_U3088), .C2(n6698), .ZN(P2_U3300) );
  INV_X1 U15592 ( .A(n13552), .ZN(n13553) );
  MUX2_X1 U15593 ( .A(n13553), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XOR2_X1 U15594 ( .A(n13555), .B(n13554), .Z(n13561) );
  OAI22_X1 U15595 ( .A1(n13679), .A2(n13906), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13556), .ZN(n13557) );
  AOI21_X1 U15596 ( .B1(n6433), .B2(n14105), .A(n13557), .ZN(n13558) );
  OAI21_X1 U15597 ( .B1(n13900), .B2(n13667), .A(n13558), .ZN(n13559) );
  AOI21_X1 U15598 ( .B1(n14121), .B2(n13685), .A(n13559), .ZN(n13560) );
  OAI21_X1 U15599 ( .B1(n13561), .B2(n13688), .A(n13560), .ZN(P1_U3214) );
  AOI21_X1 U15600 ( .B1(n13563), .B2(n13562), .A(n13671), .ZN(n13568) );
  NAND2_X1 U15601 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14625)
         );
  OAI21_X1 U15602 ( .B1(n13679), .B2(n14080), .A(n14625), .ZN(n13564) );
  AOI21_X1 U15603 ( .B1(n13681), .B2(n14086), .A(n13564), .ZN(n13565) );
  OAI21_X1 U15604 ( .B1(n14085), .B2(n13683), .A(n13565), .ZN(n13566) );
  AOI21_X1 U15605 ( .B1(n14194), .B2(n13685), .A(n13566), .ZN(n13567) );
  OAI21_X1 U15606 ( .B1(n13568), .B2(n13688), .A(n13567), .ZN(P1_U3215) );
  XOR2_X1 U15607 ( .A(n13569), .B(n13570), .Z(n13576) );
  INV_X1 U15608 ( .A(n13995), .ZN(n13851) );
  NAND2_X1 U15609 ( .A1(n6433), .A2(n14132), .ZN(n13573) );
  INV_X1 U15610 ( .A(n13571), .ZN(n13970) );
  AOI22_X1 U15611 ( .A1(n13664), .A2(n13970), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13572) );
  OAI211_X1 U15612 ( .C1(n13851), .C2(n13667), .A(n13573), .B(n13572), .ZN(
        n13574) );
  AOI21_X1 U15613 ( .B1(n14144), .B2(n13685), .A(n13574), .ZN(n13575) );
  OAI21_X1 U15614 ( .B1(n13576), .B2(n13688), .A(n13575), .ZN(P1_U3216) );
  AOI21_X1 U15615 ( .B1(n13578), .B2(n13577), .A(n13688), .ZN(n13580) );
  NAND2_X1 U15616 ( .A1(n13580), .A2(n13579), .ZN(n13585) );
  OAI22_X1 U15617 ( .A1(n14723), .A2(n14720), .B1(n13581), .B2(n14722), .ZN(
        n14748) );
  AOI22_X1 U15618 ( .A1(n14748), .A2(n13582), .B1(n13685), .B2(n14753), .ZN(
        n13584) );
  MUX2_X1 U15619 ( .A(n13679), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n13583) );
  NAND3_X1 U15620 ( .A1(n13585), .A2(n13584), .A3(n13583), .ZN(P1_U3218) );
  OAI211_X1 U15621 ( .C1(n13588), .C2(n13587), .A(n13586), .B(n13645), .ZN(
        n13592) );
  NAND2_X1 U15622 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13798)
         );
  OAI21_X1 U15623 ( .B1(n13679), .B2(n14032), .A(n13798), .ZN(n13590) );
  NOR2_X1 U15624 ( .A1(n14166), .A2(n13667), .ZN(n13589) );
  AOI211_X1 U15625 ( .C1(n6433), .C2(n13996), .A(n13590), .B(n13589), .ZN(
        n13591) );
  OAI211_X1 U15626 ( .C1(n13848), .C2(n13652), .A(n13592), .B(n13591), .ZN(
        P1_U3219) );
  INV_X1 U15627 ( .A(n13593), .ZN(n13594) );
  AOI21_X1 U15628 ( .B1(n13596), .B2(n13595), .A(n13594), .ZN(n13602) );
  INV_X1 U15629 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13597) );
  OAI22_X1 U15630 ( .A1(n14002), .A2(n13679), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13597), .ZN(n13598) );
  AOI21_X1 U15631 ( .B1(n6433), .B2(n13995), .A(n13598), .ZN(n13599) );
  OAI21_X1 U15632 ( .B1(n14040), .B2(n13667), .A(n13599), .ZN(n13600) );
  AOI21_X1 U15633 ( .B1(n14154), .B2(n13685), .A(n13600), .ZN(n13601) );
  OAI21_X1 U15634 ( .B1(n13602), .B2(n13688), .A(n13601), .ZN(P1_U3223) );
  XOR2_X1 U15635 ( .A(n13604), .B(n13603), .Z(n13610) );
  INV_X1 U15636 ( .A(n14132), .ZN(n13945) );
  NAND2_X1 U15637 ( .A1(n6433), .A2(n13933), .ZN(n13607) );
  INV_X1 U15638 ( .A(n13942), .ZN(n13605) );
  AOI22_X1 U15639 ( .A1(n13664), .A2(n13605), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13606) );
  OAI211_X1 U15640 ( .C1(n13945), .C2(n13667), .A(n13607), .B(n13606), .ZN(
        n13608) );
  AOI21_X1 U15641 ( .B1(n14133), .B2(n13685), .A(n13608), .ZN(n13609) );
  OAI21_X1 U15642 ( .B1(n13610), .B2(n13688), .A(n13609), .ZN(P1_U3225) );
  AOI21_X1 U15643 ( .B1(n13612), .B2(n13611), .A(n6581), .ZN(n13618) );
  NAND2_X1 U15644 ( .A1(n13681), .A2(n13690), .ZN(n13613) );
  NAND2_X1 U15645 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14650)
         );
  OAI211_X1 U15646 ( .C1(n13679), .C2(n13614), .A(n13613), .B(n14650), .ZN(
        n13616) );
  NAND2_X1 U15647 ( .A1(n13843), .A2(n14792), .ZN(n14184) );
  NOR2_X1 U15648 ( .A1(n14184), .A2(n13621), .ZN(n13615) );
  AOI211_X1 U15649 ( .C1(n6433), .C2(n13844), .A(n13616), .B(n13615), .ZN(
        n13617) );
  OAI21_X1 U15650 ( .B1(n13618), .B2(n13688), .A(n13617), .ZN(P1_U3226) );
  XOR2_X1 U15651 ( .A(n13619), .B(n6487), .Z(n13625) );
  NAND2_X1 U15652 ( .A1(n13664), .A2(n14069), .ZN(n13620) );
  NAND2_X1 U15653 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14662)
         );
  OAI211_X1 U15654 ( .C1(n13683), .C2(n14166), .A(n13620), .B(n14662), .ZN(
        n13623) );
  NAND2_X1 U15655 ( .A1(n14070), .A2(n14792), .ZN(n14178) );
  NOR2_X1 U15656 ( .A1(n14178), .A2(n13621), .ZN(n13622) );
  AOI211_X1 U15657 ( .C1(n13681), .C2(n14064), .A(n13623), .B(n13622), .ZN(
        n13624) );
  OAI21_X1 U15658 ( .B1(n13625), .B2(n13688), .A(n13624), .ZN(P1_U3228) );
  XOR2_X1 U15659 ( .A(n13627), .B(n13626), .Z(n13633) );
  NAND2_X1 U15660 ( .A1(n6433), .A2(n13924), .ZN(n13630) );
  INV_X1 U15661 ( .A(n13628), .ZN(n13955) );
  AOI22_X1 U15662 ( .A1(n13664), .A2(n13955), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13629) );
  OAI211_X1 U15663 ( .C1(n13961), .C2(n13667), .A(n13630), .B(n13629), .ZN(
        n13631) );
  AOI21_X1 U15664 ( .B1(n14139), .B2(n13685), .A(n13631), .ZN(n13632) );
  OAI21_X1 U15665 ( .B1(n13633), .B2(n13688), .A(n13632), .ZN(P1_U3229) );
  OAI211_X1 U15666 ( .C1(n13636), .C2(n13635), .A(n13634), .B(n13645), .ZN(
        n13641) );
  OAI22_X1 U15667 ( .A1(n14018), .A2(n13679), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13637), .ZN(n13639) );
  NOR2_X1 U15668 ( .A1(n14054), .A2(n13667), .ZN(n13638) );
  AOI211_X1 U15669 ( .C1(n6433), .C2(n14017), .A(n13639), .B(n13638), .ZN(
        n13640) );
  OAI211_X1 U15670 ( .C1(n14161), .C2(n13652), .A(n13641), .B(n13640), .ZN(
        P1_U3233) );
  OAI21_X1 U15671 ( .B1(n13644), .B2(n13643), .A(n13642), .ZN(n13646) );
  NAND2_X1 U15672 ( .A1(n13646), .A2(n13645), .ZN(n13651) );
  OAI22_X1 U15673 ( .A1(n13679), .A2(n13984), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13647), .ZN(n13649) );
  NOR2_X1 U15674 ( .A1(n13823), .A2(n13667), .ZN(n13648) );
  AOI211_X1 U15675 ( .C1(n6433), .C2(n13980), .A(n13649), .B(n13648), .ZN(
        n13650) );
  OAI211_X1 U15676 ( .C1(n13652), .C2(n13852), .A(n13651), .B(n13650), .ZN(
        P1_U3235) );
  XOR2_X1 U15677 ( .A(n13654), .B(n13653), .Z(n13659) );
  NAND2_X1 U15678 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14677)
         );
  OAI21_X1 U15679 ( .B1(n13679), .B2(n14055), .A(n14677), .ZN(n13655) );
  AOI21_X1 U15680 ( .B1(n14016), .B2(n6433), .A(n13655), .ZN(n13656) );
  OAI21_X1 U15681 ( .B1(n14052), .B2(n13667), .A(n13656), .ZN(n13657) );
  AOI21_X1 U15682 ( .B1(n14174), .B2(n13685), .A(n13657), .ZN(n13658) );
  OAI21_X1 U15683 ( .B1(n13659), .B2(n13688), .A(n13658), .ZN(P1_U3238) );
  XOR2_X1 U15684 ( .A(n13661), .B(n13660), .Z(n13670) );
  NAND2_X1 U15685 ( .A1(n6433), .A2(n13925), .ZN(n13666) );
  INV_X1 U15686 ( .A(n13913), .ZN(n13663) );
  AOI22_X1 U15687 ( .A1(n13664), .A2(n13663), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13665) );
  OAI211_X1 U15688 ( .C1(n13960), .C2(n13667), .A(n13666), .B(n13665), .ZN(
        n13668) );
  AOI21_X1 U15689 ( .B1(n14126), .B2(n13685), .A(n13668), .ZN(n13669) );
  OAI21_X1 U15690 ( .B1(n13670), .B2(n13688), .A(n13669), .ZN(P1_U3240) );
  INV_X1 U15691 ( .A(n13671), .ZN(n13673) );
  NAND2_X1 U15692 ( .A1(n13673), .A2(n13672), .ZN(n13677) );
  XNOR2_X1 U15693 ( .A(n13675), .B(n13674), .ZN(n13676) );
  XNOR2_X1 U15694 ( .A(n13677), .B(n13676), .ZN(n13689) );
  NAND2_X1 U15695 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14638)
         );
  OAI21_X1 U15696 ( .B1(n13679), .B2(n13678), .A(n14638), .ZN(n13680) );
  AOI21_X1 U15697 ( .B1(n13681), .B2(n13691), .A(n13680), .ZN(n13682) );
  OAI21_X1 U15698 ( .B1(n13840), .B2(n13683), .A(n13682), .ZN(n13684) );
  AOI21_X1 U15699 ( .B1(n13686), .B2(n13685), .A(n13684), .ZN(n13687) );
  OAI21_X1 U15700 ( .B1(n13689), .B2(n13688), .A(n13687), .ZN(P1_U3241) );
  MUX2_X1 U15701 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13804), .S(n13701), .Z(
        P1_U3591) );
  MUX2_X1 U15702 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13868), .S(n13701), .Z(
        P1_U3590) );
  MUX2_X1 U15703 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13879), .S(n13701), .Z(
        P1_U3589) );
  MUX2_X1 U15704 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14105), .S(n13701), .Z(
        P1_U3588) );
  MUX2_X1 U15705 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13925), .S(n13701), .Z(
        P1_U3587) );
  MUX2_X1 U15706 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13933), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15707 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13924), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15708 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14132), .S(n13701), .Z(
        P1_U3584) );
  MUX2_X1 U15709 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13980), .S(n13701), .Z(
        P1_U3583) );
  MUX2_X1 U15710 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13995), .S(n13701), .Z(
        P1_U3582) );
  MUX2_X1 U15711 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14017), .S(n13701), .Z(
        P1_U3581) );
  MUX2_X1 U15712 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13996), .S(n13701), .Z(
        P1_U3580) );
  MUX2_X1 U15713 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14016), .S(n13701), .Z(
        P1_U3579) );
  MUX2_X1 U15714 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14065), .S(n13701), .Z(
        P1_U3578) );
  MUX2_X1 U15715 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n13844), .S(n13701), .Z(
        P1_U3577) );
  MUX2_X1 U15716 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14064), .S(n13701), .Z(
        P1_U3576) );
  MUX2_X1 U15717 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13690), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15718 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13691), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15719 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14086), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U15720 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13692), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U15721 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13693), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U15722 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13694), .S(n13701), .Z(
        P1_U3570) );
  MUX2_X1 U15723 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14683), .S(n13701), .Z(
        P1_U3569) );
  MUX2_X1 U15724 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14703), .S(n13701), .Z(
        P1_U3568) );
  MUX2_X1 U15725 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14682), .S(n13701), .Z(
        P1_U3567) );
  MUX2_X1 U15726 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14704), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U15727 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13696), .S(n13701), .Z(
        P1_U3565) );
  MUX2_X1 U15728 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13697), .S(n13701), .Z(
        P1_U3564) );
  MUX2_X1 U15729 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13698), .S(n13701), .Z(
        P1_U3563) );
  MUX2_X1 U15730 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13699), .S(n13701), .Z(
        P1_U3562) );
  MUX2_X1 U15731 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n13700), .S(n13701), .Z(
        P1_U3561) );
  MUX2_X1 U15732 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n13702), .S(n13701), .Z(
        P1_U3560) );
  NAND2_X1 U15733 ( .A1(n14377), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n13705) );
  AOI211_X1 U15734 ( .C1(n13705), .C2(n13704), .A(n13703), .B(n14665), .ZN(
        n13706) );
  INV_X1 U15735 ( .A(n13706), .ZN(n13714) );
  AOI22_X1 U15736 ( .A1(n14585), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n13713) );
  NAND2_X1 U15737 ( .A1(n14676), .A2(n13707), .ZN(n13712) );
  OAI211_X1 U15738 ( .C1(n13710), .C2(n13709), .A(n14633), .B(n13708), .ZN(
        n13711) );
  NAND4_X1 U15739 ( .A1(n13714), .A2(n13713), .A3(n13712), .A4(n13711), .ZN(
        P1_U3244) );
  NAND2_X1 U15740 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n13715) );
  OAI21_X1 U15741 ( .B1(n14679), .B2(n13716), .A(n13715), .ZN(n13717) );
  AOI21_X1 U15742 ( .B1(n6715), .B2(n14676), .A(n13717), .ZN(n13727) );
  AOI211_X1 U15743 ( .C1(n13720), .C2(n13719), .A(n13718), .B(n14665), .ZN(
        n13721) );
  INV_X1 U15744 ( .A(n13721), .ZN(n13726) );
  OAI211_X1 U15745 ( .C1(n13724), .C2(n13723), .A(n14633), .B(n13722), .ZN(
        n13725) );
  NAND3_X1 U15746 ( .A1(n13727), .A2(n13726), .A3(n13725), .ZN(P1_U3246) );
  OAI21_X1 U15747 ( .B1(n13730), .B2(n13729), .A(n13728), .ZN(n13731) );
  NAND2_X1 U15748 ( .A1(n13731), .A2(n14636), .ZN(n13740) );
  NOR2_X1 U15749 ( .A1(n14679), .A2(n14349), .ZN(n13732) );
  AOI211_X1 U15750 ( .C1(n14676), .C2(n13734), .A(n13733), .B(n13732), .ZN(
        n13739) );
  OAI211_X1 U15751 ( .C1(n13737), .C2(n13736), .A(n14633), .B(n13735), .ZN(
        n13738) );
  NAND3_X1 U15752 ( .A1(n13740), .A2(n13739), .A3(n13738), .ZN(P1_U3248) );
  AOI211_X1 U15753 ( .C1(n13743), .C2(n13742), .A(n14665), .B(n13741), .ZN(
        n13744) );
  INV_X1 U15754 ( .A(n13744), .ZN(n13754) );
  INV_X1 U15755 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n13746) );
  OAI21_X1 U15756 ( .B1(n14679), .B2(n13746), .A(n13745), .ZN(n13747) );
  AOI21_X1 U15757 ( .B1(n13748), .B2(n14676), .A(n13747), .ZN(n13753) );
  OAI211_X1 U15758 ( .C1(n13751), .C2(n13750), .A(n14633), .B(n13749), .ZN(
        n13752) );
  NAND3_X1 U15759 ( .A1(n13754), .A2(n13753), .A3(n13752), .ZN(P1_U3250) );
  MUX2_X1 U15760 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n13755), .S(n13782), .Z(
        n13758) );
  OAI21_X1 U15761 ( .B1(n13758), .B2(n13757), .A(n13781), .ZN(n13759) );
  NAND2_X1 U15762 ( .A1(n13759), .A2(n14636), .ZN(n13770) );
  AOI21_X1 U15763 ( .B1(n14585), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n13760), 
        .ZN(n13769) );
  MUX2_X1 U15764 ( .A(n10875), .B(P1_REG2_REG_12__SCAN_IN), .S(n13782), .Z(
        n13763) );
  INV_X1 U15765 ( .A(n13763), .ZN(n13764) );
  NAND2_X1 U15766 ( .A1(n13765), .A2(n13764), .ZN(n13772) );
  OAI21_X1 U15767 ( .B1(n13765), .B2(n13764), .A(n13772), .ZN(n13766) );
  NAND2_X1 U15768 ( .A1(n13766), .A2(n14633), .ZN(n13768) );
  NAND2_X1 U15769 ( .A1(n14676), .A2(n13782), .ZN(n13767) );
  NAND4_X1 U15770 ( .A1(n13770), .A2(n13769), .A3(n13768), .A4(n13767), .ZN(
        P1_U3255) );
  AOI22_X1 U15771 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n13771), .B1(n14610), 
        .B2(n11005), .ZN(n14603) );
  OAI21_X1 U15772 ( .B1(n13782), .B2(P1_REG2_REG_12__SCAN_IN), .A(n13772), 
        .ZN(n14604) );
  NOR2_X1 U15773 ( .A1(n14603), .A2(n14604), .ZN(n14602) );
  NAND2_X1 U15774 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n13783), .ZN(n13773) );
  OAI21_X1 U15775 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n13783), .A(n13773), 
        .ZN(n14620) );
  NOR2_X1 U15776 ( .A1(n14621), .A2(n14620), .ZN(n14619) );
  NAND2_X1 U15777 ( .A1(n13774), .A2(n13786), .ZN(n13775) );
  XOR2_X1 U15778 ( .A(n13774), .B(n13786), .Z(n14632) );
  NAND2_X1 U15779 ( .A1(n14632), .A2(n11296), .ZN(n14631) );
  NAND2_X1 U15780 ( .A1(n13775), .A2(n14631), .ZN(n14646) );
  XNOR2_X1 U15781 ( .A(n14649), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n14645) );
  NOR2_X1 U15782 ( .A1(n14646), .A2(n14645), .ZN(n14644) );
  AOI22_X1 U15783 ( .A1(n14661), .A2(n11358), .B1(P1_REG2_REG_17__SCAN_IN), 
        .B2(n13789), .ZN(n14654) );
  NOR2_X1 U15784 ( .A1(n14655), .A2(n14654), .ZN(n14653) );
  NOR2_X1 U15785 ( .A1(n13776), .A2(n13790), .ZN(n13777) );
  XNOR2_X1 U15786 ( .A(n13776), .B(n13790), .ZN(n14672) );
  NOR2_X1 U15787 ( .A1(n14671), .A2(n14672), .ZN(n14670) );
  XNOR2_X1 U15788 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n13778), .ZN(n13795) );
  MUX2_X1 U15789 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n13779), .S(n13783), .Z(
        n14616) );
  INV_X1 U15790 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n13780) );
  MUX2_X1 U15791 ( .A(n13780), .B(P1_REG1_REG_13__SCAN_IN), .S(n14610), .Z(
        n14606) );
  OAI21_X1 U15792 ( .B1(n13782), .B2(P1_REG1_REG_12__SCAN_IN), .A(n13781), 
        .ZN(n14607) );
  NOR2_X1 U15793 ( .A1(n14606), .A2(n14607), .ZN(n14605) );
  NAND2_X1 U15794 ( .A1(n13786), .A2(n13784), .ZN(n13787) );
  XNOR2_X1 U15795 ( .A(n13786), .B(n13785), .ZN(n14630) );
  INV_X1 U15796 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14629) );
  NAND2_X1 U15797 ( .A1(n14630), .A2(n14629), .ZN(n14628) );
  NAND2_X1 U15798 ( .A1(n13787), .A2(n14628), .ZN(n14643) );
  XNOR2_X1 U15799 ( .A(n14649), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n14642) );
  NOR2_X1 U15800 ( .A1(n14643), .A2(n14642), .ZN(n14641) );
  AOI21_X1 U15801 ( .B1(n14649), .B2(P1_REG1_REG_16__SCAN_IN), .A(n14641), 
        .ZN(n14658) );
  XNOR2_X1 U15802 ( .A(n13789), .B(n13788), .ZN(n14657) );
  NOR2_X1 U15803 ( .A1(n14658), .A2(n14657), .ZN(n14656) );
  AOI21_X1 U15804 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n14661), .A(n14656), 
        .ZN(n13791) );
  XNOR2_X1 U15805 ( .A(n13790), .B(n13791), .ZN(n14668) );
  NOR2_X1 U15806 ( .A1(n14667), .A2(n14668), .ZN(n14666) );
  NOR2_X1 U15807 ( .A1(n13791), .A2(n13790), .ZN(n13792) );
  NOR2_X1 U15808 ( .A1(n14666), .A2(n13792), .ZN(n13793) );
  XNOR2_X1 U15809 ( .A(n13793), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n13794) );
  AOI22_X1 U15810 ( .A1(n13795), .A2(n14633), .B1(n14636), .B2(n13794), .ZN(
        n13797) );
  INV_X1 U15811 ( .A(n14154), .ZN(n14006) );
  INV_X1 U15812 ( .A(n14070), .ZN(n14068) );
  NAND2_X1 U15813 ( .A1(n14068), .A2(n14067), .ZN(n14066) );
  OR2_X2 U15814 ( .A1(n14174), .A2(n14066), .ZN(n14045) );
  AND2_X2 U15815 ( .A1(n14161), .A2(n14030), .ZN(n14020) );
  NAND2_X1 U15816 ( .A1(n14006), .A2(n14020), .ZN(n14001) );
  INV_X1 U15817 ( .A(n14126), .ZN(n13915) );
  AND2_X2 U15818 ( .A1(n13939), .A2(n13915), .ZN(n13917) );
  INV_X1 U15819 ( .A(n14121), .ZN(n13905) );
  AND2_X2 U15820 ( .A1(n13917), .A2(n13905), .ZN(n13903) );
  INV_X1 U15821 ( .A(n14115), .ZN(n13886) );
  XNOR2_X1 U15822 ( .A(n13807), .B(n14098), .ZN(n13800) );
  NAND2_X1 U15823 ( .A1(n13800), .A2(n14756), .ZN(n14099) );
  NOR2_X1 U15824 ( .A1(n14691), .A2(n13801), .ZN(n13805) );
  NOR2_X1 U15825 ( .A1(n6453), .A2(n13802), .ZN(n13803) );
  NOR2_X1 U15826 ( .A1(n14720), .A2(n13803), .ZN(n13867) );
  NAND2_X1 U15827 ( .A1(n13804), .A2(n13867), .ZN(n14101) );
  NOR2_X1 U15828 ( .A1(n6442), .A2(n14101), .ZN(n13810) );
  AOI211_X1 U15829 ( .C1(n14098), .C2(n14754), .A(n13805), .B(n13810), .ZN(
        n13806) );
  OAI21_X1 U15830 ( .B1(n14099), .B2(n14695), .A(n13806), .ZN(P1_U3263) );
  OAI211_X1 U15831 ( .C1(n14103), .C2(n6968), .A(n13808), .B(n14756), .ZN(
        n14102) );
  NOR2_X1 U15832 ( .A1(n14691), .A2(n13809), .ZN(n13811) );
  AOI211_X1 U15833 ( .C1(n13812), .C2(n14754), .A(n13811), .B(n13810), .ZN(
        n13813) );
  OAI21_X1 U15834 ( .B1(n14102), .B2(n14695), .A(n13813), .ZN(P1_U3264) );
  NAND2_X1 U15835 ( .A1(n13843), .A2(n13840), .ZN(n13814) );
  INV_X1 U15836 ( .A(n13816), .ZN(n13818) );
  OR2_X1 U15837 ( .A1(n14174), .A2(n14166), .ZN(n13819) );
  NAND2_X1 U15838 ( .A1(n13820), .A2(n13819), .ZN(n14038) );
  NAND2_X1 U15839 ( .A1(n14161), .A2(n13996), .ZN(n13822) );
  NOR2_X1 U15840 ( .A1(n14154), .A2(n13823), .ZN(n13824) );
  NAND2_X1 U15841 ( .A1(n13979), .A2(n6813), .ZN(n13826) );
  NAND2_X1 U15842 ( .A1(n14149), .A2(n13851), .ZN(n13825) );
  NAND2_X1 U15843 ( .A1(n13826), .A2(n13825), .ZN(n13974) );
  NAND2_X1 U15844 ( .A1(n13974), .A2(n13973), .ZN(n13972) );
  NAND2_X1 U15845 ( .A1(n14144), .A2(n13961), .ZN(n13828) );
  OR2_X1 U15846 ( .A1(n14139), .A2(n13945), .ZN(n13830) );
  NAND2_X1 U15847 ( .A1(n13920), .A2(n13895), .ZN(n13831) );
  NAND2_X1 U15848 ( .A1(n14121), .A2(n13832), .ZN(n13833) );
  OR2_X1 U15849 ( .A1(n14115), .A2(n13899), .ZN(n13834) );
  NAND2_X1 U15850 ( .A1(n13878), .A2(n13834), .ZN(n13836) );
  NAND2_X1 U15851 ( .A1(n14115), .A2(n13899), .ZN(n13835) );
  NAND2_X1 U15852 ( .A1(n13836), .A2(n13835), .ZN(n13838) );
  XNOR2_X1 U15853 ( .A(n13838), .B(n13861), .ZN(n13839) );
  NAND2_X1 U15854 ( .A1(n13839), .A2(n14685), .ZN(n14112) );
  INV_X1 U15855 ( .A(n13845), .ZN(n13847) );
  NAND2_X1 U15856 ( .A1(n13852), .A2(n13851), .ZN(n13853) );
  NOR2_X1 U15857 ( .A1(n14144), .A2(n13980), .ZN(n13855) );
  NAND2_X1 U15858 ( .A1(n14144), .A2(n13980), .ZN(n13950) );
  INV_X1 U15859 ( .A(n14139), .ZN(n13957) );
  NAND2_X1 U15860 ( .A1(n13957), .A2(n13945), .ZN(n13856) );
  INV_X1 U15861 ( .A(n14133), .ZN(n13857) );
  XNOR2_X1 U15862 ( .A(n13862), .B(n13861), .ZN(n14104) );
  NAND2_X1 U15863 ( .A1(n14104), .A2(n14697), .ZN(n13876) );
  AOI21_X1 U15864 ( .B1(n13888), .B2(n14109), .A(n14090), .ZN(n13864) );
  NAND2_X1 U15865 ( .A1(n13864), .A2(n13863), .ZN(n14110) );
  OR2_X1 U15866 ( .A1(n6442), .A2(n14722), .ZN(n14031) );
  NOR2_X1 U15867 ( .A1(n14751), .A2(n13865), .ZN(n13866) );
  AOI21_X1 U15868 ( .B1(n6442), .B2(P1_REG2_REG_29__SCAN_IN), .A(n13866), .ZN(
        n13871) );
  NAND2_X1 U15869 ( .A1(n13868), .A2(n13867), .ZN(n14107) );
  OR2_X1 U15870 ( .A1(n14107), .A2(n13869), .ZN(n13870) );
  OAI211_X1 U15871 ( .C1(n14031), .C2(n13899), .A(n13871), .B(n13870), .ZN(
        n13872) );
  AOI21_X1 U15872 ( .B1(n14109), .B2(n14754), .A(n13872), .ZN(n13873) );
  OAI21_X1 U15873 ( .B1(n14110), .B2(n14695), .A(n13873), .ZN(n13874) );
  INV_X1 U15874 ( .A(n13874), .ZN(n13875) );
  OAI211_X1 U15875 ( .C1(n6442), .C2(n14112), .A(n13876), .B(n13875), .ZN(
        P1_U3356) );
  NAND2_X1 U15876 ( .A1(n13880), .A2(n7179), .ZN(n13881) );
  NAND2_X1 U15877 ( .A1(n13882), .A2(n13881), .ZN(n14118) );
  NAND2_X1 U15878 ( .A1(n6442), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n13883) );
  OAI21_X1 U15879 ( .B1(n14751), .B2(n13884), .A(n13883), .ZN(n13885) );
  AOI21_X1 U15880 ( .B1(n14115), .B2(n14754), .A(n13885), .ZN(n13890) );
  OR2_X1 U15881 ( .A1(n13903), .A2(n13886), .ZN(n13887) );
  NAND2_X1 U15882 ( .A1(n14114), .A2(n14759), .ZN(n13889) );
  OAI211_X1 U15883 ( .C1(n14118), .C2(n14059), .A(n13890), .B(n13889), .ZN(
        n13891) );
  INV_X1 U15884 ( .A(n13891), .ZN(n13892) );
  OAI21_X1 U15885 ( .B1(n14117), .B2(n6442), .A(n13892), .ZN(P1_U3265) );
  NAND3_X1 U15886 ( .A1(n13920), .A2(n13896), .A3(n13895), .ZN(n13897) );
  AOI21_X1 U15887 ( .B1(n13898), .B2(n13897), .A(n14744), .ZN(n13902) );
  OAI22_X1 U15888 ( .A1(n13900), .A2(n14722), .B1(n13899), .B2(n14720), .ZN(
        n13901) );
  INV_X1 U15889 ( .A(n13917), .ZN(n13904) );
  AOI211_X1 U15890 ( .C1(n14121), .C2(n13904), .A(n14090), .B(n13903), .ZN(
        n14120) );
  NOR2_X1 U15891 ( .A1(n13905), .A2(n14047), .ZN(n13909) );
  OAI22_X1 U15892 ( .A1(n14691), .A2(n13907), .B1(n13906), .B2(n14751), .ZN(
        n13908) );
  AOI211_X1 U15893 ( .C1(n14120), .C2(n14759), .A(n13909), .B(n13908), .ZN(
        n13911) );
  NAND2_X1 U15894 ( .A1(n14119), .A2(n14760), .ZN(n13910) );
  OAI211_X1 U15895 ( .C1(n6571), .C2(n6442), .A(n13911), .B(n13910), .ZN(
        P1_U3266) );
  XNOR2_X1 U15896 ( .A(n13912), .B(n13922), .ZN(n14124) );
  INV_X1 U15897 ( .A(n14124), .ZN(n13931) );
  OAI22_X1 U15898 ( .A1(n14691), .A2(n13914), .B1(n13913), .B2(n14751), .ZN(
        n13919) );
  OAI21_X1 U15899 ( .B1(n13939), .B2(n13915), .A(n14756), .ZN(n13916) );
  NOR2_X1 U15900 ( .A1(n14127), .A2(n14695), .ZN(n13918) );
  AOI211_X1 U15901 ( .C1(n14754), .C2(n14126), .A(n13919), .B(n13918), .ZN(
        n13930) );
  OAI21_X1 U15902 ( .B1(n13922), .B2(n13921), .A(n13920), .ZN(n13923) );
  NAND2_X1 U15903 ( .A1(n13923), .A2(n14685), .ZN(n14128) );
  INV_X1 U15904 ( .A(n14128), .ZN(n13928) );
  NAND2_X1 U15905 ( .A1(n13924), .A2(n14705), .ZN(n13927) );
  NAND2_X1 U15906 ( .A1(n13925), .A2(n14702), .ZN(n13926) );
  NAND2_X1 U15907 ( .A1(n13927), .A2(n13926), .ZN(n14125) );
  OAI21_X1 U15908 ( .B1(n13928), .B2(n14125), .A(n14691), .ZN(n13929) );
  OAI211_X1 U15909 ( .C1(n13931), .C2(n14059), .A(n13930), .B(n13929), .ZN(
        P1_U3267) );
  OAI21_X1 U15910 ( .B1(n6526), .B2(n13938), .A(n13932), .ZN(n13934) );
  AOI22_X1 U15911 ( .A1(n13934), .A2(n14685), .B1(n14702), .B2(n13933), .ZN(
        n14136) );
  INV_X1 U15912 ( .A(n13935), .ZN(n13936) );
  AOI21_X1 U15913 ( .B1(n13938), .B2(n13937), .A(n13936), .ZN(n14131) );
  INV_X1 U15914 ( .A(n13939), .ZN(n13941) );
  AOI21_X1 U15915 ( .B1(n13953), .B2(n14133), .A(n14090), .ZN(n13940) );
  NAND2_X1 U15916 ( .A1(n13941), .A2(n13940), .ZN(n14134) );
  NOR2_X1 U15917 ( .A1(n14751), .A2(n13942), .ZN(n13943) );
  AOI21_X1 U15918 ( .B1(n6442), .B2(P1_REG2_REG_25__SCAN_IN), .A(n13943), .ZN(
        n13944) );
  OAI21_X1 U15919 ( .B1(n14031), .B2(n13945), .A(n13944), .ZN(n13946) );
  AOI21_X1 U15920 ( .B1(n14133), .B2(n14754), .A(n13946), .ZN(n13947) );
  OAI21_X1 U15921 ( .B1(n14134), .B2(n14695), .A(n13947), .ZN(n13948) );
  AOI21_X1 U15922 ( .B1(n14131), .B2(n14697), .A(n13948), .ZN(n13949) );
  OAI21_X1 U15923 ( .B1(n6442), .B2(n14136), .A(n13949), .ZN(P1_U3268) );
  NAND2_X1 U15924 ( .A1(n13951), .A2(n13950), .ZN(n13952) );
  XNOR2_X1 U15925 ( .A(n13952), .B(n13958), .ZN(n14142) );
  INV_X1 U15926 ( .A(n13953), .ZN(n13954) );
  AOI211_X1 U15927 ( .C1(n14139), .C2(n13969), .A(n14090), .B(n13954), .ZN(
        n14138) );
  AOI22_X1 U15928 ( .A1(n6442), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n13955), 
        .B2(n14710), .ZN(n13956) );
  OAI21_X1 U15929 ( .B1(n13957), .B2(n14047), .A(n13956), .ZN(n13966) );
  AOI21_X1 U15930 ( .B1(n13959), .B2(n13958), .A(n14744), .ZN(n13964) );
  OAI22_X1 U15931 ( .A1(n13961), .A2(n14722), .B1(n13960), .B2(n14720), .ZN(
        n13962) );
  AOI21_X1 U15932 ( .B1(n13964), .B2(n13963), .A(n13962), .ZN(n14141) );
  NOR2_X1 U15933 ( .A1(n14141), .A2(n6442), .ZN(n13965) );
  AOI211_X1 U15934 ( .C1(n14138), .C2(n14759), .A(n13966), .B(n13965), .ZN(
        n13967) );
  OAI21_X1 U15935 ( .B1(n14142), .B2(n14059), .A(n13967), .ZN(P1_U3269) );
  XNOR2_X1 U15936 ( .A(n13968), .B(n13973), .ZN(n14147) );
  AOI211_X1 U15937 ( .C1(n14144), .C2(n13986), .A(n14090), .B(n6441), .ZN(
        n14143) );
  AOI22_X1 U15938 ( .A1(n6442), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n13970), 
        .B2(n14710), .ZN(n13971) );
  OAI21_X1 U15939 ( .B1(n6959), .B2(n14047), .A(n13971), .ZN(n13977) );
  OAI21_X1 U15940 ( .B1(n13974), .B2(n13973), .A(n13972), .ZN(n13975) );
  AOI222_X1 U15941 ( .A1(n14685), .A2(n13975), .B1(n14132), .B2(n14702), .C1(
        n13995), .C2(n14705), .ZN(n14146) );
  NOR2_X1 U15942 ( .A1(n14146), .A2(n6442), .ZN(n13976) );
  AOI211_X1 U15943 ( .C1(n14143), .C2(n14759), .A(n13977), .B(n13976), .ZN(
        n13978) );
  OAI21_X1 U15944 ( .B1(n14147), .B2(n14059), .A(n13978), .ZN(P1_U3270) );
  XNOR2_X1 U15945 ( .A(n13979), .B(n6813), .ZN(n13981) );
  AOI222_X1 U15946 ( .A1(n14685), .A2(n13981), .B1(n13980), .B2(n14702), .C1(
        n14017), .C2(n14705), .ZN(n14151) );
  XNOR2_X1 U15947 ( .A(n13982), .B(n6813), .ZN(n14152) );
  NAND2_X1 U15948 ( .A1(n6442), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n13983) );
  OAI21_X1 U15949 ( .B1(n14751), .B2(n13984), .A(n13983), .ZN(n13985) );
  AOI21_X1 U15950 ( .B1(n14149), .B2(n14754), .A(n13985), .ZN(n13989) );
  AOI21_X1 U15951 ( .B1(n14149), .B2(n14001), .A(n14090), .ZN(n13987) );
  AND2_X1 U15952 ( .A1(n13987), .A2(n13986), .ZN(n14148) );
  NAND2_X1 U15953 ( .A1(n14148), .A2(n14759), .ZN(n13988) );
  OAI211_X1 U15954 ( .C1(n14152), .C2(n14059), .A(n13989), .B(n13988), .ZN(
        n13990) );
  INV_X1 U15955 ( .A(n13990), .ZN(n13991) );
  OAI21_X1 U15956 ( .B1(n6442), .B2(n14151), .A(n13991), .ZN(P1_U3271) );
  XNOR2_X1 U15957 ( .A(n13993), .B(n13992), .ZN(n13994) );
  AOI222_X1 U15958 ( .A1(n13996), .A2(n14705), .B1(n13995), .B2(n14702), .C1(
        n14685), .C2(n13994), .ZN(n14156) );
  AOI21_X1 U15959 ( .B1(n13999), .B2(n13998), .A(n6808), .ZN(n14157) );
  INV_X1 U15960 ( .A(n14157), .ZN(n14008) );
  OR2_X1 U15961 ( .A1(n14006), .A2(n14020), .ZN(n14000) );
  AND3_X1 U15962 ( .A1(n14001), .A2(n14756), .A3(n14000), .ZN(n14153) );
  NAND2_X1 U15963 ( .A1(n14153), .A2(n14759), .ZN(n14005) );
  INV_X1 U15964 ( .A(n14002), .ZN(n14003) );
  AOI22_X1 U15965 ( .A1(n14003), .A2(n14710), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n6442), .ZN(n14004) );
  OAI211_X1 U15966 ( .C1(n14006), .C2(n14047), .A(n14005), .B(n14004), .ZN(
        n14007) );
  AOI21_X1 U15967 ( .B1(n14008), .B2(n14697), .A(n14007), .ZN(n14009) );
  OAI21_X1 U15968 ( .B1(n6442), .B2(n14156), .A(n14009), .ZN(P1_U3272) );
  NAND2_X1 U15969 ( .A1(n14011), .A2(n14010), .ZN(n14158) );
  NAND3_X1 U15970 ( .A1(n14159), .A2(n14158), .A3(n14697), .ZN(n14025) );
  AOI22_X1 U15971 ( .A1(n14012), .A2(n14754), .B1(n6442), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n14024) );
  INV_X1 U15972 ( .A(n14013), .ZN(n14014) );
  AOI211_X1 U15973 ( .C1(n7169), .C2(n14015), .A(n14744), .B(n14014), .ZN(
        n14164) );
  AOI22_X1 U15974 ( .A1(n14017), .A2(n14702), .B1(n14705), .B2(n14016), .ZN(
        n14160) );
  OAI21_X1 U15975 ( .B1(n14018), .B2(n14751), .A(n14160), .ZN(n14019) );
  OAI21_X1 U15976 ( .B1(n14164), .B2(n14019), .A(n14691), .ZN(n14023) );
  OAI21_X1 U15977 ( .B1(n14161), .B2(n14030), .A(n14756), .ZN(n14021) );
  NOR2_X1 U15978 ( .A1(n14021), .A2(n14020), .ZN(n14163) );
  NAND2_X1 U15979 ( .A1(n14163), .A2(n14759), .ZN(n14022) );
  NAND4_X1 U15980 ( .A1(n14025), .A2(n14024), .A3(n14023), .A4(n14022), .ZN(
        P1_U3273) );
  XOR2_X1 U15981 ( .A(n14026), .B(n14039), .Z(n14171) );
  NAND2_X1 U15982 ( .A1(n14027), .A2(n14045), .ZN(n14028) );
  NAND2_X1 U15983 ( .A1(n14028), .A2(n14756), .ZN(n14029) );
  NOR2_X1 U15984 ( .A1(n14030), .A2(n14029), .ZN(n14168) );
  INV_X1 U15985 ( .A(n14031), .ZN(n14035) );
  OAI22_X1 U15986 ( .A1(n14691), .A2(n14033), .B1(n14032), .B2(n14751), .ZN(
        n14034) );
  AOI21_X1 U15987 ( .B1(n14035), .B2(n14065), .A(n14034), .ZN(n14036) );
  OAI21_X1 U15988 ( .B1(n13848), .B2(n14047), .A(n14036), .ZN(n14037) );
  AOI21_X1 U15989 ( .B1(n14168), .B2(n14759), .A(n14037), .ZN(n14043) );
  XOR2_X1 U15990 ( .A(n14038), .B(n14039), .Z(n14041) );
  OAI22_X1 U15991 ( .A1(n14041), .A2(n14744), .B1(n14040), .B2(n14720), .ZN(
        n14169) );
  NAND2_X1 U15992 ( .A1(n14169), .A2(n14691), .ZN(n14042) );
  OAI211_X1 U15993 ( .C1(n14171), .C2(n14059), .A(n14043), .B(n14042), .ZN(
        P1_U3274) );
  XOR2_X1 U15994 ( .A(n14044), .B(n14050), .Z(n14176) );
  INV_X1 U15995 ( .A(n14045), .ZN(n14046) );
  AOI211_X1 U15996 ( .C1(n14174), .C2(n14066), .A(n14090), .B(n14046), .ZN(
        n14173) );
  INV_X1 U15997 ( .A(n14174), .ZN(n14048) );
  OAI22_X1 U15998 ( .A1(n14048), .A2(n14047), .B1(n14671), .B2(n14691), .ZN(
        n14049) );
  AOI21_X1 U15999 ( .B1(n14173), .B2(n14759), .A(n14049), .ZN(n14058) );
  XNOR2_X1 U16000 ( .A(n14051), .B(n14050), .ZN(n14053) );
  OAI222_X1 U16001 ( .A1(n14720), .A2(n14054), .B1(n14053), .B2(n14744), .C1(
        n14722), .C2(n14052), .ZN(n14172) );
  NOR2_X1 U16002 ( .A1(n14055), .A2(n14751), .ZN(n14056) );
  OAI21_X1 U16003 ( .B1(n14172), .B2(n14056), .A(n14691), .ZN(n14057) );
  OAI211_X1 U16004 ( .C1(n14176), .C2(n14059), .A(n14058), .B(n14057), .ZN(
        P1_U3275) );
  XOR2_X1 U16005 ( .A(n14061), .B(n14060), .Z(n14182) );
  XNOR2_X1 U16006 ( .A(n14062), .B(n14061), .ZN(n14063) );
  NAND2_X1 U16007 ( .A1(n14063), .A2(n14685), .ZN(n14180) );
  AOI22_X1 U16008 ( .A1(n14065), .A2(n14702), .B1(n14064), .B2(n14705), .ZN(
        n14179) );
  AOI21_X1 U16009 ( .B1(n14180), .B2(n14179), .A(n6442), .ZN(n14074) );
  OAI211_X1 U16010 ( .C1(n14068), .C2(n14067), .A(n14756), .B(n14066), .ZN(
        n14177) );
  AOI22_X1 U16011 ( .A1(n6442), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n14069), 
        .B2(n14710), .ZN(n14072) );
  NAND2_X1 U16012 ( .A1(n14070), .A2(n14754), .ZN(n14071) );
  OAI211_X1 U16013 ( .C1(n14177), .C2(n14695), .A(n14072), .B(n14071), .ZN(
        n14073) );
  AOI211_X1 U16014 ( .C1(n14182), .C2(n14697), .A(n14074), .B(n14073), .ZN(
        n14075) );
  INV_X1 U16015 ( .A(n14075), .ZN(P1_U3276) );
  AOI21_X1 U16016 ( .B1(n14078), .B2(n14077), .A(n14076), .ZN(n14191) );
  NAND2_X1 U16017 ( .A1(n14191), .A2(n14697), .ZN(n14097) );
  NAND2_X1 U16018 ( .A1(n6442), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n14079) );
  OAI21_X1 U16019 ( .B1(n14751), .B2(n14080), .A(n14079), .ZN(n14081) );
  AOI21_X1 U16020 ( .B1(n14194), .B2(n14754), .A(n14081), .ZN(n14096) );
  XNOR2_X1 U16021 ( .A(n14083), .B(n14082), .ZN(n14084) );
  NAND2_X1 U16022 ( .A1(n14084), .A2(n14685), .ZN(n14195) );
  INV_X1 U16023 ( .A(n14195), .ZN(n14089) );
  OR2_X1 U16024 ( .A1(n14085), .A2(n14720), .ZN(n14088) );
  NAND2_X1 U16025 ( .A1(n14086), .A2(n14705), .ZN(n14087) );
  NAND2_X1 U16026 ( .A1(n14088), .A2(n14087), .ZN(n14193) );
  OAI21_X1 U16027 ( .B1(n14089), .B2(n14193), .A(n14691), .ZN(n14095) );
  AOI21_X1 U16028 ( .B1(n14091), .B2(n14194), .A(n14090), .ZN(n14093) );
  AND2_X1 U16029 ( .A1(n14093), .A2(n14092), .ZN(n14192) );
  NAND2_X1 U16030 ( .A1(n14192), .A2(n14759), .ZN(n14094) );
  NAND4_X1 U16031 ( .A1(n14097), .A2(n14096), .A3(n14095), .A4(n14094), .ZN(
        P1_U3279) );
  INV_X1 U16032 ( .A(n14098), .ZN(n14100) );
  OAI211_X1 U16033 ( .C1(n14100), .C2(n14821), .A(n14099), .B(n14101), .ZN(
        n14199) );
  MUX2_X1 U16034 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14199), .S(n14839), .Z(
        P1_U3559) );
  OAI211_X1 U16035 ( .C1(n14103), .C2(n14821), .A(n14102), .B(n14101), .ZN(
        n14200) );
  MUX2_X1 U16036 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14200), .S(n14839), .Z(
        P1_U3558) );
  NAND2_X1 U16037 ( .A1(n14104), .A2(n14824), .ZN(n14113) );
  NAND2_X1 U16038 ( .A1(n14105), .A2(n14705), .ZN(n14106) );
  NAND2_X1 U16039 ( .A1(n14107), .A2(n14106), .ZN(n14108) );
  AOI21_X1 U16040 ( .B1(n14109), .B2(n14792), .A(n14108), .ZN(n14111) );
  MUX2_X1 U16041 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14201), .S(n14839), .Z(
        P1_U3557) );
  AOI21_X1 U16042 ( .B1(n14115), .B2(n14792), .A(n14114), .ZN(n14116) );
  MUX2_X1 U16043 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14202), .S(n14839), .Z(
        P1_U3556) );
  INV_X1 U16044 ( .A(n14119), .ZN(n14123) );
  AOI21_X1 U16045 ( .B1(n14121), .B2(n14792), .A(n14120), .ZN(n14122) );
  MUX2_X1 U16046 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14203), .S(n14839), .Z(
        P1_U3555) );
  NAND2_X1 U16047 ( .A1(n14124), .A2(n14824), .ZN(n14130) );
  AOI21_X1 U16048 ( .B1(n14126), .B2(n14792), .A(n14125), .ZN(n14129) );
  NAND4_X1 U16049 ( .A1(n14130), .A2(n14129), .A3(n14128), .A4(n14127), .ZN(
        n14204) );
  MUX2_X1 U16050 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14204), .S(n14839), .Z(
        P1_U3554) );
  NAND2_X1 U16051 ( .A1(n14131), .A2(n14824), .ZN(n14137) );
  AOI22_X1 U16052 ( .A1(n14133), .A2(n14792), .B1(n14705), .B2(n14132), .ZN(
        n14135) );
  NAND4_X1 U16053 ( .A1(n14137), .A2(n14136), .A3(n14135), .A4(n14134), .ZN(
        n14205) );
  MUX2_X1 U16054 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14205), .S(n14839), .Z(
        P1_U3553) );
  AOI21_X1 U16055 ( .B1(n14139), .B2(n14792), .A(n14138), .ZN(n14140) );
  OAI211_X1 U16056 ( .C1(n14142), .C2(n14197), .A(n14141), .B(n14140), .ZN(
        n14206) );
  MUX2_X1 U16057 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14206), .S(n14839), .Z(
        P1_U3552) );
  AOI21_X1 U16058 ( .B1(n14144), .B2(n14792), .A(n14143), .ZN(n14145) );
  OAI211_X1 U16059 ( .C1(n14147), .C2(n14197), .A(n14146), .B(n14145), .ZN(
        n14207) );
  MUX2_X1 U16060 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14207), .S(n14839), .Z(
        P1_U3551) );
  AOI21_X1 U16061 ( .B1(n14149), .B2(n14792), .A(n14148), .ZN(n14150) );
  OAI211_X1 U16062 ( .C1(n14152), .C2(n14197), .A(n14151), .B(n14150), .ZN(
        n14208) );
  MUX2_X1 U16063 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14208), .S(n14839), .Z(
        P1_U3550) );
  AOI21_X1 U16064 ( .B1(n14154), .B2(n14792), .A(n14153), .ZN(n14155) );
  OAI211_X1 U16065 ( .C1(n14157), .C2(n14197), .A(n14156), .B(n14155), .ZN(
        n14209) );
  MUX2_X1 U16066 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14209), .S(n14839), .Z(
        P1_U3549) );
  AND3_X1 U16067 ( .A1(n14159), .A2(n14158), .A3(n14824), .ZN(n14165) );
  OAI21_X1 U16068 ( .B1(n14161), .B2(n14821), .A(n14160), .ZN(n14162) );
  MUX2_X1 U16069 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14210), .S(n14839), .Z(
        P1_U3548) );
  OAI22_X1 U16070 ( .A1(n13848), .A2(n14821), .B1(n14166), .B2(n14722), .ZN(
        n14167) );
  NOR3_X1 U16071 ( .A1(n14169), .A2(n14168), .A3(n14167), .ZN(n14170) );
  OAI21_X1 U16072 ( .B1(n14171), .B2(n14197), .A(n14170), .ZN(n14211) );
  MUX2_X1 U16073 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14211), .S(n14839), .Z(
        P1_U3547) );
  AOI211_X1 U16074 ( .C1(n14174), .C2(n14792), .A(n14173), .B(n14172), .ZN(
        n14175) );
  OAI21_X1 U16075 ( .B1(n14176), .B2(n14197), .A(n14175), .ZN(n14212) );
  MUX2_X1 U16076 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14212), .S(n14839), .Z(
        P1_U3546) );
  NAND4_X1 U16077 ( .A1(n14180), .A2(n14179), .A3(n14178), .A4(n14177), .ZN(
        n14181) );
  AOI21_X1 U16078 ( .B1(n14182), .B2(n14824), .A(n14181), .ZN(n14183) );
  INV_X1 U16079 ( .A(n14183), .ZN(n14213) );
  MUX2_X1 U16080 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14213), .S(n14839), .Z(
        P1_U3545) );
  NAND3_X1 U16081 ( .A1(n14186), .A2(n14185), .A3(n14184), .ZN(n14187) );
  AOI211_X1 U16082 ( .C1(n14189), .C2(n14824), .A(n14188), .B(n14187), .ZN(
        n14190) );
  INV_X1 U16083 ( .A(n14190), .ZN(n14214) );
  MUX2_X1 U16084 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14214), .S(n14839), .Z(
        P1_U3544) );
  INV_X1 U16085 ( .A(n14191), .ZN(n14198) );
  AOI211_X1 U16086 ( .C1(n14194), .C2(n14792), .A(n14193), .B(n14192), .ZN(
        n14196) );
  OAI211_X1 U16087 ( .C1(n14198), .C2(n14197), .A(n14196), .B(n14195), .ZN(
        n14215) );
  MUX2_X1 U16088 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n14215), .S(n14839), .Z(
        P1_U3542) );
  MUX2_X1 U16089 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14199), .S(n14827), .Z(
        P1_U3527) );
  MUX2_X1 U16090 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14200), .S(n14827), .Z(
        P1_U3526) );
  MUX2_X1 U16091 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14201), .S(n14827), .Z(
        P1_U3525) );
  MUX2_X1 U16092 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14202), .S(n14827), .Z(
        P1_U3524) );
  MUX2_X1 U16093 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14204), .S(n14827), .Z(
        P1_U3522) );
  MUX2_X1 U16094 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14205), .S(n14827), .Z(
        P1_U3521) );
  MUX2_X1 U16095 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14206), .S(n14827), .Z(
        P1_U3520) );
  MUX2_X1 U16096 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14207), .S(n14827), .Z(
        P1_U3519) );
  MUX2_X1 U16097 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14208), .S(n14827), .Z(
        P1_U3518) );
  MUX2_X1 U16098 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14209), .S(n14827), .Z(
        P1_U3517) );
  MUX2_X1 U16099 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14210), .S(n14827), .Z(
        P1_U3516) );
  MUX2_X1 U16100 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14211), .S(n14827), .Z(
        P1_U3515) );
  MUX2_X1 U16101 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14212), .S(n14827), .Z(
        P1_U3513) );
  MUX2_X1 U16102 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14213), .S(n14827), .Z(
        P1_U3510) );
  MUX2_X1 U16103 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14214), .S(n14827), .Z(
        P1_U3507) );
  MUX2_X1 U16104 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n14215), .S(n14827), .Z(
        P1_U3501) );
  NOR4_X1 U16105 ( .A1(n14217), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n14216), .ZN(n14220) );
  NOR2_X1 U16106 ( .A1(n14372), .A2(n14218), .ZN(n14219) );
  AOI211_X1 U16107 ( .C1(n14222), .C2(n14221), .A(n14220), .B(n14219), .ZN(
        n14365) );
  AOI22_X1 U16108 ( .A1(n14335), .A2(keyinput15), .B1(n10597), .B2(keyinput10), 
        .ZN(n14223) );
  OAI221_X1 U16109 ( .B1(n14335), .B2(keyinput15), .C1(n10597), .C2(keyinput10), .A(n14223), .ZN(n14234) );
  AOI22_X1 U16110 ( .A1(n14226), .A2(keyinput2), .B1(n14225), .B2(keyinput42), 
        .ZN(n14224) );
  OAI221_X1 U16111 ( .B1(n14226), .B2(keyinput2), .C1(n14225), .C2(keyinput42), 
        .A(n14224), .ZN(n14233) );
  INV_X1 U16112 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n14228) );
  AOI22_X1 U16113 ( .A1(n13322), .A2(keyinput47), .B1(keyinput3), .B2(n14228), 
        .ZN(n14227) );
  OAI221_X1 U16114 ( .B1(n13322), .B2(keyinput47), .C1(n14228), .C2(keyinput3), 
        .A(n14227), .ZN(n14232) );
  AOI22_X1 U16115 ( .A1(n14230), .A2(keyinput58), .B1(n7806), .B2(keyinput43), 
        .ZN(n14229) );
  OAI221_X1 U16116 ( .B1(n14230), .B2(keyinput58), .C1(n7806), .C2(keyinput43), 
        .A(n14229), .ZN(n14231) );
  NOR4_X1 U16117 ( .A1(n14234), .A2(n14233), .A3(n14232), .A4(n14231), .ZN(
        n14250) );
  INV_X1 U16118 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n14236) );
  AOI22_X1 U16119 ( .A1(n14237), .A2(keyinput34), .B1(keyinput1), .B2(n14236), 
        .ZN(n14235) );
  OAI221_X1 U16120 ( .B1(n14237), .B2(keyinput34), .C1(n14236), .C2(keyinput1), 
        .A(n14235), .ZN(n14248) );
  INV_X1 U16121 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n14763) );
  AOI22_X1 U16122 ( .A1(n14763), .A2(keyinput61), .B1(n14239), .B2(keyinput6), 
        .ZN(n14238) );
  OAI221_X1 U16123 ( .B1(n14763), .B2(keyinput61), .C1(n14239), .C2(keyinput6), 
        .A(n14238), .ZN(n14247) );
  AOI22_X1 U16124 ( .A1(n14242), .A2(keyinput24), .B1(keyinput33), .B2(n14241), 
        .ZN(n14240) );
  OAI221_X1 U16125 ( .B1(n14242), .B2(keyinput24), .C1(n14241), .C2(keyinput33), .A(n14240), .ZN(n14246) );
  AOI22_X1 U16126 ( .A1(n14244), .A2(keyinput57), .B1(n14350), .B2(keyinput19), 
        .ZN(n14243) );
  OAI221_X1 U16127 ( .B1(n14244), .B2(keyinput57), .C1(n14350), .C2(keyinput19), .A(n14243), .ZN(n14245) );
  NOR4_X1 U16128 ( .A1(n14248), .A2(n14247), .A3(n14246), .A4(n14245), .ZN(
        n14249) );
  NAND2_X1 U16129 ( .A1(n14250), .A2(n14249), .ZN(n14304) );
  AOI22_X1 U16130 ( .A1(n14252), .A2(keyinput60), .B1(n14351), .B2(keyinput51), 
        .ZN(n14251) );
  OAI221_X1 U16131 ( .B1(n14252), .B2(keyinput60), .C1(n14351), .C2(keyinput51), .A(n14251), .ZN(n14262) );
  AOI22_X1 U16132 ( .A1(n15007), .A2(keyinput45), .B1(n14254), .B2(keyinput41), 
        .ZN(n14253) );
  OAI221_X1 U16133 ( .B1(n15007), .B2(keyinput45), .C1(n14254), .C2(keyinput41), .A(n14253), .ZN(n14261) );
  AOI22_X1 U16134 ( .A1(n9829), .A2(keyinput50), .B1(n8754), .B2(keyinput56), 
        .ZN(n14255) );
  OAI221_X1 U16135 ( .B1(n9829), .B2(keyinput50), .C1(n8754), .C2(keyinput56), 
        .A(n14255), .ZN(n14260) );
  AOI22_X1 U16136 ( .A1(n14258), .A2(keyinput13), .B1(n14257), .B2(keyinput16), 
        .ZN(n14256) );
  OAI221_X1 U16137 ( .B1(n14258), .B2(keyinput13), .C1(n14257), .C2(keyinput16), .A(n14256), .ZN(n14259) );
  NOR4_X1 U16138 ( .A1(n14262), .A2(n14261), .A3(n14260), .A4(n14259), .ZN(
        n14302) );
  INV_X1 U16139 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n14876) );
  AOI22_X1 U16140 ( .A1(n14264), .A2(keyinput31), .B1(n14876), .B2(keyinput52), 
        .ZN(n14263) );
  OAI221_X1 U16141 ( .B1(n14264), .B2(keyinput31), .C1(n14876), .C2(keyinput52), .A(n14263), .ZN(n14268) );
  AOI22_X1 U16142 ( .A1(n14266), .A2(keyinput23), .B1(n9053), .B2(keyinput35), 
        .ZN(n14265) );
  OAI221_X1 U16143 ( .B1(n14266), .B2(keyinput23), .C1(n9053), .C2(keyinput35), 
        .A(n14265), .ZN(n14267) );
  NOR2_X1 U16144 ( .A1(n14268), .A2(n14267), .ZN(n14301) );
  AOI22_X1 U16145 ( .A1(n10854), .A2(keyinput25), .B1(keyinput62), .B2(n9606), 
        .ZN(n14269) );
  OAI221_X1 U16146 ( .B1(n10854), .B2(keyinput25), .C1(n9606), .C2(keyinput62), 
        .A(n14269), .ZN(n14274) );
  AOI22_X1 U16147 ( .A1(n14272), .A2(keyinput55), .B1(keyinput7), .B2(n14271), 
        .ZN(n14270) );
  OAI221_X1 U16148 ( .B1(n14272), .B2(keyinput55), .C1(n14271), .C2(keyinput7), 
        .A(n14270), .ZN(n14273) );
  NOR2_X1 U16149 ( .A1(n14274), .A2(n14273), .ZN(n14300) );
  AOI22_X1 U16150 ( .A1(n7110), .A2(keyinput54), .B1(n14349), .B2(keyinput9), 
        .ZN(n14275) );
  OAI221_X1 U16151 ( .B1(n7110), .B2(keyinput54), .C1(n14349), .C2(keyinput9), 
        .A(n14275), .ZN(n14279) );
  AOI22_X1 U16152 ( .A1(n14345), .A2(keyinput30), .B1(keyinput5), .B2(n14277), 
        .ZN(n14276) );
  OAI221_X1 U16153 ( .B1(n14345), .B2(keyinput30), .C1(n14277), .C2(keyinput5), 
        .A(n14276), .ZN(n14278) );
  NOR2_X1 U16154 ( .A1(n14279), .A2(n14278), .ZN(n14298) );
  XNOR2_X1 U16155 ( .A(P1_REG0_REG_24__SCAN_IN), .B(keyinput26), .ZN(n14283)
         );
  XNOR2_X1 U16156 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput46), .ZN(n14282) );
  XNOR2_X1 U16157 ( .A(P3_REG1_REG_29__SCAN_IN), .B(keyinput59), .ZN(n14281)
         );
  XNOR2_X1 U16158 ( .A(P1_REG1_REG_1__SCAN_IN), .B(keyinput39), .ZN(n14280) );
  NAND4_X1 U16159 ( .A1(n14283), .A2(n14282), .A3(n14281), .A4(n14280), .ZN(
        n14289) );
  XNOR2_X1 U16160 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput38), .ZN(n14287) );
  XNOR2_X1 U16161 ( .A(P3_IR_REG_16__SCAN_IN), .B(keyinput29), .ZN(n14286) );
  XNOR2_X1 U16162 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput53), .ZN(n14285)
         );
  XNOR2_X1 U16163 ( .A(keyinput28), .B(P1_REG0_REG_15__SCAN_IN), .ZN(n14284)
         );
  NAND4_X1 U16164 ( .A1(n14287), .A2(n14286), .A3(n14285), .A4(n14284), .ZN(
        n14288) );
  NOR2_X1 U16165 ( .A1(n14289), .A2(n14288), .ZN(n14297) );
  AOI22_X1 U16166 ( .A1(n14291), .A2(keyinput27), .B1(n7521), .B2(keyinput20), 
        .ZN(n14290) );
  OAI221_X1 U16167 ( .B1(n14291), .B2(keyinput27), .C1(n7521), .C2(keyinput20), 
        .A(n14290), .ZN(n14295) );
  AOI22_X1 U16168 ( .A1(n14481), .A2(keyinput12), .B1(n14293), .B2(keyinput49), 
        .ZN(n14292) );
  OAI221_X1 U16169 ( .B1(n14481), .B2(keyinput12), .C1(n14293), .C2(keyinput49), .A(n14292), .ZN(n14294) );
  NOR2_X1 U16170 ( .A1(n14295), .A2(n14294), .ZN(n14296) );
  AND3_X1 U16171 ( .A1(n14298), .A2(n14297), .A3(n14296), .ZN(n14299) );
  NAND4_X1 U16172 ( .A1(n14302), .A2(n14301), .A3(n14300), .A4(n14299), .ZN(
        n14303) );
  NOR2_X1 U16173 ( .A1(n14304), .A2(n14303), .ZN(n14333) );
  AOI22_X1 U16174 ( .A1(n14306), .A2(keyinput36), .B1(keyinput37), .B2(n14671), 
        .ZN(n14305) );
  OAI221_X1 U16175 ( .B1(n14306), .B2(keyinput36), .C1(n14671), .C2(keyinput37), .A(n14305), .ZN(n14318) );
  AOI22_X1 U16176 ( .A1(n14309), .A2(keyinput18), .B1(n14308), .B2(keyinput14), 
        .ZN(n14307) );
  OAI221_X1 U16177 ( .B1(n14309), .B2(keyinput18), .C1(n14308), .C2(keyinput14), .A(n14307), .ZN(n14317) );
  INV_X1 U16178 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n14494) );
  AOI22_X1 U16179 ( .A1(n14311), .A2(keyinput44), .B1(n14494), .B2(keyinput4), 
        .ZN(n14310) );
  OAI221_X1 U16180 ( .B1(n14311), .B2(keyinput44), .C1(n14494), .C2(keyinput4), 
        .A(n14310), .ZN(n14316) );
  INV_X1 U16181 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n14313) );
  AOI22_X1 U16182 ( .A1(n14314), .A2(keyinput32), .B1(keyinput63), .B2(n14313), 
        .ZN(n14312) );
  OAI221_X1 U16183 ( .B1(n14314), .B2(keyinput32), .C1(n14313), .C2(keyinput63), .A(n14312), .ZN(n14315) );
  NOR4_X1 U16184 ( .A1(n14318), .A2(n14317), .A3(n14316), .A4(n14315), .ZN(
        n14332) );
  AOI22_X1 U16185 ( .A1(n14320), .A2(keyinput40), .B1(keyinput11), .B2(n10331), 
        .ZN(n14319) );
  OAI221_X1 U16186 ( .B1(n14320), .B2(keyinput40), .C1(n10331), .C2(keyinput11), .A(n14319), .ZN(n14330) );
  AOI22_X1 U16187 ( .A1(n14322), .A2(keyinput17), .B1(keyinput0), .B2(n14492), 
        .ZN(n14321) );
  OAI221_X1 U16188 ( .B1(n14322), .B2(keyinput17), .C1(n14492), .C2(keyinput0), 
        .A(n14321), .ZN(n14329) );
  AOI22_X1 U16189 ( .A1(n15176), .A2(keyinput48), .B1(n14334), .B2(keyinput8), 
        .ZN(n14323) );
  OAI221_X1 U16190 ( .B1(n15176), .B2(keyinput48), .C1(n14334), .C2(keyinput8), 
        .A(n14323), .ZN(n14328) );
  AOI22_X1 U16191 ( .A1(n14326), .A2(keyinput21), .B1(keyinput22), .B2(n14325), 
        .ZN(n14324) );
  OAI221_X1 U16192 ( .B1(n14326), .B2(keyinput21), .C1(n14325), .C2(keyinput22), .A(n14324), .ZN(n14327) );
  NOR4_X1 U16193 ( .A1(n14330), .A2(n14329), .A3(n14328), .A4(n14327), .ZN(
        n14331) );
  NAND3_X1 U16194 ( .A1(n14333), .A2(n14332), .A3(n14331), .ZN(n14363) );
  NOR4_X1 U16195 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_REG0_REG_15__SCAN_IN), 
        .A3(P3_REG1_REG_14__SCAN_IN), .A4(P3_REG0_REG_14__SCAN_IN), .ZN(n14348) );
  NAND4_X1 U16196 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_REG1_REG_21__SCAN_IN), 
        .A3(P3_REG0_REG_23__SCAN_IN), .A4(P1_REG3_REG_0__SCAN_IN), .ZN(n14342)
         );
  NAND3_X1 U16197 ( .A1(SI_10_), .A2(SI_0_), .A3(P1_IR_REG_18__SCAN_IN), .ZN(
        n14341) );
  NAND3_X1 U16198 ( .A1(P3_REG1_REG_29__SCAN_IN), .A2(n14335), .A3(n14334), 
        .ZN(n14339) );
  NAND4_X1 U16199 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_REG0_REG_9__SCAN_IN), 
        .A3(P2_REG0_REG_3__SCAN_IN), .A4(P1_REG0_REG_24__SCAN_IN), .ZN(n14338)
         );
  NAND4_X1 U16200 ( .A1(P2_REG0_REG_13__SCAN_IN), .A2(P1_REG2_REG_18__SCAN_IN), 
        .A3(P1_REG0_REG_11__SCAN_IN), .A4(P1_REG0_REG_2__SCAN_IN), .ZN(n14337)
         );
  NAND4_X1 U16201 ( .A1(P2_REG2_REG_23__SCAN_IN), .A2(P3_REG0_REG_15__SCAN_IN), 
        .A3(P1_REG3_REG_14__SCAN_IN), .A4(P1_REG1_REG_1__SCAN_IN), .ZN(n14336)
         );
  OR4_X1 U16202 ( .A1(n14339), .A2(n14338), .A3(n14337), .A4(n14336), .ZN(
        n14340) );
  NOR4_X1 U16203 ( .A1(P3_REG2_REG_24__SCAN_IN), .A2(n14342), .A3(n14341), 
        .A4(n14340), .ZN(n14347) );
  NAND4_X1 U16204 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_D_REG_31__SCAN_IN), .A3(
        P3_REG1_REG_25__SCAN_IN), .A4(P3_REG3_REG_0__SCAN_IN), .ZN(n14344) );
  NAND4_X1 U16205 ( .A1(P3_REG3_REG_25__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .A3(P3_DATAO_REG_20__SCAN_IN), .A4(P3_DATAO_REG_30__SCAN_IN), .ZN(
        n14343) );
  NOR2_X1 U16206 ( .A1(n14344), .A2(n14343), .ZN(n14346) );
  NAND4_X1 U16207 ( .A1(n14348), .A2(n14347), .A3(n14346), .A4(n14345), .ZN(
        n14361) );
  NOR3_X1 U16208 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(P3_ADDR_REG_6__SCAN_IN), 
        .A3(n14349), .ZN(n14354) );
  NOR4_X1 U16209 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(P2_DATAO_REG_28__SCAN_IN), .A3(n14351), .A4(n14350), .ZN(n14353) );
  NOR4_X1 U16210 ( .A1(P3_REG0_REG_30__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .A3(P1_REG3_REG_6__SCAN_IN), .A4(P3_DATAO_REG_9__SCAN_IN), .ZN(n14352)
         );
  NAND4_X1 U16211 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14354), .A3(n14353), 
        .A4(n14352), .ZN(n14360) );
  NOR4_X1 U16212 ( .A1(P3_D_REG_22__SCAN_IN), .A2(P3_REG3_REG_12__SCAN_IN), 
        .A3(P3_REG1_REG_3__SCAN_IN), .A4(P3_DATAO_REG_13__SCAN_IN), .ZN(n14358) );
  NOR4_X1 U16213 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        P3_REG2_REG_3__SCAN_IN), .A4(P3_REG2_REG_1__SCAN_IN), .ZN(n14357) );
  NOR4_X1 U16214 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_REG2_REG_8__SCAN_IN), 
        .A3(P2_REG2_REG_6__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n14356) );
  NOR4_X1 U16215 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(P1_REG2_REG_4__SCAN_IN), 
        .A3(P3_ADDR_REG_12__SCAN_IN), .A4(P2_ADDR_REG_12__SCAN_IN), .ZN(n14355) );
  NAND4_X1 U16216 ( .A1(n14358), .A2(n14357), .A3(n14356), .A4(n14355), .ZN(
        n14359) );
  NOR3_X1 U16217 ( .A1(n14361), .A2(n14360), .A3(n14359), .ZN(n14362) );
  XNOR2_X1 U16218 ( .A(n14363), .B(n14362), .ZN(n14364) );
  XNOR2_X1 U16219 ( .A(n14365), .B(n14364), .ZN(P1_U3324) );
  OAI222_X1 U16220 ( .A1(n14375), .A2(n14368), .B1(n14367), .B2(P1_U3086), 
        .C1(n14366), .C2(n14372), .ZN(P1_U3325) );
  OAI222_X1 U16221 ( .A1(n14375), .A2(n14371), .B1(n14370), .B2(P1_U3086), 
        .C1(n14369), .C2(n14372), .ZN(P1_U3326) );
  OAI222_X1 U16222 ( .A1(n6453), .A2(P1_U3086), .B1(n14375), .B2(n14374), .C1(
        n14373), .C2(n14372), .ZN(P1_U3328) );
  MUX2_X1 U16223 ( .A(n11840), .B(n14376), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16224 ( .A(n6602), .B(n14377), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3355) );
  AOI21_X1 U16225 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14380) );
  OAI21_X1 U16226 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14380), 
        .ZN(U28) );
  AOI21_X1 U16227 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14381) );
  OAI21_X1 U16228 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14381), 
        .ZN(U29) );
  OAI21_X1 U16229 ( .B1(n14384), .B2(n14383), .A(n14382), .ZN(n14385) );
  XNOR2_X1 U16230 ( .A(n14385), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  AOI21_X1 U16231 ( .B1(n14388), .B2(n14387), .A(n14386), .ZN(SUB_1596_U57) );
  OAI21_X1 U16232 ( .B1(n14391), .B2(n14390), .A(n14389), .ZN(SUB_1596_U55) );
  OAI21_X1 U16233 ( .B1(n14394), .B2(n14393), .A(n14392), .ZN(SUB_1596_U54) );
  OAI222_X1 U16234 ( .A1(n14399), .A2(n14398), .B1(n14399), .B2(n14397), .C1(
        n14396), .C2(n14395), .ZN(SUB_1596_U70) );
  OAI21_X1 U16235 ( .B1(n14402), .B2(n14401), .A(n14400), .ZN(SUB_1596_U63) );
  AOI21_X1 U16236 ( .B1(n14405), .B2(n14404), .A(n14403), .ZN(n14420) );
  OAI21_X1 U16237 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n14407), .A(n14406), 
        .ZN(n14413) );
  NOR2_X1 U16238 ( .A1(n15101), .A2(n14408), .ZN(n14412) );
  OAI21_X1 U16239 ( .B1(n15104), .B2(n14410), .A(n14409), .ZN(n14411) );
  AOI211_X1 U16240 ( .C1(n14413), .C2(n15107), .A(n14412), .B(n14411), .ZN(
        n14419) );
  NOR2_X1 U16241 ( .A1(n14415), .A2(n14414), .ZN(n14416) );
  OAI21_X1 U16242 ( .B1(n14417), .B2(n14416), .A(n15090), .ZN(n14418) );
  OAI211_X1 U16243 ( .C1(n14420), .C2(n15116), .A(n14419), .B(n14418), .ZN(
        P3_U3197) );
  AOI22_X1 U16244 ( .A1(n15000), .A2(n14421), .B1(n15082), .B2(
        P3_ADDR_REG_16__SCAN_IN), .ZN(n14437) );
  INV_X1 U16245 ( .A(n14422), .ZN(n14423) );
  NAND2_X1 U16246 ( .A1(n14424), .A2(n14423), .ZN(n14425) );
  XNOR2_X1 U16247 ( .A(n14426), .B(n14425), .ZN(n14431) );
  OAI21_X1 U16248 ( .B1(n14429), .B2(n14428), .A(n14427), .ZN(n14430) );
  AOI22_X1 U16249 ( .A1(n14431), .A2(n15090), .B1(n15107), .B2(n14430), .ZN(
        n14436) );
  NAND2_X1 U16250 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P3_U3151), .ZN(n14435)
         );
  OAI221_X1 U16251 ( .B1(n14433), .B2(n6530), .C1(n14433), .C2(n14432), .A(
        n14960), .ZN(n14434) );
  NAND4_X1 U16252 ( .A1(n14437), .A2(n14436), .A3(n14435), .A4(n14434), .ZN(
        P3_U3198) );
  AOI22_X1 U16253 ( .A1(n15000), .A2(n14438), .B1(n15082), .B2(
        P3_ADDR_REG_17__SCAN_IN), .ZN(n14453) );
  OAI21_X1 U16254 ( .B1(P3_REG1_REG_17__SCAN_IN), .B2(n14440), .A(n14439), 
        .ZN(n14445) );
  AOI211_X1 U16255 ( .C1(n14443), .C2(n14442), .A(n14441), .B(n15109), .ZN(
        n14444) );
  AOI21_X1 U16256 ( .B1(n15107), .B2(n14445), .A(n14444), .ZN(n14452) );
  INV_X1 U16257 ( .A(n14446), .ZN(n14451) );
  OAI221_X1 U16258 ( .B1(n14449), .B2(n14448), .C1(n14449), .C2(n14447), .A(
        n14960), .ZN(n14450) );
  NAND4_X1 U16259 ( .A1(n14453), .A2(n14452), .A3(n14451), .A4(n14450), .ZN(
        P3_U3199) );
  AOI22_X1 U16260 ( .A1(n15000), .A2(n14454), .B1(n15082), .B2(
        P3_ADDR_REG_18__SCAN_IN), .ZN(n14470) );
  XNOR2_X1 U16261 ( .A(n14456), .B(n14455), .ZN(n14462) );
  AOI21_X1 U16262 ( .B1(n14459), .B2(n14458), .A(n14457), .ZN(n14460) );
  NOR2_X1 U16263 ( .A1(n14460), .A2(n15109), .ZN(n14461) );
  AOI21_X1 U16264 ( .B1(n14462), .B2(n15107), .A(n14461), .ZN(n14469) );
  INV_X1 U16265 ( .A(n14463), .ZN(n14468) );
  NAND4_X1 U16266 ( .A1(n14470), .A2(n14469), .A3(n14468), .A4(n14467), .ZN(
        P3_U3200) );
  AOI22_X1 U16267 ( .A1(n14475), .A2(n14471), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n15136), .ZN(n14472) );
  NAND2_X1 U16268 ( .A1(n14473), .A2(n14472), .ZN(P3_U3203) );
  AOI21_X1 U16269 ( .B1(n14475), .B2(n15152), .A(n14474), .ZN(n14493) );
  INV_X1 U16270 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14476) );
  AOI22_X1 U16271 ( .A1(n15166), .A2(n14493), .B1(n14476), .B2(n15164), .ZN(
        P3_U3489) );
  OAI22_X1 U16272 ( .A1(n14478), .A2(n14483), .B1(n14477), .B2(n15144), .ZN(
        n14479) );
  NOR2_X1 U16273 ( .A1(n14480), .A2(n14479), .ZN(n14495) );
  AOI22_X1 U16274 ( .A1(n15166), .A2(n14495), .B1(n14481), .B2(n15164), .ZN(
        P3_U3473) );
  OAI22_X1 U16275 ( .A1(n14484), .A2(n14483), .B1(n14482), .B2(n15144), .ZN(
        n14485) );
  NOR2_X1 U16276 ( .A1(n14486), .A2(n14485), .ZN(n14497) );
  AOI22_X1 U16277 ( .A1(n15166), .A2(n14497), .B1(n8916), .B2(n15164), .ZN(
        P3_U3472) );
  AOI22_X1 U16278 ( .A1(n14488), .A2(n15150), .B1(n15152), .B2(n14487), .ZN(
        n14489) );
  AOI22_X1 U16279 ( .A1(n15166), .A2(n14498), .B1(n14491), .B2(n15164), .ZN(
        P3_U3471) );
  AOI22_X1 U16280 ( .A1(n15158), .A2(n14493), .B1(n14492), .B2(n15157), .ZN(
        P3_U3457) );
  AOI22_X1 U16281 ( .A1(n15158), .A2(n14495), .B1(n14494), .B2(n15157), .ZN(
        P3_U3432) );
  INV_X1 U16282 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14496) );
  AOI22_X1 U16283 ( .A1(n15158), .A2(n14497), .B1(n14496), .B2(n15157), .ZN(
        P3_U3429) );
  AOI22_X1 U16284 ( .A1(n15158), .A2(n14498), .B1(n8895), .B2(n15157), .ZN(
        P3_U3426) );
  OAI22_X1 U16285 ( .A1(n14499), .A2(n14519), .B1(n14518), .B2(n14520), .ZN(
        n14506) );
  NAND2_X1 U16286 ( .A1(n14501), .A2(n14500), .ZN(n14503) );
  AOI21_X1 U16287 ( .B1(n14504), .B2(n14503), .A(n14502), .ZN(n14505) );
  AOI211_X1 U16288 ( .C1(n14508), .C2(n14507), .A(n14506), .B(n14505), .ZN(
        n14510) );
  OAI211_X1 U16289 ( .C1(n14528), .C2(n14511), .A(n14510), .B(n14509), .ZN(
        P2_U3187) );
  OAI21_X1 U16290 ( .B1(n14514), .B2(n14513), .A(n14512), .ZN(n14524) );
  NOR2_X1 U16291 ( .A1(n14516), .A2(n14515), .ZN(n14522) );
  OAI22_X1 U16292 ( .A1(n14520), .A2(n14519), .B1(n14518), .B2(n14517), .ZN(
        n14521) );
  AOI211_X1 U16293 ( .C1(n14524), .C2(n14523), .A(n14522), .B(n14521), .ZN(
        n14526) );
  OAI211_X1 U16294 ( .C1(n14528), .C2(n14527), .A(n14526), .B(n14525), .ZN(
        P2_U3198) );
  OAI21_X1 U16295 ( .B1(n14530), .B2(n14922), .A(n14529), .ZN(n14532) );
  AOI211_X1 U16296 ( .C1(n14534), .C2(n14533), .A(n14532), .B(n14531), .ZN(
        n14535) );
  AOI22_X1 U16297 ( .A1(n14933), .A2(n14535), .B1(n11113), .B2(n14931), .ZN(
        P2_U3512) );
  AOI22_X1 U16298 ( .A1(n6443), .A2(n14535), .B1(n7806), .B2(n14928), .ZN(
        P2_U3469) );
  OAI211_X1 U16299 ( .C1(n14538), .C2(n14821), .A(n14537), .B(n14536), .ZN(
        n14539) );
  AOI211_X1 U16300 ( .C1(n14541), .C2(n14824), .A(n14540), .B(n14539), .ZN(
        n14553) );
  AOI22_X1 U16301 ( .A1(n14839), .A2(n14553), .B1(n14629), .B2(n14837), .ZN(
        P1_U3543) );
  OAI211_X1 U16302 ( .C1(n14544), .C2(n14821), .A(n14543), .B(n14542), .ZN(
        n14545) );
  AOI211_X1 U16303 ( .C1(n14547), .C2(n14824), .A(n14546), .B(n14545), .ZN(
        n14554) );
  AOI22_X1 U16304 ( .A1(n14839), .A2(n14554), .B1(n13780), .B2(n14837), .ZN(
        P1_U3541) );
  OAI21_X1 U16305 ( .B1(n14549), .B2(n14821), .A(n14548), .ZN(n14550) );
  AOI211_X1 U16306 ( .C1(n14552), .C2(n14824), .A(n14551), .B(n14550), .ZN(
        n14555) );
  AOI22_X1 U16307 ( .A1(n14839), .A2(n14555), .B1(n10851), .B2(n14837), .ZN(
        P1_U3539) );
  AOI22_X1 U16308 ( .A1(n14827), .A2(n14553), .B1(n11290), .B2(n14826), .ZN(
        P1_U3504) );
  AOI22_X1 U16309 ( .A1(n14827), .A2(n14554), .B1(n11010), .B2(n14826), .ZN(
        P1_U3498) );
  AOI22_X1 U16310 ( .A1(n14827), .A2(n14555), .B1(n10854), .B2(n14826), .ZN(
        P1_U3492) );
  OAI21_X1 U16311 ( .B1(n14558), .B2(n14557), .A(n14556), .ZN(n14559) );
  XNOR2_X1 U16312 ( .A(n14559), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  OAI21_X1 U16313 ( .B1(n14562), .B2(n14561), .A(n14560), .ZN(n14563) );
  XNOR2_X1 U16314 ( .A(n14563), .B(P2_ADDR_REG_12__SCAN_IN), .ZN(SUB_1596_U68)
         );
  OAI222_X1 U16315 ( .A1(n14870), .A2(n14567), .B1(n14870), .B2(n14566), .C1(
        n14565), .C2(n14564), .ZN(SUB_1596_U67) );
  OAI21_X1 U16316 ( .B1(n14570), .B2(n14569), .A(n14568), .ZN(n14571) );
  XNOR2_X1 U16317 ( .A(n14571), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  OAI222_X1 U16318 ( .A1(n14576), .A2(n14575), .B1(n14576), .B2(n14574), .C1(
        n14573), .C2(n14572), .ZN(SUB_1596_U65) );
  OAI21_X1 U16319 ( .B1(n14579), .B2(n14578), .A(n14577), .ZN(n14580) );
  XNOR2_X1 U16320 ( .A(n14580), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  OAI21_X1 U16321 ( .B1(n14582), .B2(P1_REG1_REG_0__SCAN_IN), .A(n14581), .ZN(
        n14584) );
  XNOR2_X1 U16322 ( .A(n14584), .B(n14583), .ZN(n14588) );
  AOI22_X1 U16323 ( .A1(n14585), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14586) );
  OAI21_X1 U16324 ( .B1(n14588), .B2(n14587), .A(n14586), .ZN(P1_U3243) );
  AOI211_X1 U16325 ( .C1(n14591), .C2(n14590), .A(n14669), .B(n14589), .ZN(
        n14596) );
  AOI211_X1 U16326 ( .C1(n14594), .C2(n14593), .A(n14665), .B(n14592), .ZN(
        n14595) );
  AOI211_X1 U16327 ( .C1(n14676), .C2(n14597), .A(n14596), .B(n14595), .ZN(
        n14600) );
  INV_X1 U16328 ( .A(n14598), .ZN(n14599) );
  OAI211_X1 U16329 ( .C1(n14601), .C2(n14679), .A(n14600), .B(n14599), .ZN(
        P1_U3253) );
  AOI211_X1 U16330 ( .C1(n14604), .C2(n14603), .A(n14602), .B(n14669), .ZN(
        n14609) );
  AOI211_X1 U16331 ( .C1(n14607), .C2(n14606), .A(n14605), .B(n14665), .ZN(
        n14608) );
  AOI211_X1 U16332 ( .C1(n14676), .C2(n14610), .A(n14609), .B(n14608), .ZN(
        n14612) );
  OAI211_X1 U16333 ( .C1(n14613), .C2(n14679), .A(n14612), .B(n14611), .ZN(
        P1_U3256) );
  OAI21_X1 U16334 ( .B1(n14616), .B2(n14615), .A(n14614), .ZN(n14624) );
  NOR2_X1 U16335 ( .A1(n14618), .A2(n14617), .ZN(n14623) );
  AOI211_X1 U16336 ( .C1(n14621), .C2(n14620), .A(n14619), .B(n14669), .ZN(
        n14622) );
  AOI211_X1 U16337 ( .C1(n14636), .C2(n14624), .A(n14623), .B(n14622), .ZN(
        n14626) );
  OAI211_X1 U16338 ( .C1(n14627), .C2(n14679), .A(n14626), .B(n14625), .ZN(
        P1_U3257) );
  OAI21_X1 U16339 ( .B1(n14630), .B2(n14629), .A(n14628), .ZN(n14637) );
  OAI21_X1 U16340 ( .B1(n14632), .B2(n11296), .A(n14631), .ZN(n14634) );
  AOI222_X1 U16341 ( .A1(n14637), .A2(n14636), .B1(n14635), .B2(n14676), .C1(
        n14634), .C2(n14633), .ZN(n14639) );
  OAI211_X1 U16342 ( .C1(n14640), .C2(n14679), .A(n14639), .B(n14638), .ZN(
        P1_U3258) );
  AOI211_X1 U16343 ( .C1(n14643), .C2(n14642), .A(n14665), .B(n14641), .ZN(
        n14648) );
  AOI211_X1 U16344 ( .C1(n14646), .C2(n14645), .A(n14669), .B(n14644), .ZN(
        n14647) );
  AOI211_X1 U16345 ( .C1(n14676), .C2(n14649), .A(n14648), .B(n14647), .ZN(
        n14651) );
  OAI211_X1 U16346 ( .C1(n14652), .C2(n14679), .A(n14651), .B(n14650), .ZN(
        P1_U3259) );
  INV_X1 U16347 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14664) );
  AOI211_X1 U16348 ( .C1(n14655), .C2(n14654), .A(n14653), .B(n14669), .ZN(
        n14660) );
  AOI211_X1 U16349 ( .C1(n14658), .C2(n14657), .A(n14665), .B(n14656), .ZN(
        n14659) );
  AOI211_X1 U16350 ( .C1(n14676), .C2(n14661), .A(n14660), .B(n14659), .ZN(
        n14663) );
  OAI211_X1 U16351 ( .C1(n14664), .C2(n14679), .A(n14663), .B(n14662), .ZN(
        P1_U3260) );
  AOI211_X1 U16352 ( .C1(n14668), .C2(n14667), .A(n14666), .B(n14665), .ZN(
        n14674) );
  AOI211_X1 U16353 ( .C1(n14672), .C2(n14671), .A(n14670), .B(n14669), .ZN(
        n14673) );
  AOI211_X1 U16354 ( .C1(n14676), .C2(n14675), .A(n14674), .B(n14673), .ZN(
        n14678) );
  OAI211_X1 U16355 ( .C1(n14680), .C2(n14679), .A(n14678), .B(n14677), .ZN(
        P1_U3261) );
  XNOR2_X1 U16356 ( .A(n14681), .B(n14686), .ZN(n14684) );
  AOI222_X1 U16357 ( .A1(n14685), .A2(n14684), .B1(n14683), .B2(n14702), .C1(
        n14682), .C2(n14705), .ZN(n14809) );
  XNOR2_X1 U16358 ( .A(n14687), .B(n14686), .ZN(n14811) );
  INV_X1 U16359 ( .A(n14688), .ZN(n14689) );
  OAI211_X1 U16360 ( .C1(n10753), .C2(n14714), .A(n14689), .B(n14756), .ZN(
        n14807) );
  OAI22_X1 U16361 ( .A1(n14691), .A2(n9748), .B1(n14690), .B2(n14751), .ZN(
        n14692) );
  AOI21_X1 U16362 ( .B1(n14693), .B2(n14754), .A(n14692), .ZN(n14694) );
  OAI21_X1 U16363 ( .B1(n14807), .B2(n14695), .A(n14694), .ZN(n14696) );
  AOI21_X1 U16364 ( .B1(n14811), .B2(n14697), .A(n14696), .ZN(n14698) );
  OAI21_X1 U16365 ( .B1(n6442), .B2(n14809), .A(n14698), .ZN(P1_U3285) );
  XNOR2_X1 U16366 ( .A(n14699), .B(n14700), .ZN(n14804) );
  XNOR2_X1 U16367 ( .A(n14701), .B(n14700), .ZN(n14707) );
  AOI22_X1 U16368 ( .A1(n14705), .A2(n14704), .B1(n14703), .B2(n14702), .ZN(
        n14706) );
  OAI21_X1 U16369 ( .B1(n14707), .B2(n14744), .A(n14706), .ZN(n14708) );
  AOI21_X1 U16370 ( .B1(n14804), .B2(n14749), .A(n14708), .ZN(n14801) );
  INV_X1 U16371 ( .A(n14709), .ZN(n14711) );
  AOI222_X1 U16372 ( .A1(n14712), .A2(n14754), .B1(n14711), .B2(n14710), .C1(
        P1_REG2_REG_7__SCAN_IN), .C2(n6442), .ZN(n14718) );
  INV_X1 U16373 ( .A(n14713), .ZN(n14715) );
  OAI211_X1 U16374 ( .C1(n14800), .C2(n14715), .A(n6958), .B(n14756), .ZN(
        n14799) );
  INV_X1 U16375 ( .A(n14799), .ZN(n14716) );
  AOI22_X1 U16376 ( .A1(n14804), .A2(n14760), .B1(n14759), .B2(n14716), .ZN(
        n14717) );
  OAI211_X1 U16377 ( .C1(n6442), .C2(n14801), .A(n14718), .B(n14717), .ZN(
        P1_U3286) );
  XNOR2_X1 U16378 ( .A(n14719), .B(n14724), .ZN(n14789) );
  OAI22_X1 U16379 ( .A1(n14723), .A2(n14722), .B1(n14721), .B2(n14720), .ZN(
        n14730) );
  NAND3_X1 U16380 ( .A1(n14726), .A2(n14725), .A3(n14724), .ZN(n14727) );
  AOI21_X1 U16381 ( .B1(n14728), .B2(n14727), .A(n14744), .ZN(n14729) );
  AOI211_X1 U16382 ( .C1(n14749), .C2(n14789), .A(n14730), .B(n14729), .ZN(
        n14786) );
  NAND2_X1 U16383 ( .A1(n6442), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n14731) );
  OAI21_X1 U16384 ( .B1(n14751), .B2(n14732), .A(n14731), .ZN(n14733) );
  AOI21_X1 U16385 ( .B1(n14754), .B2(n14734), .A(n14733), .ZN(n14739) );
  OAI211_X1 U16386 ( .C1(n14736), .C2(n14785), .A(n14735), .B(n14756), .ZN(
        n14784) );
  INV_X1 U16387 ( .A(n14784), .ZN(n14737) );
  AOI22_X1 U16388 ( .A1(n14789), .A2(n14760), .B1(n14759), .B2(n14737), .ZN(
        n14738) );
  OAI211_X1 U16389 ( .C1(n6442), .C2(n14786), .A(n14739), .B(n14738), .ZN(
        P1_U3288) );
  XNOR2_X1 U16390 ( .A(n14740), .B(n14742), .ZN(n14777) );
  NAND3_X1 U16391 ( .A1(n14743), .A2(n14742), .A3(n14741), .ZN(n14745) );
  AOI21_X1 U16392 ( .B1(n14746), .B2(n14745), .A(n14744), .ZN(n14747) );
  AOI211_X1 U16393 ( .C1(n14749), .C2(n14777), .A(n14748), .B(n14747), .ZN(
        n14774) );
  NAND2_X1 U16394 ( .A1(n6442), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n14750) );
  OAI21_X1 U16395 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(n14751), .A(n14750), .ZN(
        n14752) );
  AOI21_X1 U16396 ( .B1(n14754), .B2(n14753), .A(n14752), .ZN(n14762) );
  OAI211_X1 U16397 ( .C1(n14757), .C2(n14773), .A(n14756), .B(n14755), .ZN(
        n14772) );
  INV_X1 U16398 ( .A(n14772), .ZN(n14758) );
  AOI22_X1 U16399 ( .A1(n14777), .A2(n14760), .B1(n14759), .B2(n14758), .ZN(
        n14761) );
  OAI211_X1 U16400 ( .C1(n6442), .C2(n14774), .A(n14762), .B(n14761), .ZN(
        P1_U3290) );
  AND2_X1 U16401 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14765), .ZN(P1_U3294) );
  AND2_X1 U16402 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14765), .ZN(P1_U3295) );
  AND2_X1 U16403 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14765), .ZN(P1_U3296) );
  AND2_X1 U16404 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14765), .ZN(P1_U3297) );
  AND2_X1 U16405 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14765), .ZN(P1_U3298) );
  AND2_X1 U16406 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14765), .ZN(P1_U3299) );
  AND2_X1 U16407 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14765), .ZN(P1_U3300) );
  AND2_X1 U16408 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14765), .ZN(P1_U3301) );
  AND2_X1 U16409 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14765), .ZN(P1_U3302) );
  AND2_X1 U16410 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14765), .ZN(P1_U3303) );
  AND2_X1 U16411 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14765), .ZN(P1_U3304) );
  AND2_X1 U16412 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14765), .ZN(P1_U3305) );
  AND2_X1 U16413 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14765), .ZN(P1_U3306) );
  AND2_X1 U16414 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14765), .ZN(P1_U3307) );
  AND2_X1 U16415 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14765), .ZN(P1_U3308) );
  AND2_X1 U16416 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14765), .ZN(P1_U3309) );
  AND2_X1 U16417 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14765), .ZN(P1_U3310) );
  AND2_X1 U16418 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14765), .ZN(P1_U3311) );
  AND2_X1 U16419 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14765), .ZN(P1_U3312) );
  AND2_X1 U16420 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14765), .ZN(P1_U3313) );
  AND2_X1 U16421 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14765), .ZN(P1_U3314) );
  AND2_X1 U16422 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14765), .ZN(P1_U3315) );
  AND2_X1 U16423 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14765), .ZN(P1_U3316) );
  AND2_X1 U16424 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14765), .ZN(P1_U3317) );
  AND2_X1 U16425 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14765), .ZN(P1_U3318) );
  NOR2_X1 U16426 ( .A1(n14764), .A2(n14763), .ZN(P1_U3319) );
  AND2_X1 U16427 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14765), .ZN(P1_U3320) );
  AND2_X1 U16428 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14765), .ZN(P1_U3321) );
  AND2_X1 U16429 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14765), .ZN(P1_U3322) );
  AND2_X1 U16430 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14765), .ZN(P1_U3323) );
  AOI22_X1 U16431 ( .A1(n14827), .A2(n14766), .B1(n9518), .B2(n14826), .ZN(
        P1_U3462) );
  OAI211_X1 U16432 ( .C1(n14769), .C2(n14797), .A(n14768), .B(n14767), .ZN(
        n14770) );
  NOR2_X1 U16433 ( .A1(n14771), .A2(n14770), .ZN(n14828) );
  AOI22_X1 U16434 ( .A1(n14827), .A2(n14828), .B1(n9606), .B2(n14826), .ZN(
        P1_U3465) );
  OAI21_X1 U16435 ( .B1(n14773), .B2(n14821), .A(n14772), .ZN(n14776) );
  INV_X1 U16436 ( .A(n14774), .ZN(n14775) );
  AOI211_X1 U16437 ( .C1(n14805), .C2(n14777), .A(n14776), .B(n14775), .ZN(
        n14829) );
  INV_X1 U16438 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14778) );
  AOI22_X1 U16439 ( .A1(n14827), .A2(n14829), .B1(n14778), .B2(n14826), .ZN(
        P1_U3468) );
  OAI211_X1 U16440 ( .C1(n14781), .C2(n14821), .A(n14780), .B(n14779), .ZN(
        n14782) );
  AOI21_X1 U16441 ( .B1(n14824), .B2(n14783), .A(n14782), .ZN(n14831) );
  AOI22_X1 U16442 ( .A1(n14827), .A2(n14831), .B1(n10130), .B2(n14826), .ZN(
        P1_U3471) );
  OAI21_X1 U16443 ( .B1(n14785), .B2(n14821), .A(n14784), .ZN(n14788) );
  INV_X1 U16444 ( .A(n14786), .ZN(n14787) );
  AOI211_X1 U16445 ( .C1(n14805), .C2(n14789), .A(n14788), .B(n14787), .ZN(
        n14832) );
  INV_X1 U16446 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14790) );
  AOI22_X1 U16447 ( .A1(n14827), .A2(n14832), .B1(n14790), .B2(n14826), .ZN(
        P1_U3474) );
  AOI21_X1 U16448 ( .B1(n14793), .B2(n14792), .A(n14791), .ZN(n14794) );
  OAI211_X1 U16449 ( .C1(n14797), .C2(n14796), .A(n14795), .B(n14794), .ZN(
        n14798) );
  INV_X1 U16450 ( .A(n14798), .ZN(n14833) );
  AOI22_X1 U16451 ( .A1(n14827), .A2(n14833), .B1(n10235), .B2(n14826), .ZN(
        P1_U3477) );
  OAI21_X1 U16452 ( .B1(n14800), .B2(n14821), .A(n14799), .ZN(n14803) );
  INV_X1 U16453 ( .A(n14801), .ZN(n14802) );
  AOI211_X1 U16454 ( .C1(n14805), .C2(n14804), .A(n14803), .B(n14802), .ZN(
        n14834) );
  AOI22_X1 U16455 ( .A1(n14827), .A2(n14834), .B1(n10335), .B2(n14826), .ZN(
        P1_U3480) );
  INV_X1 U16456 ( .A(n14806), .ZN(n14808) );
  NAND3_X1 U16457 ( .A1(n14809), .A2(n14808), .A3(n14807), .ZN(n14810) );
  AOI21_X1 U16458 ( .B1(n14811), .B2(n14824), .A(n14810), .ZN(n14835) );
  INV_X1 U16459 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14812) );
  AOI22_X1 U16460 ( .A1(n14827), .A2(n14835), .B1(n14812), .B2(n14826), .ZN(
        P1_U3483) );
  INV_X1 U16461 ( .A(n14813), .ZN(n14818) );
  OAI21_X1 U16462 ( .B1(n14815), .B2(n14821), .A(n14814), .ZN(n14817) );
  AOI211_X1 U16463 ( .C1(n14824), .C2(n14818), .A(n14817), .B(n14816), .ZN(
        n14836) );
  AOI22_X1 U16464 ( .A1(n14827), .A2(n14836), .B1(n10734), .B2(n14826), .ZN(
        P1_U3486) );
  OAI211_X1 U16465 ( .C1(n14822), .C2(n14821), .A(n14820), .B(n14819), .ZN(
        n14823) );
  AOI21_X1 U16466 ( .B1(n14825), .B2(n14824), .A(n14823), .ZN(n14838) );
  AOI22_X1 U16467 ( .A1(n14827), .A2(n14838), .B1(n10761), .B2(n14826), .ZN(
        P1_U3489) );
  AOI22_X1 U16468 ( .A1(n14839), .A2(n14828), .B1(n9607), .B2(n14837), .ZN(
        P1_U3530) );
  AOI22_X1 U16469 ( .A1(n14839), .A2(n14829), .B1(n9773), .B2(n14837), .ZN(
        P1_U3531) );
  INV_X1 U16470 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n14830) );
  AOI22_X1 U16471 ( .A1(n14839), .A2(n14831), .B1(n14830), .B2(n14837), .ZN(
        P1_U3532) );
  AOI22_X1 U16472 ( .A1(n14839), .A2(n14832), .B1(n10169), .B2(n14837), .ZN(
        P1_U3533) );
  AOI22_X1 U16473 ( .A1(n14839), .A2(n14833), .B1(n9481), .B2(n14837), .ZN(
        P1_U3534) );
  AOI22_X1 U16474 ( .A1(n14839), .A2(n14834), .B1(n9742), .B2(n14837), .ZN(
        P1_U3535) );
  AOI22_X1 U16475 ( .A1(n14839), .A2(n14835), .B1(n10573), .B2(n14837), .ZN(
        P1_U3536) );
  AOI22_X1 U16476 ( .A1(n14839), .A2(n14836), .B1(n10729), .B2(n14837), .ZN(
        P1_U3537) );
  AOI22_X1 U16477 ( .A1(n14839), .A2(n14838), .B1(n10349), .B2(n14837), .ZN(
        P1_U3538) );
  NOR2_X1 U16478 ( .A1(n14840), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI211_X1 U16479 ( .C1(n14843), .C2(n14842), .A(n14841), .B(n14856), .ZN(
        n14844) );
  AOI211_X1 U16480 ( .C1(n14862), .C2(n14846), .A(n14845), .B(n14844), .ZN(
        n14852) );
  AOI211_X1 U16481 ( .C1(n14849), .C2(n14848), .A(n14847), .B(n14864), .ZN(
        n14850) );
  INV_X1 U16482 ( .A(n14850), .ZN(n14851) );
  OAI211_X1 U16483 ( .C1(n14871), .C2(n14853), .A(n14852), .B(n14851), .ZN(
        P2_U3218) );
  NOR2_X1 U16484 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14854), .ZN(n14860) );
  AOI211_X1 U16485 ( .C1(n14858), .C2(n14857), .A(n14856), .B(n14855), .ZN(
        n14859) );
  AOI211_X1 U16486 ( .C1(n14862), .C2(n14861), .A(n14860), .B(n14859), .ZN(
        n14869) );
  AOI211_X1 U16487 ( .C1(n14866), .C2(n14865), .A(n14864), .B(n14863), .ZN(
        n14867) );
  INV_X1 U16488 ( .A(n14867), .ZN(n14868) );
  OAI211_X1 U16489 ( .C1(n14871), .C2(n14870), .A(n14869), .B(n14868), .ZN(
        P2_U3227) );
  INV_X1 U16490 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n14874) );
  NOR2_X1 U16491 ( .A1(n14910), .A2(n14874), .ZN(P2_U3266) );
  INV_X1 U16492 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n14875) );
  NOR2_X1 U16493 ( .A1(n14910), .A2(n14875), .ZN(P2_U3267) );
  NOR2_X1 U16494 ( .A1(n14910), .A2(n14876), .ZN(P2_U3268) );
  INV_X1 U16495 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n14877) );
  NOR2_X1 U16496 ( .A1(n14910), .A2(n14877), .ZN(P2_U3269) );
  INV_X1 U16497 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n14878) );
  NOR2_X1 U16498 ( .A1(n14888), .A2(n14878), .ZN(P2_U3270) );
  INV_X1 U16499 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n14879) );
  NOR2_X1 U16500 ( .A1(n14888), .A2(n14879), .ZN(P2_U3271) );
  INV_X1 U16501 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n14880) );
  NOR2_X1 U16502 ( .A1(n14888), .A2(n14880), .ZN(P2_U3272) );
  INV_X1 U16503 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n14881) );
  NOR2_X1 U16504 ( .A1(n14888), .A2(n14881), .ZN(P2_U3273) );
  INV_X1 U16505 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n14882) );
  NOR2_X1 U16506 ( .A1(n14888), .A2(n14882), .ZN(P2_U3274) );
  INV_X1 U16507 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n14883) );
  NOR2_X1 U16508 ( .A1(n14888), .A2(n14883), .ZN(P2_U3275) );
  INV_X1 U16509 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n14884) );
  NOR2_X1 U16510 ( .A1(n14888), .A2(n14884), .ZN(P2_U3276) );
  INV_X1 U16511 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n14885) );
  NOR2_X1 U16512 ( .A1(n14888), .A2(n14885), .ZN(P2_U3277) );
  INV_X1 U16513 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n14886) );
  NOR2_X1 U16514 ( .A1(n14888), .A2(n14886), .ZN(P2_U3278) );
  INV_X1 U16515 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n14887) );
  NOR2_X1 U16516 ( .A1(n14888), .A2(n14887), .ZN(P2_U3279) );
  INV_X1 U16517 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n14889) );
  NOR2_X1 U16518 ( .A1(n14910), .A2(n14889), .ZN(P2_U3280) );
  INV_X1 U16519 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n14890) );
  NOR2_X1 U16520 ( .A1(n14910), .A2(n14890), .ZN(P2_U3281) );
  INV_X1 U16521 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n14891) );
  NOR2_X1 U16522 ( .A1(n14910), .A2(n14891), .ZN(P2_U3282) );
  INV_X1 U16523 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n14892) );
  NOR2_X1 U16524 ( .A1(n14910), .A2(n14892), .ZN(P2_U3283) );
  INV_X1 U16525 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n14893) );
  NOR2_X1 U16526 ( .A1(n14910), .A2(n14893), .ZN(P2_U3284) );
  INV_X1 U16527 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n14894) );
  NOR2_X1 U16528 ( .A1(n14910), .A2(n14894), .ZN(P2_U3285) );
  INV_X1 U16529 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n14895) );
  NOR2_X1 U16530 ( .A1(n14910), .A2(n14895), .ZN(P2_U3286) );
  INV_X1 U16531 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n14896) );
  NOR2_X1 U16532 ( .A1(n14910), .A2(n14896), .ZN(P2_U3287) );
  INV_X1 U16533 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n14897) );
  NOR2_X1 U16534 ( .A1(n14910), .A2(n14897), .ZN(P2_U3288) );
  INV_X1 U16535 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n14898) );
  NOR2_X1 U16536 ( .A1(n14910), .A2(n14898), .ZN(P2_U3289) );
  INV_X1 U16537 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n14899) );
  NOR2_X1 U16538 ( .A1(n14910), .A2(n14899), .ZN(P2_U3290) );
  INV_X1 U16539 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n14900) );
  NOR2_X1 U16540 ( .A1(n14910), .A2(n14900), .ZN(P2_U3291) );
  INV_X1 U16541 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n14901) );
  NOR2_X1 U16542 ( .A1(n14910), .A2(n14901), .ZN(P2_U3292) );
  INV_X1 U16543 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n14902) );
  NOR2_X1 U16544 ( .A1(n14910), .A2(n14902), .ZN(P2_U3293) );
  INV_X1 U16545 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n14903) );
  NOR2_X1 U16546 ( .A1(n14910), .A2(n14903), .ZN(P2_U3294) );
  INV_X1 U16547 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n14904) );
  NOR2_X1 U16548 ( .A1(n14910), .A2(n14904), .ZN(P2_U3295) );
  INV_X1 U16549 ( .A(n14905), .ZN(n14909) );
  OAI22_X1 U16550 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n14910), .B1(n14909), .B2(
        n14906), .ZN(n14907) );
  INV_X1 U16551 ( .A(n14907), .ZN(P2_U3416) );
  OAI22_X1 U16552 ( .A1(P2_D_REG_1__SCAN_IN), .A2(n14910), .B1(n14909), .B2(
        n14908), .ZN(n14911) );
  INV_X1 U16553 ( .A(n14911), .ZN(P2_U3417) );
  INV_X1 U16554 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14912) );
  AOI22_X1 U16555 ( .A1(n6443), .A2(n14913), .B1(n14912), .B2(n14928), .ZN(
        P2_U3430) );
  INV_X1 U16556 ( .A(n14914), .ZN(n14918) );
  OAI21_X1 U16557 ( .B1(n7130), .B2(n14922), .A(n14915), .ZN(n14917) );
  AOI211_X1 U16558 ( .C1(n14927), .C2(n14918), .A(n14917), .B(n14916), .ZN(
        n14930) );
  INV_X1 U16559 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n14919) );
  AOI22_X1 U16560 ( .A1(n6443), .A2(n14930), .B1(n14919), .B2(n14928), .ZN(
        P2_U3454) );
  INV_X1 U16561 ( .A(n14920), .ZN(n14926) );
  OAI21_X1 U16562 ( .B1(n14923), .B2(n14922), .A(n14921), .ZN(n14925) );
  AOI211_X1 U16563 ( .C1(n14927), .C2(n14926), .A(n14925), .B(n14924), .ZN(
        n14932) );
  INV_X1 U16564 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n14929) );
  AOI22_X1 U16565 ( .A1(n6443), .A2(n14932), .B1(n14929), .B2(n14928), .ZN(
        P2_U3460) );
  AOI22_X1 U16566 ( .A1(n14933), .A2(n14930), .B1(n9657), .B2(n14931), .ZN(
        P2_U3507) );
  AOI22_X1 U16567 ( .A1(n14933), .A2(n14932), .B1(n10115), .B2(n14931), .ZN(
        P2_U3509) );
  NOR2_X1 U16568 ( .A1(P3_U3897), .A2(n15082), .ZN(P3_U3150) );
  AOI21_X1 U16569 ( .B1(n10597), .B2(n14935), .A(n14934), .ZN(n14948) );
  AOI21_X1 U16570 ( .B1(n14938), .B2(n14937), .A(n14936), .ZN(n14940) );
  OAI22_X1 U16571 ( .A1(n14940), .A2(n15109), .B1(n14939), .B2(n15101), .ZN(
        n14941) );
  AOI211_X1 U16572 ( .C1(P3_ADDR_REG_3__SCAN_IN), .C2(n15082), .A(n14942), .B(
        n14941), .ZN(n14947) );
  OAI21_X1 U16573 ( .B1(P3_REG1_REG_3__SCAN_IN), .B2(n14944), .A(n14943), .ZN(
        n14945) );
  NAND2_X1 U16574 ( .A1(n15107), .A2(n14945), .ZN(n14946) );
  OAI211_X1 U16575 ( .C1(n14948), .C2(n15116), .A(n14947), .B(n14946), .ZN(
        P3_U3185) );
  INV_X1 U16576 ( .A(n14949), .ZN(n14953) );
  INV_X1 U16577 ( .A(n14950), .ZN(n14951) );
  AOI21_X1 U16578 ( .B1(n14953), .B2(n14952), .A(n14951), .ZN(n14954) );
  INV_X1 U16579 ( .A(n14954), .ZN(n14959) );
  OAI21_X1 U16580 ( .B1(n14957), .B2(n14956), .A(n14955), .ZN(n14958) );
  AOI22_X1 U16581 ( .A1(n14960), .A2(n14959), .B1(n15107), .B2(n14958), .ZN(
        n14966) );
  AOI21_X1 U16582 ( .B1(n14963), .B2(n14962), .A(n14961), .ZN(n14964) );
  OR2_X1 U16583 ( .A1(n14964), .A2(n15109), .ZN(n14965) );
  OAI211_X1 U16584 ( .C1(n15101), .C2(n14967), .A(n14966), .B(n14965), .ZN(
        n14968) );
  INV_X1 U16585 ( .A(n14968), .ZN(n14970) );
  OAI211_X1 U16586 ( .C1(n7117), .C2(n15104), .A(n14970), .B(n14969), .ZN(
        P3_U3186) );
  AOI21_X1 U16587 ( .B1(n10633), .B2(n14972), .A(n14971), .ZN(n14986) );
  NOR2_X1 U16588 ( .A1(n14974), .A2(n14973), .ZN(n14975) );
  XNOR2_X1 U16589 ( .A(n14976), .B(n14975), .ZN(n14978) );
  OAI22_X1 U16590 ( .A1(n14978), .A2(n15109), .B1(n14977), .B2(n15101), .ZN(
        n14979) );
  AOI211_X1 U16591 ( .C1(n15082), .C2(P3_ADDR_REG_5__SCAN_IN), .A(n14980), .B(
        n14979), .ZN(n14985) );
  OAI21_X1 U16592 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n14982), .A(n14981), .ZN(
        n14983) );
  NAND2_X1 U16593 ( .A1(n15107), .A2(n14983), .ZN(n14984) );
  OAI211_X1 U16594 ( .C1(n14986), .C2(n15116), .A(n14985), .B(n14984), .ZN(
        P3_U3187) );
  OAI21_X1 U16595 ( .B1(n14989), .B2(n14988), .A(n14987), .ZN(n15004) );
  INV_X1 U16596 ( .A(n14990), .ZN(n14991) );
  AOI21_X1 U16597 ( .B1(n14993), .B2(n14992), .A(n14991), .ZN(n15002) );
  INV_X1 U16598 ( .A(n14994), .ZN(n14999) );
  OAI21_X1 U16599 ( .B1(n14997), .B2(n14996), .A(n14995), .ZN(n14998) );
  AOI22_X1 U16600 ( .A1(n15000), .A2(n14999), .B1(n15107), .B2(n14998), .ZN(
        n15001) );
  OAI21_X1 U16601 ( .B1(n15002), .B2(n15116), .A(n15001), .ZN(n15003) );
  AOI21_X1 U16602 ( .B1(n15004), .B2(n15090), .A(n15003), .ZN(n15006) );
  OAI211_X1 U16603 ( .C1(n15104), .C2(n15007), .A(n15006), .B(n15005), .ZN(
        P3_U3188) );
  AOI21_X1 U16604 ( .B1(n15010), .B2(n15009), .A(n15008), .ZN(n15023) );
  NAND2_X1 U16605 ( .A1(n6601), .A2(n15011), .ZN(n15012) );
  XNOR2_X1 U16606 ( .A(n15013), .B(n15012), .ZN(n15015) );
  OAI22_X1 U16607 ( .A1(n15015), .A2(n15109), .B1(n15014), .B2(n15101), .ZN(
        n15016) );
  AOI211_X1 U16608 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n15082), .A(n15017), .B(
        n15016), .ZN(n15022) );
  OAI21_X1 U16609 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n15019), .A(n15018), .ZN(
        n15020) );
  NAND2_X1 U16610 ( .A1(n15020), .A2(n15107), .ZN(n15021) );
  OAI211_X1 U16611 ( .C1(n15023), .C2(n15116), .A(n15022), .B(n15021), .ZN(
        P3_U3191) );
  INV_X1 U16612 ( .A(n15024), .ZN(n15025) );
  AOI21_X1 U16613 ( .B1(n15027), .B2(n15026), .A(n15025), .ZN(n15042) );
  OAI21_X1 U16614 ( .B1(n15030), .B2(n15029), .A(n15028), .ZN(n15040) );
  NAND2_X1 U16615 ( .A1(n15082), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n15031) );
  OAI211_X1 U16616 ( .C1(n15101), .C2(n15033), .A(n15032), .B(n15031), .ZN(
        n15039) );
  AOI21_X1 U16617 ( .B1(n15036), .B2(n15035), .A(n15034), .ZN(n15037) );
  NOR2_X1 U16618 ( .A1(n15037), .A2(n15109), .ZN(n15038) );
  AOI211_X1 U16619 ( .C1(n15107), .C2(n15040), .A(n15039), .B(n15038), .ZN(
        n15041) );
  OAI21_X1 U16620 ( .B1(n15042), .B2(n15116), .A(n15041), .ZN(P3_U3192) );
  AOI21_X1 U16621 ( .B1(n12602), .B2(n15044), .A(n15043), .ZN(n15058) );
  OAI21_X1 U16622 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n15046), .A(n15045), 
        .ZN(n15051) );
  AOI21_X1 U16623 ( .B1(n15082), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n15047), 
        .ZN(n15048) );
  OAI21_X1 U16624 ( .B1(n15101), .B2(n15049), .A(n15048), .ZN(n15050) );
  AOI21_X1 U16625 ( .B1(n15051), .B2(n15107), .A(n15050), .ZN(n15057) );
  OAI21_X1 U16626 ( .B1(n15054), .B2(n15053), .A(n15052), .ZN(n15055) );
  NAND2_X1 U16627 ( .A1(n15055), .A2(n15090), .ZN(n15056) );
  OAI211_X1 U16628 ( .C1(n15058), .C2(n15116), .A(n15057), .B(n15056), .ZN(
        P3_U3193) );
  INV_X1 U16629 ( .A(n15059), .ZN(n15060) );
  AOI21_X1 U16630 ( .B1(n15062), .B2(n15061), .A(n15060), .ZN(n15076) );
  OAI21_X1 U16631 ( .B1(n15065), .B2(n15064), .A(n15063), .ZN(n15070) );
  AOI21_X1 U16632 ( .B1(n15082), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n15066), 
        .ZN(n15067) );
  OAI21_X1 U16633 ( .B1(n15101), .B2(n15068), .A(n15067), .ZN(n15069) );
  AOI21_X1 U16634 ( .B1(n15070), .B2(n15107), .A(n15069), .ZN(n15075) );
  OAI211_X1 U16635 ( .C1(n15073), .C2(n15072), .A(n15071), .B(n15090), .ZN(
        n15074) );
  OAI211_X1 U16636 ( .C1(n15076), .C2(n15116), .A(n15075), .B(n15074), .ZN(
        P3_U3194) );
  AOI21_X1 U16637 ( .B1(n12626), .B2(n15078), .A(n15077), .ZN(n15094) );
  OAI21_X1 U16638 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n15080), .A(n15079), 
        .ZN(n15086) );
  AOI21_X1 U16639 ( .B1(n15082), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n15081), 
        .ZN(n15083) );
  OAI21_X1 U16640 ( .B1(n15101), .B2(n15084), .A(n15083), .ZN(n15085) );
  AOI21_X1 U16641 ( .B1(n15086), .B2(n15107), .A(n15085), .ZN(n15093) );
  OAI21_X1 U16642 ( .B1(n15089), .B2(n15088), .A(n15087), .ZN(n15091) );
  NAND2_X1 U16643 ( .A1(n15091), .A2(n15090), .ZN(n15092) );
  OAI211_X1 U16644 ( .C1(n15094), .C2(n15116), .A(n15093), .B(n15092), .ZN(
        P3_U3195) );
  AOI21_X1 U16645 ( .B1(n15097), .B2(n15096), .A(n15095), .ZN(n15117) );
  XOR2_X1 U16646 ( .A(n15099), .B(n15098), .Z(n15108) );
  NOR2_X1 U16647 ( .A1(n15101), .A2(n15100), .ZN(n15106) );
  INV_X1 U16648 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15103) );
  OAI21_X1 U16649 ( .B1(n15104), .B2(n15103), .A(n15102), .ZN(n15105) );
  AOI211_X1 U16650 ( .C1(n15108), .C2(n15107), .A(n15106), .B(n15105), .ZN(
        n15115) );
  AOI21_X1 U16651 ( .B1(n15111), .B2(n15110), .A(n15109), .ZN(n15113) );
  NAND2_X1 U16652 ( .A1(n15113), .A2(n15112), .ZN(n15114) );
  OAI211_X1 U16653 ( .C1(n15117), .C2(n15116), .A(n15115), .B(n15114), .ZN(
        P3_U3196) );
  XNOR2_X1 U16654 ( .A(n15118), .B(n15120), .ZN(n15127) );
  OAI21_X1 U16655 ( .B1(n15121), .B2(n15120), .A(n15119), .ZN(n15142) );
  OAI22_X1 U16656 ( .A1(n9097), .A2(n12799), .B1(n15123), .B2(n15122), .ZN(
        n15124) );
  AOI21_X1 U16657 ( .B1(n15142), .B2(n15125), .A(n15124), .ZN(n15126) );
  OAI21_X1 U16658 ( .B1(n15128), .B2(n15127), .A(n15126), .ZN(n15140) );
  NOR2_X1 U16659 ( .A1(n15129), .A2(n15144), .ZN(n15141) );
  AOI22_X1 U16660 ( .A1(n15142), .A2(n15131), .B1(n15141), .B2(n15130), .ZN(
        n15132) );
  INV_X1 U16661 ( .A(n15132), .ZN(n15133) );
  AOI211_X1 U16662 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n15134), .A(n15140), .B(
        n15133), .ZN(n15135) );
  AOI22_X1 U16663 ( .A1(n15136), .A2(n6874), .B1(n15135), .B2(n12818), .ZN(
        P3_U3231) );
  AOI211_X1 U16664 ( .C1(n15150), .C2(n15139), .A(n15138), .B(n15137), .ZN(
        n15160) );
  AOI22_X1 U16665 ( .A1(n15158), .A2(n15160), .B1(n8730), .B2(n15157), .ZN(
        P3_U3393) );
  AOI211_X1 U16666 ( .C1(n15143), .C2(n15142), .A(n15141), .B(n15140), .ZN(
        n15162) );
  AOI22_X1 U16667 ( .A1(n15158), .A2(n15162), .B1(n7047), .B2(n15157), .ZN(
        P3_U3396) );
  OAI22_X1 U16668 ( .A1(n15147), .A2(n15146), .B1(n15145), .B2(n15144), .ZN(
        n15148) );
  NOR2_X1 U16669 ( .A1(n15149), .A2(n15148), .ZN(n15163) );
  AOI22_X1 U16670 ( .A1(n15158), .A2(n15163), .B1(n8856), .B2(n15157), .ZN(
        P3_U3417) );
  AND2_X1 U16671 ( .A1(n15151), .A2(n15150), .ZN(n15155) );
  AND2_X1 U16672 ( .A1(n15153), .A2(n15152), .ZN(n15154) );
  NOR3_X1 U16673 ( .A1(n15156), .A2(n15155), .A3(n15154), .ZN(n15165) );
  AOI22_X1 U16674 ( .A1(n15158), .A2(n15165), .B1(n8839), .B2(n15157), .ZN(
        P3_U3420) );
  INV_X1 U16675 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15159) );
  AOI22_X1 U16676 ( .A1(n15166), .A2(n15160), .B1(n15159), .B2(n15164), .ZN(
        P3_U3460) );
  AOI22_X1 U16677 ( .A1(n15166), .A2(n15162), .B1(n15161), .B2(n15164), .ZN(
        P3_U3461) );
  AOI22_X1 U16678 ( .A1(n15166), .A2(n15163), .B1(n8852), .B2(n15164), .ZN(
        P3_U3468) );
  AOI22_X1 U16679 ( .A1(n15166), .A2(n15165), .B1(n12583), .B2(n15164), .ZN(
        P3_U3469) );
  OAI21_X1 U16680 ( .B1(n15169), .B2(n15168), .A(n15167), .ZN(SUB_1596_U59) );
  OAI21_X1 U16681 ( .B1(n15172), .B2(n15171), .A(n15170), .ZN(SUB_1596_U58) );
  XOR2_X1 U16682 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15173), .Z(SUB_1596_U53) );
  OAI21_X1 U16683 ( .B1(n15176), .B2(n15175), .A(n15174), .ZN(n15178) );
  XNOR2_X1 U16684 ( .A(n15178), .B(n15177), .ZN(SUB_1596_U56) );
  OAI21_X1 U16685 ( .B1(n15181), .B2(n15180), .A(n15179), .ZN(n15182) );
  XNOR2_X1 U16686 ( .A(n15182), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  AOI21_X1 U16687 ( .B1(n15185), .B2(n15184), .A(n15183), .ZN(SUB_1596_U5) );
  INV_X2 U7542 ( .A(n12026), .ZN(n11873) );
  INV_X2 U7183 ( .A(n12327), .ZN(n12317) );
  CLKBUF_X2 U7193 ( .A(n6449), .Z(n6436) );
  OR2_X1 U7237 ( .A1(n13264), .A2(n13438), .ZN(n13254) );
  NOR2_X2 U7238 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7545) );
  INV_X1 U7239 ( .A(n8748), .ZN(n9089) );
  CLKBUF_X1 U7240 ( .A(n7570), .Z(n6704) );
  AND4_X2 U7254 ( .A1(n8735), .A2(n8734), .A3(n8733), .A4(n8732), .ZN(n9097)
         );
  NAND4_X1 U7304 ( .A1(n8724), .A2(n8723), .A3(n8722), .A4(n8721), .ZN(n12559)
         );
  CLKBUF_X2 U7516 ( .A(n7563), .Z(n6449) );
endmodule

