

module b15_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, 
        DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, 
        DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, 
        DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, 
        DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, 
        DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, 
        HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3621, n3622, n3623, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767;

  AOI21_X1 U3654 ( .B1(n5248), .B2(n5247), .A(n5288), .ZN(n6707) );
  XNOR2_X1 U3655 ( .A(n5257), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n7059)
         );
  AOI211_X2 U3656 ( .C1(n7508), .C2(n7071), .A(n6581), .B(n7085), .ZN(n7062)
         );
  NAND2_X1 U3657 ( .A1(n6627), .A2(n3684), .ZN(n6607) );
  INV_X1 U3658 ( .A(n5512), .ZN(n5504) );
  BUF_X1 U3659 ( .A(n5432), .Z(n3662) );
  CLKBUF_X2 U3661 ( .A(n3903), .Z(n5769) );
  CLKBUF_X2 U3662 ( .A(n3639), .Z(n3661) );
  CLKBUF_X2 U3663 ( .A(n4004), .Z(n5260) );
  BUF_X2 U3664 ( .A(n3957), .Z(n6280) );
  CLKBUF_X2 U3665 ( .A(n3847), .Z(n5591) );
  AND4_X1 U3666 ( .A1(n3907), .A2(n3906), .A3(n3905), .A4(n3904), .ZN(n3908)
         );
  AND4_X1 U3667 ( .A1(n3811), .A2(n3810), .A3(n3809), .A4(n3808), .ZN(n3854)
         );
  BUF_X2 U3669 ( .A(n4003), .Z(n3639) );
  AND2_X2 U3670 ( .A1(n3760), .A2(n5770), .ZN(n4552) );
  AND2_X2 U3671 ( .A1(n3760), .A2(n5770), .ZN(n3650) );
  BUF_X2 U3673 ( .A(n4397), .Z(n3651) );
  AND2_X1 U3675 ( .A1(n3766), .A2(n3765), .ZN(n4020) );
  INV_X1 U3677 ( .A(n7766), .ZN(n3621) );
  CLKBUF_X3 U3678 ( .A(n4032), .Z(n3660) );
  AND2_X2 U3679 ( .A1(n5770), .A2(n5762), .ZN(n4397) );
  NOR2_X2 U3680 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5799) );
  AND2_X2 U3681 ( .A1(n3765), .A2(n5762), .ZN(n3648) );
  NAND2_X1 U3682 ( .A1(n6680), .A2(n6586), .ZN(n5135) );
  AND4_X1 U3683 ( .A1(n3895), .A2(n3894), .A3(n3893), .A4(n3892), .ZN(n3896)
         );
  NAND2_X1 U3685 ( .A1(n3862), .A2(n3860), .ZN(n3836) );
  MUX2_X1 U3686 ( .A(n6571), .B(n5256), .S(n3631), .Z(n5257) );
  NAND2_X1 U3687 ( .A1(n6974), .A2(n6976), .ZN(n6975) );
  OAI21_X1 U3688 ( .B1(n5512), .B2(n7726), .A(n5925), .ZN(n5511) );
  INV_X2 U3689 ( .A(n3847), .ZN(n3956) );
  OR2_X2 U3690 ( .A1(n6736), .A2(n5287), .ZN(n6663) );
  INV_X1 U3692 ( .A(n7696), .ZN(n7679) );
  INV_X2 U3693 ( .A(n7682), .ZN(n7699) );
  AOI21_X1 U3694 ( .B1(n6685), .B2(n7421), .A(n6667), .ZN(n6668) );
  AND2_X1 U3695 ( .A1(n6833), .A2(n3732), .ZN(n6786) );
  AND2_X2 U3696 ( .A1(n3766), .A2(n5770), .ZN(n4009) );
  BUF_X2 U3697 ( .A(n4009), .Z(n3654) );
  NAND2_X2 U3699 ( .A1(n4241), .A2(n4240), .ZN(n6220) );
  NAND2_X2 U3700 ( .A1(n4256), .A2(n4255), .ZN(n6469) );
  OAI21_X2 U3701 ( .B1(n6501), .B2(n6503), .A(n4254), .ZN(n4256) );
  AOI21_X1 U3702 ( .B1(n3994), .B2(n6064), .A(n5591), .ZN(n3991) );
  OAI222_X1 U3703 ( .A1(n6260), .A2(n5438), .B1(n6256), .B2(n6219), .C1(n7193), 
        .C2(n6218), .ZN(U3464) );
  AOI21_X2 U3704 ( .B1(n6975), .B2(n5255), .A(n5254), .ZN(n6571) );
  NOR2_X2 U3705 ( .A1(n5422), .A2(n4001), .ZN(n4018) );
  INV_X1 U3706 ( .A(n3891), .ZN(n4011) );
  BUF_X2 U3707 ( .A(n3915), .Z(n3622) );
  BUF_X2 U3708 ( .A(n3915), .Z(n3623) );
  AND2_X1 U3709 ( .A1(n3765), .A2(n3760), .ZN(n3915) );
  CLKBUF_X1 U3710 ( .A(n4260), .Z(n3632) );
  XNOR2_X1 U3711 ( .A(n4245), .B(n4232), .ZN(n4331) );
  XNOR2_X1 U3712 ( .A(n4220), .B(n4204), .ZN(n4310) );
  NAND2_X1 U3714 ( .A1(n4182), .A2(n4181), .ZN(n4220) );
  INV_X1 U3715 ( .A(n7508), .ZN(n6580) );
  BUF_X1 U3716 ( .A(n5502), .Z(n3640) );
  NAND2_X1 U3717 ( .A1(n4078), .A2(n4077), .ZN(n5393) );
  AND2_X1 U3718 ( .A1(n4157), .A2(n4156), .ZN(n4159) );
  CLKBUF_X3 U3719 ( .A(n5433), .Z(n3646) );
  NAND2_X1 U3720 ( .A1(n4148), .A2(n4147), .ZN(n4157) );
  NAND2_X1 U3721 ( .A1(n7369), .A2(n6670), .ZN(n6917) );
  XNOR2_X1 U3722 ( .A(n5801), .B(n5865), .ZN(n5436) );
  NAND4_X2 U3723 ( .A1(n3795), .A2(n3794), .A3(n3793), .A4(n3792), .ZN(n3860)
         );
  CLKBUF_X3 U3724 ( .A(n3922), .Z(n3657) );
  AND2_X2 U3725 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5762) );
  INV_X2 U3726 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3725) );
  INV_X2 U3727 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4279) );
  AOI21_X1 U3728 ( .B1(n3689), .B2(n7696), .A(n3688), .ZN(n3687) );
  INV_X1 U3729 ( .A(n4705), .ZN(n6710) );
  INV_X1 U3730 ( .A(n7007), .ZN(n3625) );
  XNOR2_X1 U3731 ( .A(n6612), .B(n6611), .ZN(n7069) );
  NAND2_X1 U3732 ( .A1(n6595), .A2(n6594), .ZN(n6881) );
  NAND2_X1 U3733 ( .A1(n6591), .A2(n6590), .ZN(n6595) );
  NAND2_X1 U3734 ( .A1(n6609), .A2(n6608), .ZN(n6612) );
  AND2_X1 U3735 ( .A1(n4433), .A2(n4428), .ZN(n6491) );
  OAI21_X1 U3736 ( .B1(n6289), .B2(n6449), .A(n4427), .ZN(n4428) );
  AOI211_X1 U3737 ( .C1(n6867), .C2(n7569), .A(n6866), .B(n6865), .ZN(n6868)
         );
  NOR2_X1 U3738 ( .A1(n6720), .A2(n6721), .ZN(n5319) );
  AOI21_X1 U3739 ( .B1(n3698), .B2(n3700), .A(n3669), .ZN(n3695) );
  AND2_X1 U3740 ( .A1(n4258), .A2(n3708), .ZN(n3664) );
  AOI21_X1 U3741 ( .B1(n7395), .B2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n3713), 
        .ZN(n3712) );
  OAI21_X1 U3742 ( .B1(n6221), .B2(n3700), .A(n6269), .ZN(n3699) );
  OR2_X1 U3743 ( .A1(n6470), .A2(n3709), .ZN(n3708) );
  NAND2_X1 U3744 ( .A1(n3670), .A2(n4257), .ZN(n3709) );
  XNOR2_X1 U3745 ( .A(n4250), .B(n6222), .ZN(n6221) );
  NAND2_X1 U3746 ( .A1(n4252), .A2(n7091), .ZN(n4267) );
  NAND2_X1 U3747 ( .A1(n4301), .A2(n4300), .ZN(n5362) );
  NOR2_X1 U3748 ( .A1(n4701), .A2(n4712), .ZN(n5242) );
  NAND2_X1 U3749 ( .A1(n4276), .A2(n4275), .ZN(n5355) );
  NAND2_X1 U3750 ( .A1(n4158), .A2(n4156), .ZN(n4149) );
  NOR2_X1 U3751 ( .A1(n5564), .A2(n3638), .ZN(n6430) );
  NAND2_X1 U3752 ( .A1(n5436), .A2(n7437), .ZN(n4148) );
  NOR2_X1 U3753 ( .A1(n5564), .A2(n5452), .ZN(n6409) );
  NOR2_X1 U3754 ( .A1(n5564), .A2(n6067), .ZN(n6388) );
  NAND2_X1 U3755 ( .A1(n4092), .A2(n3702), .ZN(n5433) );
  NOR2_X1 U3756 ( .A1(n5564), .A2(n6670), .ZN(n6395) );
  NAND2_X1 U3757 ( .A1(n5406), .A2(n5405), .ZN(n5428) );
  CLKBUF_X1 U3758 ( .A(n5437), .Z(n3663) );
  MUX2_X1 U3759 ( .A(n5346), .B(n5282), .S(n5345), .Z(n5354) );
  NAND2_X1 U3760 ( .A1(n5397), .A2(n5396), .ZN(n5794) );
  AND2_X1 U3761 ( .A1(n3635), .A2(n3636), .ZN(n4049) );
  NAND2_X1 U3762 ( .A1(n3886), .A2(n3885), .ZN(n5790) );
  NOR2_X1 U3763 ( .A1(n5498), .A2(n5499), .ZN(n5491) );
  NOR2_X1 U3764 ( .A1(n4499), .A2(n7026), .ZN(n4500) );
  NOR2_X1 U3765 ( .A1(n4465), .A2(n6824), .ZN(n4481) );
  INV_X1 U3766 ( .A(n5118), .ZN(n3945) );
  NAND2_X1 U3767 ( .A1(n4044), .A2(n4242), .ZN(n4081) );
  AND3_X1 U3768 ( .A1(n5423), .A2(n3993), .A3(n3992), .ZN(n3999) );
  NAND2_X4 U3769 ( .A1(n5322), .A2(n6586), .ZN(n6587) );
  AND2_X1 U3770 ( .A1(n3746), .A2(n6680), .ZN(n5320) );
  NOR2_X1 U3771 ( .A1(n3836), .A2(n4082), .ZN(n3884) );
  CLKBUF_X2 U3772 ( .A(n3961), .Z(n3638) );
  INV_X2 U3773 ( .A(n4548), .ZN(n6660) );
  INV_X1 U3774 ( .A(n4052), .ZN(n3626) );
  NAND2_X2 U3775 ( .A1(n4064), .A2(n4063), .ZN(n4229) );
  NAND2_X2 U3776 ( .A1(n5449), .A2(n6280), .ZN(n5322) );
  CLKBUF_X1 U3777 ( .A(n3935), .Z(n5563) );
  CLKBUF_X1 U3778 ( .A(n4272), .Z(n4457) );
  OR2_X1 U3779 ( .A1(n4042), .A2(n4041), .ZN(n4083) );
  OR2_X1 U3780 ( .A1(n4031), .A2(n4030), .ZN(n4247) );
  AND2_X1 U3781 ( .A1(n4346), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4362)
         );
  CLKBUF_X2 U3782 ( .A(n4045), .Z(n5452) );
  OR2_X1 U3783 ( .A1(n3860), .A2(n7437), .ZN(n4063) );
  NOR2_X1 U3784 ( .A1(n4325), .A2(n7404), .ZN(n4346) );
  NAND4_X2 U3785 ( .A1(n3832), .A2(n3831), .A3(n3830), .A4(n3829), .ZN(n3847)
         );
  AND4_X1 U3786 ( .A1(n3914), .A2(n3913), .A3(n3912), .A4(n3911), .ZN(n3667)
         );
  NAND2_X2 U3787 ( .A1(n3897), .A2(n3896), .ZN(n3937) );
  NAND2_X2 U3788 ( .A1(n3931), .A2(n3740), .ZN(n3994) );
  AND4_X1 U3789 ( .A1(n3813), .A2(n3814), .A3(n3815), .A4(n3812), .ZN(n3832)
         );
  AND4_X1 U3790 ( .A1(n3759), .A2(n3758), .A3(n3757), .A4(n3756), .ZN(n3774)
         );
  AND4_X1 U3791 ( .A1(n3764), .A2(n3763), .A3(n3762), .A4(n3761), .ZN(n3773)
         );
  AND4_X1 U3792 ( .A1(n3787), .A2(n3786), .A3(n3785), .A4(n3784), .ZN(n3793)
         );
  AND4_X1 U3793 ( .A1(n3779), .A2(n3778), .A3(n3777), .A4(n3776), .ZN(n3795)
         );
  AND4_X1 U3794 ( .A1(n3755), .A2(n3754), .A3(n3753), .A4(n3752), .ZN(n3775)
         );
  AND4_X1 U3795 ( .A1(n3771), .A2(n3770), .A3(n3769), .A4(n3768), .ZN(n3772)
         );
  AND4_X1 U3796 ( .A1(n3819), .A2(n3818), .A3(n3817), .A4(n3816), .ZN(n3831)
         );
  AND4_X1 U3797 ( .A1(n3783), .A2(n3782), .A3(n3781), .A4(n3780), .ZN(n3794)
         );
  AND4_X1 U3798 ( .A1(n3926), .A2(n3925), .A3(n3924), .A4(n3923), .ZN(n3931)
         );
  AND4_X1 U3799 ( .A1(n3791), .A2(n3790), .A3(n3789), .A4(n3788), .ZN(n3792)
         );
  AND4_X1 U3800 ( .A1(n3919), .A2(n3918), .A3(n3917), .A4(n3916), .ZN(n3920)
         );
  AND4_X1 U3801 ( .A1(n3828), .A2(n3827), .A3(n3826), .A4(n3825), .ZN(n3829)
         );
  AND4_X1 U3802 ( .A1(n3807), .A2(n3806), .A3(n3805), .A4(n3804), .ZN(n3855)
         );
  AND4_X1 U3803 ( .A1(n3803), .A2(n3802), .A3(n3801), .A4(n3800), .ZN(n3856)
         );
  AND4_X1 U3804 ( .A1(n3799), .A2(n3798), .A3(n3797), .A4(n3796), .ZN(n3857)
         );
  AND2_X1 U3805 ( .A1(n3821), .A2(n3820), .ZN(n3823) );
  NAND2_X2 U3807 ( .A1(STATE_REG_2__SCAN_IN), .A2(n7734), .ZN(n7338) );
  NAND2_X2 U3808 ( .A1(n7734), .A2(n7737), .ZN(n7320) );
  BUF_X4 U3809 ( .A(n3921), .Z(n4689) );
  CLKBUF_X3 U3810 ( .A(n3921), .Z(n4351) );
  BUF_X2 U3811 ( .A(n4025), .Z(n5261) );
  BUF_X2 U3812 ( .A(n4020), .Z(n5259) );
  CLKBUF_X2 U3813 ( .A(n3922), .Z(n3655) );
  BUF_X4 U3814 ( .A(n4009), .Z(n3627) );
  AND2_X2 U3816 ( .A1(n3760), .A2(n5796), .ZN(n3643) );
  NAND2_X1 U3818 ( .A1(n3957), .A2(n3956), .ZN(n4073) );
  NAND2_X1 U3819 ( .A1(n3935), .A2(n3956), .ZN(n3946) );
  INV_X2 U3820 ( .A(n4073), .ZN(n3958) );
  AND2_X1 U3821 ( .A1(n3949), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3629) );
  INV_X1 U3822 ( .A(n5785), .ZN(n3630) );
  NAND2_X1 U3823 ( .A1(n3945), .A2(n3956), .ZN(n5803) );
  INV_X2 U3824 ( .A(n3937), .ZN(n5446) );
  NAND2_X1 U3825 ( .A1(n6528), .A2(n6527), .ZN(n7007) );
  INV_X2 U3826 ( .A(n4252), .ZN(n3631) );
  AND2_X2 U3827 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5796) );
  BUF_X4 U3828 ( .A(n3922), .Z(n3656) );
  NAND2_X1 U3829 ( .A1(n3706), .A2(n3703), .ZN(n7036) );
  NOR2_X2 U3830 ( .A1(n5307), .A2(n6772), .ZN(n3694) );
  NOR2_X2 U3831 ( .A1(n5490), .A2(n3691), .ZN(n5526) );
  NOR2_X2 U3832 ( .A1(n6758), .A2(n6539), .ZN(n6735) );
  NAND2_X2 U3833 ( .A1(n6833), .A2(n3633), .ZN(n6787) );
  AND2_X1 U3834 ( .A1(n3732), .A2(n6789), .ZN(n3633) );
  NAND2_X1 U3836 ( .A1(n4055), .A2(n3637), .ZN(n3635) );
  OR2_X1 U3837 ( .A1(n3626), .A2(n4079), .ZN(n3636) );
  AND2_X1 U3838 ( .A1(n4081), .A2(n4052), .ZN(n3637) );
  INV_X2 U3839 ( .A(n3983), .ZN(n3961) );
  AOI21_X2 U3840 ( .B1(n6255), .B2(n4277), .A(n5838), .ZN(n5346) );
  OAI21_X2 U3842 ( .B1(n6992), .B2(n6537), .A(n6536), .ZN(n6538) );
  XNOR2_X1 U3843 ( .A(n4180), .B(n4181), .ZN(n4309) );
  NAND2_X1 U3844 ( .A1(n5360), .A2(n5362), .ZN(n5361) );
  XNOR2_X1 U3845 ( .A(n4149), .B(n4157), .ZN(n5502) );
  NOR2_X2 U3846 ( .A1(n7000), .A2(n6999), .ZN(n6998) );
  NAND2_X1 U3847 ( .A1(n4245), .A2(n4244), .ZN(n3641) );
  NAND2_X1 U3848 ( .A1(n4245), .A2(n4244), .ZN(n3642) );
  INV_X1 U3849 ( .A(n4126), .ZN(n4158) );
  NAND2_X1 U3850 ( .A1(n4289), .A2(n4626), .ZN(n5530) );
  INV_X2 U3851 ( .A(n4292), .ZN(n5360) );
  AND2_X4 U3852 ( .A1(n3725), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3760)
         );
  NOR2_X4 U3853 ( .A1(n6723), .A2(n6712), .ZN(n6627) );
  NAND2_X2 U3854 ( .A1(n3973), .A2(n3972), .ZN(n4098) );
  INV_X2 U3855 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3720) );
  AND2_X2 U3856 ( .A1(n3760), .A2(n5796), .ZN(n3644) );
  AND2_X2 U3858 ( .A1(n3751), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3765)
         );
  INV_X2 U3859 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3751) );
  AND2_X4 U3861 ( .A1(n3720), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5770)
         );
  NOR2_X2 U3862 ( .A1(n5361), .A2(n5496), .ZN(n5487) );
  NOR2_X2 U3863 ( .A1(n6228), .A2(n4378), .ZN(n6261) );
  NAND3_X2 U3864 ( .A1(n3726), .A2(n3673), .A3(n4332), .ZN(n6228) );
  AND2_X2 U3865 ( .A1(n6563), .A2(n6737), .ZN(n6725) );
  NOR2_X2 U3866 ( .A1(n6561), .A2(n6564), .ZN(n6563) );
  NAND2_X2 U3867 ( .A1(n4019), .A2(n4002), .ZN(n4094) );
  AND2_X4 U3868 ( .A1(n3760), .A2(n3767), .ZN(n3921) );
  INV_X2 U3869 ( .A(n4011), .ZN(n4488) );
  NOR2_X2 U3870 ( .A1(n3997), .A2(n3932), .ZN(n3953) );
  AND2_X1 U3871 ( .A1(n3765), .A2(n5762), .ZN(n3647) );
  AND2_X2 U3872 ( .A1(n3765), .A2(n5762), .ZN(n5258) );
  AND2_X1 U3873 ( .A1(n3760), .A2(n5770), .ZN(n3649) );
  BUF_X4 U3874 ( .A(n4009), .Z(n3653) );
  BUF_X4 U3875 ( .A(n4032), .Z(n3659) );
  XNOR2_X1 U3876 ( .A(n4126), .B(n4156), .ZN(n5432) );
  OR2_X2 U3877 ( .A1(n5438), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4061) );
  XNOR2_X2 U3878 ( .A(n4093), .B(n4094), .ZN(n5438) );
  INV_X1 U3879 ( .A(n6004), .ZN(n3729) );
  NOR2_X1 U3880 ( .A1(n4252), .A2(n5220), .ZN(n5254) );
  OR2_X1 U3881 ( .A1(n4219), .A2(n4221), .ZN(n4218) );
  INV_X1 U3882 ( .A(n4082), .ZN(n4243) );
  NAND2_X1 U3883 ( .A1(n4074), .A2(n5591), .ZN(n4082) );
  INV_X1 U3884 ( .A(n4626), .ZN(n6659) );
  NAND2_X1 U3885 ( .A1(n5790), .A2(n7711), .ZN(n5404) );
  NOR2_X1 U3886 ( .A1(n3686), .A2(n3685), .ZN(n3684) );
  INV_X1 U3887 ( .A(n5334), .ZN(n3685) );
  NOR2_X1 U3888 ( .A1(n3674), .A2(n7033), .ZN(n3710) );
  NAND2_X1 U3890 ( .A1(n4769), .A2(n4768), .ZN(n4772) );
  INV_X1 U3891 ( .A(n4880), .ZN(n4889) );
  AND2_X1 U3892 ( .A1(n4229), .A2(n3846), .ZN(n3871) );
  AND2_X1 U3893 ( .A1(n3946), .A2(n3848), .ZN(n3872) );
  NAND2_X1 U3894 ( .A1(n3939), .A2(n4045), .ZN(n3965) );
  AND2_X1 U3895 ( .A1(n4217), .A2(n4216), .ZN(n4221) );
  INV_X1 U3896 ( .A(n4180), .ZN(n4182) );
  AOI21_X1 U3897 ( .B1(n7181), .B2(n7198), .A(n3750), .ZN(n3833) );
  NOR2_X1 U3898 ( .A1(n3837), .A2(n3749), .ZN(n3750) );
  NOR2_X1 U3899 ( .A1(n5135), .A2(EBX_REG_1__SCAN_IN), .ZN(n5128) );
  NAND2_X1 U3900 ( .A1(n6902), .A2(n6903), .ZN(n3731) );
  NAND2_X1 U3901 ( .A1(n4466), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5278) );
  NOR2_X1 U3902 ( .A1(n3680), .A2(n6828), .ZN(n3679) );
  INV_X1 U3903 ( .A(n6814), .ZN(n3680) );
  AND2_X1 U3904 ( .A1(n3709), .A2(n3677), .ZN(n3705) );
  INV_X1 U3905 ( .A(n4251), .ZN(n3700) );
  INV_X1 U3906 ( .A(n5652), .ZN(n5148) );
  INV_X1 U3907 ( .A(n4063), .ZN(n4242) );
  OR2_X1 U3908 ( .A1(n6280), .A2(n7437), .ZN(n4064) );
  AND2_X1 U3909 ( .A1(n6280), .A2(n3722), .ZN(n3721) );
  AND2_X1 U3910 ( .A1(n3952), .A2(n3951), .ZN(n3976) );
  AOI21_X1 U3911 ( .B1(n3859), .B2(n4243), .A(n5115), .ZN(n3880) );
  INV_X1 U3912 ( .A(n3957), .ZN(n3935) );
  INV_X1 U3913 ( .A(n3860), .ZN(n4045) );
  OAI21_X1 U3914 ( .B1(n7446), .B2(n6253), .A(n7177), .ZN(n5445) );
  CLKBUF_X1 U3915 ( .A(n5366), .Z(n5367) );
  CLKBUF_X1 U3916 ( .A(n4073), .Z(n7443) );
  NAND2_X1 U3917 ( .A1(n7431), .A2(n5121), .ZN(n6871) );
  AND3_X1 U3918 ( .A1(n7220), .A2(n7524), .A3(n7719), .ZN(n5121) );
  NAND2_X1 U3919 ( .A1(n6871), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6281) );
  NAND2_X1 U3920 ( .A1(n6725), .A2(n3735), .ZN(n4705) );
  NOR2_X1 U3921 ( .A1(n6711), .A2(n3736), .ZN(n3735) );
  INV_X1 U3922 ( .A(n6724), .ZN(n3736) );
  AND3_X1 U3923 ( .A1(n4345), .A2(n4344), .A3(n4343), .ZN(n6004) );
  AOI21_X1 U3924 ( .B1(n4331), .B2(n4457), .A(n4330), .ZN(n5524) );
  INV_X1 U3925 ( .A(n4318), .ZN(n4319) );
  NAND2_X1 U3926 ( .A1(n4319), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4325)
         );
  AOI21_X1 U3927 ( .B1(n3662), .B2(n4243), .A(n4123), .ZN(n7376) );
  NOR2_X1 U3928 ( .A1(n3631), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3715)
         );
  NAND2_X1 U3929 ( .A1(n3675), .A2(n4267), .ZN(n3719) );
  INV_X1 U3930 ( .A(n5254), .ZN(n3717) );
  NAND2_X1 U3931 ( .A1(n6966), .A2(n3717), .ZN(n3716) );
  NOR2_X1 U3932 ( .A1(n6966), .A2(n3719), .ZN(n6570) );
  INV_X1 U3933 ( .A(n6966), .ZN(n3718) );
  INV_X1 U3934 ( .A(n7018), .ZN(n6527) );
  XNOR2_X1 U3935 ( .A(n4252), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6470)
         );
  XNOR2_X1 U3936 ( .A(n3642), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6269)
         );
  OAI21_X1 U3937 ( .B1(n5794), .B2(n5399), .A(n7711), .ZN(n5406) );
  INV_X1 U3938 ( .A(n3671), .ZN(n4070) );
  NAND2_X1 U3939 ( .A1(n4092), .A2(n4091), .ZN(n4126) );
  NAND2_X1 U3940 ( .A1(n7437), .A2(n5445), .ZN(n5808) );
  AND2_X1 U3941 ( .A1(n7705), .A2(n5806), .ZN(n7208) );
  INV_X1 U3942 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n7437) );
  AND2_X1 U3943 ( .A1(n4908), .A2(n4907), .ZN(n4914) );
  AND2_X1 U3944 ( .A1(n6871), .A2(STATE2_REG_3__SCAN_IN), .ZN(n7688) );
  INV_X1 U3945 ( .A(n7693), .ZN(n7666) );
  NAND2_X2 U3946 ( .A1(n5304), .A2(n5303), .ZN(n7369) );
  OR3_X1 U3947 ( .A1(n5790), .A2(n7211), .A3(n6678), .ZN(n5304) );
  NAND2_X1 U3948 ( .A1(n6063), .A2(n6062), .ZN(n6952) );
  AOI21_X1 U3949 ( .B1(n6061), .B2(n7711), .A(n6060), .ZN(n6062) );
  INV_X1 U3950 ( .A(n7405), .ZN(n7415) );
  NAND2_X1 U3951 ( .A1(n6607), .A2(n3746), .ZN(n6608) );
  INV_X1 U3952 ( .A(n7251), .ZN(n6218) );
  NAND2_X1 U3953 ( .A1(n4772), .A2(n4771), .ZN(n4782) );
  NOR2_X1 U3954 ( .A1(n4799), .A2(n4798), .ZN(n4803) );
  NAND2_X1 U3955 ( .A1(n4823), .A2(n4822), .ZN(n4834) );
  NAND2_X1 U3956 ( .A1(n4846), .A2(n4845), .ZN(n4856) );
  NAND2_X1 U3957 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n5726), .ZN(n3861) );
  AND2_X1 U3958 ( .A1(n3840), .A2(n3841), .ZN(n3839) );
  AOI21_X1 U3959 ( .B1(n4889), .B2(n4888), .A(n4887), .ZN(n4890) );
  NAND2_X1 U3960 ( .A1(n4159), .A2(n4158), .ZN(n4180) );
  CLKBUF_X2 U3961 ( .A(n4104), .Z(n5266) );
  OR2_X1 U3962 ( .A1(n4193), .A2(n4192), .ZN(n4224) );
  OR2_X1 U3963 ( .A1(n4170), .A2(n4169), .ZN(n4196) );
  AND2_X1 U3964 ( .A1(n3957), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3862) );
  OR2_X1 U3965 ( .A1(n4017), .A2(n4016), .ZN(n4071) );
  INV_X1 U3966 ( .A(n4229), .ZN(n3859) );
  INV_X1 U3967 ( .A(n5112), .ZN(n3877) );
  OR2_X1 U3968 ( .A1(n3645), .A2(n6648), .ZN(n5727) );
  AOI22_X1 U3969 ( .A1(n3649), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3639), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3888) );
  NOR2_X1 U3970 ( .A1(n3938), .A2(n5449), .ZN(n3940) );
  AND2_X1 U3971 ( .A1(n3833), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3834)
         );
  NOR2_X1 U3972 ( .A1(n3994), .A2(n3957), .ZN(n3944) );
  AND2_X1 U3973 ( .A1(n6066), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4302) );
  OR2_X1 U3974 ( .A1(n6711), .A2(n5246), .ZN(n5285) );
  NOR2_X1 U3975 ( .A1(n6801), .A2(n3733), .ZN(n3732) );
  INV_X1 U3976 ( .A(n3734), .ZN(n3733) );
  AND2_X1 U3977 ( .A1(n4464), .A2(n6832), .ZN(n3734) );
  INV_X1 U3978 ( .A(n6822), .ZN(n4464) );
  NOR2_X1 U3979 ( .A1(n6794), .A2(n6905), .ZN(n6896) );
  NAND2_X1 U3980 ( .A1(n4278), .A2(n7437), .ZN(n4055) );
  AND2_X1 U3981 ( .A1(n3977), .A2(n3976), .ZN(n3975) );
  OR2_X1 U3982 ( .A1(n4114), .A2(n4113), .ZN(n4117) );
  OR2_X1 U3983 ( .A1(n4145), .A2(n4144), .ZN(n4151) );
  OR2_X1 U3984 ( .A1(n3663), .A2(n7169), .ZN(n5949) );
  OR2_X1 U3985 ( .A1(n3662), .A2(n5687), .ZN(n5917) );
  CLKBUF_X1 U3986 ( .A(n5118), .Z(n5119) );
  NAND2_X1 U3987 ( .A1(n3941), .A2(n6280), .ZN(n5111) );
  AND2_X1 U3988 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n4533), .ZN(n4534)
         );
  INV_X1 U3989 ( .A(n4532), .ZN(n4533) );
  INV_X1 U3990 ( .A(n7599), .ZN(n7618) );
  INV_X1 U3991 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6858) );
  INV_X1 U3992 ( .A(n7435), .ZN(n6682) );
  NOR2_X1 U3993 ( .A1(n5128), .A2(n5127), .ZN(n5129) );
  NOR2_X1 U3994 ( .A1(n6586), .A2(n6285), .ZN(n5127) );
  NOR2_X1 U3995 ( .A1(n6451), .A2(n6450), .ZN(n6483) );
  NOR3_X1 U3996 ( .A1(n3994), .A2(n3983), .A3(n4074), .ZN(n3947) );
  AND2_X1 U3997 ( .A1(n5369), .A2(n6682), .ZN(n7255) );
  NAND2_X1 U3998 ( .A1(n5592), .A2(n5368), .ZN(n5369) );
  OR2_X1 U3999 ( .A1(n5404), .A2(n7188), .ZN(n5368) );
  NOR2_X1 U4000 ( .A1(n5590), .A2(READY_N), .ZN(n5593) );
  OR2_X1 U4001 ( .A1(n5404), .A2(n7212), .ZN(n5592) );
  OR2_X1 U4002 ( .A1(n4649), .A2(n6727), .ZN(n4700) );
  AND2_X1 U4003 ( .A1(n6973), .A2(n5282), .ZN(n4645) );
  OR2_X1 U4004 ( .A1(n4623), .A2(n6985), .ZN(n4644) );
  NOR2_X1 U4005 ( .A1(n4570), .A2(n7001), .ZN(n4571) );
  NAND2_X1 U4006 ( .A1(n4571), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4623)
         );
  AND2_X1 U4007 ( .A1(n7683), .A2(n5282), .ZN(n4529) );
  NAND2_X1 U4008 ( .A1(n4500), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4532)
         );
  NAND2_X1 U4009 ( .A1(n4481), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4499)
         );
  NAND2_X1 U4010 ( .A1(n4448), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4465)
         );
  INV_X1 U4011 ( .A(n4434), .ZN(n4448) );
  NOR2_X1 U4012 ( .A1(n4429), .A2(n6848), .ZN(n4430) );
  NAND2_X1 U4013 ( .A1(n4430), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4434)
         );
  OR2_X1 U4014 ( .A1(n4393), .A2(n7632), .ZN(n4429) );
  CLKBUF_X1 U4015 ( .A(n6289), .Z(n6290) );
  OR2_X1 U4016 ( .A1(n4379), .A2(n7623), .ZN(n4393) );
  INV_X1 U4017 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n7632) );
  NAND2_X1 U4018 ( .A1(n4362), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4379)
         );
  INV_X1 U4019 ( .A(n6262), .ZN(n4378) );
  NAND2_X1 U4020 ( .A1(n4332), .A2(n3729), .ZN(n3727) );
  AOI21_X1 U4021 ( .B1(n4322), .B2(n4457), .A(n4321), .ZN(n5655) );
  INV_X1 U4022 ( .A(n4311), .ZN(n4312) );
  NAND2_X1 U4023 ( .A1(n4312), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4318)
         );
  CLKBUF_X1 U4024 ( .A(n5485), .Z(n5486) );
  NAND2_X1 U4025 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4293) );
  NAND2_X1 U4026 ( .A1(n5333), .A2(n6606), .ZN(n6609) );
  AND2_X1 U4027 ( .A1(n6627), .A2(n6629), .ZN(n5333) );
  NAND2_X1 U4028 ( .A1(n3694), .A2(n3693), .ZN(n6758) );
  INV_X1 U4029 ( .A(n6756), .ZN(n3693) );
  INV_X1 U4030 ( .A(n3694), .ZN(n6773) );
  AND2_X1 U4031 ( .A1(n5191), .A2(n5190), .ZN(n6897) );
  NAND2_X1 U4032 ( .A1(n6980), .A2(n4262), .ZN(n7019) );
  AND2_X1 U4033 ( .A1(n5181), .A2(n5180), .ZN(n6814) );
  AOI21_X1 U4034 ( .B1(n3664), .B2(n3705), .A(n3704), .ZN(n3703) );
  INV_X1 U4035 ( .A(n7041), .ZN(n3704) );
  AND3_X1 U4036 ( .A1(n4243), .A2(n4242), .A3(n4247), .ZN(n4244) );
  INV_X1 U4037 ( .A(n6231), .ZN(n3683) );
  NAND2_X1 U4038 ( .A1(n3682), .A2(n3681), .ZN(n6451) );
  INV_X1 U4039 ( .A(n6370), .ZN(n3681) );
  INV_X1 U4040 ( .A(n3699), .ZN(n3698) );
  CLKBUF_X1 U4041 ( .A(n6231), .Z(n6265) );
  NAND2_X1 U4042 ( .A1(n5148), .A2(n3692), .ZN(n3691) );
  INV_X1 U4043 ( .A(n5527), .ZN(n3692) );
  NAND2_X1 U4044 ( .A1(n3690), .A2(n5148), .ZN(n5654) );
  INV_X1 U4045 ( .A(n5490), .ZN(n3690) );
  NAND2_X1 U4046 ( .A1(n5579), .A2(n3712), .ZN(n3711) );
  INV_X1 U4047 ( .A(n4203), .ZN(n3713) );
  OAI21_X1 U4048 ( .B1(n7375), .B2(n7475), .A(n7376), .ZN(n4125) );
  INV_X1 U4049 ( .A(n5539), .ZN(n5534) );
  INV_X1 U4050 ( .A(n7530), .ZN(n6550) );
  NAND2_X1 U4051 ( .A1(n4086), .A2(n4085), .ZN(n5347) );
  OR2_X1 U4052 ( .A1(n6255), .A2(n4082), .ZN(n4086) );
  OR2_X1 U4053 ( .A1(n6064), .A2(n3934), .ZN(n7166) );
  NAND2_X1 U4054 ( .A1(n3883), .A2(n3882), .ZN(n3886) );
  AND2_X1 U4055 ( .A1(n3662), .A2(n5455), .ZN(n5460) );
  OR2_X1 U4056 ( .A1(n3645), .A2(n6375), .ZN(n6323) );
  OR2_X1 U4057 ( .A1(n5686), .A2(n3646), .ZN(n5512) );
  INV_X1 U4058 ( .A(n5864), .ZN(n5870) );
  INV_X1 U4059 ( .A(n3994), .ZN(n5449) );
  INV_X1 U4060 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5726) );
  INV_X1 U4061 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n5838) );
  NAND2_X1 U4062 ( .A1(n5885), .A2(n6322), .ZN(n5862) );
  INV_X1 U4063 ( .A(n6255), .ZN(n5732) );
  AOI21_X1 U4064 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5726), .A(n5808), .ZN(
        n5922) );
  INV_X1 U4065 ( .A(n5925), .ZN(n6375) );
  AND2_X1 U4066 ( .A1(n5590), .A2(n5343), .ZN(n7431) );
  INV_X1 U4067 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n7623) );
  INV_X1 U4068 ( .A(n7688), .ZN(n7633) );
  OR2_X1 U4069 ( .A1(n6279), .A2(n7696), .ZN(n7569) );
  OR2_X1 U4070 ( .A1(n6281), .A2(n5211), .ZN(n7686) );
  INV_X1 U4071 ( .A(n7686), .ZN(n7687) );
  INV_X1 U4072 ( .A(n6917), .ZN(n6914) );
  NAND2_X1 U4073 ( .A1(n4706), .A2(n5248), .ZN(n6925) );
  NAND2_X1 U4074 ( .A1(n4705), .A2(n5245), .ZN(n4706) );
  INV_X1 U4075 ( .A(n6952), .ZN(n7762) );
  AND2_X1 U4076 ( .A1(n6952), .A2(n6068), .ZN(n7763) );
  NAND2_X2 U4077 ( .A1(n6952), .A2(n6065), .ZN(n7751) );
  CLKBUF_X1 U4078 ( .A(n5705), .Z(n5617) );
  XNOR2_X1 U4079 ( .A(n5123), .B(n5122), .ZN(n6666) );
  OR2_X1 U4080 ( .A1(n5281), .A2(n5280), .ZN(n5123) );
  INV_X1 U4081 ( .A(n6925), .ZN(n6630) );
  INV_X1 U4082 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n7026) );
  INV_X1 U4083 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n7404) );
  NAND2_X1 U4084 ( .A1(n7701), .A2(n4709), .ZN(n7405) );
  CLKBUF_X1 U4085 ( .A(n5522), .Z(n5523) );
  OAI21_X1 U4086 ( .B1(n6574), .B2(n6573), .A(n6572), .ZN(n6575) );
  NAND2_X1 U4087 ( .A1(n3716), .A2(n3714), .ZN(n5222) );
  AOI21_X1 U4088 ( .B1(n3719), .B2(n3717), .A(n3715), .ZN(n3714) );
  XNOR2_X1 U4089 ( .A(n4271), .B(n4270), .ZN(n7081) );
  NAND2_X1 U4090 ( .A1(n3718), .A2(n4267), .ZN(n6955) );
  NAND2_X1 U4091 ( .A1(n6535), .A2(n3631), .ZN(n6536) );
  OAI21_X1 U4092 ( .B1(n6469), .B2(n3709), .A(n3664), .ZN(n7043) );
  NAND2_X1 U4093 ( .A1(n6469), .A2(n6470), .ZN(n3707) );
  OR2_X1 U4094 ( .A1(n7428), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7524) );
  NOR2_X1 U4095 ( .A1(n7492), .A2(n6521), .ZN(n7542) );
  NAND2_X1 U4096 ( .A1(n6220), .A2(n6221), .ZN(n3697) );
  INV_X1 U4097 ( .A(n7524), .ZN(n7544) );
  AND2_X1 U4098 ( .A1(n5428), .A2(n5413), .ZN(n7545) );
  AND2_X1 U4099 ( .A1(n5428), .A2(n5411), .ZN(n7557) );
  INV_X1 U4100 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n7193) );
  AND2_X1 U4101 ( .A1(n3662), .A2(n5466), .ZN(n5810) );
  AND2_X1 U4102 ( .A1(n5809), .A2(n5808), .ZN(n7251) );
  NOR2_X1 U4103 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n7713) );
  CLKBUF_X1 U4104 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n7181) );
  INV_X1 U4105 ( .A(n7218), .ZN(n7177) );
  INV_X1 U4106 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n7709) );
  NOR2_X1 U4107 ( .A1(n6645), .A2(n7706), .ZN(n7704) );
  INV_X1 U4108 ( .A(n6214), .ZN(n6186) );
  AOI22_X1 U4109 ( .A1(n6386), .A2(n6382), .B1(n6380), .B2(n6379), .ZN(n6448)
         );
  INV_X1 U4110 ( .A(n6374), .ZN(n6442) );
  NOR2_X1 U4111 ( .A1(n6072), .A2(n5808), .ZN(n6324) );
  NOR2_X1 U4112 ( .A1(n6071), .A2(n5808), .ZN(n6349) );
  NOR2_X1 U4113 ( .A1(n6088), .A2(n5808), .ZN(n6354) );
  NOR2_X1 U4114 ( .A1(n6091), .A2(n5808), .ZN(n6344) );
  NOR2_X1 U4115 ( .A1(n6944), .A2(n5808), .ZN(n6334) );
  NOR2_X1 U4116 ( .A1(n6086), .A2(n5808), .ZN(n6329) );
  AND2_X1 U4117 ( .A1(n5810), .A2(n6255), .ZN(n6114) );
  NOR2_X1 U4118 ( .A1(n6069), .A2(n5808), .ZN(n6360) );
  INV_X1 U4119 ( .A(n6349), .ZN(n6429) );
  INV_X1 U4120 ( .A(n6339), .ZN(n6436) );
  INV_X1 U4121 ( .A(n6354), .ZN(n6422) );
  INV_X1 U4122 ( .A(n6344), .ZN(n6415) );
  INV_X1 U4123 ( .A(n6329), .ZN(n6408) );
  INV_X1 U4124 ( .A(n6360), .ZN(n6401) );
  AND2_X1 U4125 ( .A1(n3980), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7711) );
  AOI21_X1 U4126 ( .B1(n6881), .B2(n7666), .A(n6693), .ZN(n6694) );
  OAI21_X1 U4127 ( .B1(n7069), .B2(n7693), .A(n3687), .ZN(U2797) );
  NAND2_X1 U4128 ( .A1(n6626), .A2(n3742), .ZN(n3688) );
  INV_X1 U4129 ( .A(n6922), .ZN(n3689) );
  INV_X1 U4130 ( .A(n5217), .ZN(n5218) );
  INV_X1 U4131 ( .A(n5337), .ZN(n5338) );
  OAI21_X1 U4132 ( .B1(n6705), .B2(n6917), .A(n5336), .ZN(n5337) );
  OAI21_X1 U4133 ( .B1(n6922), .B2(n7052), .A(n5291), .ZN(n5292) );
  NAND2_X2 U4134 ( .A1(n3739), .A2(n3908), .ZN(n3933) );
  OR2_X1 U4135 ( .A1(n6787), .A2(n3731), .ZN(n6901) );
  NOR2_X1 U4136 ( .A1(n5522), .A2(n3727), .ZN(n6005) );
  INV_X1 U4137 ( .A(n7033), .ZN(n4259) );
  AND2_X1 U4138 ( .A1(n3664), .A2(n3677), .ZN(n3665) );
  NAND2_X1 U4139 ( .A1(n3683), .A2(n5160), .ZN(n6264) );
  NOR2_X1 U4140 ( .A1(n7014), .A2(n3731), .ZN(n3666) );
  INV_X2 U4141 ( .A(n5592), .ZN(n5755) );
  AND2_X1 U4142 ( .A1(n5796), .A2(n5799), .ZN(n4004) );
  NAND2_X1 U4143 ( .A1(n3632), .A2(n4259), .ZN(n7024) );
  NAND2_X1 U4144 ( .A1(n6735), .A2(n6734), .ZN(n6720) );
  AND2_X1 U4145 ( .A1(n3766), .A2(n3767), .ZN(n4003) );
  NAND2_X1 U4146 ( .A1(n4061), .A2(n4060), .ZN(n4091) );
  AND2_X1 U4147 ( .A1(n3767), .A2(n5799), .ZN(n3891) );
  NAND2_X1 U4148 ( .A1(n3730), .A2(n3666), .ZN(n5107) );
  NAND4_X1 U4149 ( .A1(n3775), .A2(n3774), .A3(n3773), .A4(n3772), .ZN(n3957)
         );
  OR2_X1 U4150 ( .A1(n7395), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3668)
         );
  OAI21_X1 U4151 ( .B1(n7019), .B2(n4265), .A(n4264), .ZN(n6974) );
  AND2_X1 U4152 ( .A1(n3631), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3669)
         );
  NAND2_X1 U4153 ( .A1(n6725), .A2(n6724), .ZN(n6709) );
  NAND2_X1 U4154 ( .A1(n4252), .A2(n6514), .ZN(n3670) );
  AND4_X1 U4155 ( .A1(n3857), .A2(n3856), .A3(n3855), .A4(n3854), .ZN(n3898)
         );
  AND2_X1 U4156 ( .A1(n3765), .A2(n5799), .ZN(n4025) );
  NAND2_X1 U4157 ( .A1(n4069), .A2(n4068), .ZN(n3671) );
  INV_X1 U4158 ( .A(n6680), .ZN(n5298) );
  NAND2_X1 U4159 ( .A1(n6833), .A2(n6832), .ZN(n6820) );
  AND2_X1 U4160 ( .A1(n6518), .A2(n5179), .ZN(n6813) );
  NAND2_X1 U4161 ( .A1(n6833), .A2(n3734), .ZN(n6800) );
  NAND2_X1 U4162 ( .A1(n5579), .A2(n4203), .ZN(n7394) );
  NAND2_X1 U4163 ( .A1(n3697), .A2(n4251), .ZN(n6268) );
  NAND2_X1 U4164 ( .A1(n3696), .A2(n3695), .ZN(n6462) );
  NAND2_X1 U4165 ( .A1(n3707), .A2(n4257), .ZN(n6513) );
  AND2_X1 U4166 ( .A1(n6518), .A2(n3679), .ZN(n6795) );
  NAND2_X1 U4167 ( .A1(n3728), .A2(n4332), .ZN(n5521) );
  INV_X1 U4168 ( .A(n3965), .ZN(n5295) );
  AND2_X1 U4169 ( .A1(n3679), .A2(n6796), .ZN(n3672) );
  AND2_X1 U4170 ( .A1(n6896), .A2(n5192), .ZN(n6898) );
  INV_X1 U4171 ( .A(n5522), .ZN(n3728) );
  AND2_X1 U4172 ( .A1(n3729), .A2(n6230), .ZN(n3673) );
  NAND2_X1 U4173 ( .A1(n6518), .A2(n3672), .ZN(n6794) );
  AND2_X1 U4174 ( .A1(n4252), .A2(n7149), .ZN(n3674) );
  AND2_X1 U4175 ( .A1(n5178), .A2(n5177), .ZN(n6828) );
  NAND2_X1 U4176 ( .A1(n4252), .A2(n5321), .ZN(n3675) );
  AND2_X1 U4177 ( .A1(n3711), .A2(n3668), .ZN(n3676) );
  OR2_X1 U4178 ( .A1(n5404), .A2(n7200), .ZN(n7701) );
  INV_X1 U4179 ( .A(n7701), .ZN(n7422) );
  NAND2_X1 U4180 ( .A1(n5534), .A2(n5142), .ZN(n5498) );
  AND2_X1 U4181 ( .A1(n5526), .A2(n6008), .ZN(n6007) );
  OR2_X1 U4182 ( .A1(n4252), .A2(n7514), .ZN(n3677) );
  NAND3_X1 U4183 ( .A1(n5417), .A2(n3990), .A3(n3989), .ZN(n5423) );
  INV_X1 U4184 ( .A(n6264), .ZN(n3682) );
  NAND2_X1 U4185 ( .A1(n5491), .A2(n5492), .ZN(n5490) );
  INV_X1 U4186 ( .A(n6629), .ZN(n3686) );
  NOR2_X1 U4187 ( .A1(n5564), .A2(n3956), .ZN(n3678) );
  NAND2_X1 U4188 ( .A1(n6645), .A2(n5445), .ZN(n5564) );
  AND2_X2 U4189 ( .A1(n3720), .A2(n3751), .ZN(n3767) );
  AND2_X2 U4190 ( .A1(n4279), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3766)
         );
  NAND2_X1 U4191 ( .A1(n6220), .A2(n3698), .ZN(n3696) );
  NAND2_X1 U4192 ( .A1(n3701), .A2(n3671), .ZN(n3702) );
  NAND2_X1 U4193 ( .A1(n4062), .A2(n4091), .ZN(n3701) );
  NAND3_X1 U4194 ( .A1(n4062), .A2(n4091), .A3(n4070), .ZN(n4092) );
  NAND2_X1 U4195 ( .A1(n6469), .A2(n3665), .ZN(n3706) );
  NAND2_X1 U4196 ( .A1(n4260), .A2(n3710), .ZN(n6980) );
  NAND3_X1 U4197 ( .A1(n3711), .A2(n3668), .A3(n6052), .ZN(n4241) );
  NAND2_X1 U4198 ( .A1(n3941), .A2(n3721), .ZN(n3723) );
  INV_X1 U4199 ( .A(n3954), .ZN(n3722) );
  NAND3_X1 U4200 ( .A1(n5803), .A2(n3723), .A3(n5412), .ZN(n3949) );
  OAI211_X1 U4201 ( .C1(n7081), .C2(n7701), .A(n3724), .B(n4714), .ZN(U2958)
         );
  NAND2_X1 U4202 ( .A1(n6630), .A2(n7421), .ZN(n3724) );
  INV_X1 U4203 ( .A(n5522), .ZN(n3726) );
  INV_X1 U4204 ( .A(n6787), .ZN(n3730) );
  NOR2_X1 U4205 ( .A1(n6787), .A2(n4515), .ZN(n6900) );
  OR2_X1 U4206 ( .A1(n6570), .A2(n4269), .ZN(n4271) );
  AND2_X2 U4207 ( .A1(n3847), .A2(n3994), .ZN(n3746) );
  AOI22_X1 U4208 ( .A1(n3648), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3903), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3923) );
  OR2_X1 U4209 ( .A1(n5104), .A2(n5103), .ZN(n3737) );
  AND2_X1 U4210 ( .A1(DATAI_3_), .A2(keyinput_156), .ZN(n3738) );
  AND4_X1 U4211 ( .A1(n3902), .A2(n3901), .A3(n3900), .A4(n3899), .ZN(n3739)
         );
  AND4_X1 U4212 ( .A1(n3930), .A2(n3929), .A3(n3928), .A4(n3927), .ZN(n3740)
         );
  AND3_X1 U4213 ( .A1(n4831), .A2(n4830), .A3(n4829), .ZN(n3741) );
  OR2_X1 U4214 ( .A1(n6692), .A2(n7337), .ZN(n3742) );
  OR2_X1 U4215 ( .A1(n4252), .A2(n6529), .ZN(n3743) );
  INV_X1 U4216 ( .A(n6760), .ZN(n4610) );
  OR2_X1 U4217 ( .A1(n4895), .A2(n4894), .ZN(n3744) );
  OR2_X1 U4218 ( .A1(n7336), .A2(keyinput_199), .ZN(n3745) );
  OR2_X1 U4219 ( .A1(n7433), .A2(STATE_REG_0__SCAN_IN), .ZN(n7746) );
  NOR2_X1 U4220 ( .A1(n5795), .A2(n5794), .ZN(n7190) );
  INV_X1 U4221 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n7198) );
  OR2_X1 U4222 ( .A1(STATEBS16_REG_SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n4665) );
  AND2_X2 U4223 ( .A1(n5762), .A2(n5796), .ZN(n3903) );
  NOR4_X1 U4224 ( .A1(n4727), .A2(n4726), .A3(n4725), .A4(n4724), .ZN(n4730)
         );
  OAI22_X1 U4225 ( .A1(n4745), .A2(n4744), .B1(DATAI_17_), .B2(keyinput_142), 
        .ZN(n4746) );
  INV_X1 U4226 ( .A(n4746), .ZN(n4747) );
  OAI22_X1 U4227 ( .A1(n6950), .A2(n4752), .B1(DATAI_15_), .B2(keyinput_144), 
        .ZN(n4753) );
  INV_X1 U4228 ( .A(n4753), .ZN(n4754) );
  NOR2_X1 U4229 ( .A1(keyinput_156), .A2(DATAI_3_), .ZN(n4770) );
  NOR2_X1 U4230 ( .A1(n3738), .A2(n4770), .ZN(n4771) );
  XNOR2_X1 U4231 ( .A(n7735), .B(keyinput_164), .ZN(n4780) );
  AOI21_X1 U4232 ( .B1(n4782), .B2(n4781), .A(n4780), .ZN(n4783) );
  XNOR2_X1 U4233 ( .A(keyinput_179), .B(REIP_REG_31__SCAN_IN), .ZN(n4802) );
  OAI21_X1 U4234 ( .B1(n4803), .B2(n4802), .A(n4801), .ZN(n4806) );
  INV_X1 U4235 ( .A(keyinput_187), .ZN(n4812) );
  XNOR2_X1 U4236 ( .A(n7322), .B(n4812), .ZN(n4813) );
  NAND2_X1 U4237 ( .A1(n4814), .A2(n4813), .ZN(n4815) );
  INV_X1 U4238 ( .A(n4828), .ZN(n4829) );
  NAND2_X1 U4239 ( .A1(n7336), .A2(keyinput_199), .ZN(n4832) );
  NAND2_X1 U4240 ( .A1(n3745), .A2(n4832), .ZN(n4833) );
  AOI21_X1 U4241 ( .B1(n4834), .B2(n3741), .A(n4833), .ZN(n4836) );
  AOI22_X1 U4242 ( .A1(n4840), .A2(n4839), .B1(n7324), .B2(keyinput_205), .ZN(
        n4843) );
  NAND2_X1 U4243 ( .A1(keyinput_214), .A2(ADDRESS_REG_14__SCAN_IN), .ZN(n4852)
         );
  NAND2_X1 U4244 ( .A1(n4853), .A2(n4852), .ZN(n4854) );
  AOI21_X1 U4245 ( .B1(n4856), .B2(n4855), .A(n4854), .ZN(n4870) );
  NOR4_X1 U4246 ( .A1(n4870), .A2(n4869), .A3(n4868), .A4(n4867), .ZN(n4875)
         );
  XNOR2_X1 U4247 ( .A(DATAWIDTH_REG_7__SCAN_IN), .B(keyinput_239), .ZN(n4887)
         );
  NAND2_X1 U4248 ( .A1(n3937), .A2(n4074), .ZN(n3962) );
  XNOR2_X1 U4249 ( .A(DATAWIDTH_REG_11__SCAN_IN), .B(keyinput_243), .ZN(n4894)
         );
  OAI21_X1 U4250 ( .B1(n3860), .B2(n3937), .A(n3962), .ZN(n3963) );
  NAND2_X1 U4251 ( .A1(n3903), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3820)
         );
  NAND2_X1 U4252 ( .A1(n3937), .A2(n3983), .ZN(n3966) );
  INV_X1 U4253 ( .A(n5655), .ZN(n4323) );
  OR2_X1 U4254 ( .A1(n4215), .A2(n4214), .ZN(n4234) );
  OAI21_X1 U4255 ( .B1(n4146), .B2(n3877), .A(n3876), .ZN(n3878) );
  AOI21_X1 U4256 ( .B1(n4099), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3839), 
        .ZN(n3837) );
  OR2_X1 U4257 ( .A1(n3850), .A2(n3861), .ZN(n3852) );
  INV_X1 U4258 ( .A(keyinput_250), .ZN(n4904) );
  NAND2_X1 U4259 ( .A1(n4352), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3752)
         );
  INV_X1 U4260 ( .A(n5524), .ZN(n4332) );
  INV_X1 U4261 ( .A(n6266), .ZN(n5160) );
  INV_X1 U4262 ( .A(n5538), .ZN(n5142) );
  XNOR2_X1 U4263 ( .A(n4904), .B(DATAWIDTH_REG_18__SCAN_IN), .ZN(n4905) );
  INV_X1 U4264 ( .A(n6903), .ZN(n4515) );
  NAND2_X1 U4265 ( .A1(n4172), .A2(n4171), .ZN(n4181) );
  OR2_X1 U4266 ( .A1(n4641), .A2(n4640), .ZN(n4651) );
  INV_X1 U4267 ( .A(n7166), .ZN(n4466) );
  NOR2_X1 U4268 ( .A1(n3933), .A2(n5838), .ZN(n4283) );
  INV_X1 U4269 ( .A(n6828), .ZN(n5179) );
  AND2_X1 U4270 ( .A1(n5164), .A2(n5163), .ZN(n6370) );
  NAND2_X1 U4271 ( .A1(n4116), .A2(n4115), .ZN(n4156) );
  NAND2_X1 U4272 ( .A1(n3834), .A2(n7709), .ZN(n5115) );
  AND2_X1 U4273 ( .A1(n4906), .A2(n4905), .ZN(n4907) );
  NAND2_X1 U4274 ( .A1(n4902), .A2(n4901), .ZN(n4908) );
  AND2_X1 U4275 ( .A1(n7563), .A2(REIP_REG_5__SCAN_IN), .ZN(n7599) );
  AND2_X1 U4276 ( .A1(n5153), .A2(n5152), .ZN(n5527) );
  OR2_X1 U4277 ( .A1(n4700), .A2(n6959), .ZN(n4701) );
  INV_X1 U4278 ( .A(n5278), .ZN(n5236) );
  INV_X1 U4279 ( .A(n4283), .ZN(n4548) );
  INV_X1 U4280 ( .A(n6897), .ZN(n5192) );
  AND2_X1 U4281 ( .A1(n4252), .A2(n7516), .ZN(n7033) );
  AND2_X1 U4282 ( .A1(n5688), .A2(n3640), .ZN(n6374) );
  NAND2_X1 U4283 ( .A1(n4135), .A2(n4134), .ZN(n5865) );
  AND2_X1 U4284 ( .A1(n3663), .A2(n7169), .ZN(n5844) );
  INV_X1 U4285 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6824) );
  INV_X1 U4286 ( .A(n7677), .ZN(n7648) );
  AND2_X1 U4287 ( .A1(n5124), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5125) );
  OR3_X1 U4288 ( .A1(n6281), .A2(n5205), .A3(n5209), .ZN(n6808) );
  OR2_X1 U4289 ( .A1(n7369), .A2(n6699), .ZN(n5336) );
  AND2_X1 U4290 ( .A1(n3933), .A2(n3937), .ZN(n6066) );
  NOR2_X1 U4291 ( .A1(n4644), .A2(n6750), .ZN(n4648) );
  INV_X1 U4292 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6848) );
  NAND2_X1 U4293 ( .A1(n6593), .A2(n6592), .ZN(n6594) );
  INV_X1 U4294 ( .A(n5320), .ZN(n5332) );
  AND2_X1 U4295 ( .A1(n7032), .A2(n4261), .ZN(n4262) );
  OR2_X1 U4296 ( .A1(n5404), .A2(n5403), .ZN(n5405) );
  NOR2_X1 U4297 ( .A1(n5909), .A2(n3646), .ZN(n5733) );
  INV_X1 U4298 ( .A(n6314), .ZN(n6363) );
  OR2_X1 U4299 ( .A1(n3662), .A2(n3640), .ZN(n5909) );
  NAND2_X1 U4300 ( .A1(n3662), .A2(n5434), .ZN(n5444) );
  INV_X1 U4301 ( .A(n5808), .ZN(n5885) );
  OAI211_X1 U4302 ( .C1(n3836), .C2(n4048), .A(n4047), .B(n4046), .ZN(n4079)
         );
  OR2_X1 U4303 ( .A1(n3621), .A2(n6374), .ZN(n6376) );
  OR2_X1 U4304 ( .A1(n5634), .A2(n6255), .ZN(n6047) );
  AND2_X1 U4305 ( .A1(n7715), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3980) );
  OR2_X1 U4306 ( .A1(n6281), .A2(n6882), .ZN(n6687) );
  NAND2_X1 U4307 ( .A1(n4534), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4570)
         );
  AND2_X1 U4308 ( .A1(n6871), .A2(n5125), .ZN(n7696) );
  NOR2_X1 U4309 ( .A1(n6843), .A2(n7428), .ZN(n7677) );
  INV_X1 U4310 ( .A(n7369), .ZN(n6913) );
  INV_X1 U4311 ( .A(n6063), .ZN(n5708) );
  INV_X1 U4312 ( .A(n7420), .ZN(n7756) );
  INV_X1 U4313 ( .A(n7425), .ZN(n7409) );
  NOR2_X1 U4314 ( .A1(n4293), .A2(n6858), .ZN(n4304) );
  INV_X1 U4315 ( .A(n5319), .ZN(n6723) );
  OR2_X1 U4316 ( .A1(n7528), .A2(n6550), .ZN(n7508) );
  INV_X1 U4317 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n7715) );
  AND2_X1 U4318 ( .A1(n5790), .A2(STATE2_REG_3__SCAN_IN), .ZN(n7218) );
  OAI21_X1 U4319 ( .B1(n5889), .B2(n5888), .A(n5887), .ZN(n6002) );
  AND2_X1 U4320 ( .A1(n5733), .A2(n6255), .ZN(n6214) );
  INV_X1 U4321 ( .A(n6212), .ZN(n6365) );
  NOR2_X1 U4322 ( .A1(n5909), .A2(n5858), .ZN(n6195) );
  AND2_X1 U4323 ( .A1(n5460), .A2(n6255), .ZN(n6148) );
  INV_X1 U4324 ( .A(n5947), .ZN(n6097) );
  NAND2_X1 U4325 ( .A1(n5885), .A2(n5884), .ZN(n6384) );
  INV_X1 U4326 ( .A(n6117), .ZN(n6163) );
  OR3_X1 U4327 ( .A1(n5820), .A2(n5862), .A3(n5819), .ZN(n6110) );
  NOR2_X1 U4328 ( .A1(n6085), .A2(n5808), .ZN(n6339) );
  INV_X1 U4329 ( .A(n4665), .ZN(n5282) );
  INV_X1 U4330 ( .A(STATE_REG_2__SCAN_IN), .ZN(n7737) );
  INV_X1 U4331 ( .A(STATE_REG_1__SCAN_IN), .ZN(n7433) );
  OR2_X1 U4332 ( .A1(n5404), .A2(n5111), .ZN(n5590) );
  INV_X1 U4333 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n7726) );
  OR2_X1 U4334 ( .A1(n6687), .A2(n5126), .ZN(n7693) );
  INV_X1 U4335 ( .A(n7569), .ZN(n6879) );
  NOR2_X2 U4336 ( .A1(n7759), .A2(n7763), .ZN(n6953) );
  INV_X1 U4337 ( .A(n7255), .ZN(n7286) );
  NAND2_X1 U4338 ( .A1(n5593), .A2(n5591), .ZN(n6063) );
  NAND2_X1 U4339 ( .A1(n5925), .A2(n4707), .ZN(n7052) );
  NAND2_X1 U4340 ( .A1(n7405), .A2(n5348), .ZN(n7425) );
  INV_X1 U4341 ( .A(n7545), .ZN(n7555) );
  INV_X1 U4342 ( .A(n7557), .ZN(n7506) );
  INV_X1 U4343 ( .A(n5731), .ZN(n6217) );
  INV_X1 U4344 ( .A(n6195), .ZN(n6151) );
  NAND2_X1 U4345 ( .A1(n5460), .A2(n5732), .ZN(n6026) );
  AND2_X1 U4346 ( .A1(n5663), .A2(n5662), .ZN(n6031) );
  NAND2_X1 U4347 ( .A1(n5435), .A2(n5732), .ZN(n6095) );
  NAND2_X1 U4348 ( .A1(n5504), .A2(n6255), .ZN(n5947) );
  INV_X1 U4349 ( .A(n6324), .ZN(n6447) );
  INV_X1 U4350 ( .A(n6334), .ZN(n6394) );
  OR2_X1 U4351 ( .A1(n5686), .A2(n5858), .ZN(n6117) );
  NAND2_X1 U4352 ( .A1(n5810), .A2(n5732), .ZN(n6143) );
  AND2_X1 U4353 ( .A1(n5922), .A2(n5633), .ZN(n6051) );
  CLKBUF_X1 U4354 ( .A(n7230), .Z(n7729) );
  OAI21_X1 U4355 ( .B1(n6640), .B2(n6919), .A(n5338), .ZN(U2830) );
  NAND2_X1 U4356 ( .A1(n7193), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3748) );
  NAND2_X1 U4357 ( .A1(n3725), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3747) );
  NAND2_X1 U4358 ( .A1(n3748), .A2(n3747), .ZN(n3850) );
  NAND2_X1 U4359 ( .A1(n3852), .A2(n3748), .ZN(n3840) );
  MUX2_X1 U4360 ( .A(n4099), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n3841) );
  MUX2_X1 U4361 ( .A(n7198), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(n7181), 
        .Z(n3838) );
  INV_X1 U4362 ( .A(n3838), .ZN(n3749) );
  AOI222_X1 U4363 ( .A1(n3833), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B1(
        n3833), .B2(n7709), .C1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n7709), 
        .ZN(n5117) );
  AND2_X4 U4364 ( .A1(n3766), .A2(n5796), .ZN(n4032) );
  NAND2_X1 U4365 ( .A1(n3659), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3755)
         );
  NAND2_X1 U4366 ( .A1(n3652), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3754)
         );
  NAND2_X1 U4367 ( .A1(n4025), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3753) );
  NAND2_X1 U4368 ( .A1(n5258), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3759) );
  NAND2_X1 U4369 ( .A1(n3622), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3758) );
  NAND2_X1 U4370 ( .A1(n4351), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3757) );
  AND2_X4 U4371 ( .A1(n3767), .A2(n5762), .ZN(n3922) );
  NAND2_X1 U4372 ( .A1(n3657), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3756) );
  NAND2_X1 U4373 ( .A1(n4104), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3764) );
  NAND2_X1 U4374 ( .A1(n3650), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3763) );
  NAND2_X1 U4375 ( .A1(n3639), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3762) );
  NAND2_X1 U4376 ( .A1(n4004), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3761)
         );
  NAND2_X1 U4377 ( .A1(n4020), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3771) );
  NAND2_X1 U4378 ( .A1(n3654), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3770)
         );
  NAND2_X1 U4379 ( .A1(n3903), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3769)
         );
  NAND2_X1 U4380 ( .A1(n3891), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3768) );
  NAND2_X1 U4381 ( .A1(n3623), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3779) );
  NAND2_X1 U4382 ( .A1(n3891), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3778) );
  NAND2_X1 U4383 ( .A1(n4351), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3777) );
  NAND2_X1 U4384 ( .A1(n3654), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3776)
         );
  NAND2_X1 U4385 ( .A1(n3652), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3783)
         );
  NAND2_X1 U4386 ( .A1(n4104), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3782) );
  NAND2_X1 U4387 ( .A1(n3643), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3781)
         );
  NAND2_X1 U4388 ( .A1(n3660), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3780)
         );
  NAND2_X1 U4389 ( .A1(n4025), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3787) );
  NAND2_X1 U4390 ( .A1(n4552), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3786) );
  NAND2_X1 U4391 ( .A1(n3639), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3785) );
  NAND2_X1 U4392 ( .A1(n4004), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3784)
         );
  NAND2_X1 U4393 ( .A1(n4020), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3791) );
  NAND2_X1 U4394 ( .A1(n3648), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3790) );
  NAND2_X1 U4395 ( .A1(n3903), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3789)
         );
  NAND2_X1 U4396 ( .A1(n3656), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3788) );
  NAND2_X1 U4397 ( .A1(n5117), .A2(n4229), .ZN(n3883) );
  NAND2_X1 U4398 ( .A1(n3648), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3799) );
  NAND2_X1 U4399 ( .A1(n4020), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3798) );
  NAND2_X1 U4400 ( .A1(n3903), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3797)
         );
  NAND2_X1 U4401 ( .A1(n3655), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3796) );
  NAND2_X1 U4402 ( .A1(n4104), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3803) );
  NAND2_X1 U4403 ( .A1(n3628), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3802)
         );
  NAND2_X1 U4404 ( .A1(n4352), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3801)
         );
  NAND2_X1 U4405 ( .A1(n3658), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3800)
         );
  NAND2_X1 U4406 ( .A1(n3650), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3807) );
  NAND2_X1 U4407 ( .A1(n4025), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3806) );
  NAND2_X1 U4408 ( .A1(n3639), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3805) );
  NAND2_X1 U4409 ( .A1(n4004), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3804)
         );
  NAND2_X1 U4410 ( .A1(n3627), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3811)
         );
  NAND2_X1 U4411 ( .A1(n3623), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3810) );
  NAND2_X1 U4412 ( .A1(n3921), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3809) );
  NAND2_X1 U4413 ( .A1(n3891), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3808) );
  NAND4_X2 U4414 ( .A1(n3857), .A2(n3856), .A3(n3855), .A4(n3854), .ZN(n4074)
         );
  NAND2_X1 U4415 ( .A1(n3623), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3815) );
  NAND2_X1 U4416 ( .A1(n3653), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3814)
         );
  NAND2_X1 U4417 ( .A1(n4689), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3813) );
  NAND2_X1 U4418 ( .A1(n3891), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3812) );
  NAND2_X1 U4419 ( .A1(n3651), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3819)
         );
  NAND2_X1 U4420 ( .A1(n4104), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3818) );
  NAND2_X1 U4421 ( .A1(n3643), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3817)
         );
  NAND2_X1 U4422 ( .A1(n3659), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3816)
         );
  NAND2_X1 U4423 ( .A1(n3922), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3821) );
  NAND2_X1 U4424 ( .A1(n4020), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3822) );
  NAND2_X1 U4425 ( .A1(n3823), .A2(n3822), .ZN(n3824) );
  AOI21_X2 U4426 ( .B1(n3648), .B2(INSTQUEUE_REG_7__1__SCAN_IN), .A(n3824), 
        .ZN(n3830) );
  NAND2_X1 U4427 ( .A1(n4025), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3828) );
  NAND2_X1 U4428 ( .A1(n3650), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3827) );
  NAND2_X1 U4429 ( .A1(n3639), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3826) );
  NAND2_X1 U4430 ( .A1(n4004), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3825)
         );
  OAI22_X1 U4431 ( .A1(n5115), .A2(n3836), .B1(STATE2_REG_0__SCAN_IN), .B2(
        n7709), .ZN(n3835) );
  INV_X1 U4432 ( .A(n3835), .ZN(n3879) );
  XOR2_X1 U4433 ( .A(n3838), .B(n3837), .Z(n5112) );
  INV_X1 U4434 ( .A(n3839), .ZN(n3845) );
  INV_X1 U4435 ( .A(n3840), .ZN(n3843) );
  INV_X1 U4436 ( .A(n3841), .ZN(n3842) );
  NAND2_X1 U4437 ( .A1(n3843), .A2(n3842), .ZN(n3844) );
  NAND2_X1 U4438 ( .A1(n3845), .A2(n3844), .ZN(n5113) );
  INV_X1 U4439 ( .A(n5113), .ZN(n3846) );
  NAND2_X1 U4440 ( .A1(n3956), .A2(n4074), .ZN(n3848) );
  INV_X1 U4441 ( .A(n3872), .ZN(n3849) );
  AOI211_X1 U4442 ( .C1(n4146), .C2(n5113), .A(n3871), .B(n3849), .ZN(n3875)
         );
  NAND2_X1 U4443 ( .A1(n3850), .A2(n3861), .ZN(n3851) );
  NAND2_X1 U4444 ( .A1(n3852), .A2(n3851), .ZN(n5114) );
  INV_X1 U4445 ( .A(n3884), .ZN(n3853) );
  OAI21_X1 U4446 ( .B1(n7437), .B2(n5114), .A(n3853), .ZN(n3870) );
  AOI21_X1 U4447 ( .B1(n4146), .B2(n5114), .A(n6067), .ZN(n3858) );
  OAI21_X1 U4448 ( .B1(n3956), .B2(n3859), .A(n3858), .ZN(n3869) );
  NAND2_X1 U4449 ( .A1(n4045), .A2(n4074), .ZN(n5407) );
  INV_X1 U4450 ( .A(n5407), .ZN(n3955) );
  OAI21_X1 U4451 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5726), .A(n3861), 
        .ZN(n3863) );
  OAI21_X1 U4452 ( .B1(n3955), .B2(n3863), .A(n3862), .ZN(n3867) );
  NOR2_X1 U4453 ( .A1(n3870), .A2(n3869), .ZN(n3866) );
  INV_X1 U4454 ( .A(n3863), .ZN(n3864) );
  AOI21_X1 U4455 ( .B1(n4229), .B2(n3864), .A(n3884), .ZN(n3865) );
  AOI211_X1 U4456 ( .C1(n3872), .C2(n3867), .A(n3866), .B(n3865), .ZN(n3868)
         );
  AOI21_X1 U4457 ( .B1(n3870), .B2(n3869), .A(n3868), .ZN(n3874) );
  INV_X1 U4458 ( .A(n3871), .ZN(n3873) );
  OAI222_X1 U4459 ( .A1(n3877), .A2(n4082), .B1(n3875), .B2(n3874), .C1(n3873), 
        .C2(n3872), .ZN(n3876) );
  AOI222_X1 U4460 ( .A1(n3880), .A2(n3879), .B1(n3880), .B2(n3878), .C1(n3879), 
        .C2(n3878), .ZN(n3881) );
  INV_X1 U4461 ( .A(n3881), .ZN(n3882) );
  NAND2_X1 U4462 ( .A1(n5117), .A2(n3884), .ZN(n3885) );
  AOI22_X1 U4463 ( .A1(n4104), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4397), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4464 ( .A1(n3644), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4032), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4465 ( .A1(n4025), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4004), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3887) );
  AND4_X2 U4466 ( .A1(n3890), .A2(n3889), .A3(n3888), .A4(n3887), .ZN(n3897)
         );
  AOI22_X1 U4467 ( .A1(n3647), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3903), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4468 ( .A1(n3915), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3891), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4469 ( .A1(n4020), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3922), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4470 ( .A1(n4009), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3892) );
  NAND2_X1 U4471 ( .A1(n3937), .A2(n3898), .ZN(n3909) );
  AOI22_X1 U4472 ( .A1(n4020), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5258), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3902) );
  AOI22_X1 U4473 ( .A1(n4351), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3628), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3901) );
  AOI22_X1 U4474 ( .A1(n4552), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3639), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4475 ( .A1(n3659), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4004), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3899) );
  AOI22_X1 U4476 ( .A1(n3657), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3903), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4477 ( .A1(n3622), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3891), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4478 ( .A1(n3644), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4479 ( .A1(n3627), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4104), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3904) );
  AND2_X2 U4480 ( .A1(n3909), .A2(n3933), .ZN(n3939) );
  NAND3_X1 U4481 ( .A1(n4045), .A2(n4074), .A3(n5446), .ZN(n3910) );
  NAND2_X1 U4482 ( .A1(n3939), .A2(n3910), .ZN(n3997) );
  AOI22_X1 U4483 ( .A1(n4020), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3657), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4484 ( .A1(n3639), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4004), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4485 ( .A1(n4689), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4488), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4486 ( .A1(n3652), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4487 ( .A1(n3622), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3653), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3919) );
  AOI22_X1 U4488 ( .A1(n4552), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4489 ( .A1(n4104), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3643), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4490 ( .A1(n3648), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3903), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3916) );
  NAND2_X2 U4491 ( .A1(n3667), .A2(n3920), .ZN(n3983) );
  AOI22_X1 U4492 ( .A1(n3623), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3891), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3926) );
  AOI22_X1 U4493 ( .A1(n3653), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3925) );
  AOI22_X1 U4494 ( .A1(n4020), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3657), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3924) );
  AOI22_X1 U4495 ( .A1(n3651), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4104), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4496 ( .A1(n3643), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3659), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4497 ( .A1(n4552), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3639), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4498 ( .A1(n4025), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4004), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3927) );
  NAND2_X1 U4499 ( .A1(n3961), .A2(n3994), .ZN(n3932) );
  NAND2_X2 U4500 ( .A1(n5446), .A2(n4074), .ZN(n6064) );
  AND2_X1 U4501 ( .A1(n3933), .A2(n3860), .ZN(n3990) );
  INV_X1 U4502 ( .A(n3990), .ZN(n3934) );
  NAND2_X1 U4503 ( .A1(n7166), .A2(n5563), .ZN(n3936) );
  NAND2_X1 U4504 ( .A1(n3953), .A2(n3936), .ZN(n5761) );
  OR2_X1 U4505 ( .A1(n5761), .A2(n5407), .ZN(n7200) );
  NAND2_X1 U4506 ( .A1(n3961), .A2(n5446), .ZN(n3938) );
  NAND3_X1 U4507 ( .A1(n3940), .A2(n5295), .A3(n6064), .ZN(n5366) );
  INV_X1 U4508 ( .A(n5366), .ZN(n3941) );
  NAND2_X1 U4509 ( .A1(n7737), .A2(STATE_REG_1__SCAN_IN), .ZN(n7739) );
  NAND2_X1 U4510 ( .A1(n7433), .A2(STATE_REG_2__SCAN_IN), .ZN(n3942) );
  NAND2_X1 U4511 ( .A1(n7739), .A2(n3942), .ZN(n5203) );
  NOR2_X1 U4512 ( .A1(n5591), .A2(n5203), .ZN(n3954) );
  INV_X1 U4513 ( .A(n3966), .ZN(n3943) );
  NAND3_X1 U4514 ( .A1(n5295), .A2(n3944), .A3(n3943), .ZN(n5118) );
  INV_X1 U4515 ( .A(n3946), .ZN(n6681) );
  NAND2_X1 U4516 ( .A1(n3947), .A2(n6681), .ZN(n5758) );
  INV_X1 U4517 ( .A(n5758), .ZN(n3948) );
  NAND2_X1 U4518 ( .A1(n3948), .A2(n6066), .ZN(n5412) );
  NAND2_X1 U4519 ( .A1(n3949), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3977) );
  NAND2_X1 U4520 ( .A1(n7713), .A2(n7437), .ZN(n4708) );
  NAND2_X1 U4521 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4100) );
  NOR2_X1 U4522 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5943) );
  INV_X1 U4523 ( .A(n5943), .ZN(n3950) );
  NAND2_X1 U4524 ( .A1(n4100), .A2(n3950), .ZN(n5837) );
  OR2_X1 U4525 ( .A1(n4708), .A2(n5837), .ZN(n3952) );
  INV_X1 U4526 ( .A(n3980), .ZN(n4132) );
  NAND2_X1 U4527 ( .A1(n4132), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3951) );
  OAI21_X1 U4528 ( .B1(n3954), .B2(n4074), .A(n3953), .ZN(n3960) );
  NAND2_X1 U4529 ( .A1(n3955), .A2(n3746), .ZN(n3987) );
  NAND2_X1 U4530 ( .A1(n3965), .A2(n3958), .ZN(n3988) );
  NAND2_X1 U4531 ( .A1(n3987), .A2(n3988), .ZN(n3959) );
  NOR2_X1 U4532 ( .A1(n3960), .A2(n3959), .ZN(n3970) );
  NAND2_X1 U4533 ( .A1(n3961), .A2(n3933), .ZN(n3964) );
  NOR2_X1 U4534 ( .A1(n3964), .A2(n3963), .ZN(n3968) );
  NOR2_X1 U4535 ( .A1(n3966), .A2(n3965), .ZN(n3967) );
  OAI21_X1 U4536 ( .B1(n3968), .B2(n3967), .A(n3991), .ZN(n3969) );
  NAND2_X1 U4537 ( .A1(n3969), .A2(n5563), .ZN(n3986) );
  NAND2_X1 U4538 ( .A1(n3970), .A2(n3986), .ZN(n3971) );
  NAND2_X1 U4539 ( .A1(n3971), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3973) );
  NAND2_X1 U4540 ( .A1(n4146), .A2(n6064), .ZN(n3972) );
  NAND2_X1 U4541 ( .A1(n4098), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3974) );
  NAND2_X1 U4542 ( .A1(n3975), .A2(n3974), .ZN(n4096) );
  INV_X1 U4543 ( .A(n3976), .ZN(n3978) );
  OAI21_X1 U4544 ( .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n3978), .A(n3629), 
        .ZN(n3979) );
  NAND2_X1 U4545 ( .A1(n4098), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3982) );
  MUX2_X1 U4546 ( .A(n4708), .B(n3980), .S(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .Z(n3981) );
  NAND2_X2 U4547 ( .A1(n3982), .A2(n3981), .ZN(n4019) );
  NOR2_X1 U4548 ( .A1(n5407), .A2(n3956), .ZN(n3985) );
  NAND2_X1 U4549 ( .A1(n3983), .A2(n6280), .ZN(n3984) );
  OAI21_X1 U4550 ( .B1(n3986), .B2(n3985), .A(n3984), .ZN(n5422) );
  AND2_X1 U4551 ( .A1(n3988), .A2(n3987), .ZN(n4000) );
  NOR2_X1 U4552 ( .A1(n3983), .A2(n6280), .ZN(n5417) );
  NOR2_X1 U4553 ( .A1(n3937), .A2(n3994), .ZN(n3989) );
  NAND2_X1 U4554 ( .A1(n3991), .A2(n6280), .ZN(n3993) );
  AND2_X1 U4555 ( .A1(n7713), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3992) );
  NAND2_X1 U4556 ( .A1(n6064), .A2(n3860), .ZN(n3995) );
  NAND2_X1 U4557 ( .A1(n3995), .A2(n3994), .ZN(n3996) );
  OAI21_X1 U4558 ( .B1(n3997), .B2(n3996), .A(n5591), .ZN(n3998) );
  NAND3_X1 U4559 ( .A1(n4000), .A2(n3999), .A3(n3998), .ZN(n4001) );
  INV_X1 U4560 ( .A(n4018), .ZN(n4002) );
  AOI22_X1 U4561 ( .A1(n3628), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4562 ( .A1(n4552), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3639), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U4563 ( .A1(n5259), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3656), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U4564 ( .A1(n5261), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4004), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4005) );
  NAND4_X1 U4565 ( .A1(n4008), .A2(n4007), .A3(n4006), .A4(n4005), .ZN(n4017)
         );
  AOI22_X1 U4566 ( .A1(n3627), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4689), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U4567 ( .A1(n5266), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3643), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4014) );
  AOI22_X1 U4568 ( .A1(n3648), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U4569 ( .A1(n3623), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4488), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4012) );
  NAND4_X1 U4570 ( .A1(n4015), .A2(n4014), .A3(n4013), .A4(n4012), .ZN(n4016)
         );
  NAND2_X1 U4571 ( .A1(n4242), .A2(n4071), .ZN(n4051) );
  NAND2_X1 U4572 ( .A1(n4061), .A2(n4051), .ZN(n4050) );
  XNOR2_X2 U4573 ( .A(n4019), .B(n4018), .ZN(n4278) );
  AOI22_X1 U4574 ( .A1(n5259), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3622), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U4575 ( .A1(n3651), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U4576 ( .A1(n3650), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U4577 ( .A1(n5258), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4021) );
  NAND4_X1 U4578 ( .A1(n4024), .A2(n4023), .A3(n4022), .A4(n4021), .ZN(n4031)
         );
  AOI22_X1 U4579 ( .A1(n3653), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4689), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U4580 ( .A1(n3643), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U4581 ( .A1(n4488), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3657), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U4582 ( .A1(n5261), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4026) );
  NAND4_X1 U4583 ( .A1(n4029), .A2(n4028), .A3(n4027), .A4(n4026), .ZN(n4030)
         );
  INV_X1 U4584 ( .A(n4247), .ZN(n4043) );
  AOI22_X1 U4585 ( .A1(n4351), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4036) );
  AOI22_X1 U4586 ( .A1(n3628), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3659), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4035) );
  AOI22_X1 U4587 ( .A1(n3650), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4034) );
  AOI22_X1 U4588 ( .A1(n3622), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4488), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4033) );
  NAND4_X1 U4589 ( .A1(n4036), .A2(n4035), .A3(n4034), .A4(n4033), .ZN(n4042)
         );
  AOI22_X1 U4590 ( .A1(n3627), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3644), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U4591 ( .A1(n5259), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3655), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U4592 ( .A1(n5261), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4038) );
  AOI22_X1 U4593 ( .A1(n5258), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4037) );
  NAND4_X1 U4594 ( .A1(n4040), .A2(n4039), .A3(n4038), .A4(n4037), .ZN(n4041)
         );
  XNOR2_X1 U4595 ( .A(n4043), .B(n4083), .ZN(n4044) );
  NAND2_X1 U4596 ( .A1(n4055), .A2(n4081), .ZN(n4080) );
  INV_X1 U4597 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4048) );
  AOI21_X1 U4598 ( .B1(n5452), .B2(n4247), .A(n7437), .ZN(n4047) );
  NAND2_X1 U4599 ( .A1(n5563), .A2(n4083), .ZN(n4046) );
  NAND2_X1 U4600 ( .A1(n4242), .A2(n4247), .ZN(n4052) );
  NAND2_X1 U4601 ( .A1(n4050), .A2(n4049), .ZN(n4062) );
  INV_X1 U4602 ( .A(n4051), .ZN(n4053) );
  NOR2_X1 U4603 ( .A1(n4053), .A2(n3626), .ZN(n4056) );
  AND2_X1 U4604 ( .A1(n4081), .A2(n4056), .ZN(n4054) );
  NAND2_X1 U4605 ( .A1(n4055), .A2(n4054), .ZN(n4059) );
  INV_X1 U4606 ( .A(n4056), .ZN(n4057) );
  OR2_X1 U4607 ( .A1(n4057), .A2(n4079), .ZN(n4058) );
  NAND2_X1 U4608 ( .A1(n4059), .A2(n4058), .ZN(n4060) );
  INV_X1 U4609 ( .A(n4071), .ZN(n4065) );
  OAI22_X1 U4610 ( .A1(n4065), .A2(n4064), .B1(n4063), .B2(n4247), .ZN(n4066)
         );
  INV_X1 U4611 ( .A(n4066), .ZN(n4069) );
  INV_X1 U4612 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4067) );
  OR2_X1 U4613 ( .A1(n3836), .A2(n4067), .ZN(n4068) );
  NAND2_X1 U4614 ( .A1(n3646), .A2(n4243), .ZN(n4078) );
  NAND2_X1 U4615 ( .A1(n4083), .A2(n4071), .ZN(n4118) );
  OAI21_X1 U4616 ( .B1(n4083), .B2(n4071), .A(n4118), .ZN(n4072) );
  INV_X1 U4617 ( .A(n4072), .ZN(n4076) );
  NAND3_X1 U4618 ( .A1(n3638), .A2(n4074), .A3(n3994), .ZN(n4075) );
  AOI21_X1 U4619 ( .B1(n4076), .B2(n3958), .A(n4075), .ZN(n4077) );
  NAND2_X1 U4620 ( .A1(n5393), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4087)
         );
  MUX2_X2 U4621 ( .A(n4081), .B(n4080), .S(n4079), .Z(n6255) );
  NAND2_X1 U4622 ( .A1(n5563), .A2(n3994), .ZN(n4121) );
  OAI21_X1 U4623 ( .B1(n7443), .B2(n4083), .A(n4121), .ZN(n4084) );
  INV_X1 U4624 ( .A(n4084), .ZN(n4085) );
  NAND2_X1 U4625 ( .A1(n5347), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5394)
         );
  NAND2_X1 U4626 ( .A1(n4087), .A2(n5394), .ZN(n4090) );
  INV_X1 U4627 ( .A(n5393), .ZN(n4088) );
  NAND2_X1 U4628 ( .A1(n4088), .A2(n6653), .ZN(n4089) );
  NAND2_X1 U4629 ( .A1(n4090), .A2(n4089), .ZN(n7375) );
  INV_X1 U4630 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n7475) );
  INV_X1 U4631 ( .A(n4093), .ZN(n4095) );
  NAND2_X1 U4632 ( .A1(n4095), .A2(n4094), .ZN(n4097) );
  NAND2_X1 U4633 ( .A1(n4097), .A2(n3634), .ZN(n4129) );
  NAND2_X1 U4634 ( .A1(n4098), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4103) );
  INV_X1 U4635 ( .A(n4100), .ZN(n5911) );
  NAND2_X1 U4636 ( .A1(n5911), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5629) );
  INV_X1 U4637 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4099) );
  NAND2_X1 U4638 ( .A1(n4100), .A2(n4099), .ZN(n4101) );
  AND2_X1 U4639 ( .A1(n5629), .A2(n4101), .ZN(n5664) );
  INV_X1 U4640 ( .A(n4708), .ZN(n4133) );
  AOI22_X1 U4641 ( .A1(n5664), .A2(n4133), .B1(n4132), .B2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4102) );
  NAND2_X1 U4642 ( .A1(n4103), .A2(n4102), .ZN(n4127) );
  XNOR2_X1 U4643 ( .A(n4129), .B(n4127), .ZN(n5437) );
  NAND2_X1 U4644 ( .A1(n5437), .A2(n7437), .ZN(n4116) );
  AOI22_X1 U4645 ( .A1(n4689), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U4646 ( .A1(n3652), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3643), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U4647 ( .A1(n4552), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4106) );
  AOI22_X1 U4648 ( .A1(n3657), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4105) );
  NAND4_X1 U4649 ( .A1(n4108), .A2(n4107), .A3(n4106), .A4(n4105), .ZN(n4114)
         );
  AOI22_X1 U4650 ( .A1(n5259), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3648), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4112) );
  AOI22_X1 U4651 ( .A1(n3654), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4111) );
  INV_X1 U4652 ( .A(n4011), .ZN(n4505) );
  AOI22_X1 U4653 ( .A1(n3623), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4505), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4110) );
  AOI22_X1 U4654 ( .A1(n5261), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4109) );
  NAND4_X1 U4655 ( .A1(n4112), .A2(n4111), .A3(n4110), .A4(n4109), .ZN(n4113)
         );
  AOI22_X1 U4656 ( .A1(n4146), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4229), 
        .B2(n4117), .ZN(n4115) );
  INV_X1 U4657 ( .A(n4117), .ZN(n4119) );
  NAND2_X1 U4658 ( .A1(n4118), .A2(n4119), .ZN(n4150) );
  OAI21_X1 U4659 ( .B1(n4119), .B2(n4118), .A(n4150), .ZN(n4120) );
  NAND2_X1 U4660 ( .A1(n4120), .A2(n3958), .ZN(n4122) );
  NAND2_X1 U4661 ( .A1(n4122), .A2(n4121), .ZN(n4123) );
  NAND2_X1 U4662 ( .A1(n7375), .A2(n7475), .ZN(n4124) );
  NAND2_X1 U4663 ( .A1(n4125), .A2(n4124), .ZN(n5357) );
  INV_X1 U4664 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n5581) );
  INV_X1 U4665 ( .A(n4127), .ZN(n4128) );
  OR2_X2 U4666 ( .A1(n4129), .A2(n4128), .ZN(n5801) );
  NAND2_X1 U4667 ( .A1(n4098), .A2(n7181), .ZN(n4135) );
  INV_X1 U4668 ( .A(n5629), .ZN(n4130) );
  NAND2_X1 U4669 ( .A1(n4130), .A2(n7198), .ZN(n5439) );
  NAND2_X1 U4670 ( .A1(n5629), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4131) );
  NAND2_X1 U4671 ( .A1(n5439), .A2(n4131), .ZN(n5861) );
  AOI22_X1 U4672 ( .A1(n5861), .A2(n4133), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n4132), .ZN(n4134) );
  AOI22_X1 U4673 ( .A1(n3652), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4139) );
  AOI22_X1 U4674 ( .A1(n3644), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4138) );
  AOI22_X1 U4675 ( .A1(n3650), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4137) );
  AOI22_X1 U4676 ( .A1(n5261), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4136) );
  NAND4_X1 U4677 ( .A1(n4139), .A2(n4138), .A3(n4137), .A4(n4136), .ZN(n4145)
         );
  AOI22_X1 U4678 ( .A1(n3653), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4689), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4143) );
  AOI22_X1 U4679 ( .A1(n5259), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3656), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4142) );
  AOI22_X1 U4680 ( .A1(n3623), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4505), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4141) );
  AOI22_X1 U4681 ( .A1(n5258), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4140) );
  NAND4_X1 U4682 ( .A1(n4143), .A2(n4142), .A3(n4141), .A4(n4140), .ZN(n4144)
         );
  AOI22_X1 U4683 ( .A1(n4146), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4229), 
        .B2(n4151), .ZN(n4147) );
  NAND2_X1 U4684 ( .A1(n4150), .A2(n4151), .ZN(n4198) );
  OAI211_X1 U4685 ( .C1(n4151), .C2(n4150), .A(n4198), .B(n3958), .ZN(n4152)
         );
  INV_X1 U4686 ( .A(n4152), .ZN(n4153) );
  AOI21_X1 U4687 ( .B1(n3640), .B2(n4243), .A(n4153), .ZN(n5358) );
  OAI21_X1 U4688 ( .B1(n5357), .B2(n5581), .A(n5358), .ZN(n4155) );
  NAND2_X1 U4689 ( .A1(n5357), .A2(n5581), .ZN(n4154) );
  NAND2_X1 U4690 ( .A1(n4155), .A2(n4154), .ZN(n7382) );
  INV_X1 U4691 ( .A(n7382), .ZN(n4177) );
  INV_X1 U4692 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4160) );
  OR2_X1 U4693 ( .A1(n3836), .A2(n4160), .ZN(n4172) );
  AOI22_X1 U4694 ( .A1(n3653), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4164) );
  AOI22_X1 U4695 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n3659), .B1(n3651), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4163) );
  AOI22_X1 U4696 ( .A1(n4351), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3657), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4162) );
  AOI22_X1 U4697 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n5261), .B1(n5260), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4161) );
  NAND4_X1 U4698 ( .A1(n4164), .A2(n4163), .A3(n4162), .A4(n4161), .ZN(n4170)
         );
  AOI22_X1 U4699 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n5259), .B1(n4010), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4168) );
  AOI22_X1 U4700 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n4552), .B1(n3661), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4167) );
  AOI22_X1 U4701 ( .A1(n3648), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4166) );
  AOI22_X1 U4702 ( .A1(n4352), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4505), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4165) );
  NAND4_X1 U4703 ( .A1(n4168), .A2(n4167), .A3(n4166), .A4(n4165), .ZN(n4169)
         );
  NAND2_X1 U4704 ( .A1(n4229), .A2(n4196), .ZN(n4171) );
  NAND2_X1 U4705 ( .A1(n4309), .A2(n4243), .ZN(n4175) );
  XNOR2_X1 U4706 ( .A(n4198), .B(n4196), .ZN(n4173) );
  NAND2_X1 U4707 ( .A1(n4173), .A2(n3958), .ZN(n4174) );
  NAND2_X1 U4708 ( .A1(n4175), .A2(n4174), .ZN(n4178) );
  XNOR2_X1 U4709 ( .A(n4178), .B(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n7383)
         );
  INV_X1 U4710 ( .A(n7383), .ZN(n4176) );
  NAND2_X1 U4711 ( .A1(n4177), .A2(n4176), .ZN(n7385) );
  NAND2_X1 U4712 ( .A1(n4178), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4179)
         );
  NAND2_X1 U4713 ( .A1(n7385), .A2(n4179), .ZN(n5578) );
  INV_X1 U4714 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4183) );
  OR2_X1 U4715 ( .A1(n3836), .A2(n4183), .ZN(n4195) );
  AOI22_X1 U4716 ( .A1(n3628), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4187) );
  AOI22_X1 U4717 ( .A1(n3643), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3659), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4186) );
  AOI22_X1 U4718 ( .A1(n3650), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4185) );
  AOI22_X1 U4719 ( .A1(n5261), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4184) );
  NAND4_X1 U4720 ( .A1(n4187), .A2(n4186), .A3(n4185), .A4(n4184), .ZN(n4193)
         );
  AOI22_X1 U4721 ( .A1(n3627), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4689), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4191) );
  AOI22_X1 U4722 ( .A1(n5259), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3656), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4190) );
  AOI22_X1 U4723 ( .A1(n4010), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4505), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4189) );
  AOI22_X1 U4724 ( .A1(n5258), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4188) );
  NAND4_X1 U4725 ( .A1(n4191), .A2(n4190), .A3(n4189), .A4(n4188), .ZN(n4192)
         );
  NAND2_X1 U4726 ( .A1(n4229), .A2(n4224), .ZN(n4194) );
  NAND2_X1 U4727 ( .A1(n4195), .A2(n4194), .ZN(n4204) );
  NAND2_X1 U4728 ( .A1(n4310), .A2(n4243), .ZN(n4201) );
  INV_X1 U4729 ( .A(n4196), .ZN(n4197) );
  OR2_X1 U4730 ( .A1(n4198), .A2(n4197), .ZN(n4223) );
  XNOR2_X1 U4731 ( .A(n4223), .B(n4224), .ZN(n4199) );
  NAND2_X1 U4732 ( .A1(n4199), .A2(n3958), .ZN(n4200) );
  NAND2_X1 U4733 ( .A1(n4201), .A2(n4200), .ZN(n4202) );
  INV_X1 U4734 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n7460) );
  XNOR2_X1 U4735 ( .A(n4202), .B(n7460), .ZN(n5580) );
  NAND2_X1 U4736 ( .A1(n5578), .A2(n5580), .ZN(n5579) );
  NAND2_X1 U4737 ( .A1(n4202), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4203)
         );
  INV_X1 U4738 ( .A(n4204), .ZN(n4219) );
  INV_X1 U4739 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4205) );
  OR2_X1 U4740 ( .A1(n3836), .A2(n4205), .ZN(n4217) );
  AOI22_X1 U4741 ( .A1(n5259), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3648), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4209) );
  AOI22_X1 U4742 ( .A1(n3653), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4208) );
  AOI22_X1 U4743 ( .A1(n4552), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3651), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4207) );
  AOI22_X1 U4744 ( .A1(n4010), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3656), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4206) );
  NAND4_X1 U4745 ( .A1(n4209), .A2(n4208), .A3(n4207), .A4(n4206), .ZN(n4215)
         );
  AOI22_X1 U4746 ( .A1(n4351), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4213) );
  AOI22_X1 U4747 ( .A1(n5261), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4212) );
  AOI22_X1 U4748 ( .A1(n4505), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4211) );
  AOI22_X1 U4749 ( .A1(n3644), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4210) );
  NAND4_X1 U4750 ( .A1(n4213), .A2(n4212), .A3(n4211), .A4(n4210), .ZN(n4214)
         );
  NAND2_X1 U4751 ( .A1(n4229), .A2(n4234), .ZN(n4216) );
  OR2_X1 U4752 ( .A1(n4220), .A2(n4219), .ZN(n4222) );
  NAND2_X1 U4753 ( .A1(n4222), .A2(n4221), .ZN(n4322) );
  NAND3_X1 U4754 ( .A1(n4245), .A2(n4243), .A3(n4322), .ZN(n4228) );
  INV_X1 U4755 ( .A(n4223), .ZN(n4225) );
  NAND2_X1 U4756 ( .A1(n4225), .A2(n4224), .ZN(n4233) );
  XNOR2_X1 U4757 ( .A(n4233), .B(n4234), .ZN(n4226) );
  NAND2_X1 U4758 ( .A1(n4226), .A2(n3958), .ZN(n4227) );
  NAND2_X1 U4759 ( .A1(n4228), .A2(n4227), .ZN(n7395) );
  INV_X1 U4760 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4231) );
  NAND2_X1 U4761 ( .A1(n4229), .A2(n4247), .ZN(n4230) );
  OAI21_X1 U4762 ( .B1(n3836), .B2(n4231), .A(n4230), .ZN(n4232) );
  NAND2_X1 U4763 ( .A1(n4331), .A2(n4243), .ZN(n4238) );
  INV_X1 U4764 ( .A(n4233), .ZN(n4235) );
  NAND2_X1 U4765 ( .A1(n4235), .A2(n4234), .ZN(n4246) );
  XNOR2_X1 U4766 ( .A(n4246), .B(n4247), .ZN(n4236) );
  NAND2_X1 U4767 ( .A1(n4236), .A2(n3958), .ZN(n4237) );
  NAND2_X1 U4768 ( .A1(n4238), .A2(n4237), .ZN(n4239) );
  INV_X1 U4769 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n5149) );
  XNOR2_X1 U4770 ( .A(n4239), .B(n5149), .ZN(n6052) );
  NAND2_X1 U4771 ( .A1(n4239), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4240)
         );
  NAND2_X4 U4772 ( .A1(n4245), .A2(n4244), .ZN(n4252) );
  INV_X1 U4773 ( .A(n4246), .ZN(n4248) );
  NAND3_X1 U4774 ( .A1(n4248), .A2(n3958), .A3(n4247), .ZN(n4249) );
  NAND2_X1 U4775 ( .A1(n3641), .A2(n4249), .ZN(n4250) );
  NAND2_X1 U4776 ( .A1(n4250), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4251)
         );
  NAND2_X1 U4777 ( .A1(n4252), .A2(n7489), .ZN(n6463) );
  NAND2_X1 U4778 ( .A1(n6462), .A2(n6463), .ZN(n6501) );
  INV_X1 U4779 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n7503) );
  AND2_X1 U4780 ( .A1(n4252), .A2(n7503), .ZN(n6503) );
  INV_X1 U4781 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6506) );
  NAND2_X1 U4782 ( .A1(n3631), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6502) );
  NAND2_X1 U4783 ( .A1(n3631), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6505) );
  OAI211_X1 U4784 ( .C1(n4252), .C2(n6506), .A(n6502), .B(n6505), .ZN(n4253)
         );
  INV_X1 U4785 ( .A(n4253), .ZN(n4254) );
  NAND2_X1 U4786 ( .A1(n4252), .A2(n6506), .ZN(n4255) );
  INV_X1 U4787 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5168) );
  NAND2_X1 U4788 ( .A1(n4252), .A2(n5168), .ZN(n4257) );
  INV_X1 U4789 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6514) );
  NAND2_X1 U4790 ( .A1(n3631), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4258) );
  INV_X1 U4791 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n7514) );
  NAND2_X1 U4792 ( .A1(n4252), .A2(n7514), .ZN(n7041) );
  INV_X1 U4793 ( .A(n7036), .ZN(n4260) );
  INV_X1 U4794 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n7516) );
  NAND2_X1 U4795 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n7149) );
  NAND2_X1 U4796 ( .A1(n3631), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n7032) );
  OAI21_X1 U4797 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A(n3631), .ZN(n4261) );
  NOR2_X1 U4798 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n7122) );
  NOR2_X1 U4799 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n7150) );
  INV_X1 U4800 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6558) );
  INV_X1 U4801 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n7110) );
  AND4_X1 U4802 ( .A1(n7122), .A2(n7150), .A3(n6558), .A4(n7110), .ZN(n4263)
         );
  NOR2_X1 U4803 ( .A1(n4252), .A2(n4263), .ZN(n4265) );
  AND2_X1 U4804 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n7119) );
  AND2_X1 U4805 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n7121) );
  AND2_X1 U4806 ( .A1(n7119), .A2(n7121), .ZN(n7111) );
  AND2_X1 U4807 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6555) );
  NAND2_X1 U4808 ( .A1(n7111), .A2(n6555), .ZN(n6576) );
  NAND2_X1 U4809 ( .A1(n4252), .A2(n6576), .ZN(n4264) );
  XNOR2_X1 U4810 ( .A(n4252), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6976)
         );
  INV_X1 U4811 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n7103) );
  NAND2_X1 U4812 ( .A1(n4252), .A2(n7103), .ZN(n4266) );
  NAND2_X1 U4813 ( .A1(n6975), .A2(n4266), .ZN(n6966) );
  INV_X1 U4814 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n7091) );
  INV_X1 U4815 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5321) );
  OAI21_X1 U4816 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .A(n3631), .ZN(n4268) );
  INV_X1 U4817 ( .A(n4268), .ZN(n4269) );
  XNOR2_X1 U4818 ( .A(n4252), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4270)
         );
  NOR2_X1 U4819 ( .A1(n3937), .A2(n5838), .ZN(n4272) );
  NAND2_X1 U4820 ( .A1(n5433), .A2(n4457), .ZN(n4276) );
  AOI22_X1 U4821 ( .A1(n4283), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n5838), .ZN(n4274) );
  NAND2_X1 U4822 ( .A1(n4302), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4273) );
  AND2_X1 U4823 ( .A1(n4274), .A2(n4273), .ZN(n4275) );
  AND2_X1 U4824 ( .A1(n5446), .A2(n3933), .ZN(n4277) );
  INV_X1 U4825 ( .A(n4302), .ZN(n4298) );
  NAND2_X1 U4826 ( .A1(n4283), .A2(EAX_REG_0__SCAN_IN), .ZN(n4281) );
  NAND2_X1 U4827 ( .A1(n5838), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4280)
         );
  OAI211_X1 U4828 ( .C1(n4298), .C2(n4279), .A(n4281), .B(n4280), .ZN(n4282)
         );
  AOI21_X1 U4829 ( .B1(n4278), .B2(n4457), .A(n4282), .ZN(n5345) );
  NAND2_X1 U4830 ( .A1(n5355), .A2(n5354), .ZN(n5353) );
  NAND2_X1 U4831 ( .A1(n4302), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4288) );
  NAND2_X1 U4832 ( .A1(n5838), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4626) );
  INV_X1 U4833 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4285) );
  OAI21_X1 U4834 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n4293), .ZN(n7381) );
  NAND2_X1 U4835 ( .A1(n5282), .A2(n7381), .ZN(n4284) );
  OAI21_X1 U4836 ( .B1(n4626), .B2(n4285), .A(n4284), .ZN(n4286) );
  AOI21_X1 U4837 ( .B1(n6660), .B2(EAX_REG_2__SCAN_IN), .A(n4286), .ZN(n4287)
         );
  AND2_X1 U4838 ( .A1(n4288), .A2(n4287), .ZN(n4290) );
  NOR2_X1 U4839 ( .A1(n5353), .A2(n4290), .ZN(n4291) );
  NAND2_X1 U4840 ( .A1(n5432), .A2(n4457), .ZN(n4289) );
  NAND2_X1 U4841 ( .A1(n5353), .A2(n4290), .ZN(n5531) );
  OAI21_X1 U4842 ( .B1(n4291), .B2(n5530), .A(n5531), .ZN(n4292) );
  NAND2_X1 U4843 ( .A1(n5502), .A2(n4457), .ZN(n4301) );
  INV_X1 U4844 ( .A(n4293), .ZN(n4295) );
  INV_X1 U4845 ( .A(n4304), .ZN(n4294) );
  OAI21_X1 U4846 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n4295), .A(n4294), 
        .ZN(n6857) );
  AOI22_X1 U4847 ( .A1(n5282), .A2(n6857), .B1(n6659), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4297) );
  NAND2_X1 U4848 ( .A1(n6660), .A2(EAX_REG_3__SCAN_IN), .ZN(n4296) );
  OAI211_X1 U4849 ( .C1(n4298), .C2(n3751), .A(n4297), .B(n4296), .ZN(n4299)
         );
  INV_X1 U4850 ( .A(n4299), .ZN(n4300) );
  NAND2_X1 U4851 ( .A1(n4302), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4307) );
  INV_X1 U4852 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6302) );
  AOI21_X1 U4853 ( .B1(n6302), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4303) );
  AOI21_X1 U4854 ( .B1(n6660), .B2(EAX_REG_4__SCAN_IN), .A(n4303), .ZN(n4306)
         );
  NAND2_X1 U4855 ( .A1(n4304), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4311)
         );
  OAI21_X1 U4856 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n4304), .A(n4311), 
        .ZN(n7389) );
  NOR2_X1 U4857 ( .A1(n4665), .A2(n7389), .ZN(n4305) );
  AOI21_X1 U4858 ( .B1(n4307), .B2(n4306), .A(n4305), .ZN(n4308) );
  AOI21_X1 U4859 ( .B1(n4309), .B2(n4457), .A(n4308), .ZN(n5496) );
  NAND2_X1 U4860 ( .A1(n4310), .A2(n4457), .ZN(n4317) );
  INV_X1 U4861 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4314) );
  OAI21_X1 U4862 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n4312), .A(n4318), 
        .ZN(n7567) );
  NAND2_X1 U4863 ( .A1(n7567), .A2(n5282), .ZN(n4313) );
  OAI21_X1 U4864 ( .B1(n4314), .B2(n4626), .A(n4313), .ZN(n4315) );
  AOI21_X1 U4865 ( .B1(n6660), .B2(EAX_REG_5__SCAN_IN), .A(n4315), .ZN(n4316)
         );
  NAND2_X1 U4866 ( .A1(n4317), .A2(n4316), .ZN(n5488) );
  NAND2_X1 U4867 ( .A1(n5487), .A2(n5488), .ZN(n5485) );
  INV_X1 U4868 ( .A(n5485), .ZN(n4324) );
  INV_X1 U4869 ( .A(EAX_REG_6__SCAN_IN), .ZN(n7269) );
  OAI21_X1 U4870 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n4319), .A(n4325), 
        .ZN(n7584) );
  AOI22_X1 U4871 ( .A1(n5282), .A2(n7584), .B1(n6659), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4320) );
  OAI21_X1 U4872 ( .B1(n4548), .B2(n7269), .A(n4320), .ZN(n4321) );
  NAND2_X1 U4873 ( .A1(n4324), .A2(n4323), .ZN(n5522) );
  INV_X1 U4874 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4329) );
  INV_X1 U4875 ( .A(n4325), .ZN(n4327) );
  INV_X1 U4876 ( .A(n4346), .ZN(n4326) );
  OAI21_X1 U4877 ( .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n4327), .A(n4326), 
        .ZN(n7596) );
  AOI22_X1 U4878 ( .A1(n5282), .A2(n7596), .B1(n6659), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4328) );
  OAI21_X1 U4879 ( .B1(n4548), .B2(n4329), .A(n4328), .ZN(n4330) );
  AOI22_X1 U4880 ( .A1(n4010), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n5258), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4336) );
  AOI22_X1 U4881 ( .A1(n3652), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4335) );
  AOI22_X1 U4882 ( .A1(n4552), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4334) );
  AOI22_X1 U4883 ( .A1(n4351), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4505), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4333) );
  NAND4_X1 U4884 ( .A1(n4336), .A2(n4335), .A3(n4334), .A4(n4333), .ZN(n4342)
         );
  AOI22_X1 U4885 ( .A1(n3643), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4340) );
  AOI22_X1 U4886 ( .A1(n3654), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3656), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4339) );
  AOI22_X1 U4887 ( .A1(n5261), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4338) );
  AOI22_X1 U4888 ( .A1(n5259), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4337) );
  NAND4_X1 U4889 ( .A1(n4340), .A2(n4339), .A3(n4338), .A4(n4337), .ZN(n4341)
         );
  OAI21_X1 U4890 ( .B1(n4342), .B2(n4341), .A(n4457), .ZN(n4345) );
  XNOR2_X1 U4891 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n4346), .ZN(n7604) );
  AOI22_X1 U4892 ( .A1(n5282), .A2(n7604), .B1(n6659), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4344) );
  NAND2_X1 U4893 ( .A1(n6660), .A2(EAX_REG_8__SCAN_IN), .ZN(n4343) );
  XOR2_X1 U4894 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n4362), .Z(n7616) );
  AOI22_X1 U4895 ( .A1(n5259), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3648), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4350) );
  AOI22_X1 U4896 ( .A1(n3627), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3659), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4349) );
  AOI22_X1 U4897 ( .A1(n3650), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5261), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4348) );
  AOI22_X1 U4898 ( .A1(n4505), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3655), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4347) );
  NAND4_X1 U4899 ( .A1(n4350), .A2(n4349), .A3(n4348), .A4(n4347), .ZN(n4358)
         );
  AOI22_X1 U4900 ( .A1(n4351), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4356) );
  AOI22_X1 U4901 ( .A1(n3628), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4352), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4355) );
  AOI22_X1 U4902 ( .A1(n4010), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4354) );
  AOI22_X1 U4903 ( .A1(n3661), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4353) );
  NAND4_X1 U4904 ( .A1(n4356), .A2(n4355), .A3(n4354), .A4(n4353), .ZN(n4357)
         );
  OR2_X1 U4905 ( .A1(n4358), .A2(n4357), .ZN(n4359) );
  AOI22_X1 U4906 ( .A1(n4457), .A2(n4359), .B1(n6659), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4361) );
  NAND2_X1 U4907 ( .A1(n6660), .A2(EAX_REG_9__SCAN_IN), .ZN(n4360) );
  OAI211_X1 U4908 ( .C1(n7616), .C2(n4665), .A(n4361), .B(n4360), .ZN(n6230)
         );
  XNOR2_X1 U4909 ( .A(n4379), .B(n7623), .ZN(n7624) );
  NAND2_X1 U4910 ( .A1(n7624), .A2(n5282), .ZN(n4377) );
  AOI22_X1 U4911 ( .A1(n3653), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4689), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4366) );
  AOI22_X1 U4912 ( .A1(n3651), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4365) );
  AOI22_X1 U4913 ( .A1(n4010), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4505), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4364) );
  AOI22_X1 U4914 ( .A1(n3643), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4363) );
  NAND4_X1 U4915 ( .A1(n4366), .A2(n4365), .A3(n4364), .A4(n4363), .ZN(n4372)
         );
  AOI22_X1 U4916 ( .A1(n5266), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5261), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4370) );
  AOI22_X1 U4917 ( .A1(n4552), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4369) );
  AOI22_X1 U4918 ( .A1(n5258), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4368) );
  AOI22_X1 U4919 ( .A1(n5259), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3657), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4367) );
  NAND4_X1 U4920 ( .A1(n4370), .A2(n4369), .A3(n4368), .A4(n4367), .ZN(n4371)
         );
  OAI21_X1 U4921 ( .B1(n4372), .B2(n4371), .A(n4457), .ZN(n4375) );
  NAND2_X1 U4922 ( .A1(n6660), .A2(EAX_REG_10__SCAN_IN), .ZN(n4374) );
  NAND2_X1 U4923 ( .A1(n6659), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4373)
         );
  AND3_X1 U4924 ( .A1(n4375), .A2(n4374), .A3(n4373), .ZN(n4376) );
  NAND2_X1 U4925 ( .A1(n4377), .A2(n4376), .ZN(n6262) );
  XOR2_X1 U4926 ( .A(n7632), .B(n4393), .Z(n7638) );
  AOI22_X1 U4927 ( .A1(n5259), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4689), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4383) );
  AOI22_X1 U4928 ( .A1(n3651), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4382) );
  AOI22_X1 U4929 ( .A1(n5261), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4381) );
  AOI22_X1 U4930 ( .A1(n3644), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4380) );
  NAND4_X1 U4931 ( .A1(n4383), .A2(n4382), .A3(n4381), .A4(n4380), .ZN(n4389)
         );
  AOI22_X1 U4932 ( .A1(n4552), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4387) );
  AOI22_X1 U4933 ( .A1(n4010), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3657), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4386) );
  AOI22_X1 U4934 ( .A1(n3653), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4505), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4385) );
  AOI22_X1 U4935 ( .A1(n3648), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4384) );
  NAND4_X1 U4936 ( .A1(n4387), .A2(n4386), .A3(n4385), .A4(n4384), .ZN(n4388)
         );
  OR2_X1 U4937 ( .A1(n4389), .A2(n4388), .ZN(n4390) );
  AOI22_X1 U4938 ( .A1(n4457), .A2(n4390), .B1(n6659), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4392) );
  NAND2_X1 U4939 ( .A1(n6660), .A2(EAX_REG_11__SCAN_IN), .ZN(n4391) );
  OAI211_X1 U4940 ( .C1(n7638), .C2(n4665), .A(n4392), .B(n4391), .ZN(n6291)
         );
  NAND2_X1 U4941 ( .A1(n6261), .A2(n6291), .ZN(n6289) );
  XNOR2_X1 U4942 ( .A(n4429), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6850)
         );
  NAND2_X1 U4943 ( .A1(n6850), .A2(n5282), .ZN(n4412) );
  INV_X1 U4944 ( .A(EAX_REG_12__SCAN_IN), .ZN(n4396) );
  AOI21_X1 U4945 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n6848), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4394) );
  INV_X1 U4946 ( .A(n4394), .ZN(n4395) );
  OAI21_X1 U4947 ( .B1(n4548), .B2(n4396), .A(n4395), .ZN(n4411) );
  INV_X1 U4948 ( .A(n4457), .ZN(n4409) );
  AOI22_X1 U4949 ( .A1(n5259), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4689), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4401) );
  AOI22_X1 U4950 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n3660), .B1(n3652), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4400) );
  AOI22_X1 U4951 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n3643), .B1(n3661), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4399) );
  AOI22_X1 U4952 ( .A1(n3647), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4398) );
  NAND4_X1 U4953 ( .A1(n4401), .A2(n4400), .A3(n4399), .A4(n4398), .ZN(n4407)
         );
  AOI22_X1 U4954 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3650), .B1(n5261), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4405) );
  AOI22_X1 U4955 ( .A1(n4010), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3655), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4404) );
  AOI22_X1 U4956 ( .A1(n3653), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4505), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4403) );
  AOI22_X1 U4957 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n5266), .B1(n5260), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4402) );
  NAND4_X1 U4958 ( .A1(n4405), .A2(n4404), .A3(n4403), .A4(n4402), .ZN(n4406)
         );
  NOR2_X1 U4959 ( .A1(n4407), .A2(n4406), .ZN(n4408) );
  NOR2_X1 U4960 ( .A1(n4409), .A2(n4408), .ZN(n4410) );
  AOI21_X1 U4961 ( .B1(n4412), .B2(n4411), .A(n4410), .ZN(n6449) );
  INV_X1 U4962 ( .A(n6449), .ZN(n4425) );
  AOI22_X1 U4963 ( .A1(n3653), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4689), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4416) );
  AOI22_X1 U4964 ( .A1(n3652), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4415) );
  AOI22_X1 U4965 ( .A1(n4552), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5261), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4414) );
  AOI22_X1 U4966 ( .A1(n3657), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4413) );
  NAND4_X1 U4967 ( .A1(n4416), .A2(n4415), .A3(n4414), .A4(n4413), .ZN(n4422)
         );
  AOI22_X1 U4968 ( .A1(n5259), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5258), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4420) );
  AOI22_X1 U4969 ( .A1(n5266), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3643), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4419) );
  AOI22_X1 U4970 ( .A1(n4010), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4505), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4418) );
  AOI22_X1 U4971 ( .A1(n3661), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4417) );
  NAND4_X1 U4972 ( .A1(n4420), .A2(n4419), .A3(n4418), .A4(n4417), .ZN(n4421)
         );
  OR2_X1 U4973 ( .A1(n4422), .A2(n4421), .ZN(n4423) );
  NAND2_X1 U4974 ( .A1(n4457), .A2(n4423), .ZN(n4427) );
  INV_X1 U4975 ( .A(n4427), .ZN(n4424) );
  NAND2_X1 U4976 ( .A1(n4425), .A2(n4424), .ZN(n4426) );
  OR2_X2 U4977 ( .A1(n6289), .A2(n4426), .ZN(n4433) );
  NAND2_X1 U4978 ( .A1(n6660), .A2(EAX_REG_13__SCAN_IN), .ZN(n4432) );
  OAI21_X1 U4979 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n4430), .A(n4434), 
        .ZN(n7661) );
  AOI22_X1 U4980 ( .A1(n5282), .A2(n7661), .B1(n6659), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4431) );
  NAND2_X1 U4981 ( .A1(n4432), .A2(n4431), .ZN(n6492) );
  NAND2_X1 U4982 ( .A1(n6491), .A2(n6492), .ZN(n6495) );
  NAND2_X2 U4983 ( .A1(n6495), .A2(n4433), .ZN(n6833) );
  XOR2_X1 U4984 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n4448), .Z(n7056) );
  AOI22_X1 U4985 ( .A1(n3653), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3644), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4438) );
  AOI22_X1 U4986 ( .A1(n5261), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4437) );
  AOI22_X1 U4987 ( .A1(n5259), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3656), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4436) );
  AOI22_X1 U4988 ( .A1(n4689), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4505), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4435) );
  NAND4_X1 U4989 ( .A1(n4438), .A2(n4437), .A3(n4436), .A4(n4435), .ZN(n4444)
         );
  AOI22_X1 U4990 ( .A1(n4010), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4442) );
  AOI22_X1 U4991 ( .A1(n3652), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3659), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4441) );
  AOI22_X1 U4992 ( .A1(n5258), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4440) );
  AOI22_X1 U4993 ( .A1(n3650), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4439) );
  NAND4_X1 U4994 ( .A1(n4442), .A2(n4441), .A3(n4440), .A4(n4439), .ZN(n4443)
         );
  OR2_X1 U4995 ( .A1(n4444), .A2(n4443), .ZN(n4445) );
  AOI22_X1 U4996 ( .A1(n4457), .A2(n4445), .B1(n6659), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4447) );
  NAND2_X1 U4997 ( .A1(n6660), .A2(EAX_REG_14__SCAN_IN), .ZN(n4446) );
  OAI211_X1 U4998 ( .C1(n7056), .C2(n4665), .A(n4447), .B(n4446), .ZN(n6832)
         );
  XNOR2_X1 U4999 ( .A(n4465), .B(n6824), .ZN(n7045) );
  AOI22_X1 U5000 ( .A1(n3653), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4452) );
  AOI22_X1 U5001 ( .A1(n4552), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4451) );
  AOI22_X1 U5002 ( .A1(n4010), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3656), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4450) );
  AOI22_X1 U5003 ( .A1(n4689), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4505), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4449) );
  NAND4_X1 U5004 ( .A1(n4452), .A2(n4451), .A3(n4450), .A4(n4449), .ZN(n4459)
         );
  AOI22_X1 U5005 ( .A1(n5259), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3651), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4456) );
  AOI22_X1 U5006 ( .A1(n4352), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3659), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4455) );
  AOI22_X1 U5007 ( .A1(n3648), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4454) );
  AOI22_X1 U5008 ( .A1(n5261), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4453) );
  NAND4_X1 U5009 ( .A1(n4456), .A2(n4455), .A3(n4454), .A4(n4453), .ZN(n4458)
         );
  OAI21_X1 U5010 ( .B1(n4459), .B2(n4458), .A(n4457), .ZN(n4462) );
  NAND2_X1 U5011 ( .A1(n6660), .A2(EAX_REG_15__SCAN_IN), .ZN(n4461) );
  NAND2_X1 U5012 ( .A1(n6659), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4460)
         );
  NAND3_X1 U5013 ( .A1(n4462), .A2(n4461), .A3(n4460), .ZN(n4463) );
  AOI21_X1 U5014 ( .B1(n7045), .B2(n5282), .A(n4463), .ZN(n6822) );
  XOR2_X1 U5015 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n4481), .Z(n7038) );
  INV_X1 U5016 ( .A(n7038), .ZN(n4480) );
  AOI22_X1 U5017 ( .A1(n5259), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3627), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4470) );
  AOI22_X1 U5018 ( .A1(n5266), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3659), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4469) );
  AOI22_X1 U5019 ( .A1(n3648), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4468) );
  AOI22_X1 U5020 ( .A1(n3650), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4467) );
  NAND4_X1 U5021 ( .A1(n4470), .A2(n4469), .A3(n4468), .A4(n4467), .ZN(n4476)
         );
  AOI22_X1 U5022 ( .A1(n3628), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3644), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4474) );
  AOI22_X1 U5023 ( .A1(n5261), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4473) );
  AOI22_X1 U5024 ( .A1(n3623), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3657), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4472) );
  AOI22_X1 U5025 ( .A1(n4351), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4505), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4471) );
  NAND4_X1 U5026 ( .A1(n4474), .A2(n4473), .A3(n4472), .A4(n4471), .ZN(n4475)
         );
  NOR2_X1 U5027 ( .A1(n4476), .A2(n4475), .ZN(n4478) );
  AOI22_X1 U5028 ( .A1(n6660), .A2(EAX_REG_16__SCAN_IN), .B1(n6659), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4477) );
  OAI21_X1 U5029 ( .B1(n5278), .B2(n4478), .A(n4477), .ZN(n4479) );
  AOI21_X1 U5030 ( .B1(n4480), .B2(n5282), .A(n4479), .ZN(n6801) );
  XNOR2_X1 U5031 ( .A(n4499), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n7030)
         );
  NAND2_X1 U5032 ( .A1(n5278), .A2(n4665), .ZN(n4563) );
  AOI22_X1 U5033 ( .A1(n5259), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4487) );
  AOI22_X1 U5034 ( .A1(n3622), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3653), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4486) );
  NAND2_X1 U5035 ( .A1(n3661), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4483) );
  NAND2_X1 U5036 ( .A1(n5266), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4482)
         );
  AND3_X1 U5037 ( .A1(n4483), .A2(n4482), .A3(n4665), .ZN(n4485) );
  AOI22_X1 U5038 ( .A1(n3648), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3656), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4484) );
  NAND4_X1 U5039 ( .A1(n4487), .A2(n4486), .A3(n4485), .A4(n4484), .ZN(n4494)
         );
  AOI22_X1 U5040 ( .A1(n3649), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3643), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4492) );
  AOI22_X1 U5041 ( .A1(n3658), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4488), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4491) );
  AOI22_X1 U5042 ( .A1(n3651), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4490) );
  AOI22_X1 U5043 ( .A1(n5261), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4489) );
  NAND4_X1 U5044 ( .A1(n4492), .A2(n4491), .A3(n4490), .A4(n4489), .ZN(n4493)
         );
  OR2_X1 U5045 ( .A1(n4494), .A2(n4493), .ZN(n4497) );
  INV_X1 U5046 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4495) );
  OAI22_X1 U5047 ( .A1(n4548), .A2(n4495), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n7026), .ZN(n4496) );
  AOI21_X1 U5048 ( .B1(n4563), .B2(n4497), .A(n4496), .ZN(n4498) );
  AOI21_X1 U5049 ( .B1(n7030), .B2(n5282), .A(n4498), .ZN(n6789) );
  OAI21_X1 U5050 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n4500), .A(n4532), 
        .ZN(n7669) );
  AOI22_X1 U5051 ( .A1(n5259), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4689), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4504) );
  AOI22_X1 U5052 ( .A1(n5266), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4503) );
  AOI22_X1 U5053 ( .A1(n3650), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4502) );
  AOI22_X1 U5054 ( .A1(n5261), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4501) );
  NAND4_X1 U5055 ( .A1(n4504), .A2(n4503), .A3(n4502), .A4(n4501), .ZN(n4511)
         );
  AOI22_X1 U5056 ( .A1(n3651), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3644), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4509) );
  AOI22_X1 U5057 ( .A1(n4010), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3656), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4508) );
  AOI22_X1 U5058 ( .A1(n3653), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4505), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4507) );
  AOI22_X1 U5059 ( .A1(n5258), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4506) );
  NAND4_X1 U5060 ( .A1(n4509), .A2(n4508), .A3(n4507), .A4(n4506), .ZN(n4510)
         );
  NOR2_X1 U5061 ( .A1(n4511), .A2(n4510), .ZN(n4513) );
  AOI22_X1 U5062 ( .A1(n6660), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n5838), .ZN(n4512) );
  OAI21_X1 U5063 ( .B1(n5278), .B2(n4513), .A(n4512), .ZN(n4514) );
  MUX2_X1 U5064 ( .A(n7669), .B(n4514), .S(n4665), .Z(n6903) );
  AOI22_X1 U5065 ( .A1(n3648), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4351), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4521) );
  NAND2_X1 U5066 ( .A1(n3623), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4517) );
  NAND2_X1 U5067 ( .A1(n5261), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4516) );
  AND3_X1 U5068 ( .A1(n4517), .A2(n4516), .A3(n4665), .ZN(n4520) );
  AOI22_X1 U5069 ( .A1(n4352), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3657), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4519) );
  AOI22_X1 U5070 ( .A1(n3659), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4518) );
  NAND4_X1 U5071 ( .A1(n4521), .A2(n4520), .A3(n4519), .A4(n4518), .ZN(n4527)
         );
  AOI22_X1 U5072 ( .A1(n3650), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4525) );
  AOI22_X1 U5073 ( .A1(n5259), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4524) );
  AOI22_X1 U5074 ( .A1(n3627), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4523) );
  AOI22_X1 U5075 ( .A1(n3628), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4488), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4522) );
  NAND4_X1 U5076 ( .A1(n4525), .A2(n4524), .A3(n4523), .A4(n4522), .ZN(n4526)
         );
  OR2_X1 U5077 ( .A1(n4527), .A2(n4526), .ZN(n4528) );
  NAND2_X1 U5078 ( .A1(n4563), .A2(n4528), .ZN(n4531) );
  AOI22_X1 U5079 ( .A1(n6660), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n5838), .ZN(n4530) );
  XNOR2_X1 U5080 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n4532), .ZN(n7683)
         );
  AOI21_X1 U5081 ( .B1(n4531), .B2(n4530), .A(n4529), .ZN(n6902) );
  INV_X1 U5082 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n7011) );
  INV_X1 U5083 ( .A(n4534), .ZN(n4535) );
  NAND2_X1 U5084 ( .A1(n7011), .A2(n4535), .ZN(n4536) );
  NAND2_X1 U5085 ( .A1(n4570), .A2(n4536), .ZN(n7700) );
  INV_X1 U5086 ( .A(n7700), .ZN(n7013) );
  AOI22_X1 U5087 ( .A1(n5259), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3647), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4540) );
  AOI22_X1 U5088 ( .A1(n3654), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n5261), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4539) );
  AOI22_X1 U5089 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3649), .B1(n3661), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4538) );
  AOI22_X1 U5090 ( .A1(n4010), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4505), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4537) );
  NAND4_X1 U5091 ( .A1(n4540), .A2(n4539), .A3(n4538), .A4(n4537), .ZN(n4546)
         );
  AOI22_X1 U5092 ( .A1(n4351), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4544) );
  AOI22_X1 U5093 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n3660), .B1(n3628), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4543) );
  AOI22_X1 U5094 ( .A1(n3656), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4542) );
  AOI22_X1 U5095 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n4352), .B1(n5260), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4541) );
  NAND4_X1 U5096 ( .A1(n4544), .A2(n4543), .A3(n4542), .A4(n4541), .ZN(n4545)
         );
  OR2_X1 U5097 ( .A1(n4546), .A2(n4545), .ZN(n4550) );
  INV_X1 U5098 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4547) );
  OAI22_X1 U5099 ( .A1(n4548), .A2(n4547), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n7011), .ZN(n4549) );
  AOI21_X1 U5100 ( .B1(n5236), .B2(n4550), .A(n4549), .ZN(n4551) );
  MUX2_X1 U5101 ( .A(n7013), .B(n4551), .S(n4665), .Z(n7014) );
  AOI22_X1 U5102 ( .A1(n3653), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3649), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4556) );
  AOI22_X1 U5103 ( .A1(n5259), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4555) );
  AOI22_X1 U5104 ( .A1(n3921), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4554) );
  AOI22_X1 U5105 ( .A1(n5261), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4505), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4553) );
  NAND4_X1 U5106 ( .A1(n4556), .A2(n4555), .A3(n4554), .A4(n4553), .ZN(n4565)
         );
  AOI22_X1 U5107 ( .A1(n3648), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4562) );
  AOI22_X1 U5108 ( .A1(n4010), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4032), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4561) );
  AOI22_X1 U5109 ( .A1(n3651), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3644), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4560) );
  NAND2_X1 U5110 ( .A1(n5260), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4558)
         );
  NAND2_X1 U5111 ( .A1(n3656), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4557) );
  AND3_X1 U5112 ( .A1(n4558), .A2(n4557), .A3(n4665), .ZN(n4559) );
  NAND4_X1 U5113 ( .A1(n4562), .A2(n4561), .A3(n4560), .A4(n4559), .ZN(n4564)
         );
  OAI21_X1 U5114 ( .B1(n4565), .B2(n4564), .A(n4563), .ZN(n4567) );
  AOI22_X1 U5115 ( .A1(n6660), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n5838), .ZN(n4566) );
  NAND2_X1 U5116 ( .A1(n4567), .A2(n4566), .ZN(n4569) );
  XNOR2_X1 U5117 ( .A(n4570), .B(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n7003)
         );
  NAND2_X1 U5118 ( .A1(n7003), .A2(n5282), .ZN(n4568) );
  NAND2_X1 U5119 ( .A1(n4569), .A2(n4568), .ZN(n5110) );
  NOR2_X2 U5120 ( .A1(n5107), .A2(n5110), .ZN(n5108) );
  INV_X1 U5121 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n7001) );
  OR2_X1 U5122 ( .A1(n4571), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4572)
         );
  NAND2_X1 U5123 ( .A1(n4623), .A2(n4572), .ZN(n6993) );
  AOI22_X1 U5124 ( .A1(n4010), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4576) );
  AOI22_X1 U5125 ( .A1(n3651), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3643), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4575) );
  AOI22_X1 U5126 ( .A1(n3650), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4574) );
  AOI22_X1 U5127 ( .A1(n5259), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3657), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4573) );
  NAND4_X1 U5128 ( .A1(n4576), .A2(n4575), .A3(n4574), .A4(n4573), .ZN(n4582)
         );
  AOI22_X1 U5129 ( .A1(n3653), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3659), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4580) );
  AOI22_X1 U5130 ( .A1(n3921), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4488), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4579) );
  AOI22_X1 U5131 ( .A1(n5261), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4578) );
  AOI22_X1 U5132 ( .A1(n3647), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4577) );
  NAND4_X1 U5133 ( .A1(n4580), .A2(n4579), .A3(n4578), .A4(n4577), .ZN(n4581)
         );
  NOR2_X1 U5134 ( .A1(n4582), .A2(n4581), .ZN(n4584) );
  AOI22_X1 U5135 ( .A1(n6660), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n5838), .ZN(n4583) );
  OAI21_X1 U5136 ( .B1(n5278), .B2(n4584), .A(n4583), .ZN(n4585) );
  MUX2_X1 U5137 ( .A(n6993), .B(n4585), .S(n4665), .Z(n6770) );
  NAND2_X1 U5138 ( .A1(n5108), .A2(n6770), .ZN(n6759) );
  AOI22_X1 U5139 ( .A1(n5259), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3648), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4589) );
  AOI22_X1 U5140 ( .A1(n3628), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4588) );
  AOI22_X1 U5141 ( .A1(n3627), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3656), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4587) );
  AOI22_X1 U5142 ( .A1(n3661), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4586) );
  NAND4_X1 U5143 ( .A1(n4589), .A2(n4588), .A3(n4587), .A4(n4586), .ZN(n4595)
         );
  AOI22_X1 U5144 ( .A1(n5266), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4352), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4593) );
  AOI22_X1 U5145 ( .A1(n3650), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5261), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4592) );
  AOI22_X1 U5146 ( .A1(n4010), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4591) );
  AOI22_X1 U5147 ( .A1(n4689), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4505), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4590) );
  NAND4_X1 U5148 ( .A1(n4593), .A2(n4592), .A3(n4591), .A4(n4590), .ZN(n4594)
         );
  NOR2_X1 U5149 ( .A1(n4595), .A2(n4594), .ZN(n4611) );
  AOI22_X1 U5150 ( .A1(n4689), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4599) );
  AOI22_X1 U5151 ( .A1(n3650), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3659), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4598) );
  AOI22_X1 U5152 ( .A1(n3647), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4597) );
  AOI22_X1 U5153 ( .A1(n4010), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4505), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4596) );
  NAND4_X1 U5154 ( .A1(n4599), .A2(n4598), .A3(n4597), .A4(n4596), .ZN(n4605)
         );
  AOI22_X1 U5155 ( .A1(n3627), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3628), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4603) );
  AOI22_X1 U5156 ( .A1(n5261), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4602) );
  AOI22_X1 U5157 ( .A1(n5259), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3656), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4601) );
  AOI22_X1 U5158 ( .A1(n4352), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4600) );
  NAND4_X1 U5159 ( .A1(n4603), .A2(n4602), .A3(n4601), .A4(n4600), .ZN(n4604)
         );
  NOR2_X1 U5160 ( .A1(n4605), .A2(n4604), .ZN(n4612) );
  XOR2_X1 U5161 ( .A(n4611), .B(n4612), .Z(n4608) );
  INV_X1 U5162 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6985) );
  NAND2_X1 U5163 ( .A1(n6660), .A2(EAX_REG_23__SCAN_IN), .ZN(n4606) );
  OAI21_X1 U5164 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6985), .A(n4606), .ZN(
        n4607) );
  AOI21_X1 U5165 ( .B1(n5236), .B2(n4608), .A(n4607), .ZN(n4609) );
  XNOR2_X1 U5166 ( .A(n4623), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6987)
         );
  MUX2_X1 U5167 ( .A(n4609), .B(n6987), .S(n5282), .Z(n6760) );
  NAND2_X1 U5168 ( .A1(n6761), .A2(n4610), .ZN(n6561) );
  OR2_X1 U5169 ( .A1(n4612), .A2(n4611), .ZN(n4641) );
  AOI22_X1 U5170 ( .A1(n3652), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5261), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4616) );
  AOI22_X1 U5171 ( .A1(n5259), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4615) );
  AOI22_X1 U5172 ( .A1(n3649), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3659), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4614) );
  AOI22_X1 U5173 ( .A1(n4505), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4613) );
  NAND4_X1 U5174 ( .A1(n4616), .A2(n4615), .A3(n4614), .A4(n4613), .ZN(n4622)
         );
  AOI22_X1 U5175 ( .A1(n5258), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3644), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4620) );
  AOI22_X1 U5176 ( .A1(n3654), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4689), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4619) );
  AOI22_X1 U5177 ( .A1(n5266), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4618) );
  AOI22_X1 U5178 ( .A1(n4010), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3657), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4617) );
  NAND4_X1 U5179 ( .A1(n4620), .A2(n4619), .A3(n4618), .A4(n4617), .ZN(n4621)
         );
  OR2_X1 U5180 ( .A1(n4622), .A2(n4621), .ZN(n4639) );
  XNOR2_X1 U5181 ( .A(n4641), .B(n4639), .ZN(n4628) );
  INV_X1 U5182 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6750) );
  NAND2_X1 U5183 ( .A1(n6660), .A2(EAX_REG_24__SCAN_IN), .ZN(n4625) );
  XNOR2_X1 U5184 ( .A(n4644), .B(n6750), .ZN(n6749) );
  NAND2_X1 U5185 ( .A1(n6749), .A2(n5282), .ZN(n4624) );
  OAI211_X1 U5186 ( .C1(n4626), .C2(n6750), .A(n4625), .B(n4624), .ZN(n4627)
         );
  AOI21_X1 U5187 ( .B1(n5236), .B2(n4628), .A(n4627), .ZN(n6564) );
  AOI22_X1 U5188 ( .A1(n3628), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4632) );
  AOI22_X1 U5189 ( .A1(n3649), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5261), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4631) );
  AOI22_X1 U5190 ( .A1(n4505), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4630) );
  AOI22_X1 U5191 ( .A1(n3658), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4629) );
  NAND4_X1 U5192 ( .A1(n4632), .A2(n4631), .A3(n4630), .A4(n4629), .ZN(n4638)
         );
  AOI22_X1 U5193 ( .A1(n5259), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3647), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4636) );
  AOI22_X1 U5194 ( .A1(n3627), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4689), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4635) );
  AOI22_X1 U5195 ( .A1(n3643), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4634) );
  AOI22_X1 U5196 ( .A1(n4010), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3656), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4633) );
  NAND4_X1 U5197 ( .A1(n4636), .A2(n4635), .A3(n4634), .A4(n4633), .ZN(n4637)
         );
  NOR2_X1 U5198 ( .A1(n4638), .A2(n4637), .ZN(n4652) );
  INV_X1 U5199 ( .A(n4639), .ZN(n4640) );
  XOR2_X1 U5200 ( .A(n4652), .B(n4651), .Z(n4642) );
  NAND2_X1 U5201 ( .A1(n4642), .A2(n5236), .ZN(n4647) );
  INV_X1 U5202 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6971) );
  AOI21_X1 U5203 ( .B1(n6971), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4643) );
  AOI21_X1 U5204 ( .B1(n6660), .B2(EAX_REG_25__SCAN_IN), .A(n4643), .ZN(n4646)
         );
  XNOR2_X1 U5205 ( .A(n4648), .B(n6971), .ZN(n6973) );
  AOI21_X1 U5206 ( .B1(n4647), .B2(n4646), .A(n4645), .ZN(n6737) );
  NAND2_X1 U5207 ( .A1(n4648), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4649)
         );
  INV_X1 U5208 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6727) );
  NAND2_X1 U5209 ( .A1(n4649), .A2(n6727), .ZN(n4650) );
  NAND2_X1 U5210 ( .A1(n4700), .A2(n4650), .ZN(n6964) );
  NOR2_X1 U5211 ( .A1(n4652), .A2(n4651), .ZN(n4678) );
  AOI22_X1 U5212 ( .A1(n3652), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4656) );
  AOI22_X1 U5213 ( .A1(n3644), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4655) );
  AOI22_X1 U5214 ( .A1(n4552), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4654) );
  AOI22_X1 U5215 ( .A1(n5261), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4653) );
  NAND4_X1 U5216 ( .A1(n4656), .A2(n4655), .A3(n4654), .A4(n4653), .ZN(n4662)
         );
  AOI22_X1 U5217 ( .A1(n3654), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4689), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4660) );
  AOI22_X1 U5218 ( .A1(n5259), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3655), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4659) );
  AOI22_X1 U5219 ( .A1(n4010), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4505), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4658) );
  AOI22_X1 U5220 ( .A1(n3647), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4657) );
  NAND4_X1 U5221 ( .A1(n4660), .A2(n4659), .A3(n4658), .A4(n4657), .ZN(n4661)
         );
  OR2_X1 U5222 ( .A1(n4662), .A2(n4661), .ZN(n4677) );
  XNOR2_X1 U5223 ( .A(n4678), .B(n4677), .ZN(n4664) );
  AOI22_X1 U5224 ( .A1(n6660), .A2(EAX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n5838), .ZN(n4663) );
  OAI21_X1 U5225 ( .B1(n4664), .B2(n5278), .A(n4663), .ZN(n4666) );
  MUX2_X1 U5226 ( .A(n6964), .B(n4666), .S(n4665), .Z(n6724) );
  AOI22_X1 U5227 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n4689), .B1(n5266), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4670) );
  AOI22_X1 U5228 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3661), .B1(n3660), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4669) );
  AOI22_X1 U5229 ( .A1(n5258), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4668) );
  AOI22_X1 U5230 ( .A1(n4505), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3655), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4667) );
  NAND4_X1 U5231 ( .A1(n4670), .A2(n4669), .A3(n4668), .A4(n4667), .ZN(n4676)
         );
  AOI22_X1 U5232 ( .A1(n5259), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4674) );
  AOI22_X1 U5233 ( .A1(n3653), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3651), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4673) );
  AOI22_X1 U5234 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3649), .B1(n5261), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4672) );
  AOI22_X1 U5235 ( .A1(n4352), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4671) );
  NAND4_X1 U5236 ( .A1(n4674), .A2(n4673), .A3(n4672), .A4(n4671), .ZN(n4675)
         );
  NOR2_X1 U5237 ( .A1(n4676), .A2(n4675), .ZN(n4684) );
  NAND2_X1 U5238 ( .A1(n4678), .A2(n4677), .ZN(n4683) );
  XOR2_X1 U5239 ( .A(n4684), .B(n4683), .Z(n4681) );
  INV_X1 U5240 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n6959) );
  NAND2_X1 U5241 ( .A1(n6660), .A2(EAX_REG_27__SCAN_IN), .ZN(n4679) );
  OAI21_X1 U5242 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6959), .A(n4679), .ZN(
        n4680) );
  AOI21_X1 U5243 ( .B1(n4681), .B2(n5236), .A(n4680), .ZN(n4682) );
  XNOR2_X1 U5244 ( .A(n4700), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n6961)
         );
  MUX2_X1 U5245 ( .A(n4682), .B(n6961), .S(n5282), .Z(n6711) );
  NOR2_X1 U5246 ( .A1(n4684), .A2(n4683), .ZN(n5235) );
  AOI22_X1 U5247 ( .A1(n3652), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4688) );
  AOI22_X1 U5248 ( .A1(n4352), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4687) );
  AOI22_X1 U5249 ( .A1(n4552), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4686) );
  AOI22_X1 U5250 ( .A1(n5261), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4685) );
  NAND4_X1 U5251 ( .A1(n4688), .A2(n4687), .A3(n4686), .A4(n4685), .ZN(n4695)
         );
  AOI22_X1 U5252 ( .A1(n3627), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4689), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4693) );
  AOI22_X1 U5253 ( .A1(n5259), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3657), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4692) );
  AOI22_X1 U5254 ( .A1(n4010), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4505), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4691) );
  AOI22_X1 U5255 ( .A1(n3647), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4690) );
  NAND4_X1 U5256 ( .A1(n4693), .A2(n4692), .A3(n4691), .A4(n4690), .ZN(n4694)
         );
  OR2_X1 U5257 ( .A1(n4695), .A2(n4694), .ZN(n5234) );
  INV_X1 U5258 ( .A(n5234), .ZN(n4696) );
  XNOR2_X1 U5259 ( .A(n5235), .B(n4696), .ZN(n4699) );
  INV_X1 U5260 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4712) );
  NAND2_X1 U5261 ( .A1(n6660), .A2(EAX_REG_28__SCAN_IN), .ZN(n4697) );
  OAI21_X1 U5262 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4712), .A(n4697), .ZN(
        n4698) );
  AOI21_X1 U5263 ( .B1(n4699), .B2(n5236), .A(n4698), .ZN(n4703) );
  AND2_X1 U5264 ( .A1(n4701), .A2(n4712), .ZN(n4702) );
  NOR2_X1 U5265 ( .A1(n5242), .A2(n4702), .ZN(n6631) );
  MUX2_X1 U5266 ( .A(n4703), .B(n6631), .S(n5282), .Z(n5245) );
  INV_X1 U5267 ( .A(n5245), .ZN(n4704) );
  NAND2_X1 U5268 ( .A1(n6710), .A2(n4704), .ZN(n5248) );
  NOR2_X2 U5269 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n5925) );
  NOR2_X1 U5270 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n7715), .ZN(n5370) );
  NAND2_X1 U5271 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n5370), .ZN(n7438) );
  INV_X1 U5272 ( .A(n7438), .ZN(n4707) );
  INV_X2 U5273 ( .A(n7052), .ZN(n7421) );
  NAND2_X1 U5274 ( .A1(n6375), .A2(n4708), .ZN(n7441) );
  NAND2_X1 U5275 ( .A1(n7441), .A2(n7437), .ZN(n4709) );
  NAND2_X1 U5276 ( .A1(n7437), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4711) );
  NAND2_X1 U5277 ( .A1(n7726), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4710) );
  NAND2_X1 U5278 ( .A1(n4711), .A2(n4710), .ZN(n5348) );
  NAND2_X1 U5279 ( .A1(n5925), .A2(n7715), .ZN(n7428) );
  INV_X1 U5280 ( .A(REIP_REG_28__SCAN_IN), .ZN(n7332) );
  OR2_X1 U5281 ( .A1(n7524), .A2(n7332), .ZN(n7075) );
  OAI21_X1 U5282 ( .B1(n7405), .B2(n4712), .A(n7075), .ZN(n4713) );
  AOI21_X1 U5283 ( .B1(n7409), .B2(n6631), .A(n4713), .ZN(n4714) );
  INV_X1 U5284 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n7243) );
  INV_X1 U5285 ( .A(keyinput_246), .ZN(n4898) );
  INV_X1 U5286 ( .A(DATAWIDTH_REG_10__SCAN_IN), .ZN(n7239) );
  INV_X1 U5287 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n7238) );
  AOI22_X1 U5288 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(keyinput_240), .B1(n7238), .B2(keyinput_241), .ZN(n4715) );
  OAI221_X1 U5289 ( .B1(DATAWIDTH_REG_8__SCAN_IN), .B2(keyinput_240), .C1(
        n7238), .C2(keyinput_241), .A(n4715), .ZN(n4891) );
  INV_X1 U5290 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n7331) );
  AOI22_X1 U5291 ( .A1(ADDRESS_REG_28__SCAN_IN), .A2(keyinput_200), .B1(n7331), 
        .B2(keyinput_201), .ZN(n4716) );
  OAI221_X1 U5292 ( .B1(ADDRESS_REG_28__SCAN_IN), .B2(keyinput_200), .C1(n7331), .C2(keyinput_201), .A(n4716), .ZN(n4837) );
  INV_X1 U5293 ( .A(keyinput_190), .ZN(n4820) );
  INV_X1 U5294 ( .A(REIP_REG_20__SCAN_IN), .ZN(n7315) );
  INV_X1 U5295 ( .A(keyinput_189), .ZN(n4818) );
  INV_X1 U5296 ( .A(REIP_REG_21__SCAN_IN), .ZN(n7317) );
  INV_X1 U5297 ( .A(REIP_REG_25__SCAN_IN), .ZN(n7326) );
  INV_X1 U5298 ( .A(keyinput_185), .ZN(n4809) );
  INV_X1 U5299 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n7747) );
  OAI22_X1 U5300 ( .A1(n7747), .A2(keyinput_168), .B1(keyinput_169), .B2(
        D_C_N_REG_SCAN_IN), .ZN(n4717) );
  AOI221_X1 U5301 ( .B1(n7747), .B2(keyinput_168), .C1(D_C_N_REG_SCAN_IN), 
        .C2(keyinput_169), .A(n4717), .ZN(n4788) );
  INV_X1 U5302 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n5341) );
  INV_X1 U5303 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n7429) );
  OAI22_X1 U5304 ( .A1(n7429), .A2(keyinput_165), .B1(keyinput_166), .B2(
        ADS_N_REG_SCAN_IN), .ZN(n4718) );
  AOI221_X1 U5305 ( .B1(n7429), .B2(keyinput_165), .C1(ADS_N_REG_SCAN_IN), 
        .C2(keyinput_166), .A(n4718), .ZN(n4785) );
  INV_X1 U5306 ( .A(DATAI_11_), .ZN(n6292) );
  OAI22_X1 U5307 ( .A1(DATAI_13_), .A2(keyinput_146), .B1(keyinput_147), .B2(
        DATAI_12_), .ZN(n4719) );
  AOI221_X1 U5308 ( .B1(DATAI_13_), .B2(keyinput_146), .C1(DATAI_12_), .C2(
        keyinput_147), .A(n4719), .ZN(n4759) );
  INV_X1 U5309 ( .A(DATAI_14_), .ZN(n6954) );
  INV_X1 U5310 ( .A(keyinput_145), .ZN(n4757) );
  INV_X1 U5311 ( .A(DATAI_16_), .ZN(n7749) );
  INV_X1 U5312 ( .A(keyinput_143), .ZN(n4751) );
  INV_X1 U5313 ( .A(DATAI_27_), .ZN(n4721) );
  AOI22_X1 U5314 ( .A1(DATAI_30_), .A2(keyinput_129), .B1(n4721), .B2(
        keyinput_132), .ZN(n4720) );
  OAI221_X1 U5315 ( .B1(DATAI_30_), .B2(keyinput_129), .C1(n4721), .C2(
        keyinput_132), .A(n4720), .ZN(n4727) );
  AOI22_X1 U5316 ( .A1(DATAI_28_), .A2(keyinput_131), .B1(DATAI_31_), .B2(
        keyinput_128), .ZN(n4722) );
  OAI221_X1 U5317 ( .B1(DATAI_28_), .B2(keyinput_131), .C1(DATAI_31_), .C2(
        keyinput_128), .A(n4722), .ZN(n4726) );
  XOR2_X1 U5318 ( .A(DATAI_29_), .B(keyinput_130), .Z(n4725) );
  INV_X1 U5319 ( .A(DATAI_26_), .ZN(n4723) );
  XNOR2_X1 U5320 ( .A(keyinput_133), .B(n4723), .ZN(n4724) );
  INV_X1 U5321 ( .A(keyinput_134), .ZN(n4728) );
  MUX2_X1 U5322 ( .A(n4728), .B(keyinput_134), .S(DATAI_25_), .Z(n4729) );
  NOR2_X1 U5323 ( .A1(n4730), .A2(n4729), .ZN(n4735) );
  INV_X1 U5324 ( .A(keyinput_135), .ZN(n4731) );
  MUX2_X1 U5325 ( .A(keyinput_135), .B(n4731), .S(DATAI_24_), .Z(n4734) );
  XOR2_X1 U5326 ( .A(DATAI_23_), .B(keyinput_136), .Z(n4733) );
  XNOR2_X1 U5327 ( .A(DATAI_22_), .B(keyinput_137), .ZN(n4732) );
  OAI211_X1 U5328 ( .C1(n4735), .C2(n4734), .A(n4733), .B(n4732), .ZN(n4741)
         );
  XOR2_X1 U5329 ( .A(DATAI_21_), .B(keyinput_138), .Z(n4740) );
  INV_X1 U5330 ( .A(keyinput_140), .ZN(n4738) );
  XNOR2_X1 U5331 ( .A(DATAI_20_), .B(keyinput_139), .ZN(n4737) );
  XNOR2_X1 U5332 ( .A(keyinput_141), .B(DATAI_18_), .ZN(n4736) );
  OAI211_X1 U5333 ( .C1(n4738), .C2(DATAI_19_), .A(n4737), .B(n4736), .ZN(
        n4739) );
  AOI21_X1 U5334 ( .B1(n4741), .B2(n4740), .A(n4739), .ZN(n4742) );
  INV_X1 U5335 ( .A(n4742), .ZN(n4749) );
  INV_X1 U5336 ( .A(DATAI_19_), .ZN(n4743) );
  NOR2_X1 U5337 ( .A1(n4743), .A2(keyinput_140), .ZN(n4748) );
  INV_X1 U5338 ( .A(DATAI_17_), .ZN(n4745) );
  INV_X1 U5339 ( .A(keyinput_142), .ZN(n4744) );
  OAI21_X1 U5340 ( .B1(n4749), .B2(n4748), .A(n4747), .ZN(n4750) );
  OAI221_X1 U5341 ( .B1(DATAI_16_), .B2(keyinput_143), .C1(n7749), .C2(n4751), 
        .A(n4750), .ZN(n4755) );
  INV_X1 U5342 ( .A(DATAI_15_), .ZN(n6950) );
  INV_X1 U5343 ( .A(keyinput_144), .ZN(n4752) );
  NAND2_X1 U5344 ( .A1(n4755), .A2(n4754), .ZN(n4756) );
  OAI221_X1 U5345 ( .B1(DATAI_14_), .B2(keyinput_145), .C1(n6954), .C2(n4757), 
        .A(n4756), .ZN(n4758) );
  AOI22_X1 U5346 ( .A1(keyinput_148), .A2(n6292), .B1(n4759), .B2(n4758), .ZN(
        n4760) );
  OAI21_X1 U5347 ( .B1(n6292), .B2(keyinput_148), .A(n4760), .ZN(n4766) );
  INV_X1 U5348 ( .A(DATAI_7_), .ZN(n6069) );
  INV_X1 U5349 ( .A(DATAI_6_), .ZN(n6086) );
  OAI22_X1 U5350 ( .A1(n6069), .A2(keyinput_152), .B1(n6086), .B2(keyinput_153), .ZN(n4761) );
  AOI221_X1 U5351 ( .B1(n6069), .B2(keyinput_152), .C1(keyinput_153), .C2(
        n6086), .A(n4761), .ZN(n4765) );
  INV_X1 U5352 ( .A(DATAI_10_), .ZN(n6278) );
  OAI22_X1 U5353 ( .A1(n6278), .A2(keyinput_149), .B1(DATAI_9_), .B2(
        keyinput_150), .ZN(n4762) );
  AOI221_X1 U5354 ( .B1(n6278), .B2(keyinput_149), .C1(keyinput_150), .C2(
        DATAI_9_), .A(n4762), .ZN(n4764) );
  INV_X1 U5355 ( .A(DATAI_8_), .ZN(n6936) );
  XNOR2_X1 U5356 ( .A(n6936), .B(keyinput_151), .ZN(n4763) );
  NAND4_X1 U5357 ( .A1(n4766), .A2(n4765), .A3(n4764), .A4(n4763), .ZN(n4769)
         );
  INV_X1 U5358 ( .A(DATAI_4_), .ZN(n6091) );
  OAI22_X1 U5359 ( .A1(n6091), .A2(keyinput_155), .B1(keyinput_154), .B2(
        DATAI_5_), .ZN(n4767) );
  AOI221_X1 U5360 ( .B1(n6091), .B2(keyinput_155), .C1(DATAI_5_), .C2(
        keyinput_154), .A(n4767), .ZN(n4768) );
  INV_X1 U5361 ( .A(BS16_N), .ZN(n7228) );
  XNOR2_X1 U5362 ( .A(n7228), .B(keyinput_162), .ZN(n4779) );
  INV_X1 U5363 ( .A(READY_N), .ZN(n7442) );
  INV_X1 U5364 ( .A(DATAI_1_), .ZN(n6071) );
  AOI22_X1 U5365 ( .A1(n7442), .A2(keyinput_163), .B1(keyinput_158), .B2(n6071), .ZN(n4773) );
  OAI221_X1 U5366 ( .B1(n7442), .B2(keyinput_163), .C1(n6071), .C2(
        keyinput_158), .A(n4773), .ZN(n4778) );
  INV_X1 U5367 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n7748) );
  AOI22_X1 U5368 ( .A1(NA_N), .A2(keyinput_161), .B1(n7748), .B2(keyinput_160), 
        .ZN(n4774) );
  OAI221_X1 U5369 ( .B1(NA_N), .B2(keyinput_161), .C1(n7748), .C2(keyinput_160), .A(n4774), .ZN(n4777) );
  INV_X1 U5370 ( .A(DATAI_2_), .ZN(n6085) );
  AOI22_X1 U5371 ( .A1(DATAI_0_), .A2(keyinput_159), .B1(n6085), .B2(
        keyinput_157), .ZN(n4775) );
  OAI221_X1 U5372 ( .B1(DATAI_0_), .B2(keyinput_159), .C1(n6085), .C2(
        keyinput_157), .A(n4775), .ZN(n4776) );
  NOR4_X1 U5373 ( .A1(n4779), .A2(n4778), .A3(n4777), .A4(n4776), .ZN(n4781)
         );
  INV_X1 U5374 ( .A(HOLD), .ZN(n7735) );
  INV_X1 U5375 ( .A(n4783), .ZN(n4784) );
  AOI22_X1 U5376 ( .A1(keyinput_167), .A2(n5341), .B1(n4785), .B2(n4784), .ZN(
        n4786) );
  OAI21_X1 U5377 ( .B1(n5341), .B2(keyinput_167), .A(n4786), .ZN(n4787) );
  OAI211_X1 U5378 ( .C1(REQUESTPENDING_REG_SCAN_IN), .C2(keyinput_170), .A(
        n4788), .B(n4787), .ZN(n4789) );
  AOI21_X1 U5379 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_170), .A(
        n4789), .ZN(n4799) );
  INV_X1 U5380 ( .A(FLUSH_REG_SCAN_IN), .ZN(n7702) );
  OAI22_X1 U5381 ( .A1(n7702), .A2(keyinput_173), .B1(keyinput_174), .B2(
        W_R_N_REG_SCAN_IN), .ZN(n4790) );
  AOI221_X1 U5382 ( .B1(n7702), .B2(keyinput_173), .C1(W_R_N_REG_SCAN_IN), 
        .C2(keyinput_174), .A(n4790), .ZN(n4797) );
  INV_X1 U5383 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n7363) );
  INV_X1 U5384 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n7340) );
  OAI22_X1 U5385 ( .A1(n7363), .A2(keyinput_175), .B1(n7340), .B2(keyinput_178), .ZN(n4791) );
  AOI221_X1 U5386 ( .B1(n7363), .B2(keyinput_175), .C1(keyinput_178), .C2(
        n7340), .A(n4791), .ZN(n4796) );
  OAI22_X1 U5387 ( .A1(BYTEENABLE_REG_2__SCAN_IN), .A2(keyinput_177), .B1(
        MORE_REG_SCAN_IN), .B2(keyinput_172), .ZN(n4792) );
  AOI221_X1 U5388 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_177), .C1(
        keyinput_172), .C2(MORE_REG_SCAN_IN), .A(n4792), .ZN(n4795) );
  OAI22_X1 U5389 ( .A1(STATEBS16_REG_SCAN_IN), .A2(keyinput_171), .B1(
        keyinput_176), .B2(BYTEENABLE_REG_1__SCAN_IN), .ZN(n4793) );
  AOI221_X1 U5390 ( .B1(STATEBS16_REG_SCAN_IN), .B2(keyinput_171), .C1(
        BYTEENABLE_REG_1__SCAN_IN), .C2(keyinput_176), .A(n4793), .ZN(n4794)
         );
  NAND4_X1 U5391 ( .A1(n4797), .A2(n4796), .A3(n4795), .A4(n4794), .ZN(n4798)
         );
  OAI22_X1 U5392 ( .A1(REIP_REG_30__SCAN_IN), .A2(keyinput_180), .B1(
        keyinput_183), .B2(REIP_REG_27__SCAN_IN), .ZN(n4800) );
  AOI221_X1 U5393 ( .B1(REIP_REG_30__SCAN_IN), .B2(keyinput_180), .C1(
        REIP_REG_27__SCAN_IN), .C2(keyinput_183), .A(n4800), .ZN(n4801) );
  INV_X1 U5394 ( .A(REIP_REG_29__SCAN_IN), .ZN(n7333) );
  AOI22_X1 U5395 ( .A1(n7333), .A2(keyinput_181), .B1(keyinput_182), .B2(n7332), .ZN(n4804) );
  OAI221_X1 U5396 ( .B1(n7333), .B2(keyinput_181), .C1(n7332), .C2(
        keyinput_182), .A(n4804), .ZN(n4805) );
  OAI22_X1 U5397 ( .A1(n4806), .A2(n4805), .B1(keyinput_184), .B2(
        REIP_REG_26__SCAN_IN), .ZN(n4807) );
  AOI21_X1 U5398 ( .B1(keyinput_184), .B2(REIP_REG_26__SCAN_IN), .A(n4807), 
        .ZN(n4808) );
  AOI221_X1 U5399 ( .B1(REIP_REG_25__SCAN_IN), .B2(keyinput_185), .C1(n7326), 
        .C2(n4809), .A(n4808), .ZN(n4816) );
  INV_X1 U5400 ( .A(REIP_REG_22__SCAN_IN), .ZN(n7318) );
  INV_X1 U5401 ( .A(REIP_REG_24__SCAN_IN), .ZN(n7323) );
  AOI22_X1 U5402 ( .A1(n7318), .A2(keyinput_188), .B1(n7323), .B2(keyinput_186), .ZN(n4810) );
  OAI221_X1 U5403 ( .B1(n7318), .B2(keyinput_188), .C1(n7323), .C2(
        keyinput_186), .A(n4810), .ZN(n4811) );
  INV_X1 U5404 ( .A(n4811), .ZN(n4814) );
  INV_X1 U5405 ( .A(REIP_REG_23__SCAN_IN), .ZN(n7322) );
  OR2_X1 U5406 ( .A1(n4816), .A2(n4815), .ZN(n4817) );
  OAI221_X1 U5407 ( .B1(REIP_REG_21__SCAN_IN), .B2(n4818), .C1(n7317), .C2(
        keyinput_189), .A(n4817), .ZN(n4819) );
  OAI221_X1 U5408 ( .B1(REIP_REG_20__SCAN_IN), .B2(n4820), .C1(n7315), .C2(
        keyinput_190), .A(n4819), .ZN(n4823) );
  INV_X1 U5409 ( .A(REIP_REG_18__SCAN_IN), .ZN(n7671) );
  INV_X1 U5410 ( .A(REIP_REG_19__SCAN_IN), .ZN(n7673) );
  OAI22_X1 U5411 ( .A1(n7671), .A2(keyinput_192), .B1(n7673), .B2(keyinput_191), .ZN(n4821) );
  AOI221_X1 U5412 ( .B1(n7671), .B2(keyinput_192), .C1(keyinput_191), .C2(
        n7673), .A(n4821), .ZN(n4822) );
  INV_X1 U5413 ( .A(REIP_REG_16__SCAN_IN), .ZN(n7525) );
  AOI22_X1 U5414 ( .A1(REIP_REG_17__SCAN_IN), .A2(keyinput_193), .B1(n7525), 
        .B2(keyinput_194), .ZN(n4824) );
  OAI221_X1 U5415 ( .B1(REIP_REG_17__SCAN_IN), .B2(keyinput_193), .C1(n7525), 
        .C2(keyinput_194), .A(n4824), .ZN(n4825) );
  INV_X1 U5416 ( .A(n4825), .ZN(n4831) );
  OAI22_X1 U5417 ( .A1(BE_N_REG_2__SCAN_IN), .A2(keyinput_196), .B1(
        BE_N_REG_0__SCAN_IN), .B2(keyinput_198), .ZN(n4826) );
  AOI221_X1 U5418 ( .B1(BE_N_REG_2__SCAN_IN), .B2(keyinput_196), .C1(
        keyinput_198), .C2(BE_N_REG_0__SCAN_IN), .A(n4826), .ZN(n4830) );
  INV_X1 U5419 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n7357) );
  INV_X1 U5420 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n7339) );
  AOI22_X1 U5421 ( .A1(n7357), .A2(keyinput_197), .B1(n7339), .B2(keyinput_195), .ZN(n4827) );
  OAI221_X1 U5422 ( .B1(n7357), .B2(keyinput_197), .C1(n7339), .C2(
        keyinput_195), .A(n4827), .ZN(n4828) );
  INV_X1 U5423 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n7336) );
  INV_X1 U5424 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n7329) );
  NAND2_X1 U5425 ( .A1(n7329), .A2(keyinput_202), .ZN(n4835) );
  OAI221_X1 U5426 ( .B1(n4837), .B2(n4836), .C1(n7329), .C2(keyinput_202), .A(
        n4835), .ZN(n4840) );
  INV_X1 U5427 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n7327) );
  OAI22_X1 U5428 ( .A1(n7327), .A2(keyinput_203), .B1(ADDRESS_REG_24__SCAN_IN), 
        .B2(keyinput_204), .ZN(n4838) );
  AOI221_X1 U5429 ( .B1(n7327), .B2(keyinput_203), .C1(keyinput_204), .C2(
        ADDRESS_REG_24__SCAN_IN), .A(n4838), .ZN(n4839) );
  INV_X1 U5430 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n7324) );
  INV_X1 U5431 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n7319) );
  AOI22_X1 U5432 ( .A1(ADDRESS_REG_22__SCAN_IN), .A2(keyinput_206), .B1(n7319), 
        .B2(keyinput_207), .ZN(n4841) );
  OAI221_X1 U5433 ( .B1(ADDRESS_REG_22__SCAN_IN), .B2(keyinput_206), .C1(n7319), .C2(keyinput_207), .A(n4841), .ZN(n4842) );
  AOI221_X1 U5434 ( .B1(keyinput_205), .B2(n4843), .C1(n7324), .C2(n4843), .A(
        n4842), .ZN(n4846) );
  INV_X1 U5435 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n7314) );
  INV_X1 U5436 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n7316) );
  OAI22_X1 U5437 ( .A1(n7314), .A2(keyinput_209), .B1(n7316), .B2(keyinput_208), .ZN(n4844) );
  AOI221_X1 U5438 ( .B1(n7314), .B2(keyinput_209), .C1(keyinput_208), .C2(
        n7316), .A(n4844), .ZN(n4845) );
  INV_X1 U5439 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n7313) );
  INV_X1 U5440 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n7312) );
  AOI22_X1 U5441 ( .A1(n7313), .A2(keyinput_210), .B1(keyinput_211), .B2(n7312), .ZN(n4847) );
  OAI221_X1 U5442 ( .B1(n7313), .B2(keyinput_210), .C1(n7312), .C2(
        keyinput_211), .A(n4847), .ZN(n4850) );
  INV_X1 U5443 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n7309) );
  INV_X1 U5444 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n7310) );
  AOI22_X1 U5445 ( .A1(n7309), .A2(keyinput_213), .B1(n7310), .B2(keyinput_212), .ZN(n4848) );
  OAI221_X1 U5446 ( .B1(n7309), .B2(keyinput_213), .C1(n7310), .C2(
        keyinput_212), .A(n4848), .ZN(n4849) );
  NOR2_X1 U5447 ( .A1(n4850), .A2(n4849), .ZN(n4855) );
  INV_X1 U5448 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n7307) );
  INV_X1 U5449 ( .A(keyinput_214), .ZN(n4851) );
  NAND2_X1 U5450 ( .A1(n7307), .A2(n4851), .ZN(n4853) );
  INV_X1 U5451 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n7293) );
  INV_X1 U5452 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n7298) );
  AOI22_X1 U5453 ( .A1(n7293), .A2(keyinput_225), .B1(n7298), .B2(keyinput_222), .ZN(n4857) );
  OAI221_X1 U5454 ( .B1(n7293), .B2(keyinput_225), .C1(n7298), .C2(
        keyinput_222), .A(n4857), .ZN(n4869) );
  INV_X1 U5455 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n7294) );
  INV_X1 U5456 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n7297) );
  AOI22_X1 U5457 ( .A1(n7294), .A2(keyinput_224), .B1(keyinput_223), .B2(n7297), .ZN(n4858) );
  OAI221_X1 U5458 ( .B1(n7294), .B2(keyinput_224), .C1(n7297), .C2(
        keyinput_223), .A(n4858), .ZN(n4868) );
  OAI22_X1 U5459 ( .A1(ADDRESS_REG_10__SCAN_IN), .A2(keyinput_218), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(keyinput_219), .ZN(n4859) );
  AOI221_X1 U5460 ( .B1(ADDRESS_REG_10__SCAN_IN), .B2(keyinput_218), .C1(
        keyinput_219), .C2(ADDRESS_REG_9__SCAN_IN), .A(n4859), .ZN(n4866) );
  OAI22_X1 U5461 ( .A1(ADDRESS_REG_8__SCAN_IN), .A2(keyinput_220), .B1(
        keyinput_216), .B2(ADDRESS_REG_12__SCAN_IN), .ZN(n4860) );
  AOI221_X1 U5462 ( .B1(ADDRESS_REG_8__SCAN_IN), .B2(keyinput_220), .C1(
        ADDRESS_REG_12__SCAN_IN), .C2(keyinput_216), .A(n4860), .ZN(n4865) );
  INV_X1 U5463 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n7306) );
  INV_X1 U5464 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n7291) );
  OAI22_X1 U5465 ( .A1(n7306), .A2(keyinput_215), .B1(n7291), .B2(keyinput_226), .ZN(n4861) );
  AOI221_X1 U5466 ( .B1(n7306), .B2(keyinput_215), .C1(keyinput_226), .C2(
        n7291), .A(n4861), .ZN(n4864) );
  OAI22_X1 U5467 ( .A1(ADDRESS_REG_11__SCAN_IN), .A2(keyinput_217), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(keyinput_221), .ZN(n4862) );
  AOI221_X1 U5468 ( .B1(ADDRESS_REG_11__SCAN_IN), .B2(keyinput_217), .C1(
        keyinput_221), .C2(ADDRESS_REG_7__SCAN_IN), .A(n4862), .ZN(n4863) );
  NAND4_X1 U5469 ( .A1(n4866), .A2(n4865), .A3(n4864), .A4(n4863), .ZN(n4867)
         );
  INV_X1 U5470 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n7289) );
  INV_X1 U5471 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n7288) );
  AOI22_X1 U5472 ( .A1(n7289), .A2(keyinput_227), .B1(keyinput_228), .B2(n7288), .ZN(n4871) );
  OAI221_X1 U5473 ( .B1(n7289), .B2(keyinput_227), .C1(n7288), .C2(
        keyinput_228), .A(n4871), .ZN(n4874) );
  OAI22_X1 U5474 ( .A1(n7737), .A2(keyinput_229), .B1(n7433), .B2(keyinput_230), .ZN(n4872) );
  AOI221_X1 U5475 ( .B1(n7737), .B2(keyinput_229), .C1(keyinput_230), .C2(
        n7433), .A(n4872), .ZN(n4873) );
  OAI21_X1 U5476 ( .B1(n4875), .B2(n4874), .A(n4873), .ZN(n4879) );
  INV_X1 U5477 ( .A(STATE_REG_0__SCAN_IN), .ZN(n7736) );
  INV_X1 U5478 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n7229) );
  OAI22_X1 U5479 ( .A1(n7736), .A2(keyinput_231), .B1(n7229), .B2(keyinput_232), .ZN(n4876) );
  AOI221_X1 U5480 ( .B1(n7736), .B2(keyinput_231), .C1(keyinput_232), .C2(
        n7229), .A(n4876), .ZN(n4878) );
  INV_X1 U5481 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n7728) );
  NOR2_X1 U5482 ( .A1(n7728), .A2(keyinput_233), .ZN(n4877) );
  AOI221_X1 U5483 ( .B1(n4879), .B2(n4878), .C1(keyinput_233), .C2(n7728), .A(
        n4877), .ZN(n4880) );
  INV_X1 U5484 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n7234) );
  INV_X1 U5485 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n7235) );
  AOI22_X1 U5486 ( .A1(n7234), .A2(keyinput_237), .B1(keyinput_238), .B2(n7235), .ZN(n4881) );
  OAI221_X1 U5487 ( .B1(n7234), .B2(keyinput_237), .C1(n7235), .C2(
        keyinput_238), .A(n4881), .ZN(n4884) );
  INV_X1 U5488 ( .A(DATAWIDTH_REG_4__SCAN_IN), .ZN(n7233) );
  INV_X1 U5489 ( .A(DATAWIDTH_REG_3__SCAN_IN), .ZN(n7232) );
  AOI22_X1 U5490 ( .A1(n7233), .A2(keyinput_236), .B1(keyinput_235), .B2(n7232), .ZN(n4882) );
  OAI221_X1 U5491 ( .B1(n7233), .B2(keyinput_236), .C1(n7232), .C2(
        keyinput_235), .A(n4882), .ZN(n4883) );
  AOI211_X1 U5492 ( .C1(keyinput_234), .C2(DATAWIDTH_REG_2__SCAN_IN), .A(n4884), .B(n4883), .ZN(n4885) );
  OAI21_X1 U5493 ( .B1(keyinput_234), .B2(DATAWIDTH_REG_2__SCAN_IN), .A(n4885), 
        .ZN(n4886) );
  INV_X1 U5494 ( .A(n4886), .ZN(n4888) );
  OAI22_X1 U5495 ( .A1(keyinput_242), .A2(n7239), .B1(n4891), .B2(n4890), .ZN(
        n4892) );
  AOI21_X1 U5496 ( .B1(keyinput_242), .B2(n7239), .A(n4892), .ZN(n4896) );
  INV_X1 U5497 ( .A(DATAWIDTH_REG_13__SCAN_IN), .ZN(n7242) );
  AOI22_X1 U5498 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(keyinput_244), .B1(
        n7242), .B2(keyinput_245), .ZN(n4893) );
  OAI221_X1 U5499 ( .B1(DATAWIDTH_REG_12__SCAN_IN), .B2(keyinput_244), .C1(
        n7242), .C2(keyinput_245), .A(n4893), .ZN(n4895) );
  OR2_X1 U5500 ( .A1(n4896), .A2(n3744), .ZN(n4897) );
  OAI221_X1 U5501 ( .B1(DATAWIDTH_REG_14__SCAN_IN), .B2(keyinput_246), .C1(
        n7243), .C2(n4898), .A(n4897), .ZN(n4902) );
  INV_X1 U5502 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n7244) );
  INV_X1 U5503 ( .A(keyinput_247), .ZN(n4899) );
  OAI22_X1 U5504 ( .A1(n7244), .A2(n4899), .B1(DATAWIDTH_REG_15__SCAN_IN), 
        .B2(keyinput_247), .ZN(n4900) );
  INV_X1 U5505 ( .A(n4900), .ZN(n4901) );
  INV_X1 U5506 ( .A(DATAWIDTH_REG_16__SCAN_IN), .ZN(n7245) );
  INV_X1 U5507 ( .A(DATAWIDTH_REG_17__SCAN_IN), .ZN(n7246) );
  OAI22_X1 U5508 ( .A1(n7245), .A2(keyinput_248), .B1(n7246), .B2(keyinput_249), .ZN(n4903) );
  AOI221_X1 U5509 ( .B1(n7245), .B2(keyinput_248), .C1(keyinput_249), .C2(
        n7246), .A(n4903), .ZN(n4906) );
  INV_X1 U5510 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n7247) );
  XNOR2_X1 U5511 ( .A(n7247), .B(keyinput_251), .ZN(n4913) );
  INV_X1 U5512 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n7248) );
  XNOR2_X1 U5513 ( .A(n7248), .B(keyinput_253), .ZN(n4911) );
  INV_X1 U5514 ( .A(DATAWIDTH_REG_22__SCAN_IN), .ZN(n7249) );
  XNOR2_X1 U5515 ( .A(n7249), .B(keyinput_254), .ZN(n4910) );
  XNOR2_X1 U5516 ( .A(keyinput_252), .B(DATAWIDTH_REG_20__SCAN_IN), .ZN(n4909)
         );
  NOR3_X1 U5517 ( .A1(n4911), .A2(n4910), .A3(n4909), .ZN(n4912) );
  OAI21_X1 U5518 ( .B1(n4914), .B2(n4913), .A(n4912), .ZN(n5106) );
  XOR2_X1 U5519 ( .A(DATAI_31_), .B(keyinput_0), .Z(n4916) );
  XOR2_X1 U5520 ( .A(DATAI_30_), .B(keyinput_1), .Z(n4915) );
  NAND2_X1 U5521 ( .A1(n4916), .A2(n4915), .ZN(n4925) );
  INV_X1 U5522 ( .A(keyinput_5), .ZN(n4917) );
  XNOR2_X1 U5523 ( .A(n4917), .B(DATAI_26_), .ZN(n4922) );
  INV_X1 U5524 ( .A(keyinput_4), .ZN(n4918) );
  XNOR2_X1 U5525 ( .A(n4918), .B(DATAI_27_), .ZN(n4921) );
  XNOR2_X1 U5526 ( .A(DATAI_29_), .B(keyinput_2), .ZN(n4920) );
  XNOR2_X1 U5527 ( .A(DATAI_28_), .B(keyinput_3), .ZN(n4919) );
  NAND4_X1 U5528 ( .A1(n4922), .A2(n4921), .A3(n4920), .A4(n4919), .ZN(n4924)
         );
  XOR2_X1 U5529 ( .A(keyinput_6), .B(DATAI_25_), .Z(n4923) );
  OAI21_X1 U5530 ( .B1(n4925), .B2(n4924), .A(n4923), .ZN(n4929) );
  XOR2_X1 U5531 ( .A(keyinput_7), .B(DATAI_24_), .Z(n4928) );
  XOR2_X1 U5532 ( .A(keyinput_9), .B(DATAI_22_), .Z(n4927) );
  XOR2_X1 U5533 ( .A(keyinput_8), .B(DATAI_23_), .Z(n4926) );
  AOI211_X1 U5534 ( .C1(n4929), .C2(n4928), .A(n4927), .B(n4926), .ZN(n4935)
         );
  XOR2_X1 U5535 ( .A(keyinput_10), .B(DATAI_21_), .Z(n4934) );
  XOR2_X1 U5536 ( .A(keyinput_12), .B(DATAI_19_), .Z(n4932) );
  XOR2_X1 U5537 ( .A(keyinput_11), .B(DATAI_20_), .Z(n4931) );
  XNOR2_X1 U5538 ( .A(keyinput_13), .B(DATAI_18_), .ZN(n4930) );
  NOR3_X1 U5539 ( .A1(n4932), .A2(n4931), .A3(n4930), .ZN(n4933) );
  OAI21_X1 U5540 ( .B1(n4935), .B2(n4934), .A(n4933), .ZN(n4938) );
  XOR2_X1 U5541 ( .A(keyinput_14), .B(DATAI_17_), .Z(n4937) );
  XNOR2_X1 U5542 ( .A(keyinput_15), .B(DATAI_16_), .ZN(n4936) );
  AOI21_X1 U5543 ( .B1(n4938), .B2(n4937), .A(n4936), .ZN(n4941) );
  XOR2_X1 U5544 ( .A(keyinput_16), .B(DATAI_15_), .Z(n4940) );
  XOR2_X1 U5545 ( .A(DATAI_14_), .B(keyinput_17), .Z(n4939) );
  OAI21_X1 U5546 ( .B1(n4941), .B2(n4940), .A(n4939), .ZN(n4944) );
  XOR2_X1 U5547 ( .A(DATAI_12_), .B(keyinput_19), .Z(n4943) );
  XNOR2_X1 U5548 ( .A(DATAI_13_), .B(keyinput_18), .ZN(n4942) );
  NAND3_X1 U5549 ( .A1(n4944), .A2(n4943), .A3(n4942), .ZN(n4953) );
  XOR2_X1 U5550 ( .A(DATAI_11_), .B(keyinput_20), .Z(n4952) );
  XOR2_X1 U5551 ( .A(keyinput_25), .B(DATAI_6_), .Z(n4947) );
  XOR2_X1 U5552 ( .A(DATAI_10_), .B(keyinput_21), .Z(n4946) );
  XNOR2_X1 U5553 ( .A(DATAI_7_), .B(keyinput_24), .ZN(n4945) );
  NOR3_X1 U5554 ( .A1(n4947), .A2(n4946), .A3(n4945), .ZN(n4950) );
  XOR2_X1 U5555 ( .A(DATAI_9_), .B(keyinput_22), .Z(n4949) );
  XOR2_X1 U5556 ( .A(keyinput_23), .B(DATAI_8_), .Z(n4948) );
  NAND3_X1 U5557 ( .A1(n4950), .A2(n4949), .A3(n4948), .ZN(n4951) );
  AOI21_X1 U5558 ( .B1(n4953), .B2(n4952), .A(n4951), .ZN(n4956) );
  XOR2_X1 U5559 ( .A(keyinput_26), .B(DATAI_5_), .Z(n4955) );
  XOR2_X1 U5560 ( .A(keyinput_27), .B(DATAI_4_), .Z(n4954) );
  NOR3_X1 U5561 ( .A1(n4956), .A2(n4955), .A3(n4954), .ZN(n4968) );
  XOR2_X1 U5562 ( .A(keyinput_28), .B(DATAI_3_), .Z(n4967) );
  OAI22_X1 U5563 ( .A1(keyinput_32), .A2(MEMORYFETCH_REG_SCAN_IN), .B1(READY_N), .B2(keyinput_35), .ZN(n4964) );
  OAI22_X1 U5564 ( .A1(n7228), .A2(keyinput_34), .B1(keyinput_33), .B2(NA_N), 
        .ZN(n4963) );
  INV_X1 U5565 ( .A(DATAI_0_), .ZN(n6072) );
  NOR2_X1 U5566 ( .A1(n6072), .A2(keyinput_31), .ZN(n4962) );
  AOI22_X1 U5567 ( .A1(n7228), .A2(keyinput_34), .B1(keyinput_31), .B2(n6072), 
        .ZN(n4959) );
  AOI22_X1 U5568 ( .A1(DATAI_1_), .A2(keyinput_30), .B1(READY_N), .B2(
        keyinput_35), .ZN(n4958) );
  AOI22_X1 U5569 ( .A1(NA_N), .A2(keyinput_33), .B1(MEMORYFETCH_REG_SCAN_IN), 
        .B2(keyinput_32), .ZN(n4957) );
  AND3_X1 U5570 ( .A1(n4959), .A2(n4958), .A3(n4957), .ZN(n4960) );
  OAI21_X1 U5571 ( .B1(keyinput_30), .B2(DATAI_1_), .A(n4960), .ZN(n4961) );
  NOR4_X1 U5572 ( .A1(n4964), .A2(n4963), .A3(n4962), .A4(n4961), .ZN(n4966)
         );
  XNOR2_X1 U5573 ( .A(keyinput_29), .B(DATAI_2_), .ZN(n4965) );
  OAI211_X1 U5574 ( .C1(n4968), .C2(n4967), .A(n4966), .B(n4965), .ZN(n4972)
         );
  XOR2_X1 U5575 ( .A(HOLD), .B(keyinput_36), .Z(n4971) );
  INV_X1 U5576 ( .A(ADS_N_REG_SCAN_IN), .ZN(n7253) );
  XNOR2_X1 U5577 ( .A(n7253), .B(keyinput_38), .ZN(n4970) );
  XNOR2_X1 U5578 ( .A(READREQUEST_REG_SCAN_IN), .B(keyinput_37), .ZN(n4969) );
  AOI211_X1 U5579 ( .C1(n4972), .C2(n4971), .A(n4970), .B(n4969), .ZN(n4978)
         );
  XOR2_X1 U5580 ( .A(keyinput_39), .B(CODEFETCH_REG_SCAN_IN), .Z(n4977) );
  XOR2_X1 U5581 ( .A(keyinput_40), .B(M_IO_N_REG_SCAN_IN), .Z(n4975) );
  XOR2_X1 U5582 ( .A(D_C_N_REG_SCAN_IN), .B(keyinput_41), .Z(n4974) );
  XOR2_X1 U5583 ( .A(keyinput_42), .B(REQUESTPENDING_REG_SCAN_IN), .Z(n4973)
         );
  NOR3_X1 U5584 ( .A1(n4975), .A2(n4974), .A3(n4973), .ZN(n4976) );
  OAI21_X1 U5585 ( .B1(n4978), .B2(n4977), .A(n4976), .ZN(n4992) );
  INV_X1 U5586 ( .A(W_R_N_REG_SCAN_IN), .ZN(n7432) );
  INV_X1 U5587 ( .A(MORE_REG_SCAN_IN), .ZN(n7202) );
  AOI22_X1 U5588 ( .A1(keyinput_46), .A2(n7432), .B1(n7202), .B2(keyinput_44), 
        .ZN(n4991) );
  AOI22_X1 U5589 ( .A1(FLUSH_REG_SCAN_IN), .A2(keyinput_45), .B1(keyinput_48), 
        .B2(BYTEENABLE_REG_1__SCAN_IN), .ZN(n4990) );
  INV_X1 U5590 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n7356) );
  INV_X1 U5591 ( .A(keyinput_43), .ZN(n4984) );
  OAI22_X1 U5592 ( .A1(STATEBS16_REG_SCAN_IN), .A2(keyinput_43), .B1(
        BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_48), .ZN(n4982) );
  OAI22_X1 U5593 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_50), .B1(
        FLUSH_REG_SCAN_IN), .B2(keyinput_45), .ZN(n4981) );
  OAI22_X1 U5594 ( .A1(n7432), .A2(keyinput_46), .B1(n7202), .B2(keyinput_44), 
        .ZN(n4980) );
  OAI22_X1 U5595 ( .A1(n7363), .A2(keyinput_47), .B1(n7356), .B2(keyinput_49), 
        .ZN(n4979) );
  NOR4_X1 U5596 ( .A1(n4982), .A2(n4981), .A3(n4980), .A4(n4979), .ZN(n4983)
         );
  OAI21_X1 U5597 ( .B1(n7726), .B2(n4984), .A(n4983), .ZN(n4988) );
  INV_X1 U5598 ( .A(keyinput_50), .ZN(n4986) );
  INV_X1 U5599 ( .A(keyinput_47), .ZN(n4985) );
  OAI22_X1 U5600 ( .A1(n7340), .A2(n4986), .B1(n4985), .B2(
        BYTEENABLE_REG_0__SCAN_IN), .ZN(n4987) );
  AOI211_X1 U5601 ( .C1(keyinput_49), .C2(n7356), .A(n4988), .B(n4987), .ZN(
        n4989) );
  NAND4_X1 U5602 ( .A1(n4992), .A2(n4991), .A3(n4990), .A4(n4989), .ZN(n4999)
         );
  XOR2_X1 U5603 ( .A(REIP_REG_31__SCAN_IN), .B(keyinput_51), .Z(n4998) );
  XOR2_X1 U5604 ( .A(REIP_REG_30__SCAN_IN), .B(keyinput_52), .Z(n4996) );
  XOR2_X1 U5605 ( .A(REIP_REG_28__SCAN_IN), .B(keyinput_54), .Z(n4995) );
  XOR2_X1 U5606 ( .A(REIP_REG_27__SCAN_IN), .B(keyinput_55), .Z(n4994) );
  XNOR2_X1 U5607 ( .A(REIP_REG_29__SCAN_IN), .B(keyinput_53), .ZN(n4993) );
  NAND4_X1 U5608 ( .A1(n4996), .A2(n4995), .A3(n4994), .A4(n4993), .ZN(n4997)
         );
  AOI21_X1 U5609 ( .B1(n4999), .B2(n4998), .A(n4997), .ZN(n5002) );
  XOR2_X1 U5610 ( .A(REIP_REG_26__SCAN_IN), .B(keyinput_56), .Z(n5001) );
  XNOR2_X1 U5611 ( .A(REIP_REG_25__SCAN_IN), .B(keyinput_57), .ZN(n5000) );
  OAI21_X1 U5612 ( .B1(n5002), .B2(n5001), .A(n5000), .ZN(n5008) );
  XOR2_X1 U5613 ( .A(REIP_REG_24__SCAN_IN), .B(keyinput_58), .Z(n5005) );
  XNOR2_X1 U5614 ( .A(REIP_REG_22__SCAN_IN), .B(keyinput_60), .ZN(n5004) );
  XNOR2_X1 U5615 ( .A(REIP_REG_23__SCAN_IN), .B(keyinput_59), .ZN(n5003) );
  NOR3_X1 U5616 ( .A1(n5005), .A2(n5004), .A3(n5003), .ZN(n5007) );
  XOR2_X1 U5617 ( .A(REIP_REG_21__SCAN_IN), .B(keyinput_61), .Z(n5006) );
  AOI21_X1 U5618 ( .B1(n5008), .B2(n5007), .A(n5006), .ZN(n5012) );
  XNOR2_X1 U5619 ( .A(keyinput_62), .B(REIP_REG_20__SCAN_IN), .ZN(n5011) );
  XOR2_X1 U5620 ( .A(REIP_REG_18__SCAN_IN), .B(keyinput_64), .Z(n5010) );
  XOR2_X1 U5621 ( .A(REIP_REG_19__SCAN_IN), .B(keyinput_63), .Z(n5009) );
  OAI211_X1 U5622 ( .C1(n5012), .C2(n5011), .A(n5010), .B(n5009), .ZN(n5020)
         );
  XOR2_X1 U5623 ( .A(BE_N_REG_2__SCAN_IN), .B(keyinput_68), .Z(n5019) );
  XOR2_X1 U5624 ( .A(REIP_REG_16__SCAN_IN), .B(keyinput_66), .Z(n5018) );
  XOR2_X1 U5625 ( .A(keyinput_65), .B(REIP_REG_17__SCAN_IN), .Z(n5016) );
  XOR2_X1 U5626 ( .A(keyinput_69), .B(BE_N_REG_1__SCAN_IN), .Z(n5015) );
  XOR2_X1 U5627 ( .A(keyinput_67), .B(BE_N_REG_3__SCAN_IN), .Z(n5014) );
  INV_X1 U5628 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n7361) );
  XNOR2_X1 U5629 ( .A(n7361), .B(keyinput_70), .ZN(n5013) );
  NOR4_X1 U5630 ( .A1(n5016), .A2(n5015), .A3(n5014), .A4(n5013), .ZN(n5017)
         );
  NAND4_X1 U5631 ( .A1(n5020), .A2(n5019), .A3(n5018), .A4(n5017), .ZN(n5024)
         );
  XOR2_X1 U5632 ( .A(ADDRESS_REG_29__SCAN_IN), .B(keyinput_71), .Z(n5023) );
  XOR2_X1 U5633 ( .A(keyinput_73), .B(ADDRESS_REG_27__SCAN_IN), .Z(n5022) );
  INV_X1 U5634 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n7334) );
  XNOR2_X1 U5635 ( .A(n7334), .B(keyinput_72), .ZN(n5021) );
  AOI211_X1 U5636 ( .C1(n5024), .C2(n5023), .A(n5022), .B(n5021), .ZN(n5028)
         );
  XNOR2_X1 U5637 ( .A(ADDRESS_REG_26__SCAN_IN), .B(keyinput_74), .ZN(n5027) );
  XOR2_X1 U5638 ( .A(ADDRESS_REG_24__SCAN_IN), .B(keyinput_76), .Z(n5026) );
  XNOR2_X1 U5639 ( .A(keyinput_75), .B(ADDRESS_REG_25__SCAN_IN), .ZN(n5025) );
  OAI211_X1 U5640 ( .C1(n5028), .C2(n5027), .A(n5026), .B(n5025), .ZN(n5035)
         );
  XOR2_X1 U5641 ( .A(ADDRESS_REG_23__SCAN_IN), .B(keyinput_77), .Z(n5034) );
  XOR2_X1 U5642 ( .A(ADDRESS_REG_19__SCAN_IN), .B(keyinput_81), .Z(n5032) );
  XNOR2_X1 U5643 ( .A(keyinput_80), .B(ADDRESS_REG_20__SCAN_IN), .ZN(n5031) );
  XNOR2_X1 U5644 ( .A(keyinput_78), .B(ADDRESS_REG_22__SCAN_IN), .ZN(n5030) );
  XNOR2_X1 U5645 ( .A(keyinput_79), .B(ADDRESS_REG_21__SCAN_IN), .ZN(n5029) );
  NAND4_X1 U5646 ( .A1(n5032), .A2(n5031), .A3(n5030), .A4(n5029), .ZN(n5033)
         );
  AOI21_X1 U5647 ( .B1(n5035), .B2(n5034), .A(n5033), .ZN(n5042) );
  XOR2_X1 U5648 ( .A(ADDRESS_REG_16__SCAN_IN), .B(keyinput_84), .Z(n5039) );
  XOR2_X1 U5649 ( .A(ADDRESS_REG_15__SCAN_IN), .B(keyinput_85), .Z(n5038) );
  XOR2_X1 U5650 ( .A(ADDRESS_REG_18__SCAN_IN), .B(keyinput_82), .Z(n5037) );
  XNOR2_X1 U5651 ( .A(keyinput_83), .B(ADDRESS_REG_17__SCAN_IN), .ZN(n5036) );
  NAND4_X1 U5652 ( .A1(n5039), .A2(n5038), .A3(n5037), .A4(n5036), .ZN(n5041)
         );
  XOR2_X1 U5653 ( .A(keyinput_86), .B(ADDRESS_REG_14__SCAN_IN), .Z(n5040) );
  OAI21_X1 U5654 ( .B1(n5042), .B2(n5041), .A(n5040), .ZN(n5065) );
  INV_X1 U5655 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n7299) );
  AOI22_X1 U5656 ( .A1(keyinput_93), .A2(n7299), .B1(n7297), .B2(keyinput_95), 
        .ZN(n5055) );
  AOI22_X1 U5657 ( .A1(keyinput_96), .A2(n7294), .B1(n7293), .B2(keyinput_97), 
        .ZN(n5054) );
  INV_X1 U5658 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n7301) );
  AOI22_X1 U5659 ( .A1(n7301), .A2(keyinput_91), .B1(ADDRESS_REG_12__SCAN_IN), 
        .B2(keyinput_88), .ZN(n5053) );
  OAI22_X1 U5660 ( .A1(n7294), .A2(keyinput_96), .B1(n7291), .B2(keyinput_98), 
        .ZN(n5044) );
  OAI22_X1 U5661 ( .A1(n7301), .A2(keyinput_91), .B1(n7297), .B2(keyinput_95), 
        .ZN(n5043) );
  NOR2_X1 U5662 ( .A1(n5044), .A2(n5043), .ZN(n5048) );
  OAI22_X1 U5663 ( .A1(ADDRESS_REG_13__SCAN_IN), .A2(keyinput_87), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(keyinput_88), .ZN(n5046) );
  OAI22_X1 U5664 ( .A1(n7299), .A2(keyinput_93), .B1(n7293), .B2(keyinput_97), 
        .ZN(n5045) );
  NOR2_X1 U5665 ( .A1(n5046), .A2(n5045), .ZN(n5047) );
  NAND2_X1 U5666 ( .A1(n5048), .A2(n5047), .ZN(n5049) );
  AOI21_X1 U5667 ( .B1(keyinput_87), .B2(ADDRESS_REG_13__SCAN_IN), .A(n5049), 
        .ZN(n5051) );
  NAND2_X1 U5668 ( .A1(n7291), .A2(keyinput_98), .ZN(n5050) );
  AND2_X1 U5669 ( .A1(n5051), .A2(n5050), .ZN(n5052) );
  NAND4_X1 U5670 ( .A1(n5055), .A2(n5054), .A3(n5053), .A4(n5052), .ZN(n5061)
         );
  XOR2_X1 U5671 ( .A(ADDRESS_REG_11__SCAN_IN), .B(keyinput_89), .Z(n5057) );
  XNOR2_X1 U5672 ( .A(keyinput_92), .B(ADDRESS_REG_8__SCAN_IN), .ZN(n5056) );
  NAND2_X1 U5673 ( .A1(n5057), .A2(n5056), .ZN(n5060) );
  XNOR2_X1 U5674 ( .A(ADDRESS_REG_6__SCAN_IN), .B(keyinput_94), .ZN(n5059) );
  XNOR2_X1 U5675 ( .A(ADDRESS_REG_10__SCAN_IN), .B(keyinput_90), .ZN(n5058) );
  NOR4_X1 U5676 ( .A1(n5061), .A2(n5060), .A3(n5059), .A4(n5058), .ZN(n5064)
         );
  XOR2_X1 U5677 ( .A(keyinput_100), .B(ADDRESS_REG_0__SCAN_IN), .Z(n5063) );
  XNOR2_X1 U5678 ( .A(ADDRESS_REG_1__SCAN_IN), .B(keyinput_99), .ZN(n5062) );
  AOI211_X1 U5679 ( .C1(n5065), .C2(n5064), .A(n5063), .B(n5062), .ZN(n5068)
         );
  XOR2_X1 U5680 ( .A(STATE_REG_2__SCAN_IN), .B(keyinput_101), .Z(n5067) );
  XOR2_X1 U5681 ( .A(STATE_REG_1__SCAN_IN), .B(keyinput_102), .Z(n5066) );
  NOR3_X1 U5682 ( .A1(n5068), .A2(n5067), .A3(n5066), .ZN(n5071) );
  XOR2_X1 U5683 ( .A(STATE_REG_0__SCAN_IN), .B(keyinput_103), .Z(n5070) );
  XNOR2_X1 U5684 ( .A(DATAWIDTH_REG_0__SCAN_IN), .B(keyinput_104), .ZN(n5069)
         );
  NOR3_X1 U5685 ( .A1(n5071), .A2(n5070), .A3(n5069), .ZN(n5073) );
  XOR2_X1 U5686 ( .A(keyinput_105), .B(DATAWIDTH_REG_1__SCAN_IN), .Z(n5072) );
  NOR2_X1 U5687 ( .A1(n5073), .A2(n5072), .ZN(n5079) );
  AOI22_X1 U5688 ( .A1(n7234), .A2(keyinput_109), .B1(keyinput_110), .B2(n7235), .ZN(n5074) );
  OAI221_X1 U5689 ( .B1(n7234), .B2(keyinput_109), .C1(n7235), .C2(
        keyinput_110), .A(n5074), .ZN(n5078) );
  INV_X1 U5690 ( .A(DATAWIDTH_REG_2__SCAN_IN), .ZN(n7231) );
  AOI22_X1 U5691 ( .A1(n7232), .A2(keyinput_107), .B1(keyinput_106), .B2(n7231), .ZN(n5075) );
  OAI221_X1 U5692 ( .B1(n7232), .B2(keyinput_107), .C1(n7231), .C2(
        keyinput_106), .A(n5075), .ZN(n5077) );
  XNOR2_X1 U5693 ( .A(DATAWIDTH_REG_4__SCAN_IN), .B(keyinput_108), .ZN(n5076)
         );
  NOR4_X1 U5694 ( .A1(n5079), .A2(n5078), .A3(n5077), .A4(n5076), .ZN(n5083)
         );
  INV_X1 U5695 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n7236) );
  XNOR2_X1 U5696 ( .A(n7236), .B(keyinput_111), .ZN(n5082) );
  XOR2_X1 U5697 ( .A(DATAWIDTH_REG_9__SCAN_IN), .B(keyinput_113), .Z(n5081) );
  XNOR2_X1 U5698 ( .A(keyinput_112), .B(DATAWIDTH_REG_8__SCAN_IN), .ZN(n5080)
         );
  OAI211_X1 U5699 ( .C1(n5083), .C2(n5082), .A(n5081), .B(n5080), .ZN(n5089)
         );
  XNOR2_X1 U5700 ( .A(keyinput_114), .B(DATAWIDTH_REG_10__SCAN_IN), .ZN(n5088)
         );
  XOR2_X1 U5701 ( .A(DATAWIDTH_REG_13__SCAN_IN), .B(keyinput_117), .Z(n5086)
         );
  XNOR2_X1 U5702 ( .A(keyinput_116), .B(DATAWIDTH_REG_12__SCAN_IN), .ZN(n5085)
         );
  XNOR2_X1 U5703 ( .A(keyinput_115), .B(DATAWIDTH_REG_11__SCAN_IN), .ZN(n5084)
         );
  NAND3_X1 U5704 ( .A1(n5086), .A2(n5085), .A3(n5084), .ZN(n5087) );
  AOI21_X1 U5705 ( .B1(n5089), .B2(n5088), .A(n5087), .ZN(n5092) );
  XOR2_X1 U5706 ( .A(keyinput_118), .B(DATAWIDTH_REG_14__SCAN_IN), .Z(n5091)
         );
  XOR2_X1 U5707 ( .A(keyinput_119), .B(DATAWIDTH_REG_15__SCAN_IN), .Z(n5090)
         );
  OAI21_X1 U5708 ( .B1(n5092), .B2(n5091), .A(n5090), .ZN(n5096) );
  XOR2_X1 U5709 ( .A(DATAWIDTH_REG_18__SCAN_IN), .B(keyinput_122), .Z(n5095)
         );
  XNOR2_X1 U5710 ( .A(keyinput_121), .B(DATAWIDTH_REG_17__SCAN_IN), .ZN(n5094)
         );
  XNOR2_X1 U5711 ( .A(keyinput_120), .B(DATAWIDTH_REG_16__SCAN_IN), .ZN(n5093)
         );
  NAND4_X1 U5712 ( .A1(n5096), .A2(n5095), .A3(n5094), .A4(n5093), .ZN(n5102)
         );
  XOR2_X1 U5713 ( .A(keyinput_123), .B(DATAWIDTH_REG_19__SCAN_IN), .Z(n5101)
         );
  XOR2_X1 U5714 ( .A(DATAWIDTH_REG_20__SCAN_IN), .B(keyinput_124), .Z(n5099)
         );
  XNOR2_X1 U5715 ( .A(DATAWIDTH_REG_22__SCAN_IN), .B(keyinput_126), .ZN(n5098)
         );
  XNOR2_X1 U5716 ( .A(DATAWIDTH_REG_21__SCAN_IN), .B(keyinput_125), .ZN(n5097)
         );
  NAND3_X1 U5717 ( .A1(n5099), .A2(n5098), .A3(n5097), .ZN(n5100) );
  AOI21_X1 U5718 ( .B1(n5102), .B2(n5101), .A(n5100), .ZN(n5104) );
  XNOR2_X1 U5719 ( .A(keyinput_255), .B(keyinput_127), .ZN(n5103) );
  XOR2_X1 U5720 ( .A(DATAWIDTH_REG_23__SCAN_IN), .B(keyinput_255), .Z(n5105)
         );
  NAND3_X1 U5721 ( .A1(n5106), .A2(n3737), .A3(n5105), .ZN(n5219) );
  BUF_X1 U5722 ( .A(n5108), .Z(n5109) );
  AOI21_X1 U5723 ( .B1(n5110), .B2(n5107), .A(n5109), .ZN(n6941) );
  NOR3_X1 U5724 ( .A1(n5114), .A2(n5113), .A3(n5112), .ZN(n5116) );
  OAI21_X1 U5725 ( .B1(n5117), .B2(n5116), .A(n5115), .ZN(n6674) );
  INV_X1 U5726 ( .A(n7711), .ZN(n7211) );
  NOR2_X1 U5727 ( .A1(n5119), .A2(n7211), .ZN(n5120) );
  NAND2_X1 U5728 ( .A1(n6674), .A2(n5120), .ZN(n5343) );
  NOR2_X1 U5729 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n7446) );
  NAND3_X1 U5730 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), 
        .A3(n7446), .ZN(n7220) );
  NAND2_X1 U5731 ( .A1(n5282), .A2(n5370), .ZN(n7719) );
  NAND2_X1 U5732 ( .A1(n5242), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5281)
         );
  INV_X1 U5733 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5280) );
  INV_X1 U5734 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5122) );
  INV_X1 U5735 ( .A(n6666), .ZN(n5124) );
  INV_X1 U5736 ( .A(EBX_REG_31__SCAN_IN), .ZN(n6882) );
  AND2_X4 U5737 ( .A1(n6280), .A2(n5591), .ZN(n6680) );
  NAND2_X1 U5738 ( .A1(n7442), .A2(n7726), .ZN(n5209) );
  NAND2_X1 U5739 ( .A1(n6680), .A2(n5209), .ZN(n5126) );
  NAND2_X1 U5740 ( .A1(n5298), .A2(n3746), .ZN(n5130) );
  INV_X4 U5741 ( .A(n3746), .ZN(n6586) );
  OAI211_X1 U5742 ( .C1(INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n6587), .A(n5130), 
        .B(n5129), .ZN(n5134) );
  INV_X1 U5743 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5131) );
  OR2_X1 U5744 ( .A1(n5322), .A2(n5131), .ZN(n5133) );
  NAND2_X1 U5745 ( .A1(n3746), .A2(n5131), .ZN(n5132) );
  NAND2_X1 U5746 ( .A1(n5133), .A2(n5132), .ZN(n5390) );
  XNOR2_X1 U5747 ( .A(n5134), .B(n5390), .ZN(n5352) );
  AOI21_X1 U5748 ( .B1(n5352), .B2(n6680), .A(n5134), .ZN(n5533) );
  MUX2_X1 U5749 ( .A(n5327), .B(n6586), .S(EBX_REG_2__SCAN_IN), .Z(n5136) );
  OAI21_X1 U5750 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6587), .A(n5136), 
        .ZN(n5535) );
  INV_X1 U5751 ( .A(n5535), .ZN(n5137) );
  NAND2_X1 U5752 ( .A1(n5533), .A2(n5137), .ZN(n5539) );
  INV_X1 U5753 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6856) );
  NAND2_X1 U5754 ( .A1(n5320), .A2(n6856), .ZN(n5141) );
  NAND2_X1 U5755 ( .A1(n5322), .A2(n5581), .ZN(n5139) );
  NAND2_X1 U5756 ( .A1(n6680), .A2(n6856), .ZN(n5138) );
  NAND3_X1 U5757 ( .A1(n5139), .A2(n6586), .A3(n5138), .ZN(n5140) );
  AND2_X1 U5758 ( .A1(n5141), .A2(n5140), .ZN(n5538) );
  MUX2_X1 U5759 ( .A(n5327), .B(n6586), .S(EBX_REG_4__SCAN_IN), .Z(n5143) );
  OAI21_X1 U5760 ( .B1(INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n6587), .A(n5143), 
        .ZN(n5499) );
  NAND2_X1 U5761 ( .A1(n5322), .A2(n7460), .ZN(n5145) );
  INV_X1 U5762 ( .A(EBX_REG_5__SCAN_IN), .ZN(n7565) );
  NAND2_X1 U5763 ( .A1(n6680), .A2(n7565), .ZN(n5144) );
  NAND3_X1 U5764 ( .A1(n5145), .A2(n6586), .A3(n5144), .ZN(n5146) );
  OAI21_X1 U5765 ( .B1(n5332), .B2(EBX_REG_5__SCAN_IN), .A(n5146), .ZN(n5492)
         );
  MUX2_X1 U5766 ( .A(n5327), .B(n6586), .S(EBX_REG_6__SCAN_IN), .Z(n5147) );
  OAI21_X1 U5767 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n6587), .A(n5147), 
        .ZN(n5652) );
  INV_X1 U5768 ( .A(EBX_REG_7__SCAN_IN), .ZN(n7586) );
  NAND2_X1 U5769 ( .A1(n5320), .A2(n7586), .ZN(n5153) );
  NAND2_X1 U5770 ( .A1(n5322), .A2(n5149), .ZN(n5151) );
  NAND2_X1 U5771 ( .A1(n6680), .A2(n7586), .ZN(n5150) );
  NAND3_X1 U5772 ( .A1(n5151), .A2(n6586), .A3(n5150), .ZN(n5152) );
  MUX2_X1 U5773 ( .A(n5327), .B(n6586), .S(EBX_REG_8__SCAN_IN), .Z(n5154) );
  OAI21_X1 U5774 ( .B1(n6587), .B2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n5154), 
        .ZN(n5155) );
  INV_X1 U5775 ( .A(n5155), .ZN(n6008) );
  INV_X1 U5776 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n7482) );
  NAND2_X1 U5777 ( .A1(n5322), .A2(n7482), .ZN(n5157) );
  INV_X1 U5778 ( .A(EBX_REG_9__SCAN_IN), .ZN(n7611) );
  NAND2_X1 U5779 ( .A1(n6680), .A2(n7611), .ZN(n5156) );
  NAND3_X1 U5780 ( .A1(n5157), .A2(n6586), .A3(n5156), .ZN(n5158) );
  OAI21_X1 U5781 ( .B1(n5332), .B2(EBX_REG_9__SCAN_IN), .A(n5158), .ZN(n6232)
         );
  NAND2_X1 U5782 ( .A1(n6007), .A2(n6232), .ZN(n6231) );
  MUX2_X1 U5783 ( .A(n5327), .B(n6586), .S(EBX_REG_10__SCAN_IN), .Z(n5159) );
  OAI21_X1 U5784 ( .B1(n6587), .B2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n5159), 
        .ZN(n6266) );
  INV_X1 U5785 ( .A(EBX_REG_11__SCAN_IN), .ZN(n7635) );
  NAND2_X1 U5786 ( .A1(n5320), .A2(n7635), .ZN(n5164) );
  NAND2_X1 U5787 ( .A1(n5322), .A2(n7503), .ZN(n5162) );
  NAND2_X1 U5788 ( .A1(n6680), .A2(n7635), .ZN(n5161) );
  NAND3_X1 U5789 ( .A1(n5162), .A2(n6586), .A3(n5161), .ZN(n5163) );
  INV_X1 U5790 ( .A(n5327), .ZN(n5193) );
  INV_X1 U5791 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6453) );
  NAND2_X1 U5792 ( .A1(n5193), .A2(n6453), .ZN(n5167) );
  NAND2_X1 U5793 ( .A1(n6680), .A2(n6453), .ZN(n5165) );
  OAI211_X1 U5794 ( .C1(n3746), .C2(n6506), .A(n5165), .B(n5322), .ZN(n5166)
         );
  NAND2_X1 U5795 ( .A1(n5167), .A2(n5166), .ZN(n6450) );
  NAND2_X1 U5796 ( .A1(n5322), .A2(n5168), .ZN(n5170) );
  INV_X1 U5797 ( .A(EBX_REG_13__SCAN_IN), .ZN(n7650) );
  NAND2_X1 U5798 ( .A1(n6680), .A2(n7650), .ZN(n5169) );
  NAND3_X1 U5799 ( .A1(n5170), .A2(n6586), .A3(n5169), .ZN(n5171) );
  OAI21_X1 U5800 ( .B1(n5332), .B2(EBX_REG_13__SCAN_IN), .A(n5171), .ZN(n6482)
         );
  NAND2_X1 U5801 ( .A1(n6483), .A2(n6482), .ZN(n6516) );
  MUX2_X1 U5802 ( .A(n5327), .B(n6586), .S(EBX_REG_14__SCAN_IN), .Z(n5173) );
  INV_X1 U5803 ( .A(n6587), .ZN(n5416) );
  NAND2_X1 U5804 ( .A1(n5416), .A2(n6514), .ZN(n5172) );
  NAND2_X1 U5805 ( .A1(n5173), .A2(n5172), .ZN(n6517) );
  NOR2_X2 U5806 ( .A1(n6516), .A2(n6517), .ZN(n6518) );
  INV_X1 U5807 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5174) );
  NAND2_X1 U5808 ( .A1(n5320), .A2(n5174), .ZN(n5178) );
  NAND2_X1 U5809 ( .A1(n5322), .A2(n7514), .ZN(n5176) );
  NAND2_X1 U5810 ( .A1(n6680), .A2(n5174), .ZN(n5175) );
  NAND3_X1 U5811 ( .A1(n5176), .A2(n6586), .A3(n5175), .ZN(n5177) );
  MUX2_X1 U5812 ( .A(n5327), .B(n6586), .S(EBX_REG_16__SCAN_IN), .Z(n5181) );
  OR2_X1 U5813 ( .A1(n6587), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5180)
         );
  INV_X1 U5814 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n7539) );
  NAND2_X1 U5815 ( .A1(n5322), .A2(n7539), .ZN(n5183) );
  INV_X1 U5816 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6909) );
  NAND2_X1 U5817 ( .A1(n6680), .A2(n6909), .ZN(n5182) );
  NAND3_X1 U5818 ( .A1(n5183), .A2(n6586), .A3(n5182), .ZN(n5184) );
  OAI21_X1 U5819 ( .B1(n5332), .B2(EBX_REG_17__SCAN_IN), .A(n5184), .ZN(n6796)
         );
  MUX2_X1 U5820 ( .A(n5327), .B(n6586), .S(EBX_REG_18__SCAN_IN), .Z(n5185) );
  OAI21_X1 U5821 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n6587), .A(n5185), 
        .ZN(n6905) );
  INV_X1 U5822 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5187) );
  NAND2_X1 U5823 ( .A1(n5320), .A2(n5187), .ZN(n5191) );
  NAND2_X1 U5824 ( .A1(n6586), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U5825 ( .A1(n5322), .A2(n5186), .ZN(n5189) );
  NAND2_X1 U5826 ( .A1(n6680), .A2(n5187), .ZN(n5188) );
  NAND2_X1 U5827 ( .A1(n5189), .A2(n5188), .ZN(n5190) );
  INV_X1 U5828 ( .A(EBX_REG_20__SCAN_IN), .ZN(n7368) );
  NAND2_X1 U5829 ( .A1(n5193), .A2(n7368), .ZN(n5197) );
  NAND2_X1 U5830 ( .A1(n6680), .A2(n7368), .ZN(n5195) );
  NAND2_X1 U5831 ( .A1(n6586), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5194) );
  NAND3_X1 U5832 ( .A1(n5195), .A2(n5322), .A3(n5194), .ZN(n5196) );
  AND2_X1 U5833 ( .A1(n5197), .A2(n5196), .ZN(n7143) );
  AND2_X2 U5834 ( .A1(n6898), .A2(n7143), .ZN(n7145) );
  NAND2_X1 U5835 ( .A1(n6586), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U5836 ( .A1(n5322), .A2(n5198), .ZN(n5200) );
  NAND2_X1 U5837 ( .A1(n6680), .A2(n6895), .ZN(n5199) );
  NAND2_X1 U5838 ( .A1(n5200), .A2(n5199), .ZN(n5201) );
  OAI21_X1 U5839 ( .B1(n5332), .B2(EBX_REG_21__SCAN_IN), .A(n5201), .ZN(n5202)
         );
  NAND2_X1 U5840 ( .A1(n7145), .A2(n5202), .ZN(n5307) );
  OAI21_X1 U5841 ( .B1(n7145), .B2(n5202), .A(n5307), .ZN(n7139) );
  INV_X1 U5842 ( .A(REIP_REG_17__SCAN_IN), .ZN(n7311) );
  NAND2_X1 U5843 ( .A1(n5203), .A2(n7736), .ZN(n7435) );
  AND2_X1 U5844 ( .A1(n6280), .A2(n6682), .ZN(n5204) );
  NOR2_X1 U5845 ( .A1(n6680), .A2(n5204), .ZN(n5205) );
  INV_X1 U5846 ( .A(n6808), .ZN(n6876) );
  NAND3_X1 U5847 ( .A1(REIP_REG_6__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_8__SCAN_IN), .ZN(n7620) );
  INV_X1 U5848 ( .A(REIP_REG_11__SCAN_IN), .ZN(n7640) );
  INV_X1 U5849 ( .A(REIP_REG_10__SCAN_IN), .ZN(n7631) );
  INV_X1 U5850 ( .A(REIP_REG_9__SCAN_IN), .ZN(n7619) );
  NOR4_X1 U5851 ( .A1(n7620), .A2(n7640), .A3(n7631), .A4(n7619), .ZN(n6846)
         );
  NAND4_X1 U5852 ( .A1(n6846), .A2(REIP_REG_13__SCAN_IN), .A3(
        REIP_REG_12__SCAN_IN), .A4(REIP_REG_14__SCAN_IN), .ZN(n6809) );
  INV_X1 U5853 ( .A(REIP_REG_15__SCAN_IN), .ZN(n7308) );
  NAND3_X1 U5854 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .A3(
        REIP_REG_3__SCAN_IN), .ZN(n6294) );
  INV_X1 U5855 ( .A(REIP_REG_4__SCAN_IN), .ZN(n7292) );
  NOR2_X1 U5856 ( .A1(n6294), .A2(n7292), .ZN(n6806) );
  NAND2_X1 U5857 ( .A1(n6806), .A2(REIP_REG_5__SCAN_IN), .ZN(n6842) );
  NOR4_X1 U5858 ( .A1(n6809), .A2(n7525), .A3(n7308), .A4(n6842), .ZN(n5206)
         );
  NAND2_X1 U5859 ( .A1(n6876), .A2(n5206), .ZN(n6791) );
  NOR2_X1 U5860 ( .A1(n7311), .A2(n6791), .ZN(n7672) );
  NAND2_X1 U5861 ( .A1(REIP_REG_18__SCAN_IN), .A2(n7672), .ZN(n7674) );
  NOR2_X1 U5862 ( .A1(n7673), .A2(n7674), .ZN(n7691) );
  NAND3_X1 U5863 ( .A1(n7691), .A2(REIP_REG_20__SCAN_IN), .A3(n7317), .ZN(
        n6782) );
  INV_X1 U5864 ( .A(n6871), .ZN(n6843) );
  NAND2_X1 U5865 ( .A1(n5206), .A2(REIP_REG_17__SCAN_IN), .ZN(n6613) );
  NOR2_X1 U5866 ( .A1(n6843), .A2(n6613), .ZN(n6790) );
  NOR3_X1 U5867 ( .A1(n7315), .A2(n7671), .A3(n7673), .ZN(n5207) );
  NAND2_X1 U5868 ( .A1(n6790), .A2(n5207), .ZN(n5208) );
  NAND2_X1 U5869 ( .A1(n6808), .A2(n6871), .ZN(n7598) );
  AND2_X1 U5870 ( .A1(n5208), .A2(n7598), .ZN(n7692) );
  NOR2_X1 U5871 ( .A1(n7435), .A2(n5209), .ZN(n7213) );
  OR2_X1 U5872 ( .A1(n7443), .A2(n7213), .ZN(n6686) );
  NAND3_X1 U5873 ( .A1(n6280), .A2(n6882), .A3(n5209), .ZN(n5210) );
  AND2_X1 U5874 ( .A1(n6686), .A2(n5210), .ZN(n5211) );
  AND2_X1 U5875 ( .A1(n6666), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5212) );
  AND2_X2 U5876 ( .A1(n6871), .A2(n5212), .ZN(n7682) );
  AOI22_X1 U5877 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n7688), .B1(n7682), 
        .B2(n7003), .ZN(n5213) );
  OAI21_X1 U5878 ( .B1(n6895), .B2(n7686), .A(n5213), .ZN(n5214) );
  AOI21_X1 U5879 ( .B1(n7692), .B2(REIP_REG_21__SCAN_IN), .A(n5214), .ZN(n5215) );
  OAI211_X1 U5880 ( .C1(n7693), .C2(n7139), .A(n6782), .B(n5215), .ZN(n5216)
         );
  AOI21_X1 U5881 ( .B1(n6941), .B2(n7696), .A(n5216), .ZN(n5217) );
  XNOR2_X1 U5882 ( .A(n5219), .B(n5218), .ZN(U2806) );
  INV_X1 U5883 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n7076) );
  NAND2_X1 U5884 ( .A1(n7076), .A2(n5321), .ZN(n7072) );
  NOR2_X1 U5885 ( .A1(n7072), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5220)
         );
  INV_X1 U5886 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6581) );
  XNOR2_X1 U5887 ( .A(n4252), .B(n6581), .ZN(n5221) );
  XNOR2_X1 U5888 ( .A(n5222), .B(n5221), .ZN(n6604) );
  INV_X1 U5889 ( .A(n6604), .ZN(n5223) );
  NAND2_X1 U5890 ( .A1(n5223), .A2(n7422), .ZN(n5253) );
  AOI22_X1 U5891 ( .A1(n3921), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5227) );
  AOI22_X1 U5892 ( .A1(n4552), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5226) );
  AOI22_X1 U5893 ( .A1(n4010), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3655), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n5225) );
  AOI22_X1 U5894 ( .A1(n3660), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5224) );
  NAND4_X1 U5895 ( .A1(n5227), .A2(n5226), .A3(n5225), .A4(n5224), .ZN(n5233)
         );
  AOI22_X1 U5896 ( .A1(n3653), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3651), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5231) );
  AOI22_X1 U5897 ( .A1(n3644), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n5261), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5230) );
  AOI22_X1 U5898 ( .A1(n5258), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5229) );
  AOI22_X1 U5899 ( .A1(n5259), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4505), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5228) );
  NAND4_X1 U5900 ( .A1(n5231), .A2(n5230), .A3(n5229), .A4(n5228), .ZN(n5232)
         );
  NOR2_X1 U5901 ( .A1(n5233), .A2(n5232), .ZN(n5274) );
  NAND2_X1 U5902 ( .A1(n5235), .A2(n5234), .ZN(n5273) );
  XOR2_X1 U5903 ( .A(n5274), .B(n5273), .Z(n5237) );
  NAND2_X1 U5904 ( .A1(n5237), .A2(n5236), .ZN(n5240) );
  INV_X1 U5905 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5241) );
  AOI21_X1 U5906 ( .B1(n5241), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n5238) );
  AOI21_X1 U5907 ( .B1(n6660), .B2(EAX_REG_29__SCAN_IN), .A(n5238), .ZN(n5239)
         );
  NAND2_X1 U5908 ( .A1(n5240), .A2(n5239), .ZN(n5244) );
  XNOR2_X1 U5909 ( .A(n5242), .B(n5241), .ZN(n6696) );
  NAND2_X1 U5910 ( .A1(n6696), .A2(n5282), .ZN(n5243) );
  NAND2_X1 U5911 ( .A1(n5244), .A2(n5243), .ZN(n5247) );
  OR2_X1 U5912 ( .A1(n5247), .A2(n5245), .ZN(n5246) );
  NOR2_X2 U5913 ( .A1(n6709), .A2(n5285), .ZN(n5288) );
  INV_X1 U5914 ( .A(n6696), .ZN(n5250) );
  NOR2_X1 U5915 ( .A1(n7524), .A2(n7333), .ZN(n6601) );
  AOI21_X1 U5916 ( .B1(n7415), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n6601), 
        .ZN(n5249) );
  OAI21_X1 U5917 ( .B1(n7425), .B2(n5250), .A(n5249), .ZN(n5251) );
  AOI21_X1 U5918 ( .B1(n6707), .B2(n7421), .A(n5251), .ZN(n5252) );
  NAND2_X1 U5919 ( .A1(n5253), .A2(n5252), .ZN(U2957) );
  NAND2_X1 U5920 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6578) );
  AND2_X1 U5921 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6598) );
  NAND2_X1 U5922 ( .A1(n6598), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n7063) );
  OAI21_X1 U5923 ( .B1(n6578), .B2(n7063), .A(n4252), .ZN(n5255) );
  NAND2_X1 U5924 ( .A1(n6571), .A2(n6581), .ZN(n5256) );
  NAND2_X1 U5925 ( .A1(n7059), .A2(n7422), .ZN(n5294) );
  AOI22_X1 U5926 ( .A1(n5259), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5258), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n5265) );
  AOI22_X1 U5927 ( .A1(n4352), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5264) );
  AOI22_X1 U5928 ( .A1(n3622), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4488), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5263) );
  AOI22_X1 U5929 ( .A1(n5261), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5260), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5262) );
  NAND4_X1 U5930 ( .A1(n5265), .A2(n5264), .A3(n5263), .A4(n5262), .ZN(n5272)
         );
  AOI22_X1 U5931 ( .A1(n3627), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5270) );
  AOI22_X1 U5932 ( .A1(n3628), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5269) );
  AOI22_X1 U5933 ( .A1(n4552), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5268) );
  AOI22_X1 U5934 ( .A1(n3657), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5769), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5267) );
  NAND4_X1 U5935 ( .A1(n5270), .A2(n5269), .A3(n5268), .A4(n5267), .ZN(n5271)
         );
  NOR2_X1 U5936 ( .A1(n5272), .A2(n5271), .ZN(n5276) );
  NOR2_X1 U5937 ( .A1(n5274), .A2(n5273), .ZN(n5275) );
  XOR2_X1 U5938 ( .A(n5276), .B(n5275), .Z(n5279) );
  AOI22_X1 U5939 ( .A1(n6660), .A2(EAX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n5838), .ZN(n5277) );
  OAI21_X1 U5940 ( .B1(n5279), .B2(n5278), .A(n5277), .ZN(n5283) );
  XNOR2_X1 U5941 ( .A(n5281), .B(n5280), .ZN(n6621) );
  MUX2_X1 U5942 ( .A(n5283), .B(n6621), .S(n5282), .Z(n5289) );
  INV_X1 U5943 ( .A(n6725), .ZN(n6736) );
  INV_X1 U5944 ( .A(n5289), .ZN(n5284) );
  NOR2_X1 U5945 ( .A1(n5285), .A2(n5284), .ZN(n5286) );
  NAND2_X1 U5946 ( .A1(n6724), .A2(n5286), .ZN(n5287) );
  OAI21_X2 U5947 ( .B1(n5289), .B2(n5288), .A(n6663), .ZN(n6922) );
  INV_X1 U5948 ( .A(REIP_REG_30__SCAN_IN), .ZN(n7337) );
  NOR2_X1 U5949 ( .A1(n7524), .A2(n7337), .ZN(n7065) );
  NOR2_X1 U5950 ( .A1(n7425), .A2(n6621), .ZN(n5290) );
  AOI211_X1 U5951 ( .C1(n7415), .C2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n7065), 
        .B(n5290), .ZN(n5291) );
  INV_X1 U5952 ( .A(n5292), .ZN(n5293) );
  NAND2_X1 U5953 ( .A1(n5294), .A2(n5293), .ZN(U2956) );
  INV_X1 U5954 ( .A(n6707), .ZN(n6640) );
  NAND2_X1 U5955 ( .A1(n6064), .A2(n6280), .ZN(n5296) );
  OAI22_X1 U5956 ( .A1(n5295), .A2(n5296), .B1(n7443), .B2(n6064), .ZN(n5419)
         );
  OR2_X1 U5957 ( .A1(n5761), .A2(n5419), .ZN(n5297) );
  NAND2_X1 U5958 ( .A1(n5297), .A2(n5119), .ZN(n5396) );
  NOR2_X1 U5959 ( .A1(n7166), .A2(n5298), .ZN(n5299) );
  NAND2_X1 U5960 ( .A1(n5396), .A2(n5299), .ZN(n6678) );
  INV_X1 U5961 ( .A(n3933), .ZN(n6670) );
  NAND4_X1 U5962 ( .A1(n6670), .A2(n5452), .A3(n7711), .A4(n3937), .ZN(n6059)
         );
  INV_X1 U5963 ( .A(n6059), .ZN(n5302) );
  INV_X1 U5964 ( .A(n5322), .ZN(n5301) );
  AND2_X1 U5965 ( .A1(n6067), .A2(n5591), .ZN(n5300) );
  NAND4_X1 U5966 ( .A1(n5302), .A2(n3638), .A3(n5301), .A4(n5300), .ZN(n5303)
         );
  NAND2_X2 U5967 ( .A1(n7369), .A2(n3933), .ZN(n6919) );
  INV_X1 U5968 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6531) );
  INV_X1 U5969 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6894) );
  NAND2_X1 U5970 ( .A1(n6680), .A2(n6894), .ZN(n5305) );
  OAI211_X1 U5971 ( .C1(n3746), .C2(n6531), .A(n5305), .B(n5322), .ZN(n5306)
         );
  OAI21_X1 U5972 ( .B1(n5327), .B2(EBX_REG_22__SCAN_IN), .A(n5306), .ZN(n6772)
         );
  INV_X1 U5973 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6891) );
  NAND2_X1 U5974 ( .A1(n5320), .A2(n6891), .ZN(n5311) );
  NAND2_X1 U5975 ( .A1(n5322), .A2(n7110), .ZN(n5309) );
  NAND2_X1 U5976 ( .A1(n6680), .A2(n6891), .ZN(n5308) );
  NAND3_X1 U5977 ( .A1(n5309), .A2(n6586), .A3(n5308), .ZN(n5310) );
  AND2_X1 U5978 ( .A1(n5311), .A2(n5310), .ZN(n6756) );
  INV_X1 U5979 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5312) );
  NAND2_X1 U5980 ( .A1(n6680), .A2(n5312), .ZN(n5313) );
  OAI211_X1 U5981 ( .C1(n3746), .C2(n6558), .A(n5313), .B(n5322), .ZN(n5314)
         );
  OAI21_X1 U5982 ( .B1(n5327), .B2(EBX_REG_24__SCAN_IN), .A(n5314), .ZN(n6539)
         );
  OAI21_X1 U5983 ( .B1(n3746), .B2(n7103), .A(n5322), .ZN(n5315) );
  OAI21_X1 U5984 ( .B1(EBX_REG_25__SCAN_IN), .B2(n5298), .A(n5315), .ZN(n5317)
         );
  INV_X1 U5985 ( .A(EBX_REG_25__SCAN_IN), .ZN(n6887) );
  NAND2_X1 U5986 ( .A1(n5320), .A2(n6887), .ZN(n5316) );
  NAND2_X1 U5987 ( .A1(n5317), .A2(n5316), .ZN(n6734) );
  MUX2_X1 U5988 ( .A(n5327), .B(n6586), .S(EBX_REG_26__SCAN_IN), .Z(n5318) );
  OAI21_X1 U5989 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n6587), .A(n5318), 
        .ZN(n6721) );
  INV_X1 U5990 ( .A(EBX_REG_27__SCAN_IN), .ZN(n6713) );
  NAND2_X1 U5991 ( .A1(n5320), .A2(n6713), .ZN(n5326) );
  NAND2_X1 U5992 ( .A1(n5322), .A2(n5321), .ZN(n5324) );
  NAND2_X1 U5993 ( .A1(n6680), .A2(n6713), .ZN(n5323) );
  NAND3_X1 U5994 ( .A1(n5324), .A2(n6586), .A3(n5323), .ZN(n5325) );
  AND2_X1 U5995 ( .A1(n5326), .A2(n5325), .ZN(n6712) );
  MUX2_X1 U5996 ( .A(n5327), .B(n6586), .S(EBX_REG_28__SCAN_IN), .Z(n5329) );
  OR2_X1 U5997 ( .A1(n6587), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5328)
         );
  AND2_X1 U5998 ( .A1(n5329), .A2(n5328), .ZN(n6629) );
  OR2_X1 U5999 ( .A1(n6587), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5331)
         );
  INV_X1 U6000 ( .A(EBX_REG_29__SCAN_IN), .ZN(n6699) );
  NAND2_X1 U6001 ( .A1(n6680), .A2(n6699), .ZN(n5330) );
  NAND2_X1 U6002 ( .A1(n5331), .A2(n5330), .ZN(n6605) );
  OAI22_X1 U6003 ( .A1(n6605), .A2(n3746), .B1(n5332), .B2(EBX_REG_29__SCAN_IN), .ZN(n5334) );
  OR2_X1 U6004 ( .A1(n5333), .A2(n5334), .ZN(n5335) );
  NAND2_X1 U6005 ( .A1(n6607), .A2(n5335), .ZN(n6705) );
  INV_X1 U6006 ( .A(n5790), .ZN(n6679) );
  NAND2_X1 U6007 ( .A1(n6674), .A2(n3945), .ZN(n5339) );
  AOI22_X1 U6008 ( .A1(n6679), .A2(n3946), .B1(n5111), .B2(n5339), .ZN(n6684)
         );
  AND2_X1 U6009 ( .A1(n6684), .A2(n7711), .ZN(n5342) );
  INV_X1 U6010 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n7724) );
  NAND3_X1 U6011 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n7446), .A3(n7724), .ZN(
        n5340) );
  OAI21_X1 U6012 ( .B1(n5342), .B2(n5341), .A(n5340), .ZN(U2790) );
  INV_X1 U6013 ( .A(n5343), .ZN(n5344) );
  OAI211_X1 U6014 ( .C1(n5344), .C2(n7748), .A(n5590), .B(n7428), .ZN(U2788)
         );
  XNOR2_X1 U6015 ( .A(n5346), .B(n5345), .ZN(n5392) );
  OAI21_X1 U6016 ( .B1(n5347), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n5394), 
        .ZN(n7551) );
  NAND2_X1 U6017 ( .A1(n7544), .A2(REIP_REG_0__SCAN_IN), .ZN(n7552) );
  OAI21_X1 U6018 ( .B1(n7415), .B2(n5348), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5349) );
  OAI211_X1 U6019 ( .C1(n7551), .C2(n7701), .A(n7552), .B(n5349), .ZN(n5350)
         );
  AOI21_X1 U6020 ( .B1(n7421), .B2(n5392), .A(n5350), .ZN(n5351) );
  INV_X1 U6021 ( .A(n5351), .ZN(U2986) );
  XNOR2_X1 U6022 ( .A(n5352), .B(n6680), .ZN(n5427) );
  INV_X1 U6023 ( .A(n5427), .ZN(n5356) );
  INV_X1 U6024 ( .A(EBX_REG_1__SCAN_IN), .ZN(n6285) );
  OAI21_X1 U6025 ( .B1(n5355), .B2(n5354), .A(n5353), .ZN(n7370) );
  OAI222_X1 U6026 ( .A1(n5356), .A2(n6917), .B1(n6285), .B2(n7369), .C1(n7370), 
        .C2(n6919), .ZN(U2858) );
  XNOR2_X1 U6027 ( .A(n5358), .B(n5581), .ZN(n5359) );
  XNOR2_X1 U6028 ( .A(n5357), .B(n5359), .ZN(n5984) );
  OAI21_X1 U6029 ( .B1(n5360), .B2(n5362), .A(n5361), .ZN(n6089) );
  INV_X1 U6030 ( .A(n6089), .ZN(n6867) );
  NAND2_X1 U6031 ( .A1(n7544), .A2(REIP_REG_3__SCAN_IN), .ZN(n5978) );
  NAND2_X1 U6032 ( .A1(n7415), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5363)
         );
  OAI211_X1 U6033 ( .C1(n7425), .C2(n6857), .A(n5978), .B(n5363), .ZN(n5364)
         );
  AOI21_X1 U6034 ( .B1(n6867), .B2(n7421), .A(n5364), .ZN(n5365) );
  OAI21_X1 U6035 ( .B1(n5984), .B2(n7701), .A(n5365), .ZN(U2983) );
  INV_X1 U6036 ( .A(EAX_REG_21__SCAN_IN), .ZN(n5372) );
  OR2_X1 U6037 ( .A1(n5367), .A2(n7443), .ZN(n7212) );
  OR2_X1 U6038 ( .A1(n5119), .A2(n3956), .ZN(n7188) );
  NAND2_X1 U6039 ( .A1(n7255), .A2(n6280), .ZN(n6244) );
  NAND2_X1 U6040 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5370), .ZN(n7210) );
  INV_X2 U6041 ( .A(n7210), .ZN(n7284) );
  NOR2_X4 U6042 ( .A1(n7284), .A2(n7255), .ZN(n7252) );
  AOI22_X1 U6043 ( .A1(n7284), .A2(UWORD_REG_5__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n5371) );
  OAI21_X1 U6044 ( .B1(n5372), .B2(n6244), .A(n5371), .ZN(U2902) );
  INV_X1 U6045 ( .A(EAX_REG_22__SCAN_IN), .ZN(n5374) );
  AOI22_X1 U6046 ( .A1(n7284), .A2(UWORD_REG_6__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n5373) );
  OAI21_X1 U6047 ( .B1(n5374), .B2(n6244), .A(n5373), .ZN(U2901) );
  INV_X1 U6048 ( .A(EAX_REG_25__SCAN_IN), .ZN(n5376) );
  AOI22_X1 U6049 ( .A1(n7284), .A2(UWORD_REG_9__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n5375) );
  OAI21_X1 U6050 ( .B1(n5376), .B2(n6244), .A(n5375), .ZN(U2898) );
  AOI22_X1 U6051 ( .A1(n7284), .A2(UWORD_REG_4__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n5377) );
  OAI21_X1 U6052 ( .B1(n4547), .B2(n6244), .A(n5377), .ZN(U2903) );
  INV_X1 U6053 ( .A(EAX_REG_28__SCAN_IN), .ZN(n5379) );
  AOI22_X1 U6054 ( .A1(n7284), .A2(UWORD_REG_12__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n5378) );
  OAI21_X1 U6055 ( .B1(n5379), .B2(n6244), .A(n5378), .ZN(U2895) );
  INV_X1 U6056 ( .A(EAX_REG_27__SCAN_IN), .ZN(n5381) );
  AOI22_X1 U6057 ( .A1(n7284), .A2(UWORD_REG_11__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n5380) );
  OAI21_X1 U6058 ( .B1(n5381), .B2(n6244), .A(n5380), .ZN(U2896) );
  INV_X1 U6059 ( .A(EAX_REG_26__SCAN_IN), .ZN(n5383) );
  AOI22_X1 U6060 ( .A1(n7284), .A2(UWORD_REG_10__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n5382) );
  OAI21_X1 U6061 ( .B1(n5383), .B2(n6244), .A(n5382), .ZN(U2897) );
  INV_X1 U6062 ( .A(EAX_REG_23__SCAN_IN), .ZN(n5385) );
  AOI22_X1 U6063 ( .A1(n7284), .A2(UWORD_REG_7__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n5384) );
  OAI21_X1 U6064 ( .B1(n5385), .B2(n6244), .A(n5384), .ZN(U2900) );
  INV_X1 U6065 ( .A(EAX_REG_29__SCAN_IN), .ZN(n5387) );
  AOI22_X1 U6066 ( .A1(n7284), .A2(UWORD_REG_13__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n5386) );
  OAI21_X1 U6067 ( .B1(n5387), .B2(n6244), .A(n5386), .ZN(U2894) );
  INV_X1 U6068 ( .A(EAX_REG_24__SCAN_IN), .ZN(n5389) );
  AOI22_X1 U6069 ( .A1(n7284), .A2(UWORD_REG_8__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n5388) );
  OAI21_X1 U6070 ( .B1(n5389), .B2(n6244), .A(n5388), .ZN(U2899) );
  INV_X1 U6071 ( .A(n5390), .ZN(n5391) );
  OAI21_X1 U6072 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n6587), .A(n5391), 
        .ZN(n7554) );
  INV_X1 U6073 ( .A(n5392), .ZN(n6312) );
  OAI222_X1 U6074 ( .A1(n7554), .A2(n6917), .B1(n7369), .B2(n5131), .C1(n6919), 
        .C2(n6312), .ZN(U2859) );
  XOR2_X1 U6075 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .B(n5394), .Z(n5395) );
  XNOR2_X1 U6076 ( .A(n5393), .B(n5395), .ZN(n7371) );
  INV_X1 U6077 ( .A(n7371), .ZN(n5431) );
  OR3_X1 U6078 ( .A1(n5790), .A2(n3956), .A3(n7166), .ZN(n5397) );
  NAND2_X1 U6079 ( .A1(n5591), .A2(n7435), .ZN(n5398) );
  AND2_X1 U6080 ( .A1(n7442), .A2(n6674), .ZN(n5784) );
  AND3_X1 U6081 ( .A1(n5398), .A2(n3983), .A3(n5784), .ZN(n5399) );
  OAI21_X1 U6082 ( .B1(n5591), .B2(n6682), .A(n7442), .ZN(n5401) );
  OAI21_X1 U6083 ( .B1(n6066), .B2(n5563), .A(n3638), .ZN(n5400) );
  OAI21_X1 U6084 ( .B1(n5367), .B2(n5401), .A(n5400), .ZN(n5402) );
  INV_X1 U6085 ( .A(n5402), .ZN(n5403) );
  AND2_X1 U6086 ( .A1(n3946), .A2(n5407), .ZN(n5410) );
  OAI22_X1 U6087 ( .A1(n5367), .A2(n5298), .B1(n5412), .B2(n5452), .ZN(n5408)
         );
  INV_X1 U6088 ( .A(n5408), .ZN(n5409) );
  OAI211_X1 U6089 ( .C1(n5761), .C2(n5410), .A(n5409), .B(n3630), .ZN(n5411)
         );
  OAI21_X1 U6090 ( .B1(n5412), .B2(n3860), .A(n7212), .ZN(n5413) );
  INV_X1 U6091 ( .A(n5428), .ZN(n5414) );
  NAND2_X1 U6092 ( .A1(n5414), .A2(n7524), .ZN(n7560) );
  INV_X1 U6093 ( .A(n6678), .ZN(n5415) );
  NOR2_X1 U6095 ( .A1(n3953), .A2(n5416), .ZN(n5420) );
  NAND2_X1 U6096 ( .A1(n5417), .A2(n5591), .ZN(n5791) );
  OAI21_X1 U6097 ( .B1(n3638), .B2(n6066), .A(n5791), .ZN(n5418) );
  OR3_X1 U6098 ( .A1(n5420), .A2(n5419), .A3(n5418), .ZN(n5421) );
  NOR2_X1 U6099 ( .A1(n5422), .A2(n5421), .ZN(n5760) );
  NAND2_X1 U6100 ( .A1(n5760), .A2(n5423), .ZN(n5424) );
  NAND2_X1 U6101 ( .A1(n5428), .A2(n5424), .ZN(n6475) );
  NAND2_X1 U6102 ( .A1(n7530), .A2(n6475), .ZN(n6471) );
  INV_X1 U6103 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n7562) );
  NAND2_X1 U6104 ( .A1(n6471), .A2(n7562), .ZN(n7553) );
  INV_X1 U6105 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6653) );
  AOI21_X1 U6106 ( .B1(n7560), .B2(n7553), .A(n6653), .ZN(n5426) );
  INV_X1 U6107 ( .A(REIP_REG_1__SCAN_IN), .ZN(n7353) );
  NOR2_X1 U6108 ( .A1(n7524), .A2(n7353), .ZN(n5425) );
  AOI211_X1 U6109 ( .C1(n7545), .C2(n5427), .A(n5426), .B(n5425), .ZN(n5430)
         );
  INV_X1 U6110 ( .A(n7188), .ZN(n6646) );
  NAND2_X1 U6111 ( .A1(n5428), .A2(n6646), .ZN(n7561) );
  NAND2_X1 U6112 ( .A1(n7561), .A2(n6475), .ZN(n7528) );
  NAND2_X1 U6113 ( .A1(n7562), .A2(n7561), .ZN(n5583) );
  NAND3_X1 U6114 ( .A1(n7508), .A2(n5583), .A3(n6653), .ZN(n5429) );
  OAI211_X1 U6115 ( .C1(n5431), .C2(n7506), .A(n5430), .B(n5429), .ZN(U3017)
         );
  AND2_X1 U6116 ( .A1(n7421), .A2(DATAI_22_), .ZN(n5966) );
  INV_X1 U6117 ( .A(n5966), .ZN(n6404) );
  INV_X1 U6118 ( .A(n4157), .ZN(n5465) );
  AND2_X1 U6119 ( .A1(n3646), .A2(n5465), .ZN(n5434) );
  INV_X1 U6120 ( .A(n5444), .ZN(n5435) );
  NOR2_X1 U6121 ( .A1(n7715), .A2(n5838), .ZN(n6253) );
  INV_X1 U6122 ( .A(n4278), .ZN(n6648) );
  INV_X1 U6123 ( .A(n5727), .ZN(n5914) );
  INV_X1 U6124 ( .A(n5438), .ZN(n7169) );
  INV_X1 U6125 ( .A(n5439), .ZN(n5570) );
  AOI21_X1 U6126 ( .B1(n5914), .B2(n5844), .A(n5570), .ZN(n5443) );
  NOR2_X1 U6127 ( .A1(n5444), .A2(n7726), .ZN(n5812) );
  NOR2_X1 U6128 ( .A1(n5812), .A2(n6375), .ZN(n5441) );
  NAND3_X1 U6129 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n7198), .ZN(n5658) );
  AOI22_X1 U6130 ( .A1(n5443), .A2(n5441), .B1(n6375), .B2(n5658), .ZN(n5440)
         );
  NAND2_X1 U6131 ( .A1(n5922), .A2(n5440), .ZN(n5569) );
  INV_X1 U6132 ( .A(n5441), .ZN(n5442) );
  OAI22_X1 U6133 ( .A1(n5443), .A2(n5442), .B1(n5838), .B2(n5658), .ZN(n5568)
         );
  AOI22_X1 U6134 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n5569), .B1(n6329), 
        .B2(n5568), .ZN(n5448) );
  NOR2_X2 U6135 ( .A1(n5444), .A2(n5732), .ZN(n6028) );
  NAND2_X1 U6136 ( .A1(n7421), .A2(DATAI_30_), .ZN(n5964) );
  INV_X1 U6137 ( .A(n5964), .ZN(n6406) );
  NAND2_X1 U6138 ( .A1(n7437), .A2(STATE2_REG_3__SCAN_IN), .ZN(n7722) );
  INV_X1 U6139 ( .A(n7722), .ZN(n6645) );
  NOR2_X2 U6140 ( .A1(n5564), .A2(n5446), .ZN(n6402) );
  AOI22_X1 U6141 ( .A1(n6028), .A2(n6406), .B1(n6402), .B2(n5570), .ZN(n5447)
         );
  OAI211_X1 U6142 ( .C1(n6404), .C2(n6095), .A(n5448), .B(n5447), .ZN(U3082)
         );
  AND2_X1 U6143 ( .A1(n7421), .A2(DATAI_19_), .ZN(n5960) );
  INV_X1 U6144 ( .A(n5960), .ZN(n6418) );
  INV_X1 U6145 ( .A(DATAI_3_), .ZN(n6088) );
  AOI22_X1 U6146 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n5569), .B1(n6354), 
        .B2(n5568), .ZN(n5451) );
  NAND2_X1 U6147 ( .A1(n7421), .A2(DATAI_27_), .ZN(n5958) );
  INV_X1 U6148 ( .A(n5958), .ZN(n6420) );
  NOR2_X1 U6149 ( .A1(n5564), .A2(n5449), .ZN(n6416) );
  AOI22_X1 U6150 ( .A1(n6028), .A2(n6420), .B1(n6416), .B2(n5570), .ZN(n5450)
         );
  OAI211_X1 U6151 ( .C1(n6418), .C2(n6095), .A(n5451), .B(n5450), .ZN(U3079)
         );
  AND2_X1 U6152 ( .A1(n7421), .A2(DATAI_20_), .ZN(n5954) );
  INV_X1 U6153 ( .A(n5954), .ZN(n6411) );
  AOI22_X1 U6154 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n5569), .B1(n6344), 
        .B2(n5568), .ZN(n5454) );
  NAND2_X1 U6155 ( .A1(n7421), .A2(DATAI_28_), .ZN(n5952) );
  INV_X1 U6156 ( .A(n5952), .ZN(n6413) );
  AOI22_X1 U6157 ( .A1(n6028), .A2(n6413), .B1(n6409), .B2(n5570), .ZN(n5453)
         );
  OAI211_X1 U6158 ( .C1(n6411), .C2(n6095), .A(n5454), .B(n5453), .ZN(U3080)
         );
  AND2_X1 U6159 ( .A1(n7421), .A2(DATAI_23_), .ZN(n5972) );
  INV_X1 U6160 ( .A(n5972), .ZN(n6397) );
  NOR2_X1 U6161 ( .A1(n3646), .A2(n4157), .ZN(n5455) );
  AOI21_X1 U6162 ( .B1(n5460), .B2(STATEBS16_REG_SCAN_IN), .A(n6375), .ZN(
        n5457) );
  NAND2_X1 U6163 ( .A1(n3663), .A2(n5438), .ZN(n5864) );
  NAND3_X1 U6164 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n7198), .A3(n7193), .ZN(n5859) );
  NOR2_X1 U6165 ( .A1(n5726), .A2(n5859), .ZN(n5565) );
  AOI21_X1 U6166 ( .B1(n5914), .B2(n5870), .A(n5565), .ZN(n5459) );
  AOI22_X1 U6167 ( .A1(n5457), .A2(n5459), .B1(n6375), .B2(n5859), .ZN(n5456)
         );
  NAND2_X1 U6168 ( .A1(n5922), .A2(n5456), .ZN(n5562) );
  INV_X1 U6169 ( .A(n5457), .ZN(n5458) );
  OAI22_X1 U6170 ( .A1(n5459), .A2(n5458), .B1(n5838), .B2(n5859), .ZN(n5561)
         );
  AOI22_X1 U6171 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n5562), .B1(n6360), 
        .B2(n5561), .ZN(n5462) );
  NAND2_X1 U6172 ( .A1(n7421), .A2(DATAI_31_), .ZN(n5970) );
  INV_X1 U6173 ( .A(n5970), .ZN(n6399) );
  AOI22_X1 U6174 ( .A1(n6148), .A2(n6399), .B1(n6395), .B2(n5565), .ZN(n5461)
         );
  OAI211_X1 U6175 ( .C1(n6397), .C2(n6026), .A(n5462), .B(n5461), .ZN(U3067)
         );
  AOI22_X1 U6176 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n5562), .B1(n6329), 
        .B2(n5561), .ZN(n5464) );
  AOI22_X1 U6177 ( .A1(n6148), .A2(n6406), .B1(n6402), .B2(n5565), .ZN(n5463)
         );
  OAI211_X1 U6178 ( .C1(n6404), .C2(n6026), .A(n5464), .B(n5463), .ZN(U3066)
         );
  NOR2_X1 U6179 ( .A1(n3646), .A2(n5465), .ZN(n5466) );
  AOI21_X1 U6180 ( .B1(n5810), .B2(STATEBS16_REG_SCAN_IN), .A(n6375), .ZN(
        n5468) );
  AND2_X1 U6181 ( .A1(n4278), .A2(n3645), .ZN(n5684) );
  NAND3_X1 U6182 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n7193), .ZN(n5818) );
  NOR2_X1 U6183 ( .A1(n5726), .A2(n5818), .ZN(n5575) );
  AOI21_X1 U6184 ( .B1(n5684), .B2(n5870), .A(n5575), .ZN(n5470) );
  AOI22_X1 U6185 ( .A1(n5468), .A2(n5470), .B1(n6375), .B2(n5818), .ZN(n5467)
         );
  NAND2_X1 U6186 ( .A1(n5922), .A2(n5467), .ZN(n5574) );
  INV_X1 U6187 ( .A(n5468), .ZN(n5469) );
  OAI22_X1 U6188 ( .A1(n5470), .A2(n5469), .B1(n5838), .B2(n5818), .ZN(n5573)
         );
  AOI22_X1 U6189 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n5574), .B1(n6354), 
        .B2(n5573), .ZN(n5472) );
  AOI22_X1 U6190 ( .A1(n6114), .A2(n6420), .B1(n6416), .B2(n5575), .ZN(n5471)
         );
  OAI211_X1 U6191 ( .C1(n6418), .C2(n6143), .A(n5472), .B(n5471), .ZN(U3127)
         );
  AOI22_X1 U6192 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n5574), .B1(n6360), 
        .B2(n5573), .ZN(n5474) );
  AOI22_X1 U6193 ( .A1(n6114), .A2(n6399), .B1(n6395), .B2(n5575), .ZN(n5473)
         );
  OAI211_X1 U6194 ( .C1(n6397), .C2(n6143), .A(n5474), .B(n5473), .ZN(U3131)
         );
  AOI22_X1 U6195 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n5574), .B1(n6329), 
        .B2(n5573), .ZN(n5476) );
  AOI22_X1 U6196 ( .A1(n6114), .A2(n6406), .B1(n6402), .B2(n5575), .ZN(n5475)
         );
  OAI211_X1 U6197 ( .C1(n6404), .C2(n6143), .A(n5476), .B(n5475), .ZN(U3130)
         );
  AOI22_X1 U6198 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n5562), .B1(n6344), 
        .B2(n5561), .ZN(n5478) );
  AOI22_X1 U6199 ( .A1(n6148), .A2(n6413), .B1(n6409), .B2(n5565), .ZN(n5477)
         );
  OAI211_X1 U6200 ( .C1(n6411), .C2(n6026), .A(n5478), .B(n5477), .ZN(U3064)
         );
  AOI22_X1 U6201 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n5574), .B1(n6344), 
        .B2(n5573), .ZN(n5480) );
  AOI22_X1 U6202 ( .A1(n6114), .A2(n6413), .B1(n6409), .B2(n5575), .ZN(n5479)
         );
  OAI211_X1 U6203 ( .C1(n6411), .C2(n6143), .A(n5480), .B(n5479), .ZN(U3128)
         );
  AOI22_X1 U6204 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n5562), .B1(n6354), 
        .B2(n5561), .ZN(n5482) );
  AOI22_X1 U6205 ( .A1(n6148), .A2(n6420), .B1(n6416), .B2(n5565), .ZN(n5481)
         );
  OAI211_X1 U6206 ( .C1(n6418), .C2(n6026), .A(n5482), .B(n5481), .ZN(U3063)
         );
  AOI22_X1 U6207 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n5569), .B1(n6360), 
        .B2(n5568), .ZN(n5484) );
  AOI22_X1 U6208 ( .A1(n6028), .A2(n6399), .B1(n6395), .B2(n5570), .ZN(n5483)
         );
  OAI211_X1 U6209 ( .C1(n6397), .C2(n6095), .A(n5484), .B(n5483), .ZN(U3083)
         );
  OR2_X1 U6210 ( .A1(n5487), .A2(n5488), .ZN(n5489) );
  AND2_X1 U6211 ( .A1(n5486), .A2(n5489), .ZN(n7570) );
  INV_X1 U6212 ( .A(n6919), .ZN(n7366) );
  OR2_X1 U6213 ( .A1(n5491), .A2(n5492), .ZN(n5493) );
  NAND2_X1 U6214 ( .A1(n5490), .A2(n5493), .ZN(n7564) );
  OAI22_X1 U6215 ( .A1(n7564), .A2(n6917), .B1(n7565), .B2(n7369), .ZN(n5494)
         );
  AOI21_X1 U6216 ( .B1(n7570), .B2(n7366), .A(n5494), .ZN(n5495) );
  INV_X1 U6217 ( .A(n5495), .ZN(U2854) );
  AND2_X1 U6218 ( .A1(n5361), .A2(n5496), .ZN(n5497) );
  OR2_X1 U6219 ( .A1(n5497), .A2(n5487), .ZN(n6293) );
  AND2_X1 U6220 ( .A1(n5498), .A2(n5499), .ZN(n5500) );
  NOR2_X1 U6221 ( .A1(n5491), .A2(n5500), .ZN(n7450) );
  AOI22_X1 U6222 ( .A1(n7450), .A2(n6914), .B1(n6913), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n5501) );
  OAI21_X1 U6223 ( .B1(n6293), .B2(n6919), .A(n5501), .ZN(U2855) );
  INV_X1 U6224 ( .A(n3662), .ZN(n5503) );
  NAND2_X1 U6225 ( .A1(n3640), .A2(n5503), .ZN(n5686) );
  NOR2_X1 U6226 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n7198), .ZN(n5942)
         );
  NAND2_X1 U6227 ( .A1(n5942), .A2(n7193), .ZN(n5509) );
  INV_X1 U6228 ( .A(n5509), .ZN(n5508) );
  INV_X1 U6229 ( .A(n5511), .ZN(n5506) );
  INV_X1 U6230 ( .A(n5949), .ZN(n5505) );
  NOR2_X1 U6231 ( .A1(n5726), .A2(n5509), .ZN(n5626) );
  AOI21_X1 U6232 ( .B1(n5684), .B2(n5505), .A(n5626), .ZN(n5510) );
  NAND2_X1 U6233 ( .A1(n5506), .A2(n5510), .ZN(n5507) );
  OAI211_X1 U6234 ( .C1(n5925), .C2(n5508), .A(n5922), .B(n5507), .ZN(n5625)
         );
  OAI22_X1 U6235 ( .A1(n5511), .A2(n5510), .B1(n5838), .B2(n5509), .ZN(n5624)
         );
  AOI22_X1 U6236 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n5625), .B1(n6360), 
        .B2(n5624), .ZN(n5514) );
  AOI22_X1 U6237 ( .A1(n3621), .A2(n5972), .B1(n5626), .B2(n6395), .ZN(n5513)
         );
  OAI211_X1 U6238 ( .C1(n5947), .C2(n5970), .A(n5514), .B(n5513), .ZN(U3099)
         );
  AOI22_X1 U6239 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n5625), .B1(n6329), 
        .B2(n5624), .ZN(n5516) );
  AOI22_X1 U6240 ( .A1(n3621), .A2(n5966), .B1(n5626), .B2(n6402), .ZN(n5515)
         );
  OAI211_X1 U6241 ( .C1(n5947), .C2(n5964), .A(n5516), .B(n5515), .ZN(U3098)
         );
  AOI22_X1 U6242 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5625), .B1(n6344), 
        .B2(n5624), .ZN(n5518) );
  AOI22_X1 U6243 ( .A1(n3621), .A2(n5954), .B1(n5626), .B2(n6409), .ZN(n5517)
         );
  OAI211_X1 U6244 ( .C1(n5947), .C2(n5952), .A(n5518), .B(n5517), .ZN(U3096)
         );
  AOI22_X1 U6245 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n5625), .B1(n6354), 
        .B2(n5624), .ZN(n5520) );
  AOI22_X1 U6246 ( .A1(n3621), .A2(n5960), .B1(n5626), .B2(n6416), .ZN(n5519)
         );
  OAI211_X1 U6247 ( .C1(n5947), .C2(n5958), .A(n5520), .B(n5519), .ZN(U3095)
         );
  NAND2_X1 U6248 ( .A1(n5523), .A2(n5524), .ZN(n5525) );
  AND2_X1 U6249 ( .A1(n5521), .A2(n5525), .ZN(n7592) );
  INV_X1 U6250 ( .A(n7592), .ZN(n6070) );
  AND2_X1 U6251 ( .A1(n5654), .A2(n5527), .ZN(n5528) );
  NOR2_X1 U6252 ( .A1(n5526), .A2(n5528), .ZN(n7585) );
  AOI22_X1 U6253 ( .A1(n7585), .A2(n6914), .B1(n6913), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n5529) );
  OAI21_X1 U6254 ( .B1(n6070), .B2(n6919), .A(n5529), .ZN(U2852) );
  NOR2_X1 U6255 ( .A1(n5530), .A2(n5531), .ZN(n5532) );
  NOR2_X1 U6256 ( .A1(n5360), .A2(n5532), .ZN(n7378) );
  INV_X1 U6257 ( .A(n7378), .ZN(n6880) );
  INV_X1 U6258 ( .A(n5533), .ZN(n5536) );
  AOI21_X1 U6259 ( .B1(n5536), .B2(n5535), .A(n5534), .ZN(n7468) );
  AOI22_X1 U6260 ( .A1(n6914), .A2(n7468), .B1(n6913), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n5537) );
  OAI21_X1 U6261 ( .B1(n6880), .B2(n6919), .A(n5537), .ZN(U2857) );
  NAND2_X1 U6262 ( .A1(n5539), .A2(n5538), .ZN(n5540) );
  NAND2_X1 U6263 ( .A1(n5498), .A2(n5540), .ZN(n6862) );
  INV_X1 U6264 ( .A(n6862), .ZN(n5541) );
  AOI22_X1 U6265 ( .A1(n6914), .A2(n5541), .B1(n6913), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n5542) );
  OAI21_X1 U6266 ( .B1(n6089), .B2(n6919), .A(n5542), .ZN(U2856) );
  AND2_X1 U6267 ( .A1(n7421), .A2(DATAI_17_), .ZN(n6175) );
  INV_X1 U6268 ( .A(n6175), .ZN(n6425) );
  AOI22_X1 U6269 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n5574), .B1(n6349), 
        .B2(n5573), .ZN(n5544) );
  NAND2_X1 U6270 ( .A1(n7421), .A2(DATAI_25_), .ZN(n6173) );
  INV_X1 U6271 ( .A(n6173), .ZN(n6427) );
  NOR2_X1 U6272 ( .A1(n5564), .A2(n3956), .ZN(n6423) );
  AOI22_X1 U6273 ( .A1(n6114), .A2(n6427), .B1(n3678), .B2(n5575), .ZN(n5543)
         );
  OAI211_X1 U6274 ( .C1(n6425), .C2(n6143), .A(n5544), .B(n5543), .ZN(U3125)
         );
  AND2_X1 U6275 ( .A1(n7421), .A2(DATAI_18_), .ZN(n6181) );
  INV_X1 U6276 ( .A(n6181), .ZN(n6432) );
  AOI22_X1 U6277 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n5569), .B1(n6339), 
        .B2(n5568), .ZN(n5546) );
  NAND2_X1 U6278 ( .A1(n7421), .A2(DATAI_26_), .ZN(n6179) );
  INV_X1 U6279 ( .A(n6179), .ZN(n6434) );
  AOI22_X1 U6280 ( .A1(n6028), .A2(n6434), .B1(n6430), .B2(n5570), .ZN(n5545)
         );
  OAI211_X1 U6281 ( .C1(n6432), .C2(n6095), .A(n5546), .B(n5545), .ZN(U3078)
         );
  AOI22_X1 U6282 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n5574), .B1(n6339), 
        .B2(n5573), .ZN(n5548) );
  AOI22_X1 U6283 ( .A1(n6114), .A2(n6434), .B1(n6430), .B2(n5575), .ZN(n5547)
         );
  OAI211_X1 U6284 ( .C1(n6432), .C2(n6143), .A(n5548), .B(n5547), .ZN(U3126)
         );
  AND2_X1 U6285 ( .A1(n7421), .A2(DATAI_21_), .ZN(n6188) );
  INV_X1 U6286 ( .A(n6188), .ZN(n6390) );
  INV_X1 U6287 ( .A(DATAI_5_), .ZN(n6944) );
  AOI22_X1 U6288 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n5569), .B1(n6334), 
        .B2(n5568), .ZN(n5550) );
  NAND2_X1 U6289 ( .A1(n7421), .A2(DATAI_29_), .ZN(n6185) );
  INV_X1 U6290 ( .A(n6185), .ZN(n6392) );
  AOI22_X1 U6291 ( .A1(n6028), .A2(n6392), .B1(n7767), .B2(n5570), .ZN(n5549)
         );
  OAI211_X1 U6292 ( .C1(n6390), .C2(n6095), .A(n5550), .B(n5549), .ZN(U3081)
         );
  AOI22_X1 U6293 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n5574), .B1(n6334), 
        .B2(n5573), .ZN(n5552) );
  AOI22_X1 U6294 ( .A1(n6114), .A2(n6392), .B1(n7767), .B2(n5575), .ZN(n5551)
         );
  OAI211_X1 U6295 ( .C1(n6390), .C2(n6143), .A(n5552), .B(n5551), .ZN(U3129)
         );
  AOI22_X1 U6296 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n5569), .B1(n6349), 
        .B2(n5568), .ZN(n5554) );
  AOI22_X1 U6297 ( .A1(n6028), .A2(n6427), .B1(n3678), .B2(n5570), .ZN(n5553)
         );
  OAI211_X1 U6298 ( .C1(n6425), .C2(n6095), .A(n5554), .B(n5553), .ZN(U3077)
         );
  AOI22_X1 U6299 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n5562), .B1(n6334), 
        .B2(n5561), .ZN(n5556) );
  AOI22_X1 U6300 ( .A1(n6148), .A2(n6392), .B1(n7767), .B2(n5565), .ZN(n5555)
         );
  OAI211_X1 U6301 ( .C1(n6390), .C2(n6026), .A(n5556), .B(n5555), .ZN(U3065)
         );
  AOI22_X1 U6302 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n5562), .B1(n6339), 
        .B2(n5561), .ZN(n5558) );
  AOI22_X1 U6303 ( .A1(n6148), .A2(n6434), .B1(n6430), .B2(n5565), .ZN(n5557)
         );
  OAI211_X1 U6304 ( .C1(n6432), .C2(n6026), .A(n5558), .B(n5557), .ZN(U3062)
         );
  AOI22_X1 U6305 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n5562), .B1(n6349), 
        .B2(n5561), .ZN(n5560) );
  AOI22_X1 U6306 ( .A1(n6148), .A2(n6427), .B1(n3678), .B2(n5565), .ZN(n5559)
         );
  OAI211_X1 U6307 ( .C1(n6425), .C2(n6026), .A(n5560), .B(n5559), .ZN(U3061)
         );
  AND2_X1 U6308 ( .A1(n7421), .A2(DATAI_16_), .ZN(n6196) );
  INV_X1 U6309 ( .A(n6196), .ZN(n6441) );
  AOI22_X1 U6310 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n5562), .B1(n6324), 
        .B2(n5561), .ZN(n5567) );
  NAND2_X1 U6311 ( .A1(n7421), .A2(DATAI_24_), .ZN(n6193) );
  INV_X1 U6312 ( .A(n6193), .ZN(n6445) );
  NOR2_X1 U6313 ( .A1(n5564), .A2(n5563), .ZN(n6439) );
  AOI22_X1 U6314 ( .A1(n6148), .A2(n6445), .B1(n6439), .B2(n5565), .ZN(n5566)
         );
  OAI211_X1 U6315 ( .C1(n6441), .C2(n6026), .A(n5567), .B(n5566), .ZN(U3060)
         );
  AOI22_X1 U6316 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n5569), .B1(n6324), 
        .B2(n5568), .ZN(n5572) );
  AOI22_X1 U6317 ( .A1(n6028), .A2(n6445), .B1(n6439), .B2(n5570), .ZN(n5571)
         );
  OAI211_X1 U6318 ( .C1(n6441), .C2(n6095), .A(n5572), .B(n5571), .ZN(U3076)
         );
  AOI22_X1 U6319 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n5574), .B1(n6324), 
        .B2(n5573), .ZN(n5577) );
  AOI22_X1 U6320 ( .A1(n6114), .A2(n6445), .B1(n6439), .B2(n5575), .ZN(n5576)
         );
  OAI211_X1 U6321 ( .C1(n6441), .C2(n6143), .A(n5577), .B(n5576), .ZN(U3124)
         );
  OAI21_X1 U6322 ( .B1(n5578), .B2(n5580), .A(n5579), .ZN(n7390) );
  INV_X1 U6323 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n5582) );
  NOR2_X1 U6324 ( .A1(n5582), .A2(n5581), .ZN(n7456) );
  OAI21_X1 U6325 ( .B1(n6653), .B2(n7562), .A(n7475), .ZN(n7473) );
  NAND2_X1 U6326 ( .A1(n7456), .A2(n7473), .ZN(n7459) );
  NAND2_X1 U6327 ( .A1(n7528), .A2(n5583), .ZN(n7474) );
  NAND2_X1 U6328 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5979) );
  INV_X1 U6329 ( .A(n5979), .ZN(n5584) );
  NAND2_X1 U6330 ( .A1(n7456), .A2(n5584), .ZN(n6053) );
  OAI22_X1 U6331 ( .A1(n7530), .A2(n7459), .B1(n7474), .B2(n6053), .ZN(n5586)
         );
  NOR2_X1 U6332 ( .A1(n7460), .A2(n7459), .ZN(n5585) );
  OAI21_X1 U6333 ( .B1(n6475), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n7560), 
        .ZN(n7526) );
  AOI21_X1 U6334 ( .B1(n7528), .B2(n5979), .A(n7526), .ZN(n7469) );
  OAI21_X1 U6335 ( .B1(n6580), .B2(n5585), .A(n7469), .ZN(n7457) );
  OAI21_X1 U6336 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n5586), .A(n7457), 
        .ZN(n5589) );
  INV_X1 U6337 ( .A(n7564), .ZN(n5587) );
  AOI22_X1 U6338 ( .A1(n7545), .A2(n5587), .B1(n7544), .B2(REIP_REG_5__SCAN_IN), .ZN(n5588) );
  OAI211_X1 U6339 ( .C1(n7390), .C2(n7506), .A(n5589), .B(n5588), .ZN(U3013)
         );
  NAND2_X1 U6340 ( .A1(n5708), .A2(DATAI_10_), .ZN(n5720) );
  NOR2_X1 U6341 ( .A1(n5593), .A2(n5755), .ZN(n5705) );
  AOI22_X1 U6342 ( .A1(n5755), .A2(EAX_REG_26__SCAN_IN), .B1(n5617), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U6343 ( .A1(n5720), .A2(n5594), .ZN(U2934) );
  NAND2_X1 U6344 ( .A1(n5708), .A2(DATAI_1_), .ZN(n5614) );
  AOI22_X1 U6345 ( .A1(n5755), .A2(EAX_REG_1__SCAN_IN), .B1(n5617), .B2(
        LWORD_REG_1__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U6346 ( .A1(n5614), .A2(n5595), .ZN(U2940) );
  NAND2_X1 U6347 ( .A1(n5708), .A2(DATAI_11_), .ZN(n5714) );
  AOI22_X1 U6348 ( .A1(n5755), .A2(EAX_REG_27__SCAN_IN), .B1(n5617), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n5596) );
  NAND2_X1 U6349 ( .A1(n5714), .A2(n5596), .ZN(U2935) );
  NAND2_X1 U6350 ( .A1(n5708), .A2(DATAI_13_), .ZN(n5707) );
  AOI22_X1 U6351 ( .A1(n5755), .A2(EAX_REG_29__SCAN_IN), .B1(n5617), .B2(
        UWORD_REG_13__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U6352 ( .A1(n5707), .A2(n5597), .ZN(U2937) );
  NAND2_X1 U6353 ( .A1(n5708), .A2(DATAI_0_), .ZN(n5609) );
  AOI22_X1 U6354 ( .A1(n5755), .A2(EAX_REG_0__SCAN_IN), .B1(n5617), .B2(
        LWORD_REG_0__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U6355 ( .A1(n5609), .A2(n5598), .ZN(U2939) );
  NAND2_X1 U6356 ( .A1(n5708), .A2(DATAI_4_), .ZN(n5619) );
  AOI22_X1 U6357 ( .A1(n5755), .A2(EAX_REG_4__SCAN_IN), .B1(n5617), .B2(
        LWORD_REG_4__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U6358 ( .A1(n5619), .A2(n5599), .ZN(U2943) );
  AOI22_X1 U6359 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n5625), .B1(n6324), 
        .B2(n5624), .ZN(n5601) );
  AOI22_X1 U6360 ( .A1(n3621), .A2(n6196), .B1(n6439), .B2(n5626), .ZN(n5600)
         );
  OAI211_X1 U6361 ( .C1(n5947), .C2(n6193), .A(n5601), .B(n5600), .ZN(U3092)
         );
  NAND2_X1 U6362 ( .A1(n5708), .A2(DATAI_6_), .ZN(n5616) );
  AOI22_X1 U6363 ( .A1(n5755), .A2(EAX_REG_6__SCAN_IN), .B1(n5617), .B2(
        LWORD_REG_6__SCAN_IN), .ZN(n5602) );
  NAND2_X1 U6364 ( .A1(n5616), .A2(n5602), .ZN(U2945) );
  NAND2_X1 U6365 ( .A1(n5708), .A2(DATAI_8_), .ZN(n5605) );
  AOI22_X1 U6366 ( .A1(n5755), .A2(EAX_REG_24__SCAN_IN), .B1(n5617), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n5603) );
  NAND2_X1 U6367 ( .A1(n5605), .A2(n5603), .ZN(U2932) );
  AOI22_X1 U6368 ( .A1(n5755), .A2(EAX_REG_8__SCAN_IN), .B1(n5617), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n5604) );
  NAND2_X1 U6369 ( .A1(n5605), .A2(n5604), .ZN(U2947) );
  NAND2_X1 U6370 ( .A1(n5708), .A2(DATAI_5_), .ZN(n5757) );
  AOI22_X1 U6371 ( .A1(n5755), .A2(EAX_REG_21__SCAN_IN), .B1(n5617), .B2(
        UWORD_REG_5__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U6372 ( .A1(n5757), .A2(n5606), .ZN(U2929) );
  INV_X1 U6373 ( .A(DATAI_9_), .ZN(n6252) );
  OR2_X1 U6374 ( .A1(n6063), .A2(n6252), .ZN(n5724) );
  AOI22_X1 U6375 ( .A1(n5755), .A2(EAX_REG_25__SCAN_IN), .B1(n5617), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n5607) );
  NAND2_X1 U6376 ( .A1(n5724), .A2(n5607), .ZN(U2933) );
  AOI22_X1 U6377 ( .A1(n5755), .A2(EAX_REG_16__SCAN_IN), .B1(n5617), .B2(
        UWORD_REG_0__SCAN_IN), .ZN(n5608) );
  NAND2_X1 U6378 ( .A1(n5609), .A2(n5608), .ZN(U2924) );
  NAND2_X1 U6379 ( .A1(n5708), .A2(DATAI_3_), .ZN(n5716) );
  AOI22_X1 U6380 ( .A1(n5755), .A2(EAX_REG_19__SCAN_IN), .B1(n5617), .B2(
        UWORD_REG_3__SCAN_IN), .ZN(n5610) );
  NAND2_X1 U6381 ( .A1(n5716), .A2(n5610), .ZN(U2927) );
  NAND2_X1 U6382 ( .A1(n5708), .A2(DATAI_2_), .ZN(n5718) );
  AOI22_X1 U6383 ( .A1(n5755), .A2(EAX_REG_18__SCAN_IN), .B1(n5617), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U6384 ( .A1(n5718), .A2(n5611), .ZN(U2926) );
  NAND2_X1 U6385 ( .A1(n5708), .A2(DATAI_7_), .ZN(n5754) );
  AOI22_X1 U6386 ( .A1(n5755), .A2(EAX_REG_23__SCAN_IN), .B1(n5617), .B2(
        UWORD_REG_7__SCAN_IN), .ZN(n5612) );
  NAND2_X1 U6387 ( .A1(n5754), .A2(n5612), .ZN(U2931) );
  AOI22_X1 U6388 ( .A1(n5755), .A2(EAX_REG_17__SCAN_IN), .B1(n5617), .B2(
        UWORD_REG_1__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U6389 ( .A1(n5614), .A2(n5613), .ZN(U2925) );
  AOI22_X1 U6390 ( .A1(n5755), .A2(EAX_REG_22__SCAN_IN), .B1(n5617), .B2(
        UWORD_REG_6__SCAN_IN), .ZN(n5615) );
  NAND2_X1 U6391 ( .A1(n5616), .A2(n5615), .ZN(U2930) );
  AOI22_X1 U6392 ( .A1(n5755), .A2(EAX_REG_20__SCAN_IN), .B1(n5617), .B2(
        UWORD_REG_4__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U6393 ( .A1(n5619), .A2(n5618), .ZN(U2928) );
  AOI22_X1 U6394 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n5625), .B1(n6349), 
        .B2(n5624), .ZN(n5621) );
  AOI22_X1 U6395 ( .A1(n3621), .A2(n6175), .B1(n5626), .B2(n3678), .ZN(n5620)
         );
  OAI211_X1 U6396 ( .C1(n5947), .C2(n6173), .A(n5621), .B(n5620), .ZN(U3093)
         );
  AOI22_X1 U6397 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n5625), .B1(n6334), 
        .B2(n5624), .ZN(n5623) );
  AOI22_X1 U6398 ( .A1(n3621), .A2(n6188), .B1(n5626), .B2(n7767), .ZN(n5622)
         );
  OAI211_X1 U6399 ( .C1(n5947), .C2(n6185), .A(n5623), .B(n5622), .ZN(U3097)
         );
  AOI22_X1 U6400 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n5625), .B1(n6339), 
        .B2(n5624), .ZN(n5628) );
  AOI22_X1 U6401 ( .A1(n3621), .A2(n6181), .B1(n5626), .B2(n6430), .ZN(n5627)
         );
  OAI211_X1 U6402 ( .C1(n5947), .C2(n6179), .A(n5628), .B(n5627), .ZN(U3094)
         );
  NOR2_X1 U6403 ( .A1(n5629), .A2(n7198), .ZN(n6045) );
  AOI21_X1 U6404 ( .B1(n5684), .B2(n5844), .A(n6045), .ZN(n5635) );
  AND2_X1 U6405 ( .A1(n3646), .A2(n4157), .ZN(n5630) );
  NAND2_X1 U6406 ( .A1(n3662), .A2(n5630), .ZN(n5634) );
  INV_X1 U6407 ( .A(n5634), .ZN(n5631) );
  NAND2_X1 U6408 ( .A1(n5925), .A2(n7726), .ZN(n6313) );
  OAI21_X1 U6409 ( .B1(n5631), .B2(n7052), .A(n6313), .ZN(n5632) );
  NAND3_X1 U6410 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5836) );
  AOI22_X1 U6411 ( .A1(n5635), .A2(n5632), .B1(n6375), .B2(n5836), .ZN(n5633)
         );
  INV_X1 U6412 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n5639) );
  NOR2_X2 U6413 ( .A1(n5634), .A2(n5732), .ZN(n6140) );
  OAI22_X1 U6414 ( .A1(n5635), .A2(n6375), .B1(n5836), .B2(n5838), .ZN(n6044)
         );
  AOI22_X1 U6415 ( .A1(n6409), .A2(n6045), .B1(n6344), .B2(n6044), .ZN(n5636)
         );
  OAI21_X1 U6416 ( .B1(n6411), .B2(n6047), .A(n5636), .ZN(n5637) );
  AOI21_X1 U6417 ( .B1(n6413), .B2(n6140), .A(n5637), .ZN(n5638) );
  OAI21_X1 U6418 ( .B1(n6051), .B2(n5639), .A(n5638), .ZN(U3144) );
  INV_X1 U6419 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5643) );
  AOI22_X1 U6420 ( .A1(n6402), .A2(n6045), .B1(n6329), .B2(n6044), .ZN(n5640)
         );
  OAI21_X1 U6421 ( .B1(n6404), .B2(n6047), .A(n5640), .ZN(n5641) );
  AOI21_X1 U6422 ( .B1(n6406), .B2(n6140), .A(n5641), .ZN(n5642) );
  OAI21_X1 U6423 ( .B1(n6051), .B2(n5643), .A(n5642), .ZN(U3146) );
  INV_X1 U6424 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5647) );
  AOI22_X1 U6425 ( .A1(n6395), .A2(n6045), .B1(n6360), .B2(n6044), .ZN(n5644)
         );
  OAI21_X1 U6426 ( .B1(n6397), .B2(n6047), .A(n5644), .ZN(n5645) );
  AOI21_X1 U6427 ( .B1(n6399), .B2(n6140), .A(n5645), .ZN(n5646) );
  OAI21_X1 U6428 ( .B1(n6051), .B2(n5647), .A(n5646), .ZN(U3147) );
  INV_X1 U6429 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n5651) );
  AOI22_X1 U6430 ( .A1(n6416), .A2(n6045), .B1(n6354), .B2(n6044), .ZN(n5648)
         );
  OAI21_X1 U6431 ( .B1(n6418), .B2(n6047), .A(n5648), .ZN(n5649) );
  AOI21_X1 U6432 ( .B1(n6420), .B2(n6140), .A(n5649), .ZN(n5650) );
  OAI21_X1 U6433 ( .B1(n6051), .B2(n5651), .A(n5650), .ZN(U3143) );
  NAND2_X1 U6434 ( .A1(n5490), .A2(n5652), .ZN(n5653) );
  NAND2_X1 U6435 ( .A1(n5654), .A2(n5653), .ZN(n7575) );
  INV_X1 U6436 ( .A(EBX_REG_6__SCAN_IN), .ZN(n7577) );
  AOI21_X1 U6437 ( .B1(n5655), .B2(n5486), .A(n3728), .ZN(n7580) );
  INV_X1 U6438 ( .A(n7580), .ZN(n6087) );
  OAI222_X1 U6439 ( .A1(n7575), .A2(n6917), .B1(n7577), .B2(n7369), .C1(n6087), 
        .C2(n6919), .ZN(U2853) );
  NAND2_X1 U6440 ( .A1(n3645), .A2(n5925), .ZN(n5950) );
  INV_X1 U6441 ( .A(n5950), .ZN(n5845) );
  NOR2_X1 U6442 ( .A1(n5844), .A2(n6375), .ZN(n5841) );
  INV_X1 U6443 ( .A(n6026), .ZN(n5656) );
  OAI21_X1 U6444 ( .B1(n5656), .B2(n6028), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5657) );
  OAI21_X1 U6445 ( .B1(n5845), .B2(n5841), .A(n5657), .ZN(n5663) );
  NOR2_X1 U6446 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5658), .ZN(n6024)
         );
  INV_X1 U6447 ( .A(n5837), .ZN(n5860) );
  NAND2_X1 U6448 ( .A1(n5860), .A2(n7198), .ZN(n6321) );
  NAND2_X1 U6449 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6321), .ZN(n6318) );
  INV_X1 U6450 ( .A(n5664), .ZN(n5659) );
  NAND2_X1 U6451 ( .A1(n5659), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6322) );
  INV_X1 U6452 ( .A(n5862), .ZN(n5660) );
  OAI211_X1 U6453 ( .C1(n7724), .C2(n6024), .A(n6318), .B(n5660), .ZN(n5661)
         );
  INV_X1 U6454 ( .A(n5661), .ZN(n5662) );
  INV_X1 U6455 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5669) );
  INV_X1 U6456 ( .A(n5844), .ZN(n5665) );
  NAND2_X1 U6457 ( .A1(n5664), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5884) );
  OAI22_X1 U6458 ( .A1(n5665), .A2(n6323), .B1(n6321), .B2(n5884), .ZN(n6023)
         );
  AOI22_X1 U6459 ( .A1(n6416), .A2(n6024), .B1(n6354), .B2(n6023), .ZN(n5666)
         );
  OAI21_X1 U6460 ( .B1(n5958), .B2(n6026), .A(n5666), .ZN(n5667) );
  AOI21_X1 U6461 ( .B1(n5960), .B2(n6028), .A(n5667), .ZN(n5668) );
  OAI21_X1 U6462 ( .B1(n6031), .B2(n5669), .A(n5668), .ZN(U3071) );
  INV_X1 U6463 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5673) );
  AOI22_X1 U6464 ( .A1(n6409), .A2(n6024), .B1(n6344), .B2(n6023), .ZN(n5670)
         );
  OAI21_X1 U6465 ( .B1(n5952), .B2(n6026), .A(n5670), .ZN(n5671) );
  AOI21_X1 U6466 ( .B1(n5954), .B2(n6028), .A(n5671), .ZN(n5672) );
  OAI21_X1 U6467 ( .B1(n6031), .B2(n5673), .A(n5672), .ZN(U3072) );
  INV_X1 U6468 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5677) );
  AOI22_X1 U6469 ( .A1(n6395), .A2(n6024), .B1(n6360), .B2(n6023), .ZN(n5674)
         );
  OAI21_X1 U6470 ( .B1(n5970), .B2(n6026), .A(n5674), .ZN(n5675) );
  AOI21_X1 U6471 ( .B1(n5972), .B2(n6028), .A(n5675), .ZN(n5676) );
  OAI21_X1 U6472 ( .B1(n6031), .B2(n5677), .A(n5676), .ZN(U3075) );
  INV_X1 U6473 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5681) );
  AOI22_X1 U6474 ( .A1(n6402), .A2(n6024), .B1(n6329), .B2(n6023), .ZN(n5678)
         );
  OAI21_X1 U6475 ( .B1(n5964), .B2(n6026), .A(n5678), .ZN(n5679) );
  AOI21_X1 U6476 ( .B1(n5966), .B2(n6028), .A(n5679), .ZN(n5680) );
  OAI21_X1 U6477 ( .B1(n6031), .B2(n5681), .A(n5680), .ZN(U3074) );
  INV_X1 U6478 ( .A(n5686), .ZN(n5813) );
  INV_X1 U6479 ( .A(n3646), .ZN(n5682) );
  NOR2_X1 U6480 ( .A1(n5682), .A2(n7726), .ZN(n5975) );
  AOI21_X1 U6481 ( .B1(n5813), .B2(n5975), .A(n6375), .ZN(n5691) );
  OR2_X1 U6482 ( .A1(n3663), .A2(n5438), .ZN(n6377) );
  INV_X1 U6483 ( .A(n6377), .ZN(n5913) );
  NAND2_X1 U6484 ( .A1(n5911), .A2(n5942), .ZN(n6161) );
  INV_X1 U6485 ( .A(n6161), .ZN(n5683) );
  AOI21_X1 U6486 ( .B1(n5684), .B2(n5913), .A(n5683), .ZN(n5690) );
  INV_X1 U6487 ( .A(n5690), .ZN(n5685) );
  NAND2_X1 U6488 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n5942), .ZN(n6381) );
  INV_X1 U6489 ( .A(n6381), .ZN(n5693) );
  AOI22_X1 U6490 ( .A1(n5691), .A2(n5685), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5693), .ZN(n6167) );
  NAND2_X1 U6491 ( .A1(n3646), .A2(n5732), .ZN(n5858) );
  NAND2_X1 U6492 ( .A1(n3646), .A2(n6255), .ZN(n5687) );
  INV_X1 U6493 ( .A(n5917), .ZN(n5688) );
  INV_X1 U6494 ( .A(n6416), .ZN(n5932) );
  OAI22_X1 U6495 ( .A1(n6442), .A2(n5958), .B1(n5932), .B2(n6161), .ZN(n5689)
         );
  AOI21_X1 U6496 ( .B1(n5960), .B2(n6163), .A(n5689), .ZN(n5695) );
  NAND2_X1 U6497 ( .A1(n5691), .A2(n5690), .ZN(n5692) );
  OAI211_X1 U6498 ( .C1(n5925), .C2(n5693), .A(n5692), .B(n5922), .ZN(n6164)
         );
  NAND2_X1 U6499 ( .A1(n6164), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n5694)
         );
  OAI211_X1 U6500 ( .C1(n6167), .C2(n6422), .A(n5695), .B(n5694), .ZN(U3111)
         );
  INV_X1 U6501 ( .A(n6395), .ZN(n5928) );
  OAI22_X1 U6502 ( .A1(n6442), .A2(n5970), .B1(n5928), .B2(n6161), .ZN(n5696)
         );
  AOI21_X1 U6503 ( .B1(n5972), .B2(n6163), .A(n5696), .ZN(n5698) );
  NAND2_X1 U6504 ( .A1(n6164), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n5697)
         );
  OAI211_X1 U6505 ( .C1(n6167), .C2(n6401), .A(n5698), .B(n5697), .ZN(U3115)
         );
  INV_X1 U6506 ( .A(n6409), .ZN(n5918) );
  OAI22_X1 U6507 ( .A1(n6442), .A2(n5952), .B1(n5918), .B2(n6161), .ZN(n5699)
         );
  AOI21_X1 U6508 ( .B1(n5954), .B2(n6163), .A(n5699), .ZN(n5701) );
  NAND2_X1 U6509 ( .A1(n6164), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n5700)
         );
  OAI211_X1 U6510 ( .C1(n6167), .C2(n6415), .A(n5701), .B(n5700), .ZN(U3112)
         );
  INV_X1 U6511 ( .A(n6402), .ZN(n5936) );
  OAI22_X1 U6512 ( .A1(n6442), .A2(n5964), .B1(n5936), .B2(n6161), .ZN(n5702)
         );
  AOI21_X1 U6513 ( .B1(n5966), .B2(n6163), .A(n5702), .ZN(n5704) );
  NAND2_X1 U6514 ( .A1(n6164), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n5703)
         );
  OAI211_X1 U6515 ( .C1(n6167), .C2(n6408), .A(n5704), .B(n5703), .ZN(U3114)
         );
  AOI22_X1 U6516 ( .A1(n5755), .A2(EAX_REG_13__SCAN_IN), .B1(n5705), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n5706) );
  NAND2_X1 U6517 ( .A1(n5707), .A2(n5706), .ZN(U2952) );
  NAND2_X1 U6518 ( .A1(n5708), .A2(DATAI_14_), .ZN(n5712) );
  AOI22_X1 U6519 ( .A1(n5755), .A2(EAX_REG_30__SCAN_IN), .B1(n5705), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n5709) );
  NAND2_X1 U6520 ( .A1(n5712), .A2(n5709), .ZN(U2938) );
  INV_X1 U6521 ( .A(DATAI_12_), .ZN(n6468) );
  OR2_X1 U6522 ( .A1(n6063), .A2(n6468), .ZN(n5722) );
  AOI22_X1 U6523 ( .A1(n5755), .A2(EAX_REG_12__SCAN_IN), .B1(n5705), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n5710) );
  NAND2_X1 U6524 ( .A1(n5722), .A2(n5710), .ZN(U2951) );
  AOI22_X1 U6525 ( .A1(n5755), .A2(EAX_REG_14__SCAN_IN), .B1(n5705), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U6526 ( .A1(n5712), .A2(n5711), .ZN(U2953) );
  AOI22_X1 U6527 ( .A1(n5755), .A2(EAX_REG_11__SCAN_IN), .B1(n5705), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n5713) );
  NAND2_X1 U6528 ( .A1(n5714), .A2(n5713), .ZN(U2950) );
  AOI22_X1 U6529 ( .A1(n5755), .A2(EAX_REG_3__SCAN_IN), .B1(n5705), .B2(
        LWORD_REG_3__SCAN_IN), .ZN(n5715) );
  NAND2_X1 U6530 ( .A1(n5716), .A2(n5715), .ZN(U2942) );
  AOI22_X1 U6531 ( .A1(n5755), .A2(EAX_REG_2__SCAN_IN), .B1(n5705), .B2(
        LWORD_REG_2__SCAN_IN), .ZN(n5717) );
  NAND2_X1 U6532 ( .A1(n5718), .A2(n5717), .ZN(U2941) );
  AOI22_X1 U6533 ( .A1(n5755), .A2(EAX_REG_10__SCAN_IN), .B1(n5705), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n5719) );
  NAND2_X1 U6534 ( .A1(n5720), .A2(n5719), .ZN(U2949) );
  AOI22_X1 U6535 ( .A1(n5755), .A2(EAX_REG_28__SCAN_IN), .B1(n5705), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n5721) );
  NAND2_X1 U6536 ( .A1(n5722), .A2(n5721), .ZN(U2936) );
  AOI22_X1 U6537 ( .A1(n5755), .A2(EAX_REG_9__SCAN_IN), .B1(n5705), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n5723) );
  NAND2_X1 U6538 ( .A1(n5724), .A2(n5723), .ZN(U2948) );
  NOR2_X1 U6539 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5915) );
  NAND2_X1 U6540 ( .A1(n5915), .A2(n7193), .ZN(n5725) );
  NOR2_X1 U6541 ( .A1(n5726), .A2(n5725), .ZN(n6209) );
  NOR2_X1 U6542 ( .A1(n5727), .A2(n5949), .ZN(n5734) );
  AOI21_X1 U6543 ( .B1(n5733), .B2(STATEBS16_REG_SCAN_IN), .A(n5734), .ZN(
        n5728) );
  AOI21_X1 U6544 ( .B1(n5728), .B2(n5838), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n5730) );
  AOI21_X1 U6545 ( .B1(n5915), .B2(n7193), .A(n5838), .ZN(n5735) );
  INV_X1 U6546 ( .A(n5735), .ZN(n5729) );
  OAI211_X1 U6547 ( .C1(n6209), .C2(n5730), .A(n5885), .B(n5729), .ZN(n5731)
         );
  INV_X1 U6548 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n5740) );
  NAND2_X1 U6549 ( .A1(n5733), .A2(n5732), .ZN(n6212) );
  OAI21_X1 U6550 ( .B1(n6209), .B2(n5734), .A(n7724), .ZN(n5736) );
  AOI21_X1 U6551 ( .B1(n5838), .B2(n5736), .A(n5735), .ZN(n6210) );
  AOI22_X1 U6552 ( .A1(n6210), .A2(n6354), .B1(n6416), .B2(n6209), .ZN(n5737)
         );
  OAI21_X1 U6553 ( .B1(n6418), .B2(n6212), .A(n5737), .ZN(n5738) );
  AOI21_X1 U6554 ( .B1(n6420), .B2(n6214), .A(n5738), .ZN(n5739) );
  OAI21_X1 U6555 ( .B1(n6217), .B2(n5740), .A(n5739), .ZN(U3031) );
  INV_X1 U6556 ( .A(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n5744) );
  AOI22_X1 U6557 ( .A1(n6210), .A2(n6344), .B1(n6409), .B2(n6209), .ZN(n5741)
         );
  OAI21_X1 U6558 ( .B1(n6186), .B2(n5952), .A(n5741), .ZN(n5742) );
  AOI21_X1 U6559 ( .B1(n5954), .B2(n6365), .A(n5742), .ZN(n5743) );
  OAI21_X1 U6560 ( .B1(n6217), .B2(n5744), .A(n5743), .ZN(U3032) );
  INV_X1 U6561 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n5748) );
  AOI22_X1 U6562 ( .A1(n6210), .A2(n6329), .B1(n6402), .B2(n6209), .ZN(n5745)
         );
  OAI21_X1 U6563 ( .B1(n6186), .B2(n5964), .A(n5745), .ZN(n5746) );
  AOI21_X1 U6564 ( .B1(n5966), .B2(n6365), .A(n5746), .ZN(n5747) );
  OAI21_X1 U6565 ( .B1(n6217), .B2(n5748), .A(n5747), .ZN(U3034) );
  INV_X1 U6566 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5752) );
  AOI22_X1 U6567 ( .A1(n6210), .A2(n6360), .B1(n6395), .B2(n6209), .ZN(n5749)
         );
  OAI21_X1 U6568 ( .B1(n6186), .B2(n5970), .A(n5749), .ZN(n5750) );
  AOI21_X1 U6569 ( .B1(n5972), .B2(n6365), .A(n5750), .ZN(n5751) );
  OAI21_X1 U6570 ( .B1(n6217), .B2(n5752), .A(n5751), .ZN(U3035) );
  AOI22_X1 U6571 ( .A1(n5755), .A2(EAX_REG_7__SCAN_IN), .B1(n5705), .B2(
        LWORD_REG_7__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U6572 ( .A1(n5754), .A2(n5753), .ZN(U2946) );
  AOI22_X1 U6573 ( .A1(n5755), .A2(EAX_REG_5__SCAN_IN), .B1(n5617), .B2(
        LWORD_REG_5__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U6574 ( .A1(n5757), .A2(n5756), .ZN(U2944) );
  AND3_X1 U6575 ( .A1(n5758), .A2(n5367), .A3(n5803), .ZN(n5759) );
  NAND2_X1 U6576 ( .A1(n5760), .A2(n5759), .ZN(n7168) );
  NAND2_X1 U6577 ( .A1(n3645), .A2(n7168), .ZN(n5776) );
  NAND2_X1 U6578 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5763) );
  NAND2_X1 U6579 ( .A1(n6646), .A2(n5763), .ZN(n5767) );
  NOR2_X1 U6580 ( .A1(n5761), .A2(n3946), .ZN(n5783) );
  INV_X1 U6581 ( .A(n5783), .ZN(n6673) );
  NAND2_X1 U6582 ( .A1(n6673), .A2(n6678), .ZN(n5780) );
  INV_X1 U6583 ( .A(n5762), .ZN(n7164) );
  NAND2_X1 U6584 ( .A1(n7164), .A2(n3720), .ZN(n5765) );
  INV_X1 U6585 ( .A(n5763), .ZN(n5764) );
  AOI22_X1 U6586 ( .A1(n5780), .A2(n5765), .B1(n6646), .B2(n5764), .ZN(n5766)
         );
  MUX2_X1 U6587 ( .A(n5767), .B(n5766), .S(n3751), .Z(n5774) );
  AOI21_X1 U6588 ( .B1(n5762), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n7181), 
        .ZN(n5768) );
  NOR2_X1 U6589 ( .A1(n5769), .A2(n5768), .ZN(n7176) );
  INV_X1 U6590 ( .A(n5423), .ZN(n5772) );
  AND2_X1 U6591 ( .A1(n7164), .A2(n5770), .ZN(n5771) );
  AOI21_X1 U6592 ( .B1(n7176), .B2(n5772), .A(n5771), .ZN(n5773) );
  AND2_X1 U6593 ( .A1(n5774), .A2(n5773), .ZN(n5775) );
  NAND2_X1 U6594 ( .A1(n5776), .A2(n5775), .ZN(n7183) );
  NAND2_X1 U6595 ( .A1(n3663), .A2(n7168), .ZN(n5782) );
  XNOR2_X1 U6596 ( .A(n5762), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5779)
         );
  XNOR2_X1 U6597 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5777) );
  OAI22_X1 U6598 ( .A1(n7188), .A2(n5777), .B1(n5423), .B2(n5779), .ZN(n5778)
         );
  AOI21_X1 U6599 ( .B1(n5780), .B2(n5779), .A(n5778), .ZN(n5781) );
  NAND2_X1 U6600 ( .A1(n5782), .A2(n5781), .ZN(n7185) );
  NAND2_X1 U6601 ( .A1(n5790), .A2(n5783), .ZN(n5787) );
  INV_X1 U6602 ( .A(n5803), .ZN(n5785) );
  NAND2_X1 U6603 ( .A1(n5785), .A2(n5784), .ZN(n5786) );
  NAND2_X1 U6604 ( .A1(n5787), .A2(n5786), .ZN(n6061) );
  NOR2_X1 U6605 ( .A1(n6680), .A2(n6682), .ZN(n5788) );
  OAI22_X1 U6606 ( .A1(n7188), .A2(n7435), .B1(n5788), .B2(n5367), .ZN(n5789)
         );
  NAND3_X1 U6607 ( .A1(n5790), .A2(n7442), .A3(n5789), .ZN(n5792) );
  NAND2_X1 U6608 ( .A1(n5792), .A2(n5791), .ZN(n5793) );
  OR2_X1 U6609 ( .A1(n6061), .A2(n5793), .ZN(n5795) );
  INV_X1 U6610 ( .A(n7190), .ZN(n7184) );
  NAND4_X1 U6611 ( .A1(n7183), .A2(n7715), .A3(n7185), .A4(n7184), .ZN(n5798)
         );
  MUX2_X1 U6612 ( .A(n7702), .B(n7190), .S(n7715), .Z(n5805) );
  NAND2_X1 U6613 ( .A1(n5805), .A2(n5796), .ZN(n5797) );
  NAND2_X1 U6614 ( .A1(n5798), .A2(n5797), .ZN(n7206) );
  INV_X1 U6615 ( .A(n5799), .ZN(n7165) );
  NAND2_X1 U6616 ( .A1(n7206), .A2(n7165), .ZN(n5807) );
  INV_X1 U6617 ( .A(n5865), .ZN(n5800) );
  NOR2_X1 U6618 ( .A1(n5801), .A2(n5800), .ZN(n5802) );
  XNOR2_X1 U6619 ( .A(n5802), .B(n7709), .ZN(n6297) );
  NOR2_X1 U6620 ( .A1(n3630), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U6621 ( .A1(n6297), .A2(n5804), .ZN(n7705) );
  NAND2_X1 U6622 ( .A1(n5805), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5806) );
  NAND2_X1 U6623 ( .A1(n5807), .A2(n7208), .ZN(n7221) );
  NAND2_X1 U6624 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6253), .ZN(n7721) );
  INV_X1 U6625 ( .A(n7721), .ZN(n6642) );
  OAI21_X1 U6626 ( .B1(n7221), .B2(FLUSH_REG_SCAN_IN), .A(n6642), .ZN(n5809)
         );
  OAI21_X1 U6627 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n7715), .A(n6218), .ZN(
        n6260) );
  INV_X1 U6628 ( .A(n3645), .ZN(n6378) );
  NAND2_X1 U6629 ( .A1(n6218), .A2(n5925), .ZN(n6256) );
  INV_X1 U6630 ( .A(n5810), .ZN(n5811) );
  NAND2_X1 U6631 ( .A1(n5811), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5814) );
  AOI211_X1 U6632 ( .C1(n3640), .C2(n5814), .A(n5813), .B(n5812), .ZN(n5815)
         );
  OAI222_X1 U6633 ( .A1(n6260), .A2(n6378), .B1(n6218), .B2(n7198), .C1(n6256), 
        .C2(n5815), .ZN(U3462) );
  INV_X1 U6634 ( .A(n6114), .ZN(n5816) );
  AOI21_X1 U6635 ( .B1(n5816), .B2(n6117), .A(n7726), .ZN(n5817) );
  AOI211_X1 U6636 ( .C1(n5870), .C2(n5865), .A(n6375), .B(n5817), .ZN(n5820)
         );
  NOR2_X1 U6637 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5818), .ZN(n5821)
         );
  NAND2_X1 U6638 ( .A1(n5861), .A2(n5837), .ZN(n5948) );
  NAND2_X1 U6639 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5948), .ZN(n5944) );
  OAI21_X1 U6640 ( .B1(n5821), .B2(n7724), .A(n5944), .ZN(n5819) );
  NAND2_X1 U6641 ( .A1(n6110), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5825)
         );
  INV_X1 U6642 ( .A(n5821), .ZN(n6112) );
  INV_X1 U6643 ( .A(n5948), .ZN(n5822) );
  INV_X1 U6644 ( .A(n5884), .ZN(n5869) );
  AOI22_X1 U6645 ( .A1(n5845), .A2(n5870), .B1(n5822), .B2(n5869), .ZN(n6111)
         );
  OAI22_X1 U6646 ( .A1(n5932), .A2(n6112), .B1(n6111), .B2(n6422), .ZN(n5823)
         );
  AOI21_X1 U6647 ( .B1(n5960), .B2(n6114), .A(n5823), .ZN(n5824) );
  OAI211_X1 U6648 ( .C1(n6117), .C2(n5958), .A(n5825), .B(n5824), .ZN(U3119)
         );
  NAND2_X1 U6649 ( .A1(n6110), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5828)
         );
  OAI22_X1 U6650 ( .A1(n5936), .A2(n6112), .B1(n6111), .B2(n6408), .ZN(n5826)
         );
  AOI21_X1 U6651 ( .B1(n5966), .B2(n6114), .A(n5826), .ZN(n5827) );
  OAI211_X1 U6652 ( .C1(n6117), .C2(n5964), .A(n5828), .B(n5827), .ZN(U3122)
         );
  NAND2_X1 U6653 ( .A1(n6110), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5831)
         );
  OAI22_X1 U6654 ( .A1(n5918), .A2(n6112), .B1(n6111), .B2(n6415), .ZN(n5829)
         );
  AOI21_X1 U6655 ( .B1(n5954), .B2(n6114), .A(n5829), .ZN(n5830) );
  OAI211_X1 U6656 ( .C1(n6117), .C2(n5952), .A(n5831), .B(n5830), .ZN(U3120)
         );
  NAND2_X1 U6657 ( .A1(n6110), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5834)
         );
  OAI22_X1 U6658 ( .A1(n5928), .A2(n6112), .B1(n6111), .B2(n6401), .ZN(n5832)
         );
  AOI21_X1 U6659 ( .B1(n5972), .B2(n6114), .A(n5832), .ZN(n5833) );
  OAI211_X1 U6660 ( .C1(n6117), .C2(n5970), .A(n5834), .B(n5833), .ZN(U3123)
         );
  AOI22_X1 U6661 ( .A1(n5755), .A2(EAX_REG_15__SCAN_IN), .B1(n5617), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n5835) );
  OAI21_X1 U6662 ( .B1(n6063), .B2(n6950), .A(n5835), .ZN(U2954) );
  OR2_X1 U6663 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5836), .ZN(n6138)
         );
  NOR2_X1 U6664 ( .A1(n5837), .A2(n7198), .ZN(n6379) );
  NOR2_X1 U6665 ( .A1(n6379), .A2(n5838), .ZN(n6383) );
  AOI211_X1 U6666 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6138), .A(n6383), .B(
        n5862), .ZN(n5843) );
  INV_X1 U6667 ( .A(n6323), .ZN(n5871) );
  INV_X1 U6668 ( .A(n6143), .ZN(n5839) );
  OAI21_X1 U6669 ( .B1(n5839), .B2(n6140), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5840) );
  OAI21_X1 U6670 ( .B1(n5871), .B2(n5841), .A(n5840), .ZN(n5842) );
  NAND2_X1 U6671 ( .A1(n5843), .A2(n5842), .ZN(n6136) );
  NAND2_X1 U6672 ( .A1(n6136), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5848)
         );
  AOI22_X1 U6673 ( .A1(n5845), .A2(n5844), .B1(n6379), .B2(n5869), .ZN(n6137)
         );
  OAI22_X1 U6674 ( .A1(n5928), .A2(n6138), .B1(n6137), .B2(n6401), .ZN(n5846)
         );
  AOI21_X1 U6675 ( .B1(n5972), .B2(n6140), .A(n5846), .ZN(n5847) );
  OAI211_X1 U6676 ( .C1(n6143), .C2(n5970), .A(n5848), .B(n5847), .ZN(U3139)
         );
  NAND2_X1 U6677 ( .A1(n6136), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5851)
         );
  OAI22_X1 U6678 ( .A1(n5936), .A2(n6138), .B1(n6137), .B2(n6408), .ZN(n5849)
         );
  AOI21_X1 U6679 ( .B1(n5966), .B2(n6140), .A(n5849), .ZN(n5850) );
  OAI211_X1 U6680 ( .C1(n6143), .C2(n5964), .A(n5851), .B(n5850), .ZN(U3138)
         );
  NAND2_X1 U6681 ( .A1(n6136), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5854)
         );
  OAI22_X1 U6682 ( .A1(n5918), .A2(n6138), .B1(n6137), .B2(n6415), .ZN(n5852)
         );
  AOI21_X1 U6683 ( .B1(n5954), .B2(n6140), .A(n5852), .ZN(n5853) );
  OAI211_X1 U6684 ( .C1(n6143), .C2(n5952), .A(n5854), .B(n5853), .ZN(U3136)
         );
  NAND2_X1 U6685 ( .A1(n6136), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5857)
         );
  OAI22_X1 U6686 ( .A1(n5932), .A2(n6138), .B1(n6137), .B2(n6422), .ZN(n5855)
         );
  AOI21_X1 U6687 ( .B1(n5960), .B2(n6140), .A(n5855), .ZN(n5856) );
  OAI211_X1 U6688 ( .C1(n6143), .C2(n5958), .A(n5857), .B(n5856), .ZN(U3135)
         );
  OR2_X1 U6689 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5859), .ZN(n6146)
         );
  OR2_X1 U6690 ( .A1(n5861), .A2(n5860), .ZN(n5868) );
  AND2_X1 U6691 ( .A1(n5868), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5886) );
  AOI211_X1 U6692 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6146), .A(n5886), .B(
        n5862), .ZN(n5867) );
  OAI21_X1 U6693 ( .B1(n6195), .B2(n6148), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5863) );
  OAI211_X1 U6694 ( .C1(n5865), .C2(n5864), .A(n5863), .B(n5925), .ZN(n5866)
         );
  NAND2_X1 U6695 ( .A1(n5867), .A2(n5866), .ZN(n6144) );
  NAND2_X1 U6696 ( .A1(n6144), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5874) );
  INV_X1 U6697 ( .A(n5868), .ZN(n5891) );
  AOI22_X1 U6698 ( .A1(n5871), .A2(n5870), .B1(n5891), .B2(n5869), .ZN(n6145)
         );
  OAI22_X1 U6699 ( .A1(n5932), .A2(n6146), .B1(n6145), .B2(n6422), .ZN(n5872)
         );
  AOI21_X1 U6700 ( .B1(n5960), .B2(n6148), .A(n5872), .ZN(n5873) );
  OAI211_X1 U6701 ( .C1(n6151), .C2(n5958), .A(n5874), .B(n5873), .ZN(U3055)
         );
  NAND2_X1 U6702 ( .A1(n6144), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5877) );
  OAI22_X1 U6703 ( .A1(n5928), .A2(n6146), .B1(n6145), .B2(n6401), .ZN(n5875)
         );
  AOI21_X1 U6704 ( .B1(n5972), .B2(n6148), .A(n5875), .ZN(n5876) );
  OAI211_X1 U6705 ( .C1(n6151), .C2(n5970), .A(n5877), .B(n5876), .ZN(U3059)
         );
  NAND2_X1 U6706 ( .A1(n6144), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5880) );
  OAI22_X1 U6707 ( .A1(n5936), .A2(n6146), .B1(n6145), .B2(n6408), .ZN(n5878)
         );
  AOI21_X1 U6708 ( .B1(n5966), .B2(n6148), .A(n5878), .ZN(n5879) );
  OAI211_X1 U6709 ( .C1(n6151), .C2(n5964), .A(n5880), .B(n5879), .ZN(U3058)
         );
  NAND2_X1 U6710 ( .A1(n6144), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5883) );
  OAI22_X1 U6711 ( .A1(n5918), .A2(n6146), .B1(n6145), .B2(n6415), .ZN(n5881)
         );
  AOI21_X1 U6712 ( .B1(n5954), .B2(n6148), .A(n5881), .ZN(n5882) );
  OAI211_X1 U6713 ( .C1(n6151), .C2(n5952), .A(n5883), .B(n5882), .ZN(U3056)
         );
  AOI21_X1 U6714 ( .B1(n6186), .B2(n6047), .A(n7726), .ZN(n5889) );
  NAND2_X1 U6715 ( .A1(n5949), .A2(n5925), .ZN(n5941) );
  AND2_X1 U6716 ( .A1(n5950), .A2(n5941), .ZN(n5888) );
  NAND2_X1 U6717 ( .A1(n5943), .A2(n5915), .ZN(n5890) );
  AOI211_X1 U6718 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5890), .A(n5886), .B(
        n6384), .ZN(n5887) );
  NAND2_X1 U6719 ( .A1(n6214), .A2(n5960), .ZN(n5894) );
  INV_X1 U6720 ( .A(n5890), .ZN(n5998) );
  INV_X1 U6721 ( .A(n6322), .ZN(n6380) );
  NAND2_X1 U6722 ( .A1(n5891), .A2(n6380), .ZN(n5892) );
  OAI21_X1 U6723 ( .B1(n6323), .B2(n5949), .A(n5892), .ZN(n5997) );
  AOI22_X1 U6724 ( .A1(n6416), .A2(n5998), .B1(n6354), .B2(n5997), .ZN(n5893)
         );
  OAI211_X1 U6725 ( .C1(n6047), .C2(n5958), .A(n5894), .B(n5893), .ZN(n5895)
         );
  AOI21_X1 U6726 ( .B1(n6002), .B2(INSTQUEUE_REG_0__3__SCAN_IN), .A(n5895), 
        .ZN(n5896) );
  INV_X1 U6727 ( .A(n5896), .ZN(U3023) );
  NAND2_X1 U6728 ( .A1(n6214), .A2(n5966), .ZN(n5898) );
  AOI22_X1 U6729 ( .A1(n6402), .A2(n5998), .B1(n6329), .B2(n5997), .ZN(n5897)
         );
  OAI211_X1 U6730 ( .C1(n6047), .C2(n5964), .A(n5898), .B(n5897), .ZN(n5899)
         );
  AOI21_X1 U6731 ( .B1(n6002), .B2(INSTQUEUE_REG_0__6__SCAN_IN), .A(n5899), 
        .ZN(n5900) );
  INV_X1 U6732 ( .A(n5900), .ZN(U3026) );
  NAND2_X1 U6733 ( .A1(n6214), .A2(n5954), .ZN(n5902) );
  AOI22_X1 U6734 ( .A1(n6409), .A2(n5998), .B1(n6344), .B2(n5997), .ZN(n5901)
         );
  OAI211_X1 U6735 ( .C1(n6047), .C2(n5952), .A(n5902), .B(n5901), .ZN(n5903)
         );
  AOI21_X1 U6736 ( .B1(n6002), .B2(INSTQUEUE_REG_0__4__SCAN_IN), .A(n5903), 
        .ZN(n5904) );
  INV_X1 U6737 ( .A(n5904), .ZN(U3024) );
  NAND2_X1 U6738 ( .A1(n6214), .A2(n5972), .ZN(n5906) );
  AOI22_X1 U6739 ( .A1(n6395), .A2(n5998), .B1(n6360), .B2(n5997), .ZN(n5905)
         );
  OAI211_X1 U6740 ( .C1(n6047), .C2(n5970), .A(n5906), .B(n5905), .ZN(n5907)
         );
  AOI21_X1 U6741 ( .B1(n6002), .B2(INSTQUEUE_REG_0__7__SCAN_IN), .A(n5907), 
        .ZN(n5908) );
  INV_X1 U6742 ( .A(n5908), .ZN(U3027) );
  INV_X1 U6743 ( .A(n5909), .ZN(n5910) );
  AOI21_X1 U6744 ( .B1(n5910), .B2(n5975), .A(n6375), .ZN(n5921) );
  NAND2_X1 U6745 ( .A1(n5911), .A2(n5915), .ZN(n6191) );
  INV_X1 U6746 ( .A(n6191), .ZN(n5912) );
  AOI21_X1 U6747 ( .B1(n5914), .B2(n5913), .A(n5912), .ZN(n5920) );
  INV_X1 U6748 ( .A(n5920), .ZN(n5916) );
  NAND2_X1 U6749 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n5915), .ZN(n6316) );
  INV_X1 U6750 ( .A(n6316), .ZN(n5924) );
  AOI22_X1 U6751 ( .A1(n5921), .A2(n5916), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5924), .ZN(n6200) );
  NOR2_X1 U6752 ( .A1(n3640), .A2(n5917), .ZN(n6314) );
  OAI22_X1 U6753 ( .A1(n6363), .A2(n5952), .B1(n5918), .B2(n6191), .ZN(n5919)
         );
  AOI21_X1 U6754 ( .B1(n5954), .B2(n6195), .A(n5919), .ZN(n5927) );
  NAND2_X1 U6755 ( .A1(n5921), .A2(n5920), .ZN(n5923) );
  OAI211_X1 U6756 ( .C1(n5925), .C2(n5924), .A(n5923), .B(n5922), .ZN(n6197)
         );
  NAND2_X1 U6757 ( .A1(n6197), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n5926) );
  OAI211_X1 U6758 ( .C1(n6200), .C2(n6415), .A(n5927), .B(n5926), .ZN(U3048)
         );
  OAI22_X1 U6759 ( .A1(n6363), .A2(n5970), .B1(n5928), .B2(n6191), .ZN(n5929)
         );
  AOI21_X1 U6760 ( .B1(n5972), .B2(n6195), .A(n5929), .ZN(n5931) );
  NAND2_X1 U6761 ( .A1(n6197), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5930) );
  OAI211_X1 U6762 ( .C1(n6200), .C2(n6401), .A(n5931), .B(n5930), .ZN(U3051)
         );
  OAI22_X1 U6763 ( .A1(n6363), .A2(n5958), .B1(n5932), .B2(n6191), .ZN(n5933)
         );
  AOI21_X1 U6764 ( .B1(n5960), .B2(n6195), .A(n5933), .ZN(n5935) );
  NAND2_X1 U6765 ( .A1(n6197), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n5934) );
  OAI211_X1 U6766 ( .C1(n6200), .C2(n6422), .A(n5935), .B(n5934), .ZN(U3047)
         );
  OAI22_X1 U6767 ( .A1(n6363), .A2(n5964), .B1(n5936), .B2(n6191), .ZN(n5937)
         );
  AOI21_X1 U6768 ( .B1(n5966), .B2(n6195), .A(n5937), .ZN(n5939) );
  NAND2_X1 U6769 ( .A1(n6197), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5938) );
  OAI211_X1 U6770 ( .C1(n6200), .C2(n6408), .A(n5939), .B(n5938), .ZN(U3050)
         );
  AOI21_X1 U6771 ( .B1(n5947), .B2(n6095), .A(n7726), .ZN(n5940) );
  AOI21_X1 U6772 ( .B1(n6323), .B2(n5941), .A(n5940), .ZN(n5946) );
  AND2_X1 U6773 ( .A1(n5943), .A2(n5942), .ZN(n6093) );
  OAI21_X1 U6774 ( .B1(n7724), .B2(n6093), .A(n5944), .ZN(n5945) );
  NOR3_X2 U6775 ( .A1(n5946), .A2(n6384), .A3(n5945), .ZN(n6100) );
  INV_X1 U6776 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5956) );
  OAI22_X1 U6777 ( .A1(n5950), .A2(n5949), .B1(n6322), .B2(n5948), .ZN(n6092)
         );
  AOI22_X1 U6778 ( .A1(n6409), .A2(n6093), .B1(n6344), .B2(n6092), .ZN(n5951)
         );
  OAI21_X1 U6779 ( .B1(n5952), .B2(n6095), .A(n5951), .ZN(n5953) );
  AOI21_X1 U6780 ( .B1(n6097), .B2(n5954), .A(n5953), .ZN(n5955) );
  OAI21_X1 U6781 ( .B1(n6100), .B2(n5956), .A(n5955), .ZN(U3088) );
  INV_X1 U6782 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5962) );
  AOI22_X1 U6783 ( .A1(n6416), .A2(n6093), .B1(n6354), .B2(n6092), .ZN(n5957)
         );
  OAI21_X1 U6784 ( .B1(n5958), .B2(n6095), .A(n5957), .ZN(n5959) );
  AOI21_X1 U6785 ( .B1(n6097), .B2(n5960), .A(n5959), .ZN(n5961) );
  OAI21_X1 U6786 ( .B1(n6100), .B2(n5962), .A(n5961), .ZN(U3087) );
  INV_X1 U6787 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5968) );
  AOI22_X1 U6788 ( .A1(n6402), .A2(n6093), .B1(n6329), .B2(n6092), .ZN(n5963)
         );
  OAI21_X1 U6789 ( .B1(n5964), .B2(n6095), .A(n5963), .ZN(n5965) );
  AOI21_X1 U6790 ( .B1(n6097), .B2(n5966), .A(n5965), .ZN(n5967) );
  OAI21_X1 U6791 ( .B1(n6100), .B2(n5968), .A(n5967), .ZN(U3090) );
  INV_X1 U6792 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5974) );
  AOI22_X1 U6793 ( .A1(n6395), .A2(n6093), .B1(n6360), .B2(n6092), .ZN(n5969)
         );
  OAI21_X1 U6794 ( .B1(n5970), .B2(n6095), .A(n5969), .ZN(n5971) );
  AOI21_X1 U6795 ( .B1(n6097), .B2(n5972), .A(n5971), .ZN(n5973) );
  OAI21_X1 U6796 ( .B1(n6100), .B2(n5974), .A(n5973), .ZN(U3091) );
  INV_X1 U6797 ( .A(n3663), .ZN(n5977) );
  XNOR2_X1 U6798 ( .A(n5975), .B(n3662), .ZN(n5976) );
  OAI222_X1 U6799 ( .A1(n6218), .A2(n4099), .B1(n6260), .B2(n5977), .C1(n6256), 
        .C2(n5976), .ZN(U3463) );
  OAI21_X1 U6800 ( .B1(n7530), .B2(n7473), .A(n7469), .ZN(n7452) );
  OAI21_X1 U6801 ( .B1(n7555), .B2(n6862), .A(n5978), .ZN(n5982) );
  OAI21_X1 U6802 ( .B1(n7474), .B2(n5979), .A(n7530), .ZN(n7461) );
  NAND2_X1 U6803 ( .A1(n7461), .A2(n7473), .ZN(n5980) );
  NOR2_X1 U6804 ( .A1(n5980), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n5981)
         );
  AOI211_X1 U6805 ( .C1(n7452), .C2(INSTADDRPOINTER_REG_3__SCAN_IN), .A(n5982), 
        .B(n5981), .ZN(n5983) );
  OAI21_X1 U6806 ( .B1(n5984), .B2(n7506), .A(n5983), .ZN(U3015) );
  NAND2_X1 U6807 ( .A1(n6214), .A2(n6181), .ZN(n5986) );
  AOI22_X1 U6808 ( .A1(n6430), .A2(n5998), .B1(n6339), .B2(n5997), .ZN(n5985)
         );
  OAI211_X1 U6809 ( .C1(n6047), .C2(n6179), .A(n5986), .B(n5985), .ZN(n5987)
         );
  AOI21_X1 U6810 ( .B1(n6002), .B2(INSTQUEUE_REG_0__2__SCAN_IN), .A(n5987), 
        .ZN(n5988) );
  INV_X1 U6811 ( .A(n5988), .ZN(U3022) );
  NAND2_X1 U6812 ( .A1(n6214), .A2(n6175), .ZN(n5990) );
  AOI22_X1 U6813 ( .A1(n3678), .A2(n5998), .B1(n6349), .B2(n5997), .ZN(n5989)
         );
  OAI211_X1 U6814 ( .C1(n6047), .C2(n6173), .A(n5990), .B(n5989), .ZN(n5991)
         );
  AOI21_X1 U6815 ( .B1(n6002), .B2(INSTQUEUE_REG_0__1__SCAN_IN), .A(n5991), 
        .ZN(n5992) );
  INV_X1 U6816 ( .A(n5992), .ZN(U3021) );
  NAND2_X1 U6817 ( .A1(n6214), .A2(n6196), .ZN(n5994) );
  AOI22_X1 U6818 ( .A1(n6439), .A2(n5998), .B1(n6324), .B2(n5997), .ZN(n5993)
         );
  OAI211_X1 U6819 ( .C1(n6047), .C2(n6193), .A(n5994), .B(n5993), .ZN(n5995)
         );
  AOI21_X1 U6820 ( .B1(n6002), .B2(INSTQUEUE_REG_0__0__SCAN_IN), .A(n5995), 
        .ZN(n5996) );
  INV_X1 U6821 ( .A(n5996), .ZN(U3020) );
  NAND2_X1 U6822 ( .A1(n6214), .A2(n6188), .ZN(n6000) );
  AOI22_X1 U6823 ( .A1(n7767), .A2(n5998), .B1(n6334), .B2(n5997), .ZN(n5999)
         );
  OAI211_X1 U6824 ( .C1(n6047), .C2(n6185), .A(n6000), .B(n5999), .ZN(n6001)
         );
  AOI21_X1 U6825 ( .B1(n6002), .B2(INSTQUEUE_REG_0__5__SCAN_IN), .A(n6001), 
        .ZN(n6003) );
  INV_X1 U6826 ( .A(n6003), .ZN(U3025) );
  AND2_X1 U6827 ( .A1(n5521), .A2(n6004), .ZN(n6006) );
  OR2_X1 U6828 ( .A1(n6006), .A2(n6005), .ZN(n7605) );
  INV_X1 U6829 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6010) );
  NOR2_X1 U6830 ( .A1(n5526), .A2(n6008), .ZN(n6009) );
  OR2_X1 U6831 ( .A1(n6007), .A2(n6009), .ZN(n6224) );
  OAI222_X1 U6832 ( .A1(n7605), .A2(n6919), .B1(n7369), .B2(n6010), .C1(n6224), 
        .C2(n6917), .ZN(U2851) );
  INV_X1 U6833 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n6014) );
  AOI22_X1 U6834 ( .A1(n6423), .A2(n6024), .B1(n6349), .B2(n6023), .ZN(n6011)
         );
  OAI21_X1 U6835 ( .B1(n6173), .B2(n6026), .A(n6011), .ZN(n6012) );
  AOI21_X1 U6836 ( .B1(n6175), .B2(n6028), .A(n6012), .ZN(n6013) );
  OAI21_X1 U6837 ( .B1(n6031), .B2(n6014), .A(n6013), .ZN(U3069) );
  INV_X1 U6838 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n6018) );
  AOI22_X1 U6839 ( .A1(n6430), .A2(n6024), .B1(n6339), .B2(n6023), .ZN(n6015)
         );
  OAI21_X1 U6840 ( .B1(n6179), .B2(n6026), .A(n6015), .ZN(n6016) );
  AOI21_X1 U6841 ( .B1(n6181), .B2(n6028), .A(n6016), .ZN(n6017) );
  OAI21_X1 U6842 ( .B1(n6031), .B2(n6018), .A(n6017), .ZN(U3070) );
  INV_X1 U6843 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n6022) );
  AOI22_X1 U6844 ( .A1(n6439), .A2(n6024), .B1(n6324), .B2(n6023), .ZN(n6019)
         );
  OAI21_X1 U6845 ( .B1(n6193), .B2(n6026), .A(n6019), .ZN(n6020) );
  AOI21_X1 U6846 ( .B1(n6196), .B2(n6028), .A(n6020), .ZN(n6021) );
  OAI21_X1 U6847 ( .B1(n6031), .B2(n6022), .A(n6021), .ZN(U3068) );
  INV_X1 U6848 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n6030) );
  AOI22_X1 U6849 ( .A1(n6388), .A2(n6024), .B1(n6334), .B2(n6023), .ZN(n6025)
         );
  OAI21_X1 U6850 ( .B1(n6185), .B2(n6026), .A(n6025), .ZN(n6027) );
  AOI21_X1 U6851 ( .B1(n6188), .B2(n6028), .A(n6027), .ZN(n6029) );
  OAI21_X1 U6852 ( .B1(n6031), .B2(n6030), .A(n6029), .ZN(U3073) );
  INV_X1 U6853 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n6035) );
  AOI22_X1 U6854 ( .A1(n6388), .A2(n6045), .B1(n6334), .B2(n6044), .ZN(n6032)
         );
  OAI21_X1 U6855 ( .B1(n6390), .B2(n6047), .A(n6032), .ZN(n6033) );
  AOI21_X1 U6856 ( .B1(n6392), .B2(n6140), .A(n6033), .ZN(n6034) );
  OAI21_X1 U6857 ( .B1(n6051), .B2(n6035), .A(n6034), .ZN(U3145) );
  INV_X1 U6858 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n6039) );
  AOI22_X1 U6859 ( .A1(n6423), .A2(n6045), .B1(n6349), .B2(n6044), .ZN(n6036)
         );
  OAI21_X1 U6860 ( .B1(n6425), .B2(n6047), .A(n6036), .ZN(n6037) );
  AOI21_X1 U6861 ( .B1(n6427), .B2(n6140), .A(n6037), .ZN(n6038) );
  OAI21_X1 U6862 ( .B1(n6051), .B2(n6039), .A(n6038), .ZN(U3141) );
  INV_X1 U6863 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n6043) );
  AOI22_X1 U6864 ( .A1(n6430), .A2(n6045), .B1(n6339), .B2(n6044), .ZN(n6040)
         );
  OAI21_X1 U6865 ( .B1(n6432), .B2(n6047), .A(n6040), .ZN(n6041) );
  AOI21_X1 U6866 ( .B1(n6434), .B2(n6140), .A(n6041), .ZN(n6042) );
  OAI21_X1 U6867 ( .B1(n6051), .B2(n6043), .A(n6042), .ZN(U3142) );
  INV_X1 U6868 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n6050) );
  AOI22_X1 U6869 ( .A1(n6439), .A2(n6045), .B1(n6324), .B2(n6044), .ZN(n6046)
         );
  OAI21_X1 U6870 ( .B1(n6441), .B2(n6047), .A(n6046), .ZN(n6048) );
  AOI21_X1 U6871 ( .B1(n6445), .B2(n6140), .A(n6048), .ZN(n6049) );
  OAI21_X1 U6872 ( .B1(n6051), .B2(n6050), .A(n6049), .ZN(U3140) );
  XNOR2_X1 U6873 ( .A(n3676), .B(n6052), .ZN(n7399) );
  INV_X1 U6874 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n7466) );
  NOR3_X1 U6875 ( .A1(n7466), .A2(n7460), .A3(n7459), .ZN(n6478) );
  NOR3_X1 U6876 ( .A1(n7466), .A2(n7460), .A3(n6053), .ZN(n6474) );
  INV_X1 U6877 ( .A(n6474), .ZN(n6054) );
  AOI21_X1 U6878 ( .B1(n7528), .B2(n6054), .A(n7526), .ZN(n6270) );
  OAI21_X1 U6879 ( .B1(n6478), .B2(n7530), .A(n6270), .ZN(n6271) );
  NAND2_X1 U6880 ( .A1(n6478), .A2(n7461), .ZN(n6273) );
  NAND2_X1 U6881 ( .A1(n7585), .A2(n7545), .ZN(n6056) );
  INV_X1 U6882 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6055) );
  OR2_X1 U6883 ( .A1(n7524), .A2(n6055), .ZN(n7402) );
  OAI211_X1 U6884 ( .C1(n6273), .C2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6056), 
        .B(n7402), .ZN(n6057) );
  AOI21_X1 U6885 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n6271), .A(n6057), 
        .ZN(n6058) );
  OAI21_X1 U6886 ( .B1(n7399), .B2(n7506), .A(n6058), .ZN(U3011) );
  NOR2_X1 U6887 ( .A1(n5758), .A2(n6059), .ZN(n6060) );
  NAND2_X1 U6888 ( .A1(n6064), .A2(n3933), .ZN(n6065) );
  AND2_X1 U6889 ( .A1(n6952), .A2(n6066), .ZN(n7759) );
  AND2_X1 U6890 ( .A1(n6067), .A2(n3933), .ZN(n6068) );
  OAI222_X1 U6891 ( .A1(n6070), .A2(n7751), .B1(n6953), .B2(n6069), .C1(n6952), 
        .C2(n4329), .ZN(U2884) );
  INV_X1 U6892 ( .A(EAX_REG_1__SCAN_IN), .ZN(n7259) );
  OAI222_X1 U6893 ( .A1(n7370), .A2(n7751), .B1(n6953), .B2(n6071), .C1(n6952), 
        .C2(n7259), .ZN(U2890) );
  INV_X1 U6894 ( .A(EAX_REG_0__SCAN_IN), .ZN(n7257) );
  OAI222_X1 U6895 ( .A1(n6952), .A2(n7257), .B1(n7751), .B2(n6312), .C1(n6072), 
        .C2(n6953), .ZN(U2891) );
  INV_X1 U6896 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n6076) );
  AOI22_X1 U6897 ( .A1(n6423), .A2(n6093), .B1(n6349), .B2(n6092), .ZN(n6073)
         );
  OAI21_X1 U6898 ( .B1(n6173), .B2(n6095), .A(n6073), .ZN(n6074) );
  AOI21_X1 U6899 ( .B1(n6097), .B2(n6175), .A(n6074), .ZN(n6075) );
  OAI21_X1 U6900 ( .B1(n6100), .B2(n6076), .A(n6075), .ZN(U3085) );
  INV_X1 U6901 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n6080) );
  AOI22_X1 U6902 ( .A1(n6430), .A2(n6093), .B1(n6339), .B2(n6092), .ZN(n6077)
         );
  OAI21_X1 U6903 ( .B1(n6179), .B2(n6095), .A(n6077), .ZN(n6078) );
  AOI21_X1 U6904 ( .B1(n6097), .B2(n6181), .A(n6078), .ZN(n6079) );
  OAI21_X1 U6905 ( .B1(n6100), .B2(n6080), .A(n6079), .ZN(U3086) );
  INV_X1 U6906 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n6084) );
  AOI22_X1 U6907 ( .A1(n6439), .A2(n6093), .B1(n6324), .B2(n6092), .ZN(n6081)
         );
  OAI21_X1 U6908 ( .B1(n6193), .B2(n6095), .A(n6081), .ZN(n6082) );
  AOI21_X1 U6909 ( .B1(n6097), .B2(n6196), .A(n6082), .ZN(n6083) );
  OAI21_X1 U6910 ( .B1(n6100), .B2(n6084), .A(n6083), .ZN(U3084) );
  INV_X1 U6911 ( .A(EAX_REG_2__SCAN_IN), .ZN(n7261) );
  OAI222_X1 U6912 ( .A1(n6880), .A2(n7751), .B1(n6085), .B2(n6953), .C1(n6952), 
        .C2(n7261), .ZN(U2889) );
  OAI222_X1 U6913 ( .A1(n6087), .A2(n7751), .B1(n6086), .B2(n6953), .C1(n7269), 
        .C2(n6952), .ZN(U2885) );
  INV_X1 U6914 ( .A(EAX_REG_3__SCAN_IN), .ZN(n7263) );
  OAI222_X1 U6915 ( .A1(n6089), .A2(n7751), .B1(n6088), .B2(n6953), .C1(n6952), 
        .C2(n7263), .ZN(U2888) );
  INV_X1 U6916 ( .A(n7570), .ZN(n6090) );
  INV_X1 U6917 ( .A(EAX_REG_5__SCAN_IN), .ZN(n7267) );
  OAI222_X1 U6918 ( .A1(n6090), .A2(n7751), .B1(n6944), .B2(n6953), .C1(n6952), 
        .C2(n7267), .ZN(U2886) );
  INV_X1 U6919 ( .A(EAX_REG_4__SCAN_IN), .ZN(n7265) );
  OAI222_X1 U6920 ( .A1(n6293), .A2(n7751), .B1(n6091), .B2(n6953), .C1(n7265), 
        .C2(n6952), .ZN(U2887) );
  INV_X1 U6921 ( .A(EAX_REG_8__SCAN_IN), .ZN(n7272) );
  OAI222_X1 U6922 ( .A1(n7605), .A2(n7751), .B1(n6936), .B2(n6953), .C1(n6952), 
        .C2(n7272), .ZN(U2883) );
  INV_X1 U6923 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n6099) );
  AOI22_X1 U6924 ( .A1(n6388), .A2(n6093), .B1(n6334), .B2(n6092), .ZN(n6094)
         );
  OAI21_X1 U6925 ( .B1(n6185), .B2(n6095), .A(n6094), .ZN(n6096) );
  AOI21_X1 U6926 ( .B1(n6097), .B2(n6188), .A(n6096), .ZN(n6098) );
  OAI21_X1 U6927 ( .B1(n6100), .B2(n6099), .A(n6098), .ZN(U3089) );
  NAND2_X1 U6928 ( .A1(n6110), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n6103)
         );
  INV_X1 U6929 ( .A(n6430), .ZN(n6178) );
  OAI22_X1 U6930 ( .A1(n6178), .A2(n6112), .B1(n6111), .B2(n6436), .ZN(n6101)
         );
  AOI21_X1 U6931 ( .B1(n6181), .B2(n6114), .A(n6101), .ZN(n6102) );
  OAI211_X1 U6932 ( .C1(n6117), .C2(n6179), .A(n6103), .B(n6102), .ZN(U3118)
         );
  NAND2_X1 U6933 ( .A1(n6110), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n6106)
         );
  INV_X1 U6934 ( .A(n6388), .ZN(n6168) );
  OAI22_X1 U6935 ( .A1(n6168), .A2(n6112), .B1(n6111), .B2(n6394), .ZN(n6104)
         );
  AOI21_X1 U6936 ( .B1(n6188), .B2(n6114), .A(n6104), .ZN(n6105) );
  OAI211_X1 U6937 ( .C1(n6117), .C2(n6185), .A(n6106), .B(n6105), .ZN(U3121)
         );
  NAND2_X1 U6938 ( .A1(n6110), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n6109)
         );
  INV_X1 U6939 ( .A(n6423), .ZN(n6172) );
  OAI22_X1 U6940 ( .A1(n6172), .A2(n6112), .B1(n6111), .B2(n6429), .ZN(n6107)
         );
  AOI21_X1 U6941 ( .B1(n6175), .B2(n6114), .A(n6107), .ZN(n6108) );
  OAI211_X1 U6942 ( .C1(n6117), .C2(n6173), .A(n6109), .B(n6108), .ZN(U3117)
         );
  NAND2_X1 U6943 ( .A1(n6110), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n6116)
         );
  INV_X1 U6944 ( .A(n6439), .ZN(n6192) );
  OAI22_X1 U6945 ( .A1(n6192), .A2(n6112), .B1(n6111), .B2(n6447), .ZN(n6113)
         );
  AOI21_X1 U6946 ( .B1(n6196), .B2(n6114), .A(n6113), .ZN(n6115) );
  OAI211_X1 U6947 ( .C1(n6117), .C2(n6193), .A(n6116), .B(n6115), .ZN(U3116)
         );
  NAND2_X1 U6948 ( .A1(n6136), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n6120)
         );
  OAI22_X1 U6949 ( .A1(n6168), .A2(n6138), .B1(n6137), .B2(n6394), .ZN(n6118)
         );
  AOI21_X1 U6950 ( .B1(n6188), .B2(n6140), .A(n6118), .ZN(n6119) );
  OAI211_X1 U6951 ( .C1(n6143), .C2(n6185), .A(n6120), .B(n6119), .ZN(U3137)
         );
  NAND2_X1 U6952 ( .A1(n6136), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n6123)
         );
  OAI22_X1 U6953 ( .A1(n6172), .A2(n6138), .B1(n6137), .B2(n6429), .ZN(n6121)
         );
  AOI21_X1 U6954 ( .B1(n6175), .B2(n6140), .A(n6121), .ZN(n6122) );
  OAI211_X1 U6955 ( .C1(n6143), .C2(n6173), .A(n6123), .B(n6122), .ZN(U3133)
         );
  NAND2_X1 U6956 ( .A1(n6136), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n6126)
         );
  OAI22_X1 U6957 ( .A1(n6178), .A2(n6138), .B1(n6137), .B2(n6436), .ZN(n6124)
         );
  AOI21_X1 U6958 ( .B1(n6181), .B2(n6140), .A(n6124), .ZN(n6125) );
  OAI211_X1 U6959 ( .C1(n6143), .C2(n6179), .A(n6126), .B(n6125), .ZN(U3134)
         );
  NAND2_X1 U6960 ( .A1(n6144), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n6129) );
  OAI22_X1 U6961 ( .A1(n6172), .A2(n6146), .B1(n6145), .B2(n6429), .ZN(n6127)
         );
  AOI21_X1 U6962 ( .B1(n6175), .B2(n6148), .A(n6127), .ZN(n6128) );
  OAI211_X1 U6963 ( .C1(n6151), .C2(n6173), .A(n6129), .B(n6128), .ZN(U3053)
         );
  NAND2_X1 U6964 ( .A1(n6144), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n6132) );
  OAI22_X1 U6965 ( .A1(n6168), .A2(n6146), .B1(n6145), .B2(n6394), .ZN(n6130)
         );
  AOI21_X1 U6966 ( .B1(n6188), .B2(n6148), .A(n6130), .ZN(n6131) );
  OAI211_X1 U6967 ( .C1(n6151), .C2(n6185), .A(n6132), .B(n6131), .ZN(U3057)
         );
  NAND2_X1 U6968 ( .A1(n6144), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n6135) );
  OAI22_X1 U6969 ( .A1(n6178), .A2(n6146), .B1(n6145), .B2(n6436), .ZN(n6133)
         );
  AOI21_X1 U6970 ( .B1(n6181), .B2(n6148), .A(n6133), .ZN(n6134) );
  OAI211_X1 U6971 ( .C1(n6151), .C2(n6179), .A(n6135), .B(n6134), .ZN(U3054)
         );
  NAND2_X1 U6972 ( .A1(n6136), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n6142)
         );
  OAI22_X1 U6973 ( .A1(n6192), .A2(n6138), .B1(n6137), .B2(n6447), .ZN(n6139)
         );
  AOI21_X1 U6974 ( .B1(n6196), .B2(n6140), .A(n6139), .ZN(n6141) );
  OAI211_X1 U6975 ( .C1(n6143), .C2(n6193), .A(n6142), .B(n6141), .ZN(U3132)
         );
  NAND2_X1 U6976 ( .A1(n6144), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n6150) );
  OAI22_X1 U6977 ( .A1(n6192), .A2(n6146), .B1(n6145), .B2(n6447), .ZN(n6147)
         );
  AOI21_X1 U6978 ( .B1(n6196), .B2(n6148), .A(n6147), .ZN(n6149) );
  OAI211_X1 U6979 ( .C1(n6151), .C2(n6193), .A(n6150), .B(n6149), .ZN(U3052)
         );
  OAI22_X1 U6980 ( .A1(n6442), .A2(n6179), .B1(n6178), .B2(n6161), .ZN(n6152)
         );
  AOI21_X1 U6981 ( .B1(n6181), .B2(n6163), .A(n6152), .ZN(n6154) );
  NAND2_X1 U6982 ( .A1(n6164), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n6153)
         );
  OAI211_X1 U6983 ( .C1(n6167), .C2(n6436), .A(n6154), .B(n6153), .ZN(U3110)
         );
  OAI22_X1 U6984 ( .A1(n6442), .A2(n6173), .B1(n6172), .B2(n6161), .ZN(n6155)
         );
  AOI21_X1 U6985 ( .B1(n6175), .B2(n6163), .A(n6155), .ZN(n6157) );
  NAND2_X1 U6986 ( .A1(n6164), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n6156)
         );
  OAI211_X1 U6987 ( .C1(n6167), .C2(n6429), .A(n6157), .B(n6156), .ZN(U3109)
         );
  OAI22_X1 U6988 ( .A1(n6442), .A2(n6193), .B1(n6192), .B2(n6161), .ZN(n6158)
         );
  AOI21_X1 U6989 ( .B1(n6196), .B2(n6163), .A(n6158), .ZN(n6160) );
  NAND2_X1 U6990 ( .A1(n6164), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n6159)
         );
  OAI211_X1 U6991 ( .C1(n6167), .C2(n6447), .A(n6160), .B(n6159), .ZN(U3108)
         );
  OAI22_X1 U6992 ( .A1(n6442), .A2(n6185), .B1(n6168), .B2(n6161), .ZN(n6162)
         );
  AOI21_X1 U6993 ( .B1(n6188), .B2(n6163), .A(n6162), .ZN(n6166) );
  NAND2_X1 U6994 ( .A1(n6164), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n6165)
         );
  OAI211_X1 U6995 ( .C1(n6167), .C2(n6394), .A(n6166), .B(n6165), .ZN(U3113)
         );
  OAI22_X1 U6996 ( .A1(n6363), .A2(n6185), .B1(n6168), .B2(n6191), .ZN(n6169)
         );
  AOI21_X1 U6997 ( .B1(n6188), .B2(n6195), .A(n6169), .ZN(n6171) );
  NAND2_X1 U6998 ( .A1(n6197), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n6170) );
  OAI211_X1 U6999 ( .C1(n6200), .C2(n6394), .A(n6171), .B(n6170), .ZN(U3049)
         );
  OAI22_X1 U7000 ( .A1(n6363), .A2(n6173), .B1(n6172), .B2(n6191), .ZN(n6174)
         );
  AOI21_X1 U7001 ( .B1(n6175), .B2(n6195), .A(n6174), .ZN(n6177) );
  NAND2_X1 U7002 ( .A1(n6197), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n6176) );
  OAI211_X1 U7003 ( .C1(n6200), .C2(n6429), .A(n6177), .B(n6176), .ZN(U3045)
         );
  OAI22_X1 U7004 ( .A1(n6363), .A2(n6179), .B1(n6178), .B2(n6191), .ZN(n6180)
         );
  AOI21_X1 U7005 ( .B1(n6181), .B2(n6195), .A(n6180), .ZN(n6183) );
  NAND2_X1 U7006 ( .A1(n6197), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n6182) );
  OAI211_X1 U7007 ( .C1(n6200), .C2(n6436), .A(n6183), .B(n6182), .ZN(U3046)
         );
  INV_X1 U7008 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n6190) );
  AOI22_X1 U7009 ( .A1(n6210), .A2(n6334), .B1(n6388), .B2(n6209), .ZN(n6184)
         );
  OAI21_X1 U7010 ( .B1(n6186), .B2(n6185), .A(n6184), .ZN(n6187) );
  AOI21_X1 U7011 ( .B1(n6188), .B2(n6365), .A(n6187), .ZN(n6189) );
  OAI21_X1 U7012 ( .B1(n6217), .B2(n6190), .A(n6189), .ZN(U3033) );
  OAI22_X1 U7013 ( .A1(n6363), .A2(n6193), .B1(n6192), .B2(n6191), .ZN(n6194)
         );
  AOI21_X1 U7014 ( .B1(n6196), .B2(n6195), .A(n6194), .ZN(n6199) );
  NAND2_X1 U7015 ( .A1(n6197), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n6198) );
  OAI211_X1 U7016 ( .C1(n6200), .C2(n6447), .A(n6199), .B(n6198), .ZN(U3044)
         );
  INV_X1 U7017 ( .A(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n6204) );
  AOI22_X1 U7018 ( .A1(n6210), .A2(n6349), .B1(n6423), .B2(n6209), .ZN(n6201)
         );
  OAI21_X1 U7019 ( .B1(n6425), .B2(n6212), .A(n6201), .ZN(n6202) );
  AOI21_X1 U7020 ( .B1(n6427), .B2(n6214), .A(n6202), .ZN(n6203) );
  OAI21_X1 U7021 ( .B1(n6217), .B2(n6204), .A(n6203), .ZN(U3029) );
  INV_X1 U7022 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n6208) );
  AOI22_X1 U7023 ( .A1(n6210), .A2(n6339), .B1(n6430), .B2(n6209), .ZN(n6205)
         );
  OAI21_X1 U7024 ( .B1(n6432), .B2(n6212), .A(n6205), .ZN(n6206) );
  AOI21_X1 U7025 ( .B1(n6434), .B2(n6214), .A(n6206), .ZN(n6207) );
  OAI21_X1 U7026 ( .B1(n6217), .B2(n6208), .A(n6207), .ZN(U3030) );
  INV_X1 U7027 ( .A(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n6216) );
  AOI22_X1 U7028 ( .A1(n6210), .A2(n6324), .B1(n6439), .B2(n6209), .ZN(n6211)
         );
  OAI21_X1 U7029 ( .B1(n6441), .B2(n6212), .A(n6211), .ZN(n6213) );
  AOI21_X1 U7030 ( .B1(n6445), .B2(n6214), .A(n6213), .ZN(n6215) );
  OAI21_X1 U7031 ( .B1(n6217), .B2(n6216), .A(n6215), .ZN(U3028) );
  XNOR2_X1 U7032 ( .A(n3646), .B(STATEBS16_REG_SCAN_IN), .ZN(n6219) );
  XNOR2_X1 U7033 ( .A(n6220), .B(n6221), .ZN(n6251) );
  INV_X1 U7034 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6222) );
  AOI21_X1 U7035 ( .B1(n6222), .B2(n5149), .A(n6273), .ZN(n6223) );
  NAND2_X1 U7036 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6473) );
  AOI22_X1 U7037 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n6271), .B1(n6223), 
        .B2(n6473), .ZN(n6227) );
  INV_X1 U7038 ( .A(n6224), .ZN(n7600) );
  INV_X1 U7039 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6225) );
  NOR2_X1 U7040 ( .A1(n7524), .A2(n6225), .ZN(n6246) );
  AOI21_X1 U7041 ( .B1(n7600), .B2(n7545), .A(n6246), .ZN(n6226) );
  OAI211_X1 U7042 ( .C1(n6251), .C2(n7506), .A(n6227), .B(n6226), .ZN(U3010)
         );
  INV_X1 U7043 ( .A(n6228), .ZN(n6229) );
  OAI21_X1 U7044 ( .B1(n6005), .B2(n6230), .A(n6228), .ZN(n7614) );
  OR2_X1 U7045 ( .A1(n6007), .A2(n6232), .ZN(n6233) );
  NAND2_X1 U7046 ( .A1(n6265), .A2(n6233), .ZN(n7610) );
  OAI22_X1 U7047 ( .A1(n7610), .A2(n6917), .B1(n7611), .B2(n7369), .ZN(n6234)
         );
  INV_X1 U7048 ( .A(n6234), .ZN(n6235) );
  OAI21_X1 U7049 ( .B1(n7614), .B2(n6919), .A(n6235), .ZN(U2850) );
  INV_X1 U7050 ( .A(EAX_REG_18__SCAN_IN), .ZN(n6237) );
  AOI22_X1 U7051 ( .A1(n7284), .A2(UWORD_REG_2__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n6236) );
  OAI21_X1 U7052 ( .B1(n6237), .B2(n6244), .A(n6236), .ZN(U2905) );
  INV_X1 U7053 ( .A(EAX_REG_19__SCAN_IN), .ZN(n6239) );
  AOI22_X1 U7054 ( .A1(n7284), .A2(UWORD_REG_3__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n6238) );
  OAI21_X1 U7055 ( .B1(n6239), .B2(n6244), .A(n6238), .ZN(U2904) );
  INV_X1 U7056 ( .A(EAX_REG_16__SCAN_IN), .ZN(n6241) );
  AOI22_X1 U7057 ( .A1(n7284), .A2(UWORD_REG_0__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n6240) );
  OAI21_X1 U7058 ( .B1(n6241), .B2(n6244), .A(n6240), .ZN(U2907) );
  AOI22_X1 U7059 ( .A1(n7284), .A2(UWORD_REG_1__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n6242) );
  OAI21_X1 U7060 ( .B1(n4495), .B2(n6244), .A(n6242), .ZN(U2906) );
  INV_X1 U7061 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6245) );
  AOI22_X1 U7062 ( .A1(n7284), .A2(UWORD_REG_14__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n6243) );
  OAI21_X1 U7063 ( .B1(n6245), .B2(n6244), .A(n6243), .ZN(U2893) );
  AOI21_X1 U7064 ( .B1(n7415), .B2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6246), 
        .ZN(n6248) );
  OR2_X1 U7065 ( .A1(n7425), .A2(n7604), .ZN(n6247) );
  OAI211_X1 U7066 ( .C1(n7605), .C2(n7052), .A(n6248), .B(n6247), .ZN(n6249)
         );
  INV_X1 U7067 ( .A(n6249), .ZN(n6250) );
  OAI21_X1 U7068 ( .B1(n6251), .B2(n7701), .A(n6250), .ZN(U2978) );
  INV_X1 U7069 ( .A(EAX_REG_9__SCAN_IN), .ZN(n7274) );
  OAI222_X1 U7070 ( .A1(n7614), .A2(n7751), .B1(n6953), .B2(n6252), .C1(n6952), 
        .C2(n7274), .ZN(U2882) );
  INV_X1 U7071 ( .A(n6253), .ZN(n6254) );
  NOR3_X1 U7072 ( .A1(n7251), .A2(n7221), .A3(n6254), .ZN(n6258) );
  NOR2_X1 U7073 ( .A1(n6256), .A2(n6255), .ZN(n6257) );
  AOI211_X1 U7074 ( .C1(n7251), .C2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n6258), .B(n6257), .ZN(n6259) );
  OAI21_X1 U7075 ( .B1(n6648), .B2(n6260), .A(n6259), .ZN(U3465) );
  NOR2_X1 U7076 ( .A1(n6229), .A2(n6262), .ZN(n6263) );
  OR2_X1 U7077 ( .A1(n6261), .A2(n6263), .ZN(n7625) );
  AOI21_X1 U7078 ( .B1(n6266), .B2(n6265), .A(n3682), .ZN(n7621) );
  AOI22_X1 U7079 ( .A1(n7621), .A2(n6914), .B1(EBX_REG_10__SCAN_IN), .B2(n6913), .ZN(n6267) );
  OAI21_X1 U7080 ( .B1(n7625), .B2(n6919), .A(n6267), .ZN(U2849) );
  XNOR2_X1 U7081 ( .A(n6268), .B(n6269), .ZN(n6461) );
  INV_X1 U7082 ( .A(n6270), .ZN(n6272) );
  OAI22_X1 U7083 ( .A1(n7508), .A2(n6272), .B1(n6271), .B2(n6473), .ZN(n7488)
         );
  INV_X1 U7084 ( .A(n7488), .ZN(n6276) );
  OR2_X1 U7085 ( .A1(n7524), .A2(n7619), .ZN(n6456) );
  NOR2_X1 U7086 ( .A1(n6473), .A2(n6273), .ZN(n7483) );
  NAND2_X1 U7087 ( .A1(n7482), .A2(n7483), .ZN(n6274) );
  OAI211_X1 U7088 ( .C1(n7610), .C2(n7555), .A(n6456), .B(n6274), .ZN(n6275)
         );
  AOI21_X1 U7089 ( .B1(n6276), .B2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n6275), 
        .ZN(n6277) );
  OAI21_X1 U7090 ( .B1(n6461), .B2(n7506), .A(n6277), .ZN(U3009) );
  INV_X1 U7091 ( .A(EAX_REG_10__SCAN_IN), .ZN(n7276) );
  OAI222_X1 U7092 ( .A1(n7625), .A2(n7751), .B1(n6278), .B2(n6953), .C1(n6952), 
        .C2(n7276), .ZN(U2881) );
  NOR2_X1 U7093 ( .A1(n6281), .A2(n3946), .ZN(n6279) );
  OR3_X1 U7094 ( .A1(n6281), .A2(n3956), .A3(n6280), .ZN(n6307) );
  OAI22_X1 U7095 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6808), .B1(n6307), .B2(n5438), .ZN(n6287) );
  AOI22_X1 U7096 ( .A1(n7688), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6843), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n6284) );
  INV_X1 U7097 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6282) );
  NAND2_X1 U7098 ( .A1(n7682), .A2(n6282), .ZN(n6283) );
  OAI211_X1 U7099 ( .C1(n6285), .C2(n7686), .A(n6284), .B(n6283), .ZN(n6286)
         );
  AOI211_X1 U7100 ( .C1(n7666), .C2(n5352), .A(n6287), .B(n6286), .ZN(n6288)
         );
  OAI21_X1 U7101 ( .B1(n7370), .B2(n6879), .A(n6288), .ZN(U2826) );
  OAI21_X1 U7102 ( .B1(n6261), .B2(n6291), .A(n6290), .ZN(n6369) );
  INV_X1 U7103 ( .A(EAX_REG_11__SCAN_IN), .ZN(n7278) );
  OAI222_X1 U7104 ( .A1(n6369), .A2(n7751), .B1(n6953), .B2(n6292), .C1(n6952), 
        .C2(n7278), .ZN(U2880) );
  INV_X1 U7105 ( .A(n6293), .ZN(n7386) );
  NOR2_X1 U7106 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6294), .ZN(n6295) );
  AOI22_X1 U7107 ( .A1(n7687), .A2(EBX_REG_4__SCAN_IN), .B1(n6876), .B2(n6295), 
        .ZN(n6301) );
  NAND2_X1 U7108 ( .A1(n7666), .A2(n7450), .ZN(n6300) );
  INV_X1 U7109 ( .A(n7389), .ZN(n6296) );
  AOI21_X1 U7110 ( .B1(n7682), .B2(n6296), .A(n7677), .ZN(n6299) );
  INV_X1 U7111 ( .A(n6307), .ZN(n6874) );
  NAND2_X1 U7112 ( .A1(n6297), .A2(n6874), .ZN(n6298) );
  NAND4_X1 U7113 ( .A1(n6301), .A2(n6300), .A3(n6299), .A4(n6298), .ZN(n6304)
         );
  INV_X1 U7114 ( .A(REIP_REG_3__SCAN_IN), .ZN(n7290) );
  NAND3_X1 U7115 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .A3(
        n6871), .ZN(n6864) );
  OAI21_X1 U7116 ( .B1(n7290), .B2(n6864), .A(n7598), .ZN(n6863) );
  OAI22_X1 U7117 ( .A1(n6302), .A2(n7633), .B1(n7292), .B2(n6863), .ZN(n6303)
         );
  AOI211_X1 U7118 ( .C1(n7386), .C2(n7569), .A(n6304), .B(n6303), .ZN(n6305)
         );
  INV_X1 U7119 ( .A(n6305), .ZN(U2823) );
  OAI21_X1 U7120 ( .B1(n7682), .B2(n7688), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n6306) );
  OAI21_X1 U7121 ( .B1(n6307), .B2(n6648), .A(n6306), .ZN(n6310) );
  INV_X1 U7122 ( .A(n7598), .ZN(n6844) );
  INV_X1 U7123 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6308) );
  OAI22_X1 U7124 ( .A1(n6844), .A2(n6308), .B1(n7693), .B2(n7554), .ZN(n6309)
         );
  AOI211_X1 U7125 ( .C1(n7687), .C2(EBX_REG_0__SCAN_IN), .A(n6310), .B(n6309), 
        .ZN(n6311) );
  OAI21_X1 U7126 ( .B1(n6879), .B2(n6312), .A(n6311), .ZN(U2827) );
  OAI21_X1 U7127 ( .B1(n6365), .B2(n6314), .A(n6313), .ZN(n6315) );
  OAI21_X1 U7128 ( .B1(n3645), .B2(n6377), .A(n6315), .ZN(n6317) );
  NOR2_X1 U7129 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6316), .ZN(n6361)
         );
  AOI21_X1 U7130 ( .B1(n6317), .B2(n7724), .A(n6361), .ZN(n6320) );
  INV_X1 U7131 ( .A(n6318), .ZN(n6319) );
  NOR3_X2 U7132 ( .A1(n6320), .A2(n6384), .A3(n6319), .ZN(n6368) );
  INV_X1 U7133 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n6328) );
  OAI22_X1 U7134 ( .A1(n6323), .A2(n6377), .B1(n6322), .B2(n6321), .ZN(n6359)
         );
  AOI22_X1 U7135 ( .A1(n6439), .A2(n6361), .B1(n6324), .B2(n6359), .ZN(n6325)
         );
  OAI21_X1 U7136 ( .B1(n6441), .B2(n6363), .A(n6325), .ZN(n6326) );
  AOI21_X1 U7137 ( .B1(n6365), .B2(n6445), .A(n6326), .ZN(n6327) );
  OAI21_X1 U7138 ( .B1(n6368), .B2(n6328), .A(n6327), .ZN(U3036) );
  INV_X1 U7139 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n6333) );
  AOI22_X1 U7140 ( .A1(n6402), .A2(n6361), .B1(n6329), .B2(n6359), .ZN(n6330)
         );
  OAI21_X1 U7141 ( .B1(n6363), .B2(n6404), .A(n6330), .ZN(n6331) );
  AOI21_X1 U7142 ( .B1(n6406), .B2(n6365), .A(n6331), .ZN(n6332) );
  OAI21_X1 U7143 ( .B1(n6368), .B2(n6333), .A(n6332), .ZN(U3042) );
  INV_X1 U7144 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n6338) );
  AOI22_X1 U7145 ( .A1(n7767), .A2(n6361), .B1(n6334), .B2(n6359), .ZN(n6335)
         );
  OAI21_X1 U7146 ( .B1(n6363), .B2(n6390), .A(n6335), .ZN(n6336) );
  AOI21_X1 U7147 ( .B1(n6392), .B2(n6365), .A(n6336), .ZN(n6337) );
  OAI21_X1 U7148 ( .B1(n6368), .B2(n6338), .A(n6337), .ZN(U3041) );
  INV_X1 U7149 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n6343) );
  AOI22_X1 U7150 ( .A1(n6430), .A2(n6361), .B1(n6339), .B2(n6359), .ZN(n6340)
         );
  OAI21_X1 U7151 ( .B1(n6363), .B2(n6432), .A(n6340), .ZN(n6341) );
  AOI21_X1 U7152 ( .B1(n6434), .B2(n6365), .A(n6341), .ZN(n6342) );
  OAI21_X1 U7153 ( .B1(n6368), .B2(n6343), .A(n6342), .ZN(U3038) );
  INV_X1 U7154 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n6348) );
  AOI22_X1 U7155 ( .A1(n6409), .A2(n6361), .B1(n6344), .B2(n6359), .ZN(n6345)
         );
  OAI21_X1 U7156 ( .B1(n6363), .B2(n6411), .A(n6345), .ZN(n6346) );
  AOI21_X1 U7157 ( .B1(n6413), .B2(n6365), .A(n6346), .ZN(n6347) );
  OAI21_X1 U7158 ( .B1(n6368), .B2(n6348), .A(n6347), .ZN(U3040) );
  INV_X1 U7159 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n6353) );
  AOI22_X1 U7160 ( .A1(n3678), .A2(n6361), .B1(n6349), .B2(n6359), .ZN(n6350)
         );
  OAI21_X1 U7161 ( .B1(n6363), .B2(n6425), .A(n6350), .ZN(n6351) );
  AOI21_X1 U7162 ( .B1(n6427), .B2(n6365), .A(n6351), .ZN(n6352) );
  OAI21_X1 U7163 ( .B1(n6368), .B2(n6353), .A(n6352), .ZN(U3037) );
  INV_X1 U7164 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n6358) );
  AOI22_X1 U7165 ( .A1(n6416), .A2(n6361), .B1(n6354), .B2(n6359), .ZN(n6355)
         );
  OAI21_X1 U7166 ( .B1(n6363), .B2(n6418), .A(n6355), .ZN(n6356) );
  AOI21_X1 U7167 ( .B1(n6420), .B2(n6365), .A(n6356), .ZN(n6357) );
  OAI21_X1 U7168 ( .B1(n6368), .B2(n6358), .A(n6357), .ZN(U3039) );
  INV_X1 U7169 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n6367) );
  AOI22_X1 U7170 ( .A1(n6395), .A2(n6361), .B1(n6360), .B2(n6359), .ZN(n6362)
         );
  OAI21_X1 U7171 ( .B1(n6363), .B2(n6397), .A(n6362), .ZN(n6364) );
  AOI21_X1 U7172 ( .B1(n6399), .B2(n6365), .A(n6364), .ZN(n6366) );
  OAI21_X1 U7173 ( .B1(n6368), .B2(n6367), .A(n6366), .ZN(U3043) );
  INV_X1 U7174 ( .A(n6369), .ZN(n7639) );
  NAND2_X1 U7175 ( .A1(n6264), .A2(n6370), .ZN(n6371) );
  NAND2_X1 U7176 ( .A1(n6451), .A2(n6371), .ZN(n7634) );
  OAI22_X1 U7177 ( .A1(n7634), .A2(n6917), .B1(n7635), .B2(n7369), .ZN(n6372)
         );
  AOI21_X1 U7178 ( .B1(n7639), .B2(n7366), .A(n6372), .ZN(n6373) );
  INV_X1 U7179 ( .A(n6373), .ZN(U2848) );
  AOI21_X1 U7180 ( .B1(n6376), .B2(STATEBS16_REG_SCAN_IN), .A(n6375), .ZN(
        n6386) );
  NOR2_X1 U7181 ( .A1(n6378), .A2(n6377), .ZN(n6382) );
  NOR2_X1 U7182 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6381), .ZN(n6438)
         );
  INV_X1 U7183 ( .A(n6382), .ZN(n6385) );
  AOI211_X1 U7184 ( .C1(n6386), .C2(n6385), .A(n6384), .B(n6383), .ZN(n6387)
         );
  OAI21_X1 U7185 ( .B1(n6438), .B2(n7724), .A(n6387), .ZN(n6437) );
  AOI22_X1 U7186 ( .A1(n7767), .A2(n6438), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n6437), .ZN(n6389) );
  OAI21_X1 U7187 ( .B1(n6442), .B2(n6390), .A(n6389), .ZN(n6391) );
  AOI21_X1 U7188 ( .B1(n3621), .B2(n6392), .A(n6391), .ZN(n6393) );
  OAI21_X1 U7189 ( .B1(n6448), .B2(n6394), .A(n6393), .ZN(U3105) );
  AOI22_X1 U7190 ( .A1(n6395), .A2(n6438), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n6437), .ZN(n6396) );
  OAI21_X1 U7191 ( .B1(n6442), .B2(n6397), .A(n6396), .ZN(n6398) );
  AOI21_X1 U7192 ( .B1(n3621), .B2(n6399), .A(n6398), .ZN(n6400) );
  OAI21_X1 U7193 ( .B1(n6448), .B2(n6401), .A(n6400), .ZN(U3107) );
  AOI22_X1 U7194 ( .A1(n6402), .A2(n6438), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n6437), .ZN(n6403) );
  OAI21_X1 U7195 ( .B1(n6442), .B2(n6404), .A(n6403), .ZN(n6405) );
  AOI21_X1 U7196 ( .B1(n3621), .B2(n6406), .A(n6405), .ZN(n6407) );
  OAI21_X1 U7197 ( .B1(n6448), .B2(n6408), .A(n6407), .ZN(U3106) );
  AOI22_X1 U7198 ( .A1(n6409), .A2(n6438), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n6437), .ZN(n6410) );
  OAI21_X1 U7199 ( .B1(n6442), .B2(n6411), .A(n6410), .ZN(n6412) );
  AOI21_X1 U7200 ( .B1(n3621), .B2(n6413), .A(n6412), .ZN(n6414) );
  OAI21_X1 U7201 ( .B1(n6448), .B2(n6415), .A(n6414), .ZN(U3104) );
  AOI22_X1 U7202 ( .A1(n6416), .A2(n6438), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n6437), .ZN(n6417) );
  OAI21_X1 U7203 ( .B1(n6442), .B2(n6418), .A(n6417), .ZN(n6419) );
  AOI21_X1 U7204 ( .B1(n3621), .B2(n6420), .A(n6419), .ZN(n6421) );
  OAI21_X1 U7205 ( .B1(n6448), .B2(n6422), .A(n6421), .ZN(U3103) );
  AOI22_X1 U7206 ( .A1(n3678), .A2(n6438), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n6437), .ZN(n6424) );
  OAI21_X1 U7207 ( .B1(n6425), .B2(n6442), .A(n6424), .ZN(n6426) );
  AOI21_X1 U7208 ( .B1(n3621), .B2(n6427), .A(n6426), .ZN(n6428) );
  OAI21_X1 U7209 ( .B1(n6448), .B2(n6429), .A(n6428), .ZN(U3101) );
  AOI22_X1 U7210 ( .A1(n6430), .A2(n6438), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n6437), .ZN(n6431) );
  OAI21_X1 U7211 ( .B1(n6442), .B2(n6432), .A(n6431), .ZN(n6433) );
  AOI21_X1 U7212 ( .B1(n3621), .B2(n6434), .A(n6433), .ZN(n6435) );
  OAI21_X1 U7213 ( .B1(n6448), .B2(n6436), .A(n6435), .ZN(U3102) );
  AOI22_X1 U7214 ( .A1(n6439), .A2(n6438), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n6437), .ZN(n6440) );
  OAI21_X1 U7215 ( .B1(n6442), .B2(n6441), .A(n6440), .ZN(n6443) );
  AOI21_X1 U7216 ( .B1(n6445), .B2(n3621), .A(n6443), .ZN(n6446) );
  OAI21_X1 U7217 ( .B1(n6448), .B2(n6447), .A(n6446), .ZN(U3100) );
  XNOR2_X1 U7218 ( .A(n6290), .B(n6449), .ZN(n6855) );
  AND2_X1 U7219 ( .A1(n6451), .A2(n6450), .ZN(n6452) );
  OR2_X1 U7220 ( .A1(n6452), .A2(n6483), .ZN(n7493) );
  OAI22_X1 U7221 ( .A1(n7493), .A2(n6917), .B1(n6453), .B2(n7369), .ZN(n6454)
         );
  INV_X1 U7222 ( .A(n6454), .ZN(n6455) );
  OAI21_X1 U7223 ( .B1(n6855), .B2(n6919), .A(n6455), .ZN(U2847) );
  INV_X1 U7224 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6457) );
  OAI21_X1 U7225 ( .B1(n7405), .B2(n6457), .A(n6456), .ZN(n6459) );
  NOR2_X1 U7226 ( .A1(n7614), .A2(n7052), .ZN(n6458) );
  AOI211_X1 U7227 ( .C1(n7409), .C2(n7616), .A(n6459), .B(n6458), .ZN(n6460)
         );
  OAI21_X1 U7228 ( .B1(n6461), .B2(n7701), .A(n6460), .ZN(U2977) );
  NAND2_X1 U7229 ( .A1(n6502), .A2(n6463), .ZN(n6464) );
  XNOR2_X1 U7230 ( .A(n6462), .B(n6464), .ZN(n7485) );
  NAND2_X1 U7231 ( .A1(n7485), .A2(n7422), .ZN(n6467) );
  NOR2_X1 U7232 ( .A1(n7524), .A2(n7631), .ZN(n7480) );
  NOR2_X1 U7233 ( .A1(n7425), .A2(n7624), .ZN(n6465) );
  AOI211_X1 U7234 ( .C1(n7415), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n7480), 
        .B(n6465), .ZN(n6466) );
  OAI211_X1 U7235 ( .C1(n7052), .C2(n7625), .A(n6467), .B(n6466), .ZN(U2976)
         );
  OAI222_X1 U7236 ( .A1(n7751), .A2(n6855), .B1(n6952), .B2(n4396), .C1(n6468), 
        .C2(n6953), .ZN(U2879) );
  XNOR2_X1 U7237 ( .A(n6469), .B(n6470), .ZN(n7412) );
  INV_X1 U7238 ( .A(n7412), .ZN(n6490) );
  NAND2_X1 U7239 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6479) );
  NOR2_X1 U7240 ( .A1(n5168), .A2(n6479), .ZN(n6541) );
  INV_X1 U7241 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n7489) );
  NOR2_X1 U7242 ( .A1(n7489), .A2(n7482), .ZN(n7481) );
  OAI21_X1 U7243 ( .B1(n6580), .B2(n7481), .A(n7488), .ZN(n7507) );
  AOI21_X1 U7244 ( .B1(n6471), .B2(n6479), .A(n7507), .ZN(n6480) );
  INV_X1 U7245 ( .A(n7481), .ZN(n6472) );
  NOR2_X1 U7246 ( .A1(n6473), .A2(n6472), .ZN(n6477) );
  NAND2_X1 U7247 ( .A1(n6477), .A2(n6474), .ZN(n6542) );
  NOR3_X1 U7248 ( .A1(n6475), .A2(n6542), .A3(n7562), .ZN(n6476) );
  NOR2_X1 U7249 ( .A1(n6476), .A2(n6550), .ZN(n7490) );
  NAND2_X1 U7250 ( .A1(n6478), .A2(n6477), .ZN(n6546) );
  NOR2_X1 U7251 ( .A1(n7490), .A2(n6546), .ZN(n6521) );
  NOR2_X1 U7252 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6479), .ZN(n6485)
         );
  NAND2_X1 U7253 ( .A1(n6521), .A2(n6485), .ZN(n6481) );
  OAI211_X1 U7254 ( .C1(n6541), .C2(n7561), .A(n6480), .B(n6481), .ZN(n6525)
         );
  NAND2_X1 U7255 ( .A1(n5168), .A2(n6481), .ZN(n6488) );
  OR2_X1 U7256 ( .A1(n6483), .A2(n6482), .ZN(n6484) );
  NAND2_X1 U7257 ( .A1(n6516), .A2(n6484), .ZN(n7647) );
  NOR2_X1 U7258 ( .A1(n7561), .A2(n6542), .ZN(n7492) );
  AOI22_X1 U7259 ( .A1(n7544), .A2(REIP_REG_13__SCAN_IN), .B1(n6485), .B2(
        n7492), .ZN(n6486) );
  OAI21_X1 U7260 ( .B1(n7647), .B2(n7555), .A(n6486), .ZN(n6487) );
  AOI21_X1 U7261 ( .B1(n6525), .B2(n6488), .A(n6487), .ZN(n6489) );
  OAI21_X1 U7262 ( .B1(n6490), .B2(n7506), .A(n6489), .ZN(U3005) );
  INV_X1 U7263 ( .A(n6491), .ZN(n6494) );
  INV_X1 U7264 ( .A(n6492), .ZN(n6493) );
  NAND2_X1 U7265 ( .A1(n6494), .A2(n6493), .ZN(n6496) );
  AND2_X1 U7266 ( .A1(n6496), .A2(n6495), .ZN(n7656) );
  OAI22_X1 U7267 ( .A1(n7647), .A2(n6917), .B1(n7650), .B2(n7369), .ZN(n6497)
         );
  AOI21_X1 U7268 ( .B1(n7656), .B2(n7366), .A(n6497), .ZN(n6498) );
  INV_X1 U7269 ( .A(n6498), .ZN(U2846) );
  INV_X1 U7270 ( .A(n7656), .ZN(n6500) );
  INV_X1 U7271 ( .A(DATAI_13_), .ZN(n6499) );
  INV_X1 U7272 ( .A(EAX_REG_13__SCAN_IN), .ZN(n7281) );
  OAI222_X1 U7273 ( .A1(n6500), .A2(n7751), .B1(n6499), .B2(n6953), .C1(n6952), 
        .C2(n7281), .ZN(U2878) );
  NAND2_X1 U7274 ( .A1(n6501), .A2(n6502), .ZN(n7408) );
  INV_X1 U7275 ( .A(n6505), .ZN(n6504) );
  NOR2_X1 U7276 ( .A1(n6504), .A2(n6503), .ZN(n7407) );
  NAND2_X1 U7277 ( .A1(n7408), .A2(n7407), .ZN(n7406) );
  NAND2_X1 U7278 ( .A1(n7406), .A2(n6505), .ZN(n6508) );
  XNOR2_X1 U7279 ( .A(n4252), .B(n6506), .ZN(n6507) );
  XNOR2_X1 U7280 ( .A(n6508), .B(n6507), .ZN(n7497) );
  NAND2_X1 U7281 ( .A1(n7497), .A2(n7422), .ZN(n6512) );
  INV_X1 U7282 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6509) );
  NOR2_X1 U7283 ( .A1(n7524), .A2(n6509), .ZN(n7494) );
  NOR2_X1 U7284 ( .A1(n7405), .A2(n6848), .ZN(n6510) );
  AOI211_X1 U7285 ( .C1(n7409), .C2(n6850), .A(n7494), .B(n6510), .ZN(n6511)
         );
  OAI211_X1 U7286 ( .C1(n6855), .C2(n7052), .A(n6512), .B(n6511), .ZN(U2974)
         );
  XNOR2_X1 U7287 ( .A(n4252), .B(n6514), .ZN(n6515) );
  XNOR2_X1 U7288 ( .A(n6513), .B(n6515), .ZN(n7058) );
  INV_X1 U7289 ( .A(n6516), .ZN(n6520) );
  INV_X1 U7290 ( .A(n6517), .ZN(n6519) );
  INV_X1 U7291 ( .A(n6518), .ZN(n6827) );
  OAI21_X1 U7292 ( .B1(n6520), .B2(n6519), .A(n6827), .ZN(n6916) );
  NOR2_X1 U7293 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n7542), .ZN(n6522)
         );
  NAND2_X1 U7294 ( .A1(n6522), .A2(n6541), .ZN(n6523) );
  NAND2_X1 U7295 ( .A1(n7544), .A2(REIP_REG_14__SCAN_IN), .ZN(n7050) );
  OAI211_X1 U7296 ( .C1(n7555), .C2(n6916), .A(n6523), .B(n7050), .ZN(n6524)
         );
  AOI21_X1 U7297 ( .B1(n6525), .B2(INSTADDRPOINTER_REG_14__SCAN_IN), .A(n6524), 
        .ZN(n6526) );
  OAI21_X1 U7298 ( .B1(n7058), .B2(n7506), .A(n6526), .ZN(U3004) );
  INV_X1 U7299 ( .A(n7019), .ZN(n6528) );
  INV_X1 U7300 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n7160) );
  XNOR2_X1 U7301 ( .A(n4252), .B(n7160), .ZN(n7018) );
  INV_X1 U7302 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6529) );
  NAND2_X1 U7303 ( .A1(n3625), .A2(n3743), .ZN(n6533) );
  INV_X1 U7304 ( .A(n7119), .ZN(n7152) );
  NAND2_X1 U7305 ( .A1(n4252), .A2(n7152), .ZN(n6530) );
  NAND2_X1 U7306 ( .A1(n6533), .A2(n6530), .ZN(n7000) );
  INV_X1 U7307 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n7135) );
  XNOR2_X1 U7308 ( .A(n4252), .B(n7135), .ZN(n6999) );
  AOI21_X1 U7309 ( .B1(n3631), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n6998), 
        .ZN(n6992) );
  NOR2_X1 U7310 ( .A1(n7110), .A2(n6531), .ZN(n6532) );
  NAND2_X1 U7311 ( .A1(n4252), .A2(n6532), .ZN(n6537) );
  INV_X1 U7312 ( .A(n6533), .ZN(n6534) );
  NAND2_X1 U7313 ( .A1(n6534), .A2(n7122), .ZN(n6982) );
  NOR2_X1 U7314 ( .A1(n6982), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6535)
         );
  XNOR2_X1 U7315 ( .A(n6538), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6569)
         );
  AND2_X1 U7316 ( .A1(n6758), .A2(n6539), .ZN(n6540) );
  NOR2_X1 U7317 ( .A1(n6735), .A2(n6540), .ZN(n6888) );
  NOR2_X1 U7318 ( .A1(n7524), .A2(n7323), .ZN(n6565) );
  NOR2_X1 U7319 ( .A1(n7516), .A2(n7514), .ZN(n7148) );
  INV_X1 U7320 ( .A(n7148), .ZN(n7520) );
  NAND2_X1 U7321 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6541), .ZN(n7509) );
  NOR2_X1 U7322 ( .A1(n7520), .A2(n7509), .ZN(n6545) );
  INV_X1 U7323 ( .A(n6542), .ZN(n6543) );
  NAND2_X1 U7324 ( .A1(n6545), .A2(n6543), .ZN(n7527) );
  NOR2_X1 U7325 ( .A1(n7527), .A2(n7149), .ZN(n6552) );
  INV_X1 U7326 ( .A(n6552), .ZN(n6544) );
  OR2_X1 U7327 ( .A1(n7474), .A2(n6544), .ZN(n6548) );
  NAND2_X1 U7328 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n6545), .ZN(n7541) );
  NOR2_X1 U7329 ( .A1(n7541), .A2(n6546), .ZN(n7531) );
  NAND2_X1 U7330 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n7531), .ZN(n6549) );
  OR2_X1 U7331 ( .A1(n7530), .A2(n6549), .ZN(n6547) );
  NAND2_X1 U7332 ( .A1(n6548), .A2(n6547), .ZN(n7120) );
  NAND3_X1 U7333 ( .A1(n7120), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n7111), .ZN(n6557) );
  NAND2_X1 U7334 ( .A1(n6550), .A2(n6549), .ZN(n7141) );
  AOI21_X1 U7335 ( .B1(n7119), .B2(n7141), .A(n6580), .ZN(n6554) );
  INV_X1 U7336 ( .A(n7528), .ZN(n6553) );
  INV_X1 U7337 ( .A(n7526), .ZN(n6551) );
  OAI21_X1 U7338 ( .B1(n6553), .B2(n6552), .A(n6551), .ZN(n7140) );
  NOR2_X1 U7339 ( .A1(n6554), .A2(n7140), .ZN(n7133) );
  OAI21_X1 U7340 ( .B1(n7121), .B2(n6580), .A(n7133), .ZN(n7114) );
  AOI21_X1 U7341 ( .B1(n7474), .B2(n7530), .A(n6555), .ZN(n6556) );
  NOR2_X1 U7342 ( .A1(n7114), .A2(n6556), .ZN(n7104) );
  AOI21_X1 U7343 ( .B1(n6558), .B2(n6557), .A(n7104), .ZN(n6559) );
  AOI211_X1 U7344 ( .C1(n6888), .C2(n7545), .A(n6565), .B(n6559), .ZN(n6560)
         );
  OAI21_X1 U7345 ( .B1(n6569), .B2(n7506), .A(n6560), .ZN(U2994) );
  BUF_X1 U7346 ( .A(n6561), .Z(n6562) );
  AOI21_X1 U7347 ( .B1(n6564), .B2(n6562), .A(n6563), .ZN(n6933) );
  AOI21_X1 U7348 ( .B1(n7415), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n6565), 
        .ZN(n6566) );
  OAI21_X1 U7349 ( .B1(n6749), .B2(n7425), .A(n6566), .ZN(n6567) );
  AOI21_X1 U7350 ( .B1(n6933), .B2(n7421), .A(n6567), .ZN(n6568) );
  OAI21_X1 U7351 ( .B1(n6569), .B2(n7701), .A(n6568), .ZN(U2962) );
  INV_X1 U7352 ( .A(n6570), .ZN(n6574) );
  NAND4_X1 U7353 ( .A1(n4252), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_28__SCAN_IN), .A4(INSTADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n6573) );
  INV_X1 U7354 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n7060) );
  NAND4_X1 U7355 ( .A1(n6571), .A2(n3631), .A3(n6581), .A4(n7060), .ZN(n6572)
         );
  XNOR2_X1 U7356 ( .A(n6575), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n6669)
         );
  INV_X1 U7357 ( .A(n6576), .ZN(n6577) );
  NAND2_X1 U7358 ( .A1(n7120), .A2(n6577), .ZN(n7092) );
  NOR2_X1 U7359 ( .A1(n7092), .A2(n6578), .ZN(n7073) );
  NOR3_X1 U7360 ( .A1(n7063), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n7060), 
        .ZN(n6583) );
  INV_X1 U7361 ( .A(REIP_REG_31__SCAN_IN), .ZN(n7335) );
  NOR2_X1 U7362 ( .A1(n7524), .A2(n7335), .ZN(n6664) );
  INV_X1 U7363 ( .A(n6598), .ZN(n7071) );
  INV_X1 U7364 ( .A(n6578), .ZN(n6579) );
  OAI21_X1 U7365 ( .B1(n6580), .B2(n6579), .A(n7104), .ZN(n7085) );
  NOR2_X1 U7366 ( .A1(n7085), .A2(n7508), .ZN(n7061) );
  INV_X1 U7367 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n6652) );
  AOI211_X1 U7368 ( .C1(n7062), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n7061), .B(n6652), .ZN(n6582) );
  AOI211_X1 U7369 ( .C1(n7073), .C2(n6583), .A(n6664), .B(n6582), .ZN(n6597)
         );
  OR2_X1 U7370 ( .A1(n6587), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6585)
         );
  INV_X1 U7371 ( .A(EBX_REG_30__SCAN_IN), .ZN(n6884) );
  NAND2_X1 U7372 ( .A1(n6680), .A2(n6884), .ZN(n6584) );
  NAND2_X1 U7373 ( .A1(n6585), .A2(n6584), .ZN(n6610) );
  MUX2_X2 U7374 ( .A(n6610), .B(n6586), .S(n6607), .Z(n6591) );
  OR2_X1 U7375 ( .A1(n6587), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n6589)
         );
  NAND2_X1 U7376 ( .A1(n6680), .A2(n6882), .ZN(n6588) );
  NAND2_X1 U7377 ( .A1(n6589), .A2(n6588), .ZN(n6592) );
  INV_X1 U7378 ( .A(n6592), .ZN(n6590) );
  NOR2_X1 U7379 ( .A1(n6607), .A2(n6610), .ZN(n6593) );
  NAND2_X1 U7380 ( .A1(n6881), .A2(n7545), .ZN(n6596) );
  OAI211_X1 U7381 ( .C1(n6669), .C2(n7506), .A(n6597), .B(n6596), .ZN(U2987)
         );
  INV_X1 U7382 ( .A(n6705), .ZN(n6602) );
  AOI21_X1 U7383 ( .B1(n7073), .B2(n6598), .A(INSTADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n6599) );
  NOR2_X1 U7384 ( .A1(n7062), .A2(n6599), .ZN(n6600) );
  AOI211_X1 U7385 ( .C1(n6602), .C2(n7545), .A(n6601), .B(n6600), .ZN(n6603)
         );
  OAI21_X1 U7386 ( .B1(n6604), .B2(n7506), .A(n6603), .ZN(U2989) );
  INV_X1 U7387 ( .A(n6605), .ZN(n6606) );
  INV_X1 U7388 ( .A(n6610), .ZN(n6611) );
  NAND2_X1 U7389 ( .A1(REIP_REG_29__SCAN_IN), .A2(REIP_REG_30__SCAN_IN), .ZN(
        n6617) );
  NAND4_X1 U7390 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_23__SCAN_IN), .A3(
        REIP_REG_26__SCAN_IN), .A4(REIP_REG_25__SCAN_IN), .ZN(n6633) );
  NAND4_X1 U7391 ( .A1(REIP_REG_21__SCAN_IN), .A2(REIP_REG_20__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .A4(REIP_REG_19__SCAN_IN), .ZN(n6779) );
  NOR3_X1 U7392 ( .A1(n7318), .A2(n6613), .A3(n6779), .ZN(n6618) );
  NAND2_X1 U7393 ( .A1(n6618), .A2(n6871), .ZN(n6741) );
  OR2_X1 U7394 ( .A1(n6633), .A2(n6741), .ZN(n6614) );
  NAND2_X1 U7395 ( .A1(n7598), .A2(n6614), .ZN(n6728) );
  INV_X1 U7396 ( .A(REIP_REG_27__SCAN_IN), .ZN(n7330) );
  OR2_X1 U7397 ( .A1(n7332), .A2(n7330), .ZN(n6615) );
  NAND2_X1 U7398 ( .A1(n7598), .A2(n6615), .ZN(n6616) );
  NAND2_X1 U7399 ( .A1(n6728), .A2(n6616), .ZN(n6702) );
  AOI21_X1 U7400 ( .B1(n6876), .B2(n6617), .A(n6702), .ZN(n6692) );
  INV_X1 U7401 ( .A(n6618), .ZN(n6619) );
  NOR2_X1 U7402 ( .A1(n6808), .A2(n6619), .ZN(n6740) );
  INV_X1 U7403 ( .A(n6633), .ZN(n6620) );
  NAND2_X1 U7404 ( .A1(n6740), .A2(n6620), .ZN(n6716) );
  OR3_X1 U7405 ( .A1(n6716), .A2(n7330), .A3(n7332), .ZN(n6688) );
  INV_X1 U7406 ( .A(n6688), .ZN(n6701) );
  NAND3_X1 U7407 ( .A1(n6701), .A2(REIP_REG_29__SCAN_IN), .A3(n7337), .ZN(
        n6624) );
  INV_X1 U7408 ( .A(n6621), .ZN(n6622) );
  AOI22_X1 U7409 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n7688), .B1(n7682), 
        .B2(n6622), .ZN(n6623) );
  OAI211_X1 U7410 ( .C1(n6884), .C2(n7686), .A(n6624), .B(n6623), .ZN(n6625)
         );
  INV_X1 U7411 ( .A(n6625), .ZN(n6626) );
  INV_X1 U7412 ( .A(n5333), .ZN(n6628) );
  OAI21_X1 U7413 ( .B1(n6629), .B2(n6627), .A(n6628), .ZN(n7070) );
  NAND2_X1 U7414 ( .A1(n6630), .A2(n7696), .ZN(n6637) );
  INV_X1 U7415 ( .A(EBX_REG_28__SCAN_IN), .ZN(n6641) );
  AOI22_X1 U7416 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n7688), .B1(n7682), 
        .B2(n6631), .ZN(n6632) );
  OAI21_X1 U7417 ( .B1(n7686), .B2(n6641), .A(n6632), .ZN(n6635) );
  INV_X1 U7418 ( .A(n6740), .ZN(n6765) );
  NOR4_X1 U7419 ( .A1(n6765), .A2(REIP_REG_28__SCAN_IN), .A3(n6633), .A4(n7330), .ZN(n6634) );
  AOI211_X1 U7420 ( .C1(REIP_REG_28__SCAN_IN), .C2(n6702), .A(n6635), .B(n6634), .ZN(n6636) );
  OAI211_X1 U7421 ( .C1(n7070), .C2(n7693), .A(n6637), .B(n6636), .ZN(U2799)
         );
  AOI22_X1 U7422 ( .A1(n7759), .A2(DATAI_29_), .B1(n7762), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n6639) );
  NAND2_X1 U7423 ( .A1(n7763), .A2(DATAI_13_), .ZN(n6638) );
  OAI211_X1 U7424 ( .C1(n6640), .C2(n7751), .A(n6639), .B(n6638), .ZN(U2862)
         );
  OAI222_X1 U7425 ( .A1(n6641), .A2(n7369), .B1(n6917), .B2(n7070), .C1(n6925), 
        .C2(n6919), .ZN(U2831) );
  OR2_X1 U7426 ( .A1(n7190), .A2(n7211), .ZN(n6644) );
  NAND2_X1 U7427 ( .A1(n6642), .A2(FLUSH_REG_SCAN_IN), .ZN(n6643) );
  NAND2_X1 U7428 ( .A1(n6644), .A2(n6643), .ZN(n7706) );
  AOI21_X1 U7429 ( .B1(n6646), .B2(n7713), .A(n7704), .ZN(n6651) );
  INV_X1 U7430 ( .A(n7168), .ZN(n6647) );
  OAI22_X1 U7431 ( .A1(n6648), .A2(n6647), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n7166), .ZN(n7186) );
  OAI22_X1 U7432 ( .A1(n7177), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n7715), .ZN(n6649) );
  AOI21_X1 U7433 ( .B1(n7186), .B2(n7713), .A(n6649), .ZN(n6650) );
  OAI22_X1 U7434 ( .A1(n6651), .A2(n4279), .B1(n7704), .B2(n6650), .ZN(U3461)
         );
  AOI21_X1 U7435 ( .B1(n7218), .B2(n7164), .A(n7704), .ZN(n6658) );
  AOI22_X1 U7436 ( .A1(INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n6653), .B1(
        INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n6652), .ZN(n7171) );
  NOR3_X1 U7437 ( .A1(n7715), .A2(n7562), .A3(n7171), .ZN(n6656) );
  NOR3_X1 U7438 ( .A1(n7177), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n7164), 
        .ZN(n6655) );
  AOI211_X1 U7439 ( .C1(n7185), .C2(n7713), .A(n6656), .B(n6655), .ZN(n6657)
         );
  OAI22_X1 U7440 ( .A1(n6658), .A2(n3720), .B1(n7704), .B2(n6657), .ZN(U3459)
         );
  AOI22_X1 U7441 ( .A1(n6660), .A2(EAX_REG_31__SCAN_IN), .B1(n6659), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n6661) );
  INV_X1 U7442 ( .A(n6661), .ZN(n6662) );
  XNOR2_X2 U7443 ( .A(n6663), .B(n6662), .ZN(n6685) );
  AOI21_X1 U7444 ( .B1(n7415), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n6664), 
        .ZN(n6665) );
  OAI21_X1 U7445 ( .B1(n6666), .B2(n7425), .A(n6665), .ZN(n6667) );
  OAI21_X1 U7446 ( .B1(n6669), .B2(n7701), .A(n6668), .ZN(U2955) );
  NAND3_X1 U7447 ( .A1(n6685), .A2(n6670), .A3(n6952), .ZN(n6672) );
  AOI22_X1 U7448 ( .A1(n7759), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n7762), .ZN(n6671) );
  NAND2_X1 U7449 ( .A1(n6672), .A2(n6671), .ZN(U2860) );
  NAND3_X1 U7450 ( .A1(n6673), .A2(n5111), .A3(n7200), .ZN(n6676) );
  INV_X1 U7451 ( .A(n6674), .ZN(n6675) );
  AOI22_X1 U7452 ( .A1(n6679), .A2(n6676), .B1(n3945), .B2(n6675), .ZN(n6677)
         );
  OAI21_X1 U7453 ( .B1(n6679), .B2(n6678), .A(n6677), .ZN(n7203) );
  NOR2_X1 U7454 ( .A1(n6681), .A2(n6680), .ZN(n7430) );
  INV_X1 U7455 ( .A(n7430), .ZN(n6683) );
  OAI21_X1 U7456 ( .B1(n6683), .B2(n6682), .A(n7442), .ZN(n7445) );
  NAND2_X1 U7457 ( .A1(n6684), .A2(n7445), .ZN(n7201) );
  AND2_X1 U7458 ( .A1(n7201), .A2(n7711), .ZN(n7703) );
  MUX2_X1 U7459 ( .A(MORE_REG_SCAN_IN), .B(n7203), .S(n7703), .Z(U3471) );
  INV_X1 U7460 ( .A(n6685), .ZN(n6695) );
  NOR2_X1 U7461 ( .A1(n6687), .A2(n6686), .ZN(n6690) );
  NOR4_X1 U7462 ( .A1(n6688), .A2(REIP_REG_31__SCAN_IN), .A3(n7337), .A4(n7333), .ZN(n6689) );
  AOI211_X1 U7463 ( .C1(PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n7688), .A(n6690), 
        .B(n6689), .ZN(n6691) );
  OAI21_X1 U7464 ( .B1(n6692), .B2(n7335), .A(n6691), .ZN(n6693) );
  OAI21_X1 U7465 ( .B1(n6695), .B2(n7679), .A(n6694), .ZN(U2796) );
  NAND2_X1 U7466 ( .A1(n7688), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n6698)
         );
  NAND2_X1 U7467 ( .A1(n7682), .A2(n6696), .ZN(n6697) );
  OAI211_X1 U7468 ( .C1(n7686), .C2(n6699), .A(n6698), .B(n6697), .ZN(n6700)
         );
  AOI21_X1 U7469 ( .B1(n6701), .B2(n7333), .A(n6700), .ZN(n6704) );
  NAND2_X1 U7470 ( .A1(n6702), .A2(REIP_REG_29__SCAN_IN), .ZN(n6703) );
  OAI211_X1 U7471 ( .C1(n6705), .C2(n7693), .A(n6704), .B(n6703), .ZN(n6706)
         );
  AOI21_X1 U7472 ( .B1(n6707), .B2(n7696), .A(n6706), .ZN(n6708) );
  INV_X1 U7473 ( .A(n6708), .ZN(U2798) );
  AOI21_X1 U7474 ( .B1(n6711), .B2(n6709), .A(n6710), .ZN(n6958) );
  INV_X1 U7475 ( .A(n6958), .ZN(n6928) );
  AOI21_X1 U7476 ( .B1(n6712), .B2(n6723), .A(n6627), .ZN(n7086) );
  NOR2_X1 U7477 ( .A1(n6728), .A2(n7330), .ZN(n6718) );
  AOI22_X1 U7478 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n7688), .B1(n7682), 
        .B2(n6961), .ZN(n6715) );
  OR2_X1 U7479 ( .A1(n7686), .A2(n6713), .ZN(n6714) );
  OAI211_X1 U7480 ( .C1(n6716), .C2(REIP_REG_27__SCAN_IN), .A(n6715), .B(n6714), .ZN(n6717) );
  AOI211_X1 U7481 ( .C1(n7086), .C2(n7666), .A(n6718), .B(n6717), .ZN(n6719)
         );
  OAI21_X1 U7482 ( .B1(n6928), .B2(n7679), .A(n6719), .ZN(U2800) );
  NAND2_X1 U7483 ( .A1(n6720), .A2(n6721), .ZN(n6722) );
  NAND2_X1 U7484 ( .A1(n6723), .A2(n6722), .ZN(n7098) );
  OAI21_X1 U7485 ( .B1(n6725), .B2(n6724), .A(n6709), .ZN(n6970) );
  INV_X1 U7486 ( .A(n6970), .ZN(n6726) );
  NAND2_X1 U7487 ( .A1(n6726), .A2(n7696), .ZN(n6733) );
  OAI22_X1 U7488 ( .A1(n6727), .A2(n7633), .B1(n7699), .B2(n6964), .ZN(n6731)
         );
  NOR3_X1 U7489 ( .A1(n6765), .A2(n7323), .A3(n7322), .ZN(n6746) );
  AOI21_X1 U7490 ( .B1(n6746), .B2(REIP_REG_25__SCAN_IN), .A(
        REIP_REG_26__SCAN_IN), .ZN(n6729) );
  NOR2_X1 U7491 ( .A1(n6729), .A2(n6728), .ZN(n6730) );
  AOI211_X1 U7492 ( .C1(EBX_REG_26__SCAN_IN), .C2(n7687), .A(n6731), .B(n6730), 
        .ZN(n6732) );
  OAI211_X1 U7493 ( .C1(n7098), .C2(n7693), .A(n6733), .B(n6732), .ZN(U2801)
         );
  OAI21_X1 U7494 ( .B1(n6735), .B2(n6734), .A(n6720), .ZN(n7100) );
  OAI21_X1 U7495 ( .B1(n6563), .B2(n6737), .A(n6736), .ZN(n6979) );
  INV_X1 U7496 ( .A(n6979), .ZN(n6738) );
  NAND2_X1 U7497 ( .A1(n6738), .A2(n7696), .ZN(n6748) );
  AOI22_X1 U7498 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n7688), .B1(n7682), 
        .B2(n6973), .ZN(n6739) );
  OAI21_X1 U7499 ( .B1(n7686), .B2(n6887), .A(n6739), .ZN(n6745) );
  NAND3_X1 U7500 ( .A1(n6740), .A2(REIP_REG_23__SCAN_IN), .A3(n7323), .ZN(
        n6752) );
  INV_X1 U7501 ( .A(n6741), .ZN(n6742) );
  NAND2_X1 U7502 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6742), .ZN(n6743) );
  NAND2_X1 U7503 ( .A1(n7598), .A2(n6743), .ZN(n6764) );
  AOI21_X1 U7504 ( .B1(n6752), .B2(n6764), .A(n7326), .ZN(n6744) );
  AOI211_X1 U7505 ( .C1(n6746), .C2(n7326), .A(n6745), .B(n6744), .ZN(n6747)
         );
  OAI211_X1 U7506 ( .C1(n7100), .C2(n7693), .A(n6748), .B(n6747), .ZN(U2802)
         );
  INV_X1 U7507 ( .A(n6933), .ZN(n6890) );
  OAI22_X1 U7508 ( .A1(n6750), .A2(n7633), .B1(n7699), .B2(n6749), .ZN(n6751)
         );
  AOI21_X1 U7509 ( .B1(n7687), .B2(EBX_REG_24__SCAN_IN), .A(n6751), .ZN(n6753)
         );
  OAI211_X1 U7510 ( .C1(n6764), .C2(n7323), .A(n6753), .B(n6752), .ZN(n6754)
         );
  AOI21_X1 U7511 ( .B1(n6888), .B2(n7666), .A(n6754), .ZN(n6755) );
  OAI21_X1 U7512 ( .B1(n6890), .B2(n7679), .A(n6755), .ZN(U2803) );
  NAND2_X1 U7513 ( .A1(n6773), .A2(n6756), .ZN(n6757) );
  NAND2_X1 U7514 ( .A1(n6758), .A2(n6757), .ZN(n7117) );
  INV_X1 U7515 ( .A(n6759), .ZN(n6761) );
  OAI21_X1 U7516 ( .B1(n6761), .B2(n4610), .A(n6562), .ZN(n6990) );
  INV_X1 U7517 ( .A(n6990), .ZN(n6762) );
  NAND2_X1 U7518 ( .A1(n6762), .A2(n7696), .ZN(n6769) );
  INV_X1 U7519 ( .A(n6987), .ZN(n6763) );
  OAI22_X1 U7520 ( .A1(n6985), .A2(n7633), .B1(n7699), .B2(n6763), .ZN(n6767)
         );
  AOI21_X1 U7521 ( .B1(n6765), .B2(n7322), .A(n6764), .ZN(n6766) );
  AOI211_X1 U7522 ( .C1(n7687), .C2(EBX_REG_23__SCAN_IN), .A(n6767), .B(n6766), 
        .ZN(n6768) );
  OAI211_X1 U7523 ( .C1(n7117), .C2(n7693), .A(n6769), .B(n6768), .ZN(U2804)
         );
  OAI21_X1 U7524 ( .B1(n5109), .B2(n6770), .A(n6759), .ZN(n6997) );
  NAND2_X1 U7525 ( .A1(n7672), .A2(n7318), .ZN(n6780) );
  INV_X1 U7526 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6771) );
  OAI22_X1 U7527 ( .A1(n6771), .A2(n7633), .B1(n7699), .B2(n6993), .ZN(n6777)
         );
  INV_X1 U7528 ( .A(n5307), .ZN(n6775) );
  INV_X1 U7529 ( .A(n6772), .ZN(n6774) );
  OAI21_X1 U7530 ( .B1(n6775), .B2(n6774), .A(n6773), .ZN(n7128) );
  NOR2_X1 U7531 ( .A1(n7128), .A2(n7693), .ZN(n6776) );
  AOI211_X1 U7532 ( .C1(EBX_REG_22__SCAN_IN), .C2(n7687), .A(n6777), .B(n6776), 
        .ZN(n6778) );
  OAI21_X1 U7533 ( .B1(n6780), .B2(n6779), .A(n6778), .ZN(n6784) );
  INV_X1 U7534 ( .A(n7692), .ZN(n6781) );
  AOI21_X1 U7535 ( .B1(n6782), .B2(n6781), .A(n7318), .ZN(n6783) );
  NOR2_X1 U7536 ( .A1(n6784), .A2(n6783), .ZN(n6785) );
  OAI21_X1 U7537 ( .B1(n6997), .B2(n7679), .A(n6785), .ZN(U2805) );
  INV_X1 U7538 ( .A(n6787), .ZN(n6788) );
  OAI21_X1 U7539 ( .B1(n6789), .B2(n6786), .A(n6787), .ZN(n7027) );
  NOR2_X1 U7540 ( .A1(n6844), .A2(n6790), .ZN(n7670) );
  NAND2_X1 U7541 ( .A1(n7311), .A2(n6791), .ZN(n6793) );
  OAI22_X1 U7542 ( .A1(n7026), .A2(n7633), .B1(n6909), .B2(n7686), .ZN(n6792)
         );
  AOI211_X1 U7543 ( .C1(n7670), .C2(n6793), .A(n7677), .B(n6792), .ZN(n6799)
         );
  OR2_X1 U7544 ( .A1(n6795), .A2(n6796), .ZN(n6797) );
  AND2_X1 U7545 ( .A1(n6794), .A2(n6797), .ZN(n7533) );
  AOI22_X1 U7546 ( .A1(n7533), .A2(n7666), .B1(n7682), .B2(n7030), .ZN(n6798)
         );
  OAI211_X1 U7547 ( .C1(n7027), .C2(n7679), .A(n6799), .B(n6798), .ZN(U2810)
         );
  AND2_X1 U7548 ( .A1(n6800), .A2(n6801), .ZN(n6802) );
  OR2_X1 U7549 ( .A1(n6802), .A2(n6786), .ZN(n7752) );
  INV_X1 U7550 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6812) );
  INV_X1 U7551 ( .A(n6809), .ZN(n6805) );
  INV_X1 U7552 ( .A(n6842), .ZN(n6803) );
  OR2_X1 U7553 ( .A1(n6808), .A2(n6803), .ZN(n6804) );
  AND2_X1 U7554 ( .A1(n6804), .A2(n6871), .ZN(n7574) );
  OAI21_X1 U7555 ( .B1(n6805), .B2(n6844), .A(n7574), .ZN(n6835) );
  INV_X1 U7556 ( .A(n6806), .ZN(n6807) );
  NOR2_X1 U7557 ( .A1(n6808), .A2(n6807), .ZN(n7563) );
  NOR2_X1 U7558 ( .A1(n6809), .A2(n7618), .ZN(n6826) );
  XOR2_X1 U7559 ( .A(n7525), .B(n7308), .Z(n6810) );
  AOI22_X1 U7560 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6835), .B1(n6826), .B2(
        n6810), .ZN(n6811) );
  OAI211_X1 U7561 ( .C1(n7633), .C2(n6812), .A(n6811), .B(n7648), .ZN(n6818)
         );
  NOR2_X1 U7562 ( .A1(n6813), .A2(n6814), .ZN(n6815) );
  OR2_X1 U7563 ( .A1(n6795), .A2(n6815), .ZN(n7515) );
  AOI22_X1 U7564 ( .A1(n7687), .A2(EBX_REG_16__SCAN_IN), .B1(n7682), .B2(n7038), .ZN(n6816) );
  OAI21_X1 U7565 ( .B1(n7515), .B2(n7693), .A(n6816), .ZN(n6817) );
  NOR2_X1 U7566 ( .A1(n6818), .A2(n6817), .ZN(n6819) );
  OAI21_X1 U7567 ( .B1(n7752), .B2(n7679), .A(n6819), .ZN(U2811) );
  INV_X1 U7568 ( .A(n6800), .ZN(n6821) );
  AOI21_X1 U7569 ( .B1(n6822), .B2(n6820), .A(n6821), .ZN(n7047) );
  INV_X1 U7570 ( .A(n7047), .ZN(n6951) );
  AOI22_X1 U7571 ( .A1(EBX_REG_15__SCAN_IN), .A2(n7687), .B1(
        REIP_REG_15__SCAN_IN), .B2(n6835), .ZN(n6823) );
  OAI211_X1 U7572 ( .C1(n7633), .C2(n6824), .A(n6823), .B(n7648), .ZN(n6825)
         );
  AOI21_X1 U7573 ( .B1(n6826), .B2(n7308), .A(n6825), .ZN(n6831) );
  AOI21_X1 U7574 ( .B1(n6828), .B2(n6827), .A(n6813), .ZN(n7510) );
  INV_X1 U7575 ( .A(n7045), .ZN(n6829) );
  AOI22_X1 U7576 ( .A1(n7510), .A2(n7666), .B1(n7682), .B2(n6829), .ZN(n6830)
         );
  OAI211_X1 U7577 ( .C1(n6951), .C2(n7679), .A(n6831), .B(n6830), .ZN(U2812)
         );
  OAI21_X1 U7578 ( .B1(n6833), .B2(n6832), .A(n6820), .ZN(n7053) );
  INV_X1 U7579 ( .A(n6916), .ZN(n6840) );
  INV_X1 U7580 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n7051) );
  NAND2_X1 U7581 ( .A1(n7682), .A2(n7056), .ZN(n6834) );
  OAI211_X1 U7582 ( .C1(n7633), .C2(n7051), .A(n6834), .B(n7648), .ZN(n6839)
         );
  NAND2_X1 U7583 ( .A1(n6846), .A2(n7599), .ZN(n6849) );
  INV_X1 U7584 ( .A(n6849), .ZN(n7646) );
  NAND3_X1 U7585 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .A3(
        n7646), .ZN(n6837) );
  AOI22_X1 U7586 ( .A1(EBX_REG_14__SCAN_IN), .A2(n7687), .B1(
        REIP_REG_14__SCAN_IN), .B2(n6835), .ZN(n6836) );
  OAI21_X1 U7587 ( .B1(REIP_REG_14__SCAN_IN), .B2(n6837), .A(n6836), .ZN(n6838) );
  AOI211_X1 U7588 ( .C1(n6840), .C2(n7666), .A(n6839), .B(n6838), .ZN(n6841)
         );
  OAI21_X1 U7589 ( .B1(n7053), .B2(n7679), .A(n6841), .ZN(U2813) );
  NOR2_X1 U7590 ( .A1(n6843), .A2(n6842), .ZN(n6845) );
  AOI21_X1 U7591 ( .B1(n6846), .B2(n6845), .A(n6844), .ZN(n7657) );
  AOI22_X1 U7592 ( .A1(EBX_REG_12__SCAN_IN), .A2(n7687), .B1(
        REIP_REG_12__SCAN_IN), .B2(n7657), .ZN(n6847) );
  OAI211_X1 U7593 ( .C1(n7633), .C2(n6848), .A(n6847), .B(n7648), .ZN(n6853)
         );
  NOR2_X1 U7594 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6849), .ZN(n7658) );
  INV_X1 U7595 ( .A(n6850), .ZN(n6851) );
  OAI22_X1 U7596 ( .A1(n7493), .A2(n7693), .B1(n6851), .B2(n7699), .ZN(n6852)
         );
  NOR3_X1 U7597 ( .A1(n6853), .A2(n7658), .A3(n6852), .ZN(n6854) );
  OAI21_X1 U7598 ( .B1(n6855), .B2(n7679), .A(n6854), .ZN(U2815) );
  NOR2_X1 U7599 ( .A1(n7686), .A2(n6856), .ZN(n6860) );
  OAI22_X1 U7600 ( .A1(n6858), .A2(n7633), .B1(n7699), .B2(n6857), .ZN(n6859)
         );
  AOI211_X1 U7601 ( .C1(n6874), .C2(n3645), .A(n6860), .B(n6859), .ZN(n6861)
         );
  OAI21_X1 U7602 ( .B1(n7693), .B2(n6862), .A(n6861), .ZN(n6866) );
  AOI21_X1 U7603 ( .B1(n7290), .B2(n6864), .A(n6863), .ZN(n6865) );
  INV_X1 U7604 ( .A(n6868), .ZN(U2824) );
  INV_X1 U7605 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6870) );
  AOI22_X1 U7606 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n7688), .B1(n7666), 
        .B2(n7468), .ZN(n6869) );
  OAI21_X1 U7607 ( .B1(n6871), .B2(n6870), .A(n6869), .ZN(n6873) );
  NOR2_X1 U7608 ( .A1(n7699), .A2(n7381), .ZN(n6872) );
  AOI211_X1 U7609 ( .C1(n6874), .C2(n3663), .A(n6873), .B(n6872), .ZN(n6878)
         );
  MUX2_X1 U7610 ( .A(REIP_REG_2__SCAN_IN), .B(n6870), .S(REIP_REG_1__SCAN_IN), 
        .Z(n6875) );
  AOI22_X1 U7611 ( .A1(n7687), .A2(EBX_REG_2__SCAN_IN), .B1(n6876), .B2(n6875), 
        .ZN(n6877) );
  OAI211_X1 U7612 ( .C1(n6880), .C2(n6879), .A(n6878), .B(n6877), .ZN(U2825)
         );
  INV_X1 U7613 ( .A(n6881), .ZN(n6883) );
  OAI22_X1 U7614 ( .A1(n6883), .A2(n6917), .B1(n6882), .B2(n7369), .ZN(U2828)
         );
  OAI222_X1 U7615 ( .A1(n6884), .A2(n7369), .B1(n6917), .B2(n7069), .C1(n6919), 
        .C2(n6922), .ZN(U2829) );
  AOI22_X1 U7616 ( .A1(n7086), .A2(n6914), .B1(n6913), .B2(EBX_REG_27__SCAN_IN), .ZN(n6885) );
  OAI21_X1 U7617 ( .B1(n6928), .B2(n6919), .A(n6885), .ZN(U2832) );
  INV_X1 U7618 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6886) );
  OAI222_X1 U7619 ( .A1(n6886), .A2(n7369), .B1(n6917), .B2(n7098), .C1(n6970), 
        .C2(n6919), .ZN(U2833) );
  OAI222_X1 U7620 ( .A1(n7100), .A2(n6917), .B1(n6887), .B2(n7369), .C1(n6979), 
        .C2(n6919), .ZN(U2834) );
  AOI22_X1 U7621 ( .A1(n6888), .A2(n6914), .B1(n6913), .B2(EBX_REG_24__SCAN_IN), .ZN(n6889) );
  OAI21_X1 U7622 ( .B1(n6890), .B2(n6919), .A(n6889), .ZN(U2835) );
  OAI22_X1 U7623 ( .A1(n7117), .A2(n6917), .B1(n6891), .B2(n7369), .ZN(n6892)
         );
  INV_X1 U7624 ( .A(n6892), .ZN(n6893) );
  OAI21_X1 U7625 ( .B1(n6990), .B2(n6919), .A(n6893), .ZN(U2836) );
  OAI222_X1 U7626 ( .A1(n6894), .A2(n7369), .B1(n6917), .B2(n7128), .C1(n6997), 
        .C2(n6919), .ZN(U2837) );
  INV_X1 U7627 ( .A(EBX_REG_21__SCAN_IN), .ZN(n6895) );
  INV_X1 U7628 ( .A(n6941), .ZN(n7006) );
  OAI222_X1 U7629 ( .A1(n6917), .A2(n7139), .B1(n7369), .B2(n6895), .C1(n7006), 
        .C2(n6919), .ZN(U2838) );
  INV_X1 U7630 ( .A(n6896), .ZN(n6907) );
  AND2_X1 U7631 ( .A1(n6907), .A2(n6897), .ZN(n6899) );
  OR2_X1 U7632 ( .A1(n6899), .A2(n6898), .ZN(n7678) );
  OAI21_X1 U7633 ( .B1(n6900), .B2(n6902), .A(n6901), .ZN(n7680) );
  OAI222_X1 U7634 ( .A1(n7678), .A2(n6917), .B1(n7369), .B2(n5187), .C1(n6919), 
        .C2(n7680), .ZN(U2840) );
  NOR2_X1 U7635 ( .A1(n6788), .A2(n6903), .ZN(n6904) );
  OR2_X1 U7636 ( .A1(n6900), .A2(n6904), .ZN(n7420) );
  NAND2_X1 U7637 ( .A1(n6794), .A2(n6905), .ZN(n6906) );
  AND2_X1 U7638 ( .A1(n6907), .A2(n6906), .ZN(n7665) );
  AOI22_X1 U7639 ( .A1(n7665), .A2(n6914), .B1(EBX_REG_18__SCAN_IN), .B2(n6913), .ZN(n6908) );
  OAI21_X1 U7640 ( .B1(n7420), .B2(n6919), .A(n6908), .ZN(U2841) );
  NOR2_X1 U7641 ( .A1(n7369), .A2(n6909), .ZN(n6910) );
  AOI21_X1 U7642 ( .B1(n7533), .B2(n6914), .A(n6910), .ZN(n6911) );
  OAI21_X1 U7643 ( .B1(n7027), .B2(n6919), .A(n6911), .ZN(U2842) );
  INV_X1 U7644 ( .A(EBX_REG_16__SCAN_IN), .ZN(n6912) );
  OAI222_X1 U7645 ( .A1(n7515), .A2(n6917), .B1(n6912), .B2(n7369), .C1(n7752), 
        .C2(n6919), .ZN(U2843) );
  AOI22_X1 U7646 ( .A1(n7510), .A2(n6914), .B1(n6913), .B2(EBX_REG_15__SCAN_IN), .ZN(n6915) );
  OAI21_X1 U7647 ( .B1(n6951), .B2(n6919), .A(n6915), .ZN(U2844) );
  INV_X1 U7648 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6918) );
  OAI222_X1 U7649 ( .A1(n7053), .A2(n6919), .B1(n7369), .B2(n6918), .C1(n6917), 
        .C2(n6916), .ZN(U2845) );
  AOI22_X1 U7650 ( .A1(n7759), .A2(DATAI_30_), .B1(n7762), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n6921) );
  NAND2_X1 U7651 ( .A1(n7763), .A2(DATAI_14_), .ZN(n6920) );
  OAI211_X1 U7652 ( .C1(n6922), .C2(n7751), .A(n6921), .B(n6920), .ZN(U2861)
         );
  AOI22_X1 U7653 ( .A1(n7759), .A2(DATAI_28_), .B1(n7762), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n6924) );
  NAND2_X1 U7654 ( .A1(n7763), .A2(DATAI_12_), .ZN(n6923) );
  OAI211_X1 U7655 ( .C1(n6925), .C2(n7751), .A(n6924), .B(n6923), .ZN(U2863)
         );
  AOI22_X1 U7656 ( .A1(n7759), .A2(DATAI_27_), .B1(n7762), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6927) );
  NAND2_X1 U7657 ( .A1(n7763), .A2(DATAI_11_), .ZN(n6926) );
  OAI211_X1 U7658 ( .C1(n6928), .C2(n7751), .A(n6927), .B(n6926), .ZN(U2864)
         );
  AOI22_X1 U7659 ( .A1(n7759), .A2(DATAI_26_), .B1(n7762), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n6930) );
  NAND2_X1 U7660 ( .A1(n7763), .A2(DATAI_10_), .ZN(n6929) );
  OAI211_X1 U7661 ( .C1(n6970), .C2(n7751), .A(n6930), .B(n6929), .ZN(U2865)
         );
  AOI22_X1 U7662 ( .A1(n7759), .A2(DATAI_25_), .B1(n7762), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6932) );
  NAND2_X1 U7663 ( .A1(n7763), .A2(DATAI_9_), .ZN(n6931) );
  OAI211_X1 U7664 ( .C1(n6979), .C2(n7751), .A(n6932), .B(n6931), .ZN(U2866)
         );
  INV_X1 U7665 ( .A(n7763), .ZN(n6945) );
  INV_X1 U7666 ( .A(n7751), .ZN(n7760) );
  NAND2_X1 U7667 ( .A1(n6933), .A2(n7760), .ZN(n6935) );
  AOI22_X1 U7668 ( .A1(n7759), .A2(DATAI_24_), .B1(n7762), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n6934) );
  OAI211_X1 U7669 ( .C1(n6945), .C2(n6936), .A(n6935), .B(n6934), .ZN(U2867)
         );
  AOI22_X1 U7670 ( .A1(n7759), .A2(DATAI_23_), .B1(n7762), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n6938) );
  NAND2_X1 U7671 ( .A1(n7763), .A2(DATAI_7_), .ZN(n6937) );
  OAI211_X1 U7672 ( .C1(n6990), .C2(n7751), .A(n6938), .B(n6937), .ZN(U2868)
         );
  AOI22_X1 U7673 ( .A1(n7759), .A2(DATAI_22_), .B1(n7762), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n6940) );
  NAND2_X1 U7674 ( .A1(n7763), .A2(DATAI_6_), .ZN(n6939) );
  OAI211_X1 U7675 ( .C1(n6997), .C2(n7751), .A(n6940), .B(n6939), .ZN(U2869)
         );
  NAND2_X1 U7676 ( .A1(n6941), .A2(n7760), .ZN(n6943) );
  AOI22_X1 U7677 ( .A1(n7759), .A2(DATAI_21_), .B1(n7762), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n6942) );
  OAI211_X1 U7678 ( .C1(n6945), .C2(n6944), .A(n6943), .B(n6942), .ZN(U2870)
         );
  AOI22_X1 U7679 ( .A1(n7759), .A2(DATAI_19_), .B1(n7762), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n6947) );
  NAND2_X1 U7680 ( .A1(n7763), .A2(DATAI_3_), .ZN(n6946) );
  OAI211_X1 U7681 ( .C1(n7680), .C2(n7751), .A(n6947), .B(n6946), .ZN(U2872)
         );
  AOI22_X1 U7682 ( .A1(n7759), .A2(DATAI_17_), .B1(n7762), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6949) );
  NAND2_X1 U7683 ( .A1(n7763), .A2(DATAI_1_), .ZN(n6948) );
  OAI211_X1 U7684 ( .C1(n7027), .C2(n7751), .A(n6949), .B(n6948), .ZN(U2874)
         );
  INV_X1 U7685 ( .A(EAX_REG_15__SCAN_IN), .ZN(n7287) );
  OAI222_X1 U7686 ( .A1(n6951), .A2(n7751), .B1(n6950), .B2(n6953), .C1(n6952), 
        .C2(n7287), .ZN(U2876) );
  INV_X1 U7687 ( .A(EAX_REG_14__SCAN_IN), .ZN(n7283) );
  OAI222_X1 U7688 ( .A1(n7053), .A2(n7751), .B1(n6954), .B2(n6953), .C1(n6952), 
        .C2(n7283), .ZN(U2877) );
  NOR2_X1 U7689 ( .A1(n4252), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6956)
         );
  MUX2_X1 U7690 ( .A(n4252), .B(n6956), .S(n6955), .Z(n6957) );
  XNOR2_X1 U7691 ( .A(n6957), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n7089)
         );
  NAND2_X1 U7692 ( .A1(n6958), .A2(n7421), .ZN(n6963) );
  NOR2_X1 U7693 ( .A1(n7524), .A2(n7330), .ZN(n7084) );
  NOR2_X1 U7694 ( .A1(n7405), .A2(n6959), .ZN(n6960) );
  AOI211_X1 U7695 ( .C1(n6961), .C2(n7409), .A(n7084), .B(n6960), .ZN(n6962)
         );
  OAI211_X1 U7696 ( .C1(n7089), .C2(n7701), .A(n6963), .B(n6962), .ZN(U2959)
         );
  INV_X1 U7697 ( .A(REIP_REG_26__SCAN_IN), .ZN(n7328) );
  NOR2_X1 U7698 ( .A1(n7524), .A2(n7328), .ZN(n7094) );
  NOR2_X1 U7699 ( .A1(n7425), .A2(n6964), .ZN(n6965) );
  AOI211_X1 U7700 ( .C1(n7415), .C2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n7094), 
        .B(n6965), .ZN(n6969) );
  XNOR2_X1 U7701 ( .A(n4252), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6967)
         );
  XNOR2_X1 U7702 ( .A(n6966), .B(n6967), .ZN(n7090) );
  NAND2_X1 U7703 ( .A1(n7090), .A2(n7422), .ZN(n6968) );
  OAI211_X1 U7704 ( .C1(n6970), .C2(n7052), .A(n6969), .B(n6968), .ZN(U2960)
         );
  OAI22_X1 U7705 ( .A1(n7405), .A2(n6971), .B1(n7524), .B2(n7326), .ZN(n6972)
         );
  AOI21_X1 U7706 ( .B1(n7409), .B2(n6973), .A(n6972), .ZN(n6978) );
  OAI21_X1 U7707 ( .B1(n6974), .B2(n6976), .A(n6975), .ZN(n7099) );
  NAND2_X1 U7708 ( .A1(n7099), .A2(n7422), .ZN(n6977) );
  OAI211_X1 U7709 ( .C1(n6979), .C2(n7052), .A(n6978), .B(n6977), .ZN(U2961)
         );
  INV_X1 U7710 ( .A(n6980), .ZN(n6981) );
  NAND2_X1 U7711 ( .A1(n6981), .A2(n7111), .ZN(n6983) );
  MUX2_X1 U7712 ( .A(n6983), .B(n6982), .S(n3631), .Z(n6984) );
  XNOR2_X1 U7713 ( .A(n6984), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n7109)
         );
  NAND2_X1 U7714 ( .A1(n7109), .A2(n7422), .ZN(n6989) );
  NOR2_X1 U7715 ( .A1(n7524), .A2(n7322), .ZN(n7113) );
  NOR2_X1 U7716 ( .A1(n7405), .A2(n6985), .ZN(n6986) );
  AOI211_X1 U7717 ( .C1(n7409), .C2(n6987), .A(n7113), .B(n6986), .ZN(n6988)
         );
  OAI211_X1 U7718 ( .C1(n7052), .C2(n6990), .A(n6989), .B(n6988), .ZN(U2963)
         );
  XNOR2_X1 U7719 ( .A(n4252), .B(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6991)
         );
  XNOR2_X1 U7720 ( .A(n6992), .B(n6991), .ZN(n7118) );
  NAND2_X1 U7721 ( .A1(n7118), .A2(n7422), .ZN(n6996) );
  NOR2_X1 U7722 ( .A1(n7524), .A2(n7318), .ZN(n7124) );
  NOR2_X1 U7723 ( .A1(n7425), .A2(n6993), .ZN(n6994) );
  AOI211_X1 U7724 ( .C1(n7415), .C2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n7124), 
        .B(n6994), .ZN(n6995) );
  OAI211_X1 U7725 ( .C1(n7052), .C2(n6997), .A(n6996), .B(n6995), .ZN(U2964)
         );
  INV_X1 U7726 ( .A(n6998), .ZN(n7130) );
  NAND2_X1 U7727 ( .A1(n7000), .A2(n6999), .ZN(n7129) );
  NAND3_X1 U7728 ( .A1(n7130), .A2(n7422), .A3(n7129), .ZN(n7005) );
  NAND2_X1 U7729 ( .A1(n7544), .A2(REIP_REG_21__SCAN_IN), .ZN(n7132) );
  OAI21_X1 U7730 ( .B1(n7405), .B2(n7001), .A(n7132), .ZN(n7002) );
  AOI21_X1 U7731 ( .B1(n7409), .B2(n7003), .A(n7002), .ZN(n7004) );
  OAI211_X1 U7732 ( .C1(n7006), .C2(n7052), .A(n7005), .B(n7004), .ZN(U2965)
         );
  NAND2_X1 U7733 ( .A1(n4252), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n7008) );
  MUX2_X1 U7734 ( .A(n4252), .B(n7008), .S(n7007), .Z(n7009) );
  XOR2_X1 U7735 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .B(n7009), .Z(n7155) );
  NOR2_X1 U7736 ( .A1(n7524), .A2(n7315), .ZN(n7147) );
  INV_X1 U7737 ( .A(n7147), .ZN(n7010) );
  OAI21_X1 U7738 ( .B1(n7405), .B2(n7011), .A(n7010), .ZN(n7012) );
  AOI21_X1 U7739 ( .B1(n7409), .B2(n7013), .A(n7012), .ZN(n7017) );
  NAND2_X1 U7740 ( .A1(n6901), .A2(n7014), .ZN(n7015) );
  AND2_X1 U7741 ( .A1(n5107), .A2(n7015), .ZN(n7761) );
  NAND2_X1 U7742 ( .A1(n7761), .A2(n7421), .ZN(n7016) );
  OAI211_X1 U7743 ( .C1(n7155), .C2(n7701), .A(n7017), .B(n7016), .ZN(U2966)
         );
  AOI21_X1 U7744 ( .B1(n7019), .B2(n7018), .A(n3625), .ZN(n7163) );
  INV_X1 U7745 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n7020) );
  OR2_X1 U7746 ( .A1(n7524), .A2(n7673), .ZN(n7158) );
  OAI21_X1 U7747 ( .B1(n7405), .B2(n7020), .A(n7158), .ZN(n7022) );
  NOR2_X1 U7748 ( .A1(n7680), .A2(n7052), .ZN(n7021) );
  AOI211_X1 U7749 ( .C1(n7409), .C2(n7683), .A(n7022), .B(n7021), .ZN(n7023)
         );
  OAI21_X1 U7750 ( .B1(n7163), .B2(n7701), .A(n7023), .ZN(U2967) );
  NAND2_X1 U7751 ( .A1(n7024), .A2(n7032), .ZN(n7418) );
  XNOR2_X1 U7752 ( .A(n4252), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n7025)
         );
  XNOR2_X1 U7753 ( .A(n7418), .B(n7025), .ZN(n7532) );
  OAI22_X1 U7754 ( .A1(n7405), .A2(n7026), .B1(n7524), .B2(n7311), .ZN(n7029)
         );
  NOR2_X1 U7755 ( .A1(n7027), .A2(n7052), .ZN(n7028) );
  AOI211_X1 U7756 ( .C1(n7409), .C2(n7030), .A(n7029), .B(n7028), .ZN(n7031)
         );
  OAI21_X1 U7757 ( .B1(n7532), .B2(n7701), .A(n7031), .ZN(U2969) );
  INV_X1 U7758 ( .A(n7032), .ZN(n7034) );
  NOR2_X1 U7759 ( .A1(n7034), .A2(n7033), .ZN(n7035) );
  XNOR2_X1 U7760 ( .A(n7036), .B(n7035), .ZN(n7519) );
  NAND2_X1 U7761 ( .A1(n7519), .A2(n7422), .ZN(n7040) );
  OAI22_X1 U7762 ( .A1(n7405), .A2(n6812), .B1(n7525), .B2(n7524), .ZN(n7037)
         );
  AOI21_X1 U7763 ( .B1(n7409), .B2(n7038), .A(n7037), .ZN(n7039) );
  OAI211_X1 U7764 ( .C1(n7052), .C2(n7752), .A(n7040), .B(n7039), .ZN(U2970)
         );
  NAND2_X1 U7765 ( .A1(n3677), .A2(n7041), .ZN(n7042) );
  XNOR2_X1 U7766 ( .A(n7043), .B(n7042), .ZN(n7511) );
  INV_X1 U7767 ( .A(n7511), .ZN(n7049) );
  AOI22_X1 U7768 ( .A1(n7415), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n7544), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n7044) );
  OAI21_X1 U7769 ( .B1(n7045), .B2(n7425), .A(n7044), .ZN(n7046) );
  AOI21_X1 U7770 ( .B1(n7047), .B2(n7421), .A(n7046), .ZN(n7048) );
  OAI21_X1 U7771 ( .B1(n7049), .B2(n7701), .A(n7048), .ZN(U2971) );
  OAI21_X1 U7772 ( .B1(n7405), .B2(n7051), .A(n7050), .ZN(n7055) );
  NOR2_X1 U7773 ( .A1(n7053), .A2(n7052), .ZN(n7054) );
  AOI211_X1 U7774 ( .C1(n7409), .C2(n7056), .A(n7055), .B(n7054), .ZN(n7057)
         );
  OAI21_X1 U7775 ( .B1(n7701), .B2(n7058), .A(n7057), .ZN(U2972) );
  NAND2_X1 U7776 ( .A1(n7059), .A2(n7557), .ZN(n7068) );
  NOR3_X1 U7777 ( .A1(n7062), .A2(n7061), .A3(n7060), .ZN(n7066) );
  INV_X1 U7778 ( .A(n7073), .ZN(n7082) );
  NOR3_X1 U7779 ( .A1(n7082), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n7063), 
        .ZN(n7064) );
  NOR3_X1 U7780 ( .A1(n7066), .A2(n7065), .A3(n7064), .ZN(n7067) );
  OAI211_X1 U7781 ( .C1(n7069), .C2(n7555), .A(n7068), .B(n7067), .ZN(U2988)
         );
  INV_X1 U7782 ( .A(n7070), .ZN(n7079) );
  INV_X1 U7783 ( .A(n7085), .ZN(n7077) );
  NAND3_X1 U7784 ( .A1(n7073), .A2(n7072), .A3(n7071), .ZN(n7074) );
  OAI211_X1 U7785 ( .C1(n7077), .C2(n7076), .A(n7075), .B(n7074), .ZN(n7078)
         );
  AOI21_X1 U7786 ( .B1(n7079), .B2(n7545), .A(n7078), .ZN(n7080) );
  OAI21_X1 U7787 ( .B1(n7081), .B2(n7506), .A(n7080), .ZN(U2990) );
  NOR2_X1 U7788 ( .A1(n7082), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n7083)
         );
  AOI211_X1 U7789 ( .C1(n7085), .C2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n7084), .B(n7083), .ZN(n7088) );
  NAND2_X1 U7790 ( .A1(n7086), .A2(n7545), .ZN(n7087) );
  OAI211_X1 U7791 ( .C1(n7089), .C2(n7506), .A(n7088), .B(n7087), .ZN(U2991)
         );
  NAND2_X1 U7792 ( .A1(n7090), .A2(n7557), .ZN(n7097) );
  OR2_X1 U7793 ( .A1(n7092), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n7101)
         );
  AOI21_X1 U7794 ( .B1(n7104), .B2(n7101), .A(n7091), .ZN(n7095) );
  NOR3_X1 U7795 ( .A1(n7092), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n7103), 
        .ZN(n7093) );
  NOR3_X1 U7796 ( .A1(n7095), .A2(n7094), .A3(n7093), .ZN(n7096) );
  OAI211_X1 U7797 ( .C1(n7555), .C2(n7098), .A(n7097), .B(n7096), .ZN(U2992)
         );
  INV_X1 U7798 ( .A(n7099), .ZN(n7108) );
  INV_X1 U7799 ( .A(n7100), .ZN(n7106) );
  NAND2_X1 U7800 ( .A1(n7544), .A2(REIP_REG_25__SCAN_IN), .ZN(n7102) );
  OAI211_X1 U7801 ( .C1(n7104), .C2(n7103), .A(n7102), .B(n7101), .ZN(n7105)
         );
  AOI21_X1 U7802 ( .B1(n7106), .B2(n7545), .A(n7105), .ZN(n7107) );
  OAI21_X1 U7803 ( .B1(n7108), .B2(n7506), .A(n7107), .ZN(U2993) );
  NAND2_X1 U7804 ( .A1(n7109), .A2(n7557), .ZN(n7116) );
  AND3_X1 U7805 ( .A1(n7120), .A2(n7111), .A3(n7110), .ZN(n7112) );
  AOI211_X1 U7806 ( .C1(n7114), .C2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n7113), .B(n7112), .ZN(n7115) );
  OAI211_X1 U7807 ( .C1(n7555), .C2(n7117), .A(n7116), .B(n7115), .ZN(U2995)
         );
  NAND2_X1 U7808 ( .A1(n7118), .A2(n7557), .ZN(n7127) );
  INV_X1 U7809 ( .A(n7133), .ZN(n7125) );
  NAND2_X1 U7810 ( .A1(n7120), .A2(n7119), .ZN(n7131) );
  NOR3_X1 U7811 ( .A1(n7131), .A2(n7122), .A3(n7121), .ZN(n7123) );
  AOI211_X1 U7812 ( .C1(n7125), .C2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n7124), .B(n7123), .ZN(n7126) );
  OAI211_X1 U7813 ( .C1(n7555), .C2(n7128), .A(n7127), .B(n7126), .ZN(U2996)
         );
  NAND3_X1 U7814 ( .A1(n7130), .A2(n7557), .A3(n7129), .ZN(n7138) );
  INV_X1 U7815 ( .A(n7131), .ZN(n7136) );
  OAI21_X1 U7816 ( .B1(n7133), .B2(n7135), .A(n7132), .ZN(n7134) );
  AOI21_X1 U7817 ( .B1(n7136), .B2(n7135), .A(n7134), .ZN(n7137) );
  OAI211_X1 U7818 ( .C1(n7555), .C2(n7139), .A(n7138), .B(n7137), .ZN(U2997)
         );
  INV_X1 U7819 ( .A(n7140), .ZN(n7142) );
  NAND2_X1 U7820 ( .A1(n7142), .A2(n7141), .ZN(n7156) );
  NOR2_X1 U7821 ( .A1(n6898), .A2(n7143), .ZN(n7144) );
  OR2_X1 U7822 ( .A1(n7145), .A2(n7144), .ZN(n7694) );
  NOR2_X1 U7823 ( .A1(n7694), .A2(n7555), .ZN(n7146) );
  AOI211_X1 U7824 ( .C1(INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n7156), .A(n7147), .B(n7146), .ZN(n7154) );
  NOR2_X1 U7825 ( .A1(n7542), .A2(n7509), .ZN(n7521) );
  NAND2_X1 U7826 ( .A1(n7148), .A2(n7521), .ZN(n7537) );
  NOR2_X1 U7827 ( .A1(n7537), .A2(n7149), .ZN(n7161) );
  INV_X1 U7828 ( .A(n7150), .ZN(n7151) );
  NAND3_X1 U7829 ( .A1(n7161), .A2(n7152), .A3(n7151), .ZN(n7153) );
  OAI211_X1 U7830 ( .C1(n7155), .C2(n7506), .A(n7154), .B(n7153), .ZN(U2998)
         );
  NAND2_X1 U7831 ( .A1(n7156), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n7157) );
  OAI211_X1 U7832 ( .C1(n7678), .C2(n7555), .A(n7158), .B(n7157), .ZN(n7159)
         );
  AOI21_X1 U7833 ( .B1(n7161), .B2(n7160), .A(n7159), .ZN(n7162) );
  OAI21_X1 U7834 ( .B1(n7163), .B2(n7506), .A(n7162), .ZN(U2999) );
  NAND2_X1 U7835 ( .A1(n7165), .A2(n7164), .ZN(n7170) );
  OAI22_X1 U7836 ( .A1(n7188), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(n7170), .B2(n7166), .ZN(n7167) );
  AOI21_X1 U7837 ( .B1(n7169), .B2(n7168), .A(n7167), .ZN(n7189) );
  INV_X1 U7838 ( .A(n7713), .ZN(n7179) );
  INV_X1 U7839 ( .A(n7170), .ZN(n7173) );
  NOR2_X1 U7840 ( .A1(n7715), .A2(n7562), .ZN(n7172) );
  AOI22_X1 U7841 ( .A1(n7218), .A2(n7173), .B1(n7172), .B2(n7171), .ZN(n7174)
         );
  OAI21_X1 U7842 ( .B1(n7189), .B2(n7179), .A(n7174), .ZN(n7175) );
  MUX2_X1 U7843 ( .A(n7175), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(n7704), 
        .Z(U3460) );
  INV_X1 U7844 ( .A(n7183), .ZN(n7180) );
  INV_X1 U7845 ( .A(n7176), .ZN(n7178) );
  OAI22_X1 U7846 ( .A1(n7180), .A2(n7179), .B1(n7178), .B2(n7177), .ZN(n7182)
         );
  MUX2_X1 U7847 ( .A(n7182), .B(n7181), .S(n7704), .Z(U3456) );
  AND2_X1 U7848 ( .A1(n7184), .A2(n7183), .ZN(n7199) );
  NAND2_X1 U7849 ( .A1(n7184), .A2(n7185), .ZN(n7196) );
  INV_X1 U7850 ( .A(n7186), .ZN(n7187) );
  OAI211_X1 U7851 ( .C1(n4279), .C2(n7188), .A(n7187), .B(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n7194) );
  INV_X1 U7852 ( .A(n7194), .ZN(n7191) );
  OAI22_X1 U7853 ( .A1(n7191), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n7190), .B2(n7189), .ZN(n7192) );
  OAI21_X1 U7854 ( .B1(n7194), .B2(n7193), .A(n7192), .ZN(n7195) );
  AOI222_X1 U7855 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n7196), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n7195), .C1(n7196), .C2(n7195), 
        .ZN(n7197) );
  AOI222_X1 U7856 ( .A1(n7199), .A2(n7198), .B1(n7199), .B2(n7197), .C1(n7198), 
        .C2(n7197), .ZN(n7209) );
  INV_X1 U7857 ( .A(n7200), .ZN(n7205) );
  AOI21_X1 U7858 ( .B1(n7702), .B2(n7202), .A(n7201), .ZN(n7204) );
  NOR4_X1 U7859 ( .A1(n7206), .A2(n7205), .A3(n7204), .A4(n7203), .ZN(n7207)
         );
  OAI211_X1 U7860 ( .C1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n7209), .A(n7208), .B(n7207), .ZN(n7224) );
  OAI22_X1 U7861 ( .A1(n7224), .A2(n7211), .B1(n7442), .B2(n7210), .ZN(n7216)
         );
  INV_X1 U7862 ( .A(n7212), .ZN(n7214) );
  NAND2_X1 U7863 ( .A1(n7214), .A2(n7213), .ZN(n7215) );
  NAND2_X1 U7864 ( .A1(n7216), .A2(n7215), .ZN(n7723) );
  INV_X1 U7865 ( .A(n7723), .ZN(n7217) );
  AOI211_X1 U7866 ( .C1(n7446), .C2(n7218), .A(STATE2_REG_0__SCAN_IN), .B(
        n7217), .ZN(n7219) );
  INV_X1 U7867 ( .A(n7219), .ZN(n7227) );
  INV_X1 U7868 ( .A(n7220), .ZN(n7223) );
  NOR2_X1 U7869 ( .A1(n7221), .A2(n7721), .ZN(n7222) );
  AOI211_X1 U7870 ( .C1(n7224), .C2(n7711), .A(n7223), .B(n7222), .ZN(n7226)
         );
  OAI21_X1 U7871 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n7442), .A(n7723), .ZN(
        n7225) );
  NAND2_X1 U7872 ( .A1(n7225), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7716) );
  NAND3_X1 U7873 ( .A1(n7227), .A2(n7226), .A3(n7716), .ZN(U3148) );
  INV_X2 U7874 ( .A(n7746), .ZN(n7734) );
  AND2_X1 U7875 ( .A1(STATE_REG_0__SCAN_IN), .A2(n7739), .ZN(n7254) );
  NOR2_X1 U7876 ( .A1(n7734), .A2(n7254), .ZN(n7230) );
  INV_X1 U7877 ( .A(n7230), .ZN(n7250) );
  NAND2_X1 U7878 ( .A1(n7737), .A2(n7736), .ZN(n7427) );
  AOI21_X1 U7879 ( .B1(n7228), .B2(n7427), .A(n7250), .ZN(n7725) );
  AOI21_X1 U7880 ( .B1(n7229), .B2(n7250), .A(n7725), .ZN(U3451) );
  NOR2_X1 U7881 ( .A1(n7729), .A2(n7231), .ZN(U3180) );
  NOR2_X1 U7882 ( .A1(n7729), .A2(n7232), .ZN(U3179) );
  NOR2_X1 U7883 ( .A1(n7729), .A2(n7233), .ZN(U3178) );
  NOR2_X1 U7884 ( .A1(n7729), .A2(n7234), .ZN(U3177) );
  NOR2_X1 U7885 ( .A1(n7729), .A2(n7235), .ZN(U3176) );
  NOR2_X1 U7886 ( .A1(n7729), .A2(n7236), .ZN(U3175) );
  INV_X1 U7887 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n7237) );
  NOR2_X1 U7888 ( .A1(n7729), .A2(n7237), .ZN(U3174) );
  NOR2_X1 U7889 ( .A1(n7729), .A2(n7238), .ZN(U3173) );
  NOR2_X1 U7890 ( .A1(n7729), .A2(n7239), .ZN(U3172) );
  INV_X1 U7891 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n7240) );
  NOR2_X1 U7892 ( .A1(n7729), .A2(n7240), .ZN(U3171) );
  INV_X1 U7893 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n7241) );
  NOR2_X1 U7894 ( .A1(n7729), .A2(n7241), .ZN(U3170) );
  NOR2_X1 U7895 ( .A1(n7729), .A2(n7242), .ZN(U3169) );
  NOR2_X1 U7896 ( .A1(n7729), .A2(n7243), .ZN(U3168) );
  NOR2_X1 U7897 ( .A1(n7729), .A2(n7244), .ZN(U3167) );
  NOR2_X1 U7898 ( .A1(n7729), .A2(n7245), .ZN(U3166) );
  NOR2_X1 U7899 ( .A1(n7729), .A2(n7246), .ZN(U3165) );
  AND2_X1 U7900 ( .A1(n7250), .A2(DATAWIDTH_REG_18__SCAN_IN), .ZN(U3164) );
  NOR2_X1 U7901 ( .A1(n7729), .A2(n7247), .ZN(U3163) );
  AND2_X1 U7902 ( .A1(n7250), .A2(DATAWIDTH_REG_20__SCAN_IN), .ZN(U3162) );
  NOR2_X1 U7903 ( .A1(n7729), .A2(n7248), .ZN(U3161) );
  NOR2_X1 U7904 ( .A1(n7729), .A2(n7249), .ZN(U3160) );
  AND2_X1 U7905 ( .A1(n7250), .A2(DATAWIDTH_REG_23__SCAN_IN), .ZN(U3159) );
  AND2_X1 U7906 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n7250), .ZN(U3158) );
  AND2_X1 U7907 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n7250), .ZN(U3157) );
  AND2_X1 U7908 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n7250), .ZN(U3156) );
  AND2_X1 U7909 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n7250), .ZN(U3155) );
  AND2_X1 U7910 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n7250), .ZN(U3154) );
  AND2_X1 U7911 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n7250), .ZN(U3153) );
  AND2_X1 U7912 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n7250), .ZN(U3152) );
  AND2_X1 U7913 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n7250), .ZN(U3151) );
  AND2_X1 U7914 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n7251), .ZN(U3019)
         );
  AND2_X1 U7915 ( .A1(n7252), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI21_X1 U7916 ( .B1(n7254), .B2(n7253), .A(n7734), .ZN(U2789) );
  AOI22_X1 U7917 ( .A1(n7284), .A2(LWORD_REG_0__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n7256) );
  OAI21_X1 U7918 ( .B1(n7257), .B2(n7286), .A(n7256), .ZN(U2923) );
  AOI22_X1 U7919 ( .A1(n7284), .A2(LWORD_REG_1__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n7258) );
  OAI21_X1 U7920 ( .B1(n7259), .B2(n7286), .A(n7258), .ZN(U2922) );
  AOI22_X1 U7921 ( .A1(n7284), .A2(LWORD_REG_2__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n7260) );
  OAI21_X1 U7922 ( .B1(n7261), .B2(n7286), .A(n7260), .ZN(U2921) );
  AOI22_X1 U7923 ( .A1(n7284), .A2(LWORD_REG_3__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n7262) );
  OAI21_X1 U7924 ( .B1(n7263), .B2(n7286), .A(n7262), .ZN(U2920) );
  AOI22_X1 U7925 ( .A1(n7284), .A2(LWORD_REG_4__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n7264) );
  OAI21_X1 U7926 ( .B1(n7265), .B2(n7286), .A(n7264), .ZN(U2919) );
  AOI22_X1 U7927 ( .A1(n7284), .A2(LWORD_REG_5__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n7266) );
  OAI21_X1 U7928 ( .B1(n7267), .B2(n7286), .A(n7266), .ZN(U2918) );
  AOI22_X1 U7929 ( .A1(n7284), .A2(LWORD_REG_6__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n7268) );
  OAI21_X1 U7930 ( .B1(n7269), .B2(n7286), .A(n7268), .ZN(U2917) );
  AOI22_X1 U7931 ( .A1(n7284), .A2(LWORD_REG_7__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n7270) );
  OAI21_X1 U7932 ( .B1(n4329), .B2(n7286), .A(n7270), .ZN(U2916) );
  AOI22_X1 U7933 ( .A1(n7284), .A2(LWORD_REG_8__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n7271) );
  OAI21_X1 U7934 ( .B1(n7272), .B2(n7286), .A(n7271), .ZN(U2915) );
  AOI22_X1 U7935 ( .A1(n7284), .A2(LWORD_REG_9__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n7273) );
  OAI21_X1 U7936 ( .B1(n7274), .B2(n7286), .A(n7273), .ZN(U2914) );
  AOI22_X1 U7937 ( .A1(n7284), .A2(LWORD_REG_10__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n7275) );
  OAI21_X1 U7938 ( .B1(n7276), .B2(n7286), .A(n7275), .ZN(U2913) );
  AOI22_X1 U7939 ( .A1(n7284), .A2(LWORD_REG_11__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n7277) );
  OAI21_X1 U7940 ( .B1(n7278), .B2(n7286), .A(n7277), .ZN(U2912) );
  AOI22_X1 U7941 ( .A1(n7284), .A2(LWORD_REG_12__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n7279) );
  OAI21_X1 U7942 ( .B1(n4396), .B2(n7286), .A(n7279), .ZN(U2911) );
  AOI22_X1 U7943 ( .A1(n7284), .A2(LWORD_REG_13__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n7280) );
  OAI21_X1 U7944 ( .B1(n7281), .B2(n7286), .A(n7280), .ZN(U2910) );
  AOI22_X1 U7945 ( .A1(n7284), .A2(LWORD_REG_14__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n7282) );
  OAI21_X1 U7946 ( .B1(n7283), .B2(n7286), .A(n7282), .ZN(U2909) );
  AOI22_X1 U7947 ( .A1(n7284), .A2(LWORD_REG_15__SCAN_IN), .B1(n7252), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n7285) );
  OAI21_X1 U7948 ( .B1(n7287), .B2(n7286), .A(n7285), .ZN(U2908) );
  OAI222_X1 U7949 ( .A1(n7320), .A2(n6870), .B1(n7288), .B2(n7734), .C1(n7353), 
        .C2(n7338), .ZN(U3184) );
  OAI222_X1 U7950 ( .A1(n7320), .A2(n7290), .B1(n7289), .B2(n7734), .C1(n6870), 
        .C2(n7338), .ZN(U3185) );
  OAI222_X1 U7951 ( .A1(n7320), .A2(n7292), .B1(n7291), .B2(n7734), .C1(n7290), 
        .C2(n7338), .ZN(U3186) );
  INV_X1 U7952 ( .A(REIP_REG_5__SCAN_IN), .ZN(n7295) );
  OAI222_X1 U7953 ( .A1(n7320), .A2(n7295), .B1(n7293), .B2(n7734), .C1(n7292), 
        .C2(n7338), .ZN(U3187) );
  INV_X1 U7954 ( .A(REIP_REG_6__SCAN_IN), .ZN(n7296) );
  OAI222_X1 U7955 ( .A1(n7338), .A2(n7295), .B1(n7294), .B2(n7734), .C1(n7296), 
        .C2(n7320), .ZN(U3188) );
  OAI222_X1 U7956 ( .A1(n7320), .A2(n6055), .B1(n7297), .B2(n7734), .C1(n7296), 
        .C2(n7338), .ZN(U3189) );
  OAI222_X1 U7957 ( .A1(n7320), .A2(n6225), .B1(n7298), .B2(n7734), .C1(n6055), 
        .C2(n7338), .ZN(U3190) );
  OAI222_X1 U7958 ( .A1(n7320), .A2(n7619), .B1(n7299), .B2(n7734), .C1(n6225), 
        .C2(n7338), .ZN(U3191) );
  INV_X1 U7959 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n7300) );
  OAI222_X1 U7960 ( .A1(n7338), .A2(n7619), .B1(n7300), .B2(n7734), .C1(n7631), 
        .C2(n7320), .ZN(U3192) );
  OAI222_X1 U7961 ( .A1(n7338), .A2(n7631), .B1(n7301), .B2(n7734), .C1(n7640), 
        .C2(n7320), .ZN(U3193) );
  INV_X1 U7962 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n7302) );
  OAI222_X1 U7963 ( .A1(n7320), .A2(n6509), .B1(n7302), .B2(n7734), .C1(n7640), 
        .C2(n7338), .ZN(U3194) );
  INV_X1 U7964 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n7303) );
  INV_X1 U7965 ( .A(REIP_REG_13__SCAN_IN), .ZN(n7645) );
  OAI222_X1 U7966 ( .A1(n7338), .A2(n6509), .B1(n7303), .B2(n7734), .C1(n7645), 
        .C2(n7320), .ZN(U3195) );
  INV_X1 U7967 ( .A(REIP_REG_14__SCAN_IN), .ZN(n7305) );
  INV_X1 U7968 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n7304) );
  OAI222_X1 U7969 ( .A1(n7320), .A2(n7305), .B1(n7304), .B2(n7734), .C1(n7645), 
        .C2(n7338), .ZN(U3196) );
  OAI222_X1 U7970 ( .A1(n7320), .A2(n7308), .B1(n7306), .B2(n7734), .C1(n7305), 
        .C2(n7338), .ZN(U3197) );
  OAI222_X1 U7971 ( .A1(n7338), .A2(n7308), .B1(n7307), .B2(n7734), .C1(n7525), 
        .C2(n7320), .ZN(U3198) );
  OAI222_X1 U7972 ( .A1(n7320), .A2(n7311), .B1(n7309), .B2(n7734), .C1(n7525), 
        .C2(n7338), .ZN(U3199) );
  OAI222_X1 U7973 ( .A1(n7338), .A2(n7311), .B1(n7310), .B2(n7734), .C1(n7671), 
        .C2(n7320), .ZN(U3200) );
  OAI222_X1 U7974 ( .A1(n7320), .A2(n7673), .B1(n7312), .B2(n7734), .C1(n7671), 
        .C2(n7338), .ZN(U3201) );
  OAI222_X1 U7975 ( .A1(n7338), .A2(n7673), .B1(n7313), .B2(n7734), .C1(n7315), 
        .C2(n7320), .ZN(U3202) );
  OAI222_X1 U7976 ( .A1(n7338), .A2(n7315), .B1(n7314), .B2(n7734), .C1(n7317), 
        .C2(n7320), .ZN(U3203) );
  OAI222_X1 U7977 ( .A1(n7338), .A2(n7317), .B1(n7316), .B2(n7734), .C1(n7318), 
        .C2(n7320), .ZN(U3204) );
  OAI222_X1 U7978 ( .A1(n7320), .A2(n7322), .B1(n7319), .B2(n7734), .C1(n7318), 
        .C2(n7338), .ZN(U3205) );
  INV_X1 U7979 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n7321) );
  OAI222_X1 U7980 ( .A1(n7338), .A2(n7322), .B1(n7321), .B2(n7734), .C1(n7323), 
        .C2(n7320), .ZN(U3206) );
  OAI222_X1 U7981 ( .A1(n7320), .A2(n7326), .B1(n7324), .B2(n7734), .C1(n7323), 
        .C2(n7338), .ZN(U3207) );
  INV_X1 U7982 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n7325) );
  OAI222_X1 U7983 ( .A1(n7338), .A2(n7326), .B1(n7325), .B2(n7734), .C1(n7328), 
        .C2(n7320), .ZN(U3208) );
  OAI222_X1 U7984 ( .A1(n7338), .A2(n7328), .B1(n7327), .B2(n7734), .C1(n7330), 
        .C2(n7320), .ZN(U3209) );
  OAI222_X1 U7985 ( .A1(n7338), .A2(n7330), .B1(n7329), .B2(n7734), .C1(n7332), 
        .C2(n7320), .ZN(U3210) );
  OAI222_X1 U7986 ( .A1(n7338), .A2(n7332), .B1(n7331), .B2(n7734), .C1(n7333), 
        .C2(n7320), .ZN(U3211) );
  OAI222_X1 U7987 ( .A1(n7320), .A2(n7337), .B1(n7334), .B2(n7734), .C1(n7333), 
        .C2(n7338), .ZN(U3212) );
  OAI222_X1 U7988 ( .A1(n7338), .A2(n7337), .B1(n7336), .B2(n7734), .C1(n7335), 
        .C2(n7320), .ZN(U3213) );
  AOI22_X1 U7989 ( .A1(n7734), .A2(n7340), .B1(n7339), .B2(n7746), .ZN(U3445)
         );
  AOI221_X1 U7990 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(REIP_REG_1__SCAN_IN), 
        .C1(REIP_REG_0__SCAN_IN), .C2(REIP_REG_1__SCAN_IN), .A(
        DATAWIDTH_REG_1__SCAN_IN), .ZN(n7351) );
  NOR4_X1 U7991 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(
        DATAWIDTH_REG_31__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_29__SCAN_IN), .ZN(n7344) );
  NOR4_X1 U7992 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n7343) );
  NOR4_X1 U7993 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_24__SCAN_IN), .ZN(n7342) );
  NOR4_X1 U7994 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_27__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_25__SCAN_IN), .ZN(n7341) );
  NAND4_X1 U7995 ( .A1(n7344), .A2(n7343), .A3(n7342), .A4(n7341), .ZN(n7350)
         );
  NOR4_X1 U7996 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_10__SCAN_IN), .ZN(n7348) );
  AOI211_X1 U7997 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_21__SCAN_IN), .B(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n7347) );
  NOR4_X1 U7998 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), .A3(DATAWIDTH_REG_2__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(n7346) );
  NOR4_X1 U7999 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_9__SCAN_IN), .ZN(n7345) );
  NAND4_X1 U8000 ( .A1(n7348), .A2(n7347), .A3(n7346), .A4(n7345), .ZN(n7349)
         );
  NOR2_X1 U8001 ( .A1(n7350), .A2(n7349), .ZN(n7364) );
  MUX2_X1 U8002 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(n7351), .S(n7364), .Z(
        U2795) );
  OAI22_X1 U8003 ( .A1(n7746), .A2(BYTEENABLE_REG_2__SCAN_IN), .B1(
        BE_N_REG_2__SCAN_IN), .B2(n7734), .ZN(n7352) );
  INV_X1 U8004 ( .A(n7352), .ZN(U3446) );
  AOI21_X1 U8005 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n7354) );
  OAI221_X1 U8006 ( .B1(REIP_REG_1__SCAN_IN), .B2(n7354), .C1(n7353), .C2(
        REIP_REG_0__SCAN_IN), .A(n7364), .ZN(n7355) );
  OAI21_X1 U8007 ( .B1(n7364), .B2(n7356), .A(n7355), .ZN(U3468) );
  INV_X1 U8008 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n7360) );
  AOI22_X1 U8009 ( .A1(n7734), .A2(n7360), .B1(n7357), .B2(n7746), .ZN(U3447)
         );
  NOR3_X1 U8010 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(REIP_REG_0__SCAN_IN), .ZN(n7358) );
  OAI21_X1 U8011 ( .B1(REIP_REG_1__SCAN_IN), .B2(n7358), .A(n7364), .ZN(n7359)
         );
  OAI21_X1 U8012 ( .B1(n7364), .B2(n7360), .A(n7359), .ZN(U2794) );
  AOI22_X1 U8013 ( .A1(n7734), .A2(n7363), .B1(n7361), .B2(n7746), .ZN(U3448)
         );
  OAI21_X1 U8014 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n7364), .ZN(n7362) );
  OAI21_X1 U8015 ( .B1(n7364), .B2(n7363), .A(n7362), .ZN(U3469) );
  NOR2_X1 U8016 ( .A1(n7694), .A2(n6917), .ZN(n7365) );
  AOI21_X1 U8017 ( .B1(n7761), .B2(n7366), .A(n7365), .ZN(n7367) );
  OAI21_X1 U8018 ( .B1(n7369), .B2(n7368), .A(n7367), .ZN(U2839) );
  AOI22_X1 U8019 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n7415), .B1(n7544), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n7374) );
  INV_X1 U8020 ( .A(n7370), .ZN(n7372) );
  AOI22_X1 U8021 ( .A1(n7372), .A2(n7421), .B1(n7371), .B2(n7422), .ZN(n7373)
         );
  OAI211_X1 U8022 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n7425), .A(n7374), 
        .B(n7373), .ZN(U2985) );
  AOI22_X1 U8023 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n7415), .B1(n7544), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n7380) );
  XNOR2_X1 U8024 ( .A(n7375), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n7377)
         );
  XNOR2_X1 U8025 ( .A(n7377), .B(n7376), .ZN(n7471) );
  AOI22_X1 U8026 ( .A1(n7378), .A2(n7421), .B1(n7471), .B2(n7422), .ZN(n7379)
         );
  OAI211_X1 U8027 ( .C1(n7425), .C2(n7381), .A(n7380), .B(n7379), .ZN(U2984)
         );
  AOI22_X1 U8028 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n7415), .B1(n7544), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n7388) );
  NAND2_X1 U8029 ( .A1(n7382), .A2(n7383), .ZN(n7384) );
  AND2_X1 U8030 ( .A1(n7385), .A2(n7384), .ZN(n7451) );
  AOI22_X1 U8031 ( .A1(n7422), .A2(n7451), .B1(n7386), .B2(n7421), .ZN(n7387)
         );
  OAI211_X1 U8032 ( .C1(n7425), .C2(n7389), .A(n7388), .B(n7387), .ZN(U2982)
         );
  AOI22_X1 U8033 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n7415), .B1(n7544), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n7393) );
  INV_X1 U8034 ( .A(n7390), .ZN(n7391) );
  AOI22_X1 U8035 ( .A1(n7391), .A2(n7422), .B1(n7421), .B2(n7570), .ZN(n7392)
         );
  OAI211_X1 U8036 ( .C1(n7425), .C2(n7567), .A(n7393), .B(n7392), .ZN(U2981)
         );
  AOI22_X1 U8037 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n7415), .B1(n7544), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n7398) );
  XNOR2_X1 U8038 ( .A(n7395), .B(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n7396)
         );
  XNOR2_X1 U8039 ( .A(n7394), .B(n7396), .ZN(n7463) );
  AOI22_X1 U8040 ( .A1(n7421), .A2(n7580), .B1(n7463), .B2(n7422), .ZN(n7397)
         );
  OAI211_X1 U8041 ( .C1(n7425), .C2(n7584), .A(n7398), .B(n7397), .ZN(U2980)
         );
  INV_X1 U8042 ( .A(n7399), .ZN(n7401) );
  INV_X1 U8043 ( .A(n7596), .ZN(n7400) );
  AOI222_X1 U8044 ( .A1(n7401), .A2(n7422), .B1(n7400), .B2(n7409), .C1(n7421), 
        .C2(n7592), .ZN(n7403) );
  OAI211_X1 U8045 ( .C1(n7405), .C2(n7404), .A(n7403), .B(n7402), .ZN(U2979)
         );
  OAI21_X1 U8046 ( .B1(n7408), .B2(n7407), .A(n7406), .ZN(n7505) );
  AOI22_X1 U8047 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n7415), .B1(n7544), 
        .B2(REIP_REG_11__SCAN_IN), .ZN(n7411) );
  AOI22_X1 U8048 ( .A1(n7639), .A2(n7421), .B1(n7409), .B2(n7638), .ZN(n7410)
         );
  OAI211_X1 U8049 ( .C1(n7701), .C2(n7505), .A(n7411), .B(n7410), .ZN(U2975)
         );
  AOI22_X1 U8050 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n7415), .B1(n7544), 
        .B2(REIP_REG_13__SCAN_IN), .ZN(n7414) );
  AOI22_X1 U8051 ( .A1(n7412), .A2(n7422), .B1(n7421), .B2(n7656), .ZN(n7413)
         );
  OAI211_X1 U8052 ( .C1(n7425), .C2(n7661), .A(n7414), .B(n7413), .ZN(U2973)
         );
  AOI22_X1 U8053 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n7415), .B1(n7544), 
        .B2(REIP_REG_18__SCAN_IN), .ZN(n7424) );
  NAND2_X1 U8054 ( .A1(n3631), .A2(n7539), .ZN(n7417) );
  NAND2_X1 U8055 ( .A1(n4252), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n7416) );
  OAI22_X1 U8056 ( .A1(n7418), .A2(n7417), .B1(n7024), .B2(n7416), .ZN(n7419)
         );
  XOR2_X1 U8057 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .B(n7419), .Z(n7546) );
  AOI22_X1 U8058 ( .A1(n7546), .A2(n7422), .B1(n7421), .B2(n7756), .ZN(n7423)
         );
  OAI211_X1 U8059 ( .C1(n7425), .C2(n7669), .A(n7424), .B(n7423), .ZN(U2968)
         );
  NOR2_X1 U8060 ( .A1(n7734), .A2(D_C_N_REG_SCAN_IN), .ZN(n7426) );
  AOI22_X1 U8061 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n7734), .B1(n7427), .B2(
        n7426), .ZN(U2791) );
  INV_X1 U8062 ( .A(n7431), .ZN(n7440) );
  OAI221_X1 U8063 ( .B1(n7431), .B2(n7430), .C1(n7429), .C2(n7440), .A(n7428), 
        .ZN(U3474) );
  AOI22_X1 U8064 ( .A1(n7734), .A2(READREQUEST_REG_SCAN_IN), .B1(n7432), .B2(
        n7746), .ZN(U3470) );
  NOR2_X1 U8065 ( .A1(n7737), .A2(n7735), .ZN(n7731) );
  AOI22_X1 U8066 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        STATE_REG_0__SCAN_IN), .B2(REQUESTPENDING_REG_SCAN_IN), .ZN(n7436) );
  NOR2_X1 U8067 ( .A1(n7433), .A2(n7442), .ZN(n7741) );
  INV_X1 U8068 ( .A(n7741), .ZN(n7434) );
  OAI211_X1 U8069 ( .C1(n7731), .C2(n7436), .A(n7435), .B(n7434), .ZN(U3182)
         );
  NOR2_X1 U8070 ( .A1(n7437), .A2(READY_N), .ZN(n7712) );
  OAI21_X1 U8071 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n7712), .A(n7721), .ZN(
        n7439) );
  OAI21_X1 U8072 ( .B1(n7446), .B2(n7439), .A(n7438), .ZN(U3150) );
  INV_X1 U8073 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7730) );
  AOI211_X1 U8074 ( .C1(n7284), .C2(n7442), .A(n7441), .B(n7440), .ZN(n7449)
         );
  OAI21_X1 U8075 ( .B1(n7443), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n7444) );
  OAI21_X1 U8076 ( .B1(n7445), .B2(n7444), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n7448) );
  NOR2_X1 U8077 ( .A1(n7449), .A2(n7446), .ZN(n7447) );
  AOI22_X1 U8078 ( .A1(n7730), .A2(n7449), .B1(n7448), .B2(n7447), .ZN(U3472)
         );
  OAI211_X1 U8079 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n7461), .B(n7473), .ZN(n7455) );
  AOI22_X1 U8080 ( .A1(n7545), .A2(n7450), .B1(n7544), .B2(REIP_REG_4__SCAN_IN), .ZN(n7454) );
  AOI22_X1 U8081 ( .A1(n7452), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .B1(n7451), 
        .B2(n7557), .ZN(n7453) );
  OAI211_X1 U8082 ( .C1(n7456), .C2(n7455), .A(n7454), .B(n7453), .ZN(U3014)
         );
  INV_X1 U8083 ( .A(n7457), .ZN(n7467) );
  INV_X1 U8084 ( .A(n7575), .ZN(n7458) );
  AOI22_X1 U8085 ( .A1(n7458), .A2(n7545), .B1(n7544), .B2(REIP_REG_6__SCAN_IN), .ZN(n7465) );
  NOR3_X1 U8086 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n7460), .A3(n7459), 
        .ZN(n7462) );
  AOI22_X1 U8087 ( .A1(n7463), .A2(n7557), .B1(n7462), .B2(n7461), .ZN(n7464)
         );
  OAI211_X1 U8088 ( .C1(n7467), .C2(n7466), .A(n7465), .B(n7464), .ZN(U3012)
         );
  AOI22_X1 U8089 ( .A1(n7545), .A2(n7468), .B1(n7544), .B2(REIP_REG_2__SCAN_IN), .ZN(n7479) );
  NAND2_X1 U8090 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n7470) );
  OAI21_X1 U8091 ( .B1(n7530), .B2(n7470), .A(n7469), .ZN(n7472) );
  AOI22_X1 U8092 ( .A1(n7472), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n7557), 
        .B2(n7471), .ZN(n7478) );
  OR2_X1 U8093 ( .A1(n7530), .A2(n7473), .ZN(n7477) );
  INV_X1 U8094 ( .A(n7474), .ZN(n7540) );
  NAND3_X1 U8095 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n7540), .A3(n7475), 
        .ZN(n7476) );
  NAND4_X1 U8096 ( .A1(n7479), .A2(n7478), .A3(n7477), .A4(n7476), .ZN(U3016)
         );
  AOI21_X1 U8097 ( .B1(n7621), .B2(n7545), .A(n7480), .ZN(n7487) );
  AOI21_X1 U8098 ( .B1(n7489), .B2(n7482), .A(n7481), .ZN(n7484) );
  AOI22_X1 U8099 ( .A1(n7485), .A2(n7557), .B1(n7484), .B2(n7483), .ZN(n7486)
         );
  OAI211_X1 U8100 ( .C1(n7489), .C2(n7488), .A(n7487), .B(n7486), .ZN(U3008)
         );
  INV_X1 U8101 ( .A(n7490), .ZN(n7491) );
  AOI221_X1 U8102 ( .B1(n7492), .B2(n7503), .C1(n7491), .C2(n7503), .A(n7507), 
        .ZN(n7500) );
  INV_X1 U8103 ( .A(n7493), .ZN(n7495) );
  AOI21_X1 U8104 ( .B1(n7495), .B2(n7545), .A(n7494), .ZN(n7499) );
  NOR3_X1 U8105 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n7542), .A3(n7503), 
        .ZN(n7496) );
  AOI21_X1 U8106 ( .B1(n7557), .B2(n7497), .A(n7496), .ZN(n7498) );
  OAI211_X1 U8107 ( .C1(n7500), .C2(n6506), .A(n7499), .B(n7498), .ZN(U3006)
         );
  INV_X1 U8108 ( .A(n7542), .ZN(n7502) );
  OAI22_X1 U8109 ( .A1(n7634), .A2(n7555), .B1(n7640), .B2(n7524), .ZN(n7501)
         );
  AOI221_X1 U8110 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n7507), .C1(
        n7503), .C2(n7502), .A(n7501), .ZN(n7504) );
  OAI21_X1 U8111 ( .B1(n7506), .B2(n7505), .A(n7504), .ZN(U3007) );
  AOI21_X1 U8112 ( .B1(n7509), .B2(n7508), .A(n7507), .ZN(n7517) );
  AOI22_X1 U8113 ( .A1(REIP_REG_15__SCAN_IN), .A2(n7544), .B1(n7521), .B2(
        n7514), .ZN(n7513) );
  AOI22_X1 U8114 ( .A1(n7511), .A2(n7557), .B1(n7545), .B2(n7510), .ZN(n7512)
         );
  OAI211_X1 U8115 ( .C1(n7517), .C2(n7514), .A(n7513), .B(n7512), .ZN(U3003)
         );
  OAI22_X1 U8116 ( .A1(n7517), .A2(n7516), .B1(n7555), .B2(n7515), .ZN(n7518)
         );
  AOI21_X1 U8117 ( .B1(n7519), .B2(n7557), .A(n7518), .ZN(n7523) );
  OAI211_X1 U8118 ( .C1(INSTADDRPOINTER_REG_16__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A(n7521), .B(n7520), .ZN(n7522) );
  OAI211_X1 U8119 ( .C1(n7525), .C2(n7524), .A(n7523), .B(n7522), .ZN(U3002)
         );
  AOI21_X1 U8120 ( .B1(n7528), .B2(n7527), .A(n7526), .ZN(n7529) );
  OAI21_X1 U8121 ( .B1(n7531), .B2(n7530), .A(n7529), .ZN(n7538) );
  AOI22_X1 U8122 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n7538), .B1(n7544), .B2(REIP_REG_17__SCAN_IN), .ZN(n7536) );
  INV_X1 U8123 ( .A(n7532), .ZN(n7534) );
  AOI22_X1 U8124 ( .A1(n7534), .A2(n7557), .B1(n7545), .B2(n7533), .ZN(n7535)
         );
  OAI211_X1 U8125 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n7537), .A(n7536), .B(n7535), .ZN(U3001) );
  AOI21_X1 U8126 ( .B1(n7540), .B2(n7539), .A(n7538), .ZN(n7550) );
  INV_X1 U8127 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n7549) );
  NOR3_X1 U8128 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n7542), .A3(n7541), 
        .ZN(n7543) );
  AOI21_X1 U8129 ( .B1(REIP_REG_18__SCAN_IN), .B2(n7544), .A(n7543), .ZN(n7548) );
  AOI22_X1 U8130 ( .A1(n7546), .A2(n7557), .B1(n7545), .B2(n7665), .ZN(n7547)
         );
  OAI211_X1 U8131 ( .C1(n7550), .C2(n7549), .A(n7548), .B(n7547), .ZN(U3000)
         );
  INV_X1 U8132 ( .A(n7551), .ZN(n7558) );
  OAI211_X1 U8133 ( .C1(n7555), .C2(n7554), .A(n7553), .B(n7552), .ZN(n7556)
         );
  AOI21_X1 U8134 ( .B1(n7558), .B2(n7557), .A(n7556), .ZN(n7559) );
  OAI221_X1 U8135 ( .B1(n7562), .B2(n7561), .C1(n7562), .C2(n7560), .A(n7559), 
        .ZN(U3018) );
  NOR2_X1 U8136 ( .A1(n7563), .A2(REIP_REG_5__SCAN_IN), .ZN(n7573) );
  OAI22_X1 U8137 ( .A1(n7565), .A2(n7686), .B1(n7693), .B2(n7564), .ZN(n7566)
         );
  AOI211_X1 U8138 ( .C1(n7688), .C2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n7677), 
        .B(n7566), .ZN(n7572) );
  INV_X1 U8139 ( .A(n7567), .ZN(n7568) );
  AOI22_X1 U8140 ( .A1(n7570), .A2(n7569), .B1(n7568), .B2(n7682), .ZN(n7571)
         );
  OAI211_X1 U8141 ( .C1(n7573), .C2(n7574), .A(n7572), .B(n7571), .ZN(U2822)
         );
  INV_X1 U8142 ( .A(n7574), .ZN(n7597) );
  NOR2_X1 U8143 ( .A1(REIP_REG_6__SCAN_IN), .A2(n7618), .ZN(n7593) );
  NOR2_X1 U8144 ( .A1(n7693), .A2(n7575), .ZN(n7579) );
  NAND2_X1 U8145 ( .A1(n7688), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n7576)
         );
  OAI211_X1 U8146 ( .C1(n7686), .C2(n7577), .A(n7648), .B(n7576), .ZN(n7578)
         );
  AOI211_X1 U8147 ( .C1(n7580), .C2(n7696), .A(n7579), .B(n7578), .ZN(n7581)
         );
  INV_X1 U8148 ( .A(n7581), .ZN(n7582) );
  AOI211_X1 U8149 ( .C1(n7597), .C2(REIP_REG_6__SCAN_IN), .A(n7593), .B(n7582), 
        .ZN(n7583) );
  OAI21_X1 U8150 ( .B1(n7584), .B2(n7699), .A(n7583), .ZN(U2821) );
  INV_X1 U8151 ( .A(n7585), .ZN(n7590) );
  NAND3_X1 U8152 ( .A1(REIP_REG_6__SCAN_IN), .A2(n7599), .A3(n6055), .ZN(n7589) );
  NOR2_X1 U8153 ( .A1(n7686), .A2(n7586), .ZN(n7587) );
  AOI211_X1 U8154 ( .C1(n7688), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n7677), 
        .B(n7587), .ZN(n7588) );
  OAI211_X1 U8155 ( .C1(n7693), .C2(n7590), .A(n7589), .B(n7588), .ZN(n7591)
         );
  AOI21_X1 U8156 ( .B1(n7696), .B2(n7592), .A(n7591), .ZN(n7595) );
  OAI21_X1 U8157 ( .B1(n7597), .B2(n7593), .A(REIP_REG_7__SCAN_IN), .ZN(n7594)
         );
  OAI211_X1 U8158 ( .C1(n7699), .C2(n7596), .A(n7595), .B(n7594), .ZN(U2820)
         );
  AOI21_X1 U8159 ( .B1(n7620), .B2(n7598), .A(n7597), .ZN(n7630) );
  NAND3_X1 U8160 ( .A1(REIP_REG_6__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        n7599), .ZN(n7602) );
  AOI22_X1 U8161 ( .A1(EBX_REG_8__SCAN_IN), .A2(n7687), .B1(n7666), .B2(n7600), 
        .ZN(n7601) );
  OAI21_X1 U8162 ( .B1(REIP_REG_8__SCAN_IN), .B2(n7602), .A(n7601), .ZN(n7603)
         );
  AOI211_X1 U8163 ( .C1(n7688), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n7677), 
        .B(n7603), .ZN(n7608) );
  OAI22_X1 U8164 ( .A1(n7605), .A2(n7679), .B1(n7604), .B2(n7699), .ZN(n7606)
         );
  INV_X1 U8165 ( .A(n7606), .ZN(n7607) );
  OAI211_X1 U8166 ( .C1(n7630), .C2(n6225), .A(n7608), .B(n7607), .ZN(U2819)
         );
  NOR2_X1 U8167 ( .A1(n7620), .A2(n7618), .ZN(n7609) );
  NAND2_X1 U8168 ( .A1(n7609), .A2(n7619), .ZN(n7629) );
  OAI22_X1 U8169 ( .A1(n7611), .A2(n7686), .B1(n7693), .B2(n7610), .ZN(n7612)
         );
  AOI211_X1 U8170 ( .C1(n7688), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n7677), 
        .B(n7612), .ZN(n7613) );
  OAI211_X1 U8171 ( .C1(n7614), .C2(n7679), .A(n7629), .B(n7613), .ZN(n7615)
         );
  AOI21_X1 U8172 ( .B1(n7616), .B2(n7682), .A(n7615), .ZN(n7617) );
  OAI21_X1 U8173 ( .B1(n7630), .B2(n7619), .A(n7617), .ZN(U2818) );
  NOR3_X1 U8174 ( .A1(n7620), .A2(n7619), .A3(n7618), .ZN(n7641) );
  AOI22_X1 U8175 ( .A1(n7666), .A2(n7621), .B1(n7641), .B2(n7631), .ZN(n7622)
         );
  OAI211_X1 U8176 ( .C1(n7633), .C2(n7623), .A(n7622), .B(n7648), .ZN(n7627)
         );
  OAI22_X1 U8177 ( .A1(n7625), .A2(n7679), .B1(n7624), .B2(n7699), .ZN(n7626)
         );
  AOI211_X1 U8178 ( .C1(EBX_REG_10__SCAN_IN), .C2(n7687), .A(n7627), .B(n7626), 
        .ZN(n7628) );
  OAI221_X1 U8179 ( .B1(n7631), .B2(n7630), .C1(n7631), .C2(n7629), .A(n7628), 
        .ZN(U2817) );
  OAI21_X1 U8180 ( .B1(n7633), .B2(n7632), .A(n7648), .ZN(n7637) );
  OAI22_X1 U8181 ( .A1(n7635), .A2(n7686), .B1(n7693), .B2(n7634), .ZN(n7636)
         );
  AOI211_X1 U8182 ( .C1(REIP_REG_11__SCAN_IN), .C2(n7657), .A(n7637), .B(n7636), .ZN(n7644) );
  AOI22_X1 U8183 ( .A1(n7639), .A2(n7696), .B1(n7682), .B2(n7638), .ZN(n7643)
         );
  NAND3_X1 U8184 ( .A1(REIP_REG_10__SCAN_IN), .A2(n7641), .A3(n7640), .ZN(
        n7642) );
  NAND3_X1 U8185 ( .A1(n7644), .A2(n7643), .A3(n7642), .ZN(U2816) );
  NAND3_X1 U8186 ( .A1(REIP_REG_12__SCAN_IN), .A2(n7646), .A3(n7645), .ZN(
        n7654) );
  INV_X1 U8187 ( .A(n7647), .ZN(n7652) );
  NAND2_X1 U8188 ( .A1(n7688), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n7649)
         );
  OAI211_X1 U8189 ( .C1(n7686), .C2(n7650), .A(n7649), .B(n7648), .ZN(n7651)
         );
  AOI21_X1 U8190 ( .B1(n7652), .B2(n7666), .A(n7651), .ZN(n7653) );
  NAND2_X1 U8191 ( .A1(n7654), .A2(n7653), .ZN(n7655) );
  AOI21_X1 U8192 ( .B1(n7656), .B2(n7696), .A(n7655), .ZN(n7660) );
  OAI21_X1 U8193 ( .B1(n7658), .B2(n7657), .A(REIP_REG_13__SCAN_IN), .ZN(n7659) );
  OAI211_X1 U8194 ( .C1(n7699), .C2(n7661), .A(n7660), .B(n7659), .ZN(U2814)
         );
  AOI22_X1 U8195 ( .A1(EBX_REG_18__SCAN_IN), .A2(n7687), .B1(
        REIP_REG_18__SCAN_IN), .B2(n7670), .ZN(n7663) );
  NAND2_X1 U8196 ( .A1(n7672), .A2(n7671), .ZN(n7662) );
  NAND2_X1 U8197 ( .A1(n7663), .A2(n7662), .ZN(n7664) );
  AOI211_X1 U8198 ( .C1(n7688), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n7677), 
        .B(n7664), .ZN(n7668) );
  AOI22_X1 U8199 ( .A1(n7756), .A2(n7696), .B1(n7666), .B2(n7665), .ZN(n7667)
         );
  OAI211_X1 U8200 ( .C1(n7669), .C2(n7699), .A(n7668), .B(n7667), .ZN(U2809)
         );
  AOI21_X1 U8201 ( .B1(n7672), .B2(n7671), .A(n7670), .ZN(n7675) );
  AOI22_X1 U8202 ( .A1(REIP_REG_19__SCAN_IN), .A2(n7675), .B1(n7674), .B2(
        n7673), .ZN(n7676) );
  AOI211_X1 U8203 ( .C1(n7688), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n7677), 
        .B(n7676), .ZN(n7685) );
  OAI22_X1 U8204 ( .A1(n7680), .A2(n7679), .B1(n7693), .B2(n7678), .ZN(n7681)
         );
  AOI21_X1 U8205 ( .B1(n7683), .B2(n7682), .A(n7681), .ZN(n7684) );
  OAI211_X1 U8206 ( .C1(n5187), .C2(n7686), .A(n7685), .B(n7684), .ZN(U2808)
         );
  AOI22_X1 U8207 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n7688), .B1(
        EBX_REG_20__SCAN_IN), .B2(n7687), .ZN(n7689) );
  INV_X1 U8208 ( .A(n7689), .ZN(n7690) );
  AOI221_X1 U8209 ( .B1(REIP_REG_20__SCAN_IN), .B2(n7692), .C1(n7691), .C2(
        n7692), .A(n7690), .ZN(n7698) );
  NOR2_X1 U8210 ( .A1(n7694), .A2(n7693), .ZN(n7695) );
  AOI21_X1 U8211 ( .B1(n7761), .B2(n7696), .A(n7695), .ZN(n7697) );
  OAI211_X1 U8212 ( .C1(n7700), .C2(n7699), .A(n7698), .B(n7697), .ZN(U2807)
         );
  OAI21_X1 U8213 ( .B1(n7703), .B2(n7702), .A(n7701), .ZN(U2793) );
  INV_X1 U8214 ( .A(n7704), .ZN(n7710) );
  INV_X1 U8215 ( .A(n7705), .ZN(n7707) );
  NAND3_X1 U8216 ( .A1(n7707), .A2(n7724), .A3(n7706), .ZN(n7708) );
  OAI21_X1 U8217 ( .B1(n7710), .B2(n7709), .A(n7708), .ZN(U3455) );
  AOI21_X1 U8218 ( .B1(n7713), .B2(n7712), .A(n7711), .ZN(n7714) );
  INV_X1 U8219 ( .A(n7714), .ZN(n7718) );
  AOI21_X1 U8220 ( .B1(n7716), .B2(n7723), .A(n7715), .ZN(n7717) );
  AOI21_X1 U8221 ( .B1(n7723), .B2(n7718), .A(n7717), .ZN(n7720) );
  NAND2_X1 U8222 ( .A1(n7720), .A2(n7719), .ZN(U3149) );
  OAI211_X1 U8223 ( .C1(n7724), .C2(n7723), .A(n7722), .B(n7721), .ZN(U3453)
         );
  INV_X1 U8224 ( .A(n7725), .ZN(n7727) );
  OAI21_X1 U8225 ( .B1(n7729), .B2(n7726), .A(n7727), .ZN(U2792) );
  OAI21_X1 U8226 ( .B1(n7729), .B2(n7728), .A(n7727), .ZN(U3452) );
  AOI211_X1 U8227 ( .C1(STATE_REG_1__SCAN_IN), .C2(HOLD), .A(n7731), .B(n7730), 
        .ZN(n7733) );
  NOR2_X1 U8228 ( .A1(n7741), .A2(n7736), .ZN(n7745) );
  INV_X1 U8229 ( .A(NA_N), .ZN(n7740) );
  OAI21_X1 U8230 ( .B1(n7740), .B2(STATE_REG_1__SCAN_IN), .A(
        STATE_REG_2__SCAN_IN), .ZN(n7744) );
  INV_X1 U8231 ( .A(n7744), .ZN(n7732) );
  OAI22_X1 U8232 ( .A1(n7734), .A2(n7733), .B1(n7745), .B2(n7732), .ZN(U3181)
         );
  AOI211_X1 U8233 ( .C1(REQUESTPENDING_REG_SCAN_IN), .C2(n7737), .A(n7736), 
        .B(n7735), .ZN(n7738) );
  OAI221_X1 U8234 ( .B1(n7739), .B2(READY_N), .C1(n7739), .C2(n7740), .A(n7738), .ZN(n7743) );
  NAND4_X1 U8235 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(STATE_REG_0__SCAN_IN), 
        .A3(n7741), .A4(n7740), .ZN(n7742) );
  OAI211_X1 U8236 ( .C1(n7745), .C2(n7744), .A(n7743), .B(n7742), .ZN(U3183)
         );
  AOI22_X1 U8237 ( .A1(n7734), .A2(n7748), .B1(n7747), .B2(n7746), .ZN(U3473)
         );
  INV_X1 U8238 ( .A(n7759), .ZN(n7750) );
  OAI22_X1 U8239 ( .A1(n7752), .A2(n7751), .B1(n7750), .B2(n7749), .ZN(n7753)
         );
  INV_X1 U8240 ( .A(n7753), .ZN(n7755) );
  AOI22_X1 U8241 ( .A1(n7763), .A2(DATAI_0_), .B1(n7762), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n7754) );
  NAND2_X1 U8242 ( .A1(n7755), .A2(n7754), .ZN(U2875) );
  AOI22_X1 U8243 ( .A1(n7756), .A2(n7760), .B1(DATAI_18_), .B2(n7759), .ZN(
        n7758) );
  AOI22_X1 U8244 ( .A1(n7763), .A2(DATAI_2_), .B1(n7762), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n7757) );
  NAND2_X1 U8245 ( .A1(n7758), .A2(n7757), .ZN(U2873) );
  AOI22_X1 U8246 ( .A1(n7761), .A2(n7760), .B1(n7759), .B2(DATAI_20_), .ZN(
        n7765) );
  AOI22_X1 U8247 ( .A1(n7763), .A2(DATAI_4_), .B1(n7762), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n7764) );
  NAND2_X1 U8248 ( .A1(n7765), .A2(n7764), .ZN(U2871) );
  CLKBUF_X3 U3815 ( .A(n4397), .Z(n3628) );
  CLKBUF_X2 U3672 ( .A(n4397), .Z(n3652) );
  AND2_X1 U3857 ( .A1(n3760), .A2(n5796), .ZN(n4352) );
  INV_X1 U3660 ( .A(n3836), .ZN(n4146) );
  BUF_X1 U3668 ( .A(n4032), .Z(n3658) );
  AND2_X1 U3674 ( .A1(n5770), .A2(n5799), .ZN(n4104) );
  CLKBUF_X1 U3676 ( .A(n4096), .Z(n3634) );
  CLKBUF_X1 U3684 ( .A(n5135), .Z(n5327) );
  NAND2_X1 U3691 ( .A1(n5428), .A2(n5415), .ZN(n7530) );
  CLKBUF_X1 U3698 ( .A(n5436), .Z(n3645) );
  OR2_X1 U3713 ( .A1(n5512), .A2(n6255), .ZN(n7766) );
  OR2_X4 U3806 ( .A1(n4220), .A2(n4218), .ZN(n4245) );
  NAND2_X1 U3817 ( .A1(n4096), .A2(n3979), .ZN(n4093) );
  NOR2_X1 U3835 ( .A1(n5564), .A2(n6067), .ZN(n7767) );
  CLKBUF_X1 U3841 ( .A(n3898), .Z(n6067) );
  CLKBUF_X1 U3860 ( .A(n3622), .Z(n4010) );
endmodule

