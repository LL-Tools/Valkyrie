

module b17_C_SARLock_k_64_6 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, U355, U356, U357, U358, 
        U359, U360, U361, U362, U363, U364, U366, U367, U368, U369, U370, U371, 
        U372, U373, U374, U375, U347, U348, U349, U350, U351, U352, U353, U354, 
        U365, U376, U247, U246, U245, U244, U243, U242, U241, U240, U239, U238, 
        U237, U236, U235, U234, U233, U232, U231, U230, U229, U228, U227, U226, 
        U225, U224, U223, U222, U221, U220, U219, U218, U217, U216, U251, U252, 
        U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, 
        U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, 
        U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274, 
        P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, 
        P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, 
        P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, 
        P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, 
        P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, 
        P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, 
        P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, 
        P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, 
        P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, 
        P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, 
        P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, 
        P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, 
        P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, 
        P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, 
        P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, 
        P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, 
        P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, 
        P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, 
        P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, 
        P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, 
        P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, 
        P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, 
        P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, 
        P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, 
        P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, 
        P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, 
        P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, 
        P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, 
        P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, 
        P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, 
        P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, 
        P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, 
        P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, 
        P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, 
        P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, 
        P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, 
        P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, 
        P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, 
        P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, 
        P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, 
        P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, 
        P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, 
        P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, 
        P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, 
        P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, 
        P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, 
        P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, 
        P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, 
        P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, 
        P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, 
        P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, 
        P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, 
        P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, 
        P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, 
        P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, 
        P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, 
        P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, 
        P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, 
        P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, 
        P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, 
        P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, 
        P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, 
        P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, 
        P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, 
        P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, 
        P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, 
        P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, 
        P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, 
        P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, 
        P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, 
        P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, 
        P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, 
        P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, 
        P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, 
        P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, 
        P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, 
        P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, 
        P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, 
        P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, 
        P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, 
        P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, 
        P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, 
        P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, 
        P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, 
        P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, 
        P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, 
        P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, 
        P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, 
        P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, 
        P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, 
        P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, 
        P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, 
        P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, 
        P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, 
        P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, 
        P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, 
        P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, 
        P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, 
        P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, 
        P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, 
        P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, 
        P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, 
        P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, 
        P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, 
        P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, 
        P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, 
        P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, 
        P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, 
        P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, 
        P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, 
        P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, 
        P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, 
        P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, 
        P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, 
        P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, 
        P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, 
        P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, 
        P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, 
        P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, 
        P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, 
        P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, 
        P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, 
        P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, 
        P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, 
        P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, 
        P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, 
        P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, 
        P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, 
        P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, 
        P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, 
        P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, 
        P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, 
        P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, 
        P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, 
        P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, 
        P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, 
        P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, 
        P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, 
        P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, 
        P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, 
        P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, 
        P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, 
        P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, 
        P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, 
        P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, 
        P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, 
        P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, 
        P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, 
        P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, 
        P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, 
        P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, 
        P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, 
        P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, 
        P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, 
        P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, 
        P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, 
        P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, 
        P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, 
        P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, 
        P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, 
        P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, 
        P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, 
        P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, 
        P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, 
        P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, 
        P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, 
        P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, 
        P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, 
        P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, 
        P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, 
        P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, 
        P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, 
        P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, 
        P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, 
        P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, 
        P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, 
        P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, 
        P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, 
        P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, 
        P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, 
        P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9610,
         n9611, n9612, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
         n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
         n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
         n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
         n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
         n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
         n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
         n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
         n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123,
         n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
         n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
         n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
         n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
         n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
         n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
         n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
         n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411,
         n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
         n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
         n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18946, n18947, n18948,
         n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956,
         n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
         n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972,
         n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
         n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988,
         n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996,
         n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
         n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
         n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020,
         n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028,
         n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
         n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044,
         n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
         n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
         n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
         n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076,
         n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
         n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
         n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100,
         n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
         n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
         n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
         n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132,
         n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140,
         n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
         n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
         n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
         n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172,
         n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
         n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
         n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
         n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204,
         n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212,
         n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
         n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
         n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236,
         n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244,
         n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
         n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260,
         n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
         n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276,
         n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284,
         n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292,
         n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
         n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308,
         n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316,
         n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
         n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332,
         n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340,
         n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348,
         n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
         n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364,
         n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372,
         n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380,
         n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388,
         n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
         n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404,
         n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412,
         n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420,
         n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428,
         n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436,
         n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
         n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452,
         n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460,
         n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468,
         n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476,
         n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484,
         n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492,
         n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500,
         n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508,
         n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
         n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524,
         n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532,
         n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540,
         n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548,
         n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556,
         n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564,
         n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572,
         n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580,
         n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
         n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596,
         n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604,
         n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612,
         n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620,
         n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628,
         n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636,
         n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644,
         n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
         n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
         n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668,
         n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676,
         n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684,
         n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692,
         n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700,
         n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708,
         n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716,
         n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724,
         n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732,
         n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740,
         n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748,
         n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756,
         n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764,
         n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772,
         n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780,
         n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788,
         n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796,
         n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
         n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812,
         n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820,
         n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
         n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836,
         n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844,
         n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852,
         n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860,
         n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868,
         n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
         n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884,
         n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892,
         n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900,
         n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908,
         n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916,
         n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924,
         n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932,
         n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
         n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
         n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956,
         n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964,
         n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972,
         n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980,
         n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988,
         n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996,
         n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004,
         n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012,
         n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
         n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028,
         n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036,
         n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044,
         n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052,
         n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060,
         n20061, n20062, n20063, n20064, n20066, n20067, n20068, n20069,
         n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077,
         n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085,
         n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093,
         n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
         n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109,
         n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117,
         n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125,
         n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133,
         n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141,
         n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149,
         n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157,
         n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165,
         n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
         n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181,
         n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189,
         n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197,
         n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205,
         n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213,
         n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221,
         n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229,
         n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237,
         n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245,
         n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253,
         n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261,
         n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269,
         n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277,
         n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285,
         n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293,
         n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301,
         n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309,
         n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317,
         n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325,
         n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333,
         n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341,
         n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349,
         n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357,
         n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365,
         n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373,
         n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381,
         n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389,
         n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397,
         n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405,
         n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413,
         n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421,
         n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429,
         n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437,
         n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445,
         n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453,
         n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461,
         n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469,
         n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477,
         n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485,
         n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493,
         n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501,
         n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509,
         n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517,
         n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525,
         n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533,
         n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541,
         n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549,
         n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557,
         n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565,
         n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573,
         n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581,
         n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589,
         n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597,
         n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605,
         n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613,
         n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621,
         n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
         n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637,
         n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645,
         n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653,
         n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661,
         n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669,
         n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
         n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685,
         n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693,
         n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701,
         n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709,
         n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717,
         n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725,
         n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733,
         n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741,
         n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
         n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757,
         n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765,
         n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773,
         n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781,
         n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789,
         n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797,
         n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805,
         n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813,
         n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
         n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829,
         n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837,
         n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845,
         n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853,
         n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861,
         n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869,
         n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877,
         n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885,
         n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
         n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901,
         n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909,
         n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917,
         n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925,
         n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933,
         n20934;

  INV_X1 U11044 ( .A(n17518), .ZN(n17738) );
  AOI21_X1 U11045 ( .B1(n14074), .B2(n14084), .A(n14073), .ZN(n14367) );
  INV_X2 U11046 ( .A(n20036), .ZN(n10704) );
  CLKBUF_X2 U11047 ( .A(n10496), .Z(n9611) );
  INV_X2 U11048 ( .A(n12901), .ZN(n9927) );
  AND2_X2 U11049 ( .A1(n20074), .A2(n20080), .ZN(n10677) );
  XNOR2_X1 U11050 ( .A(n10824), .B(n10823), .ZN(n17712) );
  AND2_X1 U11051 ( .A1(n13271), .A2(n13245), .ZN(n13545) );
  INV_X1 U11052 ( .A(n16910), .ZN(n17087) );
  OAI21_X1 U11053 ( .B1(n9780), .B2(n17736), .A(n9779), .ZN(n10824) );
  BUF_X2 U11054 ( .A(n10741), .Z(n17105) );
  OR2_X1 U11055 ( .A1(n10376), .A2(n10120), .ZN(n10335) );
  CLKBUF_X2 U11056 ( .A(n11753), .Z(n14967) );
  AND2_X1 U11057 ( .A1(n14903), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12057) );
  NAND2_X1 U11058 ( .A1(n10259), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10327) );
  CLKBUF_X2 U11059 ( .A(n10223), .Z(n11515) );
  INV_X2 U11060 ( .A(n9645), .ZN(n17104) );
  CLKBUF_X2 U11061 ( .A(n10761), .Z(n17081) );
  CLKBUF_X1 U11062 ( .A(n10867), .Z(n16954) );
  NAND2_X1 U11063 ( .A1(n13352), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11851) );
  NOR2_X1 U11064 ( .A1(n10573), .A2(n13440), .ZN(n12636) );
  NAND2_X2 U11065 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13810) );
  CLKBUF_X2 U11066 ( .A(n10175), .Z(n9615) );
  CLKBUF_X2 U11067 ( .A(n10185), .Z(n11510) );
  NAND4_X1 U11068 ( .A1(n10174), .A2(n10173), .A3(n10172), .A4(n10171), .ZN(
        n13390) );
  NAND2_X1 U11069 ( .A1(n13315), .A2(n11778), .ZN(n11904) );
  AND4_X1 U11070 ( .A1(n10202), .A2(n10201), .A3(n10200), .A4(n10199), .ZN(
        n10218) );
  AND2_X1 U11071 ( .A1(n10134), .A2(n10136), .ZN(n10342) );
  NAND2_X1 U11072 ( .A1(n11682), .A2(n11681), .ZN(n11768) );
  AND2_X1 U11073 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10136) );
  INV_X1 U11074 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9816) );
  CLKBUF_X2 U11075 ( .A(n11755), .Z(n9601) );
  XNOR2_X1 U11076 ( .A(n10474), .B(n10473), .ZN(n11117) );
  AND2_X1 U11077 ( .A1(n12961), .A2(n10134), .ZN(n10223) );
  NAND2_X1 U11078 ( .A1(n12635), .A2(n20092), .ZN(n12325) );
  OR2_X1 U11079 ( .A1(n12528), .A2(n15640), .ZN(n12524) );
  INV_X1 U11080 ( .A(n11851), .ZN(n11838) );
  NAND2_X1 U11081 ( .A1(n11706), .A2(n9827), .ZN(n11789) );
  NAND2_X1 U11082 ( .A1(n12536), .A2(n13342), .ZN(n15591) );
  AND4_X1 U11083 ( .A1(n10124), .A2(n10123), .A3(n10122), .A4(n10121), .ZN(
        n10174) );
  AND2_X1 U11084 ( .A1(n9606), .A2(n11637), .ZN(n14867) );
  NAND2_X1 U11085 ( .A1(n13820), .A2(n13819), .ZN(n10024) );
  NAND2_X1 U11086 ( .A1(n12772), .A2(n13002), .ZN(n12690) );
  AND2_X1 U11087 ( .A1(n13271), .A2(n13270), .ZN(n19569) );
  INV_X1 U11088 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11637) );
  NOR2_X1 U11090 ( .A1(n18136), .A2(n16776), .ZN(n10984) );
  INV_X1 U11091 ( .A(n19961), .ZN(n19950) );
  NOR2_X2 U11092 ( .A1(n14095), .A2(n14096), .ZN(n14082) );
  OR2_X1 U11093 ( .A1(n9655), .A2(n11050), .ZN(n10683) );
  INV_X1 U11094 ( .A(n10677), .ZN(n12817) );
  NOR2_X1 U11096 ( .A1(n15004), .A2(n15003), .ZN(n15002) );
  NAND2_X1 U11097 ( .A1(n11590), .A2(n11589), .ZN(n12901) );
  INV_X2 U11098 ( .A(n11773), .ZN(n12772) );
  AND2_X1 U11099 ( .A1(n13625), .A2(n13624), .ZN(n13646) );
  INV_X1 U11100 ( .A(n11798), .ZN(n14935) );
  INV_X1 U11101 ( .A(n17240), .ZN(n18136) );
  NAND2_X1 U11102 ( .A1(n10829), .A2(n16339), .ZN(n17677) );
  NAND2_X1 U11103 ( .A1(n17964), .A2(n18552), .ZN(n17883) );
  AOI221_X1 U11104 ( .B1(n17964), .B2(n17930), .C1(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n17930), .A(n9612), .ZN(
        n17932) );
  OAI21_X1 U11105 ( .B1(n14120), .B2(n14110), .A(n14109), .ZN(n14390) );
  CLKBUF_X3 U11106 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n16257) );
  NAND3_X2 U11107 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11670) );
  OR2_X1 U11108 ( .A1(n10732), .A2(n18560), .ZN(n9599) );
  OR2_X2 U11109 ( .A1(n14919), .A2(n14918), .ZN(n9600) );
  NOR2_X2 U11110 ( .A1(n17725), .A2(n17727), .ZN(n17708) );
  AND2_X2 U11111 ( .A1(n13215), .A2(n9673), .ZN(n13625) );
  AOI21_X2 U11112 ( .B1(n15857), .B2(n15856), .A(n18600), .ZN(n17151) );
  NOR2_X2 U11113 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n10848), .ZN(
        n16340) );
  AND2_X4 U11114 ( .A1(n11947), .A2(n11737), .ZN(n11752) );
  BUF_X2 U11115 ( .A(n11755), .Z(n9602) );
  BUF_X2 U11116 ( .A(n11755), .Z(n9603) );
  AND2_X1 U11117 ( .A1(n11948), .A2(n11737), .ZN(n11755) );
  NAND3_X1 U11118 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9604) );
  INV_X4 U11119 ( .A(n11670), .ZN(n14903) );
  NOR2_X2 U11120 ( .A1(n17780), .A2(n15842), .ZN(n16319) );
  NAND2_X1 U11121 ( .A1(n13352), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9605) );
  NOR2_X1 U11122 ( .A1(n17720), .A2(n17719), .ZN(n17718) );
  INV_X4 U11123 ( .A(n11765), .ZN(n11798) );
  AND2_X1 U11124 ( .A1(n12546), .A2(n15573), .ZN(n9606) );
  AND2_X2 U11125 ( .A1(n12546), .A2(n15573), .ZN(n9607) );
  AND2_X1 U11126 ( .A1(n12546), .A2(n15573), .ZN(n11946) );
  INV_X2 U11127 ( .A(n13267), .ZN(n19157) );
  AND3_X1 U11128 ( .A1(n13271), .A2(n13224), .A3(n13267), .ZN(n13669) );
  AND2_X2 U11129 ( .A1(n13286), .A2(n13267), .ZN(n15629) );
  INV_X1 U11133 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9610) );
  NAND2_X1 U11134 ( .A1(n15043), .A2(n9710), .ZN(n15031) );
  NOR2_X2 U11135 ( .A1(n14986), .A2(n14958), .ZN(n14982) );
  AND2_X4 U11136 ( .A1(n11937), .A2(n11737), .ZN(n11756) );
  AND2_X4 U11137 ( .A1(n11937), .A2(n16257), .ZN(n11754) );
  INV_X1 U11138 ( .A(n10006), .ZN(n13660) );
  NOR2_X1 U11139 ( .A1(n17703), .A2(n18019), .ZN(n17702) );
  AND2_X1 U11140 ( .A1(n11845), .A2(n11844), .ZN(n12819) );
  NOR2_X1 U11141 ( .A1(n18750), .A2(n17407), .ZN(n17408) );
  OR2_X1 U11142 ( .A1(n16462), .A2(n18753), .ZN(n15759) );
  NAND2_X1 U11143 ( .A1(n11931), .A2(n12510), .ZN(n12440) );
  INV_X1 U11144 ( .A(n10261), .ZN(n12624) );
  AND2_X1 U11145 ( .A1(n10250), .A2(n20105), .ZN(n10262) );
  INV_X1 U11146 ( .A(n11768), .ZN(n11794) );
  INV_X1 U11147 ( .A(n20092), .ZN(n12634) );
  AND4_X1 U11148 ( .A1(n10238), .A2(n10237), .A3(n10236), .A4(n10235), .ZN(
        n10239) );
  AND4_X1 U11149 ( .A1(n10210), .A2(n10209), .A3(n10208), .A4(n10207), .ZN(
        n10216) );
  INV_X4 U11150 ( .A(n17103), .ZN(n17067) );
  CLKBUF_X2 U11151 ( .A(n10278), .Z(n11538) );
  CLKBUF_X2 U11152 ( .A(n10852), .Z(n9618) );
  CLKBUF_X3 U11153 ( .A(n10852), .Z(n9614) );
  CLKBUF_X2 U11154 ( .A(n10342), .Z(n11533) );
  BUF_X2 U11155 ( .A(n10273), .Z(n11539) );
  INV_X2 U11156 ( .A(n18069), .ZN(n9612) );
  AND2_X1 U11157 ( .A1(n14643), .A2(n10135), .ZN(n10273) );
  INV_X1 U11158 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10725) );
  AOI211_X1 U11159 ( .C1(n15318), .C2(n19156), .A(n15317), .B(n15316), .ZN(
        n15319) );
  NAND2_X1 U11160 ( .A1(n9956), .A2(n9953), .ZN(n9951) );
  OAI21_X1 U11161 ( .B1(n15264), .B2(n15196), .A(n15263), .ZN(n15782) );
  XNOR2_X1 U11162 ( .A(n9852), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9886) );
  NAND2_X1 U11163 ( .A1(n15488), .A2(n15460), .ZN(n16179) );
  NOR2_X1 U11164 ( .A1(n15168), .A2(n15167), .ZN(n15157) );
  NAND2_X1 U11165 ( .A1(n13950), .A2(n9814), .ZN(n15358) );
  AOI21_X1 U11166 ( .B1(n10014), .B2(n9627), .A(n9667), .ZN(n15168) );
  NAND2_X1 U11167 ( .A1(n14363), .A2(n9823), .ZN(n14355) );
  NAND2_X1 U11168 ( .A1(n9855), .A2(n9854), .ZN(n14354) );
  AOI211_X1 U11169 ( .C1(n15976), .C2(n14393), .A(n14392), .B(n14391), .ZN(
        n14394) );
  NAND2_X1 U11170 ( .A1(n14085), .A2(n14084), .ZN(n14375) );
  AND2_X1 U11171 ( .A1(n10044), .A2(n10511), .ZN(n14363) );
  AND2_X1 U11172 ( .A1(n9965), .A2(n9963), .ZN(n15241) );
  OAI21_X1 U11173 ( .B1(n14379), .B2(n10045), .A(n14437), .ZN(n10044) );
  NAND2_X1 U11174 ( .A1(n9770), .A2(n9768), .ZN(n12343) );
  NAND2_X1 U11175 ( .A1(n13851), .A2(n13850), .ZN(n10025) );
  NAND2_X1 U11176 ( .A1(n15009), .A2(n15008), .ZN(n15007) );
  NAND2_X1 U11177 ( .A1(n13692), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13940) );
  NAND2_X1 U11178 ( .A1(n9769), .A2(n9767), .ZN(n9768) );
  AND2_X1 U11179 ( .A1(n9765), .A2(n9764), .ZN(n9770) );
  NAND2_X1 U11180 ( .A1(n13691), .A2(n13690), .ZN(n13692) );
  AOI21_X1 U11181 ( .B1(n9761), .B2(n13842), .A(n9760), .ZN(n9759) );
  XNOR2_X1 U11182 ( .A(n13946), .B(n15555), .ZN(n15544) );
  AND2_X1 U11183 ( .A1(n9913), .A2(n9914), .ZN(n17416) );
  NAND2_X1 U11184 ( .A1(n9862), .A2(n10506), .ZN(n14450) );
  INV_X1 U11185 ( .A(n13945), .ZN(n13947) );
  NAND2_X1 U11186 ( .A1(n15025), .A2(n15024), .ZN(n15023) );
  INV_X1 U11187 ( .A(n15031), .ZN(n14883) );
  NAND2_X1 U11188 ( .A1(n9824), .A2(n10052), .ZN(n9864) );
  CLKBUF_X1 U11189 ( .A(n13941), .Z(n13945) );
  NAND2_X1 U11190 ( .A1(n9786), .A2(n9785), .ZN(n9789) );
  NAND3_X1 U11191 ( .A1(n13569), .A2(n13683), .A3(n13905), .ZN(n9831) );
  NAND2_X1 U11192 ( .A1(n9825), .A2(n15988), .ZN(n13606) );
  AND3_X1 U11193 ( .A1(n9861), .A2(n9679), .A3(n10050), .ZN(n9863) );
  AND2_X1 U11194 ( .A1(n9790), .A2(n9749), .ZN(n9785) );
  NAND2_X1 U11195 ( .A1(n9758), .A2(n13566), .ZN(n13683) );
  OR2_X1 U11196 ( .A1(n17452), .A2(n17797), .ZN(n9786) );
  NOR2_X1 U11197 ( .A1(n10505), .A2(n14455), .ZN(n10506) );
  NAND2_X1 U11198 ( .A1(n9848), .A2(n10471), .ZN(n15991) );
  NOR2_X1 U11199 ( .A1(n10009), .A2(n9847), .ZN(n9846) );
  XNOR2_X1 U11200 ( .A(n13489), .B(n13304), .ZN(n13484) );
  AND2_X1 U11201 ( .A1(n14457), .A2(n15962), .ZN(n15953) );
  OR2_X1 U11202 ( .A1(n13775), .A2(n10503), .ZN(n10505) );
  AOI21_X1 U11203 ( .B1(n10052), .B2(n10051), .A(n9664), .ZN(n10050) );
  AND2_X1 U11204 ( .A1(n9925), .A2(n9923), .ZN(n14694) );
  OR2_X1 U11205 ( .A1(n15980), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15956) );
  OR2_X1 U11206 ( .A1(n15980), .A2(n10501), .ZN(n15963) );
  OR2_X1 U11207 ( .A1(n15980), .A2(n10716), .ZN(n13777) );
  NAND4_X1 U11208 ( .A1(n10104), .A2(n13301), .A3(n13300), .A4(n10118), .ZN(
        n13490) );
  NAND2_X1 U11209 ( .A1(n20016), .A2(n20015), .ZN(n20014) );
  XNOR2_X1 U11210 ( .A(n10449), .B(n16104), .ZN(n16001) );
  AND4_X1 U11211 ( .A1(n13258), .A2(n13257), .A3(n13256), .A4(n13255), .ZN(
        n13281) );
  AND4_X1 U11212 ( .A1(n13295), .A2(n13294), .A3(n13293), .A4(n13292), .ZN(
        n13301) );
  NAND2_X1 U11213 ( .A1(n13099), .A2(n13098), .ZN(n13155) );
  INV_X1 U11214 ( .A(n17755), .ZN(n17768) );
  NAND2_X1 U11215 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17689), .ZN(
        n11028) );
  INV_X1 U11216 ( .A(n10441), .ZN(n10439) );
  INV_X1 U11217 ( .A(n9947), .ZN(n12833) );
  OR2_X2 U11218 ( .A1(n18539), .A2(n18600), .ZN(n16463) );
  AND2_X1 U11219 ( .A1(n9784), .A2(n17952), .ZN(n17676) );
  BUF_X2 U11220 ( .A(n13271), .Z(n15615) );
  OR2_X2 U11221 ( .A1(n13146), .A2(n10058), .ZN(n15494) );
  AND2_X1 U11222 ( .A1(n9778), .A2(n9670), .ZN(n10838) );
  CLKBUF_X1 U11223 ( .A(n20926), .Z(n17297) );
  CLKBUF_X1 U11224 ( .A(n12845), .Z(n12898) );
  AND2_X1 U11225 ( .A1(n11062), .A2(n10368), .ZN(n10369) );
  INV_X1 U11226 ( .A(n12819), .ZN(n9960) );
  AND2_X1 U11227 ( .A1(n10043), .A2(n9693), .ZN(n11057) );
  AND2_X1 U11228 ( .A1(n12611), .A2(n12596), .ZN(n13252) );
  OR2_X1 U11229 ( .A1(n11842), .A2(n11843), .ZN(n11845) );
  NAND2_X1 U11230 ( .A1(n10990), .A2(n18542), .ZN(n15765) );
  AND2_X1 U11231 ( .A1(n10336), .A2(n9818), .ZN(n9817) );
  AND2_X1 U11232 ( .A1(n10368), .A2(n10367), .ZN(n11058) );
  NOR2_X1 U11233 ( .A1(n12025), .A2(n12024), .ZN(n12048) );
  OAI211_X1 U11234 ( .C1(n15834), .C2(n20395), .A(n10335), .B(n10334), .ZN(
        n10336) );
  CLKBUF_X2 U11235 ( .A(n11826), .Z(n11914) );
  OR2_X1 U11236 ( .A1(n10365), .A2(n10366), .ZN(n10368) );
  NOR2_X1 U11237 ( .A1(n11594), .A2(n11585), .ZN(n11586) );
  OAI21_X1 U11238 ( .B1(n18114), .B2(n10989), .A(n10988), .ZN(n18546) );
  AOI21_X1 U11239 ( .B1(n13333), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n11809), 
        .ZN(n11810) );
  AND2_X1 U11240 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n11010), .ZN(
        n11011) );
  NAND2_X1 U11241 ( .A1(n10256), .A2(n9731), .ZN(n9730) );
  OR2_X1 U11242 ( .A1(n10981), .A2(n10980), .ZN(n10987) );
  NOR2_X1 U11243 ( .A1(n17285), .A2(n10820), .ZN(n10822) );
  NOR2_X1 U11244 ( .A1(n16834), .A2(n12346), .ZN(n16327) );
  AND2_X1 U11245 ( .A1(n11808), .A2(n12434), .ZN(n11771) );
  AOI21_X1 U11246 ( .B1(n10318), .B2(n20649), .A(n10317), .ZN(n10361) );
  OR2_X1 U11247 ( .A1(n12626), .A2(n12946), .ZN(n10246) );
  INV_X1 U11248 ( .A(n11991), .ZN(n12270) );
  AND2_X1 U11249 ( .A1(n12684), .A2(n11777), .ZN(n13352) );
  CLKBUF_X1 U11250 ( .A(n12558), .Z(n16276) );
  AND2_X2 U11251 ( .A1(n12020), .A2(n11933), .ZN(n11995) );
  INV_X1 U11252 ( .A(n10936), .ZN(n18114) );
  AND2_X1 U11253 ( .A1(n10251), .A2(n10262), .ZN(n10702) );
  NAND2_X1 U11254 ( .A1(n10245), .A2(n12636), .ZN(n12626) );
  CLKBUF_X1 U11255 ( .A(n10586), .Z(n12766) );
  OR2_X1 U11256 ( .A1(n12899), .A2(n10252), .ZN(n14637) );
  INV_X1 U11257 ( .A(n9902), .ZN(n17291) );
  NOR2_X1 U11258 ( .A1(n14262), .A2(n10243), .ZN(n10245) );
  AND3_X1 U11259 ( .A1(n9905), .A2(n10768), .A3(n10769), .ZN(n10815) );
  CLKBUF_X1 U11260 ( .A(n11797), .Z(n12700) );
  NOR2_X1 U11261 ( .A1(n12690), .A2(n13916), .ZN(n11788) );
  NAND3_X1 U11262 ( .A1(n10902), .A2(n10901), .A3(n10900), .ZN(n17154) );
  NOR2_X1 U11263 ( .A1(n10933), .A2(n10932), .ZN(n18101) );
  NAND2_X1 U11264 ( .A1(n12634), .A2(n20105), .ZN(n14262) );
  OR2_X1 U11265 ( .A1(n10759), .A2(n9903), .ZN(n9902) );
  INV_X1 U11266 ( .A(n11792), .ZN(n11787) );
  CLKBUF_X1 U11267 ( .A(n11800), .Z(n19181) );
  INV_X2 U11268 ( .A(U212), .ZN(n16399) );
  INV_X1 U11269 ( .A(n20098), .ZN(n12633) );
  OR2_X1 U11270 ( .A1(n10311), .A2(n10310), .ZN(n10478) );
  NAND2_X1 U11271 ( .A1(n11644), .A2(n11643), .ZN(n11800) );
  INV_X2 U11272 ( .A(n18134), .ZN(n18478) );
  NAND2_X1 U11273 ( .A1(n11705), .A2(n11704), .ZN(n13436) );
  NAND2_X1 U11274 ( .A1(n11693), .A2(n11692), .ZN(n13345) );
  NAND2_X1 U11275 ( .A1(n11657), .A2(n11656), .ZN(n11792) );
  OR2_X2 U11276 ( .A1(n10160), .A2(n10159), .ZN(n20092) );
  OR2_X2 U11277 ( .A1(n16411), .A2(n16357), .ZN(n16413) );
  AND3_X1 U11278 ( .A1(n10183), .A2(n10182), .A3(n10184), .ZN(n9622) );
  AND4_X1 U11279 ( .A1(n10133), .A2(n10132), .A3(n10131), .A4(n10130), .ZN(
        n10172) );
  AND4_X1 U11280 ( .A1(n10128), .A2(n10127), .A3(n10126), .A4(n10125), .ZN(
        n10173) );
  AND4_X1 U11281 ( .A1(n10206), .A2(n10205), .A3(n10204), .A4(n10203), .ZN(
        n10217) );
  NAND2_X1 U11282 ( .A1(n11667), .A2(n11666), .ZN(n11668) );
  NAND2_X1 U11283 ( .A1(n11662), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11669) );
  NOR2_X2 U11284 ( .A1(n13387), .A2(n15947), .ZN(n13388) );
  NAND2_X1 U11285 ( .A1(n9656), .A2(n11655), .ZN(n11656) );
  AND2_X1 U11286 ( .A1(n10177), .A2(n10176), .ZN(n10183) );
  INV_X2 U11287 ( .A(n12081), .ZN(n14868) );
  NAND2_X2 U11288 ( .A1(n18761), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18691) );
  NAND2_X2 U11289 ( .A1(n18761), .A2(n18631), .ZN(n18687) );
  AND3_X1 U11290 ( .A1(n11633), .A2(n11632), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11636) );
  AND4_X1 U11291 ( .A1(n11665), .A2(n11664), .A3(n11663), .A4(n11637), .ZN(
        n11667) );
  AND4_X1 U11292 ( .A1(n11661), .A2(n11660), .A3(n11659), .A4(n11658), .ZN(
        n11662) );
  AND4_X1 U11293 ( .A1(n10222), .A2(n10221), .A3(n10220), .A4(n10219), .ZN(
        n10242) );
  AND2_X1 U11294 ( .A1(n11646), .A2(n11645), .ZN(n11649) );
  INV_X2 U11295 ( .A(n12097), .ZN(n14861) );
  BUF_X2 U11296 ( .A(n10741), .Z(n17021) );
  AND4_X1 U11297 ( .A1(n11715), .A2(n11714), .A3(n11713), .A4(n11712), .ZN(
        n11716) );
  BUF_X2 U11298 ( .A(n10186), .Z(n11516) );
  INV_X2 U11299 ( .A(n16445), .ZN(U215) );
  AND2_X2 U11300 ( .A1(n9601), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12056) );
  BUF_X2 U11301 ( .A(n11754), .Z(n14966) );
  NOR2_X1 U11302 ( .A1(n18710), .A2(n18613), .ZN(n18747) );
  NAND2_X2 U11303 ( .A1(n19780), .A2(n19733), .ZN(n19787) );
  INV_X2 U11304 ( .A(n15722), .ZN(n15741) );
  BUF_X2 U11305 ( .A(n16928), .Z(n17101) );
  NOR2_X1 U11306 ( .A1(n9911), .A2(n10733), .ZN(n10760) );
  NOR2_X1 U11307 ( .A1(n10727), .A2(n10734), .ZN(n10761) );
  OR2_X1 U11308 ( .A1(n10732), .A2(n10733), .ZN(n17007) );
  BUF_X2 U11309 ( .A(n10225), .Z(n9619) );
  INV_X2 U11310 ( .A(n16451), .ZN(n16453) );
  NAND2_X1 U11311 ( .A1(n10725), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10734) );
  NAND2_X1 U11312 ( .A1(n9743), .A2(n10723), .ZN(n16825) );
  AND2_X1 U11313 ( .A1(n11631), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11936) );
  NAND3_X2 U11314 ( .A1(n18763), .A2(n12414), .A3(n18762), .ZN(n18069) );
  AND2_X1 U11315 ( .A1(n19853), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11809) );
  CLKBUF_X3 U11316 ( .A(n10725), .Z(n18717) );
  NAND2_X2 U11317 ( .A1(n19853), .A2(n19812), .ZN(n18921) );
  AND2_X2 U11318 ( .A1(n11948), .A2(n16257), .ZN(n11753) );
  NAND2_X1 U11319 ( .A1(n20898), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10733) );
  AND2_X1 U11320 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11947) );
  AND2_X1 U11321 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12546) );
  NAND2_X1 U11322 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18560) );
  NOR2_X2 U11323 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11948) );
  INV_X2 U11324 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10080) );
  NOR2_X2 U11325 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10135) );
  AND2_X2 U11326 ( .A1(n12607), .A2(n12606), .ZN(n12610) );
  INV_X2 U11327 ( .A(n15722), .ZN(n9616) );
  XNOR2_X2 U11328 ( .A(n14899), .B(n9700), .ZN(n15004) );
  NAND2_X2 U11329 ( .A1(n15007), .A2(n14896), .ZN(n14899) );
  INV_X2 U11330 ( .A(n17666), .ZN(n17678) );
  AND2_X2 U11331 ( .A1(n14756), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12053) );
  NOR2_X2 U11332 ( .A1(n9738), .A2(n9737), .ZN(n13465) );
  NAND2_X1 U11333 ( .A1(n10474), .A2(n10486), .ZN(n10496) );
  NAND2_X1 U11334 ( .A1(n9741), .A2(n10369), .ZN(n10403) );
  OAI22_X2 U11335 ( .A1(n17954), .A2(n17768), .B1(n12354), .B2(n17952), .ZN(
        n17642) );
  NAND2_X1 U11336 ( .A1(n17759), .A2(n17278), .ZN(n12354) );
  INV_X1 U11337 ( .A(n17066), .ZN(n9617) );
  INV_X4 U11338 ( .A(n9647), .ZN(n17089) );
  AND2_X2 U11339 ( .A1(n19865), .A2(n19416), .ZN(n12279) );
  NOR2_X4 U11340 ( .A1(n14236), .A2(n14235), .ZN(n14226) );
  AND2_X1 U11341 ( .A1(n10135), .A2(n14642), .ZN(n10185) );
  BUF_X4 U11342 ( .A(n10225), .Z(n9620) );
  AND2_X1 U11343 ( .A1(n14642), .A2(n10136), .ZN(n10225) );
  NOR2_X4 U11344 ( .A1(n18559), .A2(n18566), .ZN(n17964) );
  AND2_X1 U11345 ( .A1(n10129), .A2(n12961), .ZN(n9621) );
  NOR2_X4 U11346 ( .A1(n15660), .A2(n16463), .ZN(n17755) );
  NOR2_X1 U11347 ( .A1(n10734), .A2(n10733), .ZN(n10852) );
  NAND2_X1 U11348 ( .A1(n9757), .A2(n13682), .ZN(n13941) );
  INV_X1 U11349 ( .A(n13685), .ZN(n13682) );
  INV_X1 U11350 ( .A(n13683), .ZN(n9757) );
  AND2_X1 U11351 ( .A1(n11794), .A2(n13436), .ZN(n13342) );
  NOR2_X1 U11352 ( .A1(n20927), .A2(n10826), .ZN(n10829) );
  NAND2_X1 U11353 ( .A1(n14679), .A2(n14680), .ZN(n14684) );
  NAND2_X1 U11354 ( .A1(n14787), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12089) );
  INV_X1 U11355 ( .A(n15159), .ZN(n9847) );
  INV_X1 U11356 ( .A(n18109), .ZN(n10981) );
  NAND2_X1 U11357 ( .A1(n18119), .A2(n18127), .ZN(n10980) );
  INV_X1 U11358 ( .A(n13414), .ZN(n11140) );
  NAND2_X1 U11359 ( .A1(n10463), .A2(n10442), .ZN(n9851) );
  INV_X1 U11360 ( .A(n13444), .ZN(n11375) );
  INV_X1 U11361 ( .A(n13803), .ZN(n9895) );
  OR2_X1 U11362 ( .A1(n10662), .A2(n12817), .ZN(n10680) );
  NAND2_X1 U11363 ( .A1(n12936), .A2(n10375), .ZN(n10401) );
  INV_X2 U11364 ( .A(n12255), .ZN(n14862) );
  NAND2_X1 U11365 ( .A1(n9973), .A2(n15414), .ZN(n9972) );
  INV_X1 U11366 ( .A(n13948), .ZN(n9973) );
  NOR2_X1 U11367 ( .A1(n9975), .A2(n15544), .ZN(n9974) );
  NAND2_X1 U11368 ( .A1(n15282), .A2(n15414), .ZN(n9975) );
  NAND2_X1 U11369 ( .A1(n15157), .A2(n15159), .ZN(n13976) );
  NAND3_X1 U11370 ( .A1(n10026), .A2(n10025), .A3(n9839), .ZN(n9838) );
  NOR2_X1 U11371 ( .A1(n9633), .A2(n15276), .ZN(n9839) );
  AND2_X1 U11372 ( .A1(n9678), .A2(n10004), .ZN(n10003) );
  INV_X1 U11373 ( .A(n13710), .ZN(n10004) );
  AND2_X1 U11374 ( .A1(n11955), .A2(n13826), .ZN(n11991) );
  NOR2_X1 U11375 ( .A1(n14935), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11955) );
  INV_X1 U11376 ( .A(n13110), .ZN(n9990) );
  NAND3_X1 U11377 ( .A1(n9812), .A2(n9813), .A3(n13585), .ZN(n13937) );
  INV_X1 U11378 ( .A(n13658), .ZN(n9812) );
  NAND2_X1 U11379 ( .A1(n10027), .A2(n13700), .ZN(n13821) );
  AND2_X1 U11380 ( .A1(n13342), .A2(n11776), .ZN(n11777) );
  NOR2_X1 U11381 ( .A1(n17698), .A2(n10828), .ZN(n10831) );
  NAND2_X1 U11382 ( .A1(n9624), .A2(n9659), .ZN(n9780) );
  XNOR2_X1 U11383 ( .A(n10817), .B(n11001), .ZN(n10818) );
  OAI21_X1 U11384 ( .B1(n17748), .B2(n17747), .A(n9665), .ZN(n9910) );
  AND2_X1 U11385 ( .A1(n14437), .A2(n14499), .ZN(n9823) );
  NAND2_X1 U11386 ( .A1(n10506), .A2(n10052), .ZN(n9860) );
  NAND2_X1 U11387 ( .A1(n13606), .A2(n10490), .ZN(n10053) );
  NOR2_X1 U11388 ( .A1(n18810), .A2(n9937), .ZN(n9933) );
  AND2_X1 U11389 ( .A1(n13216), .A2(n13213), .ZN(n13214) );
  AND2_X1 U11390 ( .A1(n11587), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12823) );
  XNOR2_X1 U11391 ( .A(n15579), .B(n12787), .ZN(n12786) );
  OR2_X1 U11392 ( .A1(n12551), .A2(n9810), .ZN(n9756) );
  NOR2_X2 U11393 ( .A1(n10734), .A2(n18560), .ZN(n16928) );
  OAI21_X1 U11394 ( .B1(n14983), .B2(n18965), .A(n12315), .ZN(n12316) );
  AOI21_X1 U11395 ( .B1(n15066), .B2(n18907), .A(n12314), .ZN(n12315) );
  AND2_X1 U11396 ( .A1(n13565), .A2(n13564), .ZN(n13566) );
  NAND2_X1 U11397 ( .A1(n11838), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n11839) );
  AOI22_X1 U11398 ( .A1(n14756), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11713) );
  OR2_X1 U11399 ( .A1(n10956), .A2(n10957), .ZN(n10949) );
  NAND2_X1 U11400 ( .A1(n10702), .A2(n12635), .ZN(n10577) );
  OR2_X1 U11401 ( .A1(n10284), .A2(n10283), .ZN(n10357) );
  AND3_X1 U11402 ( .A1(n11768), .A2(n13436), .A3(n13345), .ZN(n9827) );
  INV_X1 U11403 ( .A(n13980), .ZN(n10008) );
  NAND2_X1 U11404 ( .A1(n13681), .A2(n13680), .ZN(n13685) );
  NOR2_X1 U11405 ( .A1(n12065), .A2(n12064), .ZN(n12066) );
  OR2_X1 U11406 ( .A1(n12060), .A2(n12059), .ZN(n12065) );
  NAND2_X1 U11407 ( .A1(n14967), .A2(n11637), .ZN(n12097) );
  NAND2_X1 U11408 ( .A1(n13287), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n13288) );
  NAND2_X1 U11409 ( .A1(n13674), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n13290) );
  NAND2_X1 U11410 ( .A1(n13249), .A2(n13264), .ZN(n10006) );
  AND3_X1 U11411 ( .A1(n11708), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n11707), .ZN(n11711) );
  NAND2_X1 U11412 ( .A1(n11731), .A2(n11723), .ZN(n11739) );
  INV_X1 U11413 ( .A(n10890), .ZN(n9752) );
  NAND2_X1 U11414 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n9751) );
  NOR2_X1 U11415 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11552) );
  AND2_X1 U11416 ( .A1(n11410), .A2(n9681), .ZN(n10088) );
  NAND2_X1 U11417 ( .A1(n11261), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11527) );
  NAND2_X1 U11418 ( .A1(n13741), .A2(n10081), .ZN(n14239) );
  NOR2_X1 U11419 ( .A1(n10083), .A2(n10082), .ZN(n10081) );
  INV_X1 U11420 ( .A(n14251), .ZN(n10082) );
  AND2_X1 U11421 ( .A1(n11216), .A2(n10091), .ZN(n10090) );
  OR2_X1 U11422 ( .A1(n13733), .A2(n13748), .ZN(n10091) );
  AND2_X1 U11423 ( .A1(n11092), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11101) );
  NAND2_X1 U11424 ( .A1(n12741), .A2(n10325), .ZN(n10374) );
  INV_X1 U11425 ( .A(n11170), .ZN(n11241) );
  INV_X1 U11426 ( .A(n11552), .ZN(n13444) );
  NAND2_X1 U11427 ( .A1(n14379), .A2(n14507), .ZN(n10511) );
  NAND2_X1 U11428 ( .A1(n14437), .A2(n10507), .ZN(n10040) );
  OR2_X1 U11429 ( .A1(n9632), .A2(n14437), .ZN(n10036) );
  NAND2_X1 U11430 ( .A1(n14232), .A2(n14229), .ZN(n9891) );
  INV_X1 U11431 ( .A(n13745), .ZN(n9896) );
  INV_X1 U11432 ( .A(n10462), .ZN(n10086) );
  OAI21_X1 U11433 ( .B1(n9851), .B2(n10484), .A(n10448), .ZN(n10449) );
  OR2_X1 U11434 ( .A1(n10677), .A2(n10674), .ZN(n10639) );
  AND2_X1 U11435 ( .A1(n9900), .A2(n12842), .ZN(n9899) );
  INV_X1 U11436 ( .A(n13100), .ZN(n9900) );
  INV_X1 U11437 ( .A(n20762), .ZN(n10479) );
  OR2_X1 U11438 ( .A1(n10295), .A2(n10294), .ZN(n10319) );
  OR2_X1 U11439 ( .A1(n10352), .A2(n10351), .ZN(n10353) );
  AND2_X2 U11440 ( .A1(n9816), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12961) );
  NAND2_X1 U11441 ( .A1(n9819), .A2(n10338), .ZN(n9818) );
  NAND2_X1 U11442 ( .A1(n12956), .A2(n20649), .ZN(n10394) );
  NOR2_X1 U11443 ( .A1(n9869), .A2(n9702), .ZN(n9867) );
  OR2_X1 U11444 ( .A1(n13858), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n13902) );
  NOR2_X1 U11445 ( .A1(n13860), .A2(n9872), .ZN(n9871) );
  INV_X1 U11446 ( .A(n9873), .ZN(n9872) );
  OR2_X1 U11447 ( .A1(n13864), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n13865) );
  NOR2_X1 U11448 ( .A1(n9876), .A2(n13873), .ZN(n9875) );
  INV_X1 U11449 ( .A(n9877), .ZN(n9876) );
  NAND2_X1 U11450 ( .A1(n13839), .A2(n11866), .ZN(n13847) );
  AND2_X1 U11451 ( .A1(n13833), .A2(n18918), .ZN(n13839) );
  NAND2_X1 U11452 ( .A1(n12303), .A2(n12302), .ZN(n13085) );
  NAND2_X1 U11453 ( .A1(n12301), .A2(n13826), .ZN(n12303) );
  NAND2_X1 U11454 ( .A1(n14967), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12255) );
  NAND2_X1 U11455 ( .A1(n14966), .A2(n11637), .ZN(n12081) );
  AND2_X1 U11456 ( .A1(n14935), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12776) );
  INV_X1 U11457 ( .A(n12393), .ZN(n10072) );
  OR2_X1 U11458 ( .A1(n11989), .A2(n11990), .ZN(n10066) );
  NAND2_X1 U11459 ( .A1(n9977), .A2(n9972), .ZN(n9967) );
  INV_X1 U11460 ( .A(n14698), .ZN(n10078) );
  AND2_X1 U11461 ( .A1(n16221), .A2(n15778), .ZN(n10076) );
  INV_X1 U11462 ( .A(n13649), .ZN(n10005) );
  AND2_X1 U11463 ( .A1(n10020), .A2(n13845), .ZN(n9834) );
  NAND2_X1 U11464 ( .A1(n13822), .A2(n10021), .ZN(n9761) );
  NOR2_X1 U11465 ( .A1(n15289), .A2(n10022), .ZN(n10021) );
  INV_X1 U11466 ( .A(n15548), .ZN(n10022) );
  INV_X1 U11467 ( .A(n9761), .ZN(n10020) );
  INV_X1 U11468 ( .A(n13939), .ZN(n9968) );
  INV_X1 U11469 ( .A(n13035), .ZN(n9992) );
  NAND2_X1 U11470 ( .A1(n13569), .A2(n13683), .ZN(n13586) );
  OR2_X1 U11471 ( .A1(n13586), .A2(n13597), .ZN(n13936) );
  NAND2_X1 U11472 ( .A1(n12552), .A2(n11836), .ZN(n12820) );
  OAI22_X1 U11473 ( .A1(n12584), .A2(P2_EBX_REG_1__SCAN_IN), .B1(n12575), .B2(
        n13916), .ZN(n12590) );
  INV_X1 U11474 ( .A(n11821), .ZN(n11822) );
  INV_X1 U11475 ( .A(n13436), .ZN(n13316) );
  NOR2_X1 U11476 ( .A1(n13269), .A2(n13252), .ZN(n13268) );
  INV_X1 U11477 ( .A(n10809), .ZN(n17103) );
  AND2_X1 U11478 ( .A1(n10837), .A2(n17564), .ZN(n9784) );
  XOR2_X1 U11479 ( .A(n17285), .B(n10820), .Z(n10821) );
  AOI211_X1 U11480 ( .C1(n18114), .C2(n10944), .A(n10943), .B(n10942), .ZN(
        n10988) );
  NAND2_X1 U11481 ( .A1(n17240), .A2(n10936), .ZN(n10995) );
  NAND2_X1 U11482 ( .A1(n12704), .A2(n12620), .ZN(n13448) );
  AND2_X1 U11483 ( .A1(n10595), .A2(n10594), .ZN(n12843) );
  OR2_X1 U11484 ( .A1(n19975), .A2(n12817), .ZN(n10595) );
  OR2_X1 U11485 ( .A1(n12800), .A2(n12950), .ZN(n12804) );
  INV_X1 U11486 ( .A(n20105), .ZN(n12765) );
  AND2_X1 U11487 ( .A1(n14353), .A2(n11564), .ZN(n11575) );
  OR2_X1 U11488 ( .A1(n11502), .A2(n20810), .ZN(n11507) );
  NAND2_X1 U11489 ( .A1(n13206), .A2(n9684), .ZN(n9737) );
  INV_X1 U11490 ( .A(n13464), .ZN(n10085) );
  NAND2_X1 U11491 ( .A1(n14378), .A2(n14387), .ZN(n14379) );
  OAI21_X1 U11492 ( .B1(n14417), .B2(n14369), .A(n14437), .ZN(n14387) );
  OR2_X1 U11493 ( .A1(n9646), .A2(n10661), .ZN(n14148) );
  NAND2_X1 U11494 ( .A1(n9864), .A2(n9863), .ZN(n9862) );
  OR2_X1 U11495 ( .A1(n14248), .A2(n14247), .ZN(n14250) );
  NAND2_X1 U11496 ( .A1(n15991), .A2(n15989), .ZN(n9825) );
  NOR2_X1 U11497 ( .A1(n14258), .A2(n14257), .ZN(n13210) );
  NAND2_X1 U11498 ( .A1(n13158), .A2(n10402), .ZN(n20016) );
  AND2_X1 U11499 ( .A1(n10581), .A2(n12763), .ZN(n10705) );
  NAND2_X1 U11500 ( .A1(n14718), .A2(n13815), .ZN(n13818) );
  OR2_X1 U11501 ( .A1(n13141), .A2(n19177), .ZN(n13917) );
  NOR2_X1 U11502 ( .A1(n13913), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n13919) );
  INV_X2 U11503 ( .A(n11787), .ZN(n13916) );
  NAND2_X1 U11504 ( .A1(n13902), .A2(n13917), .ZN(n12390) );
  OR2_X1 U11505 ( .A1(n9927), .A2(n18818), .ZN(n9936) );
  NAND2_X1 U11506 ( .A1(n13865), .A2(n13917), .ZN(n13870) );
  AND2_X1 U11507 ( .A1(n12249), .A2(n12248), .ZN(n16238) );
  INV_X1 U11508 ( .A(n9600), .ZN(n9956) );
  NAND3_X1 U11509 ( .A1(n9600), .A2(n9720), .A3(n9958), .ZN(n9955) );
  NAND2_X1 U11510 ( .A1(n14883), .A2(n9709), .ZN(n14884) );
  AND2_X1 U11511 ( .A1(n13342), .A2(n12548), .ZN(n12685) );
  NAND2_X1 U11512 ( .A1(n11601), .A2(n9711), .ZN(n11594) );
  NAND2_X1 U11513 ( .A1(n11601), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11600) );
  NAND2_X1 U11514 ( .A1(n11604), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11605) );
  NAND2_X1 U11515 ( .A1(n11612), .A2(n9941), .ZN(n11608) );
  NAND2_X1 U11516 ( .A1(n9842), .A2(n9841), .ZN(n15138) );
  AOI21_X1 U11517 ( .B1(n9844), .B2(n9722), .A(n10007), .ZN(n9841) );
  NAND2_X1 U11518 ( .A1(n15157), .A2(n9843), .ZN(n9842) );
  INV_X1 U11519 ( .A(n13975), .ZN(n10007) );
  INV_X1 U11520 ( .A(n9988), .ZN(n9986) );
  AND2_X1 U11521 ( .A1(n15027), .A2(n9715), .ZN(n14708) );
  INV_X1 U11522 ( .A(n14707), .ZN(n9997) );
  NAND2_X1 U11523 ( .A1(n9865), .A2(n13929), .ZN(n10018) );
  INV_X1 U11524 ( .A(n16129), .ZN(n9865) );
  NAND2_X1 U11525 ( .A1(n10013), .A2(n10019), .ZN(n10012) );
  NAND2_X1 U11526 ( .A1(n10016), .A2(n15386), .ZN(n10015) );
  NAND2_X1 U11527 ( .A1(n9838), .A2(n9837), .ZN(n10014) );
  NOR2_X1 U11528 ( .A1(n9626), .A2(n13900), .ZN(n9837) );
  INV_X1 U11529 ( .A(n9685), .ZN(n10016) );
  AND2_X1 U11530 ( .A1(n9838), .A2(n13899), .ZN(n15385) );
  NAND2_X1 U11531 ( .A1(n15039), .A2(n15040), .ZN(n15042) );
  NAND2_X1 U11532 ( .A1(n16237), .A2(n10076), .ZN(n15780) );
  NAND2_X1 U11533 ( .A1(n13628), .A2(n9678), .ZN(n13711) );
  NOR2_X1 U11534 ( .A1(n13527), .A2(n13526), .ZN(n13628) );
  OR2_X1 U11535 ( .A1(n13218), .A2(n13403), .ZN(n13527) );
  AND2_X1 U11536 ( .A1(n10024), .A2(n9686), .ZN(n15546) );
  NAND2_X1 U11537 ( .A1(n13944), .A2(n13943), .ZN(n15282) );
  INV_X1 U11538 ( .A(n13699), .ZN(n13684) );
  INV_X1 U11539 ( .A(n13936), .ZN(n13686) );
  NAND2_X1 U11540 ( .A1(n13584), .A2(n13591), .ZN(n9813) );
  NAND2_X1 U11541 ( .A1(n13493), .A2(n13492), .ZN(n13585) );
  NAND2_X1 U11542 ( .A1(n12912), .A2(n10067), .ZN(n13498) );
  NOR2_X1 U11543 ( .A1(n12049), .A2(n10070), .ZN(n10067) );
  CLKBUF_X1 U11544 ( .A(n13333), .Z(n15587) );
  AOI21_X1 U11545 ( .B1(n19157), .B2(n12823), .A(n12775), .ZN(n12785) );
  AND3_X1 U11546 ( .A1(n13268), .A2(n13267), .A3(n13271), .ZN(n19422) );
  AND2_X1 U11547 ( .A1(n13271), .A2(n13254), .ZN(n19453) );
  INV_X1 U11548 ( .A(n13826), .ZN(n19177) );
  OR2_X1 U11549 ( .A1(n19445), .A2(n19834), .ZN(n19565) );
  OR2_X1 U11550 ( .A1(n19813), .A2(n19814), .ZN(n19798) );
  INV_X1 U11551 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19852) );
  NOR2_X1 U11552 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n15616), .ZN(n16297) );
  NOR2_X1 U11553 ( .A1(n10982), .A2(n18593), .ZN(n16462) );
  OAI21_X1 U11554 ( .B1(n10964), .B2(n10966), .A(n10963), .ZN(n16461) );
  NOR2_X1 U11555 ( .A1(n18743), .A2(n18101), .ZN(n12428) );
  AOI211_X1 U11556 ( .C1(n17110), .C2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n10899), .B(n10898), .ZN(n10900) );
  NOR2_X1 U11557 ( .A1(n10766), .A2(n9906), .ZN(n9905) );
  NAND2_X1 U11558 ( .A1(n10991), .A2(n15765), .ZN(n15854) );
  INV_X1 U11559 ( .A(n17952), .ZN(n17644) );
  AOI21_X1 U11560 ( .B1(n11029), .B2(n11028), .A(n11027), .ZN(n17675) );
  INV_X1 U11561 ( .A(n9788), .ZN(n9787) );
  AND2_X1 U11562 ( .A1(n9787), .A2(n9789), .ZN(n10848) );
  NAND2_X1 U11563 ( .A1(n16342), .A2(n17564), .ZN(n9913) );
  INV_X1 U11564 ( .A(n16340), .ZN(n9914) );
  AND2_X1 U11565 ( .A1(n17451), .A2(n10114), .ZN(n9790) );
  OR2_X1 U11566 ( .A1(n17465), .A2(n17564), .ZN(n17451) );
  NAND2_X1 U11567 ( .A1(n17928), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17599) );
  OR2_X1 U11568 ( .A1(n18543), .A2(n18541), .ZN(n11034) );
  NAND2_X1 U11569 ( .A1(n17698), .A2(n9775), .ZN(n9772) );
  INV_X1 U11570 ( .A(n10830), .ZN(n9775) );
  NAND2_X1 U11571 ( .A1(n9774), .A2(n9661), .ZN(n9773) );
  INV_X1 U11572 ( .A(n17698), .ZN(n9774) );
  INV_X1 U11573 ( .A(n9910), .ZN(n10819) );
  INV_X1 U11574 ( .A(n17736), .ZN(n9782) );
  INV_X1 U11575 ( .A(n17722), .ZN(n9781) );
  NOR2_X1 U11576 ( .A1(n10969), .A2(n10935), .ZN(n15768) );
  INV_X1 U11577 ( .A(n16461), .ZN(n18536) );
  NOR2_X2 U11578 ( .A1(n10862), .A2(n10861), .ZN(n18750) );
  INV_X1 U11579 ( .A(n13448), .ZN(n20757) );
  AND2_X1 U11580 ( .A1(n14353), .A2(n14263), .ZN(n14344) );
  AND2_X1 U11581 ( .A1(n12800), .A2(n12328), .ZN(n20019) );
  INV_X1 U11582 ( .A(n20019), .ZN(n20030) );
  NAND2_X1 U11583 ( .A1(n9822), .A2(n9853), .ZN(n9852) );
  NAND2_X1 U11584 ( .A1(n14354), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9853) );
  NAND2_X1 U11585 ( .A1(n14355), .A2(n14489), .ZN(n9822) );
  XNOR2_X1 U11586 ( .A(n10682), .B(n10681), .ZN(n14202) );
  XNOR2_X1 U11587 ( .A(n9919), .B(n9918), .ZN(n11745) );
  INV_X1 U11588 ( .A(n14662), .ZN(n9918) );
  NAND2_X1 U11589 ( .A1(n9920), .A2(n12901), .ZN(n9919) );
  AND2_X1 U11590 ( .A1(n9926), .A2(n9924), .ZN(n9923) );
  INV_X1 U11591 ( .A(n15154), .ZN(n9924) );
  NAND2_X1 U11592 ( .A1(n18817), .A2(n9933), .ZN(n9932) );
  INV_X1 U11593 ( .A(n13530), .ZN(n9959) );
  INV_X1 U11594 ( .A(n19834), .ZN(n13421) );
  XNOR2_X1 U11595 ( .A(n14022), .B(n14021), .ZN(n14983) );
  NAND2_X1 U11596 ( .A1(n15299), .A2(n15300), .ZN(n10057) );
  NAND2_X1 U11597 ( .A1(n14684), .A2(n14683), .ZN(n15301) );
  OR2_X1 U11598 ( .A1(n15303), .A2(n16248), .ZN(n10055) );
  XNOR2_X1 U11599 ( .A(n9762), .B(n13981), .ZN(n15320) );
  NAND2_X1 U11600 ( .A1(n15321), .A2(n9663), .ZN(n9762) );
  INV_X1 U11601 ( .A(n19136), .ZN(n19155) );
  INV_X1 U11602 ( .A(n19166), .ZN(n19131) );
  INV_X1 U11603 ( .A(n19159), .ZN(n16228) );
  INV_X1 U11604 ( .A(n19814), .ZN(n19824) );
  INV_X1 U11605 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19811) );
  NAND2_X1 U11606 ( .A1(n12693), .A2(n12692), .ZN(n15579) );
  INV_X1 U11607 ( .A(n19385), .ZN(n19367) );
  INV_X1 U11608 ( .A(n18951), .ZN(n19713) );
  OR2_X1 U11609 ( .A1(n16503), .A2(n9794), .ZN(n9804) );
  NAND2_X1 U11610 ( .A1(n9801), .A2(n9800), .ZN(n9799) );
  OR2_X1 U11611 ( .A1(n16501), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n9800) );
  NAND2_X1 U11612 ( .A1(n9802), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n9801) );
  OR2_X1 U11613 ( .A1(n16495), .A2(n16841), .ZN(n9802) );
  NAND2_X1 U11614 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n16842), .ZN(n16827) );
  NAND2_X1 U11615 ( .A1(n18569), .A2(n17151), .ZN(n20928) );
  OAI21_X1 U11616 ( .B1(n12352), .B2(n17768), .A(n12351), .ZN(n12356) );
  OAI21_X1 U11617 ( .B1(n17792), .B2(n17678), .A(n9747), .ZN(n9746) );
  NAND2_X1 U11618 ( .A1(n9612), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n9747) );
  NOR2_X1 U11619 ( .A1(n17278), .A2(n17767), .ZN(n17666) );
  INV_X1 U11620 ( .A(n17759), .ZN(n17767) );
  NAND2_X1 U11621 ( .A1(n9763), .A2(n9771), .ZN(n9769) );
  OAI21_X1 U11622 ( .B1(n12352), .B2(n18079), .A(n11045), .ZN(n11046) );
  AND4_X1 U11623 ( .A1(n13558), .A2(n13557), .A3(n13556), .A4(n13555), .ZN(
        n13561) );
  INV_X1 U11624 ( .A(n10533), .ZN(n10520) );
  AOI22_X1 U11625 ( .A1(n11827), .A2(P2_REIP_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11782) );
  AND3_X1 U11626 ( .A1(n13663), .A2(n13662), .A3(n13661), .ZN(n13678) );
  AOI22_X1 U11627 ( .A1(n13660), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13256) );
  INV_X1 U11628 ( .A(n11904), .ZN(n11827) );
  AOI21_X1 U11629 ( .B1(n9607), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11646) );
  NAND2_X1 U11630 ( .A1(n9850), .A2(n12988), .ZN(n10441) );
  NOR2_X1 U11631 ( .A1(n10403), .A2(n9742), .ZN(n9850) );
  INV_X1 U11632 ( .A(n10425), .ZN(n9742) );
  AND2_X1 U11633 ( .A1(n10437), .A2(n10436), .ZN(n10440) );
  AND2_X1 U11634 ( .A1(n14449), .A2(n10042), .ZN(n10041) );
  INV_X1 U11635 ( .A(n10440), .ZN(n10438) );
  INV_X1 U11636 ( .A(n10318), .ZN(n10047) );
  INV_X1 U11637 ( .A(n10382), .ZN(n10314) );
  AOI21_X1 U11638 ( .B1(n20442), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n10516), .ZN(n10524) );
  NAND2_X1 U11639 ( .A1(n10259), .A2(n9731), .ZN(n9729) );
  AND2_X2 U11640 ( .A1(n12805), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10129) );
  AND2_X2 U11641 ( .A1(n10080), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10134) );
  OR2_X1 U11642 ( .A1(n10392), .A2(n10391), .ZN(n10444) );
  NOR2_X1 U11643 ( .A1(n12402), .A2(n9870), .ZN(n9869) );
  NOR2_X1 U11644 ( .A1(n13861), .A2(n9874), .ZN(n9873) );
  INV_X1 U11645 ( .A(n13869), .ZN(n9874) );
  NOR2_X1 U11646 ( .A1(n13852), .A2(n9878), .ZN(n9877) );
  NOR2_X1 U11647 ( .A1(n16257), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14758) );
  INV_X1 U11648 ( .A(n14884), .ZN(n9948) );
  INV_X1 U11649 ( .A(n13568), .ZN(n9758) );
  NAND2_X1 U11650 ( .A1(n11841), .A2(n10106), .ZN(n11842) );
  NAND2_X1 U11651 ( .A1(n11914), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11841) );
  OR2_X1 U11652 ( .A1(n12041), .A2(n12040), .ZN(n12299) );
  AOI22_X1 U11653 ( .A1(n14756), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9606), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11632) );
  NAND2_X1 U11654 ( .A1(n10760), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n9792) );
  NAND2_X1 U11655 ( .A1(n10761), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n9791) );
  AND2_X1 U11656 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n10827), .ZN(
        n10828) );
  NOR2_X1 U11657 ( .A1(n17291), .A2(n17300), .ZN(n10817) );
  AOI21_X1 U11658 ( .B1(n18575), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n10948), .ZN(n10957) );
  NAND2_X1 U11659 ( .A1(n10723), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10727) );
  OAI21_X1 U11660 ( .B1(n10256), .B2(n10259), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n10376) );
  NAND2_X1 U11661 ( .A1(n11249), .A2(n10084), .ZN(n10083) );
  INV_X1 U11662 ( .A(n14177), .ZN(n10084) );
  INV_X1 U11663 ( .A(n14163), .ZN(n10089) );
  NOR2_X1 U11664 ( .A1(n11281), .A2(n15906), .ZN(n11315) );
  INV_X1 U11665 ( .A(n13802), .ZN(n11249) );
  INV_X1 U11666 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11123) );
  NAND2_X1 U11667 ( .A1(n10087), .A2(n12988), .ZN(n10424) );
  INV_X1 U11668 ( .A(n10403), .ZN(n10087) );
  AND2_X1 U11669 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11079), .ZN(
        n11092) );
  INV_X1 U11670 ( .A(n14111), .ZN(n9893) );
  NAND2_X1 U11671 ( .A1(n14424), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10508) );
  INV_X1 U11672 ( .A(n10498), .ZN(n9861) );
  OR2_X1 U11673 ( .A1(n15980), .A2(n14610), .ZN(n10504) );
  OR2_X1 U11674 ( .A1(n15980), .A2(n10500), .ZN(n14466) );
  OR2_X1 U11675 ( .A1(n15980), .A2(n10499), .ZN(n14470) );
  INV_X1 U11676 ( .A(n10490), .ZN(n10051) );
  INV_X1 U11677 ( .A(n13606), .ZN(n9824) );
  OR2_X1 U11678 ( .A1(n10459), .A2(n10458), .ZN(n10476) );
  NAND2_X1 U11679 ( .A1(n10299), .A2(n10298), .ZN(n10324) );
  NAND2_X1 U11680 ( .A1(n11057), .A2(n20080), .ZN(n10299) );
  NAND2_X1 U11681 ( .A1(n10674), .A2(n10662), .ZN(n10586) );
  NAND2_X1 U11682 ( .A1(n10048), .A2(n10046), .ZN(n11069) );
  AOI21_X1 U11683 ( .B1(n10256), .B2(n10049), .A(n10047), .ZN(n10046) );
  NAND2_X1 U11684 ( .A1(n10259), .A2(n10049), .ZN(n10048) );
  NOR2_X1 U11685 ( .A1(n12805), .A2(n20649), .ZN(n10049) );
  OR2_X1 U11686 ( .A1(n20074), .A2(n20649), .ZN(n10381) );
  OR2_X1 U11687 ( .A1(n13390), .A2(n20649), .ZN(n10382) );
  AND2_X1 U11688 ( .A1(n10559), .A2(n10530), .ZN(n10558) );
  NAND2_X1 U11689 ( .A1(n10382), .A2(n10381), .ZN(n10550) );
  NAND2_X1 U11690 ( .A1(n20182), .A2(n10270), .ZN(n10340) );
  INV_X1 U11691 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20475) );
  OR2_X1 U11692 ( .A1(n11733), .A2(n11732), .ZN(n11726) );
  INV_X1 U11693 ( .A(n10103), .ZN(n9928) );
  OR2_X1 U11694 ( .A1(n14733), .A2(n9927), .ZN(n9929) );
  NAND2_X1 U11695 ( .A1(n13840), .A2(n9877), .ZN(n13875) );
  NAND2_X1 U11696 ( .A1(n13840), .A2(n13846), .ZN(n13853) );
  NOR2_X1 U11697 ( .A1(n13570), .A2(n9879), .ZN(n13833) );
  NAND2_X1 U11698 ( .A1(n9881), .A2(n9880), .ZN(n9879) );
  INV_X1 U11699 ( .A(n9882), .ZN(n9881) );
  NAND2_X1 U11700 ( .A1(n13115), .A2(n9884), .ZN(n9883) );
  INV_X1 U11701 ( .A(n12919), .ZN(n9884) );
  OR2_X1 U11702 ( .A1(n9883), .A2(n13140), .ZN(n9882) );
  OR2_X1 U11703 ( .A1(n11954), .A2(n11953), .ZN(n12307) );
  CLKBUF_X1 U11704 ( .A(n9601), .Z(n14968) );
  CLKBUF_X1 U11705 ( .A(n14756), .Z(n14971) );
  AND2_X1 U11706 ( .A1(n14726), .A2(n14710), .ZN(n10079) );
  INV_X1 U11707 ( .A(n15421), .ZN(n10073) );
  AND3_X1 U11708 ( .A1(n12106), .A2(n12105), .A3(n12104), .ZN(n13679) );
  NOR2_X1 U11709 ( .A1(n15172), .A2(n9939), .ZN(n9938) );
  INV_X1 U11710 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n9939) );
  AND2_X1 U11711 ( .A1(n9630), .A2(n11582), .ZN(n9941) );
  AND2_X1 U11712 ( .A1(n11614), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11612) );
  NAND2_X1 U11713 ( .A1(n9945), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9944) );
  INV_X1 U11714 ( .A(n9946), .ZN(n9945) );
  NAND2_X1 U11715 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n9946) );
  INV_X1 U11716 ( .A(n14672), .ZN(n10000) );
  NAND2_X1 U11717 ( .A1(n9845), .A2(n9629), .ZN(n9843) );
  NAND2_X1 U11718 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n9988) );
  OR2_X1 U11719 ( .A1(n14718), .A2(n13905), .ZN(n13923) );
  INV_X1 U11720 ( .A(n14729), .ZN(n9998) );
  AND2_X1 U11721 ( .A1(n15019), .A2(n12404), .ZN(n9999) );
  INV_X1 U11722 ( .A(n15386), .ZN(n9840) );
  NAND2_X1 U11723 ( .A1(n9980), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9979) );
  INV_X1 U11724 ( .A(n9981), .ZN(n9980) );
  AND2_X1 U11725 ( .A1(n15247), .A2(n13868), .ZN(n15197) );
  AND2_X1 U11726 ( .A1(n9995), .A2(n9994), .ZN(n9993) );
  INV_X1 U11727 ( .A(n13183), .ZN(n9994) );
  NOR2_X1 U11728 ( .A1(n13172), .A2(n9996), .ZN(n9995) );
  INV_X1 U11729 ( .A(n13070), .ZN(n9996) );
  NAND2_X1 U11730 ( .A1(n10064), .A2(n13995), .ZN(n10063) );
  INV_X1 U11731 ( .A(n13147), .ZN(n10064) );
  OR2_X1 U11732 ( .A1(n10060), .A2(n10059), .ZN(n10058) );
  INV_X1 U11733 ( .A(n15504), .ZN(n10059) );
  OAI21_X1 U11734 ( .B1(n13935), .B2(n13688), .A(n13687), .ZN(n13689) );
  INV_X1 U11735 ( .A(n13937), .ZN(n13935) );
  INV_X1 U11736 ( .A(n18942), .ZN(n9830) );
  AND2_X1 U11737 ( .A1(n13490), .A2(n13488), .ZN(n9836) );
  NOR2_X1 U11738 ( .A1(n13086), .A2(n13085), .ZN(n13480) );
  NAND2_X1 U11739 ( .A1(n12067), .A2(n12066), .ZN(n12074) );
  INV_X1 U11740 ( .A(n13082), .ZN(n10070) );
  NAND2_X1 U11741 ( .A1(n12820), .A2(n12819), .ZN(n12821) );
  AND2_X1 U11742 ( .A1(n12019), .A2(n12018), .ZN(n12575) );
  INV_X1 U11743 ( .A(n11813), .ZN(n9755) );
  NAND2_X1 U11744 ( .A1(n12782), .A2(n12781), .ZN(n12784) );
  NAND2_X1 U11745 ( .A1(n13269), .A2(n12823), .ZN(n12782) );
  NAND2_X1 U11746 ( .A1(n12784), .A2(n12783), .ZN(n12834) );
  INV_X1 U11747 ( .A(n13259), .ZN(n13286) );
  NOR2_X1 U11748 ( .A1(n13269), .A2(n13248), .ZN(n13264) );
  NAND2_X1 U11749 ( .A1(n11718), .A2(n11717), .ZN(n11766) );
  NAND3_X1 U11750 ( .A1(n19812), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19604), 
        .ZN(n13239) );
  OR2_X1 U11751 ( .A1(n9911), .A2(n18560), .ZN(n9647) );
  INV_X1 U11752 ( .A(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n20912) );
  AOI22_X1 U11753 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n17021), .ZN(n9904) );
  NAND2_X1 U11754 ( .A1(n9908), .A2(n9907), .ZN(n9906) );
  INV_X1 U11755 ( .A(n10767), .ZN(n9908) );
  NAND2_X1 U11756 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n9907) );
  OAI211_X1 U11757 ( .C1(n18107), .C2(n9645), .A(n9792), .B(n9791), .ZN(n10767) );
  NOR2_X1 U11758 ( .A1(n18724), .A2(n10726), .ZN(n10809) );
  OR2_X1 U11759 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n13810), .ZN(
        n10726) );
  NAND2_X1 U11760 ( .A1(n17477), .A2(n17507), .ZN(n17508) );
  OAI21_X1 U11761 ( .B1(n10829), .B2(n16339), .A(n17677), .ZN(n10830) );
  INV_X1 U11762 ( .A(n10828), .ZN(n9777) );
  XNOR2_X1 U11763 ( .A(n11000), .B(n9902), .ZN(n10816) );
  NAND2_X1 U11764 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n10724), .ZN(
        n10732) );
  OR2_X1 U11765 ( .A1(n9750), .A2(n10889), .ZN(n10937) );
  NAND2_X1 U11766 ( .A1(n9752), .A2(n9660), .ZN(n9750) );
  OR2_X1 U11767 ( .A1(n10727), .A2(n13810), .ZN(n16940) );
  NAND2_X1 U11768 ( .A1(n14082), .A2(n10092), .ZN(n10094) );
  NOR2_X1 U11769 ( .A1(n14074), .A2(n10093), .ZN(n10092) );
  INV_X1 U11770 ( .A(n14083), .ZN(n10093) );
  AND2_X1 U11771 ( .A1(n14357), .A2(n11552), .ZN(n11553) );
  NAND2_X1 U11772 ( .A1(n11467), .A2(n11466), .ZN(n11502) );
  INV_X1 U11773 ( .A(n11465), .ZN(n11467) );
  AND2_X1 U11774 ( .A1(n14414), .A2(n11552), .ZN(n11426) );
  NAND2_X1 U11775 ( .A1(n11404), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11406) );
  INV_X1 U11776 ( .A(n11403), .ZN(n11404) );
  OR2_X1 U11777 ( .A1(n14419), .A2(n13444), .ZN(n11408) );
  AND2_X1 U11778 ( .A1(n14226), .A2(n9681), .ZN(n14150) );
  AND2_X1 U11779 ( .A1(n11358), .A2(n11357), .ZN(n14218) );
  OR2_X1 U11780 ( .A1(n15862), .A2(n13444), .ZN(n11357) );
  AND2_X1 U11781 ( .A1(n14226), .A2(n14227), .ZN(n14217) );
  AND2_X1 U11782 ( .A1(n11315), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11316) );
  AND2_X1 U11783 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n11316), .ZN(
        n11353) );
  NAND2_X1 U11784 ( .A1(n9740), .A2(n11299), .ZN(n14236) );
  INV_X1 U11785 ( .A(n14241), .ZN(n11299) );
  OR2_X1 U11786 ( .A1(n15952), .A2(n13444), .ZN(n11321) );
  CLKBUF_X1 U11787 ( .A(n14239), .Z(n14240) );
  NAND2_X1 U11788 ( .A1(n11268), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11281) );
  AND2_X1 U11789 ( .A1(n11250), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11268) );
  INV_X1 U11790 ( .A(n13742), .ZN(n9733) );
  NAND2_X1 U11791 ( .A1(n13741), .A2(n11249), .ZN(n13800) );
  INV_X1 U11792 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n20864) );
  AND2_X1 U11793 ( .A1(n11172), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11173) );
  NOR2_X1 U11794 ( .A1(n11167), .A2(n19906), .ZN(n11172) );
  AND3_X1 U11795 ( .A1(n11139), .A2(n11138), .A3(n11137), .ZN(n13414) );
  NOR2_X1 U11796 ( .A1(n11119), .A2(n11123), .ZN(n11141) );
  INV_X1 U11797 ( .A(n9738), .ZN(n13207) );
  AND2_X1 U11798 ( .A1(n11101), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11105) );
  NAND2_X1 U11799 ( .A1(n9739), .A2(n11100), .ZN(n13167) );
  INV_X1 U11800 ( .A(n13156), .ZN(n11100) );
  INV_X1 U11801 ( .A(n13155), .ZN(n9739) );
  AOI21_X1 U11802 ( .B1(n11113), .B2(n11241), .A(n11112), .ZN(n13166) );
  INV_X1 U11803 ( .A(n9851), .ZN(n11113) );
  NAND2_X1 U11804 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11080) );
  NAND2_X1 U11805 ( .A1(n12841), .A2(n11078), .ZN(n13099) );
  OAI21_X1 U11806 ( .B1(n12984), .B2(n10484), .A(n10373), .ZN(n12937) );
  NAND2_X1 U11807 ( .A1(n10096), .A2(n11077), .ZN(n12841) );
  NOR2_X1 U11808 ( .A1(n10510), .A2(n14499), .ZN(n9854) );
  INV_X1 U11809 ( .A(n10511), .ZN(n9855) );
  INV_X1 U11810 ( .A(n14506), .ZN(n10045) );
  AND2_X1 U11811 ( .A1(n14136), .A2(n9705), .ZN(n14091) );
  INV_X1 U11812 ( .A(n14092), .ZN(n9892) );
  NAND2_X1 U11813 ( .A1(n14136), .A2(n9643), .ZN(n14103) );
  NAND2_X1 U11814 ( .A1(n14136), .A2(n14129), .ZN(n14128) );
  NOR2_X1 U11815 ( .A1(n14148), .A2(n14137), .ZN(n14136) );
  INV_X1 U11816 ( .A(n10039), .ZN(n10035) );
  NAND2_X1 U11817 ( .A1(n14450), .A2(n10036), .ZN(n9826) );
  OAI21_X1 U11818 ( .B1(n9611), .B2(n14572), .A(n10040), .ZN(n10039) );
  NAND2_X1 U11819 ( .A1(n9890), .A2(n9889), .ZN(n9888) );
  INV_X1 U11820 ( .A(n14220), .ZN(n9889) );
  INV_X1 U11821 ( .A(n9891), .ZN(n9890) );
  NOR3_X1 U11822 ( .A1(n14250), .A2(n14242), .A3(n10648), .ZN(n14234) );
  NOR2_X1 U11823 ( .A1(n14250), .A2(n14242), .ZN(n14243) );
  AND2_X1 U11824 ( .A1(n9638), .A2(n14182), .ZN(n9894) );
  NAND2_X1 U11825 ( .A1(n13797), .A2(n9676), .ZN(n13804) );
  NAND2_X1 U11826 ( .A1(n13797), .A2(n10632), .ZN(n13754) );
  AND2_X1 U11827 ( .A1(n13735), .A2(n13736), .ZN(n13797) );
  NOR2_X1 U11828 ( .A1(n13521), .A2(n13520), .ZN(n13735) );
  NAND2_X1 U11829 ( .A1(n10053), .A2(n10052), .ZN(n15979) );
  OR2_X1 U11830 ( .A1(n13470), .A2(n13469), .ZN(n13521) );
  OR2_X1 U11831 ( .A1(n13417), .A2(n13416), .ZN(n13470) );
  NOR2_X1 U11832 ( .A1(n10608), .A2(n10607), .ZN(n14257) );
  INV_X1 U11833 ( .A(n10423), .ZN(n10034) );
  NAND2_X1 U11834 ( .A1(n12843), .A2(n9897), .ZN(n14258) );
  AND2_X1 U11835 ( .A1(n9899), .A2(n9672), .ZN(n9897) );
  INV_X1 U11836 ( .A(n13170), .ZN(n9901) );
  NAND2_X1 U11837 ( .A1(n12843), .A2(n9898), .ZN(n13178) );
  AND2_X1 U11838 ( .A1(n9899), .A2(n13179), .ZN(n9898) );
  AND2_X1 U11839 ( .A1(n12843), .A2(n9899), .ZN(n13180) );
  NAND2_X1 U11840 ( .A1(n12843), .A2(n12842), .ZN(n13101) );
  XNOR2_X1 U11841 ( .A(n10401), .B(n20052), .ZN(n13160) );
  NAND2_X1 U11842 ( .A1(n13160), .A2(n13159), .ZN(n13158) );
  AND2_X1 U11843 ( .A1(n12812), .A2(n12810), .ZN(n20034) );
  AND2_X1 U11844 ( .A1(n10706), .A2(n14624), .ZN(n20033) );
  NAND2_X1 U11845 ( .A1(n10705), .A2(n12638), .ZN(n20056) );
  AND2_X1 U11846 ( .A1(n20034), .A2(n20056), .ZN(n16009) );
  AND2_X1 U11847 ( .A1(n10593), .A2(n10592), .ZN(n12768) );
  AND2_X1 U11848 ( .A1(n20652), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11556) );
  CLKBUF_X1 U11849 ( .A(n10300), .Z(n12958) );
  NAND2_X1 U11850 ( .A1(n12624), .A2(n12631), .ZN(n9728) );
  INV_X1 U11851 ( .A(n10338), .ZN(n9821) );
  OR2_X1 U11852 ( .A1(n13379), .A2(n13378), .ZN(n20180) );
  OR2_X1 U11853 ( .A1(n12986), .A2(n20510), .ZN(n20372) );
  AOI221_X1 U11854 ( .B1(n20760), .B2(n14657), .C1(n16122), .C2(n14657), .A(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n20117) );
  AND2_X1 U11855 ( .A1(n12986), .A2(n20739), .ZN(n20312) );
  AND2_X1 U11856 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20117), .ZN(n20104) );
  INV_X1 U11857 ( .A(n20117), .ZN(n20224) );
  NAND2_X1 U11858 ( .A1(n11765), .A2(n19860), .ZN(n11931) );
  OR2_X1 U11859 ( .A1(n12374), .A2(n9927), .ZN(n9922) );
  NAND2_X1 U11860 ( .A1(n9922), .A2(n9921), .ZN(n9920) );
  INV_X1 U11861 ( .A(n15144), .ZN(n9921) );
  NOR2_X1 U11862 ( .A1(n13818), .A2(n12376), .ZN(n13926) );
  OR2_X1 U11863 ( .A1(n9927), .A2(n9928), .ZN(n9926) );
  OR2_X1 U11864 ( .A1(n14733), .A2(n9927), .ZN(n9925) );
  AND2_X1 U11866 ( .A1(n9929), .A2(n9928), .ZN(n14712) );
  INV_X1 U11867 ( .A(n9929), .ZN(n14713) );
  NAND2_X1 U11868 ( .A1(n9868), .A2(n9866), .ZN(n13914) );
  OR2_X1 U11869 ( .A1(n12390), .A2(n9702), .ZN(n9868) );
  AND2_X1 U11870 ( .A1(n13870), .A2(n9871), .ZN(n13856) );
  NAND2_X1 U11871 ( .A1(n13870), .A2(n13869), .ZN(n13872) );
  AND2_X1 U11872 ( .A1(n13840), .A2(n9875), .ZN(n13879) );
  NAND2_X1 U11873 ( .A1(n13847), .A2(n13917), .ZN(n13840) );
  OR2_X1 U11874 ( .A1(n13570), .A2(n9882), .ZN(n13824) );
  AND2_X1 U11875 ( .A1(n13480), .A2(n13479), .ZN(n13572) );
  NAND2_X1 U11876 ( .A1(n13572), .A2(n13571), .ZN(n13570) );
  CLKBUF_X1 U11877 ( .A(n12434), .Z(n19050) );
  INV_X1 U11878 ( .A(n10066), .ZN(n12583) );
  CLKBUF_X1 U11879 ( .A(n11931), .Z(n12581) );
  AND2_X1 U11880 ( .A1(n13187), .A2(n13186), .ZN(n13213) );
  AND2_X1 U11881 ( .A1(n13076), .A2(n13074), .ZN(n13186) );
  AND2_X1 U11882 ( .A1(n13061), .A2(n13060), .ZN(n13074) );
  NOR2_X1 U11884 ( .A1(n19865), .A2(n13826), .ZN(n11933) );
  NOR2_X1 U11885 ( .A1(n14684), .A2(n12296), .ZN(n14030) );
  NOR2_X1 U11886 ( .A1(n14987), .A2(n9954), .ZN(n9953) );
  INV_X1 U11887 ( .A(n14992), .ZN(n9954) );
  NAND2_X1 U11888 ( .A1(n15100), .A2(n9699), .ZN(n14700) );
  AND2_X1 U11889 ( .A1(n15100), .A2(n14726), .ZN(n14724) );
  AND2_X1 U11890 ( .A1(n15448), .A2(n9703), .ZN(n15389) );
  NAND2_X1 U11891 ( .A1(n15043), .A2(n9697), .ZN(n15035) );
  NAND2_X1 U11892 ( .A1(n15448), .A2(n9696), .ZN(n15424) );
  NAND2_X1 U11893 ( .A1(n15448), .A2(n15118), .ZN(n15422) );
  AND2_X1 U11894 ( .A1(n15043), .A2(n14844), .ZN(n15046) );
  AND2_X1 U11895 ( .A1(n12276), .A2(n12275), .ZN(n15449) );
  NOR2_X1 U11896 ( .A1(n15450), .A2(n15449), .ZN(n15448) );
  OR2_X1 U11897 ( .A1(n13146), .A2(n10063), .ZN(n15530) );
  NAND2_X1 U11898 ( .A1(n10065), .A2(n11994), .ZN(n12697) );
  NAND2_X1 U11899 ( .A1(n10066), .A2(n11991), .ZN(n10065) );
  AND2_X1 U11900 ( .A1(n12697), .A2(n12696), .ZN(n12699) );
  INV_X1 U11901 ( .A(n19864), .ZN(n19055) );
  AND2_X1 U11902 ( .A1(n16271), .A2(n19708), .ZN(n12435) );
  INV_X1 U11903 ( .A(n12370), .ZN(n15064) );
  AND2_X1 U11904 ( .A1(n11583), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11601) );
  NOR2_X1 U11905 ( .A1(n11605), .A2(n15206), .ZN(n11603) );
  OR2_X1 U11906 ( .A1(n9974), .A2(n9964), .ZN(n9963) );
  NAND2_X1 U11907 ( .A1(n13940), .A2(n9966), .ZN(n9965) );
  NAND2_X1 U11908 ( .A1(n11612), .A2(n11581), .ZN(n11629) );
  AND2_X1 U11909 ( .A1(n13069), .A2(n9993), .ZN(n13220) );
  NAND2_X1 U11910 ( .A1(n9991), .A2(n9628), .ZN(n13063) );
  OR2_X1 U11911 ( .A1(n11617), .A2(n9942), .ZN(n11621) );
  NAND2_X1 U11912 ( .A1(n9943), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9942) );
  INV_X1 U11913 ( .A(n9944), .ZN(n9943) );
  NOR2_X1 U11914 ( .A1(n11617), .A2(n9944), .ZN(n11622) );
  OR2_X1 U11915 ( .A1(n11617), .A2(n9946), .ZN(n11619) );
  NOR2_X1 U11916 ( .A1(n11617), .A2(n20876), .ZN(n11620) );
  NOR2_X1 U11917 ( .A1(n13034), .A2(n13035), .ZN(n13033) );
  AND2_X1 U11918 ( .A1(n12821), .A2(n11845), .ZN(n13009) );
  NAND2_X1 U11919 ( .A1(n13009), .A2(n13008), .ZN(n13034) );
  NAND2_X1 U11920 ( .A1(n11616), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11615) );
  NOR2_X1 U11921 ( .A1(n11615), .A2(n19128), .ZN(n11618) );
  AND2_X1 U11922 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11616) );
  NOR2_X1 U11923 ( .A1(n15298), .A2(n9988), .ZN(n9987) );
  OR3_X1 U11924 ( .A1(n13931), .A2(n13905), .A3(n9989), .ZN(n14007) );
  AND2_X1 U11925 ( .A1(n15100), .A2(n9706), .ZN(n14679) );
  INV_X1 U11926 ( .A(n12380), .ZN(n10077) );
  AND2_X1 U11927 ( .A1(n9721), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9815) );
  INV_X1 U11928 ( .A(n9979), .ZN(n9978) );
  NAND2_X1 U11929 ( .A1(n15027), .A2(n9698), .ZN(n14727) );
  INV_X1 U11930 ( .A(n10018), .ZN(n10010) );
  NAND2_X1 U11931 ( .A1(n13950), .A2(n9815), .ZN(n15180) );
  NAND2_X1 U11932 ( .A1(n15027), .A2(n9999), .ZN(n15018) );
  AND2_X1 U11933 ( .A1(n15027), .A2(n12404), .ZN(n15020) );
  NOR2_X1 U11934 ( .A1(n15219), .A2(n9979), .ZN(n15184) );
  NOR2_X1 U11935 ( .A1(n9648), .A2(n15028), .ZN(n15027) );
  NAND2_X1 U11936 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n9981) );
  AND2_X1 U11937 ( .A1(n10003), .A2(n10002), .ZN(n10001) );
  INV_X1 U11938 ( .A(n15057), .ZN(n10002) );
  NAND2_X1 U11939 ( .A1(n13950), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15219) );
  NAND2_X1 U11940 ( .A1(n13628), .A2(n10003), .ZN(n15056) );
  NAND2_X1 U11941 ( .A1(n16237), .A2(n10074), .ZN(n15450) );
  AND2_X1 U11942 ( .A1(n10076), .A2(n10075), .ZN(n10074) );
  INV_X1 U11943 ( .A(n15125), .ZN(n10075) );
  OR2_X1 U11944 ( .A1(n13867), .A2(n15786), .ZN(n15247) );
  INV_X1 U11945 ( .A(n15197), .ZN(n15783) );
  AND2_X1 U11946 ( .A1(n16237), .A2(n16221), .ZN(n15777) );
  NAND2_X1 U11947 ( .A1(n13849), .A2(n15492), .ZN(n10026) );
  AOI21_X1 U11948 ( .B1(n9835), .B2(n13845), .A(n13850), .ZN(n9833) );
  AND2_X1 U11949 ( .A1(n12216), .A2(n12215), .ZN(n15495) );
  INV_X1 U11950 ( .A(n13845), .ZN(n9760) );
  NAND2_X1 U11951 ( .A1(n13069), .A2(n9995), .ZN(n13184) );
  NAND2_X1 U11952 ( .A1(n10062), .A2(n10061), .ZN(n10060) );
  INV_X1 U11953 ( .A(n15531), .ZN(n10062) );
  INV_X1 U11954 ( .A(n10063), .ZN(n10061) );
  NOR2_X1 U11955 ( .A1(n13063), .A2(n13064), .ZN(n13069) );
  NAND2_X1 U11956 ( .A1(n13069), .A2(n13070), .ZN(n13173) );
  NAND2_X1 U11957 ( .A1(n10024), .A2(n10020), .ZN(n13989) );
  NAND2_X1 U11958 ( .A1(n9969), .A2(n13948), .ZN(n13987) );
  NAND2_X1 U11959 ( .A1(n9976), .A2(n9970), .ZN(n9969) );
  AND2_X1 U11960 ( .A1(n9971), .A2(n15282), .ZN(n9970) );
  INV_X1 U11961 ( .A(n15544), .ZN(n9971) );
  OAI22_X1 U11962 ( .A1(n12927), .A2(n12928), .B1(n13905), .B2(n12270), .ZN(
        n13118) );
  NAND2_X1 U11963 ( .A1(n9991), .A2(n9623), .ZN(n13109) );
  AND2_X1 U11964 ( .A1(n11979), .A2(n11978), .ZN(n13499) );
  NOR2_X1 U11965 ( .A1(n12911), .A2(n10068), .ZN(n13593) );
  NAND2_X1 U11966 ( .A1(n10071), .A2(n10069), .ZN(n10068) );
  NOR2_X1 U11967 ( .A1(n13499), .A2(n10070), .ZN(n10069) );
  INV_X1 U11968 ( .A(n12049), .ZN(n10071) );
  OR2_X1 U11969 ( .A1(n15579), .A2(n12788), .ZN(n12789) );
  NAND2_X1 U11970 ( .A1(n13313), .A2(n12523), .ZN(n16269) );
  NAND2_X1 U11971 ( .A1(n19055), .A2(n19844), .ZN(n12523) );
  AND2_X1 U11972 ( .A1(n13004), .A2(n12832), .ZN(n12837) );
  NAND2_X1 U11973 ( .A1(n12836), .A2(n12837), .ZN(n13006) );
  AND2_X1 U11974 ( .A1(n15621), .A2(n19800), .ZN(n15632) );
  OR2_X1 U11975 ( .A1(n19702), .A2(n15619), .ZN(n15621) );
  INV_X1 U11976 ( .A(n15647), .ZN(n19516) );
  OR2_X1 U11977 ( .A1(n19445), .A2(n13421), .ZN(n19597) );
  OR2_X1 U11978 ( .A1(n19813), .A2(n19824), .ZN(n19568) );
  INV_X1 U11979 ( .A(n19186), .ZN(n19172) );
  NOR2_X2 U11980 ( .A1(n15064), .A2(n13239), .ZN(n19189) );
  NOR2_X2 U11981 ( .A1(n15061), .A2(n13239), .ZN(n19190) );
  NAND2_X1 U11982 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19604), .ZN(n19186) );
  NOR2_X1 U11983 ( .A1(n10976), .A2(n17306), .ZN(n18753) );
  OR2_X1 U11984 ( .A1(n16582), .A2(n16678), .ZN(n9808) );
  INV_X1 U11985 ( .A(n18101), .ZN(n16776) );
  BUF_X1 U11986 ( .A(n17072), .Z(n17090) );
  INV_X1 U11987 ( .A(n10934), .ZN(n18569) );
  NAND2_X1 U11988 ( .A1(n16928), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10803) );
  NAND2_X1 U11989 ( .A1(n17485), .A2(n9636), .ZN(n17417) );
  NOR2_X1 U11990 ( .A1(n17456), .A2(n9806), .ZN(n9805) );
  NAND2_X1 U11991 ( .A1(n17485), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17455) );
  NAND2_X1 U11992 ( .A1(n17517), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17498) );
  NAND2_X1 U11993 ( .A1(n17592), .A2(n9637), .ZN(n17533) );
  NOR2_X1 U11994 ( .A1(n17569), .A2(n9797), .ZN(n9796) );
  INV_X1 U11995 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n9797) );
  NAND2_X1 U11996 ( .A1(n17592), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17568) );
  NOR2_X1 U11997 ( .A1(n17636), .A2(n17614), .ZN(n17592) );
  AOI21_X1 U11998 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n12345), .A(
        n18478), .ZN(n17613) );
  INV_X1 U11999 ( .A(n17925), .ZN(n17618) );
  NOR2_X1 U12000 ( .A1(n17700), .A2(n17707), .ZN(n17672) );
  NOR2_X1 U12001 ( .A1(n9767), .A2(n9726), .ZN(n9766) );
  NAND2_X1 U12002 ( .A1(n10851), .A2(n11044), .ZN(n9764) );
  NOR2_X1 U12003 ( .A1(n17677), .A2(n16342), .ZN(n16345) );
  NOR2_X1 U12004 ( .A1(n17774), .A2(n17449), .ZN(n17778) );
  OR2_X1 U12005 ( .A1(n17467), .A2(n17808), .ZN(n17449) );
  NOR2_X1 U12006 ( .A1(n17891), .A2(n11031), .ZN(n17811) );
  NAND2_X1 U12007 ( .A1(n17492), .A2(n10973), .ZN(n10845) );
  NOR2_X1 U12008 ( .A1(n17466), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17465) );
  AND3_X1 U12009 ( .A1(n10841), .A2(n10843), .A3(n10840), .ZN(n17560) );
  NAND2_X1 U12010 ( .A1(n17560), .A2(n20867), .ZN(n17559) );
  NAND2_X1 U12011 ( .A1(n17598), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17891) );
  INV_X1 U12012 ( .A(n17600), .ZN(n17585) );
  NOR2_X1 U12013 ( .A1(n17602), .A2(n17601), .ZN(n17600) );
  NOR2_X1 U12014 ( .A1(n17606), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17590) );
  NOR2_X1 U12015 ( .A1(n17676), .A2(n10832), .ZN(n17607) );
  INV_X1 U12016 ( .A(n10837), .ZN(n10832) );
  NOR2_X1 U12017 ( .A1(n11030), .A2(n17674), .ZN(n17954) );
  NAND2_X1 U12018 ( .A1(n10839), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17952) );
  OR2_X1 U12019 ( .A1(n10830), .A2(n9777), .ZN(n9776) );
  NAND2_X1 U12020 ( .A1(n9917), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9916) );
  NAND2_X1 U12021 ( .A1(n10825), .A2(n9917), .ZN(n9915) );
  INV_X1 U12022 ( .A(n17699), .ZN(n9917) );
  NOR2_X1 U12023 ( .A1(n17712), .A2(n18016), .ZN(n17711) );
  XNOR2_X1 U12024 ( .A(n9910), .B(n9909), .ZN(n17737) );
  INV_X1 U12025 ( .A(n10818), .ZN(n9909) );
  NOR2_X1 U12026 ( .A1(n17756), .A2(n10814), .ZN(n17748) );
  INV_X1 U12027 ( .A(n17988), .ZN(n18053) );
  XNOR2_X1 U12028 ( .A(n10815), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17757) );
  NOR2_X1 U12029 ( .A1(n17757), .A2(n17762), .ZN(n17756) );
  NOR2_X1 U12030 ( .A1(n10992), .A2(n15854), .ZN(n18535) );
  INV_X1 U12031 ( .A(n15759), .ZN(n10992) );
  NAND2_X1 U12032 ( .A1(n17763), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17762) );
  NOR2_X2 U12033 ( .A1(n18764), .A2(n15762), .ZN(n18566) );
  NOR2_X1 U12034 ( .A1(n10873), .A2(n10872), .ZN(n18109) );
  INV_X1 U12035 ( .A(n10937), .ZN(n18119) );
  INV_X1 U12036 ( .A(n17154), .ZN(n18124) );
  NOR2_X1 U12037 ( .A1(n10883), .A2(n10882), .ZN(n18127) );
  INV_X1 U12038 ( .A(n18142), .ZN(n18396) );
  AOI21_X1 U12039 ( .B1(n18530), .B2(n18531), .A(n9683), .ZN(n18539) );
  NOR2_X1 U12040 ( .A1(n9753), .A2(n10987), .ZN(n18593) );
  OR2_X1 U12041 ( .A1(n10995), .A2(n9668), .ZN(n9753) );
  AND2_X1 U12042 ( .A1(n14187), .A2(n13458), .ZN(n19961) );
  NAND2_X1 U12043 ( .A1(n13455), .A2(n15827), .ZN(n19924) );
  AND2_X1 U12044 ( .A1(n14187), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19962) );
  AND2_X1 U12045 ( .A1(n13455), .A2(n13442), .ZN(n19948) );
  INV_X1 U12046 ( .A(n19924), .ZN(n19972) );
  INV_X1 U12047 ( .A(n15924), .ZN(n19967) );
  INV_X1 U12048 ( .A(n19948), .ZN(n19976) );
  NAND2_X1 U12049 ( .A1(n12804), .A2(n12762), .ZN(n12764) );
  INV_X1 U12050 ( .A(n14222), .ZN(n14260) );
  INV_X1 U12051 ( .A(n14285), .ZN(n14340) );
  OR2_X1 U12052 ( .A1(n11576), .A2(n13389), .ZN(n14337) );
  INV_X1 U12053 ( .A(n14337), .ZN(n14346) );
  AND2_X1 U12054 ( .A1(n11575), .A2(n13389), .ZN(n14345) );
  AOI21_X2 U12055 ( .B1(n12803), .B2(n11563), .A(n19878), .ZN(n14353) );
  AND2_X1 U12056 ( .A1(n12795), .A2(n11562), .ZN(n11563) );
  INV_X1 U12057 ( .A(n13772), .ZN(n14352) );
  NOR2_X1 U12058 ( .A1(n19979), .A2(n20009), .ZN(n19999) );
  BUF_X1 U12059 ( .A(n19999), .Z(n20008) );
  XNOR2_X1 U12060 ( .A(n10094), .B(n14057), .ZN(n14360) );
  INV_X1 U12061 ( .A(n14447), .ZN(n15947) );
  NAND2_X1 U12062 ( .A1(n10038), .A2(n14437), .ZN(n14423) );
  OR2_X1 U12063 ( .A1(n14450), .A2(n10507), .ZN(n10038) );
  NAND2_X1 U12064 ( .A1(n10053), .A2(n10491), .ZN(n13653) );
  NAND2_X1 U12065 ( .A1(n16002), .A2(n16001), .ZN(n16000) );
  NAND2_X1 U12066 ( .A1(n20014), .A2(n10423), .ZN(n16002) );
  OR2_X1 U12067 ( .A1(n12810), .A2(n20055), .ZN(n10715) );
  CLKBUF_X1 U12068 ( .A(n12943), .Z(n12944) );
  INV_X1 U12069 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20442) );
  NAND2_X1 U12070 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n12800), .ZN(n14657) );
  INV_X1 U12071 ( .A(n20304), .ZN(n20273) );
  OR2_X1 U12072 ( .A1(n20311), .A2(n20540), .ZN(n20310) );
  INV_X1 U12073 ( .A(n20394), .ZN(n20381) );
  INV_X1 U12074 ( .A(n20631), .ZN(n20430) );
  AND2_X1 U12075 ( .A1(n20080), .A2(n20104), .ZN(n20599) );
  AND2_X1 U12076 ( .A1(n20086), .A2(n20104), .ZN(n20611) );
  AND2_X1 U12077 ( .A1(n13390), .A2(n20104), .ZN(n20617) );
  AND2_X1 U12078 ( .A1(n14320), .A2(n20117), .ZN(n20618) );
  INV_X1 U12079 ( .A(n20629), .ZN(n20642) );
  AND2_X1 U12080 ( .A1(n20648), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15834) );
  NAND2_X1 U12081 ( .A1(n9925), .A2(n9926), .ZN(n14695) );
  AND2_X1 U12082 ( .A1(n13818), .A2(n13817), .ZN(n14704) );
  NAND2_X1 U12083 ( .A1(n13917), .A2(n9658), .ZN(n14718) );
  NAND2_X1 U12084 ( .A1(n13919), .A2(n15010), .ZN(n14719) );
  AND2_X1 U12085 ( .A1(n13921), .A2(n13920), .ZN(n14737) );
  NOR2_X1 U12086 ( .A1(n15170), .A2(n14734), .ZN(n14733) );
  OR2_X1 U12087 ( .A1(n12390), .A2(n9662), .ZN(n13882) );
  NAND2_X1 U12088 ( .A1(n9927), .A2(n15222), .ZN(n9931) );
  AND2_X1 U12089 ( .A1(n18817), .A2(n9935), .ZN(n9934) );
  INV_X1 U12090 ( .A(n18810), .ZN(n9935) );
  NAND2_X1 U12091 ( .A1(n9936), .A2(n18817), .ZN(n18809) );
  NAND2_X1 U12092 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11589) );
  NAND2_X1 U12093 ( .A1(n11588), .A2(n11587), .ZN(n11590) );
  INV_X1 U12094 ( .A(n18957), .ZN(n18955) );
  INV_X1 U12095 ( .A(n18898), .ZN(n18961) );
  NOR2_X1 U12096 ( .A1(n12908), .A2(n9704), .ZN(n12915) );
  INV_X1 U12097 ( .A(n18965), .ZN(n18902) );
  AND2_X1 U12098 ( .A1(n12267), .A2(n12266), .ZN(n13530) );
  OR2_X1 U12099 ( .A1(n12229), .A2(n12228), .ZN(n13216) );
  AND2_X1 U12100 ( .A1(n9952), .A2(n9955), .ZN(n14988) );
  NAND2_X1 U12101 ( .A1(n9956), .A2(n14992), .ZN(n9952) );
  NAND2_X1 U12102 ( .A1(n15014), .A2(n15015), .ZN(n15013) );
  NAND2_X1 U12103 ( .A1(n15023), .A2(n14884), .ZN(n15014) );
  OR2_X1 U12104 ( .A1(n12687), .A2(n12686), .ZN(n12688) );
  NOR2_X1 U12105 ( .A1(n19044), .A2(n19040), .ZN(n19024) );
  INV_X1 U12106 ( .A(n18984), .ZN(n19044) );
  BUF_X1 U12108 ( .A(n19106), .Z(n19858) );
  NOR2_X1 U12109 ( .A1(n19084), .A2(n19858), .ZN(n19114) );
  INV_X1 U12110 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12904) );
  NAND2_X1 U12111 ( .A1(n18776), .A2(n12569), .ZN(n19129) );
  INV_X1 U12112 ( .A(n13269), .ZN(n13276) );
  AND2_X1 U12113 ( .A1(n19129), .A2(n12615), .ZN(n19118) );
  INV_X1 U12114 ( .A(n16192), .ZN(n19124) );
  INV_X1 U12115 ( .A(n19121), .ZN(n16160) );
  XOR2_X1 U12116 ( .A(n14024), .B(n14023), .Z(n14739) );
  OAI211_X1 U12117 ( .C1(n15160), .C2(n9989), .A(n9984), .B(n9983), .ZN(n13972) );
  NAND2_X1 U12118 ( .A1(n9985), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9984) );
  INV_X1 U12119 ( .A(n9987), .ZN(n9985) );
  AND2_X1 U12120 ( .A1(n9815), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9814) );
  XNOR2_X1 U12121 ( .A(n10018), .B(n10017), .ZN(n15176) );
  NAND2_X1 U12122 ( .A1(n10014), .A2(n10012), .ZN(n15177) );
  OAI21_X1 U12123 ( .B1(n15385), .B2(n10016), .A(n15386), .ZN(n15190) );
  NOR2_X1 U12124 ( .A1(n15219), .A2(n9981), .ZN(n16157) );
  NAND2_X1 U12125 ( .A1(n13628), .A2(n13627), .ZN(n13648) );
  NAND2_X1 U12126 ( .A1(n10024), .A2(n13822), .ZN(n15288) );
  NAND2_X1 U12127 ( .A1(n13940), .A2(n13939), .ZN(n15286) );
  OR3_X1 U12128 ( .A1(n19142), .A2(n13359), .A3(n19133), .ZN(n13701) );
  NAND2_X1 U12129 ( .A1(n9813), .A2(n13585), .ZN(n13659) );
  NOR2_X1 U12130 ( .A1(n12911), .A2(n12049), .ZN(n13083) );
  AOI211_X1 U12131 ( .C1(n13269), .C2(n19156), .A(n19139), .B(n19138), .ZN(
        n19140) );
  INV_X1 U12132 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19839) );
  OR2_X1 U12133 ( .A1(n15579), .A2(n12695), .ZN(n19834) );
  INV_X1 U12134 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19828) );
  INV_X1 U12135 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19819) );
  INV_X1 U12136 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16292) );
  XNOR2_X1 U12137 ( .A(n12777), .B(n12786), .ZN(n19814) );
  AOI21_X1 U12138 ( .B1(n13269), .B2(n15614), .A(n15597), .ZN(n16259) );
  INV_X1 U12139 ( .A(n19246), .ZN(n15642) );
  OR2_X1 U12140 ( .A1(n19309), .A2(n19516), .ZN(n19298) );
  INV_X1 U12141 ( .A(n19334), .ZN(n19324) );
  INV_X1 U12142 ( .A(n19363), .ZN(n19349) );
  OR2_X1 U12143 ( .A1(n19386), .A2(n19568), .ZN(n19385) );
  NAND2_X1 U12144 ( .A1(n13430), .A2(n13429), .ZN(n19382) );
  OAI21_X1 U12145 ( .B1(n19439), .B2(n19419), .A(n19604), .ZN(n19441) );
  AND2_X1 U12146 ( .A1(n19451), .A2(n19450), .ZN(n19460) );
  NOR2_X1 U12147 ( .A1(n19565), .A2(n19452), .ZN(n19482) );
  NOR2_X2 U12148 ( .A1(n19597), .A2(n19452), .ZN(n19474) );
  INV_X1 U12149 ( .A(n19541), .ZN(n19562) );
  INV_X1 U12150 ( .A(n19660), .ZN(n19575) );
  INV_X1 U12151 ( .A(n19666), .ZN(n19611) );
  NOR2_X1 U12152 ( .A1(n19597), .A2(n19798), .ZN(n19629) );
  OAI21_X1 U12153 ( .B1(n19608), .B2(n19607), .A(n19606), .ZN(n19636) );
  NOR2_X1 U12154 ( .A1(n19565), .A2(n19568), .ZN(n19634) );
  INV_X1 U12155 ( .A(n19707), .ZN(n19635) );
  INV_X1 U12156 ( .A(n19578), .ZN(n19657) );
  INV_X1 U12157 ( .A(n19614), .ZN(n19663) );
  AND2_X1 U12158 ( .A1(n14935), .A2(n19172), .ZN(n19661) );
  INV_X1 U12159 ( .A(n19547), .ZN(n19669) );
  INV_X1 U12160 ( .A(n19620), .ZN(n19675) );
  INV_X1 U12161 ( .A(n19624), .ZN(n19681) );
  INV_X1 U12162 ( .A(n19628), .ZN(n19687) );
  INV_X1 U12163 ( .A(n19558), .ZN(n19693) );
  NOR2_X2 U12164 ( .A1(n19565), .A2(n19798), .ZN(n19702) );
  INV_X1 U12165 ( .A(n19049), .ZN(n19708) );
  INV_X1 U12166 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n11587) );
  NOR2_X1 U12167 ( .A1(n17301), .A2(n18535), .ZN(n18765) );
  INV_X1 U12168 ( .A(n9804), .ZN(n16493) );
  OAI21_X1 U12169 ( .B1(n16545), .B2(n9794), .A(n9793), .ZN(n12426) );
  NAND2_X1 U12170 ( .A1(n9795), .A2(n17448), .ZN(n9793) );
  NOR2_X1 U12172 ( .A1(n12426), .A2(n12427), .ZN(n16481) );
  INV_X1 U12173 ( .A(n16831), .ZN(n16813) );
  NOR2_X1 U12174 ( .A1(n16545), .A2(n9794), .ZN(n16533) );
  AND2_X1 U12175 ( .A1(n9808), .A2(n17516), .ZN(n16573) );
  INV_X1 U12176 ( .A(n9808), .ZN(n16574) );
  NOR2_X1 U12177 ( .A1(n16678), .A2(n9809), .ZN(n16583) );
  AND2_X1 U12178 ( .A1(n16638), .A2(n17488), .ZN(n9809) );
  NOR2_X1 U12179 ( .A1(n16583), .A2(n17519), .ZN(n16582) );
  NOR2_X1 U12180 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16622), .ZN(n16608) );
  AOI211_X1 U12181 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n15660), .A(n18592), .B(
        n12429), .ZN(n16818) );
  NAND2_X1 U12182 ( .A1(n18592), .A2(n12428), .ZN(n16831) );
  INV_X1 U12183 ( .A(n16830), .ZN(n16841) );
  INV_X1 U12184 ( .A(n16838), .ZN(n16840) );
  NOR2_X1 U12185 ( .A1(n16623), .A2(n16979), .ZN(n16992) );
  NAND2_X1 U12186 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17032), .ZN(n17031) );
  NOR3_X2 U12187 ( .A1(n16801), .A2(n17145), .A3(n17134), .ZN(n17136) );
  NOR2_X1 U12188 ( .A1(n17363), .A2(n17185), .ZN(n17179) );
  NOR2_X1 U12189 ( .A1(n17240), .A2(n17190), .ZN(n17186) );
  NOR3_X1 U12190 ( .A1(n17357), .A2(n17231), .A3(n17203), .ZN(n17191) );
  NOR2_X1 U12191 ( .A1(n17411), .A2(n17236), .ZN(n17232) );
  NOR2_X1 U12192 ( .A1(n10740), .A2(n10739), .ZN(n20927) );
  NOR2_X1 U12193 ( .A1(n10751), .A2(n10750), .ZN(n17285) );
  INV_X1 U12195 ( .A(n20928), .ZN(n17271) );
  INV_X1 U12196 ( .A(n17342), .ZN(n17303) );
  CLKBUF_X1 U12197 ( .A(n17317), .Z(n17339) );
  CLKBUF_X1 U12199 ( .A(n17408), .Z(n17403) );
  BUF_X1 U12200 ( .A(n17398), .Z(n17407) );
  NOR2_X1 U12201 ( .A1(n17417), .A2(n17418), .ZN(n16330) );
  NOR2_X1 U12202 ( .A1(n17775), .A2(n17481), .ZN(n17436) );
  NOR2_X1 U12203 ( .A1(n17498), .A2(n17499), .ZN(n17485) );
  NOR2_X1 U12204 ( .A1(n17827), .A2(n17576), .ZN(n17497) );
  NOR2_X1 U12205 ( .A1(n17533), .A2(n17534), .ZN(n17517) );
  OR2_X1 U12206 ( .A1(n17576), .A2(n17842), .ZN(n17541) );
  NAND2_X1 U12207 ( .A1(n17873), .A2(n17642), .ZN(n17576) );
  NOR2_X1 U12208 ( .A1(n10835), .A2(n17585), .ZN(n17824) );
  INV_X1 U12209 ( .A(n12354), .ZN(n17603) );
  INV_X1 U12210 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17662) );
  INV_X1 U12211 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17727) );
  NAND2_X1 U12212 ( .A1(n17764), .A2(n17671), .ZN(n17758) );
  NAND2_X1 U12213 ( .A1(n9914), .A2(n16342), .ZN(n17429) );
  INV_X1 U12214 ( .A(n9913), .ZN(n9912) );
  NAND2_X1 U12215 ( .A1(n9786), .A2(n9790), .ZN(n17440) );
  INV_X1 U12216 ( .A(n9789), .ZN(n17439) );
  INV_X1 U12217 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18762) );
  NOR2_X1 U12218 ( .A1(n11034), .A2(n18548), .ZN(n17988) );
  NOR2_X2 U12219 ( .A1(n17883), .A2(n15660), .ZN(n18530) );
  AOI21_X1 U12220 ( .B1(n11035), .B2(n11034), .A(n18546), .ZN(n18552) );
  INV_X1 U12221 ( .A(n17982), .ZN(n17998) );
  AND2_X1 U12222 ( .A1(n9783), .A2(n9781), .ZN(n17721) );
  NAND2_X1 U12223 ( .A1(n9782), .A2(n9624), .ZN(n9783) );
  INV_X1 U12224 ( .A(n18079), .ZN(n18083) );
  INV_X1 U12225 ( .A(n18068), .ZN(n18085) );
  INV_X1 U12227 ( .A(n9886), .ZN(n12341) );
  OAI21_X1 U12228 ( .B1(n14375), .B2(n15947), .A(n9734), .ZN(P1_U2971) );
  INV_X1 U12229 ( .A(n9735), .ZN(n9734) );
  OAI21_X1 U12230 ( .B1(n14515), .B2(n20030), .A(n9736), .ZN(n9735) );
  AOI21_X1 U12231 ( .B1(n15976), .B2(n14377), .A(n14376), .ZN(n9736) );
  OAI211_X1 U12232 ( .C1(n14202), .C2(n20038), .A(n9887), .B(n9885), .ZN(
        P1_U3000) );
  NOR3_X1 U12233 ( .A1(n10722), .A2(n12336), .A3(n10721), .ZN(n9887) );
  NAND2_X1 U12234 ( .A1(n9886), .A2(n20063), .ZN(n9885) );
  INV_X1 U12235 ( .A(n12316), .ZN(n12323) );
  OR4_X1 U12236 ( .A1(n12386), .A2(n12385), .A3(n12384), .A4(n12383), .ZN(
        P2_U2827) );
  AOI211_X1 U12237 ( .C1(n19121), .C2(n15318), .A(n13985), .B(n13984), .ZN(
        n13986) );
  AOI21_X1 U12238 ( .B1(n15304), .B2(n16228), .A(n10054), .ZN(n15305) );
  OAI211_X1 U12239 ( .C1(n15301), .C2(n19136), .A(n10056), .B(n10055), .ZN(
        n10054) );
  AOI21_X1 U12240 ( .B1(n15302), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n10057), .ZN(n10056) );
  OAI21_X1 U12241 ( .B1(n19166), .B2(n15320), .A(n15319), .ZN(P2_U3018) );
  AOI21_X1 U12242 ( .B1(n9803), .B2(n16820), .A(n9799), .ZN(n16498) );
  XNOR2_X1 U12243 ( .A(n9804), .B(n16494), .ZN(n9803) );
  NOR2_X1 U12244 ( .A1(n12356), .A2(n12355), .ZN(n12357) );
  NOR2_X1 U12245 ( .A1(n10999), .A2(n12354), .ZN(n12355) );
  OAI211_X1 U12246 ( .C1(n17481), .C2(n9748), .A(n9745), .B(n9744), .ZN(
        P3_U2804) );
  NAND2_X1 U12247 ( .A1(n17786), .A2(n9749), .ZN(n9748) );
  INV_X1 U12248 ( .A(n17446), .ZN(n9744) );
  AOI21_X1 U12249 ( .B1(n17445), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n9746), .ZN(n9745) );
  AOI21_X1 U12250 ( .B1(n11047), .B2(n18071), .A(n11046), .ZN(n11048) );
  AND2_X2 U12251 ( .A1(n11937), .A2(n14757), .ZN(n11963) );
  OAI21_X1 U12252 ( .B1(n17416), .B2(n9723), .A(n17677), .ZN(n9771) );
  NAND2_X1 U12253 ( .A1(n14919), .A2(n14918), .ZN(n9958) );
  OAI211_X1 U12254 ( .C1(n9831), .C2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n9635), .B(n9828), .ZN(n13694) );
  INV_X2 U12255 ( .A(n19872), .ZN(n19780) );
  INV_X1 U12256 ( .A(n10496), .ZN(n10510) );
  BUF_X1 U12257 ( .A(n10230), .Z(n11304) );
  INV_X1 U12258 ( .A(n20080), .ZN(n12946) );
  NAND2_X1 U12259 ( .A1(n13517), .A2(n13733), .ZN(n13732) );
  INV_X1 U12261 ( .A(n11752), .ZN(n14941) );
  AND2_X1 U12262 ( .A1(n9992), .A2(n12925), .ZN(n9623) );
  OR2_X1 U12263 ( .A1(n10819), .A2(n10818), .ZN(n9624) );
  NAND2_X1 U12264 ( .A1(n14226), .A2(n9677), .ZN(n14161) );
  AND2_X1 U12265 ( .A1(n9623), .A2(n9990), .ZN(n9625) );
  OR2_X1 U12266 ( .A1(n13912), .A2(n9840), .ZN(n9626) );
  AND2_X1 U12267 ( .A1(n10012), .A2(n10011), .ZN(n9627) );
  AND2_X1 U12268 ( .A1(n9625), .A2(n13048), .ZN(n9628) );
  NAND2_X1 U12269 ( .A1(n9846), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9629) );
  AND2_X1 U12270 ( .A1(n11581), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9630) );
  AND2_X1 U12271 ( .A1(n9993), .A2(n13219), .ZN(n9631) );
  AND2_X1 U12272 ( .A1(n10041), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9632) );
  BUF_X1 U12273 ( .A(n11765), .Z(n19865) );
  NAND3_X1 U12274 ( .A1(n15200), .A2(n13881), .A3(n15202), .ZN(n9633) );
  AND2_X1 U12275 ( .A1(n9776), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9634) );
  INV_X1 U12276 ( .A(n13698), .ZN(n13905) );
  BUF_X1 U12277 ( .A(n16678), .Z(n9794) );
  AND2_X1 U12278 ( .A1(n11612), .A2(n9692), .ZN(n11604) );
  INV_X1 U12279 ( .A(n15015), .ZN(n9950) );
  OR2_X1 U12280 ( .A1(n18942), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9635) );
  AND3_X1 U12281 ( .A1(n15201), .A2(n13898), .A3(n15214), .ZN(n13899) );
  AND2_X1 U12282 ( .A1(n9805), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9636) );
  AND2_X1 U12283 ( .A1(n9796), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9637) );
  AND2_X1 U12284 ( .A1(n9676), .A2(n9895), .ZN(n9638) );
  AND2_X1 U12285 ( .A1(n9938), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9639) );
  AND2_X1 U12286 ( .A1(n10086), .A2(n10438), .ZN(n9640) );
  AND2_X1 U12287 ( .A1(n10090), .A2(n9733), .ZN(n9641) );
  INV_X1 U12288 ( .A(n10851), .ZN(n9767) );
  AND2_X1 U12289 ( .A1(n14129), .A2(n9893), .ZN(n9642) );
  AND2_X1 U12290 ( .A1(n9642), .A2(n14104), .ZN(n9643) );
  AND2_X1 U12291 ( .A1(n10000), .A2(n12379), .ZN(n9644) );
  NAND2_X2 U12292 ( .A1(n19780), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n19784) );
  INV_X1 U12293 ( .A(n11980), .ZN(n12084) );
  OR2_X2 U12294 ( .A1(n18560), .A2(n13810), .ZN(n9645) );
  INV_X4 U12295 ( .A(n17007), .ZN(n17072) );
  OR3_X1 U12296 ( .A1(n14250), .A2(n14242), .A3(n9888), .ZN(n9646) );
  NAND2_X1 U12297 ( .A1(n9864), .A2(n10050), .ZN(n13774) );
  NAND2_X1 U12298 ( .A1(n13940), .A2(n9962), .ZN(n9976) );
  NAND2_X1 U12299 ( .A1(n11763), .A2(n11762), .ZN(n11765) );
  OR2_X1 U12300 ( .A1(n15042), .A2(n12391), .ZN(n9648) );
  AND2_X2 U12301 ( .A1(n12961), .A2(n14643), .ZN(n10278) );
  NAND2_X1 U12302 ( .A1(n13285), .A2(n13284), .ZN(n13489) );
  NAND2_X1 U12303 ( .A1(n13870), .A2(n9873), .ZN(n9649) );
  INV_X1 U12304 ( .A(n10770), .ZN(n10914) );
  AND2_X1 U12305 ( .A1(n13465), .A2(n13516), .ZN(n13517) );
  NOR2_X1 U12306 ( .A1(n13570), .A2(n12919), .ZN(n12920) );
  NOR2_X1 U12307 ( .A1(n15219), .A2(n15205), .ZN(n9650) );
  NAND2_X1 U12308 ( .A1(n15100), .A2(n10079), .ZN(n14697) );
  INV_X2 U12309 ( .A(n20074), .ZN(n13440) );
  AND4_X1 U12310 ( .A1(n10181), .A2(n10180), .A3(n10179), .A4(n10178), .ZN(
        n9651) );
  AND2_X1 U12311 ( .A1(n13214), .A2(n13407), .ZN(n9652) );
  AND3_X1 U12312 ( .A1(n10163), .A2(n10164), .A3(n10162), .ZN(n9653) );
  AND4_X1 U12313 ( .A1(n10806), .A2(n10805), .A3(n10804), .A4(n10803), .ZN(
        n9654) );
  OR2_X1 U12314 ( .A1(n12758), .A2(n10261), .ZN(n9655) );
  AND3_X1 U12315 ( .A1(n11652), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n11651), .ZN(n9656) );
  AND2_X1 U12316 ( .A1(n10129), .A2(n12961), .ZN(n10175) );
  AND2_X1 U12317 ( .A1(n10449), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9657) );
  INV_X1 U12318 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18724) );
  NAND2_X1 U12319 ( .A1(n9976), .A2(n15282), .ZN(n15543) );
  NAND2_X1 U12320 ( .A1(n14450), .A2(n14449), .ZN(n14432) );
  OR2_X1 U12321 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n14719), .ZN(n9658) );
  NAND2_X1 U12322 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n10821), .ZN(
        n9659) );
  NAND2_X1 U12323 ( .A1(n9836), .A2(n13489), .ZN(n13543) );
  AND3_X1 U12324 ( .A1(n10892), .A2(n10891), .A3(n9751), .ZN(n9660) );
  AND2_X1 U12325 ( .A1(n10830), .A2(n9777), .ZN(n9661) );
  AND3_X1 U12326 ( .A1(n13858), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n19177), .ZN(
        n9662) );
  OAI21_X1 U12327 ( .B1(n11825), .B2(n9754), .A(n11810), .ZN(n11811) );
  INV_X1 U12328 ( .A(n13912), .ZN(n10019) );
  BUF_X1 U12329 ( .A(n11787), .Z(n13826) );
  INV_X1 U12330 ( .A(n13842), .ZN(n9835) );
  OR2_X1 U12331 ( .A1(n13979), .A2(n13978), .ZN(n9663) );
  AND2_X1 U12332 ( .A1(n15980), .A2(n16081), .ZN(n9664) );
  AND2_X1 U12333 ( .A1(n10491), .A2(n9671), .ZN(n10052) );
  OR2_X1 U12334 ( .A1(n18061), .A2(n10816), .ZN(n9665) );
  AND2_X1 U12335 ( .A1(n9912), .A2(n9914), .ZN(n9666) );
  INV_X1 U12336 ( .A(n13396), .ZN(n10244) );
  AND2_X1 U12337 ( .A1(n11800), .A2(n11801), .ZN(n11797) );
  INV_X1 U12338 ( .A(n9811), .ZN(n15242) );
  NAND2_X1 U12339 ( .A1(n15241), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9811) );
  AND2_X1 U12340 ( .A1(n11069), .A2(n11067), .ZN(n10270) );
  INV_X1 U12341 ( .A(n10270), .ZN(n9819) );
  INV_X1 U12342 ( .A(n9845), .ZN(n9844) );
  OAI21_X1 U12343 ( .B1(n9846), .B2(n9722), .A(n10008), .ZN(n9845) );
  AND2_X1 U12344 ( .A1(n10010), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9667) );
  INV_X1 U12345 ( .A(n13260), .ZN(n13224) );
  OAI21_X1 U12347 ( .B1(n10024), .B2(n9835), .A(n9759), .ZN(n15491) );
  NAND2_X1 U12348 ( .A1(n10026), .A2(n10025), .ZN(n15273) );
  OR2_X1 U12349 ( .A1(n17154), .A2(n18101), .ZN(n9668) );
  AND2_X1 U12350 ( .A1(n12790), .A2(n12789), .ZN(n9669) );
  OR2_X1 U12351 ( .A1(n10831), .A2(n10830), .ZN(n9670) );
  OR2_X1 U12352 ( .A1(n9611), .A2(n16081), .ZN(n9671) );
  AND2_X1 U12353 ( .A1(n13179), .A2(n9901), .ZN(n9672) );
  AND2_X1 U12354 ( .A1(n9652), .A2(n9959), .ZN(n9673) );
  OR2_X1 U12355 ( .A1(n17564), .A2(n17655), .ZN(n9674) );
  INV_X1 U12356 ( .A(n15283), .ZN(n9977) );
  AND2_X1 U12357 ( .A1(n13942), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15283) );
  OR2_X1 U12358 ( .A1(n12122), .A2(n12121), .ZN(n13698) );
  NAND2_X1 U12359 ( .A1(n20115), .A2(n10340), .ZN(n12997) );
  XNOR2_X1 U12360 ( .A(n12974), .B(n20218), .ZN(n12956) );
  AND2_X1 U12361 ( .A1(n10705), .A2(n10585), .ZN(n20063) );
  AND2_X1 U12362 ( .A1(n11612), .A2(n9630), .ZN(n11606) );
  OR2_X1 U12363 ( .A1(n10260), .A2(n9728), .ZN(n11561) );
  BUF_X1 U12364 ( .A(n11914), .Z(n11927) );
  NAND2_X1 U12365 ( .A1(n13646), .A2(n13645), .ZN(n13726) );
  NAND2_X1 U12366 ( .A1(n13517), .A2(n10090), .ZN(n13739) );
  NOR2_X1 U12367 ( .A1(n13740), .A2(n10083), .ZN(n14176) );
  NOR2_X1 U12368 ( .A1(n11621), .A2(n11579), .ZN(n11614) );
  AND2_X1 U12369 ( .A1(n14136), .A2(n9642), .ZN(n9675) );
  NAND2_X1 U12370 ( .A1(n17559), .A2(n17677), .ZN(n17477) );
  INV_X1 U12371 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12805) );
  AND2_X1 U12372 ( .A1(n10632), .A2(n9896), .ZN(n9676) );
  AND2_X1 U12373 ( .A1(n14218), .A2(n14227), .ZN(n9677) );
  NAND2_X1 U12374 ( .A1(n13207), .A2(n13206), .ZN(n13205) );
  AND2_X1 U12375 ( .A1(n13628), .A2(n10001), .ZN(n15039) );
  AND2_X1 U12376 ( .A1(n13627), .A2(n10005), .ZN(n9678) );
  AND2_X1 U12377 ( .A1(n13779), .A2(n10495), .ZN(n9679) );
  OR3_X1 U12378 ( .A1(n14250), .A2(n14242), .A3(n9891), .ZN(n9680) );
  AND2_X1 U12379 ( .A1(n9677), .A2(n10089), .ZN(n9681) );
  OAI21_X1 U12380 ( .B1(P1_EBX_REG_1__SCAN_IN), .B2(n10680), .A(n10591), .ZN(
        n10594) );
  NOR2_X1 U12381 ( .A1(n13146), .A2(n13147), .ZN(n9682) );
  NOR2_X1 U12382 ( .A1(n10080), .A2(n20649), .ZN(n9731) );
  AND2_X1 U12383 ( .A1(n15768), .A2(n18533), .ZN(n9683) );
  OR2_X1 U12384 ( .A1(n11974), .A2(n11973), .ZN(n13491) );
  AND2_X1 U12385 ( .A1(n10085), .A2(n11140), .ZN(n9684) );
  INV_X1 U12386 ( .A(n15289), .ZN(n10023) );
  AND2_X1 U12387 ( .A1(n13831), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15289) );
  NAND2_X1 U12388 ( .A1(n13517), .A2(n9641), .ZN(n13740) );
  NAND2_X1 U12389 ( .A1(n13906), .A2(n9982), .ZN(n9685) );
  INV_X1 U12390 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20649) );
  INV_X1 U12391 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9754) );
  INV_X1 U12392 ( .A(n18818), .ZN(n9937) );
  INV_X1 U12393 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n20876) );
  AND2_X1 U12394 ( .A1(n13822), .A2(n10023), .ZN(n9686) );
  AND2_X1 U12395 ( .A1(n9933), .A2(n15222), .ZN(n9687) );
  AND2_X1 U12396 ( .A1(n9875), .A2(n13877), .ZN(n9688) );
  AND2_X1 U12397 ( .A1(n9871), .A2(n12310), .ZN(n9689) );
  NOR2_X1 U12398 ( .A1(n16533), .A2(n17448), .ZN(n9690) );
  AND2_X1 U12399 ( .A1(n13488), .A2(n13491), .ZN(n9691) );
  AND2_X1 U12400 ( .A1(n9941), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9692) );
  NAND2_X1 U12401 ( .A1(n10314), .A2(n10357), .ZN(n9693) );
  AND2_X1 U12402 ( .A1(n10461), .A2(n10460), .ZN(n10462) );
  INV_X1 U12403 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15573) );
  INV_X1 U12405 ( .A(n15050), .ZN(n14743) );
  XOR2_X1 U12406 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n12344), .Z(
        n16678) );
  INV_X1 U12407 ( .A(n9794), .ZN(n9795) );
  INV_X1 U12408 ( .A(n13034), .ZN(n9991) );
  NAND2_X1 U12409 ( .A1(n17632), .A2(n17634), .ZN(n17606) );
  NAND2_X1 U12410 ( .A1(n13215), .A2(n9652), .ZN(n13529) );
  NAND2_X1 U12411 ( .A1(n10832), .A2(n17677), .ZN(n17647) );
  AND2_X1 U12412 ( .A1(n13797), .A2(n9638), .ZN(n9694) );
  AND2_X1 U12413 ( .A1(n11601), .A2(n9938), .ZN(n9695) );
  AND2_X1 U12414 ( .A1(n15118), .A2(n10073), .ZN(n9696) );
  AND2_X1 U12415 ( .A1(n14844), .A2(n15036), .ZN(n9697) );
  AND2_X1 U12416 ( .A1(n9999), .A2(n9998), .ZN(n9698) );
  AND2_X1 U12417 ( .A1(n10079), .A2(n10078), .ZN(n9699) );
  AND2_X1 U12418 ( .A1(n14816), .A2(n14900), .ZN(n9700) );
  AND2_X1 U12419 ( .A1(n9991), .A2(n9625), .ZN(n9701) );
  AND2_X1 U12420 ( .A1(n13916), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n9702) );
  AND2_X1 U12421 ( .A1(n11601), .A2(n9639), .ZN(n11591) );
  AND2_X1 U12422 ( .A1(n9696), .A2(n10072), .ZN(n9703) );
  INV_X1 U12423 ( .A(n13846), .ZN(n9878) );
  INV_X1 U12424 ( .A(n13901), .ZN(n9870) );
  NAND2_X1 U12425 ( .A1(n13215), .A2(n13214), .ZN(n13405) );
  INV_X1 U12426 ( .A(n13905), .ZN(n13929) );
  AND2_X1 U12427 ( .A1(n18902), .A2(n13269), .ZN(n9704) );
  AND2_X1 U12428 ( .A1(n9643), .A2(n9892), .ZN(n9705) );
  AND2_X1 U12429 ( .A1(n9699), .A2(n10077), .ZN(n9706) );
  NOR2_X1 U12430 ( .A1(n17711), .A2(n10825), .ZN(n9707) );
  AND2_X1 U12431 ( .A1(n12901), .A2(n9932), .ZN(n9708) );
  AND2_X1 U12432 ( .A1(n14881), .A2(n14880), .ZN(n9709) );
  AND2_X1 U12433 ( .A1(n9697), .A2(n14875), .ZN(n9710) );
  AND2_X1 U12434 ( .A1(n9639), .A2(n11584), .ZN(n9711) );
  AND2_X1 U12435 ( .A1(n9709), .A2(n10100), .ZN(n9712) );
  AND2_X1 U12436 ( .A1(n9869), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n9713) );
  NOR2_X1 U12437 ( .A1(n13146), .A2(n10060), .ZN(n9714) );
  AND2_X1 U12438 ( .A1(n9698), .A2(n9997), .ZN(n9715) );
  AND2_X1 U12439 ( .A1(n9703), .A2(n15388), .ZN(n9716) );
  AND2_X1 U12440 ( .A1(n9644), .A2(n14021), .ZN(n9717) );
  AND2_X1 U12441 ( .A1(n9936), .A2(n9934), .ZN(n9718) );
  INV_X1 U12442 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9743) );
  INV_X1 U12443 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n9880) );
  INV_X1 U12444 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n9806) );
  AND2_X1 U12445 ( .A1(n17485), .A2(n9805), .ZN(n9719) );
  AND2_X1 U12446 ( .A1(n9957), .A2(n14992), .ZN(n9720) );
  AND2_X1 U12447 ( .A1(n9978), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9721) );
  NAND2_X1 U12448 ( .A1(n15313), .A2(n15323), .ZN(n9722) );
  NAND2_X1 U12449 ( .A1(n16320), .A2(n10849), .ZN(n9723) );
  AND2_X1 U12450 ( .A1(n17592), .A2(n9796), .ZN(n9724) );
  INV_X1 U12451 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n9982) );
  INV_X1 U12452 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n9749) );
  AND2_X1 U12453 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n9725) );
  INV_X1 U12454 ( .A(n14571), .ZN(n10042) );
  INV_X1 U12455 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10017) );
  INV_X1 U12456 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9807) );
  INV_X1 U12457 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13130) );
  INV_X1 U12458 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n9798) );
  INV_X1 U12459 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n9989) );
  AND2_X1 U12460 ( .A1(n18708), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9726) );
  AND2_X1 U12461 ( .A1(n9987), .A2(n9989), .ZN(n9727) );
  NAND4_X1 U12462 ( .A1(n18069), .A2(n18743), .A3(n18608), .A4(n18598), .ZN(
        n16842) );
  AOI22_X2 U12463 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20109), .B1(DATAI_26_), 
        .B2(n13388), .ZN(n20610) );
  AOI22_X2 U12464 ( .A1(DATAI_17_), .A2(n13388), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n20109), .ZN(n20604) );
  AOI22_X2 U12465 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20109), .B1(DATAI_24_), 
        .B2(n13388), .ZN(n20598) );
  AOI22_X2 U12466 ( .A1(DATAI_20_), .A2(n13388), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n20109), .ZN(n20568) );
  AOI22_X2 U12467 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20109), .B1(DATAI_31_), 
        .B2(n13388), .ZN(n20647) );
  AOI22_X2 U12468 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20109), .B1(DATAI_30_), 
        .B2(n13388), .ZN(n20636) );
  OR2_X2 U12469 ( .A1(n14222), .A2(n12765), .ZN(n14254) );
  NAND2_X1 U12470 ( .A1(n12764), .A2(n12763), .ZN(n14222) );
  NOR3_X4 U12471 ( .A1(n18280), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18343) );
  NOR2_X1 U12472 ( .A1(n10260), .A2(n12325), .ZN(n10685) );
  NAND3_X1 U12473 ( .A1(n9730), .A2(n10258), .A3(n9729), .ZN(n9732) );
  OR2_X2 U12474 ( .A1(n9821), .A2(n20182), .ZN(n9820) );
  XNOR2_X2 U12475 ( .A(n9732), .B(n10327), .ZN(n20182) );
  OR2_X2 U12476 ( .A1(n13167), .A2(n11116), .ZN(n9738) );
  AND2_X2 U12477 ( .A1(n14226), .A2(n10088), .ZN(n14134) );
  INV_X1 U12478 ( .A(n14239), .ZN(n9740) );
  XNOR2_X2 U12479 ( .A(n9741), .B(n10369), .ZN(n12984) );
  XNOR2_X2 U12480 ( .A(n10356), .B(n10355), .ZN(n9741) );
  OR2_X2 U12481 ( .A1(n16825), .A2(n13810), .ZN(n15722) );
  NOR2_X2 U12482 ( .A1(n16463), .A2(n18750), .ZN(n17759) );
  AND2_X2 U12483 ( .A1(n9754), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11937) );
  NAND2_X1 U12484 ( .A1(n11813), .A2(n11823), .ZN(n12595) );
  OAI21_X2 U12485 ( .B1(n9755), .B2(n12610), .A(n11823), .ZN(n9810) );
  NAND2_X4 U12486 ( .A1(n12552), .A2(n9756), .ZN(n13269) );
  NAND2_X1 U12487 ( .A1(n15840), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9763) );
  NAND3_X1 U12488 ( .A1(n10850), .A2(n9771), .A3(n9766), .ZN(n9765) );
  NAND3_X1 U12489 ( .A1(n9773), .A2(n9776), .A3(n9772), .ZN(n17693) );
  NAND3_X1 U12490 ( .A1(n9773), .A2(n9634), .A3(n9772), .ZN(n9778) );
  INV_X1 U12491 ( .A(n9778), .ZN(n17692) );
  NAND2_X1 U12492 ( .A1(n9659), .A2(n17722), .ZN(n9779) );
  NOR2_X1 U12493 ( .A1(n17737), .A2(n18031), .ZN(n17736) );
  INV_X1 U12494 ( .A(n9783), .ZN(n17723) );
  NAND2_X1 U12495 ( .A1(n17952), .A2(n10837), .ZN(n17994) );
  NAND3_X1 U12496 ( .A1(n9787), .A2(n9789), .A3(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16342) );
  OAI21_X1 U12497 ( .B1(n17452), .B2(n17677), .A(n10847), .ZN(n9788) );
  NAND2_X2 U12498 ( .A1(n18717), .A2(n18554), .ZN(n9911) );
  NAND2_X2 U12499 ( .A1(n9810), .A2(n12551), .ZN(n12552) );
  NAND2_X1 U12500 ( .A1(n15241), .A2(n9725), .ZN(n15218) );
  NOR2_X2 U12501 ( .A1(n15358), .A2(n15336), .ZN(n15160) );
  NAND2_X2 U12502 ( .A1(n9820), .A2(n9817), .ZN(n12974) );
  NAND2_X4 U12503 ( .A1(n9651), .A2(n9622), .ZN(n20105) );
  NAND2_X2 U12504 ( .A1(n9826), .A2(n10035), .ZN(n14417) );
  NAND2_X1 U12505 ( .A1(n11788), .A2(n9827), .ZN(n12558) );
  NAND2_X4 U12506 ( .A1(n12822), .A2(n12821), .ZN(n13271) );
  NOR2_X2 U12507 ( .A1(n13277), .A2(n13269), .ZN(n19197) );
  NAND2_X1 U12508 ( .A1(n13249), .A2(n13275), .ZN(n13277) );
  NAND2_X1 U12509 ( .A1(n9831), .A2(n18942), .ZN(n13695) );
  NAND2_X1 U12510 ( .A1(n13694), .A2(n13693), .ZN(n13697) );
  NAND2_X1 U12511 ( .A1(n9831), .A2(n9829), .ZN(n9828) );
  NOR2_X1 U12512 ( .A1(n9830), .A2(n13597), .ZN(n9829) );
  NAND2_X1 U12513 ( .A1(n9832), .A2(n9833), .ZN(n13849) );
  NAND2_X1 U12514 ( .A1(n9834), .A2(n10024), .ZN(n9832) );
  NAND3_X1 U12515 ( .A1(n13489), .A2(n9691), .A3(n13490), .ZN(n13568) );
  NAND3_X1 U12516 ( .A1(n10026), .A2(n10025), .A3(n13855), .ZN(n15193) );
  NAND2_X1 U12517 ( .A1(n9849), .A2(n10032), .ZN(n9848) );
  INV_X1 U12518 ( .A(n10031), .ZN(n9849) );
  NAND2_X2 U12519 ( .A1(n10394), .A2(n10393), .ZN(n12988) );
  OAI21_X1 U12520 ( .B1(n13606), .B2(n9860), .A(n9856), .ZN(n10037) );
  NAND2_X1 U12521 ( .A1(n9859), .A2(n9857), .ZN(n9856) );
  NAND2_X1 U12522 ( .A1(n9858), .A2(n10041), .ZN(n9857) );
  INV_X1 U12523 ( .A(n10506), .ZN(n9858) );
  NAND4_X1 U12524 ( .A1(n9861), .A2(n9679), .A3(n10050), .A4(n10041), .ZN(
        n9859) );
  AOI21_X1 U12525 ( .B1(n12390), .B2(n9713), .A(n9867), .ZN(n9866) );
  NAND2_X1 U12526 ( .A1(n12390), .A2(n9869), .ZN(n13913) );
  NAND2_X1 U12527 ( .A1(n12390), .A2(n13901), .ZN(n13904) );
  NAND2_X1 U12528 ( .A1(n13870), .A2(n9689), .ZN(n13858) );
  NAND2_X1 U12529 ( .A1(n13840), .A2(n9688), .ZN(n13864) );
  OR2_X1 U12530 ( .A1(n13570), .A2(n9883), .ZN(n13141) );
  INV_X2 U12531 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10120) );
  NAND2_X1 U12532 ( .A1(n13797), .A2(n9894), .ZN(n14248) );
  NAND4_X1 U12533 ( .A1(n10756), .A2(n9904), .A3(n10757), .A4(n10758), .ZN(
        n9903) );
  INV_X2 U12534 ( .A(n10815), .ZN(n11000) );
  INV_X1 U12535 ( .A(n11001), .ZN(n17288) );
  NOR2_X1 U12536 ( .A1(n9911), .A2(n16825), .ZN(n10807) );
  NOR2_X1 U12537 ( .A1(n9911), .A2(n10727), .ZN(n10741) );
  NOR2_X1 U12538 ( .A1(n10837), .A2(n9674), .ZN(n17632) );
  OAI21_X2 U12539 ( .B1(n17712), .B2(n9916), .A(n9915), .ZN(n17698) );
  INV_X1 U12540 ( .A(n9922), .ZN(n14677) );
  INV_X1 U12541 ( .A(n9920), .ZN(n14676) );
  NAND2_X1 U12542 ( .A1(n18817), .A2(n9687), .ZN(n9930) );
  NAND2_X1 U12543 ( .A1(n9931), .A2(n9930), .ZN(n18799) );
  INV_X1 U12544 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9940) );
  OAI21_X1 U12545 ( .B1(n12784), .B2(n12783), .A(n12834), .ZN(n9947) );
  XNOR2_X1 U12546 ( .A(n12833), .B(n9669), .ZN(n19813) );
  AOI21_X2 U12547 ( .B1(n9948), .B2(n15015), .A(n9712), .ZN(n9949) );
  OAI21_X2 U12548 ( .B1(n15023), .B2(n9950), .A(n9949), .ZN(n14893) );
  XNOR2_X2 U12549 ( .A(n14893), .B(n14894), .ZN(n15009) );
  OAI21_X2 U12550 ( .B1(n9955), .B2(n14987), .A(n9951), .ZN(n14986) );
  AND3_X1 U12551 ( .A1(n9958), .A2(n9600), .A3(n9957), .ZN(n14997) );
  NAND2_X1 U12552 ( .A1(n9958), .A2(n9600), .ZN(n14999) );
  INV_X1 U12553 ( .A(n14998), .ZN(n9957) );
  AND2_X2 U12554 ( .A1(n11836), .A2(n11835), .ZN(n12551) );
  INV_X1 U12555 ( .A(n12820), .ZN(n9961) );
  NAND2_X2 U12556 ( .A1(n9961), .A2(n9960), .ZN(n12822) );
  NOR2_X1 U12557 ( .A1(n9968), .A2(n15283), .ZN(n9962) );
  INV_X1 U12558 ( .A(n9972), .ZN(n9964) );
  NOR2_X1 U12559 ( .A1(n9968), .A2(n9967), .ZN(n9966) );
  AND2_X1 U12560 ( .A1(n15160), .A2(n9987), .ZN(n15140) );
  NAND2_X1 U12561 ( .A1(n15160), .A2(n9727), .ZN(n9983) );
  AND2_X1 U12562 ( .A1(n15160), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15148) );
  NAND2_X1 U12563 ( .A1(n15160), .A2(n9986), .ZN(n15141) );
  NAND2_X1 U12564 ( .A1(n13069), .A2(n9631), .ZN(n13218) );
  NAND2_X1 U12565 ( .A1(n14693), .A2(n9644), .ZN(n14675) );
  NAND2_X1 U12566 ( .A1(n14693), .A2(n9717), .ZN(n14023) );
  NAND2_X1 U12567 ( .A1(n14693), .A2(n12379), .ZN(n14673) );
  INV_X1 U12568 ( .A(n14675), .ZN(n14022) );
  OAI22_X1 U12569 ( .A1(n13553), .A2(n13552), .B1(n13551), .B2(n10006), .ZN(
        n13554) );
  AND2_X1 U12570 ( .A1(n13978), .A2(n15323), .ZN(n10009) );
  NAND2_X1 U12571 ( .A1(n10018), .A2(n10017), .ZN(n10011) );
  NAND2_X1 U12572 ( .A1(n15189), .A2(n10015), .ZN(n10013) );
  NAND3_X1 U12573 ( .A1(n13941), .A2(n13905), .A3(n10028), .ZN(n10027) );
  AND2_X1 U12574 ( .A1(n13941), .A2(n10028), .ZN(n13699) );
  NAND2_X1 U12575 ( .A1(n13683), .A2(n13685), .ZN(n10028) );
  OAI21_X1 U12576 ( .B1(n20014), .B2(n10030), .A(n10029), .ZN(n15997) );
  AOI21_X1 U12577 ( .B1(n10034), .B2(n16001), .A(n9657), .ZN(n10029) );
  INV_X1 U12578 ( .A(n16001), .ZN(n10030) );
  OAI21_X1 U12579 ( .B1(n9657), .B2(n16001), .A(n10470), .ZN(n10031) );
  NAND2_X1 U12580 ( .A1(n20014), .A2(n10033), .ZN(n10032) );
  NOR2_X1 U12581 ( .A1(n9657), .A2(n10034), .ZN(n10033) );
  NAND2_X1 U12582 ( .A1(n10037), .A2(n9611), .ZN(n14424) );
  NAND3_X1 U12583 ( .A1(n20115), .A2(n10340), .A3(n20649), .ZN(n10043) );
  NOR2_X1 U12584 ( .A1(n12910), .A2(n12909), .ZN(n12911) );
  NAND2_X1 U12585 ( .A1(n15448), .A2(n9716), .ZN(n15391) );
  NAND3_X2 U12586 ( .A1(n10119), .A2(n9653), .A3(n10165), .ZN(n20098) );
  NAND3_X1 U12587 ( .A1(n13207), .A2(n13206), .A3(n11140), .ZN(n13412) );
  NAND2_X1 U12588 ( .A1(n10439), .A2(n10438), .ZN(n10463) );
  NAND2_X1 U12589 ( .A1(n10439), .A2(n9640), .ZN(n10474) );
  NAND2_X1 U12590 ( .A1(n14082), .A2(n14083), .ZN(n14084) );
  INV_X1 U12591 ( .A(n10094), .ZN(n14072) );
  NAND2_X1 U12592 ( .A1(n13728), .A2(n13727), .ZN(n14830) );
  INV_X1 U12593 ( .A(n13726), .ZN(n13728) );
  NAND2_X1 U12594 ( .A1(n18975), .A2(n19155), .ZN(n14031) );
  OAI21_X1 U12595 ( .B1(n12837), .B2(n12836), .A(n13006), .ZN(n19445) );
  INV_X1 U12596 ( .A(n15218), .ZN(n13950) );
  INV_X1 U12597 ( .A(n13689), .ZN(n13690) );
  OAI21_X1 U12598 ( .B1(n15591), .B2(n11587), .A(n11820), .ZN(n11821) );
  AOI21_X1 U12599 ( .B1(n13340), .B2(n11794), .A(n13344), .ZN(n11795) );
  INV_X1 U12600 ( .A(n13345), .ZN(n15640) );
  AND2_X1 U12601 ( .A1(n11801), .A2(n13345), .ZN(n11720) );
  OAI21_X1 U12602 ( .B1(n12984), .B2(n11170), .A(n11055), .ZN(n11056) );
  NAND2_X1 U12603 ( .A1(n11826), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11832) );
  INV_X1 U12604 ( .A(n15043), .ZN(n15052) );
  AND2_X1 U12605 ( .A1(n16257), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14757) );
  OAI22_X1 U12606 ( .A1(n11739), .A2(n11724), .B1(n16257), .B2(n19819), .ZN(
        n11733) );
  NAND2_X1 U12607 ( .A1(n12343), .A2(n17666), .ZN(n12358) );
  NAND2_X1 U12608 ( .A1(n12343), .A2(n17982), .ZN(n11049) );
  OAI21_X1 U12609 ( .B1(n12626), .B2(n10526), .A(n10683), .ZN(n10247) );
  BUF_X4 U12610 ( .A(n10404), .Z(n11509) );
  NAND2_X1 U12611 ( .A1(n13249), .A2(n13268), .ZN(n13259) );
  INV_X1 U12612 ( .A(n11800), .ZN(n13002) );
  INV_X1 U12613 ( .A(n11792), .ZN(n11801) );
  CLKBUF_X1 U12614 ( .A(n14134), .Z(n14151) );
  NAND2_X1 U12615 ( .A1(n14134), .A2(n14135), .ZN(n14119) );
  NAND2_X1 U12616 ( .A1(n10271), .A2(n9819), .ZN(n20115) );
  AND3_X1 U12617 ( .A1(n13271), .A2(n13268), .A3(n19157), .ZN(n13287) );
  AOI22_X1 U12618 ( .A1(n13594), .A2(n13593), .B1(n11991), .B2(n12107), .ZN(
        n12927) );
  NAND2_X1 U12619 ( .A1(n12974), .A2(n10341), .ZN(n12943) );
  CLKBUF_X1 U12621 ( .A(n14108), .Z(n14120) );
  NAND2_X1 U12622 ( .A1(n14108), .A2(n14110), .ZN(n14095) );
  AND2_X1 U12623 ( .A1(n20098), .A2(n20104), .ZN(n20631) );
  NAND2_X1 U12624 ( .A1(n14072), .A2(n14057), .ZN(n11559) );
  AND2_X1 U12625 ( .A1(n14353), .A2(n12765), .ZN(n10095) );
  NAND2_X1 U12626 ( .A1(n14353), .A2(n12900), .ZN(n14285) );
  AND2_X1 U12627 ( .A1(n11056), .A2(n11078), .ZN(n10096) );
  OR2_X2 U12628 ( .A1(n10734), .A2(n16825), .ZN(n10097) );
  INV_X1 U12629 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10724) );
  AND2_X1 U12630 ( .A1(n18898), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10098) );
  OR2_X1 U12631 ( .A1(n14222), .A2(n20105), .ZN(n14259) );
  AND3_X1 U12632 ( .A1(n11689), .A2(n11688), .A3(n11637), .ZN(n10099) );
  AND2_X1 U12633 ( .A1(n15017), .A2(n14888), .ZN(n10100) );
  NOR3_X1 U12634 ( .A1(n12074), .A2(n12073), .A3(n12072), .ZN(n10101) );
  AND3_X1 U12635 ( .A1(n17939), .A2(n17602), .A3(n10835), .ZN(n10102) );
  NOR2_X1 U12636 ( .A1(n11591), .A2(n11599), .ZN(n10103) );
  INV_X1 U12637 ( .A(n18759), .ZN(n18761) );
  NOR2_X1 U12638 ( .A1(n10727), .A2(n10732), .ZN(n10867) );
  INV_X1 U12639 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19906) );
  AND3_X1 U12640 ( .A1(n13290), .A2(n13289), .A3(n13288), .ZN(n10104) );
  AND2_X1 U12641 ( .A1(n14868), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10105) );
  INV_X1 U12642 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10834) );
  AND2_X1 U12643 ( .A1(n11840), .A2(n11839), .ZN(n10106) );
  AND4_X1 U12644 ( .A1(n10813), .A2(n10812), .A3(n10811), .A4(n10810), .ZN(
        n10107) );
  OR2_X1 U12645 ( .A1(n14337), .A2(n16358), .ZN(n10108) );
  AND3_X1 U12646 ( .A1(n19177), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n13837), .ZN(
        n10109) );
  AND2_X1 U12647 ( .A1(n12772), .A2(n15640), .ZN(n10110) );
  AND2_X1 U12648 ( .A1(n14861), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10111) );
  AND2_X1 U12649 ( .A1(n17142), .A2(n17240), .ZN(n17146) );
  AND2_X1 U12650 ( .A1(n11635), .A2(n11634), .ZN(n10112) );
  INV_X1 U12651 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10849) );
  OR3_X1 U12652 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n17494), .ZN(n10113) );
  INV_X1 U12653 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10835) );
  INV_X1 U12654 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10833) );
  OR2_X1 U12655 ( .A1(n17677), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10114) );
  AND2_X1 U12656 ( .A1(n11577), .A2(n10108), .ZN(n10115) );
  NAND2_X1 U12657 ( .A1(n17610), .A2(n17764), .ZN(n17490) );
  AND2_X1 U12658 ( .A1(n19865), .A2(n13436), .ZN(n10116) );
  INV_X1 U12659 ( .A(n20738), .ZN(n20586) );
  NOR2_X1 U12660 ( .A1(n14027), .A2(n14037), .ZN(n10117) );
  AND3_X1 U12661 ( .A1(n13299), .A2(n13298), .A3(n13297), .ZN(n10118) );
  AND2_X2 U12662 ( .A1(n12961), .A2(n14642), .ZN(n10300) );
  INV_X1 U12663 ( .A(n11118), .ZN(n11400) );
  AND4_X1 U12664 ( .A1(n10169), .A2(n10168), .A3(n10167), .A4(n10166), .ZN(
        n10119) );
  OR2_X1 U12665 ( .A1(n10537), .A2(n10536), .ZN(n10544) );
  AND2_X1 U12666 ( .A1(n16257), .A2(n19819), .ZN(n11724) );
  OR2_X1 U12667 ( .A1(n10435), .A2(n10434), .ZN(n10465) );
  OAI211_X1 U12668 ( .C1(n12635), .C2(n20762), .A(n10698), .B(n10690), .ZN(
        n10266) );
  NAND2_X1 U12669 ( .A1(n14756), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11645) );
  AND4_X1 U12670 ( .A1(n13673), .A2(n13672), .A3(n13671), .A4(n13670), .ZN(
        n13677) );
  AOI22_X1 U12671 ( .A1(n13660), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13299) );
  AOI22_X1 U12672 ( .A1(n10523), .A2(n10522), .B1(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n20395), .ZN(n10517) );
  OR2_X1 U12673 ( .A1(n10415), .A2(n10414), .ZN(n10443) );
  OAI21_X1 U12674 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n10329), .A(
        n10328), .ZN(n10338) );
  AND2_X1 U12675 ( .A1(n11654), .A2(n11653), .ZN(n11655) );
  INV_X1 U12676 ( .A(n12004), .ZN(n12111) );
  INV_X1 U12677 ( .A(n14867), .ZN(n12083) );
  AND2_X1 U12678 ( .A1(n11683), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11687) );
  NOR2_X1 U12679 ( .A1(n10517), .A2(n10518), .ZN(n10516) );
  INV_X1 U12680 ( .A(n11429), .ZN(n11430) );
  NAND3_X1 U12681 ( .A1(n10198), .A2(n10197), .A3(n10264), .ZN(n10260) );
  NOR2_X1 U12682 ( .A1(n11931), .A2(n11587), .ZN(n11778) );
  NAND2_X1 U12683 ( .A1(n13916), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n12302) );
  INV_X1 U12684 ( .A(n14894), .ZN(n14895) );
  NOR2_X1 U12685 ( .A1(n15640), .A2(n11787), .ZN(n11775) );
  AND2_X1 U12686 ( .A1(n11726), .A2(n11725), .ZN(n11735) );
  NAND2_X1 U12687 ( .A1(n12011), .A2(n12010), .ZN(n12012) );
  INV_X1 U12688 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10723) );
  NAND2_X1 U12689 ( .A1(n10244), .A2(n20086), .ZN(n10573) );
  NAND2_X1 U12690 ( .A1(n11430), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11431) );
  AND2_X1 U12691 ( .A1(n11353), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11354) );
  INV_X1 U12692 ( .A(n11051), .ZN(n11118) );
  INV_X1 U12693 ( .A(n10353), .ZN(n10395) );
  AND2_X1 U12694 ( .A1(n10578), .A2(n10689), .ZN(n12796) );
  INV_X1 U12695 ( .A(n10555), .ZN(n10559) );
  AND2_X1 U12696 ( .A1(n11736), .A2(n12304), .ZN(n12555) );
  AND2_X1 U12697 ( .A1(n13004), .A2(n13003), .ZN(n13005) );
  NAND2_X1 U12698 ( .A1(n14893), .A2(n14895), .ZN(n14896) );
  NAND2_X1 U12699 ( .A1(n11761), .A2(n11637), .ZN(n11762) );
  NOR2_X1 U12700 ( .A1(n18124), .A2(n18127), .ZN(n10945) );
  NAND2_X1 U12701 ( .A1(n17564), .A2(n20793), .ZN(n10840) );
  NOR2_X1 U12702 ( .A1(n11022), .A2(n17702), .ZN(n11025) );
  NAND2_X1 U12703 ( .A1(n10380), .A2(n10379), .ZN(n20218) );
  INV_X1 U12704 ( .A(n14152), .ZN(n11410) );
  INV_X1 U12705 ( .A(n11527), .ZN(n11549) );
  OR2_X1 U12706 ( .A1(n11507), .A2(n11506), .ZN(n12334) );
  OR2_X1 U12707 ( .A1(n11431), .A2(n14124), .ZN(n11465) );
  NAND2_X1 U12708 ( .A1(n11354), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11403) );
  AND2_X1 U12709 ( .A1(n20092), .A2(n20080), .ZN(n10530) );
  INV_X1 U12710 ( .A(n10680), .ZN(n10676) );
  NAND2_X1 U12711 ( .A1(n10677), .A2(n10662), .ZN(n10653) );
  NAND3_X1 U12712 ( .A1(n13390), .A2(n20074), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n10555) );
  AND2_X1 U12713 ( .A1(n10700), .A2(n10699), .ZN(n12948) );
  INV_X1 U12714 ( .A(n20146), .ZN(n20184) );
  INV_X1 U12715 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20395) );
  INV_X1 U12716 ( .A(n13917), .ZN(n13918) );
  INV_X1 U12717 ( .A(n15032), .ZN(n14875) );
  INV_X1 U12718 ( .A(n13729), .ZN(n13727) );
  NAND2_X1 U12719 ( .A1(n11729), .A2(n11728), .ZN(n12522) );
  OR2_X1 U12720 ( .A1(n19153), .A2(n19154), .ZN(n15552) );
  NAND2_X1 U12721 ( .A1(n13490), .A2(n13488), .ZN(n13304) );
  NAND2_X1 U12722 ( .A1(n12521), .A2(n12520), .ZN(n13313) );
  INV_X1 U12723 ( .A(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n20794) );
  NOR2_X1 U12724 ( .A1(n11024), .A2(n11028), .ZN(n11030) );
  XOR2_X1 U12725 ( .A(n20927), .B(n10826), .Z(n10827) );
  NOR2_X1 U12726 ( .A1(n10994), .A2(n10983), .ZN(n15658) );
  NOR2_X1 U12727 ( .A1(n11033), .A2(n18546), .ZN(n18542) );
  AND2_X1 U12728 ( .A1(n12639), .A2(n12640), .ZN(n12625) );
  AND2_X1 U12729 ( .A1(n10646), .A2(n10645), .ZN(n14242) );
  NAND2_X1 U12730 ( .A1(n11217), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11232) );
  OR3_X1 U12731 ( .A1(n13448), .A2(n13447), .A3(n13446), .ZN(n14187) );
  AND2_X1 U12732 ( .A1(n10624), .A2(n10623), .ZN(n13520) );
  INV_X1 U12733 ( .A(n12840), .ZN(n11077) );
  INV_X1 U12734 ( .A(n11557), .ZN(n11558) );
  OR2_X1 U12735 ( .A1(n11406), .A2(n11405), .ZN(n11429) );
  NOR2_X1 U12736 ( .A1(n11232), .A2(n15925), .ZN(n11250) );
  NOR2_X1 U12737 ( .A1(n20864), .A2(n11187), .ZN(n11217) );
  NAND2_X1 U12738 ( .A1(n11141), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11167) );
  AOI21_X1 U12739 ( .B1(n11099), .B2(n11241), .A(n11098), .ZN(n13156) );
  OR2_X1 U12740 ( .A1(n20019), .A2(n12331), .ZN(n20024) );
  AND2_X1 U12741 ( .A1(n16009), .A2(n20033), .ZN(n14601) );
  INV_X1 U12742 ( .A(n20587), .ZN(n20396) );
  INV_X1 U12743 ( .A(n20637), .ZN(n20435) );
  NOR2_X1 U12744 ( .A1(n20224), .A2(n20223), .ZN(n20549) );
  INV_X1 U12745 ( .A(n20185), .ZN(n20593) );
  INV_X1 U12746 ( .A(n12522), .ZN(n19844) );
  INV_X1 U12747 ( .A(n18975), .ZN(n14667) );
  NAND2_X1 U12748 ( .A1(n12835), .A2(n12834), .ZN(n12836) );
  INV_X1 U12749 ( .A(n15044), .ZN(n14844) );
  AND2_X1 U12750 ( .A1(n12143), .A2(n12142), .ZN(n13147) );
  AND2_X1 U12751 ( .A1(n12522), .A2(n11741), .ZN(n16271) );
  INV_X1 U12752 ( .A(n12610), .ZN(n12596) );
  AOI21_X1 U12753 ( .B1(n13930), .B2(n13929), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14008) );
  AND2_X1 U12754 ( .A1(n15257), .A2(n15256), .ZN(n15488) );
  INV_X1 U12755 ( .A(n12299), .ZN(n13302) );
  OR2_X1 U12756 ( .A1(n13357), .A2(n13335), .ZN(n16248) );
  NAND2_X1 U12757 ( .A1(n13252), .A2(n12823), .ZN(n12693) );
  OR3_X1 U12758 ( .A1(n19205), .A2(n19389), .A3(n19199), .ZN(n19244) );
  NAND2_X1 U12759 ( .A1(n19813), .A2(n19814), .ZN(n19452) );
  NOR2_X1 U12760 ( .A1(n18109), .A2(n10996), .ZN(n10982) );
  OR2_X1 U12761 ( .A1(n16502), .A2(P3_EBX_REG_29__SCAN_IN), .ZN(n16492) );
  NOR2_X1 U12762 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16698), .ZN(n16681) );
  AOI211_X1 U12763 ( .C1(n17082), .C2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n10909), .B(n10908), .ZN(n10910) );
  NOR2_X1 U12764 ( .A1(n17296), .A2(n17241), .ZN(n17272) );
  OAI21_X1 U12765 ( .B1(n15762), .B2(n15763), .A(n15659), .ZN(n15855) );
  INV_X1 U12766 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16708) );
  INV_X1 U12767 ( .A(n17477), .ZN(n17493) );
  NOR2_X1 U12768 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17564), .ZN(
        n17542) );
  NAND2_X1 U12769 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17618), .ZN(
        n17601) );
  INV_X1 U12770 ( .A(n17677), .ZN(n17564) );
  INV_X1 U12771 ( .A(n18531), .ZN(n15763) );
  INV_X1 U12772 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18575) );
  NAND2_X1 U12773 ( .A1(n10568), .A2(n10567), .ZN(n12800) );
  NOR3_X1 U12774 ( .A1(n19924), .A2(n19913), .A3(n13758), .ZN(n15933) );
  AND2_X1 U12775 ( .A1(n14187), .A2(n13449), .ZN(n19942) );
  INV_X1 U12777 ( .A(n14259), .ZN(n14223) );
  INV_X1 U12778 ( .A(n14353), .ZN(n14342) );
  NOR2_X1 U12779 ( .A1(n14342), .A2(n12900), .ZN(n13772) );
  AND2_X1 U12780 ( .A1(n12800), .A2(n12747), .ZN(n19979) );
  AND2_X1 U12781 ( .A1(n11507), .A2(n11503), .ZN(n14377) );
  INV_X1 U12782 ( .A(n14319), .ZN(n15880) );
  NAND2_X1 U12783 ( .A1(n11173), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11187) );
  NAND2_X1 U12784 ( .A1(n11105), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11119) );
  INV_X1 U12785 ( .A(n20024), .ZN(n20013) );
  AND2_X1 U12786 ( .A1(n20024), .A2(n12333), .ZN(n15976) );
  INV_X1 U12787 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10512) );
  NOR2_X1 U12788 ( .A1(n16054), .A2(n20047), .ZN(n16087) );
  INV_X1 U12789 ( .A(n20038), .ZN(n20059) );
  NAND2_X1 U12790 ( .A1(n10705), .A2(n10684), .ZN(n20038) );
  NOR2_X1 U12791 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19877) );
  INV_X1 U12792 ( .A(n20141), .ZN(n20127) );
  INV_X1 U12793 ( .A(n20177), .ZN(n20143) );
  OAI21_X1 U12794 ( .B1(n20150), .B2(n20148), .A(n20147), .ZN(n20174) );
  OAI21_X1 U12795 ( .B1(n20241), .B2(n20225), .A(n20549), .ZN(n20243) );
  INV_X1 U12796 ( .A(n20271), .ZN(n20261) );
  INV_X1 U12797 ( .A(n20310), .ZN(n20336) );
  OAI211_X1 U12798 ( .C1(n20361), .C2(n20481), .A(n20400), .B(n20346), .ZN(
        n20363) );
  OR2_X1 U12799 ( .A1(n12986), .A2(n20739), .ZN(n20473) );
  INV_X1 U12800 ( .A(n20403), .ZN(n20438) );
  NAND2_X1 U12801 ( .A1(n12986), .A2(n20510), .ZN(n20540) );
  NAND2_X1 U12802 ( .A1(n13379), .A2(n12984), .ZN(n20450) );
  AND2_X1 U12803 ( .A1(n20542), .A2(n20474), .ZN(n20536) );
  INV_X1 U12804 ( .A(n20573), .ZN(n20577) );
  OAI211_X1 U12805 ( .C1(n20574), .C2(n20550), .A(n20549), .B(n20548), .ZN(
        n20578) );
  AND2_X1 U12806 ( .A1(n13396), .A2(n20104), .ZN(n20605) );
  AND2_X1 U12807 ( .A1(n20105), .A2(n20104), .ZN(n20637) );
  INV_X1 U12808 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20648) );
  NOR2_X1 U12809 ( .A1(n18923), .A2(n13951), .ZN(n12321) );
  OR2_X1 U12810 ( .A1(n19051), .A2(n12298), .ZN(n18960) );
  INV_X1 U12811 ( .A(n18960), .ZN(n18907) );
  AND2_X1 U12812 ( .A1(n19855), .A2(n11744), .ZN(n18963) );
  INV_X1 U12813 ( .A(n15060), .ZN(n15047) );
  INV_X1 U12814 ( .A(n19014), .ZN(n19039) );
  INV_X1 U12815 ( .A(n12501), .ZN(n12674) );
  INV_X1 U12816 ( .A(n16194), .ZN(n19123) );
  AND2_X1 U12817 ( .A1(n19129), .A2(n19820), .ZN(n19121) );
  AND2_X1 U12818 ( .A1(n15490), .A2(n15489), .ZN(n16185) );
  INV_X1 U12819 ( .A(n16248), .ZN(n19156) );
  INV_X1 U12820 ( .A(n19650), .ZN(n19604) );
  NAND2_X1 U12821 ( .A1(n16269), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15616) );
  OAI21_X1 U12822 ( .B1(n15632), .B2(n15631), .A(n15630), .ZN(n19191) );
  NOR2_X2 U12823 ( .A1(n19452), .A2(n19309), .ZN(n19246) );
  NOR2_X1 U12824 ( .A1(n19452), .A2(n19386), .ZN(n19272) );
  INV_X1 U12825 ( .A(n19298), .ZN(n19302) );
  INV_X1 U12826 ( .A(n19313), .ZN(n19331) );
  NAND2_X1 U12827 ( .A1(n19445), .A2(n19834), .ZN(n19309) );
  NAND2_X1 U12828 ( .A1(n19424), .A2(n19423), .ZN(n19440) );
  INV_X1 U12829 ( .A(n19460), .ZN(n19476) );
  OAI21_X1 U12830 ( .B1(n19489), .B2(n19488), .A(n19604), .ZN(n19506) );
  NOR2_X2 U12831 ( .A1(n19597), .A2(n19516), .ZN(n19537) );
  AND2_X1 U12832 ( .A1(n19813), .A2(n19824), .ZN(n15647) );
  INV_X1 U12833 ( .A(n19591), .ZN(n19593) );
  INV_X1 U12834 ( .A(n19690), .ZN(n19625) );
  INV_X1 U12835 ( .A(n19260), .ZN(n19679) );
  INV_X1 U12836 ( .A(n18765), .ZN(n18743) );
  AOI21_X1 U12837 ( .B1(n10960), .B2(n10959), .A(n10958), .ZN(n18531) );
  NOR2_X1 U12838 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16598), .ZN(n16584) );
  NOR2_X1 U12839 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16645), .ZN(n16631) );
  NOR2_X1 U12840 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16668), .ZN(n16656) );
  NOR2_X1 U12841 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16722), .ZN(n16704) );
  NOR2_X1 U12842 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16748), .ZN(n16725) );
  INV_X1 U12843 ( .A(n16827), .ZN(n16791) );
  INV_X1 U12844 ( .A(n18750), .ZN(n15660) );
  NOR2_X1 U12845 ( .A1(n15735), .A2(n16923), .ZN(n16905) );
  NAND2_X1 U12846 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16992), .ZN(n16977) );
  NOR2_X1 U12847 ( .A1(n17018), .A2(n17031), .ZN(n17005) );
  INV_X1 U12848 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n16801) );
  NAND4_X1 U12849 ( .A1(n15660), .A2(n16776), .A3(n15855), .A4(n18745), .ZN(
        n17145) );
  NAND2_X1 U12850 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17186), .ZN(n17185) );
  NAND2_X1 U12851 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17232), .ZN(n17231) );
  NAND3_X1 U12852 ( .A1(n10800), .A2(n10799), .A3(n10798), .ZN(n16339) );
  NAND2_X1 U12853 ( .A1(n17151), .A2(n17240), .ZN(n20926) );
  NAND2_X1 U12854 ( .A1(n17151), .A2(P3_EAX_REG_0__SCAN_IN), .ZN(n17296) );
  NOR2_X1 U12855 ( .A1(n18710), .A2(n17758), .ZN(n17532) );
  NAND2_X1 U12856 ( .A1(n10834), .A2(n10833), .ZN(n17655) );
  AOI21_X1 U12857 ( .B1(n17938), .B2(n17937), .A(n18086), .ZN(n17980) );
  INV_X1 U12858 ( .A(n18072), .ZN(n18051) );
  NAND2_X1 U12859 ( .A1(n12414), .A2(n18099), .ZN(n18142) );
  INV_X1 U12860 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18618) );
  NAND2_X1 U12861 ( .A1(n12800), .A2(n12444), .ZN(n12704) );
  INV_X1 U12862 ( .A(n19962), .ZN(n19905) );
  INV_X1 U12863 ( .A(n19942), .ZN(n19928) );
  AND2_X1 U12864 ( .A1(n19928), .A2(n13450), .ZN(n19969) );
  INV_X1 U12865 ( .A(n15992), .ZN(n19929) );
  INV_X1 U12866 ( .A(n19979), .ZN(n20011) );
  AOI21_X1 U12867 ( .B1(n20759), .B2(n20762), .A(n12704), .ZN(n12896) );
  INV_X1 U12868 ( .A(n12338), .ZN(n12339) );
  INV_X1 U12869 ( .A(n15976), .ZN(n20023) );
  INV_X1 U12870 ( .A(n20063), .ZN(n16106) );
  INV_X1 U12871 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20742) );
  INV_X1 U12872 ( .A(n20073), .ZN(n20114) );
  OR2_X1 U12873 ( .A1(n20180), .A2(n20473), .ZN(n20141) );
  OR2_X1 U12874 ( .A1(n20180), .A2(n20372), .ZN(n20177) );
  OR2_X1 U12875 ( .A1(n20180), .A2(n20540), .ZN(n20212) );
  OR2_X1 U12876 ( .A1(n20180), .A2(n20449), .ZN(n20246) );
  OR2_X1 U12877 ( .A1(n20311), .A2(n20473), .ZN(n20271) );
  OR2_X1 U12878 ( .A1(n20311), .A2(n20372), .ZN(n20304) );
  NAND2_X1 U12879 ( .A1(n20313), .A2(n20312), .ZN(n20366) );
  OR2_X1 U12880 ( .A1(n20450), .A2(n20473), .ZN(n20394) );
  OR2_X1 U12881 ( .A1(n20450), .A2(n20372), .ZN(n20441) );
  OR2_X1 U12882 ( .A1(n20450), .A2(n20540), .ZN(n20472) );
  OR2_X1 U12883 ( .A1(n20450), .A2(n20449), .ZN(n20509) );
  OR2_X1 U12884 ( .A1(n20511), .A2(n20510), .ZN(n20573) );
  NAND2_X1 U12885 ( .A1(n20542), .A2(n20541), .ZN(n20646) );
  INV_X1 U12886 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19721) );
  OR2_X1 U12887 ( .A1(n19855), .A2(n11932), .ZN(n18965) );
  INV_X1 U12888 ( .A(n18958), .ZN(n18941) );
  INV_X1 U12889 ( .A(n14743), .ZN(n15055) );
  NAND2_X1 U12890 ( .A1(n12771), .A2(n19708), .ZN(n15050) );
  AND2_X1 U12891 ( .A1(n12688), .A2(n19708), .ZN(n19014) );
  INV_X1 U12892 ( .A(n19008), .ZN(n19048) );
  INV_X1 U12893 ( .A(n19084), .ZN(n19116) );
  NAND2_X1 U12894 ( .A1(n16295), .A2(n12435), .ZN(n19051) );
  INV_X1 U12895 ( .A(n19118), .ZN(n16190) );
  OR2_X1 U12896 ( .A1(n18776), .A2(n14935), .ZN(n16194) );
  OR2_X1 U12897 ( .A1(n13357), .A2(n13332), .ZN(n19136) );
  OR2_X1 U12898 ( .A1(n13357), .A2(n19849), .ZN(n19166) );
  OR2_X1 U12899 ( .A1(n13357), .A2(n19842), .ZN(n19159) );
  AND2_X1 U12900 ( .A1(n15626), .A2(n15625), .ZN(n19195) );
  INV_X1 U12901 ( .A(n19272), .ZN(n19250) );
  NOR2_X1 U12902 ( .A1(n15650), .A2(n19650), .ZN(n19276) );
  OR2_X1 U12903 ( .A1(n19386), .A2(n19516), .ZN(n19334) );
  OR2_X1 U12904 ( .A1(n19309), .A2(n19568), .ZN(n19363) );
  INV_X1 U12905 ( .A(n19382), .ZN(n19371) );
  OR2_X1 U12906 ( .A1(n19798), .A2(n19386), .ZN(n19444) );
  INV_X1 U12907 ( .A(n19474), .ZN(n19473) );
  INV_X1 U12908 ( .A(n19482), .ZN(n19509) );
  NAND2_X1 U12909 ( .A1(n13230), .A2(n15647), .ZN(n19552) );
  NAND2_X1 U12910 ( .A1(n13229), .A2(n13228), .ZN(n19591) );
  INV_X1 U12911 ( .A(n19634), .ZN(n19632) );
  INV_X1 U12912 ( .A(n19629), .ZN(n19706) );
  AND3_X1 U12913 ( .A1(n19721), .A2(n19784), .A3(n19727), .ZN(n19866) );
  INV_X1 U12914 ( .A(n16818), .ZN(n16830) );
  NAND4_X1 U12915 ( .A1(n12428), .A2(P3_EBX_REG_31__SCAN_IN), .A3(n15660), 
        .A4(n12413), .ZN(n16838) );
  NOR2_X1 U12916 ( .A1(n16848), .A2(n16899), .ZN(n16904) );
  NOR2_X1 U12917 ( .A1(n16599), .A2(n16977), .ZN(n16966) );
  NOR2_X1 U12918 ( .A1(n16676), .A2(n15739), .ZN(n17032) );
  NOR2_X1 U12919 ( .A1(n17371), .A2(n17165), .ZN(n17164) );
  NOR2_X1 U12920 ( .A1(n17367), .A2(n17175), .ZN(n17174) );
  OR2_X1 U12921 ( .A1(n17242), .A2(n17261), .ZN(n17260) );
  NOR2_X1 U12922 ( .A1(n17241), .A2(n17281), .ZN(n17279) );
  NOR2_X1 U12923 ( .A1(n18747), .A2(n17303), .ZN(n17317) );
  NAND2_X1 U12924 ( .A1(n17343), .A2(n17302), .ZN(n17342) );
  CLKBUF_X1 U12925 ( .A(n17410), .Z(n17405) );
  INV_X1 U12926 ( .A(n17532), .ZN(n17622) );
  INV_X1 U12927 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17707) );
  OAI21_X2 U12928 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18744), .A(n16463), 
        .ZN(n17764) );
  INV_X1 U12929 ( .A(n18071), .ZN(n18086) );
  INV_X1 U12930 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18004) );
  INV_X1 U12931 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18392) );
  INV_X1 U12932 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18584) );
  INV_X1 U12933 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18107) );
  INV_X1 U12934 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20890) );
  INV_X1 U12935 ( .A(n18163), .ZN(n18528) );
  INV_X1 U12936 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n20828) );
  INV_X1 U12937 ( .A(n18697), .ZN(n18759) );
  NAND2_X1 U12938 ( .A1(n12358), .A2(n12357), .ZN(P3_U2799) );
  NAND2_X1 U12939 ( .A1(n11049), .A2(n11048), .ZN(P3_U2831) );
  AND2_X4 U12940 ( .A1(n10120), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12964) );
  AND2_X4 U12941 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14642) );
  AND2_X4 U12942 ( .A1(n12964), .A2(n14642), .ZN(n10272) );
  NAND2_X1 U12943 ( .A1(n10272), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10124) );
  AND2_X4 U12944 ( .A1(n12964), .A2(n10129), .ZN(n10161) );
  NAND2_X1 U12945 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10123) );
  NOR2_X4 U12946 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14643) );
  NAND2_X1 U12947 ( .A1(n10278), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10122) );
  AND2_X4 U12948 ( .A1(n12964), .A2(n10134), .ZN(n10301) );
  NAND2_X1 U12949 ( .A1(n10301), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10121) );
  NAND2_X1 U12950 ( .A1(n10175), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10128) );
  AND2_X2 U12951 ( .A1(n12964), .A2(n14643), .ZN(n10404) );
  BUF_X2 U12952 ( .A(n10404), .Z(n11474) );
  NAND2_X1 U12953 ( .A1(n11474), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10127) );
  AND2_X2 U12954 ( .A1(n10129), .A2(n10135), .ZN(n10230) );
  NAND2_X1 U12955 ( .A1(n11532), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10126) );
  NAND2_X1 U12956 ( .A1(n10342), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10125) );
  NAND2_X1 U12957 ( .A1(n10223), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10133) );
  AND2_X2 U12958 ( .A1(n10129), .A2(n10136), .ZN(n10224) );
  BUF_X2 U12959 ( .A(n10224), .Z(n11363) );
  NAND2_X1 U12960 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10132) );
  NAND2_X1 U12961 ( .A1(n10300), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10131) );
  NAND2_X1 U12962 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10130) );
  AND2_X2 U12963 ( .A1(n10134), .A2(n10135), .ZN(n10186) );
  NAND2_X1 U12964 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10140) );
  NAND2_X1 U12965 ( .A1(n10273), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10139) );
  NAND2_X1 U12966 ( .A1(n10185), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10138) );
  AND2_X2 U12967 ( .A1(n14643), .A2(n10136), .ZN(n10409) );
  NAND2_X1 U12968 ( .A1(n10409), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10137) );
  AOI22_X1 U12970 ( .A1(n10175), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10230), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10144) );
  AOI22_X1 U12971 ( .A1(n10223), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10143) );
  AOI22_X1 U12972 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10342), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10142) );
  BUF_X2 U12973 ( .A(n10224), .Z(n11487) );
  AOI22_X1 U12974 ( .A1(n11487), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10300), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10141) );
  NAND4_X1 U12975 ( .A1(n10144), .A2(n10143), .A3(n10142), .A4(n10141), .ZN(
        n10150) );
  AOI22_X1 U12976 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10148) );
  AOI22_X1 U12977 ( .A1(n10186), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10409), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10147) );
  AOI22_X1 U12978 ( .A1(n10273), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10185), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10146) );
  AOI22_X1 U12979 ( .A1(n10278), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10301), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10145) );
  NAND4_X1 U12980 ( .A1(n10148), .A2(n10147), .A3(n10146), .A4(n10145), .ZN(
        n10149) );
  OR2_X2 U12981 ( .A1(n10150), .A2(n10149), .ZN(n13396) );
  AOI22_X1 U12982 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10154) );
  BUF_X4 U12983 ( .A(n10230), .Z(n11532) );
  AOI22_X1 U12984 ( .A1(n11532), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10342), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10153) );
  AOI22_X1 U12985 ( .A1(n10278), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10185), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10152) );
  AOI22_X1 U12986 ( .A1(n11474), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10409), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10151) );
  NAND4_X1 U12987 ( .A1(n10154), .A2(n10153), .A3(n10152), .A4(n10151), .ZN(
        n10160) );
  AOI22_X1 U12988 ( .A1(n10223), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10158) );
  AOI22_X1 U12989 ( .A1(n10175), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10186), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10157) );
  AOI22_X1 U12990 ( .A1(n10301), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10273), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10156) );
  AOI22_X1 U12991 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10300), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10155) );
  NAND4_X1 U12992 ( .A1(n10158), .A2(n10157), .A3(n10156), .A4(n10155), .ZN(
        n10159) );
  NAND2_X1 U12993 ( .A1(n10244), .A2(n20092), .ZN(n10170) );
  AOI22_X1 U12994 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10301), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10165) );
  AOI22_X1 U12995 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11532), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10164) );
  AOI22_X1 U12996 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10342), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10163) );
  AOI22_X1 U12997 ( .A1(n10278), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10273), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10162) );
  AOI22_X1 U12998 ( .A1(n11487), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10300), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10169) );
  AOI22_X1 U12999 ( .A1(n10272), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10185), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10168) );
  AOI22_X1 U13000 ( .A1(n10186), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10409), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10167) );
  AOI22_X1 U13001 ( .A1(n10223), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10166) );
  MUX2_X1 U13002 ( .A(n13390), .B(n10170), .S(n20098), .Z(n10198) );
  AOI22_X1 U13004 ( .A1(n10175), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11532), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10184) );
  AOI22_X1 U13005 ( .A1(n11487), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10300), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10177) );
  AOI22_X1 U13006 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10342), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10176) );
  AOI22_X1 U13007 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10181) );
  AOI22_X1 U13008 ( .A1(n10278), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10301), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10180) );
  AOI22_X1 U13009 ( .A1(n10273), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10185), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10179) );
  AOI22_X1 U13010 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10409), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10178) );
  AOI22_X1 U13011 ( .A1(n10223), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10182) );
  AOI21_X1 U13012 ( .B1(n12325), .B2(n13396), .A(n12765), .ZN(n10197) );
  NAND2_X2 U13013 ( .A1(n12633), .A2(n20092), .ZN(n12899) );
  AOI22_X1 U13014 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10190) );
  AOI22_X1 U13015 ( .A1(n10278), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10301), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10189) );
  AOI22_X1 U13016 ( .A1(n10273), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10185), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10188) );
  BUF_X2 U13017 ( .A(n10186), .Z(n11540) );
  AOI22_X1 U13018 ( .A1(n11540), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10409), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10187) );
  NAND4_X1 U13019 ( .A1(n10190), .A2(n10189), .A3(n10188), .A4(n10187), .ZN(
        n10196) );
  AOI22_X1 U13020 ( .A1(n10175), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11532), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10194) );
  AOI22_X1 U13021 ( .A1(n11487), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10300), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10193) );
  AOI22_X1 U13022 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10342), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10192) );
  AOI22_X1 U13023 ( .A1(n10223), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10191) );
  NAND4_X1 U13024 ( .A1(n10194), .A2(n10193), .A3(n10192), .A4(n10191), .ZN(
        n10195) );
  OR2_X2 U13025 ( .A1(n10196), .A2(n10195), .ZN(n20086) );
  NAND2_X1 U13026 ( .A1(n12899), .A2(n20086), .ZN(n10264) );
  NAND2_X1 U13027 ( .A1(n10272), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10202) );
  NAND2_X1 U13028 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10201) );
  NAND2_X1 U13029 ( .A1(n10278), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10200) );
  NAND2_X1 U13030 ( .A1(n10301), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10199) );
  NAND2_X1 U13031 ( .A1(n11474), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10206) );
  NAND2_X1 U13032 ( .A1(n10175), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10205) );
  NAND2_X1 U13033 ( .A1(n11532), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10204) );
  NAND2_X1 U13034 ( .A1(n10342), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10203) );
  NAND2_X1 U13035 ( .A1(n10223), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10210) );
  NAND2_X1 U13036 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10209) );
  NAND2_X1 U13037 ( .A1(n10300), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10208) );
  NAND2_X1 U13038 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10207) );
  NAND2_X1 U13039 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10214) );
  NAND2_X1 U13040 ( .A1(n10273), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10213) );
  NAND2_X1 U13041 ( .A1(n10185), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10212) );
  NAND2_X1 U13042 ( .A1(n10409), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10211) );
  AND4_X2 U13043 ( .A1(n10214), .A2(n10213), .A3(n10212), .A4(n10211), .ZN(
        n10215) );
  NAND4_X4 U13044 ( .A1(n10218), .A2(n10217), .A3(n10216), .A4(n10215), .ZN(
        n20074) );
  NAND2_X1 U13045 ( .A1(n10272), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10222) );
  NAND2_X1 U13046 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10221) );
  NAND2_X1 U13047 ( .A1(n10278), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10220) );
  NAND2_X1 U13048 ( .A1(n10301), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10219) );
  NAND2_X1 U13049 ( .A1(n10223), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10229) );
  NAND2_X1 U13050 ( .A1(n11487), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10228) );
  NAND2_X1 U13051 ( .A1(n10300), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10227) );
  NAND2_X1 U13052 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10226) );
  AND4_X2 U13053 ( .A1(n10229), .A2(n10228), .A3(n10227), .A4(n10226), .ZN(
        n10241) );
  NAND2_X1 U13054 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10234) );
  NAND2_X1 U13055 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10233) );
  NAND2_X1 U13056 ( .A1(n10273), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10232) );
  NAND2_X1 U13057 ( .A1(n10185), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10231) );
  AND4_X2 U13058 ( .A1(n10234), .A2(n10233), .A3(n10232), .A4(n10231), .ZN(
        n10240) );
  NAND2_X1 U13059 ( .A1(n10186), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10238) );
  NAND2_X1 U13060 ( .A1(n11474), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10237) );
  NAND2_X1 U13061 ( .A1(n10342), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10236) );
  NAND2_X1 U13062 ( .A1(n10409), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10235) );
  NAND4_X4 U13063 ( .A1(n10242), .A2(n10241), .A3(n10240), .A4(n10239), .ZN(
        n20080) );
  NAND2_X2 U13064 ( .A1(n13440), .A2(n12946), .ZN(n10261) );
  NAND2_X1 U13065 ( .A1(n12633), .A2(n12635), .ZN(n10243) );
  NAND2_X1 U13066 ( .A1(n11561), .A2(n10246), .ZN(n10584) );
  XNOR2_X1 U13067 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n10526) );
  NOR2_X2 U13068 ( .A1(n20086), .A2(n13396), .ZN(n12947) );
  NAND2_X1 U13069 ( .A1(n12947), .A2(n12634), .ZN(n12758) );
  NAND2_X1 U13070 ( .A1(n20098), .A2(n20105), .ZN(n11050) );
  OR2_X2 U13071 ( .A1(n10584), .A2(n10247), .ZN(n10259) );
  INV_X1 U13072 ( .A(n20086), .ZN(n10248) );
  NAND2_X4 U13073 ( .A1(n10248), .A2(n20074), .ZN(n10674) );
  NAND2_X2 U13074 ( .A1(n20086), .A2(n20080), .ZN(n10662) );
  NAND2_X1 U13075 ( .A1(n10586), .A2(n10573), .ZN(n10693) );
  NAND2_X1 U13076 ( .A1(n13440), .A2(n20080), .ZN(n13456) );
  NAND2_X1 U13077 ( .A1(n10693), .A2(n13456), .ZN(n10249) );
  NAND2_X1 U13078 ( .A1(n12946), .A2(n20074), .ZN(n20762) );
  OR2_X1 U13079 ( .A1(n12325), .A2(n10662), .ZN(n10698) );
  NAND2_X1 U13080 ( .A1(n13396), .A2(n20074), .ZN(n10690) );
  NOR2_X1 U13081 ( .A1(n10249), .A2(n10266), .ZN(n10255) );
  OR2_X1 U13082 ( .A1(n12899), .A2(n13390), .ZN(n10251) );
  NAND2_X1 U13083 ( .A1(n12634), .A2(n20098), .ZN(n10250) );
  NAND2_X1 U13084 ( .A1(n20105), .A2(n13390), .ZN(n10252) );
  NAND2_X1 U13085 ( .A1(n10577), .A2(n14637), .ZN(n10254) );
  OAI21_X1 U13086 ( .B1(n10260), .B2(n12947), .A(n13440), .ZN(n10253) );
  NAND3_X1 U13087 ( .A1(n10255), .A2(n10254), .A3(n10253), .ZN(n10256) );
  NAND2_X1 U13088 ( .A1(n19877), .A2(n20649), .ZN(n12330) );
  NAND2_X1 U13089 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10331) );
  OAI21_X1 U13090 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n10331), .ZN(n20399) );
  OR2_X1 U13091 ( .A1(n15834), .A2(n20475), .ZN(n10326) );
  OAI21_X1 U13092 ( .B1(n12330), .B2(n20399), .A(n10326), .ZN(n10257) );
  INV_X1 U13093 ( .A(n10257), .ZN(n10258) );
  MUX2_X1 U13094 ( .A(n15834), .B(n12330), .S(n20742), .Z(n10318) );
  NAND3_X1 U13095 ( .A1(n10577), .A2(n20080), .A3(n14637), .ZN(n10269) );
  NAND2_X1 U13096 ( .A1(n10260), .A2(n12624), .ZN(n12945) );
  AND2_X1 U13097 ( .A1(n10261), .A2(n10662), .ZN(n12623) );
  INV_X1 U13098 ( .A(n10262), .ZN(n10263) );
  AOI22_X1 U13099 ( .A1(n12623), .A2(n10264), .B1(n10479), .B2(n10263), .ZN(
        n10268) );
  NAND2_X1 U13100 ( .A1(n12947), .A2(n12633), .ZN(n10696) );
  NAND4_X1 U13101 ( .A1(n10696), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n19877), 
        .A4(n13456), .ZN(n10265) );
  NOR2_X1 U13102 ( .A1(n10266), .A2(n10265), .ZN(n10267) );
  NAND4_X1 U13103 ( .A1(n10269), .A2(n12945), .A3(n10268), .A4(n10267), .ZN(
        n11067) );
  INV_X1 U13104 ( .A(n20182), .ZN(n10271) );
  AOI22_X1 U13105 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10277) );
  AOI22_X1 U13106 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11532), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10276) );
  AOI22_X1 U13107 ( .A1(n10301), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10275) );
  AOI22_X1 U13108 ( .A1(n11540), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11539), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10274) );
  NAND4_X1 U13109 ( .A1(n10277), .A2(n10276), .A3(n10275), .A4(n10274), .ZN(
        n10284) );
  AOI22_X1 U13110 ( .A1(n11487), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10300), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10282) );
  AOI22_X1 U13111 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10281) );
  AOI22_X1 U13112 ( .A1(n10278), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10280) );
  AOI22_X1 U13113 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10279) );
  NAND4_X1 U13114 ( .A1(n10282), .A2(n10281), .A3(n10280), .A4(n10279), .ZN(
        n10283) );
  AOI22_X1 U13115 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10288) );
  AOI22_X1 U13116 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10300), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10287) );
  AOI22_X1 U13117 ( .A1(n10278), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10286) );
  AOI22_X1 U13118 ( .A1(n11474), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9619), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10285) );
  NAND4_X1 U13119 ( .A1(n10288), .A2(n10287), .A3(n10286), .A4(n10285), .ZN(
        n10295) );
  AOI22_X1 U13120 ( .A1(n11532), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10223), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10293) );
  AOI22_X1 U13121 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10342), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10292) );
  AOI22_X1 U13122 ( .A1(n10301), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11539), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10291) );
  BUF_X1 U13123 ( .A(n10409), .Z(n10289) );
  AOI22_X1 U13124 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10290) );
  NAND4_X1 U13125 ( .A1(n10293), .A2(n10292), .A3(n10291), .A4(n10290), .ZN(
        n10294) );
  NAND2_X1 U13126 ( .A1(n10319), .A2(n10357), .ZN(n10396) );
  OAI211_X1 U13127 ( .C1(n10357), .C2(n10319), .A(n10479), .B(n10396), .ZN(
        n10297) );
  NOR2_X1 U13128 ( .A1(n10573), .A2(n12634), .ZN(n10296) );
  AND2_X1 U13129 ( .A1(n10297), .A2(n10296), .ZN(n10298) );
  INV_X1 U13130 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20079) );
  AOI22_X1 U13131 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11474), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10305) );
  AOI22_X1 U13132 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10300), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10304) );
  AOI22_X1 U13133 ( .A1(n10301), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10303) );
  AOI22_X1 U13134 ( .A1(n11532), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10302) );
  NAND4_X1 U13135 ( .A1(n10305), .A2(n10304), .A3(n10303), .A4(n10302), .ZN(
        n10311) );
  AOI22_X1 U13136 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10309) );
  AOI22_X1 U13137 ( .A1(n10223), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10342), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10308) );
  AOI22_X1 U13138 ( .A1(n11540), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11539), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10307) );
  AOI22_X1 U13139 ( .A1(n10278), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10306) );
  NAND4_X1 U13140 ( .A1(n10309), .A2(n10308), .A3(n10307), .A4(n10306), .ZN(
        n10310) );
  AOI21_X1 U13141 ( .B1(n12635), .B2(n10478), .A(n20649), .ZN(n10313) );
  NAND2_X1 U13142 ( .A1(n13440), .A2(n10319), .ZN(n10312) );
  OAI211_X1 U13143 ( .C1(n10555), .C2(n20079), .A(n10313), .B(n10312), .ZN(
        n10363) );
  INV_X1 U13144 ( .A(n10478), .ZN(n10487) );
  NAND2_X1 U13145 ( .A1(n10314), .A2(n10487), .ZN(n10359) );
  NAND2_X1 U13146 ( .A1(n10314), .A2(n10478), .ZN(n10485) );
  INV_X1 U13147 ( .A(n10319), .ZN(n10315) );
  MUX2_X1 U13148 ( .A(n10359), .B(n10485), .S(n10315), .Z(n10316) );
  INV_X1 U13149 ( .A(n10316), .ZN(n10317) );
  XNOR2_X1 U13150 ( .A(n10363), .B(n10361), .ZN(n20739) );
  NAND2_X1 U13151 ( .A1(n20739), .A2(n10530), .ZN(n10322) );
  NAND2_X1 U13152 ( .A1(n13440), .A2(n20086), .ZN(n10370) );
  OAI21_X1 U13153 ( .B1(n20762), .B2(n10319), .A(n10370), .ZN(n10320) );
  INV_X1 U13154 ( .A(n10320), .ZN(n10321) );
  NAND2_X1 U13155 ( .A1(n10322), .A2(n10321), .ZN(n12809) );
  NAND2_X1 U13156 ( .A1(n12809), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12808) );
  XNOR2_X1 U13157 ( .A(n10324), .B(n12808), .ZN(n12740) );
  NAND2_X1 U13158 ( .A1(n12740), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12741) );
  INV_X1 U13159 ( .A(n12808), .ZN(n10323) );
  NAND2_X1 U13160 ( .A1(n10324), .A2(n10323), .ZN(n10325) );
  INV_X1 U13161 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20067) );
  XNOR2_X1 U13162 ( .A(n10374), .B(n20067), .ZN(n12938) );
  INV_X1 U13163 ( .A(n10326), .ZN(n10329) );
  INV_X1 U13164 ( .A(n10327), .ZN(n10328) );
  INV_X1 U13165 ( .A(n12330), .ZN(n10333) );
  INV_X1 U13166 ( .A(n10331), .ZN(n10330) );
  NAND2_X1 U13167 ( .A1(n10330), .A2(n20395), .ZN(n20443) );
  NAND2_X1 U13168 ( .A1(n10331), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10332) );
  NAND2_X1 U13169 ( .A1(n20443), .A2(n10332), .ZN(n13382) );
  NAND2_X1 U13170 ( .A1(n10333), .A2(n13382), .ZN(n10334) );
  INV_X1 U13171 ( .A(n10336), .ZN(n10337) );
  AND2_X1 U13172 ( .A1(n10338), .A2(n10337), .ZN(n10339) );
  NAND2_X1 U13173 ( .A1(n10340), .A2(n10339), .ZN(n10341) );
  AOI22_X1 U13174 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11532), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10346) );
  AOI22_X1 U13175 ( .A1(n11487), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10300), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10345) );
  AOI22_X1 U13176 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10342), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10344) );
  AOI22_X1 U13177 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10343) );
  NAND4_X1 U13178 ( .A1(n10346), .A2(n10345), .A3(n10344), .A4(n10343), .ZN(
        n10352) );
  AOI22_X1 U13179 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10350) );
  AOI22_X1 U13180 ( .A1(n11538), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10301), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10349) );
  AOI22_X1 U13181 ( .A1(n11539), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10348) );
  AOI22_X1 U13182 ( .A1(n11540), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10347) );
  NAND4_X1 U13183 ( .A1(n10350), .A2(n10349), .A3(n10348), .A4(n10347), .ZN(
        n10351) );
  OAI22_X2 U13184 ( .A1(n12943), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n10395), 
        .B2(n10382), .ZN(n10356) );
  INV_X1 U13185 ( .A(n10381), .ZN(n10354) );
  AOI22_X1 U13186 ( .A1(n10559), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10354), .B2(n10353), .ZN(n10355) );
  INV_X1 U13187 ( .A(n10357), .ZN(n10360) );
  NAND2_X1 U13188 ( .A1(n10559), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10358) );
  OAI211_X1 U13189 ( .C1(n10360), .C2(n10381), .A(n10359), .B(n10358), .ZN(
        n10365) );
  INV_X1 U13190 ( .A(n10361), .ZN(n10362) );
  NAND2_X1 U13191 ( .A1(n10363), .A2(n10362), .ZN(n10364) );
  NAND2_X1 U13192 ( .A1(n10364), .A2(n10485), .ZN(n10366) );
  NAND2_X1 U13193 ( .A1(n10366), .A2(n10365), .ZN(n10367) );
  NAND2_X1 U13194 ( .A1(n11057), .A2(n11058), .ZN(n11062) );
  INV_X1 U13195 ( .A(n10530), .ZN(n10484) );
  XNOR2_X1 U13196 ( .A(n10396), .B(n10395), .ZN(n10372) );
  INV_X1 U13197 ( .A(n10370), .ZN(n10371) );
  AOI21_X1 U13198 ( .B1(n10372), .B2(n10479), .A(n10371), .ZN(n10373) );
  NAND2_X1 U13199 ( .A1(n12938), .A2(n12937), .ZN(n12936) );
  NAND2_X1 U13200 ( .A1(n10374), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10375) );
  INV_X1 U13201 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20052) );
  OR2_X1 U13202 ( .A1(n10376), .A2(n9816), .ZN(n10380) );
  NOR3_X1 U13203 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20395), .A3(
        n20475), .ZN(n20319) );
  NAND2_X1 U13204 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20319), .ZN(
        n20314) );
  NAND2_X1 U13205 ( .A1(n20442), .A2(n20314), .ZN(n10377) );
  NAND3_X1 U13206 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20585) );
  INV_X1 U13207 ( .A(n20585), .ZN(n20594) );
  NAND2_X1 U13208 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20594), .ZN(
        n20582) );
  NAND2_X1 U13209 ( .A1(n10377), .A2(n20582), .ZN(n20340) );
  OAI22_X1 U13210 ( .A1(n12330), .A2(n20340), .B1(n15834), .B2(n20442), .ZN(
        n10378) );
  INV_X1 U13211 ( .A(n10378), .ZN(n10379) );
  AOI22_X1 U13212 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10386) );
  AOI22_X1 U13213 ( .A1(n11538), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10301), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10385) );
  AOI22_X1 U13214 ( .A1(n11539), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10384) );
  AOI22_X1 U13215 ( .A1(n11540), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10383) );
  NAND4_X1 U13216 ( .A1(n10386), .A2(n10385), .A3(n10384), .A4(n10383), .ZN(
        n10392) );
  AOI22_X1 U13217 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11532), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10390) );
  AOI22_X1 U13218 ( .A1(n11487), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12958), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10389) );
  AOI22_X1 U13219 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10388) );
  INV_X1 U13220 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n20091) );
  AOI22_X1 U13221 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9619), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10387) );
  NAND4_X1 U13222 ( .A1(n10390), .A2(n10389), .A3(n10388), .A4(n10387), .ZN(
        n10391) );
  AOI22_X1 U13223 ( .A1(n10550), .A2(n10444), .B1(n10559), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10393) );
  XNOR2_X2 U13224 ( .A(n10403), .B(n12988), .ZN(n13379) );
  NAND2_X1 U13225 ( .A1(n13379), .A2(n10530), .ZN(n10400) );
  NAND2_X1 U13226 ( .A1(n10396), .A2(n10395), .ZN(n10446) );
  INV_X1 U13227 ( .A(n10444), .ZN(n10397) );
  XNOR2_X1 U13228 ( .A(n10446), .B(n10397), .ZN(n10398) );
  NAND2_X1 U13229 ( .A1(n10398), .A2(n10479), .ZN(n10399) );
  NAND2_X1 U13230 ( .A1(n10400), .A2(n10399), .ZN(n13159) );
  NAND2_X1 U13231 ( .A1(n10401), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10402) );
  AOI22_X1 U13232 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11509), .B1(
        n11516), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10408) );
  AOI22_X1 U13233 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12958), .B1(
        n11487), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10407) );
  AOI22_X1 U13234 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10406) );
  AOI22_X1 U13235 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10405) );
  NAND4_X1 U13236 ( .A1(n10408), .A2(n10407), .A3(n10406), .A4(n10405), .ZN(
        n10415) );
  AOI22_X1 U13237 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10161), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10413) );
  AOI22_X1 U13238 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n10301), .B1(
        n11538), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10412) );
  AOI22_X1 U13239 ( .A1(n11539), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10411) );
  AOI22_X1 U13240 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11532), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10410) );
  NAND4_X1 U13241 ( .A1(n10413), .A2(n10412), .A3(n10411), .A4(n10410), .ZN(
        n10414) );
  NAND2_X1 U13242 ( .A1(n10550), .A2(n10443), .ZN(n10417) );
  NAND2_X1 U13243 ( .A1(n10559), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10416) );
  NAND2_X1 U13244 ( .A1(n10417), .A2(n10416), .ZN(n10425) );
  XNOR2_X1 U13245 ( .A(n10424), .B(n10425), .ZN(n11099) );
  NAND2_X1 U13246 ( .A1(n11099), .A2(n10530), .ZN(n10421) );
  NAND2_X1 U13247 ( .A1(n10446), .A2(n10444), .ZN(n10418) );
  XNOR2_X1 U13248 ( .A(n10418), .B(n10443), .ZN(n10419) );
  NAND2_X1 U13249 ( .A1(n10419), .A2(n10479), .ZN(n10420) );
  NAND2_X1 U13250 ( .A1(n10421), .A2(n10420), .ZN(n10422) );
  INV_X1 U13251 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20044) );
  XNOR2_X1 U13252 ( .A(n10422), .B(n20044), .ZN(n20015) );
  NAND2_X1 U13253 ( .A1(n10422), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10423) );
  AOI22_X1 U13254 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11532), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10429) );
  AOI22_X1 U13255 ( .A1(n11487), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12958), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10428) );
  INV_X1 U13256 ( .A(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n20844) );
  AOI22_X1 U13257 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10427) );
  AOI22_X1 U13258 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10426) );
  NAND4_X1 U13259 ( .A1(n10429), .A2(n10428), .A3(n10427), .A4(n10426), .ZN(
        n10435) );
  AOI22_X1 U13260 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10433) );
  AOI22_X1 U13261 ( .A1(n11538), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10301), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10432) );
  AOI22_X1 U13262 ( .A1(n11539), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10431) );
  AOI22_X1 U13263 ( .A1(n11540), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10430) );
  NAND4_X1 U13264 ( .A1(n10433), .A2(n10432), .A3(n10431), .A4(n10430), .ZN(
        n10434) );
  NAND2_X1 U13265 ( .A1(n10550), .A2(n10465), .ZN(n10437) );
  NAND2_X1 U13266 ( .A1(n10559), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10436) );
  NAND2_X1 U13267 ( .A1(n10441), .A2(n10440), .ZN(n10442) );
  AND2_X1 U13268 ( .A1(n10444), .A2(n10443), .ZN(n10445) );
  NAND2_X1 U13269 ( .A1(n10446), .A2(n10445), .ZN(n10464) );
  XNOR2_X1 U13270 ( .A(n10464), .B(n10465), .ZN(n10447) );
  NAND2_X1 U13271 ( .A1(n10447), .A2(n10479), .ZN(n10448) );
  INV_X1 U13272 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16104) );
  AOI22_X1 U13273 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10453) );
  AOI22_X1 U13274 ( .A1(n11538), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10301), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10452) );
  AOI22_X1 U13275 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10451) );
  AOI22_X1 U13276 ( .A1(n11539), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10450) );
  NAND4_X1 U13277 ( .A1(n10453), .A2(n10452), .A3(n10451), .A4(n10450), .ZN(
        n10459) );
  AOI22_X1 U13278 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11474), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10457) );
  AOI22_X1 U13279 ( .A1(n11487), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12958), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10456) );
  AOI22_X1 U13280 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10455) );
  AOI22_X1 U13281 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9619), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10454) );
  NAND4_X1 U13282 ( .A1(n10457), .A2(n10456), .A3(n10455), .A4(n10454), .ZN(
        n10458) );
  NAND2_X1 U13283 ( .A1(n10550), .A2(n10476), .ZN(n10461) );
  NAND2_X1 U13284 ( .A1(n10559), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10460) );
  NAND2_X1 U13285 ( .A1(n10463), .A2(n10462), .ZN(n11104) );
  NAND3_X1 U13286 ( .A1(n10474), .A2(n10530), .A3(n11104), .ZN(n10469) );
  INV_X1 U13287 ( .A(n10464), .ZN(n10466) );
  NAND2_X1 U13288 ( .A1(n10466), .A2(n10465), .ZN(n10475) );
  XNOR2_X1 U13289 ( .A(n10475), .B(n10476), .ZN(n10467) );
  NAND2_X1 U13290 ( .A1(n10467), .A2(n10479), .ZN(n10468) );
  NAND2_X1 U13291 ( .A1(n10469), .A2(n10468), .ZN(n15995) );
  OR2_X1 U13292 ( .A1(n15995), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10470) );
  NAND2_X1 U13293 ( .A1(n15995), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10471) );
  INV_X1 U13294 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n20113) );
  NAND2_X1 U13295 ( .A1(n10550), .A2(n10478), .ZN(n10472) );
  OAI21_X1 U13296 ( .B1(n20113), .B2(n10555), .A(n10472), .ZN(n10473) );
  NAND2_X1 U13297 ( .A1(n11117), .A2(n10530), .ZN(n10482) );
  INV_X1 U13298 ( .A(n10475), .ZN(n10477) );
  NAND2_X1 U13299 ( .A1(n10477), .A2(n10476), .ZN(n10488) );
  XNOR2_X1 U13300 ( .A(n10488), .B(n10478), .ZN(n10480) );
  NAND2_X1 U13301 ( .A1(n10480), .A2(n10479), .ZN(n10481) );
  NAND2_X1 U13302 ( .A1(n10482), .A2(n10481), .ZN(n10483) );
  OR2_X1 U13303 ( .A1(n10483), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15989) );
  NAND2_X1 U13304 ( .A1(n10483), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15988) );
  NOR2_X1 U13305 ( .A1(n10485), .A2(n10484), .ZN(n10486) );
  OR3_X1 U13306 ( .A1(n10488), .A2(n10487), .A3(n20762), .ZN(n10489) );
  NAND2_X1 U13307 ( .A1(n9611), .A2(n10489), .ZN(n13604) );
  OR2_X1 U13308 ( .A1(n13604), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10490) );
  NAND2_X1 U13309 ( .A1(n13604), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10491) );
  INV_X1 U13310 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16081) );
  INV_X1 U13311 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10716) );
  NAND2_X1 U13312 ( .A1(n9611), .A2(n10716), .ZN(n10492) );
  NAND2_X1 U13313 ( .A1(n13777), .A2(n10492), .ZN(n14473) );
  INV_X1 U13314 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10499) );
  NAND2_X1 U13315 ( .A1(n15980), .A2(n10499), .ZN(n14471) );
  NAND2_X1 U13316 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10493) );
  NAND2_X1 U13317 ( .A1(n15980), .A2(n10493), .ZN(n14468) );
  NAND2_X1 U13318 ( .A1(n14471), .A2(n14468), .ZN(n10494) );
  NOR2_X1 U13319 ( .A1(n14473), .A2(n10494), .ZN(n13779) );
  INV_X1 U13320 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14610) );
  NAND2_X1 U13321 ( .A1(n15980), .A2(n14610), .ZN(n10495) );
  INV_X1 U13322 ( .A(n9611), .ZN(n14437) );
  NAND2_X1 U13323 ( .A1(n15980), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10497) );
  NAND2_X1 U13324 ( .A1(n15956), .A2(n10497), .ZN(n14457) );
  INV_X1 U13325 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10501) );
  NAND2_X1 U13326 ( .A1(n15980), .A2(n10501), .ZN(n15962) );
  OAI21_X1 U13327 ( .B1(n14437), .B2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15953), .ZN(n10498) );
  NOR2_X1 U13328 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10500) );
  NAND2_X1 U13329 ( .A1(n14470), .A2(n14466), .ZN(n13775) );
  NOR2_X1 U13330 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10502) );
  OAI21_X1 U13331 ( .B1(n10502), .B2(n9611), .A(n15963), .ZN(n10503) );
  NAND2_X1 U13332 ( .A1(n13777), .A2(n10504), .ZN(n14455) );
  XNOR2_X1 U13333 ( .A(n9611), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14449) );
  NAND3_X1 U13334 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14571) );
  INV_X1 U13335 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14438) );
  INV_X1 U13336 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16014) );
  INV_X1 U13337 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14600) );
  INV_X1 U13338 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14589) );
  NAND4_X1 U13339 ( .A1(n14438), .A2(n16014), .A3(n14600), .A4(n14589), .ZN(
        n10507) );
  AND2_X1 U13340 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14526) );
  NAND2_X1 U13341 ( .A1(n14526), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14528) );
  NAND2_X1 U13342 ( .A1(n14417), .A2(n14528), .ZN(n10509) );
  NAND2_X1 U13343 ( .A1(n10508), .A2(n9611), .ZN(n14395) );
  NAND3_X1 U13344 ( .A1(n10509), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14395), .ZN(n14378) );
  INV_X1 U13345 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14561) );
  INV_X1 U13346 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14398) );
  INV_X1 U13347 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14408) );
  NAND3_X1 U13348 ( .A1(n14561), .A2(n14398), .A3(n14408), .ZN(n14369) );
  NOR2_X1 U13349 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14506) );
  AND2_X1 U13350 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14507) );
  INV_X1 U13351 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14499) );
  XNOR2_X1 U13352 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10521) );
  NAND2_X1 U13353 ( .A1(n20742), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10533) );
  NAND2_X1 U13354 ( .A1(n10521), .A2(n10520), .ZN(n10514) );
  NAND2_X1 U13355 ( .A1(n20475), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10513) );
  NAND2_X1 U13356 ( .A1(n10514), .A2(n10513), .ZN(n10523) );
  XNOR2_X1 U13357 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10522) );
  XNOR2_X1 U13358 ( .A(n9816), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10518) );
  INV_X1 U13359 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16116) );
  INV_X1 U13360 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20072) );
  NOR2_X1 U13361 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20072), .ZN(
        n10515) );
  AOI221_X1 U13362 ( .B1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n10524), 
        .C1(n16116), .C2(n10524), .A(n10515), .ZN(n10531) );
  AOI21_X1 U13363 ( .B1(n10518), .B2(n10517), .A(n10516), .ZN(n10519) );
  INV_X1 U13364 ( .A(n10519), .ZN(n10557) );
  XNOR2_X1 U13365 ( .A(n10521), .B(n10520), .ZN(n10543) );
  XNOR2_X1 U13366 ( .A(n10523), .B(n10522), .ZN(n10549) );
  NOR3_X1 U13367 ( .A1(n10557), .A2(n10543), .A3(n10549), .ZN(n10525) );
  NAND3_X1 U13368 ( .A1(n16116), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n10524), .ZN(n10563) );
  OAI21_X1 U13369 ( .B1(n10531), .B2(n10525), .A(n10563), .ZN(n12639) );
  INV_X1 U13370 ( .A(n10526), .ZN(n10528) );
  INV_X1 U13371 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n10527) );
  NAND2_X1 U13372 ( .A1(n10528), .A2(n10527), .ZN(n15849) );
  NAND2_X1 U13373 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20659) );
  INV_X1 U13374 ( .A(n20659), .ZN(n20759) );
  AOI21_X1 U13375 ( .B1(n20080), .B2(n15849), .A(n20759), .ZN(n10529) );
  NAND2_X1 U13376 ( .A1(n12639), .A2(n10529), .ZN(n10572) );
  NAND2_X1 U13377 ( .A1(n10531), .A2(n10558), .ZN(n10568) );
  NAND2_X1 U13378 ( .A1(n10531), .A2(n10550), .ZN(n10566) );
  INV_X1 U13379 ( .A(n10558), .ZN(n10562) );
  AOI22_X1 U13380 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n12634), .B1(n10550), 
        .B2(n20080), .ZN(n10545) );
  INV_X1 U13381 ( .A(n10545), .ZN(n10532) );
  NOR2_X1 U13382 ( .A1(n10543), .A2(n10532), .ZN(n10538) );
  INV_X1 U13383 ( .A(n12325), .ZN(n12631) );
  OAI21_X1 U13384 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20742), .A(
        n10533), .ZN(n10534) );
  AOI21_X1 U13385 ( .B1(n12634), .B2(n20074), .A(n20080), .ZN(n10551) );
  AOI211_X1 U13386 ( .C1(n12631), .C2(n20074), .A(n10534), .B(n10551), .ZN(
        n10537) );
  INV_X1 U13387 ( .A(n10534), .ZN(n10535) );
  AOI21_X1 U13388 ( .B1(n10550), .B2(n10535), .A(n10558), .ZN(n10536) );
  NAND2_X1 U13389 ( .A1(n10538), .A2(n10544), .ZN(n10548) );
  INV_X1 U13390 ( .A(n10550), .ZN(n10541) );
  INV_X1 U13391 ( .A(n10551), .ZN(n10540) );
  NAND2_X1 U13392 ( .A1(n10559), .A2(n10549), .ZN(n10539) );
  OAI211_X1 U13393 ( .C1(n10541), .C2(n10549), .A(n10540), .B(n10539), .ZN(
        n10547) );
  NAND2_X1 U13394 ( .A1(n10545), .A2(n20080), .ZN(n10542) );
  OAI211_X1 U13395 ( .C1(n10545), .C2(n10544), .A(n10543), .B(n10542), .ZN(
        n10546) );
  NAND3_X1 U13396 ( .A1(n10548), .A2(n10547), .A3(n10546), .ZN(n10554) );
  INV_X1 U13397 ( .A(n10549), .ZN(n10552) );
  NAND3_X1 U13398 ( .A1(n10552), .A2(n10551), .A3(n10550), .ZN(n10553) );
  AOI22_X1 U13399 ( .A1(n10555), .A2(n10557), .B1(n10554), .B2(n10553), .ZN(
        n10556) );
  AOI21_X1 U13400 ( .B1(n10558), .B2(n10557), .A(n10556), .ZN(n10561) );
  NOR2_X1 U13401 ( .A1(n10559), .A2(n10563), .ZN(n10560) );
  OAI22_X1 U13402 ( .A1(n10563), .A2(n10562), .B1(n10561), .B2(n10560), .ZN(
        n10564) );
  AOI21_X1 U13403 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20649), .A(
        n10564), .ZN(n10565) );
  NAND2_X1 U13404 ( .A1(n10566), .A2(n10565), .ZN(n10567) );
  NAND2_X1 U13405 ( .A1(n20080), .A2(n20659), .ZN(n12703) );
  OR2_X1 U13406 ( .A1(n15849), .A2(n20759), .ZN(n12798) );
  NAND2_X1 U13407 ( .A1(n12703), .A2(n12798), .ZN(n13451) );
  INV_X1 U13408 ( .A(n13451), .ZN(n10569) );
  OAI211_X1 U13409 ( .C1(n10569), .C2(n14262), .A(n20074), .B(n11050), .ZN(
        n10570) );
  NAND2_X1 U13410 ( .A1(n12800), .A2(n10570), .ZN(n10571) );
  MUX2_X1 U13411 ( .A(n10572), .B(n10571), .S(n10244), .Z(n10580) );
  AND2_X1 U13412 ( .A1(n10685), .A2(n13440), .ZN(n12640) );
  AOI21_X1 U13413 ( .B1(n14637), .B2(n13440), .A(n10573), .ZN(n10574) );
  NAND2_X1 U13414 ( .A1(n10574), .A2(n10702), .ZN(n12327) );
  INV_X1 U13415 ( .A(n12327), .ZN(n12632) );
  OR2_X1 U13416 ( .A1(n12640), .A2(n12632), .ZN(n10578) );
  NAND2_X1 U13417 ( .A1(n12899), .A2(n20074), .ZN(n10575) );
  NAND2_X1 U13418 ( .A1(n10575), .A2(n20762), .ZN(n10576) );
  NAND2_X1 U13419 ( .A1(n10577), .A2(n10576), .ZN(n10689) );
  OR3_X1 U13420 ( .A1(n12800), .A2(n12946), .A3(n14637), .ZN(n10579) );
  NAND3_X1 U13421 ( .A1(n10580), .A2(n12796), .A3(n10579), .ZN(n10581) );
  NAND2_X1 U13422 ( .A1(n15834), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19878) );
  INV_X1 U13423 ( .A(n19878), .ZN(n12763) );
  NOR2_X1 U13424 ( .A1(n12631), .A2(n12624), .ZN(n10582) );
  OAI22_X1 U13425 ( .A1(n10582), .A2(n12327), .B1(n10683), .B2(n12635), .ZN(
        n10583) );
  OR2_X1 U13426 ( .A1(n10584), .A2(n10583), .ZN(n10585) );
  AND2_X1 U13427 ( .A1(n12817), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10587) );
  AOI21_X1 U13428 ( .B1(n12766), .B2(P1_EBX_REG_30__SCAN_IN), .A(n10587), .ZN(
        n14062) );
  INV_X1 U13429 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14641) );
  NAND2_X1 U13430 ( .A1(n10674), .A2(n14641), .ZN(n10590) );
  INV_X1 U13431 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n10588) );
  NAND2_X1 U13432 ( .A1(n10677), .A2(n10588), .ZN(n10589) );
  NAND3_X1 U13433 ( .A1(n10590), .A2(n10662), .A3(n10589), .ZN(n10591) );
  NAND2_X1 U13434 ( .A1(n10674), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n10593) );
  INV_X1 U13435 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n12769) );
  NAND2_X1 U13436 ( .A1(n10662), .A2(n12769), .ZN(n10592) );
  XNOR2_X1 U13437 ( .A(n10594), .B(n12768), .ZN(n19975) );
  NAND2_X1 U13438 ( .A1(n10674), .A2(n20067), .ZN(n10598) );
  INV_X1 U13439 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n10596) );
  NAND2_X1 U13440 ( .A1(n10677), .A2(n10596), .ZN(n10597) );
  NAND3_X1 U13441 ( .A1(n10598), .A2(n10662), .A3(n10597), .ZN(n10599) );
  OAI21_X1 U13442 ( .B1(P1_EBX_REG_2__SCAN_IN), .B2(n10680), .A(n10599), .ZN(
        n12842) );
  MUX2_X1 U13443 ( .A(n10653), .B(n10662), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n10600) );
  OAI21_X1 U13444 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n12766), .A(
        n10600), .ZN(n13100) );
  MUX2_X1 U13445 ( .A(n10680), .B(n10674), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n10603) );
  OAI21_X1 U13446 ( .B1(n10677), .B2(n20044), .A(n10639), .ZN(n10601) );
  INV_X1 U13447 ( .A(n10601), .ZN(n10602) );
  NAND2_X1 U13448 ( .A1(n10603), .A2(n10602), .ZN(n13179) );
  NAND2_X1 U13449 ( .A1(n10662), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10604) );
  OAI211_X1 U13450 ( .C1(n12817), .C2(P1_EBX_REG_5__SCAN_IN), .A(n10674), .B(
        n10604), .ZN(n10605) );
  OAI21_X1 U13451 ( .B1(n10653), .B2(P1_EBX_REG_5__SCAN_IN), .A(n10605), .ZN(
        n13170) );
  INV_X1 U13452 ( .A(n10674), .ZN(n10627) );
  MUX2_X1 U13453 ( .A(n10676), .B(n10627), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n10608) );
  INV_X1 U13454 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10606) );
  OAI21_X1 U13455 ( .B1(n10677), .B2(n10606), .A(n10639), .ZN(n10607) );
  INV_X1 U13456 ( .A(n10653), .ZN(n10670) );
  INV_X1 U13457 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n10609) );
  NAND2_X1 U13458 ( .A1(n10670), .A2(n10609), .ZN(n10613) );
  NAND2_X1 U13459 ( .A1(n10677), .A2(n10609), .ZN(n10611) );
  NAND2_X1 U13460 ( .A1(n10662), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10610) );
  NAND3_X1 U13461 ( .A1(n10611), .A2(n10674), .A3(n10610), .ZN(n10612) );
  AND2_X1 U13462 ( .A1(n10613), .A2(n10612), .ZN(n13209) );
  NAND2_X1 U13463 ( .A1(n13210), .A2(n13209), .ZN(n13417) );
  MUX2_X1 U13464 ( .A(n10676), .B(n10627), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n10616) );
  NAND2_X1 U13465 ( .A1(n12817), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10614) );
  NAND2_X1 U13466 ( .A1(n10639), .A2(n10614), .ZN(n10615) );
  NOR2_X1 U13467 ( .A1(n10616), .A2(n10615), .ZN(n13416) );
  INV_X1 U13468 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n10617) );
  NAND2_X1 U13469 ( .A1(n10677), .A2(n10617), .ZN(n10619) );
  NAND2_X1 U13470 ( .A1(n10662), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10618) );
  NAND3_X1 U13471 ( .A1(n10619), .A2(n10674), .A3(n10618), .ZN(n10620) );
  OAI21_X1 U13472 ( .B1(n10653), .B2(P1_EBX_REG_9__SCAN_IN), .A(n10620), .ZN(
        n13469) );
  INV_X1 U13473 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n20911) );
  NAND2_X1 U13474 ( .A1(n10676), .A2(n20911), .ZN(n10624) );
  NAND2_X1 U13475 ( .A1(n10674), .A2(n16074), .ZN(n10622) );
  NAND2_X1 U13476 ( .A1(n10677), .A2(n20911), .ZN(n10621) );
  NAND3_X1 U13477 ( .A1(n10622), .A2(n10662), .A3(n10621), .ZN(n10623) );
  MUX2_X1 U13478 ( .A(n10653), .B(n10662), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n10626) );
  OR2_X1 U13479 ( .A1(n12766), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10625) );
  AND2_X1 U13480 ( .A1(n10626), .A2(n10625), .ZN(n13736) );
  MUX2_X1 U13481 ( .A(n10676), .B(n10627), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n10630) );
  NAND2_X1 U13482 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n12817), .ZN(
        n10628) );
  NAND2_X1 U13483 ( .A1(n10639), .A2(n10628), .ZN(n10629) );
  NOR2_X1 U13484 ( .A1(n10630), .A2(n10629), .ZN(n13795) );
  MUX2_X1 U13485 ( .A(n10653), .B(n10662), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n10631) );
  OAI21_X1 U13486 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n12766), .A(
        n10631), .ZN(n13752) );
  NOR2_X1 U13487 ( .A1(n13795), .A2(n13752), .ZN(n10632) );
  INV_X1 U13488 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15923) );
  NAND2_X1 U13489 ( .A1(n10676), .A2(n15923), .ZN(n10636) );
  NAND2_X1 U13490 ( .A1(n10674), .A2(n14610), .ZN(n10634) );
  NAND2_X1 U13491 ( .A1(n10677), .A2(n15923), .ZN(n10633) );
  NAND3_X1 U13492 ( .A1(n10634), .A2(n10662), .A3(n10633), .ZN(n10635) );
  AND2_X1 U13493 ( .A1(n10636), .A2(n10635), .ZN(n13745) );
  MUX2_X1 U13494 ( .A(n10653), .B(n10662), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n10637) );
  OAI21_X1 U13495 ( .B1(n12766), .B2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n10637), .ZN(n13803) );
  MUX2_X1 U13496 ( .A(n10680), .B(n10674), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n10641) );
  NAND2_X1 U13497 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n12817), .ZN(
        n10638) );
  AND2_X1 U13498 ( .A1(n10639), .A2(n10638), .ZN(n10640) );
  NAND2_X1 U13499 ( .A1(n10641), .A2(n10640), .ZN(n14182) );
  MUX2_X1 U13500 ( .A(n10653), .B(n10662), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n10642) );
  OAI21_X1 U13501 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n12766), .A(
        n10642), .ZN(n14247) );
  INV_X1 U13502 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15898) );
  NAND2_X1 U13503 ( .A1(n10676), .A2(n15898), .ZN(n10646) );
  NAND2_X1 U13504 ( .A1(n10674), .A2(n16014), .ZN(n10644) );
  NAND2_X1 U13505 ( .A1(n10677), .A2(n15898), .ZN(n10643) );
  NAND3_X1 U13506 ( .A1(n10644), .A2(n10662), .A3(n10643), .ZN(n10645) );
  MUX2_X1 U13507 ( .A(n10653), .B(n10662), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n10647) );
  OAI21_X1 U13508 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n12766), .A(
        n10647), .ZN(n10648) );
  INV_X1 U13509 ( .A(n10648), .ZN(n14232) );
  MUX2_X1 U13510 ( .A(n10680), .B(n10674), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n10650) );
  NAND2_X1 U13511 ( .A1(n12817), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10649) );
  NAND2_X1 U13512 ( .A1(n10650), .A2(n10649), .ZN(n14229) );
  NAND2_X1 U13513 ( .A1(n10662), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10651) );
  OAI211_X1 U13514 ( .C1(n12817), .C2(P1_EBX_REG_21__SCAN_IN), .A(n10674), .B(
        n10651), .ZN(n10652) );
  OAI21_X1 U13515 ( .B1(n10653), .B2(P1_EBX_REG_21__SCAN_IN), .A(n10652), .ZN(
        n14220) );
  MUX2_X1 U13516 ( .A(n10653), .B(n10662), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n10655) );
  OR2_X1 U13517 ( .A1(n12766), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10654) );
  NAND2_X1 U13518 ( .A1(n10655), .A2(n10654), .ZN(n14146) );
  INV_X1 U13519 ( .A(n14146), .ZN(n10660) );
  INV_X1 U13520 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14572) );
  NAND2_X1 U13521 ( .A1(n10674), .A2(n14572), .ZN(n10658) );
  INV_X1 U13522 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n10656) );
  NAND2_X1 U13523 ( .A1(n10677), .A2(n10656), .ZN(n10657) );
  NAND3_X1 U13524 ( .A1(n10658), .A2(n10662), .A3(n10657), .ZN(n10659) );
  OAI21_X1 U13525 ( .B1(P1_EBX_REG_22__SCAN_IN), .B2(n10680), .A(n10659), .ZN(
        n14165) );
  NAND2_X1 U13526 ( .A1(n10660), .A2(n14165), .ZN(n10661) );
  INV_X1 U13527 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n10665) );
  INV_X1 U13528 ( .A(n10662), .ZN(n14060) );
  NOR2_X1 U13529 ( .A1(n12817), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n10663) );
  AOI211_X1 U13530 ( .C1(n10674), .C2(n14408), .A(n14060), .B(n10663), .ZN(
        n10664) );
  AOI21_X1 U13531 ( .B1(n10676), .B2(n10665), .A(n10664), .ZN(n14137) );
  INV_X1 U13532 ( .A(n12766), .ZN(n10672) );
  MUX2_X1 U13533 ( .A(n10670), .B(n14060), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n10666) );
  AOI21_X1 U13534 ( .B1(n10672), .B2(n14398), .A(n10666), .ZN(n14129) );
  INV_X1 U13535 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n10669) );
  INV_X1 U13536 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14529) );
  NOR2_X1 U13537 ( .A1(n12817), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n10667) );
  AOI211_X1 U13538 ( .C1(n10674), .C2(n14529), .A(n14060), .B(n10667), .ZN(
        n10668) );
  AOI21_X1 U13539 ( .B1(n10676), .B2(n10669), .A(n10668), .ZN(n14111) );
  INV_X1 U13540 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14520) );
  MUX2_X1 U13541 ( .A(n10670), .B(n14060), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n10671) );
  AOI21_X1 U13542 ( .B1(n10672), .B2(n14520), .A(n10671), .ZN(n14104) );
  INV_X1 U13543 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14087) );
  INV_X1 U13544 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14373) );
  NOR2_X1 U13545 ( .A1(n12817), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n10673) );
  AOI211_X1 U13546 ( .C1(n10674), .C2(n14373), .A(n14060), .B(n10673), .ZN(
        n10675) );
  AOI21_X1 U13547 ( .B1(n10676), .B2(n14087), .A(n10675), .ZN(n14092) );
  OR2_X1 U13548 ( .A1(n12766), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10679) );
  INV_X1 U13549 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14205) );
  NAND2_X1 U13550 ( .A1(n10677), .A2(n14205), .ZN(n10678) );
  NAND2_X1 U13551 ( .A1(n10679), .A2(n10678), .ZN(n14058) );
  OAI22_X1 U13552 ( .A1(n14058), .A2(n14060), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n10680), .ZN(n14071) );
  NAND2_X1 U13553 ( .A1(n14091), .A2(n14071), .ZN(n14070) );
  MUX2_X1 U13554 ( .A(n14062), .B(n10662), .S(n14070), .Z(n10682) );
  AOI22_X1 U13555 ( .A1(n12766), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n12817), .ZN(n10681) );
  OR2_X1 U13556 ( .A1(n12626), .A2(n20080), .ZN(n12744) );
  OAI21_X1 U13557 ( .B1(n10683), .B2(n13390), .A(n12744), .ZN(n10684) );
  INV_X1 U13558 ( .A(n13456), .ZN(n10692) );
  AND2_X1 U13559 ( .A1(n10685), .A2(n10692), .ZN(n12962) );
  NAND2_X1 U13560 ( .A1(n10705), .A2(n12962), .ZN(n12812) );
  INV_X1 U13561 ( .A(n12947), .ZN(n10686) );
  NAND2_X1 U13562 ( .A1(n10702), .A2(n10686), .ZN(n10687) );
  NAND2_X1 U13563 ( .A1(n10687), .A2(n20080), .ZN(n10688) );
  AND3_X1 U13564 ( .A1(n10689), .A2(n12945), .A3(n10688), .ZN(n12792) );
  INV_X1 U13565 ( .A(n10690), .ZN(n10691) );
  AOI21_X1 U13566 ( .B1(n10692), .B2(n12325), .A(n10691), .ZN(n10694) );
  AND2_X1 U13567 ( .A1(n10694), .A2(n10693), .ZN(n10700) );
  NAND2_X1 U13568 ( .A1(n14060), .A2(n13440), .ZN(n10695) );
  NAND4_X1 U13569 ( .A1(n12792), .A2(n10700), .A3(n10696), .A4(n10695), .ZN(
        n10697) );
  NAND2_X1 U13570 ( .A1(n10705), .A2(n10697), .ZN(n12810) );
  AND2_X1 U13571 ( .A1(n10698), .A2(n14262), .ZN(n10699) );
  NOR2_X1 U13572 ( .A1(n12899), .A2(n12946), .ZN(n10701) );
  AND2_X1 U13573 ( .A1(n10702), .A2(n10701), .ZN(n10703) );
  NAND2_X1 U13574 ( .A1(n12948), .A2(n10703), .ZN(n12950) );
  INV_X1 U13575 ( .A(n12950), .ZN(n12638) );
  INV_X1 U13576 ( .A(n16009), .ZN(n16086) );
  INV_X1 U13577 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14489) );
  OR2_X1 U13578 ( .A1(n12810), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10706) );
  OR2_X1 U13579 ( .A1(n12330), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20036) );
  OR2_X1 U13580 ( .A1(n10705), .A2(n10704), .ZN(n14624) );
  INV_X1 U13581 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n20843) );
  INV_X1 U13582 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16095) );
  NOR3_X1 U13583 ( .A1(n20843), .A2(n16095), .A3(n10606), .ZN(n16068) );
  NAND3_X1 U13584 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n16068), .ZN(n16047) );
  INV_X1 U13585 ( .A(n16047), .ZN(n16043) );
  NAND2_X1 U13586 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16043), .ZN(
        n16055) );
  NOR2_X1 U13587 ( .A1(n10499), .A2(n16055), .ZN(n10707) );
  NOR2_X1 U13588 ( .A1(n20044), .A2(n20052), .ZN(n20039) );
  NAND2_X1 U13589 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20039), .ZN(
        n16054) );
  AOI21_X1 U13590 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n16052) );
  NOR2_X1 U13591 ( .A1(n16054), .A2(n16052), .ZN(n16044) );
  AND2_X1 U13592 ( .A1(n10707), .A2(n16044), .ZN(n14568) );
  NAND2_X1 U13593 ( .A1(n20034), .A2(n14568), .ZN(n10708) );
  NAND2_X1 U13594 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20054) );
  NOR2_X1 U13595 ( .A1(n20054), .A2(n16054), .ZN(n16065) );
  NAND2_X1 U13596 ( .A1(n16065), .A2(n10707), .ZN(n14567) );
  NAND2_X1 U13597 ( .A1(n10708), .A2(n14567), .ZN(n10711) );
  INV_X1 U13598 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16018) );
  INV_X1 U13599 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10709) );
  NOR4_X1 U13600 ( .A1(n10501), .A2(n14610), .A3(n16018), .A4(n10709), .ZN(
        n16015) );
  AND2_X1 U13601 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16015), .ZN(
        n10718) );
  NAND2_X1 U13602 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n10718), .ZN(
        n14570) );
  INV_X1 U13603 ( .A(n14570), .ZN(n10710) );
  AND3_X1 U13604 ( .A1(n10711), .A2(n20033), .A3(n10710), .ZN(n14602) );
  NOR2_X1 U13605 ( .A1(n14600), .A2(n14589), .ZN(n10712) );
  AOI21_X1 U13606 ( .B1(n14602), .B2(n10712), .A(n14601), .ZN(n14583) );
  AOI21_X1 U13607 ( .B1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(n16009), .ZN(n10713) );
  NOR2_X1 U13608 ( .A1(n14583), .A2(n10713), .ZN(n14562) );
  OAI21_X1 U13609 ( .B1(n14526), .B2(n16009), .A(n14562), .ZN(n14540) );
  NAND2_X1 U13610 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10714) );
  INV_X1 U13611 ( .A(n14601), .ZN(n16066) );
  OAI21_X1 U13612 ( .B1(n14540), .B2(n10714), .A(n16066), .ZN(n14521) );
  OAI21_X1 U13613 ( .B1(n14507), .B2(n14601), .A(n14521), .ZN(n14496) );
  AOI211_X1 U13614 ( .C1(n14499), .C2(n16086), .A(n14489), .B(n14496), .ZN(
        n14487) );
  NOR3_X1 U13615 ( .A1(n14487), .A2(n14601), .A3(n10512), .ZN(n10722) );
  INV_X1 U13616 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20718) );
  NOR2_X1 U13617 ( .A1(n20036), .A2(n20718), .ZN(n12336) );
  INV_X1 U13618 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20055) );
  NAND2_X1 U13619 ( .A1(n10715), .A2(n12812), .ZN(n20066) );
  NOR2_X1 U13620 ( .A1(n10716), .A2(n14567), .ZN(n13783) );
  NAND2_X1 U13621 ( .A1(n20066), .A2(n13783), .ZN(n14547) );
  NAND2_X1 U13622 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14568), .ZN(
        n13786) );
  OR2_X1 U13623 ( .A1(n20056), .A2(n13786), .ZN(n10717) );
  NAND2_X1 U13624 ( .A1(n14547), .A2(n10717), .ZN(n16013) );
  NAND2_X1 U13625 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n10718), .ZN(
        n10719) );
  NOR2_X1 U13626 ( .A1(n14571), .A2(n10719), .ZN(n10720) );
  NAND2_X1 U13627 ( .A1(n16013), .A2(n10720), .ZN(n14527) );
  OR3_X1 U13628 ( .A1(n14527), .A2(n14528), .A3(n14529), .ZN(n14508) );
  INV_X1 U13629 ( .A(n14508), .ZN(n14518) );
  NAND3_X1 U13630 ( .A1(n14518), .A2(n14507), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14488) );
  NOR3_X1 U13631 ( .A1(n14488), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14489), .ZN(n10721) );
  NOR2_X2 U13632 ( .A1(n10732), .A2(n16825), .ZN(n10770) );
  AOI22_X1 U13633 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10731) );
  AOI22_X1 U13634 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10730) );
  INV_X2 U13635 ( .A(n17103), .ZN(n15742) );
  AOI22_X1 U13636 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n15742), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10729) );
  AOI22_X1 U13637 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10728) );
  NAND4_X1 U13638 ( .A1(n10731), .A2(n10730), .A3(n10729), .A4(n10728), .ZN(
        n10740) );
  INV_X2 U13639 ( .A(n10097), .ZN(n17110) );
  AOI22_X1 U13640 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10738) );
  INV_X2 U13641 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n20898) );
  AOI22_X1 U13642 ( .A1(n17072), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17088), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10737) );
  INV_X2 U13643 ( .A(n9599), .ZN(n17109) );
  AOI22_X1 U13644 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10736) );
  INV_X2 U13645 ( .A(n10807), .ZN(n16910) );
  INV_X2 U13646 ( .A(n16910), .ZN(n17107) );
  AOI22_X1 U13647 ( .A1(n17107), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n15741), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10735) );
  NAND4_X1 U13648 ( .A1(n10738), .A2(n10737), .A3(n10736), .A4(n10735), .ZN(
        n10739) );
  AOI22_X1 U13649 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17081), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10745) );
  INV_X2 U13650 ( .A(n10760), .ZN(n17052) );
  INV_X4 U13651 ( .A(n17052), .ZN(n17088) );
  AOI22_X1 U13652 ( .A1(n17088), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10744) );
  AOI22_X1 U13653 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9616), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10743) );
  AOI22_X1 U13654 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n15742), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10742) );
  NAND4_X1 U13655 ( .A1(n10745), .A2(n10744), .A3(n10743), .A4(n10742), .ZN(
        n10751) );
  AOI22_X1 U13656 ( .A1(n17072), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10749) );
  INV_X2 U13657 ( .A(n10097), .ZN(n17053) );
  AOI22_X1 U13658 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17053), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10748) );
  AOI22_X1 U13659 ( .A1(n17107), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10747) );
  AOI22_X1 U13660 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10770), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10746) );
  NAND4_X1 U13661 ( .A1(n10749), .A2(n10748), .A3(n10747), .A4(n10746), .ZN(
        n10750) );
  AOI22_X1 U13662 ( .A1(n15741), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10755) );
  AOI22_X1 U13663 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9618), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10754) );
  AOI22_X1 U13664 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17088), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10753) );
  AOI22_X1 U13665 ( .A1(n17107), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n15742), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10752) );
  NAND4_X1 U13666 ( .A1(n10755), .A2(n10754), .A3(n10753), .A4(n10752), .ZN(
        n10759) );
  AOI22_X1 U13667 ( .A1(n17072), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10758) );
  AOI22_X1 U13668 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10757) );
  INV_X1 U13669 ( .A(n16940), .ZN(n10808) );
  AOI22_X1 U13670 ( .A1(n10770), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10808), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10756) );
  AOI22_X1 U13671 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10769) );
  INV_X2 U13672 ( .A(n16910), .ZN(n15747) );
  AOI22_X1 U13673 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n17089), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n15747), .ZN(n10768) );
  INV_X2 U13674 ( .A(n9599), .ZN(n17082) );
  AOI22_X1 U13675 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17072), .B1(
        n10808), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10765) );
  AOI22_X1 U13676 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10770), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10764) );
  AOI22_X1 U13677 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n9618), .B1(
        n10809), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10763) );
  AOI22_X1 U13678 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n9616), .ZN(n10762) );
  NAND4_X1 U13679 ( .A1(n10765), .A2(n10764), .A3(n10763), .A4(n10762), .ZN(
        n10766) );
  AOI22_X1 U13680 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n15741), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10780) );
  AOI22_X1 U13681 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17088), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10779) );
  INV_X4 U13682 ( .A(n10914), .ZN(n17108) );
  AOI22_X1 U13683 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10771) );
  OAI21_X1 U13684 ( .B1(n9617), .B2(n20794), .A(n10771), .ZN(n10777) );
  AOI22_X1 U13685 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17081), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10775) );
  AOI22_X1 U13686 ( .A1(n17072), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15747), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U13687 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U13688 ( .A1(n17067), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10772) );
  NAND4_X1 U13689 ( .A1(n10775), .A2(n10774), .A3(n10773), .A4(n10772), .ZN(
        n10776) );
  AOI211_X1 U13690 ( .C1(n17108), .C2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n10777), .B(n10776), .ZN(n10778) );
  NAND3_X1 U13691 ( .A1(n10780), .A2(n10779), .A3(n10778), .ZN(n11001) );
  NAND2_X1 U13692 ( .A1(n10817), .A2(n11001), .ZN(n10820) );
  AOI22_X1 U13693 ( .A1(n17107), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n15741), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10790) );
  AOI22_X1 U13694 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17053), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10789) );
  INV_X2 U13695 ( .A(n16940), .ZN(n17106) );
  AOI22_X1 U13696 ( .A1(n17106), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9618), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10781) );
  OAI21_X1 U13697 ( .B1(n9645), .B2(n20890), .A(n10781), .ZN(n10787) );
  AOI22_X1 U13698 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10785) );
  AOI22_X1 U13699 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17081), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10784) );
  AOI22_X1 U13700 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10783) );
  AOI22_X1 U13701 ( .A1(n17067), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17088), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10782) );
  NAND4_X1 U13702 ( .A1(n10785), .A2(n10784), .A3(n10783), .A4(n10782), .ZN(
        n10786) );
  AOI211_X1 U13703 ( .C1(n17072), .C2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n10787), .B(n10786), .ZN(n10788) );
  NAND3_X1 U13704 ( .A1(n10790), .A2(n10789), .A3(n10788), .ZN(n11002) );
  NAND2_X1 U13705 ( .A1(n10822), .A2(n11002), .ZN(n10826) );
  AOI22_X1 U13706 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10800) );
  AOI22_X1 U13707 ( .A1(n17072), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10799) );
  AOI22_X1 U13708 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15742), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10791) );
  OAI21_X1 U13709 ( .B1(n9599), .B2(n20912), .A(n10791), .ZN(n10797) );
  INV_X2 U13710 ( .A(n17052), .ZN(n17100) );
  AOI22_X1 U13711 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10795) );
  AOI22_X1 U13712 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10794) );
  AOI22_X1 U13713 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10793) );
  AOI22_X1 U13714 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n15747), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10792) );
  NAND4_X1 U13715 ( .A1(n10795), .A2(n10794), .A3(n10793), .A4(n10792), .ZN(
        n10796) );
  AOI211_X1 U13716 ( .C1(n17101), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n10797), .B(n10796), .ZN(n10798) );
  NAND2_X1 U13717 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16321) );
  INV_X1 U13718 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16320) );
  NOR2_X1 U13719 ( .A1(n16321), .A2(n16320), .ZN(n11036) );
  INV_X1 U13720 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18104) );
  AOI22_X1 U13721 ( .A1(n10770), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17053), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10801) );
  OAI21_X1 U13722 ( .B1(n9645), .B2(n18104), .A(n10801), .ZN(n10802) );
  INV_X1 U13723 ( .A(n10802), .ZN(n10806) );
  AOI22_X1 U13724 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10805) );
  AOI22_X1 U13725 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10804) );
  AOI22_X1 U13726 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10807), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10813) );
  AOI22_X1 U13727 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10808), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10812) );
  AOI22_X1 U13728 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10811) );
  AOI22_X1 U13729 ( .A1(n17072), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10809), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10810) );
  NAND2_X2 U13730 ( .A1(n9654), .A2(n10107), .ZN(n17763) );
  INV_X1 U13731 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18709) );
  NOR2_X1 U13732 ( .A1(n11000), .A2(n18709), .ZN(n10814) );
  INV_X1 U13733 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18061) );
  XNOR2_X1 U13734 ( .A(n18061), .B(n10816), .ZN(n17747) );
  INV_X1 U13735 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18031) );
  XNOR2_X1 U13736 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n10821), .ZN(
        n17722) );
  INV_X1 U13737 ( .A(n11002), .ZN(n17283) );
  XOR2_X1 U13738 ( .A(n17283), .B(n10822), .Z(n10823) );
  NOR2_X1 U13739 ( .A1(n10824), .A2(n10823), .ZN(n10825) );
  INV_X1 U13740 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18016) );
  XNOR2_X1 U13741 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n10827), .ZN(
        n17699) );
  INV_X1 U13742 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17694) );
  NAND2_X1 U13743 ( .A1(n10838), .A2(n18004), .ZN(n10837) );
  INV_X1 U13744 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17634) );
  INV_X1 U13745 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17939) );
  INV_X1 U13746 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17602) );
  NAND2_X1 U13747 ( .A1(n17590), .A2(n10102), .ZN(n10836) );
  NAND2_X1 U13748 ( .A1(n10836), .A2(n17677), .ZN(n10843) );
  INV_X1 U13749 ( .A(n10838), .ZN(n10839) );
  NAND2_X1 U13750 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17958) );
  INV_X1 U13751 ( .A(n17958), .ZN(n17922) );
  NAND2_X1 U13752 ( .A1(n17922), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17936) );
  NOR2_X1 U13753 ( .A1(n17936), .A2(n17939), .ZN(n17942) );
  INV_X1 U13754 ( .A(n17942), .ZN(n17905) );
  INV_X1 U13755 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17909) );
  NOR2_X1 U13756 ( .A1(n17905), .A2(n17909), .ZN(n17907) );
  NAND2_X1 U13757 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17907), .ZN(
        n17889) );
  NOR2_X1 U13758 ( .A1(n10835), .A2(n17889), .ZN(n17873) );
  NAND2_X1 U13759 ( .A1(n17607), .A2(n17873), .ZN(n10842) );
  NAND2_X1 U13760 ( .A1(n10842), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10841) );
  INV_X1 U13761 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n20793) );
  INV_X1 U13762 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n20867) );
  NAND2_X1 U13763 ( .A1(n10843), .A2(n10842), .ZN(n17492) );
  NOR2_X1 U13764 ( .A1(n20793), .A2(n20867), .ZN(n17551) );
  INV_X1 U13765 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17540) );
  INV_X1 U13766 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17522) );
  NOR2_X1 U13767 ( .A1(n17540), .A2(n17522), .ZN(n17844) );
  NAND3_X1 U13768 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n17844), .ZN(n17834) );
  INV_X1 U13769 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17833) );
  NOR2_X1 U13770 ( .A1(n17834), .A2(n17833), .ZN(n16336) );
  NAND3_X1 U13771 ( .A1(n17551), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n16336), .ZN(n11031) );
  INV_X1 U13772 ( .A(n11031), .ZN(n10973) );
  NAND2_X1 U13773 ( .A1(n17542), .A2(n17540), .ZN(n10844) );
  NOR2_X1 U13774 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n10844), .ZN(
        n17509) );
  INV_X1 U13775 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17511) );
  NAND2_X1 U13776 ( .A1(n17509), .A2(n17511), .ZN(n17494) );
  NAND2_X1 U13777 ( .A1(n10845), .A2(n10113), .ZN(n10846) );
  NAND2_X1 U13778 ( .A1(n17477), .A2(n10846), .ZN(n17466) );
  NAND2_X1 U13779 ( .A1(n17551), .A2(n17492), .ZN(n17507) );
  NAND2_X1 U13780 ( .A1(n16336), .A2(n17508), .ZN(n17478) );
  INV_X1 U13781 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17818) );
  NOR3_X1 U13782 ( .A1(n17465), .A2(n17478), .A3(n17818), .ZN(n17452) );
  INV_X1 U13783 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17797) );
  NAND2_X1 U13784 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17774) );
  NAND2_X1 U13785 ( .A1(n17564), .A2(n17774), .ZN(n10847) );
  NAND2_X1 U13786 ( .A1(n11036), .A2(n16345), .ZN(n10850) );
  NAND2_X1 U13787 ( .A1(n17564), .A2(n10850), .ZN(n15840) );
  INV_X1 U13788 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18708) );
  AOI22_X1 U13789 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17677), .B1(
        n17564), .B2(n18708), .ZN(n10851) );
  NOR2_X1 U13790 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18708), .ZN(
        n11044) );
  INV_X1 U13791 ( .A(n16339), .ZN(n17278) );
  AOI22_X1 U13792 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n15741), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10856) );
  AOI22_X1 U13793 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10855) );
  AOI22_X1 U13794 ( .A1(n17104), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10854) );
  AOI22_X1 U13795 ( .A1(n17067), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17088), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10853) );
  NAND4_X1 U13796 ( .A1(n10856), .A2(n10855), .A3(n10854), .A4(n10853), .ZN(
        n10862) );
  AOI22_X1 U13797 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10860) );
  BUF_X2 U13798 ( .A(n10867), .Z(n17117) );
  AOI22_X1 U13799 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10859) );
  AOI22_X1 U13800 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17087), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10858) );
  AOI22_X1 U13801 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10857) );
  NAND4_X1 U13802 ( .A1(n10860), .A2(n10859), .A3(n10858), .A4(n10857), .ZN(
        n10861) );
  AOI22_X1 U13803 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10866) );
  AOI22_X1 U13804 ( .A1(n17106), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10865) );
  AOI22_X1 U13805 ( .A1(n17072), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10864) );
  AOI22_X1 U13806 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10863) );
  NAND4_X1 U13807 ( .A1(n10866), .A2(n10865), .A3(n10864), .A4(n10863), .ZN(
        n10873) );
  AOI22_X1 U13808 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17101), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10871) );
  AOI22_X1 U13809 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17088), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10870) );
  AOI22_X1 U13810 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15741), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10869) );
  AOI22_X1 U13811 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17087), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10868) );
  NAND4_X1 U13812 ( .A1(n10871), .A2(n10870), .A3(n10869), .A4(n10868), .ZN(
        n10872) );
  NOR2_X1 U13813 ( .A1(n18750), .A2(n10981), .ZN(n10968) );
  AOI22_X1 U13814 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9616), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10877) );
  AOI22_X1 U13815 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17081), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10876) );
  AOI22_X1 U13816 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10875) );
  AOI22_X1 U13817 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n15742), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10874) );
  NAND4_X1 U13818 ( .A1(n10877), .A2(n10876), .A3(n10875), .A4(n10874), .ZN(
        n10883) );
  AOI22_X1 U13819 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17088), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10881) );
  AOI22_X1 U13820 ( .A1(n16928), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17072), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10880) );
  AOI22_X1 U13821 ( .A1(n15747), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9618), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10879) );
  AOI22_X1 U13822 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10878) );
  NAND4_X1 U13823 ( .A1(n10881), .A2(n10880), .A3(n10879), .A4(n10878), .ZN(
        n10882) );
  INV_X1 U13824 ( .A(n18127), .ZN(n10977) );
  NAND2_X1 U13825 ( .A1(n10968), .A2(n10977), .ZN(n10969) );
  AOI22_X1 U13826 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17081), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10892) );
  AOI22_X1 U13827 ( .A1(n16928), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10891) );
  INV_X1 U13828 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18122) );
  AOI22_X1 U13829 ( .A1(n17088), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10884) );
  OAI21_X1 U13830 ( .B1(n16910), .B2(n18122), .A(n10884), .ZN(n10890) );
  AOI22_X1 U13831 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10888) );
  AOI22_X1 U13832 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n15741), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10887) );
  AOI22_X1 U13833 ( .A1(n17106), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10886) );
  AOI22_X1 U13834 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17072), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10885) );
  NAND4_X1 U13835 ( .A1(n10888), .A2(n10887), .A3(n10886), .A4(n10885), .ZN(
        n10889) );
  AOI22_X1 U13836 ( .A1(n16928), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17088), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10902) );
  AOI22_X1 U13837 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17072), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10901) );
  INV_X2 U13838 ( .A(n9647), .ZN(n17066) );
  AOI22_X1 U13839 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10893) );
  OAI21_X1 U13840 ( .B1(n16910), .B2(n20890), .A(n10893), .ZN(n10899) );
  AOI22_X1 U13841 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10897) );
  AOI22_X1 U13842 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10896) );
  AOI22_X1 U13843 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9616), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10895) );
  AOI22_X1 U13844 ( .A1(n17067), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10894) );
  NAND4_X1 U13845 ( .A1(n10897), .A2(n10896), .A3(n10895), .A4(n10894), .ZN(
        n10898) );
  NAND2_X1 U13846 ( .A1(n18127), .A2(n17154), .ZN(n10934) );
  AOI22_X1 U13847 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10912) );
  AOI22_X1 U13848 ( .A1(n16928), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10911) );
  AOI22_X1 U13849 ( .A1(n17072), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17088), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10903) );
  OAI21_X1 U13850 ( .B1(n10097), .B2(n20912), .A(n10903), .ZN(n10909) );
  AOI22_X1 U13851 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15741), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10907) );
  AOI22_X1 U13852 ( .A1(n15747), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10906) );
  AOI22_X1 U13853 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10905) );
  AOI22_X1 U13854 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n15742), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10904) );
  NAND4_X1 U13855 ( .A1(n10907), .A2(n10906), .A3(n10905), .A4(n10904), .ZN(
        n10908) );
  NAND3_X2 U13856 ( .A1(n10912), .A2(n10911), .A3(n10910), .ZN(n17240) );
  AOI22_X1 U13857 ( .A1(n17107), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17081), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10923) );
  AOI22_X1 U13858 ( .A1(n15741), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9618), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10922) );
  AOI22_X1 U13859 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17110), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10913) );
  OAI21_X1 U13860 ( .B1(n10914), .B2(n20794), .A(n10913), .ZN(n10920) );
  AOI22_X1 U13861 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10918) );
  AOI22_X1 U13862 ( .A1(n17072), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10917) );
  AOI22_X1 U13863 ( .A1(n16928), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10916) );
  AOI22_X1 U13864 ( .A1(n17067), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17088), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10915) );
  NAND4_X1 U13865 ( .A1(n10918), .A2(n10917), .A3(n10916), .A4(n10915), .ZN(
        n10919) );
  AOI211_X1 U13866 ( .C1(n17117), .C2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n10920), .B(n10919), .ZN(n10921) );
  NAND3_X1 U13867 ( .A1(n10923), .A2(n10922), .A3(n10921), .ZN(n10936) );
  AOI21_X1 U13868 ( .B1(n10937), .B2(n10934), .A(n10995), .ZN(n10978) );
  AOI22_X1 U13869 ( .A1(n16928), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10927) );
  AOI22_X1 U13870 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9616), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10926) );
  AOI22_X1 U13871 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10925) );
  AOI22_X1 U13872 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10924) );
  NAND4_X1 U13873 ( .A1(n10927), .A2(n10926), .A3(n10925), .A4(n10924), .ZN(
        n10933) );
  AOI22_X1 U13874 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17088), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10931) );
  AOI22_X1 U13875 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9618), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10930) );
  AOI22_X1 U13876 ( .A1(n17072), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10929) );
  AOI22_X1 U13877 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17087), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10928) );
  NAND4_X1 U13878 ( .A1(n10931), .A2(n10930), .A3(n10929), .A4(n10928), .ZN(
        n10932) );
  NOR2_X1 U13879 ( .A1(n16776), .A2(n18750), .ZN(n10976) );
  NOR2_X1 U13880 ( .A1(n10976), .A2(n10981), .ZN(n10940) );
  NAND2_X1 U13881 ( .A1(n18124), .A2(n10977), .ZN(n10983) );
  NAND3_X1 U13882 ( .A1(n10978), .A2(n10940), .A3(n10983), .ZN(n10935) );
  INV_X1 U13883 ( .A(n15768), .ZN(n18534) );
  NOR2_X1 U13884 ( .A1(n18136), .A2(n18569), .ZN(n15858) );
  NAND2_X1 U13885 ( .A1(n18750), .A2(n16776), .ZN(n10975) );
  NOR2_X1 U13886 ( .A1(n15858), .A2(n10975), .ZN(n10985) );
  INV_X1 U13887 ( .A(n10935), .ZN(n10946) );
  INV_X1 U13888 ( .A(n10984), .ZN(n10944) );
  INV_X1 U13889 ( .A(n10945), .ZN(n10939) );
  AOI21_X1 U13890 ( .B1(n18109), .B2(n18101), .A(n18569), .ZN(n10938) );
  AOI21_X1 U13891 ( .B1(n10980), .B2(n10939), .A(n10938), .ZN(n10943) );
  NOR2_X1 U13892 ( .A1(n18136), .A2(n10945), .ZN(n10941) );
  OAI22_X1 U13893 ( .A1(n18119), .A2(n10941), .B1(n10945), .B2(n10940), .ZN(
        n10942) );
  NAND4_X1 U13894 ( .A1(n18114), .A2(n18119), .A3(n10984), .A4(n10945), .ZN(
        n10996) );
  AOI21_X1 U13895 ( .B1(n10946), .B2(n10988), .A(n10982), .ZN(n10947) );
  NOR2_X1 U13896 ( .A1(n10985), .A2(n10947), .ZN(n15761) );
  INV_X1 U13897 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18580) );
  OAI22_X1 U13898 ( .A1(n18717), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18580), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10956) );
  OAI22_X1 U13899 ( .A1(n9610), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n18575), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10961) );
  NAND2_X1 U13900 ( .A1(n18392), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10962) );
  NOR2_X1 U13901 ( .A1(n10961), .A2(n10962), .ZN(n10948) );
  OAI21_X1 U13902 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18717), .A(
        n10949), .ZN(n10950) );
  OAI22_X1 U13903 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18584), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n10950), .ZN(n10952) );
  NOR2_X1 U13904 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18584), .ZN(
        n10951) );
  NAND2_X1 U13905 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10950), .ZN(
        n10953) );
  AOI22_X1 U13906 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n10952), .B1(
        n10951), .B2(n10953), .ZN(n10960) );
  OAI21_X1 U13907 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18392), .A(
        n10962), .ZN(n10965) );
  NOR2_X1 U13908 ( .A1(n10961), .A2(n10965), .ZN(n10959) );
  AOI21_X1 U13909 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n10953), .A(
        n10952), .ZN(n10954) );
  AOI21_X1 U13910 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18584), .A(
        n10954), .ZN(n10963) );
  NAND2_X1 U13911 ( .A1(n10957), .A2(n10956), .ZN(n10955) );
  OAI211_X1 U13912 ( .C1(n10957), .C2(n10956), .A(n10960), .B(n10955), .ZN(
        n10966) );
  NAND2_X1 U13913 ( .A1(n10963), .A2(n10966), .ZN(n10958) );
  NAND2_X1 U13914 ( .A1(n18109), .A2(n17154), .ZN(n10986) );
  INV_X1 U13915 ( .A(n10986), .ZN(n10971) );
  XNOR2_X1 U13916 ( .A(n10962), .B(n10961), .ZN(n10964) );
  NOR2_X1 U13917 ( .A1(n10966), .A2(n10965), .ZN(n12342) );
  INV_X1 U13918 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18629) );
  NOR2_X2 U13919 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18618), .ZN(n18697) );
  OAI211_X1 U13920 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18629), .B(n18691), .ZN(n18748) );
  OAI21_X1 U13921 ( .B1(n18109), .B2(n15660), .A(n18748), .ZN(n10967) );
  NAND2_X1 U13922 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18751) );
  OAI21_X1 U13923 ( .B1(n10968), .B2(n10967), .A(n18751), .ZN(n16459) );
  OAI22_X1 U13924 ( .A1(n12342), .A2(n10969), .B1(n10971), .B2(n16459), .ZN(
        n10970) );
  AOI22_X1 U13925 ( .A1(n18531), .A2(n10971), .B1(n18536), .B2(n10970), .ZN(
        n10972) );
  INV_X1 U13926 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18710) );
  NAND2_X1 U13927 ( .A1(n18710), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18605) );
  NOR2_X1 U13928 ( .A1(n18605), .A2(n18762), .ZN(n18745) );
  INV_X1 U13929 ( .A(n18745), .ZN(n18600) );
  AOI21_X2 U13930 ( .B1(n15761), .B2(n10972), .A(n18600), .ZN(n18071) );
  NOR3_X2 U13931 ( .A1(n17278), .A2(n18534), .A3(n18086), .ZN(n17982) );
  NAND3_X1 U13932 ( .A1(n11036), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n18708), .ZN(n10998) );
  INV_X1 U13933 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17467) );
  NAND2_X1 U13934 ( .A1(n17942), .A2(n17644), .ZN(n17925) );
  NAND2_X1 U13935 ( .A1(n10973), .A2(n17824), .ZN(n17808) );
  INV_X1 U13936 ( .A(n17778), .ZN(n17424) );
  INV_X1 U13937 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15843) );
  NAND2_X1 U13938 ( .A1(n11036), .A2(n17778), .ZN(n16311) );
  OAI21_X1 U13939 ( .B1(n15843), .B2(n16311), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10974) );
  OAI21_X1 U13940 ( .B1(n10998), .B2(n17424), .A(n10974), .ZN(n12353) );
  INV_X1 U13941 ( .A(n12353), .ZN(n10999) );
  NAND2_X1 U13942 ( .A1(n15768), .A2(n17278), .ZN(n17995) );
  INV_X1 U13943 ( .A(n10975), .ZN(n17306) );
  INV_X1 U13944 ( .A(n18753), .ZN(n18764) );
  NOR2_X1 U13945 ( .A1(n18119), .A2(n10977), .ZN(n18544) );
  NAND3_X1 U13946 ( .A1(n18109), .A2(n10978), .A3(n18544), .ZN(n15762) );
  INV_X1 U13947 ( .A(n18566), .ZN(n18035) );
  AOI21_X1 U13948 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18058) );
  NAND3_X1 U13949 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17992) );
  NOR2_X1 U13950 ( .A1(n18058), .A2(n17992), .ZN(n17986) );
  INV_X1 U13951 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18019) );
  NOR3_X1 U13952 ( .A1(n17694), .A2(n18019), .A3(n18004), .ZN(n10979) );
  NAND2_X1 U13953 ( .A1(n17986), .A2(n10979), .ZN(n17904) );
  NAND2_X1 U13954 ( .A1(n17551), .A2(n17873), .ZN(n17552) );
  NOR2_X1 U13955 ( .A1(n17904), .A2(n17552), .ZN(n17864) );
  NAND2_X1 U13956 ( .A1(n16336), .A2(n17864), .ZN(n11040) );
  NAND2_X1 U13957 ( .A1(n18593), .A2(n15660), .ZN(n10991) );
  INV_X1 U13958 ( .A(n10996), .ZN(n10990) );
  NAND2_X1 U13959 ( .A1(n18109), .A2(n18114), .ZN(n10994) );
  NAND3_X1 U13960 ( .A1(n18750), .A2(n10984), .A3(n15658), .ZN(n10993) );
  NAND3_X1 U13961 ( .A1(n10993), .A2(n15759), .A3(n10991), .ZN(n11033) );
  AOI21_X1 U13962 ( .B1(n10987), .B2(n10986), .A(n10985), .ZN(n10989) );
  NAND2_X2 U13963 ( .A1(n18535), .A2(n10993), .ZN(n18559) );
  INV_X1 U13964 ( .A(n10994), .ZN(n18543) );
  AND2_X1 U13965 ( .A1(n15660), .A2(n10995), .ZN(n18541) );
  NAND2_X1 U13966 ( .A1(n18542), .A2(n10996), .ZN(n18548) );
  OAI21_X1 U13967 ( .B1(n18559), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18053), .ZN(n17991) );
  NAND2_X1 U13968 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18032) );
  NOR2_X1 U13969 ( .A1(n18032), .A2(n17992), .ZN(n17987) );
  NAND3_X1 U13970 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n17987), .ZN(n17978) );
  NOR2_X1 U13971 ( .A1(n18004), .A2(n17978), .ZN(n17921) );
  NAND2_X1 U13972 ( .A1(n17873), .A2(n17921), .ZN(n17863) );
  INV_X1 U13973 ( .A(n17551), .ZN(n17867) );
  OR2_X1 U13974 ( .A1(n17867), .A2(n17834), .ZN(n17827) );
  NOR2_X1 U13975 ( .A1(n17863), .A2(n17827), .ZN(n17771) );
  NAND2_X1 U13976 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17771), .ZN(
        n11037) );
  OAI22_X1 U13977 ( .A1(n18035), .A2(n11040), .B1(n17991), .B2(n11037), .ZN(
        n10997) );
  NAND2_X1 U13978 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17794) );
  INV_X1 U13979 ( .A(n17794), .ZN(n17773) );
  NAND2_X1 U13980 ( .A1(n10997), .A2(n17773), .ZN(n17796) );
  OR2_X1 U13981 ( .A1(n17774), .A2(n17796), .ZN(n15773) );
  OAI22_X1 U13982 ( .A1(n10999), .A2(n17995), .B1(n10998), .B2(n15773), .ZN(
        n11047) );
  NAND2_X1 U13983 ( .A1(n17763), .A2(n11000), .ZN(n11004) );
  NAND2_X1 U13984 ( .A1(n17291), .A2(n11004), .ZN(n11003) );
  NAND2_X1 U13985 ( .A1(n11003), .A2(n11001), .ZN(n11012) );
  NOR2_X1 U13986 ( .A1(n17285), .A2(n11012), .ZN(n11015) );
  NAND2_X1 U13987 ( .A1(n11015), .A2(n11002), .ZN(n11019) );
  NOR2_X1 U13988 ( .A1(n20927), .A2(n11019), .ZN(n11023) );
  NAND2_X1 U13989 ( .A1(n11023), .A2(n16339), .ZN(n11024) );
  XNOR2_X1 U13990 ( .A(n17288), .B(n11003), .ZN(n11010) );
  XOR2_X1 U13991 ( .A(n17291), .B(n11004), .Z(n11008) );
  NOR2_X1 U13992 ( .A1(n11008), .A2(n18061), .ZN(n11009) );
  INV_X1 U13993 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18727) );
  NOR2_X1 U13994 ( .A1(n17300), .A2(n18727), .ZN(n11007) );
  INV_X1 U13995 ( .A(n17763), .ZN(n11006) );
  NAND3_X1 U13996 ( .A1(n11006), .A2(n17300), .A3(n18727), .ZN(n11005) );
  OAI221_X1 U13997 ( .B1(n11007), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n11006), .C2(n17300), .A(n11005), .ZN(n17746) );
  XNOR2_X1 U13998 ( .A(n18061), .B(n11008), .ZN(n17745) );
  NOR2_X1 U13999 ( .A1(n17746), .A2(n17745), .ZN(n17744) );
  NOR2_X2 U14000 ( .A1(n11009), .A2(n17744), .ZN(n17735) );
  XNOR2_X1 U14001 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n11010), .ZN(
        n17734) );
  NOR2_X2 U14002 ( .A1(n17735), .A2(n17734), .ZN(n17733) );
  NOR2_X2 U14003 ( .A1(n11011), .A2(n17733), .ZN(n11013) );
  INV_X1 U14004 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18041) );
  NOR2_X1 U14005 ( .A1(n11013), .A2(n18041), .ZN(n11014) );
  XNOR2_X1 U14006 ( .A(n11012), .B(n17285), .ZN(n17720) );
  XNOR2_X1 U14007 ( .A(n18041), .B(n11013), .ZN(n17719) );
  NOR2_X2 U14008 ( .A1(n11014), .A2(n17718), .ZN(n11016) );
  XOR2_X1 U14009 ( .A(n11015), .B(n17283), .Z(n11017) );
  NOR2_X1 U14010 ( .A1(n11016), .A2(n11017), .ZN(n11018) );
  XNOR2_X1 U14011 ( .A(n11017), .B(n11016), .ZN(n17710) );
  NOR2_X2 U14012 ( .A1(n18016), .A2(n17710), .ZN(n17709) );
  NOR2_X2 U14013 ( .A1(n11018), .A2(n17709), .ZN(n11020) );
  XNOR2_X1 U14014 ( .A(n20927), .B(n11019), .ZN(n11021) );
  NOR2_X1 U14015 ( .A1(n11020), .A2(n11021), .ZN(n11022) );
  XNOR2_X1 U14016 ( .A(n11021), .B(n11020), .ZN(n17703) );
  XNOR2_X1 U14017 ( .A(n11023), .B(n16339), .ZN(n11026) );
  NAND2_X1 U14018 ( .A1(n11025), .A2(n11026), .ZN(n17689) );
  INV_X1 U14019 ( .A(n11024), .ZN(n11029) );
  OR2_X1 U14020 ( .A1(n11026), .A2(n11025), .ZN(n17690) );
  OAI21_X1 U14021 ( .B1(n11029), .B2(n11028), .A(n17690), .ZN(n11027) );
  NOR2_X2 U14022 ( .A1(n17675), .A2(n18004), .ZN(n17674) );
  NOR2_X2 U14023 ( .A1(n17954), .A2(n17905), .ZN(n17928) );
  NOR2_X2 U14024 ( .A1(n17602), .A2(n17599), .ZN(n17598) );
  NAND2_X1 U14025 ( .A1(n17811), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17450) );
  NOR2_X2 U14026 ( .A1(n17450), .A2(n17774), .ZN(n16318) );
  NAND3_X1 U14027 ( .A1(n16318), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n11036), .ZN(n11032) );
  XOR2_X1 U14028 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n11032), .Z(
        n12352) );
  INV_X1 U14029 ( .A(n11033), .ZN(n11035) );
  NAND2_X1 U14030 ( .A1(n18530), .A2(n18071), .ZN(n18079) );
  INV_X1 U14031 ( .A(n17883), .ZN(n17990) );
  NOR2_X1 U14032 ( .A1(n17990), .A2(n18086), .ZN(n18076) );
  INV_X1 U14033 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18688) );
  NOR2_X1 U14034 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18763) );
  INV_X1 U14035 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n12414) );
  NOR2_X1 U14036 ( .A1(n18688), .A2(n18069), .ZN(n12350) );
  INV_X1 U14037 ( .A(n11036), .ZN(n15842) );
  NAND2_X1 U14038 ( .A1(n18076), .A2(n15842), .ZN(n15844) );
  NOR2_X1 U14039 ( .A1(n17797), .A2(n17794), .ZN(n17786) );
  NAND2_X1 U14040 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17786), .ZN(
        n17775) );
  NOR2_X1 U14041 ( .A1(n18552), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18054) );
  AOI21_X1 U14042 ( .B1(n18566), .B2(n17775), .A(n18054), .ZN(n11042) );
  INV_X1 U14043 ( .A(n18552), .ZN(n18568) );
  NOR2_X1 U14044 ( .A1(n11037), .A2(n17775), .ZN(n11038) );
  NAND2_X1 U14045 ( .A1(n11038), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11039) );
  OAI21_X1 U14046 ( .B1(n18559), .B2(n18568), .A(n11039), .ZN(n11041) );
  NAND2_X1 U14047 ( .A1(n18069), .A2(n18086), .ZN(n18072) );
  NAND2_X1 U14048 ( .A1(n18566), .A2(n11040), .ZN(n17812) );
  NAND4_X1 U14049 ( .A1(n11042), .A2(n11041), .A3(n18072), .A4(n17812), .ZN(
        n16346) );
  NAND2_X1 U14050 ( .A1(n18069), .A2(n16346), .ZN(n15769) );
  AOI21_X1 U14051 ( .B1(n15844), .B2(n15769), .A(n18708), .ZN(n11043) );
  AOI211_X1 U14052 ( .C1(n11044), .C2(n18076), .A(n12350), .B(n11043), .ZN(
        n11045) );
  NAND2_X1 U14053 ( .A1(n12633), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11170) );
  INV_X1 U14054 ( .A(n11050), .ZN(n11564) );
  NAND2_X1 U14055 ( .A1(n11564), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11090) );
  XNOR2_X1 U14056 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14190) );
  INV_X2 U14057 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20652) );
  AOI21_X1 U14058 ( .B1(n11552), .B2(n14190), .A(n11556), .ZN(n11053) );
  NOR2_X2 U14059 ( .A1(n20105), .A2(n20652), .ZN(n11051) );
  NAND2_X1 U14060 ( .A1(n11400), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11052) );
  OAI211_X1 U14061 ( .C1(n11090), .C2(n10120), .A(n11053), .B(n11052), .ZN(
        n11054) );
  INV_X1 U14062 ( .A(n11054), .ZN(n11055) );
  NAND2_X1 U14063 ( .A1(n11556), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11078) );
  INV_X1 U14064 ( .A(n11057), .ZN(n11060) );
  INV_X1 U14065 ( .A(n11058), .ZN(n11059) );
  NAND2_X1 U14066 ( .A1(n11060), .A2(n11059), .ZN(n11061) );
  NAND2_X1 U14067 ( .A1(n11062), .A2(n11061), .ZN(n12986) );
  NAND2_X1 U14068 ( .A1(n12986), .A2(n11241), .ZN(n11066) );
  AOI22_X1 U14069 ( .A1(n11051), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20652), .ZN(n11064) );
  INV_X1 U14070 ( .A(n11090), .ZN(n11070) );
  NAND2_X1 U14071 ( .A1(n11070), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11063) );
  AND2_X1 U14072 ( .A1(n11064), .A2(n11063), .ZN(n11065) );
  NAND2_X1 U14073 ( .A1(n11066), .A2(n11065), .ZN(n12737) );
  INV_X1 U14074 ( .A(n11067), .ZN(n11068) );
  XNOR2_X1 U14075 ( .A(n11069), .B(n11068), .ZN(n20181) );
  NAND2_X1 U14076 ( .A1(n20181), .A2(n11241), .ZN(n11074) );
  AOI22_X1 U14077 ( .A1(n11051), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20652), .ZN(n11072) );
  NAND2_X1 U14078 ( .A1(n11070), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11071) );
  AND2_X1 U14079 ( .A1(n11072), .A2(n11071), .ZN(n11073) );
  NAND2_X1 U14080 ( .A1(n11074), .A2(n11073), .ZN(n12757) );
  OR2_X1 U14081 ( .A1(n20739), .A2(n20098), .ZN(n11075) );
  AND2_X1 U14082 ( .A1(n11075), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12756) );
  NAND2_X1 U14083 ( .A1(n12757), .A2(n12756), .ZN(n12755) );
  OR2_X1 U14084 ( .A1(n12757), .A2(n13444), .ZN(n11076) );
  NAND2_X1 U14085 ( .A1(n12755), .A2(n11076), .ZN(n12736) );
  NAND2_X1 U14086 ( .A1(n12737), .A2(n12736), .ZN(n12840) );
  NAND2_X1 U14087 ( .A1(n13379), .A2(n11241), .ZN(n11087) );
  INV_X1 U14088 ( .A(n11080), .ZN(n11079) );
  INV_X1 U14089 ( .A(n11092), .ZN(n11094) );
  INV_X1 U14090 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11081) );
  NAND2_X1 U14091 ( .A1(n11081), .A2(n11080), .ZN(n11082) );
  NAND2_X1 U14092 ( .A1(n11094), .A2(n11082), .ZN(n13508) );
  AOI22_X1 U14093 ( .A1(n13508), .A2(n11375), .B1(n11556), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11084) );
  NAND2_X1 U14094 ( .A1(n11400), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11083) );
  OAI211_X1 U14095 ( .C1(n11090), .C2(n9816), .A(n11084), .B(n11083), .ZN(
        n11085) );
  INV_X1 U14096 ( .A(n11085), .ZN(n11086) );
  NAND2_X1 U14097 ( .A1(n11087), .A2(n11086), .ZN(n13098) );
  NAND2_X1 U14098 ( .A1(n20652), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11089) );
  NAND2_X1 U14099 ( .A1(n11400), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11088) );
  OAI211_X1 U14100 ( .C1(n11090), .C2(n16116), .A(n11089), .B(n11088), .ZN(
        n11091) );
  NAND2_X1 U14101 ( .A1(n11091), .A2(n13444), .ZN(n11097) );
  INV_X1 U14102 ( .A(n11101), .ZN(n11107) );
  INV_X1 U14103 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11093) );
  NAND2_X1 U14104 ( .A1(n11094), .A2(n11093), .ZN(n11095) );
  NAND2_X1 U14105 ( .A1(n11107), .A2(n11095), .ZN(n20022) );
  NAND2_X1 U14106 ( .A1(n20022), .A2(n11375), .ZN(n11096) );
  NAND2_X1 U14107 ( .A1(n11097), .A2(n11096), .ZN(n11098) );
  OAI21_X1 U14108 ( .B1(n11105), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n11119), .ZN(n19937) );
  AOI22_X1 U14109 ( .A1(n19937), .A2(n11375), .B1(n11556), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11102) );
  OAI21_X1 U14110 ( .B1(n11118), .B2(n19997), .A(n11102), .ZN(n11103) );
  AOI21_X1 U14111 ( .B1(n11104), .B2(n11241), .A(n11103), .ZN(n14256) );
  INV_X1 U14112 ( .A(n14256), .ZN(n11115) );
  INV_X1 U14113 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n11111) );
  INV_X1 U14114 ( .A(n11105), .ZN(n11109) );
  INV_X1 U14115 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11106) );
  NAND2_X1 U14116 ( .A1(n11107), .A2(n11106), .ZN(n11108) );
  NAND2_X1 U14117 ( .A1(n11109), .A2(n11108), .ZN(n16008) );
  AOI22_X1 U14118 ( .A1(n16008), .A2(n11375), .B1(n11556), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11110) );
  OAI21_X1 U14119 ( .B1(n11118), .B2(n11111), .A(n11110), .ZN(n11112) );
  INV_X1 U14120 ( .A(n13166), .ZN(n11114) );
  NAND2_X1 U14121 ( .A1(n11115), .A2(n11114), .ZN(n11116) );
  NAND2_X1 U14122 ( .A1(n11117), .A2(n11241), .ZN(n11126) );
  INV_X1 U14123 ( .A(n11556), .ZN(n12987) );
  INV_X1 U14124 ( .A(n11119), .ZN(n11121) );
  INV_X1 U14125 ( .A(n11141), .ZN(n11120) );
  OAI21_X1 U14126 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n11121), .A(
        n11120), .ZN(n19927) );
  NAND2_X1 U14127 ( .A1(n19927), .A2(n11375), .ZN(n11122) );
  OAI21_X1 U14128 ( .B1(n11123), .B2(n12987), .A(n11122), .ZN(n11124) );
  AOI21_X1 U14129 ( .B1(n11400), .B2(P1_EAX_REG_7__SCAN_IN), .A(n11124), .ZN(
        n11125) );
  NAND2_X1 U14130 ( .A1(n11126), .A2(n11125), .ZN(n13206) );
  AOI22_X1 U14131 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10301), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11130) );
  AOI22_X1 U14132 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11516), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11129) );
  AOI22_X1 U14133 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11128) );
  AOI22_X1 U14134 ( .A1(n11539), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11127) );
  NAND4_X1 U14135 ( .A1(n11130), .A2(n11129), .A3(n11128), .A4(n11127), .ZN(
        n11136) );
  AOI22_X1 U14136 ( .A1(n10272), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11538), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11134) );
  AOI22_X1 U14137 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12958), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11133) );
  AOI22_X1 U14138 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11132) );
  AOI22_X1 U14139 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9619), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11131) );
  NAND4_X1 U14140 ( .A1(n11134), .A2(n11133), .A3(n11132), .A4(n11131), .ZN(
        n11135) );
  OAI21_X1 U14141 ( .B1(n11136), .B2(n11135), .A(n11241), .ZN(n11139) );
  NAND2_X1 U14142 ( .A1(n11400), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11138) );
  XNOR2_X1 U14143 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n11141), .ZN(
        n19911) );
  AOI22_X1 U14144 ( .A1(n11375), .A2(n19911), .B1(n11556), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11137) );
  XNOR2_X1 U14145 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n11167), .ZN(
        n19900) );
  INV_X1 U14146 ( .A(n19900), .ZN(n11156) );
  AOI22_X1 U14147 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10301), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11145) );
  AOI22_X1 U14148 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11515), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11144) );
  AOI22_X1 U14149 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11143) );
  AOI22_X1 U14150 ( .A1(n11540), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11539), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11142) );
  NAND4_X1 U14151 ( .A1(n11145), .A2(n11144), .A3(n11143), .A4(n11142), .ZN(
        n11151) );
  AOI22_X1 U14152 ( .A1(n10272), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11538), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11149) );
  AOI22_X1 U14153 ( .A1(n11487), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12958), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11148) );
  AOI22_X1 U14154 ( .A1(n11510), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11147) );
  AOI22_X1 U14155 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11146) );
  NAND4_X1 U14156 ( .A1(n11149), .A2(n11148), .A3(n11147), .A4(n11146), .ZN(
        n11150) );
  OAI21_X1 U14157 ( .B1(n11151), .B2(n11150), .A(n11241), .ZN(n11154) );
  NAND2_X1 U14158 ( .A1(n11400), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11153) );
  NAND2_X1 U14159 ( .A1(n11556), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11152) );
  NAND3_X1 U14160 ( .A1(n11154), .A2(n11153), .A3(n11152), .ZN(n11155) );
  AOI21_X1 U14161 ( .B1(n11156), .B2(n11375), .A(n11155), .ZN(n13464) );
  AOI22_X1 U14162 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11160) );
  AOI22_X1 U14163 ( .A1(n11538), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11516), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11159) );
  AOI22_X1 U14164 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11158) );
  AOI22_X1 U14165 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11157) );
  NAND4_X1 U14166 ( .A1(n11160), .A2(n11159), .A3(n11158), .A4(n11157), .ZN(
        n11166) );
  AOI22_X1 U14167 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12958), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11164) );
  AOI22_X1 U14168 ( .A1(n10301), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11163) );
  AOI22_X1 U14169 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11539), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11162) );
  AOI22_X1 U14170 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11161) );
  NAND4_X1 U14171 ( .A1(n11164), .A2(n11163), .A3(n11162), .A4(n11161), .ZN(
        n11165) );
  NOR2_X1 U14172 ( .A1(n11166), .A2(n11165), .ZN(n11171) );
  XNOR2_X1 U14173 ( .A(n11172), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14481) );
  NAND2_X1 U14174 ( .A1(n14481), .A2(n11375), .ZN(n11169) );
  AOI22_X1 U14175 ( .A1(n11051), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n11556), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11168) );
  OAI211_X1 U14176 ( .C1(n11171), .C2(n11170), .A(n11169), .B(n11168), .ZN(
        n13516) );
  NAND2_X1 U14177 ( .A1(n11400), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n11175) );
  OAI21_X1 U14178 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11173), .A(
        n11187), .ZN(n15987) );
  AOI22_X1 U14179 ( .A1(n11375), .A2(n15987), .B1(n11556), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11174) );
  NAND2_X1 U14180 ( .A1(n11175), .A2(n11174), .ZN(n13733) );
  AOI22_X1 U14181 ( .A1(n11538), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10301), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11179) );
  AOI22_X1 U14182 ( .A1(n11487), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12958), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11178) );
  AOI22_X1 U14183 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11177) );
  AOI22_X1 U14184 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11176) );
  NAND4_X1 U14185 ( .A1(n11179), .A2(n11178), .A3(n11177), .A4(n11176), .ZN(
        n11185) );
  AOI22_X1 U14186 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11183) );
  AOI22_X1 U14187 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11532), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11182) );
  AOI22_X1 U14188 ( .A1(n11539), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11181) );
  AOI22_X1 U14189 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11180) );
  NAND4_X1 U14190 ( .A1(n11183), .A2(n11182), .A3(n11181), .A4(n11180), .ZN(
        n11184) );
  OR2_X1 U14191 ( .A1(n11185), .A2(n11184), .ZN(n11186) );
  AND2_X1 U14192 ( .A1(n11241), .A2(n11186), .ZN(n13748) );
  AOI21_X1 U14193 ( .B1(n20864), .B2(n11187), .A(n11217), .ZN(n15975) );
  OR2_X1 U14194 ( .A1(n15975), .A2(n13444), .ZN(n11202) );
  AOI22_X1 U14195 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11191) );
  AOI22_X1 U14196 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n11509), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11190) );
  AOI22_X1 U14197 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n9615), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11189) );
  AOI22_X1 U14198 ( .A1(n11538), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11188) );
  NAND4_X1 U14199 ( .A1(n11191), .A2(n11190), .A3(n11189), .A4(n11188), .ZN(
        n11197) );
  AOI22_X1 U14200 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12958), .B1(
        n11487), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11195) );
  AOI22_X1 U14201 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10301), .B1(
        n11539), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11194) );
  AOI22_X1 U14202 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11532), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11193) );
  AOI22_X1 U14203 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11192) );
  NAND4_X1 U14204 ( .A1(n11195), .A2(n11194), .A3(n11193), .A4(n11192), .ZN(
        n11196) );
  OAI21_X1 U14205 ( .B1(n11197), .B2(n11196), .A(n11241), .ZN(n11200) );
  NAND2_X1 U14206 ( .A1(n11400), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n11199) );
  NAND2_X1 U14207 ( .A1(n11556), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11198) );
  AND3_X1 U14208 ( .A1(n11200), .A2(n11199), .A3(n11198), .ZN(n11201) );
  NAND2_X1 U14209 ( .A1(n11202), .A2(n11201), .ZN(n13768) );
  INV_X1 U14210 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n13757) );
  XNOR2_X1 U14211 ( .A(n13757), .B(n11217), .ZN(n14475) );
  AOI22_X1 U14212 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11206) );
  AOI22_X1 U14213 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11515), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11205) );
  AOI22_X1 U14214 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11204) );
  AOI22_X1 U14215 ( .A1(n11539), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11203) );
  NAND4_X1 U14216 ( .A1(n11206), .A2(n11205), .A3(n11204), .A4(n11203), .ZN(
        n11212) );
  AOI22_X1 U14217 ( .A1(n11538), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10301), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11210) );
  AOI22_X1 U14218 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12958), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11209) );
  AOI22_X1 U14219 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11208) );
  AOI22_X1 U14220 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(n9620), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11207) );
  NAND4_X1 U14221 ( .A1(n11210), .A2(n11209), .A3(n11208), .A4(n11207), .ZN(
        n11211) );
  OR2_X1 U14222 ( .A1(n11212), .A2(n11211), .ZN(n11213) );
  AOI22_X1 U14223 ( .A1(n11241), .A2(n11213), .B1(n11556), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11215) );
  NAND2_X1 U14224 ( .A1(n11400), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11214) );
  OAI211_X1 U14225 ( .C1(n14475), .C2(n13444), .A(n11215), .B(n11214), .ZN(
        n13751) );
  AND2_X1 U14226 ( .A1(n13768), .A2(n13751), .ZN(n11216) );
  XNOR2_X1 U14227 ( .A(n11232), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15922) );
  INV_X1 U14228 ( .A(n15922), .ZN(n13791) );
  AOI22_X1 U14229 ( .A1(n11538), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10301), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11221) );
  AOI22_X1 U14230 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11515), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11220) );
  AOI22_X1 U14231 ( .A1(n11540), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11219) );
  AOI22_X1 U14232 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11218) );
  NAND4_X1 U14233 ( .A1(n11221), .A2(n11220), .A3(n11219), .A4(n11218), .ZN(
        n11227) );
  AOI22_X1 U14234 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11225) );
  AOI22_X1 U14235 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12958), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11224) );
  AOI22_X1 U14236 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11539), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11223) );
  AOI22_X1 U14237 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9619), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11222) );
  NAND4_X1 U14238 ( .A1(n11225), .A2(n11224), .A3(n11223), .A4(n11222), .ZN(
        n11226) );
  OAI21_X1 U14239 ( .B1(n11227), .B2(n11226), .A(n11241), .ZN(n11230) );
  NAND2_X1 U14240 ( .A1(n11400), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11229) );
  NAND2_X1 U14241 ( .A1(n11556), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11228) );
  NAND3_X1 U14242 ( .A1(n11230), .A2(n11229), .A3(n11228), .ZN(n11231) );
  AOI21_X1 U14243 ( .B1(n13791), .B2(n11375), .A(n11231), .ZN(n13742) );
  INV_X1 U14244 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n15925) );
  XOR2_X1 U14245 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n11250), .Z(
        n15966) );
  INV_X1 U14246 ( .A(n15966), .ZN(n11248) );
  AOI22_X1 U14247 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10301), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11236) );
  AOI22_X1 U14248 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11474), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11235) );
  AOI22_X1 U14249 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11515), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11234) );
  AOI22_X1 U14250 ( .A1(n11538), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11233) );
  NAND4_X1 U14251 ( .A1(n11236), .A2(n11235), .A3(n11234), .A4(n11233), .ZN(
        n11243) );
  AOI22_X1 U14252 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12958), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11240) );
  AOI22_X1 U14253 ( .A1(n10272), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11539), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11239) );
  AOI22_X1 U14254 ( .A1(n11540), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11238) );
  AOI22_X1 U14255 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11237) );
  NAND4_X1 U14256 ( .A1(n11240), .A2(n11239), .A3(n11238), .A4(n11237), .ZN(
        n11242) );
  OAI21_X1 U14257 ( .B1(n11243), .B2(n11242), .A(n11241), .ZN(n11246) );
  NAND2_X1 U14258 ( .A1(n11400), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11245) );
  NAND2_X1 U14259 ( .A1(n11556), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11244) );
  NAND3_X1 U14260 ( .A1(n11246), .A2(n11245), .A3(n11244), .ZN(n11247) );
  AOI21_X1 U14261 ( .B1(n11248), .B2(n11375), .A(n11247), .ZN(n13802) );
  INV_X1 U14262 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n14460) );
  XNOR2_X1 U14263 ( .A(n11268), .B(n14460), .ZN(n14462) );
  NAND2_X1 U14264 ( .A1(n14462), .A2(n11375), .ZN(n11267) );
  AOI22_X1 U14265 ( .A1(n10301), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11532), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11254) );
  AOI22_X1 U14266 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11253) );
  AOI22_X1 U14267 ( .A1(n10272), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11539), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11252) );
  AOI22_X1 U14268 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11251) );
  NAND4_X1 U14269 ( .A1(n11254), .A2(n11253), .A3(n11252), .A4(n11251), .ZN(
        n11263) );
  AOI22_X1 U14270 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10300), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11260) );
  NAND2_X1 U14271 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11256) );
  NAND2_X1 U14272 ( .A1(n11538), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11255) );
  AND3_X1 U14273 ( .A1(n11256), .A2(n11255), .A3(n13444), .ZN(n11259) );
  AOI22_X1 U14274 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11258) );
  AOI22_X1 U14275 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9619), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11257) );
  NAND4_X1 U14276 ( .A1(n11260), .A2(n11259), .A3(n11258), .A4(n11257), .ZN(
        n11262) );
  INV_X1 U14277 ( .A(n14637), .ZN(n11261) );
  NAND2_X1 U14278 ( .A1(n11527), .A2(n13444), .ZN(n11370) );
  OAI21_X1 U14279 ( .B1(n11263), .B2(n11262), .A(n11370), .ZN(n11265) );
  AOI22_X1 U14280 ( .A1(n11051), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20652), .ZN(n11264) );
  NAND2_X1 U14281 ( .A1(n11265), .A2(n11264), .ZN(n11266) );
  NAND2_X1 U14282 ( .A1(n11267), .A2(n11266), .ZN(n14177) );
  XNOR2_X1 U14283 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11281), .ZN(
        n15958) );
  AOI22_X1 U14284 ( .A1(n11051), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n11556), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11280) );
  AOI22_X1 U14285 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10301), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11272) );
  AOI22_X1 U14286 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11532), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11271) );
  AOI22_X1 U14287 ( .A1(n11538), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11270) );
  AOI22_X1 U14288 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11269) );
  NAND4_X1 U14289 ( .A1(n11272), .A2(n11271), .A3(n11270), .A4(n11269), .ZN(
        n11278) );
  AOI22_X1 U14290 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10300), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11276) );
  AOI22_X1 U14291 ( .A1(n11540), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11275) );
  AOI22_X1 U14292 ( .A1(n10272), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11539), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11274) );
  AOI22_X1 U14293 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9619), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11273) );
  NAND4_X1 U14294 ( .A1(n11276), .A2(n11275), .A3(n11274), .A4(n11273), .ZN(
        n11277) );
  OAI21_X1 U14295 ( .B1(n11278), .B2(n11277), .A(n11549), .ZN(n11279) );
  OAI211_X1 U14296 ( .C1(n15958), .C2(n13444), .A(n11280), .B(n11279), .ZN(
        n14251) );
  INV_X1 U14297 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15906) );
  INV_X1 U14298 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11282) );
  XNOR2_X1 U14299 ( .A(n11315), .B(n11282), .ZN(n14451) );
  NAND2_X1 U14300 ( .A1(n14451), .A2(n11375), .ZN(n11298) );
  AOI22_X1 U14301 ( .A1(n11538), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10186), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11286) );
  AOI22_X1 U14302 ( .A1(n10272), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11285) );
  AOI22_X1 U14303 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11539), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11284) );
  AOI22_X1 U14304 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10409), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11283) );
  NAND4_X1 U14305 ( .A1(n11286), .A2(n11285), .A3(n11284), .A4(n11283), .ZN(
        n11294) );
  AOI22_X1 U14306 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9615), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11292) );
  AOI22_X1 U14307 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10300), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11291) );
  NAND2_X1 U14308 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11288) );
  NAND2_X1 U14309 ( .A1(n10301), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11287) );
  AND3_X1 U14310 ( .A1(n11288), .A2(n11287), .A3(n13444), .ZN(n11290) );
  AOI22_X1 U14311 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9619), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11289) );
  NAND4_X1 U14312 ( .A1(n11292), .A2(n11291), .A3(n11290), .A4(n11289), .ZN(
        n11293) );
  OAI21_X1 U14313 ( .B1(n11294), .B2(n11293), .A(n11370), .ZN(n11296) );
  AOI22_X1 U14314 ( .A1(n11051), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20652), .ZN(n11295) );
  NAND2_X1 U14315 ( .A1(n11296), .A2(n11295), .ZN(n11297) );
  NAND2_X1 U14316 ( .A1(n11298), .A2(n11297), .ZN(n14241) );
  AOI22_X1 U14317 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11303) );
  AOI22_X1 U14318 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11515), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11302) );
  AOI22_X1 U14319 ( .A1(n10301), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11301) );
  AOI22_X1 U14320 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10409), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11300) );
  NAND4_X1 U14321 ( .A1(n11303), .A2(n11302), .A3(n11301), .A4(n11300), .ZN(
        n11310) );
  AOI22_X1 U14322 ( .A1(n11487), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12958), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11308) );
  AOI22_X1 U14323 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11516), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11307) );
  AOI22_X1 U14324 ( .A1(n11538), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11539), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11306) );
  AOI22_X1 U14325 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10225), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11305) );
  NAND4_X1 U14326 ( .A1(n11308), .A2(n11307), .A3(n11306), .A4(n11305), .ZN(
        n11309) );
  NOR2_X1 U14327 ( .A1(n11310), .A2(n11309), .ZN(n11314) );
  NAND2_X1 U14328 ( .A1(n20652), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11311) );
  NAND2_X1 U14329 ( .A1(n13444), .A2(n11311), .ZN(n11312) );
  AOI21_X1 U14330 ( .B1(n11400), .B2(P1_EAX_REG_19__SCAN_IN), .A(n11312), .ZN(
        n11313) );
  OAI21_X1 U14331 ( .B1(n11527), .B2(n11314), .A(n11313), .ZN(n11322) );
  INV_X1 U14332 ( .A(n11353), .ZN(n11320) );
  INV_X1 U14333 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11318) );
  INV_X1 U14334 ( .A(n11316), .ZN(n11317) );
  NAND2_X1 U14335 ( .A1(n11318), .A2(n11317), .ZN(n11319) );
  NAND2_X1 U14336 ( .A1(n11320), .A2(n11319), .ZN(n15952) );
  NAND2_X1 U14337 ( .A1(n11322), .A2(n11321), .ZN(n14235) );
  AOI22_X1 U14338 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12958), .B1(
        n11515), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11328) );
  AOI21_X1 U14339 ( .B1(n11510), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A(
        n11375), .ZN(n11324) );
  NAND2_X1 U14340 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11323) );
  AND2_X1 U14341 ( .A1(n11324), .A2(n11323), .ZN(n11327) );
  AOI22_X1 U14342 ( .A1(n10272), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11326) );
  AOI22_X1 U14343 ( .A1(n11538), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11325) );
  NAND4_X1 U14344 ( .A1(n11328), .A2(n11327), .A3(n11326), .A4(n11325), .ZN(
        n11334) );
  AOI22_X1 U14345 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n11509), .B1(
        n11532), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11332) );
  AOI22_X1 U14346 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n9615), .B1(
        n10301), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11331) );
  AOI22_X1 U14347 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11330) );
  AOI22_X1 U14348 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n11533), .B1(
        n11539), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11329) );
  NAND4_X1 U14349 ( .A1(n11332), .A2(n11331), .A3(n11330), .A4(n11329), .ZN(
        n11333) );
  OR2_X1 U14350 ( .A1(n11334), .A2(n11333), .ZN(n11335) );
  NAND2_X1 U14351 ( .A1(n11370), .A2(n11335), .ZN(n11338) );
  AOI22_X1 U14352 ( .A1(n11051), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20652), .ZN(n11337) );
  INV_X1 U14353 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15883) );
  XNOR2_X1 U14354 ( .A(n11353), .B(n15883), .ZN(n15874) );
  AND2_X1 U14355 ( .A1(n15874), .A2(n11375), .ZN(n11336) );
  AOI21_X1 U14356 ( .B1(n11338), .B2(n11337), .A(n11336), .ZN(n14227) );
  AOI22_X1 U14357 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11342) );
  AOI22_X1 U14358 ( .A1(n11538), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10301), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11341) );
  AOI22_X1 U14359 ( .A1(n11532), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11515), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11340) );
  AOI22_X1 U14360 ( .A1(n11540), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11339) );
  NAND4_X1 U14361 ( .A1(n11342), .A2(n11341), .A3(n11340), .A4(n11339), .ZN(
        n11348) );
  AOI22_X1 U14362 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10300), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11346) );
  AOI22_X1 U14363 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11345) );
  AOI22_X1 U14364 ( .A1(n11539), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11344) );
  AOI22_X1 U14365 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n9620), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11343) );
  NAND4_X1 U14366 ( .A1(n11346), .A2(n11345), .A3(n11344), .A4(n11343), .ZN(
        n11347) );
  NOR2_X1 U14367 ( .A1(n11348), .A2(n11347), .ZN(n11352) );
  INV_X1 U14368 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20515) );
  OAI21_X1 U14369 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20515), .A(
        n20652), .ZN(n11349) );
  INV_X1 U14370 ( .A(n11349), .ZN(n11350) );
  AOI21_X1 U14371 ( .B1(n11400), .B2(P1_EAX_REG_21__SCAN_IN), .A(n11350), .ZN(
        n11351) );
  OAI21_X1 U14372 ( .B1(n11527), .B2(n11352), .A(n11351), .ZN(n11358) );
  INV_X1 U14373 ( .A(n11354), .ZN(n11355) );
  INV_X1 U14374 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15864) );
  NAND2_X1 U14375 ( .A1(n11355), .A2(n15864), .ZN(n11356) );
  NAND2_X1 U14376 ( .A1(n11403), .A2(n11356), .ZN(n15862) );
  AOI22_X1 U14377 ( .A1(n11538), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11474), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11362) );
  AOI22_X1 U14378 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10186), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11361) );
  AOI22_X1 U14379 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11539), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11360) );
  AOI22_X1 U14380 ( .A1(n11510), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10409), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11359) );
  NAND4_X1 U14381 ( .A1(n11362), .A2(n11361), .A3(n11360), .A4(n11359), .ZN(
        n11372) );
  AOI22_X1 U14382 ( .A1(n10301), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11532), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11369) );
  AOI22_X1 U14383 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10300), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11368) );
  NAND2_X1 U14384 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11365) );
  NAND2_X1 U14385 ( .A1(n10272), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11364) );
  AND3_X1 U14386 ( .A1(n11365), .A2(n11364), .A3(n13444), .ZN(n11367) );
  AOI22_X1 U14387 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11366) );
  NAND4_X1 U14388 ( .A1(n11369), .A2(n11368), .A3(n11367), .A4(n11366), .ZN(
        n11371) );
  OAI21_X1 U14389 ( .B1(n11372), .B2(n11371), .A(n11370), .ZN(n11374) );
  AOI22_X1 U14390 ( .A1(n11051), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20652), .ZN(n11373) );
  NAND2_X1 U14391 ( .A1(n11374), .A2(n11373), .ZN(n11377) );
  XNOR2_X1 U14392 ( .A(n11403), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14426) );
  NAND2_X1 U14393 ( .A1(n14426), .A2(n11375), .ZN(n11376) );
  NAND2_X1 U14394 ( .A1(n11377), .A2(n11376), .ZN(n14163) );
  AOI22_X1 U14395 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12958), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11381) );
  AOI22_X1 U14396 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11380) );
  AOI22_X1 U14397 ( .A1(n11538), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11539), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11379) );
  AOI22_X1 U14398 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9619), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11378) );
  NAND4_X1 U14399 ( .A1(n11381), .A2(n11380), .A3(n11379), .A4(n11378), .ZN(
        n11387) );
  AOI22_X1 U14400 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11385) );
  AOI22_X1 U14401 ( .A1(n11532), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11515), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11384) );
  AOI22_X1 U14402 ( .A1(n10301), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11383) );
  AOI22_X1 U14403 ( .A1(n11540), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11382) );
  NAND4_X1 U14404 ( .A1(n11385), .A2(n11384), .A3(n11383), .A4(n11382), .ZN(
        n11386) );
  NOR2_X1 U14405 ( .A1(n11387), .A2(n11386), .ZN(n11411) );
  AOI22_X1 U14406 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11391) );
  AOI22_X1 U14407 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12958), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11390) );
  AOI22_X1 U14408 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11389) );
  AOI22_X1 U14409 ( .A1(n11532), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11388) );
  NAND4_X1 U14410 ( .A1(n11391), .A2(n11390), .A3(n11389), .A4(n11388), .ZN(
        n11397) );
  AOI22_X1 U14411 ( .A1(n11538), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10301), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U14412 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11394) );
  AOI22_X1 U14413 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11539), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11393) );
  AOI22_X1 U14414 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11392) );
  NAND4_X1 U14415 ( .A1(n11395), .A2(n11394), .A3(n11393), .A4(n11392), .ZN(
        n11396) );
  NOR2_X1 U14416 ( .A1(n11397), .A2(n11396), .ZN(n11412) );
  XNOR2_X1 U14417 ( .A(n11411), .B(n11412), .ZN(n11402) );
  NAND2_X1 U14418 ( .A1(n20652), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11398) );
  NAND2_X1 U14419 ( .A1(n13444), .A2(n11398), .ZN(n11399) );
  AOI21_X1 U14420 ( .B1(n11400), .B2(P1_EAX_REG_23__SCAN_IN), .A(n11399), .ZN(
        n11401) );
  OAI21_X1 U14421 ( .B1(n11527), .B2(n11402), .A(n11401), .ZN(n11409) );
  INV_X1 U14422 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11405) );
  NAND2_X1 U14423 ( .A1(n11406), .A2(n11405), .ZN(n11407) );
  NAND2_X1 U14424 ( .A1(n11429), .A2(n11407), .ZN(n14419) );
  NAND2_X1 U14425 ( .A1(n11409), .A2(n11408), .ZN(n14152) );
  NOR2_X1 U14426 ( .A1(n11412), .A2(n11411), .ZN(n11444) );
  AOI22_X1 U14427 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11532), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11416) );
  AOI22_X1 U14428 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12958), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11415) );
  AOI22_X1 U14429 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11414) );
  AOI22_X1 U14430 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9619), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11413) );
  NAND4_X1 U14431 ( .A1(n11416), .A2(n11415), .A3(n11414), .A4(n11413), .ZN(
        n11422) );
  AOI22_X1 U14432 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11420) );
  AOI22_X1 U14433 ( .A1(n11538), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10301), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11419) );
  AOI22_X1 U14434 ( .A1(n11539), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11418) );
  INV_X1 U14435 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n20085) );
  AOI22_X1 U14436 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11417) );
  NAND4_X1 U14437 ( .A1(n11420), .A2(n11419), .A3(n11418), .A4(n11417), .ZN(
        n11421) );
  OR2_X1 U14438 ( .A1(n11422), .A2(n11421), .ZN(n11443) );
  INV_X1 U14439 ( .A(n11443), .ZN(n11423) );
  XNOR2_X1 U14440 ( .A(n11444), .B(n11423), .ZN(n11424) );
  NAND2_X1 U14441 ( .A1(n11424), .A2(n11549), .ZN(n11428) );
  INV_X1 U14442 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14410) );
  AOI21_X1 U14443 ( .B1(n14410), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11425) );
  AOI21_X1 U14444 ( .B1(n11400), .B2(P1_EAX_REG_24__SCAN_IN), .A(n11425), .ZN(
        n11427) );
  XNOR2_X1 U14445 ( .A(n11429), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14414) );
  AOI21_X1 U14446 ( .B1(n11428), .B2(n11427), .A(n11426), .ZN(n14135) );
  INV_X1 U14447 ( .A(n11431), .ZN(n11432) );
  INV_X1 U14448 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14124) );
  OAI21_X1 U14449 ( .B1(n11432), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n11465), .ZN(n14401) );
  AOI22_X1 U14450 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11538), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11436) );
  AOI22_X1 U14451 ( .A1(n11487), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12958), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11435) );
  AOI22_X1 U14452 ( .A1(n11510), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11434) );
  AOI22_X1 U14453 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9619), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11433) );
  NAND4_X1 U14454 ( .A1(n11436), .A2(n11435), .A3(n11434), .A4(n11433), .ZN(
        n11442) );
  AOI22_X1 U14455 ( .A1(n10272), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10301), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11440) );
  AOI22_X1 U14456 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11509), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11439) );
  AOI22_X1 U14457 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11515), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11438) );
  AOI22_X1 U14458 ( .A1(n11540), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11539), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11437) );
  NAND4_X1 U14459 ( .A1(n11440), .A2(n11439), .A3(n11438), .A4(n11437), .ZN(
        n11441) );
  NOR2_X1 U14460 ( .A1(n11442), .A2(n11441), .ZN(n11460) );
  NAND2_X1 U14461 ( .A1(n11444), .A2(n11443), .ZN(n11459) );
  XNOR2_X1 U14462 ( .A(n11460), .B(n11459), .ZN(n11447) );
  AOI21_X1 U14463 ( .B1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20652), .A(
        n11552), .ZN(n11446) );
  NAND2_X1 U14464 ( .A1(n11051), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n11445) );
  OAI211_X1 U14465 ( .C1(n11447), .C2(n11527), .A(n11446), .B(n11445), .ZN(
        n11448) );
  OAI21_X1 U14466 ( .B1(n13444), .B2(n14401), .A(n11448), .ZN(n14121) );
  NOR2_X2 U14467 ( .A1(n14119), .A2(n14121), .ZN(n14108) );
  AOI22_X1 U14468 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11452) );
  AOI22_X1 U14469 ( .A1(n11538), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10301), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11451) );
  AOI22_X1 U14470 ( .A1(n11539), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11450) );
  AOI22_X1 U14471 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10409), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11449) );
  NAND4_X1 U14472 ( .A1(n11452), .A2(n11451), .A3(n11450), .A4(n11449), .ZN(
        n11458) );
  AOI22_X1 U14473 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11532), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11456) );
  AOI22_X1 U14474 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12958), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11455) );
  AOI22_X1 U14475 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11454) );
  AOI22_X1 U14476 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11453) );
  NAND4_X1 U14477 ( .A1(n11456), .A2(n11455), .A3(n11454), .A4(n11453), .ZN(
        n11457) );
  OR2_X1 U14478 ( .A1(n11458), .A2(n11457), .ZN(n11481) );
  NOR2_X1 U14479 ( .A1(n11460), .A2(n11459), .ZN(n11482) );
  XOR2_X1 U14480 ( .A(n11481), .B(n11482), .Z(n11461) );
  NAND2_X1 U14481 ( .A1(n11461), .A2(n11549), .ZN(n11464) );
  INV_X1 U14482 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14389) );
  NOR2_X1 U14483 ( .A1(n14389), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11462) );
  AOI211_X1 U14484 ( .C1(n11400), .C2(P1_EAX_REG_26__SCAN_IN), .A(n11552), .B(
        n11462), .ZN(n11463) );
  XOR2_X1 U14485 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B(n11467), .Z(
        n14393) );
  AOI22_X1 U14486 ( .A1(n11464), .A2(n11463), .B1(n11552), .B2(n14393), .ZN(
        n14110) );
  INV_X1 U14487 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14099) );
  OAI21_X1 U14488 ( .B1(n11465), .B2(n14389), .A(n14099), .ZN(n11468) );
  AND2_X1 U14489 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11466) );
  NAND2_X1 U14490 ( .A1(n11468), .A2(n11502), .ZN(n14382) );
  AOI22_X1 U14491 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10301), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11473) );
  AOI22_X1 U14492 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12958), .B1(
        n11487), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11472) );
  AOI22_X1 U14493 ( .A1(n11538), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10186), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11471) );
  AOI22_X1 U14494 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9619), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11470) );
  NAND4_X1 U14495 ( .A1(n11473), .A2(n11472), .A3(n11471), .A4(n11470), .ZN(
        n11480) );
  AOI22_X1 U14496 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n9615), .B1(
        n11474), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11478) );
  AOI22_X1 U14497 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11515), .B1(
        n11532), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11477) );
  AOI22_X1 U14498 ( .A1(n10272), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11476) );
  AOI22_X1 U14499 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11539), .B1(
        n10409), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11475) );
  NAND4_X1 U14500 ( .A1(n11478), .A2(n11477), .A3(n11476), .A4(n11475), .ZN(
        n11479) );
  NOR2_X1 U14501 ( .A1(n11480), .A2(n11479), .ZN(n11499) );
  NAND2_X1 U14502 ( .A1(n11482), .A2(n11481), .ZN(n11498) );
  XNOR2_X1 U14503 ( .A(n11499), .B(n11498), .ZN(n11485) );
  AOI21_X1 U14504 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20652), .A(
        n11552), .ZN(n11484) );
  NAND2_X1 U14505 ( .A1(n11051), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n11483) );
  OAI211_X1 U14506 ( .C1(n11485), .C2(n11527), .A(n11484), .B(n11483), .ZN(
        n11486) );
  OAI21_X1 U14507 ( .B1(n13444), .B2(n14382), .A(n11486), .ZN(n14096) );
  AOI22_X1 U14508 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11532), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11491) );
  AOI22_X1 U14509 ( .A1(n11487), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12958), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11490) );
  AOI22_X1 U14510 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11489) );
  AOI22_X1 U14511 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11488) );
  NAND4_X1 U14512 ( .A1(n11491), .A2(n11490), .A3(n11489), .A4(n11488), .ZN(
        n11497) );
  AOI22_X1 U14513 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11495) );
  AOI22_X1 U14514 ( .A1(n10278), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10301), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11494) );
  AOI22_X1 U14515 ( .A1(n11539), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11493) );
  INV_X1 U14516 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20097) );
  AOI22_X1 U14517 ( .A1(n11540), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10409), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11492) );
  NAND4_X1 U14518 ( .A1(n11495), .A2(n11494), .A3(n11493), .A4(n11492), .ZN(
        n11496) );
  OR2_X1 U14519 ( .A1(n11497), .A2(n11496), .ZN(n11523) );
  NOR2_X1 U14520 ( .A1(n11499), .A2(n11498), .ZN(n11524) );
  XOR2_X1 U14521 ( .A(n11523), .B(n11524), .Z(n11500) );
  NAND2_X1 U14522 ( .A1(n11500), .A2(n11549), .ZN(n11505) );
  INV_X1 U14523 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n20810) );
  NOR2_X1 U14524 ( .A1(n20810), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11501) );
  AOI211_X1 U14525 ( .C1(n11400), .C2(P1_EAX_REG_28__SCAN_IN), .A(n11552), .B(
        n11501), .ZN(n11504) );
  NAND2_X1 U14526 ( .A1(n11502), .A2(n20810), .ZN(n11503) );
  AOI22_X1 U14527 ( .A1(n11505), .A2(n11504), .B1(n11552), .B2(n14377), .ZN(
        n14083) );
  INV_X1 U14528 ( .A(n11507), .ZN(n11508) );
  INV_X1 U14529 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11506) );
  OAI21_X1 U14530 ( .B1(n11508), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n12334), .ZN(n14365) );
  AOI22_X1 U14531 ( .A1(n11487), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12958), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11514) );
  AOI22_X1 U14532 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11513) );
  AOI22_X1 U14533 ( .A1(n10301), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11512) );
  AOI22_X1 U14534 ( .A1(n11532), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10225), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11511) );
  NAND4_X1 U14535 ( .A1(n11514), .A2(n11513), .A3(n11512), .A4(n11511), .ZN(
        n11522) );
  AOI22_X1 U14536 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11520) );
  AOI22_X1 U14537 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11515), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11519) );
  AOI22_X1 U14538 ( .A1(n11538), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11539), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11518) );
  AOI22_X1 U14539 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10409), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11517) );
  NAND4_X1 U14540 ( .A1(n11520), .A2(n11519), .A3(n11518), .A4(n11517), .ZN(
        n11521) );
  NOR2_X1 U14541 ( .A1(n11522), .A2(n11521), .ZN(n11531) );
  NAND2_X1 U14542 ( .A1(n11524), .A2(n11523), .ZN(n11530) );
  XNOR2_X1 U14543 ( .A(n11531), .B(n11530), .ZN(n11528) );
  AOI21_X1 U14544 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20652), .A(
        n11552), .ZN(n11526) );
  NAND2_X1 U14545 ( .A1(n11051), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n11525) );
  OAI211_X1 U14546 ( .C1(n11528), .C2(n11527), .A(n11526), .B(n11525), .ZN(
        n11529) );
  OAI21_X1 U14547 ( .B1(n13444), .B2(n14365), .A(n11529), .ZN(n14074) );
  NOR2_X1 U14548 ( .A1(n11531), .A2(n11530), .ZN(n11548) );
  AOI22_X1 U14549 ( .A1(n9615), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11532), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11537) );
  AOI22_X1 U14550 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12958), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U14551 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11510), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11535) );
  AOI22_X1 U14552 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9619), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11534) );
  NAND4_X1 U14553 ( .A1(n11537), .A2(n11536), .A3(n11535), .A4(n11534), .ZN(
        n11546) );
  AOI22_X1 U14554 ( .A1(n10161), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10272), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11544) );
  AOI22_X1 U14555 ( .A1(n11538), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10301), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11543) );
  AOI22_X1 U14556 ( .A1(n11540), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11539), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11542) );
  AOI22_X1 U14557 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10409), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11541) );
  NAND4_X1 U14558 ( .A1(n11544), .A2(n11543), .A3(n11542), .A4(n11541), .ZN(
        n11545) );
  NOR2_X1 U14559 ( .A1(n11546), .A2(n11545), .ZN(n11547) );
  XNOR2_X1 U14560 ( .A(n11548), .B(n11547), .ZN(n11550) );
  NAND2_X1 U14561 ( .A1(n11550), .A2(n11549), .ZN(n11555) );
  INV_X1 U14562 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n20880) );
  OAI21_X1 U14563 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20880), .A(n13444), 
        .ZN(n11551) );
  AOI21_X1 U14564 ( .B1(n11400), .B2(P1_EAX_REG_30__SCAN_IN), .A(n11551), .ZN(
        n11554) );
  XNOR2_X1 U14565 ( .A(n12334), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14357) );
  AOI21_X1 U14566 ( .B1(n11555), .B2(n11554), .A(n11553), .ZN(n14057) );
  AOI22_X1 U14567 ( .A1(n11051), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n11556), .ZN(n11557) );
  XNOR2_X2 U14568 ( .A(n11559), .B(n11558), .ZN(n14043) );
  NAND2_X1 U14569 ( .A1(n12632), .A2(n12624), .ZN(n12949) );
  OAI21_X1 U14570 ( .B1(n12703), .B2(n12626), .A(n12949), .ZN(n11560) );
  NAND2_X1 U14571 ( .A1(n12800), .A2(n11560), .ZN(n12803) );
  INV_X1 U14572 ( .A(n11561), .ZN(n16113) );
  NAND3_X1 U14573 ( .A1(n12639), .A2(n16113), .A3(n20659), .ZN(n12795) );
  NAND3_X1 U14574 ( .A1(n12765), .A2(n12635), .A3(n20098), .ZN(n12759) );
  OR2_X1 U14575 ( .A1(n9655), .A2(n12759), .ZN(n11562) );
  NAND2_X1 U14576 ( .A1(n14043), .A2(n10095), .ZN(n11578) );
  NOR4_X1 U14577 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n11568) );
  NOR4_X1 U14578 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_17__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n11567) );
  NOR4_X1 U14579 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(
        P1_ADDRESS_REG_6__SCAN_IN), .A3(P1_ADDRESS_REG_5__SCAN_IN), .A4(
        P1_ADDRESS_REG_4__SCAN_IN), .ZN(n11566) );
  NOR4_X1 U14580 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(
        P1_ADDRESS_REG_10__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n11565) );
  AND4_X1 U14581 ( .A1(n11568), .A2(n11567), .A3(n11566), .A4(n11565), .ZN(
        n11573) );
  NOR4_X1 U14582 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_2__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n11571) );
  NOR4_X1 U14583 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_22__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n11570) );
  NOR4_X1 U14584 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n11569) );
  INV_X1 U14585 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20671) );
  AND4_X1 U14586 ( .A1(n11571), .A2(n11570), .A3(n11569), .A4(n20671), .ZN(
        n11572) );
  NAND2_X1 U14587 ( .A1(n11573), .A2(n11572), .ZN(n11574) );
  AND2_X2 U14588 ( .A1(n11574), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n13387)
         );
  INV_X1 U14589 ( .A(n13387), .ZN(n13389) );
  AOI22_X1 U14590 ( .A1(n14345), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14342), .ZN(n11577) );
  INV_X1 U14591 ( .A(n11575), .ZN(n11576) );
  INV_X1 U14592 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16358) );
  NAND2_X1 U14593 ( .A1(n11578), .A2(n10115), .ZN(P1_U2873) );
  INV_X1 U14594 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16212) );
  INV_X1 U14595 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19128) );
  NAND2_X1 U14596 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n11618), .ZN(
        n11617) );
  INV_X1 U14597 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16199) );
  INV_X1 U14598 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16205) );
  OR2_X1 U14599 ( .A1(n16199), .A2(n16205), .ZN(n11579) );
  INV_X1 U14600 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11580) );
  INV_X1 U14601 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18886) );
  NOR2_X1 U14602 ( .A1(n11580), .A2(n18886), .ZN(n11611) );
  AND2_X1 U14603 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n11611), .ZN(
        n11581) );
  INV_X1 U14604 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11610) );
  AND2_X1 U14605 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11582) );
  INV_X1 U14606 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15233) );
  INV_X1 U14607 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15206) );
  NAND2_X1 U14608 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n11603), .ZN(
        n11602) );
  INV_X1 U14609 ( .A(n11602), .ZN(n11583) );
  INV_X1 U14610 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15172) );
  AND2_X1 U14611 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11592) );
  AND2_X1 U14612 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n11592), .ZN(
        n11584) );
  INV_X1 U14613 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n11585) );
  XNOR2_X1 U14614 ( .A(n11594), .B(n11585), .ZN(n14662) );
  XNOR2_X1 U14615 ( .A(n11586), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14035) );
  INV_X1 U14616 ( .A(n14035), .ZN(n11588) );
  NAND2_X1 U14617 ( .A1(n11591), .A2(n11592), .ZN(n11596) );
  INV_X1 U14618 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15142) );
  NAND2_X1 U14619 ( .A1(n11596), .A2(n15142), .ZN(n11593) );
  AND2_X1 U14620 ( .A1(n11594), .A2(n11593), .ZN(n15144) );
  AND2_X1 U14621 ( .A1(n11591), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11597) );
  OR2_X1 U14622 ( .A1(n11597), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11595) );
  NAND2_X1 U14623 ( .A1(n11596), .A2(n11595), .ZN(n13983) );
  INV_X1 U14624 ( .A(n13983), .ZN(n12375) );
  INV_X1 U14625 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15151) );
  INV_X1 U14626 ( .A(n11591), .ZN(n11598) );
  AOI21_X1 U14627 ( .B1(n15151), .B2(n11598), .A(n11597), .ZN(n15154) );
  NOR2_X1 U14628 ( .A1(n9695), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11599) );
  AOI21_X1 U14629 ( .B1(n15172), .B2(n11600), .A(n9695), .ZN(n15170) );
  OAI21_X1 U14630 ( .B1(n11601), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n11600), .ZN(n15179) );
  INV_X1 U14631 ( .A(n15179), .ZN(n16135) );
  INV_X1 U14632 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n20877) );
  AOI21_X1 U14633 ( .B1(n11602), .B2(n20877), .A(n11601), .ZN(n15188) );
  OAI21_X1 U14634 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n11603), .A(
        n11602), .ZN(n16166) );
  INV_X1 U14635 ( .A(n16166), .ZN(n15794) );
  AOI21_X1 U14636 ( .B1(n15206), .B2(n11605), .A(n11603), .ZN(n15208) );
  OAI21_X1 U14637 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n11604), .A(
        n11605), .ZN(n15222) );
  INV_X1 U14638 ( .A(n15222), .ZN(n18800) );
  AOI21_X1 U14639 ( .B1(n15233), .B2(n11608), .A(n11604), .ZN(n18810) );
  NAND2_X1 U14640 ( .A1(n11606), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11607) );
  INV_X1 U14641 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18819) );
  NAND2_X1 U14642 ( .A1(n11607), .A2(n18819), .ZN(n11609) );
  NAND2_X1 U14643 ( .A1(n11609), .A2(n11608), .ZN(n18818) );
  AOI21_X1 U14644 ( .B1(n11610), .B2(n11629), .A(n11606), .ZN(n18844) );
  INV_X1 U14645 ( .A(n11612), .ZN(n11627) );
  NOR2_X1 U14646 ( .A1(n18886), .A2(n11627), .ZN(n11626) );
  AND2_X1 U14647 ( .A1(n11612), .A2(n11611), .ZN(n11630) );
  INV_X1 U14648 ( .A(n11630), .ZN(n11613) );
  OAI21_X1 U14649 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n11626), .A(
        n11613), .ZN(n18865) );
  INV_X1 U14650 ( .A(n18865), .ZN(n11628) );
  OAI21_X1 U14651 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n11614), .A(
        n11627), .ZN(n18888) );
  INV_X1 U14652 ( .A(n18888), .ZN(n11625) );
  NOR2_X1 U14653 ( .A1(n16205), .A2(n11621), .ZN(n11623) );
  AOI21_X1 U14654 ( .B1(n16205), .B2(n11621), .A(n11623), .ZN(n18916) );
  AOI21_X1 U14655 ( .B1(n16212), .B2(n11619), .A(n11622), .ZN(n16206) );
  AOI21_X1 U14656 ( .B1(n20876), .B2(n11617), .A(n11620), .ZN(n16213) );
  AOI21_X1 U14657 ( .B1(n19128), .B2(n11615), .A(n11618), .ZN(n19117) );
  AOI21_X1 U14658 ( .B1(n13130), .B2(n12904), .A(n11616), .ZN(n12903) );
  AOI22_X1 U14659 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n11587), .ZN(n13196) );
  AOI22_X1 U14660 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n13130), .B2(n11587), .ZN(
        n13125) );
  NAND2_X1 U14661 ( .A1(n13196), .A2(n13125), .ZN(n13124) );
  NOR2_X1 U14662 ( .A1(n12903), .A2(n13124), .ZN(n13080) );
  OAI21_X1 U14663 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11616), .A(
        n11615), .ZN(n13369) );
  NAND2_X1 U14664 ( .A1(n13080), .A2(n13369), .ZN(n18968) );
  NOR2_X1 U14665 ( .A1(n19117), .A2(n18968), .ZN(n18944) );
  OAI21_X1 U14666 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n11618), .A(
        n11617), .ZN(n18947) );
  NAND2_X1 U14667 ( .A1(n18944), .A2(n18947), .ZN(n12922) );
  NOR2_X1 U14668 ( .A1(n16213), .A2(n12922), .ZN(n13112) );
  OAI21_X1 U14669 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n11620), .A(
        n11619), .ZN(n15292) );
  NAND2_X1 U14670 ( .A1(n13112), .A2(n15292), .ZN(n13143) );
  NOR2_X1 U14671 ( .A1(n16206), .A2(n13143), .ZN(n18932) );
  OAI21_X1 U14672 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n11622), .A(
        n11621), .ZN(n18934) );
  NAND2_X1 U14673 ( .A1(n18932), .A2(n18934), .ZN(n18915) );
  NOR2_X1 U14674 ( .A1(n18916), .A2(n18915), .ZN(n18910) );
  INV_X1 U14675 ( .A(n11623), .ZN(n11624) );
  AOI21_X1 U14676 ( .B1(n16199), .B2(n11624), .A(n11614), .ZN(n16191) );
  INV_X1 U14677 ( .A(n16191), .ZN(n18913) );
  NAND2_X1 U14678 ( .A1(n18910), .A2(n18913), .ZN(n18887) );
  NOR2_X1 U14679 ( .A1(n11625), .A2(n18887), .ZN(n18878) );
  AOI21_X1 U14680 ( .B1(n18886), .B2(n11627), .A(n11626), .ZN(n18880) );
  INV_X1 U14681 ( .A(n18880), .ZN(n15278) );
  NAND2_X1 U14682 ( .A1(n18878), .A2(n15278), .ZN(n18863) );
  NOR2_X1 U14683 ( .A1(n11628), .A2(n18863), .ZN(n18853) );
  OAI21_X1 U14684 ( .B1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n11630), .A(
        n11629), .ZN(n18854) );
  NAND2_X1 U14685 ( .A1(n18853), .A2(n18854), .ZN(n18842) );
  NOR2_X1 U14686 ( .A1(n18844), .A2(n18842), .ZN(n18832) );
  XNOR2_X1 U14687 ( .A(n11606), .B(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n18841) );
  NAND2_X1 U14688 ( .A1(n18832), .A2(n18841), .ZN(n18830) );
  NAND2_X1 U14689 ( .A1(n12901), .A2(n18830), .ZN(n18817) );
  NOR2_X1 U14690 ( .A1(n9927), .A2(n18799), .ZN(n12389) );
  NOR2_X1 U14691 ( .A1(n15208), .A2(n12389), .ZN(n12388) );
  NOR2_X1 U14692 ( .A1(n9927), .A2(n12388), .ZN(n15792) );
  NOR2_X1 U14693 ( .A1(n15794), .A2(n15792), .ZN(n15793) );
  NOR2_X1 U14694 ( .A1(n9927), .A2(n15793), .ZN(n12401) );
  NOR2_X1 U14695 ( .A1(n15188), .A2(n12401), .ZN(n12400) );
  NOR2_X1 U14696 ( .A1(n9927), .A2(n12400), .ZN(n16134) );
  NOR2_X1 U14697 ( .A1(n16135), .A2(n16134), .ZN(n16133) );
  NOR2_X1 U14698 ( .A1(n9927), .A2(n16133), .ZN(n14734) );
  NOR2_X1 U14699 ( .A1(n9927), .A2(n14694), .ZN(n12373) );
  NOR2_X1 U14700 ( .A1(n12375), .A2(n12373), .ZN(n12374) );
  INV_X1 U14701 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n12437) );
  NOR4_X4 U14702 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .A4(n12437), .ZN(n18951) );
  AOI22_X1 U14703 ( .A1(n11754), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14903), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11633) );
  INV_X1 U14704 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11631) );
  INV_X2 U14705 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11737) );
  AND2_X4 U14706 ( .A1(n11936), .A2(n11737), .ZN(n14756) );
  AOI22_X1 U14707 ( .A1(n11756), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11635) );
  AOI22_X1 U14708 ( .A1(n11753), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11634) );
  NAND2_X1 U14709 ( .A1(n11636), .A2(n10112), .ZN(n11644) );
  AOI22_X1 U14710 ( .A1(n11754), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14903), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11639) );
  AOI22_X1 U14711 ( .A1(n11753), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11638) );
  AND3_X1 U14712 ( .A1(n11639), .A2(n11638), .A3(n11637), .ZN(n11642) );
  AOI22_X1 U14713 ( .A1(n11756), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9603), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11641) );
  AOI22_X1 U14714 ( .A1(n14756), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11640) );
  NAND3_X1 U14715 ( .A1(n11642), .A2(n11641), .A3(n11640), .ZN(n11643) );
  AOI22_X1 U14716 ( .A1(n11753), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11650) );
  AOI22_X1 U14717 ( .A1(n11756), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9603), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11648) );
  AOI22_X1 U14718 ( .A1(n11754), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14903), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11647) );
  NAND4_X1 U14719 ( .A1(n11650), .A2(n11649), .A3(n11648), .A4(n11647), .ZN(
        n11657) );
  AOI22_X1 U14720 ( .A1(n11754), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14903), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11652) );
  AOI22_X1 U14721 ( .A1(n11753), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11651) );
  AOI22_X1 U14722 ( .A1(n11756), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11654) );
  AOI22_X1 U14723 ( .A1(n14756), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9606), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11653) );
  NAND2_X1 U14724 ( .A1(n11800), .A2(n11792), .ZN(n11791) );
  AOI22_X1 U14725 ( .A1(n11756), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9603), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11661) );
  AOI22_X1 U14726 ( .A1(n11754), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14903), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11660) );
  AOI22_X1 U14727 ( .A1(n14756), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9606), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11659) );
  AOI22_X1 U14728 ( .A1(n11753), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11658) );
  AOI22_X1 U14729 ( .A1(n11754), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14903), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11665) );
  AOI22_X1 U14730 ( .A1(n14756), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11664) );
  AOI22_X1 U14731 ( .A1(n11753), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11663) );
  AOI22_X1 U14732 ( .A1(n11756), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11666) );
  NAND2_X2 U14733 ( .A1(n11669), .A2(n11668), .ZN(n11773) );
  NOR2_X1 U14734 ( .A1(n11791), .A2(n11773), .ZN(n11706) );
  AOI22_X1 U14735 ( .A1(n11754), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14756), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11674) );
  AOI22_X1 U14736 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11673) );
  AOI22_X1 U14737 ( .A1(n11756), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11672) );
  AOI22_X1 U14738 ( .A1(n14903), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11671) );
  NAND4_X1 U14739 ( .A1(n11674), .A2(n11673), .A3(n11672), .A4(n11671), .ZN(
        n11675) );
  NAND2_X1 U14740 ( .A1(n11675), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11682) );
  AOI22_X1 U14741 ( .A1(n11756), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U14742 ( .A1(n11754), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14756), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U14743 ( .A1(n14903), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11677) );
  AOI22_X1 U14744 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11676) );
  NAND4_X1 U14745 ( .A1(n11679), .A2(n11678), .A3(n11677), .A4(n11676), .ZN(
        n11680) );
  NAND2_X1 U14746 ( .A1(n11680), .A2(n11637), .ZN(n11681) );
  AOI22_X1 U14747 ( .A1(n9603), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14903), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U14748 ( .A1(n11753), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11686) );
  AOI22_X1 U14749 ( .A1(n11754), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11685) );
  AOI22_X1 U14750 ( .A1(n11756), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14756), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11684) );
  NAND4_X1 U14751 ( .A1(n11687), .A2(n11686), .A3(n11685), .A4(n11684), .ZN(
        n11693) );
  AOI22_X1 U14752 ( .A1(n14903), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11689) );
  AOI22_X1 U14753 ( .A1(n11756), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11688) );
  AOI22_X1 U14754 ( .A1(n11754), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14756), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11691) );
  AOI22_X1 U14755 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11690) );
  NAND3_X1 U14756 ( .A1(n10099), .A2(n11691), .A3(n11690), .ZN(n11692) );
  AOI22_X1 U14757 ( .A1(n11754), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14756), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U14758 ( .A1(n11756), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9601), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11697) );
  AOI22_X1 U14759 ( .A1(n14903), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U14760 ( .A1(n11753), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11694) );
  AND3_X1 U14761 ( .A1(n11695), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n11694), .ZN(n11696) );
  NAND3_X1 U14762 ( .A1(n11698), .A2(n11697), .A3(n11696), .ZN(n11705) );
  AOI22_X1 U14763 ( .A1(n11754), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14903), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11703) );
  AOI22_X1 U14764 ( .A1(n14756), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11700) );
  AOI22_X1 U14765 ( .A1(n11756), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11699) );
  AND3_X1 U14766 ( .A1(n11700), .A2(n11637), .A3(n11699), .ZN(n11702) );
  AOI22_X1 U14767 ( .A1(n11753), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11701) );
  NAND3_X1 U14768 ( .A1(n11703), .A2(n11702), .A3(n11701), .ZN(n11704) );
  INV_X1 U14769 ( .A(n11789), .ZN(n11719) );
  AOI22_X1 U14770 ( .A1(n14903), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9606), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11708) );
  AOI22_X1 U14771 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11707) );
  AOI22_X1 U14772 ( .A1(n11756), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11710) );
  AOI22_X1 U14773 ( .A1(n11754), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14756), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11709) );
  NAND3_X1 U14774 ( .A1(n11711), .A2(n11710), .A3(n11709), .ZN(n11718) );
  AOI22_X1 U14775 ( .A1(n11754), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14903), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U14776 ( .A1(n11756), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9603), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11714) );
  AOI22_X1 U14777 ( .A1(n11753), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11712) );
  NAND2_X1 U14778 ( .A1(n11716), .A2(n11637), .ZN(n11717) );
  NAND2_X1 U14779 ( .A1(n11719), .A2(n19860), .ZN(n11746) );
  NAND3_X1 U14780 ( .A1(n11720), .A2(n13316), .A3(n11794), .ZN(n11721) );
  NOR2_X2 U14781 ( .A1(n11721), .A2(n12690), .ZN(n12549) );
  NAND2_X1 U14782 ( .A1(n12549), .A2(n13344), .ZN(n12434) );
  NAND2_X1 U14783 ( .A1(n11746), .A2(n12434), .ZN(n11807) );
  MUX2_X1 U14784 ( .A(n19828), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n11730) );
  NAND2_X1 U14785 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19839), .ZN(
        n12505) );
  INV_X1 U14786 ( .A(n12505), .ZN(n11722) );
  NAND2_X1 U14787 ( .A1(n11730), .A2(n11722), .ZN(n11731) );
  NAND2_X1 U14788 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n19828), .ZN(
        n11723) );
  XNOR2_X1 U14789 ( .A(n11637), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11732) );
  NAND2_X1 U14790 ( .A1(n19811), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11725) );
  NAND2_X1 U14791 ( .A1(n16292), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11727) );
  NAND2_X1 U14792 ( .A1(n11735), .A2(n11727), .ZN(n11729) );
  INV_X1 U14793 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16286) );
  NAND2_X1 U14794 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16286), .ZN(
        n11728) );
  INV_X1 U14795 ( .A(n11730), .ZN(n12506) );
  NAND2_X1 U14796 ( .A1(n12506), .A2(n12505), .ZN(n12554) );
  AND2_X1 U14797 ( .A1(n12554), .A2(n11731), .ZN(n12507) );
  XNOR2_X1 U14798 ( .A(n11733), .B(n11732), .ZN(n12300) );
  INV_X1 U14799 ( .A(n12300), .ZN(n11736) );
  NOR2_X1 U14800 ( .A1(n16292), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11734) );
  NAND2_X1 U14801 ( .A1(n11735), .A2(n11734), .ZN(n12304) );
  XNOR2_X1 U14802 ( .A(n11737), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11738) );
  XNOR2_X1 U14803 ( .A(n11739), .B(n11738), .ZN(n12504) );
  NAND2_X1 U14804 ( .A1(n12555), .A2(n12504), .ZN(n12562) );
  INV_X1 U14805 ( .A(n12562), .ZN(n11740) );
  NAND2_X1 U14806 ( .A1(n12507), .A2(n11740), .ZN(n11741) );
  NAND2_X1 U14807 ( .A1(n12437), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11742) );
  OR2_X1 U14808 ( .A1(n11742), .A2(n19852), .ZN(n19049) );
  NAND2_X1 U14809 ( .A1(n11807), .A2(n12435), .ZN(n19855) );
  NAND2_X1 U14810 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19852), .ZN(n13431) );
  NOR2_X1 U14811 ( .A1(n11742), .A2(n13431), .ZN(n16293) );
  NOR2_X1 U14812 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19853) );
  NOR2_X2 U14813 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19812) );
  NAND2_X1 U14814 ( .A1(n18921), .A2(n19713), .ZN(n11743) );
  NOR2_X1 U14815 ( .A1(n16293), .A2(n11743), .ZN(n11744) );
  NOR2_X2 U14816 ( .A1(n18963), .A2(n19416), .ZN(n18957) );
  AOI22_X1 U14817 ( .A1(n11745), .A2(n18951), .B1(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18957), .ZN(n12324) );
  INV_X1 U14818 ( .A(n11746), .ZN(n12317) );
  AOI22_X1 U14819 ( .A1(n11756), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9603), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11750) );
  AOI22_X1 U14820 ( .A1(n14756), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9606), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11749) );
  AOI22_X1 U14821 ( .A1(n11753), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11748) );
  AOI22_X1 U14822 ( .A1(n11754), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14903), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11747) );
  NAND4_X1 U14823 ( .A1(n11750), .A2(n11749), .A3(n11748), .A4(n11747), .ZN(
        n11751) );
  NAND2_X1 U14824 ( .A1(n11751), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11763) );
  AOI22_X1 U14825 ( .A1(n14756), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11760) );
  AOI22_X1 U14826 ( .A1(n11753), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11759) );
  AOI22_X1 U14827 ( .A1(n11754), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14903), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11758) );
  AOI22_X1 U14828 ( .A1(n11756), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9603), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11757) );
  NAND4_X1 U14829 ( .A1(n11760), .A2(n11759), .A3(n11758), .A4(n11757), .ZN(
        n11761) );
  NAND2_X1 U14830 ( .A1(n12317), .A2(n11798), .ZN(n12297) );
  NAND2_X1 U14831 ( .A1(n11766), .A2(n11798), .ZN(n12510) );
  INV_X1 U14832 ( .A(n12510), .ZN(n12548) );
  NOR2_X1 U14833 ( .A1(n12690), .A2(n13826), .ZN(n11764) );
  NAND2_X1 U14834 ( .A1(n12685), .A2(n11764), .ZN(n11808) );
  INV_X2 U14835 ( .A(n11766), .ZN(n19860) );
  NOR2_X1 U14836 ( .A1(n11791), .A2(n19860), .ZN(n11767) );
  OR2_X1 U14837 ( .A1(n11767), .A2(n11768), .ZN(n11770) );
  NAND2_X1 U14838 ( .A1(n11793), .A2(n11768), .ZN(n11769) );
  AND4_X2 U14839 ( .A1(n12440), .A2(n10110), .A3(n11770), .A4(n11769), .ZN(
        n12536) );
  NAND3_X1 U14840 ( .A1(n12297), .A2(n11771), .A3(n15591), .ZN(n11772) );
  AND2_X2 U14841 ( .A1(n11772), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11826) );
  AND2_X1 U14842 ( .A1(n13002), .A2(n11773), .ZN(n11774) );
  NAND2_X1 U14843 ( .A1(n11775), .A2(n11774), .ZN(n13340) );
  INV_X1 U14844 ( .A(n13340), .ZN(n12684) );
  INV_X1 U14845 ( .A(n11931), .ZN(n11776) );
  INV_X1 U14846 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n12306) );
  INV_X1 U14847 ( .A(n11789), .ZN(n13315) );
  INV_X4 U14848 ( .A(n11904), .ZN(n14017) );
  NAND2_X1 U14849 ( .A1(n14017), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11780) );
  NAND2_X1 U14850 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11779) );
  OAI211_X1 U14851 ( .C1(n14020), .C2(n12306), .A(n11780), .B(n11779), .ZN(
        n11781) );
  AOI21_X1 U14852 ( .B1(n11927), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n11781), .ZN(n13035) );
  NAND2_X1 U14853 ( .A1(n11826), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11786) );
  INV_X1 U14854 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n11783) );
  OAI21_X1 U14855 ( .B1(n9605), .B2(n11783), .A(n11782), .ZN(n11784) );
  INV_X1 U14856 ( .A(n11784), .ZN(n11785) );
  NAND2_X1 U14857 ( .A1(n11786), .A2(n11785), .ZN(n11812) );
  NAND2_X1 U14858 ( .A1(n12558), .A2(n10116), .ZN(n11790) );
  NAND2_X1 U14859 ( .A1(n11790), .A2(n11789), .ZN(n12537) );
  OAI21_X1 U14860 ( .B1(n11792), .B2(n11800), .A(n11791), .ZN(n12528) );
  INV_X1 U14861 ( .A(n11797), .ZN(n11793) );
  NAND2_X1 U14862 ( .A1(n11793), .A2(n15640), .ZN(n12525) );
  NAND3_X1 U14863 ( .A1(n12524), .A2(n12525), .A3(n12772), .ZN(n13336) );
  NAND2_X1 U14864 ( .A1(n13336), .A2(n11768), .ZN(n11796) );
  NAND2_X1 U14865 ( .A1(n11796), .A2(n11795), .ZN(n11799) );
  NAND2_X1 U14866 ( .A1(n11793), .A2(n11798), .ZN(n13339) );
  NAND2_X1 U14867 ( .A1(n11799), .A2(n13339), .ZN(n11805) );
  OAI211_X1 U14868 ( .C1(n12700), .C2(n11794), .A(n13436), .B(n12772), .ZN(
        n11804) );
  MUX2_X1 U14869 ( .A(n11801), .B(n13345), .S(n11800), .Z(n11803) );
  INV_X1 U14870 ( .A(n12549), .ZN(n11802) );
  OAI211_X1 U14871 ( .C1(n11804), .C2(n11803), .A(n11802), .B(n13344), .ZN(
        n13349) );
  OAI211_X1 U14872 ( .C1(n12537), .C2(n13344), .A(n11805), .B(n13349), .ZN(
        n11806) );
  NAND2_X2 U14873 ( .A1(n11806), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11825) );
  INV_X1 U14874 ( .A(n11807), .ZN(n16270) );
  NAND2_X1 U14875 ( .A1(n16270), .A2(n11808), .ZN(n13333) );
  OR2_X2 U14876 ( .A1(n11812), .A2(n11811), .ZN(n11823) );
  NAND2_X1 U14877 ( .A1(n11811), .A2(n11812), .ZN(n11813) );
  NAND2_X1 U14878 ( .A1(n11826), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11819) );
  INV_X1 U14879 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13199) );
  NAND2_X1 U14880 ( .A1(n11827), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11816) );
  AND2_X1 U14881 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11814) );
  NOR2_X1 U14882 ( .A1(n19853), .A2(n11814), .ZN(n11815) );
  OAI211_X1 U14883 ( .C1(n9605), .C2(n13199), .A(n11816), .B(n11815), .ZN(
        n11817) );
  INV_X1 U14884 ( .A(n11817), .ZN(n11818) );
  NAND3_X1 U14885 ( .A1(n11825), .A2(n11819), .A3(n11818), .ZN(n12607) );
  NAND2_X1 U14886 ( .A1(n19853), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11820) );
  OAI211_X1 U14887 ( .C1(n11825), .C2(n15573), .A(n11822), .B(n11851), .ZN(
        n12606) );
  AOI21_X1 U14888 ( .B1(n11587), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n11824) );
  OAI21_X1 U14889 ( .B1(n11825), .B2(n11737), .A(n11824), .ZN(n11834) );
  INV_X1 U14890 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n11829) );
  AOI22_X1 U14891 ( .A1(n11827), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11828) );
  OAI21_X1 U14892 ( .B1(n11851), .B2(n11829), .A(n11828), .ZN(n11830) );
  INV_X1 U14893 ( .A(n11830), .ZN(n11831) );
  NAND2_X1 U14894 ( .A1(n11832), .A2(n11831), .ZN(n11833) );
  OR2_X2 U14895 ( .A1(n11834), .A2(n11833), .ZN(n11836) );
  NAND2_X1 U14896 ( .A1(n11834), .A2(n11833), .ZN(n11835) );
  NAND2_X1 U14897 ( .A1(n19853), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11837) );
  OAI21_X1 U14898 ( .B1(n11825), .B2(n11637), .A(n11837), .ZN(n11843) );
  AOI22_X1 U14899 ( .A1(n14017), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11840) );
  INV_X1 U14900 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n12838) );
  NAND2_X1 U14901 ( .A1(n11843), .A2(n11842), .ZN(n11844) );
  INV_X1 U14902 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n11848) );
  NAND2_X1 U14903 ( .A1(n11927), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11847) );
  AOI22_X1 U14904 ( .A1(n14017), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11846) );
  OAI211_X1 U14905 ( .C1(n14020), .C2(n11848), .A(n11847), .B(n11846), .ZN(
        n13008) );
  INV_X1 U14906 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n12929) );
  NAND2_X1 U14907 ( .A1(n11927), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11850) );
  AOI22_X1 U14908 ( .A1(n14017), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11849) );
  OAI211_X1 U14909 ( .C1(n14020), .C2(n12929), .A(n11850), .B(n11849), .ZN(
        n12925) );
  INV_X1 U14910 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12308) );
  AOI22_X1 U14911 ( .A1(n14017), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11852) );
  OAI21_X1 U14912 ( .B1(n14020), .B2(n12308), .A(n11852), .ZN(n11853) );
  AOI21_X1 U14913 ( .B1(n11927), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n11853), .ZN(n13110) );
  INV_X1 U14914 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n13151) );
  NAND2_X1 U14915 ( .A1(n11914), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11855) );
  AOI22_X1 U14916 ( .A1(n14017), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11854) );
  OAI211_X1 U14917 ( .C1(n13151), .C2(n14020), .A(n11855), .B(n11854), .ZN(
        n13048) );
  NAND2_X1 U14918 ( .A1(n14017), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11857) );
  NAND2_X1 U14919 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11856) );
  OAI211_X1 U14920 ( .C1(n14020), .C2(n9880), .A(n11857), .B(n11856), .ZN(
        n11858) );
  AOI21_X1 U14921 ( .B1(n11927), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n11858), .ZN(n13064) );
  NAND2_X1 U14922 ( .A1(n11914), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11863) );
  INV_X1 U14923 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n18918) );
  NAND2_X1 U14924 ( .A1(n14017), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11860) );
  NAND2_X1 U14925 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11859) );
  OAI211_X1 U14926 ( .C1(n14020), .C2(n18918), .A(n11860), .B(n11859), .ZN(
        n11861) );
  INV_X1 U14927 ( .A(n11861), .ZN(n11862) );
  NAND2_X1 U14928 ( .A1(n11863), .A2(n11862), .ZN(n13070) );
  INV_X1 U14929 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n11866) );
  NAND2_X1 U14930 ( .A1(n14017), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11865) );
  NAND2_X1 U14931 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11864) );
  OAI211_X1 U14932 ( .C1(n14020), .C2(n11866), .A(n11865), .B(n11864), .ZN(
        n11867) );
  AOI21_X1 U14933 ( .B1(n11927), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n11867), .ZN(n13172) );
  INV_X1 U14934 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n18889) );
  NAND2_X1 U14935 ( .A1(n14017), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11869) );
  NAND2_X1 U14936 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11868) );
  OAI211_X1 U14937 ( .C1(n14020), .C2(n18889), .A(n11869), .B(n11868), .ZN(
        n11870) );
  AOI21_X1 U14938 ( .B1(n11927), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n11870), .ZN(n13183) );
  INV_X1 U14939 ( .A(n11914), .ZN(n11922) );
  INV_X1 U14940 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n20796) );
  AOI22_X1 U14941 ( .A1(n14017), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11872) );
  NAND2_X1 U14942 ( .A1(n11838), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11871) );
  OAI211_X1 U14943 ( .C1(n11922), .C2(n20796), .A(n11872), .B(n11871), .ZN(
        n13219) );
  INV_X1 U14944 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n11875) );
  NAND2_X1 U14945 ( .A1(n14017), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11874) );
  NAND2_X1 U14946 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11873) );
  OAI211_X1 U14947 ( .C1(n14020), .C2(n11875), .A(n11874), .B(n11873), .ZN(
        n11876) );
  AOI21_X1 U14948 ( .B1(n11927), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n11876), .ZN(n13403) );
  INV_X1 U14949 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n11879) );
  NAND2_X1 U14950 ( .A1(n14017), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11878) );
  NAND2_X1 U14951 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11877) );
  OAI211_X1 U14952 ( .C1(n14020), .C2(n11879), .A(n11878), .B(n11877), .ZN(
        n11880) );
  AOI21_X1 U14953 ( .B1(n11914), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n11880), .ZN(n13526) );
  INV_X1 U14954 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15786) );
  AOI22_X1 U14955 ( .A1(n14017), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n11882) );
  NAND2_X1 U14956 ( .A1(n11838), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11881) );
  OAI211_X1 U14957 ( .C1(n11922), .C2(n15786), .A(n11882), .B(n11881), .ZN(
        n13627) );
  INV_X1 U14958 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n11885) );
  NAND2_X1 U14959 ( .A1(n14017), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11884) );
  NAND2_X1 U14960 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11883) );
  OAI211_X1 U14961 ( .C1(n14020), .C2(n11885), .A(n11884), .B(n11883), .ZN(
        n11886) );
  AOI21_X1 U14962 ( .B1(n11927), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11886), .ZN(n13649) );
  INV_X1 U14963 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n18820) );
  NAND2_X1 U14964 ( .A1(n14017), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11888) );
  NAND2_X1 U14965 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11887) );
  OAI211_X1 U14966 ( .C1(n14020), .C2(n18820), .A(n11888), .B(n11887), .ZN(
        n11889) );
  AOI21_X1 U14967 ( .B1(n11914), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n11889), .ZN(n13710) );
  INV_X1 U14968 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n11892) );
  NAND2_X1 U14969 ( .A1(n14017), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11891) );
  NAND2_X1 U14970 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11890) );
  OAI211_X1 U14971 ( .C1(n14020), .C2(n11892), .A(n11891), .B(n11890), .ZN(
        n11893) );
  AOI21_X1 U14972 ( .B1(n11927), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n11893), .ZN(n15057) );
  INV_X1 U14973 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15419) );
  AOI22_X1 U14974 ( .A1(n14017), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n11895) );
  NAND2_X1 U14975 ( .A1(n11838), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11894) );
  OAI211_X1 U14976 ( .C1(n11922), .C2(n15419), .A(n11895), .B(n11894), .ZN(
        n15040) );
  INV_X1 U14977 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n11898) );
  NAND2_X1 U14978 ( .A1(n14017), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11897) );
  NAND2_X1 U14979 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11896) );
  OAI211_X1 U14980 ( .C1(n14020), .C2(n11898), .A(n11897), .B(n11896), .ZN(
        n11899) );
  AOI21_X1 U14981 ( .B1(n11927), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n11899), .ZN(n12391) );
  INV_X1 U14982 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n15796) );
  NAND2_X1 U14983 ( .A1(n14017), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11901) );
  NAND2_X1 U14984 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11900) );
  OAI211_X1 U14985 ( .C1(n14020), .C2(n15796), .A(n11901), .B(n11900), .ZN(
        n11902) );
  AOI21_X1 U14986 ( .B1(n11927), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n11902), .ZN(n15028) );
  NAND2_X1 U14987 ( .A1(n11914), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11908) );
  INV_X1 U14988 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n11903) );
  NOR2_X1 U14989 ( .A1(n14020), .A2(n11903), .ZN(n11906) );
  INV_X1 U14990 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20860) );
  OAI22_X1 U14991 ( .A1(n11904), .A2(n20860), .B1(n12437), .B2(n20877), .ZN(
        n11905) );
  NOR2_X1 U14992 ( .A1(n11906), .A2(n11905), .ZN(n11907) );
  NAND2_X1 U14993 ( .A1(n11908), .A2(n11907), .ZN(n12404) );
  AOI22_X1 U14994 ( .A1(n14017), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n11910) );
  NAND2_X1 U14995 ( .A1(n11838), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11909) );
  OAI211_X1 U14996 ( .C1(n11922), .C2(n10017), .A(n11910), .B(n11909), .ZN(
        n15019) );
  INV_X1 U14997 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n15010) );
  NAND2_X1 U14998 ( .A1(n14017), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11912) );
  NAND2_X1 U14999 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11911) );
  OAI211_X1 U15000 ( .C1(n14020), .C2(n15010), .A(n11912), .B(n11911), .ZN(
        n11913) );
  AOI21_X1 U15001 ( .B1(n11914), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n11913), .ZN(n14729) );
  INV_X1 U15002 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n14717) );
  NAND2_X1 U15003 ( .A1(n14017), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11916) );
  NAND2_X1 U15004 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11915) );
  OAI211_X1 U15005 ( .C1(n14020), .C2(n14717), .A(n11916), .B(n11915), .ZN(
        n11917) );
  AOI21_X1 U15006 ( .B1(n11927), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11917), .ZN(n14707) );
  INV_X1 U15007 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15323) );
  AOI22_X1 U15008 ( .A1(n14017), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11919) );
  NAND2_X1 U15009 ( .A1(n11838), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11918) );
  OAI211_X1 U15010 ( .C1(n11922), .C2(n15323), .A(n11919), .B(n11918), .ZN(
        n14691) );
  AND2_X2 U15011 ( .A1(n14708), .A2(n14691), .ZN(n14693) );
  INV_X1 U15012 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15313) );
  AOI22_X1 U15013 ( .A1(n14017), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11921) );
  NAND2_X1 U15014 ( .A1(n11838), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11920) );
  OAI211_X1 U15015 ( .C1(n11922), .C2(n15313), .A(n11921), .B(n11920), .ZN(
        n12379) );
  INV_X1 U15016 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n11925) );
  NAND2_X1 U15017 ( .A1(n14017), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11924) );
  NAND2_X1 U15018 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11923) );
  OAI211_X1 U15019 ( .C1(n14020), .C2(n11925), .A(n11924), .B(n11923), .ZN(
        n11926) );
  AOI21_X1 U15020 ( .B1(n11927), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n11926), .ZN(n14672) );
  INV_X1 U15021 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n11930) );
  NAND2_X1 U15022 ( .A1(n11927), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11929) );
  AOI22_X1 U15023 ( .A1(n14017), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11928) );
  OAI211_X1 U15024 ( .C1(n14020), .C2(n11930), .A(n11929), .B(n11928), .ZN(
        n14021) );
  NAND2_X1 U15025 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19859) );
  INV_X1 U15026 ( .A(n19859), .ZN(n19717) );
  NOR2_X1 U15027 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19717), .ZN(n12318) );
  NAND2_X1 U15028 ( .A1(n11776), .A2(n12318), .ZN(n11932) );
  NOR2_X1 U15029 ( .A1(n11773), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12020) );
  NAND2_X1 U15030 ( .A1(n11995), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11935) );
  AND2_X1 U15031 ( .A1(n11773), .A2(n19416), .ZN(n12000) );
  AOI22_X1 U15032 ( .A1(n12137), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n12279), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11934) );
  AND2_X1 U15033 ( .A1(n11935), .A2(n11934), .ZN(n12296) );
  INV_X2 U15034 ( .A(n12089), .ZN(n12144) );
  AOI22_X1 U15035 ( .A1(n12053), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12144), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11945) );
  INV_X2 U15036 ( .A(n14941), .ZN(n14972) );
  AND2_X2 U15037 ( .A1(n14972), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12004) );
  INV_X1 U15038 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11940) );
  AND2_X1 U15039 ( .A1(n11936), .A2(n14758), .ZN(n11964) );
  NAND2_X1 U15040 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11939) );
  NAND2_X1 U15041 ( .A1(n11963), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11938) );
  OAI211_X1 U15042 ( .C1(n12111), .C2(n11940), .A(n11939), .B(n11938), .ZN(
        n11941) );
  INV_X1 U15043 ( .A(n11941), .ZN(n11944) );
  AOI22_X1 U15044 ( .A1(n14861), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14862), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11943) );
  AOI22_X1 U15045 ( .A1(n12056), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12057), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11942) );
  NAND4_X1 U15046 ( .A1(n11945), .A2(n11944), .A3(n11943), .A4(n11942), .ZN(
        n11954) );
  AND2_X1 U15047 ( .A1(n14903), .A2(n11637), .ZN(n11980) );
  AOI22_X1 U15048 ( .A1(n14867), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11952) );
  AND2_X1 U15049 ( .A1(n11936), .A2(n14757), .ZN(n12026) );
  AND2_X1 U15050 ( .A1(n14758), .A2(n11947), .ZN(n12027) );
  AOI22_X1 U15051 ( .A1(n12026), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12027), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11951) );
  AND2_X1 U15052 ( .A1(n11937), .A2(n14758), .ZN(n12003) );
  AND2_X1 U15053 ( .A1(n11948), .A2(n14758), .ZN(n11958) );
  AOI22_X1 U15054 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11950) );
  NAND2_X1 U15055 ( .A1(n14868), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11949) );
  NAND4_X1 U15056 ( .A1(n11952), .A2(n11951), .A3(n11950), .A4(n11949), .ZN(
        n11953) );
  INV_X1 U15057 ( .A(n12307), .ZN(n13563) );
  NAND2_X1 U15058 ( .A1(n11995), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11957) );
  INV_X1 U15059 ( .A(n12000), .ZN(n12044) );
  AOI22_X1 U15060 ( .A1(n12137), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n12279), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11956) );
  OAI211_X1 U15061 ( .C1(n13563), .C2(n12270), .A(n11957), .B(n11956), .ZN(
        n13594) );
  AOI22_X1 U15062 ( .A1(n12053), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U15063 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n12026), .B1(
        n12027), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11961) );
  AOI22_X1 U15064 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12003), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11960) );
  NAND2_X1 U15065 ( .A1(n14868), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11959) );
  NAND4_X1 U15066 ( .A1(n11962), .A2(n11961), .A3(n11960), .A4(n11959), .ZN(
        n11974) );
  AOI22_X1 U15067 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12057), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11972) );
  INV_X1 U15068 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11967) );
  NAND2_X1 U15069 ( .A1(n11963), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11966) );
  NAND2_X1 U15070 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11965) );
  OAI211_X1 U15071 ( .C1(n12097), .C2(n11967), .A(n11966), .B(n11965), .ZN(
        n11968) );
  INV_X1 U15072 ( .A(n11968), .ZN(n11971) );
  AOI22_X1 U15073 ( .A1(n12056), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14867), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11970) );
  AOI22_X1 U15074 ( .A1(n14862), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11969) );
  NAND4_X1 U15075 ( .A1(n11972), .A2(n11971), .A3(n11970), .A4(n11969), .ZN(
        n11973) );
  INV_X1 U15076 ( .A(n13491), .ZN(n13542) );
  NAND2_X1 U15077 ( .A1(n12000), .A2(P2_EAX_REG_4__SCAN_IN), .ZN(n11976) );
  NAND2_X1 U15078 ( .A1(n12282), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11975) );
  OAI211_X1 U15079 ( .C1(n12270), .C2(n13542), .A(n11976), .B(n11975), .ZN(
        n11977) );
  INV_X1 U15080 ( .A(n11977), .ZN(n11979) );
  NAND2_X1 U15081 ( .A1(n11995), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11978) );
  AOI22_X1 U15082 ( .A1(n14867), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12057), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11984) );
  AOI22_X1 U15083 ( .A1(n12053), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12056), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11983) );
  AOI22_X1 U15084 ( .A1(n14868), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14861), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11982) );
  AOI22_X1 U15085 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11981) );
  NAND4_X1 U15086 ( .A1(n11984), .A2(n11983), .A3(n11982), .A4(n11981), .ZN(
        n11990) );
  AOI22_X1 U15087 ( .A1(n12026), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12003), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11988) );
  AOI22_X1 U15088 ( .A1(n12027), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11987) );
  AOI22_X1 U15089 ( .A1(n11963), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11964), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11986) );
  AOI22_X1 U15090 ( .A1(n14862), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11985) );
  NAND4_X1 U15091 ( .A1(n11988), .A2(n11987), .A3(n11986), .A4(n11985), .ZN(
        n11989) );
  AND2_X1 U15092 ( .A1(n19839), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11992) );
  NAND2_X1 U15093 ( .A1(n12700), .A2(n12279), .ZN(n12042) );
  OAI21_X1 U15094 ( .B1(n12020), .B2(n11992), .A(n12042), .ZN(n11993) );
  INV_X1 U15095 ( .A(n11993), .ZN(n11994) );
  INV_X1 U15096 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18788) );
  NAND2_X1 U15097 ( .A1(n11995), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11999) );
  NAND2_X1 U15098 ( .A1(n11773), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n11997) );
  AOI21_X1 U15099 ( .B1(n14935), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11996) );
  AND2_X1 U15100 ( .A1(n11997), .A2(n11996), .ZN(n11998) );
  NAND2_X1 U15101 ( .A1(n11999), .A2(n11998), .ZN(n12696) );
  INV_X1 U15102 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19734) );
  NAND2_X1 U15103 ( .A1(n11995), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n12002) );
  INV_X1 U15104 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19150) );
  AOI22_X1 U15105 ( .A1(n12000), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12282), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12001) );
  NAND2_X1 U15106 ( .A1(n12002), .A2(n12001), .ZN(n12023) );
  XNOR2_X1 U15107 ( .A(n12699), .B(n12023), .ZN(n13040) );
  AOI22_X1 U15108 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12003), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12009) );
  NAND2_X1 U15109 ( .A1(n12056), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12008) );
  NAND2_X1 U15110 ( .A1(n12004), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12007) );
  INV_X1 U15111 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12005) );
  OR2_X1 U15112 ( .A1(n12255), .A2(n12005), .ZN(n12006) );
  NAND4_X1 U15113 ( .A1(n12009), .A2(n12008), .A3(n12007), .A4(n12006), .ZN(
        n12013) );
  NAND2_X1 U15114 ( .A1(n12053), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12011) );
  NAND2_X1 U15115 ( .A1(n11980), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12010) );
  NOR4_X1 U15116 ( .A1(n12013), .A2(n10111), .A3(n10105), .A4(n12012), .ZN(
        n12019) );
  AOI22_X1 U15117 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n14867), .B1(
        n12057), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U15118 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n11963), .B1(
        n12027), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12016) );
  AOI22_X1 U15119 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n11964), .B1(
        n12026), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12015) );
  NAND2_X1 U15120 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12014) );
  AND4_X1 U15121 ( .A1(n12017), .A2(n12016), .A3(n12015), .A4(n12014), .ZN(
        n12018) );
  NAND2_X1 U15122 ( .A1(n11793), .A2(n12020), .ZN(n12022) );
  NAND2_X1 U15123 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12021) );
  OAI211_X1 U15124 ( .C1(n12270), .C2(n12575), .A(n12022), .B(n12021), .ZN(
        n13039) );
  NOR2_X1 U15125 ( .A1(n13040), .A2(n13039), .ZN(n12025) );
  NOR2_X1 U15126 ( .A1(n12699), .A2(n12023), .ZN(n12024) );
  AOI22_X1 U15127 ( .A1(n12053), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14867), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12031) );
  AOI22_X1 U15128 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n12026), .B1(
        n12027), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12030) );
  AOI22_X1 U15129 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n12003), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12029) );
  NAND2_X1 U15130 ( .A1(n14868), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n12028) );
  NAND4_X1 U15131 ( .A1(n12031), .A2(n12030), .A3(n12029), .A4(n12028), .ZN(
        n12041) );
  AOI22_X1 U15132 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12057), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12039) );
  INV_X1 U15133 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12034) );
  NAND2_X1 U15134 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n12033) );
  NAND2_X1 U15135 ( .A1(n11963), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n12032) );
  OAI211_X1 U15136 ( .C1(n12255), .C2(n12034), .A(n12033), .B(n12032), .ZN(
        n12035) );
  INV_X1 U15137 ( .A(n12035), .ZN(n12038) );
  AOI22_X1 U15138 ( .A1(n12056), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12037) );
  AOI22_X1 U15139 ( .A1(n14861), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12036) );
  NAND4_X1 U15140 ( .A1(n12039), .A2(n12038), .A3(n12037), .A4(n12036), .ZN(
        n12040) );
  NAND2_X1 U15141 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12043) );
  OAI211_X1 U15142 ( .C1(n12270), .C2(n13302), .A(n12043), .B(n12042), .ZN(
        n12047) );
  XNOR2_X1 U15143 ( .A(n12048), .B(n12047), .ZN(n12910) );
  INV_X1 U15144 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19736) );
  NAND2_X1 U15145 ( .A1(n11995), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12046) );
  BUF_X1 U15146 ( .A(n12279), .Z(n12282) );
  AOI22_X1 U15147 ( .A1(n12000), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n12282), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12045) );
  NAND2_X1 U15148 ( .A1(n12046), .A2(n12045), .ZN(n12909) );
  NOR2_X1 U15149 ( .A1(n12048), .A2(n12047), .ZN(n12049) );
  NAND2_X1 U15150 ( .A1(n11995), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U15151 ( .A1(n12282), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12077) );
  INV_X1 U15152 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12051) );
  INV_X1 U15153 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12050) );
  OAI22_X1 U15154 ( .A1(n12051), .A2(n12083), .B1(n12084), .B2(n12050), .ZN(
        n12052) );
  INV_X1 U15155 ( .A(n12052), .ZN(n12067) );
  INV_X1 U15156 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12055) );
  INV_X1 U15157 ( .A(n12053), .ZN(n12088) );
  INV_X1 U15158 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12054) );
  OAI22_X1 U15159 ( .A1(n12055), .A2(n12088), .B1(n12089), .B2(n12054), .ZN(
        n12060) );
  INV_X1 U15160 ( .A(n12056), .ZN(n12093) );
  INV_X1 U15161 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12058) );
  INV_X1 U15162 ( .A(n12057), .ZN(n12091) );
  INV_X1 U15163 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19176) );
  OAI22_X1 U15164 ( .A1(n12093), .A2(n12058), .B1(n12091), .B2(n19176), .ZN(
        n12059) );
  INV_X1 U15165 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12063) );
  NAND2_X1 U15166 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n12062) );
  NAND2_X1 U15167 ( .A1(n11963), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12061) );
  OAI211_X1 U15168 ( .C1(n12111), .C2(n12063), .A(n12062), .B(n12061), .ZN(
        n12064) );
  INV_X1 U15169 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13266) );
  AOI22_X1 U15170 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n12026), .B1(
        n12027), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12069) );
  AOI22_X1 U15171 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12003), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12068) );
  OAI211_X1 U15172 ( .C1(n13266), .C2(n12081), .A(n12069), .B(n12068), .ZN(
        n12073) );
  INV_X1 U15173 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12071) );
  INV_X1 U15174 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12070) );
  OAI22_X1 U15175 ( .A1(n12071), .A2(n12097), .B1(n12255), .B2(n12070), .ZN(
        n12072) );
  OR2_X1 U15176 ( .A1(n12270), .A2(n10101), .ZN(n12076) );
  NAND2_X1 U15177 ( .A1(n12137), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12075) );
  NAND4_X1 U15178 ( .A1(n12078), .A2(n12077), .A3(n12076), .A4(n12075), .ZN(
        n13082) );
  INV_X1 U15179 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U15180 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n12026), .B1(
        n12027), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12080) );
  AOI22_X1 U15181 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n12003), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12079) );
  OAI211_X1 U15182 ( .C1(n12082), .C2(n12081), .A(n12080), .B(n12079), .ZN(
        n12086) );
  INV_X1 U15183 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13666) );
  INV_X1 U15184 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13664) );
  OAI22_X1 U15185 ( .A1(n13666), .A2(n12084), .B1(n12083), .B2(n13664), .ZN(
        n12085) );
  NOR2_X1 U15186 ( .A1(n12086), .A2(n12085), .ZN(n12106) );
  INV_X1 U15187 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12090) );
  INV_X1 U15188 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12087) );
  OAI22_X1 U15189 ( .A1(n12090), .A2(n12089), .B1(n12088), .B2(n12087), .ZN(
        n12095) );
  INV_X1 U15190 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12092) );
  INV_X1 U15191 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19185) );
  OAI22_X1 U15192 ( .A1(n12093), .A2(n12092), .B1(n12091), .B2(n19185), .ZN(
        n12094) );
  NOR2_X1 U15193 ( .A1(n12095), .A2(n12094), .ZN(n12105) );
  INV_X1 U15194 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12098) );
  INV_X1 U15195 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12096) );
  OAI22_X1 U15196 ( .A1(n12098), .A2(n12097), .B1(n12255), .B2(n12096), .ZN(
        n12103) );
  INV_X1 U15197 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12101) );
  NAND2_X1 U15198 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n12100) );
  NAND2_X1 U15199 ( .A1(n11963), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12099) );
  OAI211_X1 U15200 ( .C1(n12111), .C2(n12101), .A(n12100), .B(n12099), .ZN(
        n12102) );
  NOR2_X1 U15201 ( .A1(n12103), .A2(n12102), .ZN(n12104) );
  INV_X1 U15202 ( .A(n13679), .ZN(n12107) );
  AOI222_X1 U15203 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n11995), .B1(n12279), 
        .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(P2_EAX_REG_6__SCAN_IN), 
        .C2(n12137), .ZN(n12928) );
  AOI22_X1 U15204 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n14861), .B1(
        n14862), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12116) );
  AOI22_X1 U15205 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12056), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12115) );
  AOI22_X1 U15206 ( .A1(n14868), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12057), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12114) );
  INV_X1 U15207 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12110) );
  NAND2_X1 U15208 ( .A1(n11963), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12109) );
  NAND2_X1 U15209 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n12108) );
  OAI211_X1 U15210 ( .C1(n12111), .C2(n12110), .A(n12109), .B(n12108), .ZN(
        n12112) );
  INV_X1 U15211 ( .A(n12112), .ZN(n12113) );
  NAND4_X1 U15212 ( .A1(n12116), .A2(n12115), .A3(n12114), .A4(n12113), .ZN(
        n12122) );
  AOI22_X1 U15213 ( .A1(n12053), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12120) );
  AOI22_X1 U15214 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n12026), .B1(
        n12027), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12119) );
  AOI22_X1 U15215 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n12003), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12118) );
  NAND2_X1 U15216 ( .A1(n14867), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12117) );
  NAND4_X1 U15217 ( .A1(n12120), .A2(n12119), .A3(n12118), .A4(n12117), .ZN(
        n12121) );
  NAND2_X1 U15218 ( .A1(n11995), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n12124) );
  AOI22_X1 U15219 ( .A1(n12000), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n12282), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12123) );
  NAND2_X1 U15220 ( .A1(n12124), .A2(n12123), .ZN(n13119) );
  NAND2_X1 U15221 ( .A1(n13118), .A2(n13119), .ZN(n13146) );
  AOI22_X1 U15222 ( .A1(n11963), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11964), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12126) );
  NAND2_X1 U15223 ( .A1(n14861), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12125) );
  AND2_X1 U15224 ( .A1(n12126), .A2(n12125), .ZN(n12130) );
  AOI22_X1 U15225 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12056), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12129) );
  AOI22_X1 U15226 ( .A1(n14862), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12128) );
  AOI22_X1 U15227 ( .A1(n12053), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12057), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12127) );
  NAND4_X1 U15228 ( .A1(n12130), .A2(n12129), .A3(n12128), .A4(n12127), .ZN(
        n12136) );
  AOI22_X1 U15229 ( .A1(n14867), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12134) );
  AOI22_X1 U15230 ( .A1(n12026), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12027), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U15231 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12132) );
  NAND2_X1 U15232 ( .A1(n14868), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12131) );
  NAND4_X1 U15233 ( .A1(n12134), .A2(n12133), .A3(n12132), .A4(n12131), .ZN(
        n12135) );
  OR2_X1 U15234 ( .A1(n12136), .A2(n12135), .ZN(n13054) );
  INV_X1 U15235 ( .A(n13054), .ZN(n12140) );
  INV_X1 U15236 ( .A(n12044), .ZN(n12137) );
  NAND2_X1 U15237 ( .A1(n12137), .A2(P2_EAX_REG_8__SCAN_IN), .ZN(n12139) );
  NAND2_X1 U15238 ( .A1(n12282), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12138) );
  OAI211_X1 U15239 ( .C1(n12270), .C2(n12140), .A(n12139), .B(n12138), .ZN(
        n12141) );
  INV_X1 U15240 ( .A(n12141), .ZN(n12143) );
  NAND2_X1 U15241 ( .A1(n11995), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12142) );
  NAND2_X1 U15242 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12148) );
  NAND2_X1 U15243 ( .A1(n12053), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12147) );
  NAND2_X1 U15244 ( .A1(n12057), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12146) );
  NAND2_X1 U15245 ( .A1(n12056), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12145) );
  NAND4_X1 U15246 ( .A1(n12148), .A2(n12147), .A3(n12146), .A4(n12145), .ZN(
        n12155) );
  AOI22_X1 U15247 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11964), .B1(
        n11963), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12153) );
  NAND2_X1 U15248 ( .A1(n12004), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12152) );
  NAND2_X1 U15249 ( .A1(n14861), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12151) );
  INV_X1 U15250 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12149) );
  OR2_X1 U15251 ( .A1(n12255), .A2(n12149), .ZN(n12150) );
  NAND4_X1 U15252 ( .A1(n12153), .A2(n12152), .A3(n12151), .A4(n12150), .ZN(
        n12154) );
  NOR2_X1 U15253 ( .A1(n12155), .A2(n12154), .ZN(n12161) );
  AOI22_X1 U15254 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n11980), .B1(
        n14867), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12159) );
  AOI22_X1 U15255 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12026), .B1(
        n12027), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12158) );
  AOI22_X1 U15256 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12003), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12157) );
  NAND2_X1 U15257 ( .A1(n14868), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12156) );
  AND4_X1 U15258 ( .A1(n12159), .A2(n12158), .A3(n12157), .A4(n12156), .ZN(
        n12160) );
  AND2_X1 U15259 ( .A1(n12161), .A2(n12160), .ZN(n13059) );
  NAND2_X1 U15260 ( .A1(n11995), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12163) );
  AOI22_X1 U15261 ( .A1(n12137), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12279), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12162) );
  OAI211_X1 U15262 ( .C1(n13059), .C2(n12270), .A(n12163), .B(n12162), .ZN(
        n13995) );
  AOI22_X1 U15263 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n14861), .B1(
        n12056), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12170) );
  AOI22_X1 U15264 ( .A1(n12053), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12057), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12169) );
  AOI22_X1 U15265 ( .A1(n14862), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12168) );
  NAND2_X1 U15266 ( .A1(n12004), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n12166) );
  NAND2_X1 U15267 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n12165) );
  NAND2_X1 U15268 ( .A1(n11963), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12164) );
  AND3_X1 U15269 ( .A1(n12166), .A2(n12165), .A3(n12164), .ZN(n12167) );
  NAND4_X1 U15270 ( .A1(n12170), .A2(n12169), .A3(n12168), .A4(n12167), .ZN(
        n12176) );
  AOI22_X1 U15271 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14867), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12174) );
  AOI22_X1 U15272 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n12026), .B1(
        n12027), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12173) );
  AOI22_X1 U15273 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12003), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12172) );
  NAND2_X1 U15274 ( .A1(n14868), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12171) );
  NAND4_X1 U15275 ( .A1(n12174), .A2(n12173), .A3(n12172), .A4(n12171), .ZN(
        n12175) );
  NOR2_X1 U15276 ( .A1(n12176), .A2(n12175), .ZN(n13073) );
  AOI22_X1 U15277 ( .A1(n12000), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12279), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12177) );
  OAI21_X1 U15278 ( .B1(n13073), .B2(n12270), .A(n12177), .ZN(n12178) );
  AOI21_X1 U15279 ( .B1(P2_REIP_REG_10__SCAN_IN), .B2(n11995), .A(n12178), 
        .ZN(n15531) );
  NAND2_X1 U15280 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12182) );
  NAND2_X1 U15281 ( .A1(n12053), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n12181) );
  NAND2_X1 U15282 ( .A1(n12057), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12180) );
  NAND2_X1 U15283 ( .A1(n12056), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12179) );
  AND4_X1 U15284 ( .A1(n12182), .A2(n12181), .A3(n12180), .A4(n12179), .ZN(
        n12194) );
  AOI22_X1 U15285 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n11964), .B1(
        n11963), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12187) );
  NAND2_X1 U15286 ( .A1(n12004), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n12186) );
  NAND2_X1 U15287 ( .A1(n14861), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12185) );
  INV_X1 U15288 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12183) );
  OR2_X1 U15289 ( .A1(n12255), .A2(n12183), .ZN(n12184) );
  AND4_X1 U15290 ( .A1(n12187), .A2(n12186), .A3(n12185), .A4(n12184), .ZN(
        n12193) );
  NAND2_X1 U15291 ( .A1(n14868), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n12190) );
  AOI22_X1 U15292 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12026), .B1(
        n12027), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U15293 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12003), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12188) );
  AND3_X1 U15294 ( .A1(n12190), .A2(n12189), .A3(n12188), .ZN(n12192) );
  AOI22_X1 U15295 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n11980), .B1(
        n14867), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12191) );
  NAND4_X1 U15296 ( .A1(n12194), .A2(n12193), .A3(n12192), .A4(n12191), .ZN(
        n13190) );
  AOI22_X1 U15297 ( .A1(n11995), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n11991), 
        .B2(n13190), .ZN(n12196) );
  AOI22_X1 U15298 ( .A1(n12000), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12279), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12195) );
  NAND2_X1 U15299 ( .A1(n12196), .A2(n12195), .ZN(n15504) );
  AOI22_X1 U15300 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12144), .B1(
        n12053), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12204) );
  INV_X1 U15301 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12199) );
  NAND2_X1 U15302 ( .A1(n11963), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12198) );
  NAND2_X1 U15303 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n12197) );
  OAI211_X1 U15304 ( .C1(n12255), .C2(n12199), .A(n12198), .B(n12197), .ZN(
        n12200) );
  INV_X1 U15305 ( .A(n12200), .ZN(n12203) );
  AOI22_X1 U15306 ( .A1(n14861), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12202) );
  AOI22_X1 U15307 ( .A1(n12056), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12057), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12201) );
  NAND4_X1 U15308 ( .A1(n12204), .A2(n12203), .A3(n12202), .A4(n12201), .ZN(
        n12210) );
  AOI22_X1 U15309 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n14867), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12208) );
  AOI22_X1 U15310 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12026), .B1(
        n12027), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12207) );
  AOI22_X1 U15311 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12003), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12206) );
  NAND2_X1 U15312 ( .A1(n14868), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12205) );
  NAND4_X1 U15313 ( .A1(n12208), .A2(n12207), .A3(n12206), .A4(n12205), .ZN(
        n12209) );
  OR2_X1 U15314 ( .A1(n12210), .A2(n12209), .ZN(n13189) );
  INV_X1 U15315 ( .A(n13189), .ZN(n12213) );
  NAND2_X1 U15316 ( .A1(n12137), .A2(P2_EAX_REG_12__SCAN_IN), .ZN(n12212) );
  NAND2_X1 U15317 ( .A1(n12279), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12211) );
  OAI211_X1 U15318 ( .C1(n12270), .C2(n12213), .A(n12212), .B(n12211), .ZN(
        n12214) );
  INV_X1 U15319 ( .A(n12214), .ZN(n12216) );
  NAND2_X1 U15320 ( .A1(n11995), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12215) );
  NOR2_X2 U15321 ( .A1(n15494), .A2(n15495), .ZN(n15477) );
  AOI22_X1 U15322 ( .A1(n12053), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12144), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12223) );
  NAND2_X1 U15323 ( .A1(n12004), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n12219) );
  NAND2_X1 U15324 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n12218) );
  NAND2_X1 U15325 ( .A1(n11963), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12217) );
  AND3_X1 U15326 ( .A1(n12219), .A2(n12218), .A3(n12217), .ZN(n12222) );
  AOI22_X1 U15327 ( .A1(n14862), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14861), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12221) );
  AOI22_X1 U15328 ( .A1(n12056), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12057), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12220) );
  NAND4_X1 U15329 ( .A1(n12223), .A2(n12222), .A3(n12221), .A4(n12220), .ZN(
        n12229) );
  AOI22_X1 U15330 ( .A1(n14867), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12227) );
  AOI22_X1 U15331 ( .A1(n12026), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12027), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U15332 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12225) );
  NAND2_X1 U15333 ( .A1(n14868), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12224) );
  NAND4_X1 U15334 ( .A1(n12227), .A2(n12226), .A3(n12225), .A4(n12224), .ZN(
        n12228) );
  INV_X1 U15335 ( .A(n13216), .ZN(n12232) );
  NAND2_X1 U15336 ( .A1(n11995), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n12231) );
  AOI22_X1 U15337 ( .A1(n12137), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12279), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12230) );
  OAI211_X1 U15338 ( .C1(n12232), .C2(n12270), .A(n12231), .B(n12230), .ZN(
        n15478) );
  NAND2_X1 U15339 ( .A1(n15477), .A2(n15478), .ZN(n15476) );
  AOI22_X1 U15340 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n11964), .B1(
        n11963), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12234) );
  NAND2_X1 U15341 ( .A1(n14861), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12233) );
  AND2_X1 U15342 ( .A1(n12234), .A2(n12233), .ZN(n12238) );
  AOI22_X1 U15343 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12056), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12237) );
  AOI22_X1 U15344 ( .A1(n14862), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12236) );
  AOI22_X1 U15345 ( .A1(n12053), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12057), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12235) );
  NAND4_X1 U15346 ( .A1(n12238), .A2(n12237), .A3(n12236), .A4(n12235), .ZN(
        n12244) );
  AOI22_X1 U15347 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n14867), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12242) );
  AOI22_X1 U15348 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12026), .B1(
        n12027), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12241) );
  AOI22_X1 U15349 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12003), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12240) );
  NAND2_X1 U15350 ( .A1(n14868), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12239) );
  NAND4_X1 U15351 ( .A1(n12242), .A2(n12241), .A3(n12240), .A4(n12239), .ZN(
        n12243) );
  NOR2_X1 U15352 ( .A1(n12244), .A2(n12243), .ZN(n13406) );
  NAND2_X1 U15353 ( .A1(n12000), .A2(P2_EAX_REG_14__SCAN_IN), .ZN(n12246) );
  NAND2_X1 U15354 ( .A1(n12279), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12245) );
  OAI211_X1 U15355 ( .C1(n12270), .C2(n13406), .A(n12246), .B(n12245), .ZN(
        n12247) );
  INV_X1 U15356 ( .A(n12247), .ZN(n12249) );
  NAND2_X1 U15357 ( .A1(n11995), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n12248) );
  NOR2_X2 U15358 ( .A1(n15476), .A2(n16238), .ZN(n16237) );
  NAND2_X1 U15359 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12253) );
  NAND2_X1 U15360 ( .A1(n12053), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n12252) );
  NAND2_X1 U15361 ( .A1(n12057), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12251) );
  NAND2_X1 U15362 ( .A1(n12056), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12250) );
  NAND4_X1 U15363 ( .A1(n12253), .A2(n12252), .A3(n12251), .A4(n12250), .ZN(
        n12261) );
  AOI22_X1 U15364 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n11964), .B1(
        n11963), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12259) );
  NAND2_X1 U15365 ( .A1(n12004), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12258) );
  NAND2_X1 U15366 ( .A1(n14861), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12257) );
  INV_X1 U15367 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12254) );
  OR2_X1 U15368 ( .A1(n12255), .A2(n12254), .ZN(n12256) );
  NAND4_X1 U15369 ( .A1(n12259), .A2(n12258), .A3(n12257), .A4(n12256), .ZN(
        n12260) );
  NOR2_X1 U15370 ( .A1(n12261), .A2(n12260), .ZN(n12267) );
  AOI22_X1 U15371 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n11980), .B1(
        n14867), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U15372 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n12026), .B1(
        n12027), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12264) );
  AOI22_X1 U15373 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12003), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12263) );
  NAND2_X1 U15374 ( .A1(n14868), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12262) );
  AND4_X1 U15375 ( .A1(n12265), .A2(n12264), .A3(n12263), .A4(n12262), .ZN(
        n12266) );
  NAND2_X1 U15376 ( .A1(n11995), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n12269) );
  AOI22_X1 U15377 ( .A1(n12000), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12279), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12268) );
  OAI211_X1 U15378 ( .C1(n13530), .C2(n12270), .A(n12269), .B(n12268), .ZN(
        n16221) );
  NAND2_X1 U15379 ( .A1(n11995), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n12272) );
  AOI22_X1 U15380 ( .A1(n12137), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12279), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12271) );
  NAND2_X1 U15381 ( .A1(n12272), .A2(n12271), .ZN(n15778) );
  NAND2_X1 U15382 ( .A1(n11995), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U15383 ( .A1(n12000), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12282), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12273) );
  AND2_X1 U15384 ( .A1(n12274), .A2(n12273), .ZN(n15125) );
  NAND2_X1 U15385 ( .A1(n11995), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n12276) );
  AOI22_X1 U15386 ( .A1(n12000), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12279), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12275) );
  NAND2_X1 U15387 ( .A1(n11995), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12278) );
  AOI22_X1 U15388 ( .A1(n12137), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12279), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12277) );
  NAND2_X1 U15389 ( .A1(n12278), .A2(n12277), .ZN(n15118) );
  INV_X1 U15390 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n12659) );
  INV_X1 U15391 ( .A(n12279), .ZN(n12292) );
  OAI22_X1 U15392 ( .A1(n12044), .A2(n12659), .B1(n12292), .B2(n15419), .ZN(
        n12280) );
  AOI21_X1 U15393 ( .B1(n11995), .B2(P2_REIP_REG_20__SCAN_IN), .A(n12280), 
        .ZN(n15421) );
  INV_X1 U15394 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n19073) );
  INV_X1 U15395 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15205) );
  OAI22_X1 U15396 ( .A1(n12044), .A2(n19073), .B1(n12292), .B2(n15205), .ZN(
        n12281) );
  AOI21_X1 U15397 ( .B1(n11995), .B2(P2_REIP_REG_21__SCAN_IN), .A(n12281), 
        .ZN(n12393) );
  NAND2_X1 U15398 ( .A1(n11995), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12284) );
  AOI22_X1 U15399 ( .A1(n12137), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12282), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12283) );
  NAND2_X1 U15400 ( .A1(n12284), .A2(n12283), .ZN(n15388) );
  INV_X1 U15401 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n19070) );
  INV_X1 U15402 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n13910) );
  OAI22_X1 U15403 ( .A1(n12044), .A2(n19070), .B1(n12292), .B2(n13910), .ZN(
        n12285) );
  AOI21_X1 U15404 ( .B1(n11995), .B2(P2_REIP_REG_23__SCAN_IN), .A(n12285), 
        .ZN(n12406) );
  OR2_X2 U15405 ( .A1(n15391), .A2(n12406), .ZN(n15098) );
  INV_X1 U15406 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n15101) );
  OAI22_X1 U15407 ( .A1(n12044), .A2(n15101), .B1(n12292), .B2(n10017), .ZN(
        n12286) );
  AOI21_X1 U15408 ( .B1(n11995), .B2(P2_REIP_REG_24__SCAN_IN), .A(n12286), 
        .ZN(n15097) );
  NOR2_X4 U15409 ( .A1(n15098), .A2(n15097), .ZN(n15100) );
  NAND2_X1 U15410 ( .A1(n11995), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12288) );
  AOI22_X1 U15411 ( .A1(n12000), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12279), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12287) );
  NAND2_X1 U15412 ( .A1(n12288), .A2(n12287), .ZN(n14726) );
  NAND2_X1 U15413 ( .A1(n11995), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12290) );
  AOI22_X1 U15414 ( .A1(n12137), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12279), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12289) );
  NAND2_X1 U15415 ( .A1(n12290), .A2(n12289), .ZN(n14710) );
  INV_X1 U15416 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n19063) );
  OAI22_X1 U15417 ( .A1(n12044), .A2(n19063), .B1(n12292), .B2(n15323), .ZN(
        n12291) );
  AOI21_X1 U15418 ( .B1(n11995), .B2(P2_REIP_REG_27__SCAN_IN), .A(n12291), 
        .ZN(n14698) );
  INV_X1 U15419 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n19061) );
  OAI22_X1 U15420 ( .A1(n12044), .A2(n19061), .B1(n12292), .B2(n15313), .ZN(
        n12293) );
  AOI21_X1 U15421 ( .B1(n11995), .B2(P2_REIP_REG_28__SCAN_IN), .A(n12293), 
        .ZN(n12380) );
  NAND2_X1 U15422 ( .A1(n11995), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n12295) );
  AOI22_X1 U15423 ( .A1(n12000), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n12279), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12294) );
  NAND2_X1 U15424 ( .A1(n12295), .A2(n12294), .ZN(n14680) );
  AOI21_X1 U15425 ( .B1(n12296), .B2(n14684), .A(n14030), .ZN(n15066) );
  INV_X1 U15426 ( .A(n12297), .ZN(n16295) );
  NAND2_X1 U15427 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19721), .ZN(n19872) );
  NOR2_X1 U15428 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n18774) );
  INV_X1 U15429 ( .A(n18774), .ZN(n19727) );
  NAND2_X1 U15430 ( .A1(n19866), .A2(n19859), .ZN(n13312) );
  NOR2_X1 U15431 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n13312), .ZN(n16294) );
  INV_X1 U15432 ( .A(n16294), .ZN(n12298) );
  MUX2_X1 U15433 ( .A(n12299), .B(n12504), .S(n12581), .Z(n12557) );
  MUX2_X1 U15434 ( .A(n12557), .B(n11829), .S(n13916), .Z(n12589) );
  NAND2_X1 U15435 ( .A1(n13916), .A2(n13199), .ZN(n12584) );
  NAND2_X1 U15436 ( .A1(n12589), .A2(n12590), .ZN(n13086) );
  MUX2_X1 U15437 ( .A(n10101), .B(n12300), .S(n12581), .Z(n12301) );
  MUX2_X1 U15438 ( .A(n13491), .B(n12304), .S(n12581), .Z(n12305) );
  MUX2_X1 U15439 ( .A(n12305), .B(n11848), .S(n13916), .Z(n13479) );
  MUX2_X1 U15440 ( .A(n12307), .B(n12306), .S(n19177), .Z(n13571) );
  MUX2_X1 U15441 ( .A(n13679), .B(P2_EBX_REG_6__SCAN_IN), .S(n19177), .Z(
        n12919) );
  MUX2_X1 U15442 ( .A(n13698), .B(n12308), .S(n19177), .Z(n13115) );
  AND2_X1 U15443 ( .A1(n19177), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13140) );
  NAND2_X1 U15444 ( .A1(n13916), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13846) );
  AND2_X1 U15445 ( .A1(n19177), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13852) );
  AND2_X1 U15446 ( .A1(n19177), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n13873) );
  NAND2_X1 U15447 ( .A1(n13916), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n13877) );
  NAND2_X1 U15448 ( .A1(n13916), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13869) );
  AND2_X1 U15449 ( .A1(n19177), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n13861) );
  AND2_X1 U15450 ( .A1(n19177), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n13860) );
  INV_X1 U15451 ( .A(n13860), .ZN(n12309) );
  INV_X1 U15452 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n12310) );
  NAND2_X1 U15453 ( .A1(n13916), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n13901) );
  AND2_X1 U15454 ( .A1(n19177), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12402) );
  NAND2_X1 U15455 ( .A1(n13916), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n13815) );
  AND2_X1 U15456 ( .A1(n19177), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12376) );
  NAND2_X1 U15457 ( .A1(n13916), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n13927) );
  NAND2_X1 U15458 ( .A1(n13926), .A2(n13927), .ZN(n14010) );
  NAND2_X1 U15459 ( .A1(n13916), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12311) );
  XNOR2_X1 U15460 ( .A(n14010), .B(n12311), .ZN(n13930) );
  INV_X1 U15461 ( .A(n13930), .ZN(n13931) );
  INV_X1 U15462 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n14742) );
  NOR2_X1 U15463 ( .A1(n12318), .A2(n14742), .ZN(n12312) );
  NAND2_X1 U15464 ( .A1(n11776), .A2(n12312), .ZN(n12313) );
  NOR2_X2 U15465 ( .A1(n19855), .A2(n12313), .ZN(n18958) );
  NOR2_X1 U15466 ( .A1(n13931), .A2(n18941), .ZN(n12314) );
  OR2_X1 U15467 ( .A1(n19051), .A2(n16294), .ZN(n14664) );
  AND2_X1 U15468 ( .A1(n12317), .A2(n12435), .ZN(n12447) );
  NOR2_X1 U15469 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n12318), .ZN(n12319) );
  NAND2_X1 U15470 ( .A1(n12447), .A2(n12319), .ZN(n12320) );
  NAND2_X1 U15471 ( .A1(n14664), .A2(n12320), .ZN(n18898) );
  INV_X1 U15472 ( .A(n18963), .ZN(n18923) );
  INV_X1 U15473 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n13951) );
  NOR2_X1 U15474 ( .A1(n10098), .A2(n12321), .ZN(n12322) );
  NAND3_X1 U15475 ( .A1(n12324), .A2(n12323), .A3(n12322), .ZN(P2_U2825) );
  OR2_X1 U15476 ( .A1(n12325), .A2(n19878), .ZN(n12326) );
  NOR2_X1 U15477 ( .A1(n12327), .A2(n12326), .ZN(n12328) );
  NAND3_X1 U15478 ( .A1(n20649), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16121) );
  INV_X1 U15479 ( .A(n16121), .ZN(n12329) );
  NOR2_X1 U15480 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20738) );
  INV_X1 U15481 ( .A(n20586), .ZN(n20369) );
  AND2_X1 U15482 ( .A1(n12329), .A2(n20369), .ZN(n14447) );
  NAND2_X1 U15483 ( .A1(n14043), .A2(n14447), .ZN(n12340) );
  NAND2_X1 U15484 ( .A1(n20586), .A2(n12330), .ZN(n20755) );
  AND2_X1 U15485 ( .A1(n20755), .A2(n20649), .ZN(n12331) );
  NAND2_X1 U15486 ( .A1(n20649), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15824) );
  NAND2_X1 U15487 ( .A1(n20515), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12332) );
  AND2_X1 U15488 ( .A1(n15824), .A2(n12332), .ZN(n20025) );
  INV_X1 U15489 ( .A(n20025), .ZN(n12333) );
  NOR2_X1 U15490 ( .A1(n12334), .A2(n20880), .ZN(n12335) );
  XNOR2_X1 U15491 ( .A(n12335), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13457) );
  AOI21_X1 U15492 ( .B1(n20013), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n12336), .ZN(n12337) );
  OAI21_X1 U15493 ( .B1(n20023), .B2(n13457), .A(n12337), .ZN(n12338) );
  OAI211_X1 U15494 ( .C1(n12341), .C2(n20030), .A(n12340), .B(n12339), .ZN(
        P1_U2968) );
  NOR2_X1 U15495 ( .A1(n16461), .A2(n12342), .ZN(n18533) );
  INV_X1 U15496 ( .A(n18763), .ZN(n18713) );
  NAND2_X1 U15497 ( .A1(n18762), .A2(n20828), .ZN(n16456) );
  AND2_X1 U15498 ( .A1(n18713), .A2(n16456), .ZN(n18744) );
  NAND2_X1 U15499 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17671) );
  INV_X1 U15500 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16834) );
  NAND2_X1 U15501 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17725) );
  NAND2_X1 U15502 ( .A1(n17708), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17700) );
  NAND2_X1 U15503 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17680) );
  NOR3_X1 U15504 ( .A1(n17680), .A2(n17662), .A3(n16708), .ZN(n16693) );
  INV_X1 U15505 ( .A(n16693), .ZN(n16690) );
  INV_X1 U15506 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16701) );
  NOR2_X1 U15507 ( .A1(n16690), .A2(n16701), .ZN(n16679) );
  NAND2_X1 U15508 ( .A1(n17672), .A2(n16679), .ZN(n17636) );
  NAND2_X1 U15509 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17614) );
  NAND2_X1 U15510 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17569) );
  NAND2_X1 U15511 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17534) );
  NAND2_X1 U15512 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17499) );
  NAND2_X1 U15513 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17456) );
  NAND2_X1 U15514 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17418) );
  NAND2_X1 U15515 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n16330), .ZN(
        n12346) );
  NAND2_X1 U15516 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16327), .ZN(
        n12344) );
  NOR2_X1 U15517 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18762), .ZN(n17610) );
  INV_X1 U15518 ( .A(n17490), .ZN(n12345) );
  NOR2_X1 U15519 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20828), .ZN(
        n18725) );
  NOR2_X1 U15520 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18754) );
  AOI21_X1 U15521 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n18754), .ZN(n18609) );
  OR2_X1 U15522 ( .A1(n18725), .A2(n18609), .ZN(n18099) );
  INV_X1 U15523 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18749) );
  NOR3_X1 U15524 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n18749), .ZN(n18445) );
  NAND2_X1 U15525 ( .A1(n18396), .A2(n18445), .ZN(n18134) );
  OR2_X1 U15526 ( .A1(n12346), .A2(n17613), .ZN(n16309) );
  INV_X1 U15527 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16484) );
  XOR2_X1 U15528 ( .A(n16484), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n12348) );
  NOR2_X1 U15529 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17490), .ZN(
        n16328) );
  NOR2_X1 U15530 ( .A1(n16834), .A2(n17417), .ZN(n16479) );
  NAND3_X1 U15531 ( .A1(n16479), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16477) );
  AOI22_X1 U15532 ( .A1(n17610), .A2(n16477), .B1(n18478), .B2(n12346), .ZN(
        n12347) );
  NAND2_X1 U15533 ( .A1(n12347), .A2(n17764), .ZN(n16329) );
  NOR2_X1 U15534 ( .A1(n16328), .A2(n16329), .ZN(n16308) );
  OAI22_X1 U15535 ( .A1(n16309), .A2(n12348), .B1(n16308), .B2(n16484), .ZN(
        n12349) );
  AOI211_X1 U15536 ( .C1(n17532), .C2(n9795), .A(n12350), .B(n12349), .ZN(
        n12351) );
  INV_X1 U15537 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20754) );
  NOR3_X1 U15538 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20754), .ZN(n12360) );
  NOR4_X1 U15539 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12359) );
  NAND4_X1 U15540 ( .A1(n13387), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12360), .A4(
        n12359), .ZN(U214) );
  NOR4_X1 U15541 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12364) );
  NOR4_X1 U15542 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12363) );
  NOR4_X1 U15543 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12362) );
  NOR4_X1 U15544 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12361) );
  NAND4_X1 U15545 ( .A1(n12364), .A2(n12363), .A3(n12362), .A4(n12361), .ZN(
        n12369) );
  NOR4_X1 U15546 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_19__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n12367) );
  NOR4_X1 U15547 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n12366) );
  NOR4_X1 U15548 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n12365) );
  INV_X1 U15549 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19738) );
  NAND4_X1 U15550 ( .A1(n12367), .A2(n12366), .A3(n12365), .A4(n19738), .ZN(
        n12368) );
  OAI21_X1 U15551 ( .B1(n12369), .B2(n12368), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12370) );
  INV_X2 U15552 ( .A(n15064), .ZN(n15061) );
  NOR2_X1 U15553 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12372) );
  NOR4_X1 U15554 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12371) );
  NAND4_X1 U15555 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12372), .A4(n12371), .ZN(n12387) );
  NOR2_X1 U15556 ( .A1(n15061), .A2(n12387), .ZN(n16357) );
  NAND2_X1 U15557 ( .A1(n16357), .A2(U214), .ZN(U212) );
  AOI211_X1 U15558 ( .C1(n12375), .C2(n12373), .A(n12374), .B(n19713), .ZN(
        n12386) );
  AOI21_X1 U15559 ( .B1(n12376), .B2(n13818), .A(n13926), .ZN(n13922) );
  INV_X1 U15560 ( .A(n13922), .ZN(n12377) );
  INV_X1 U15561 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19779) );
  OAI22_X1 U15562 ( .A1(n12377), .A2(n18941), .B1(n19779), .B2(n18923), .ZN(
        n12385) );
  AOI22_X1 U15563 ( .A1(n18898), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n18957), .ZN(n12378) );
  INV_X1 U15564 ( .A(n12378), .ZN(n12384) );
  OAI21_X1 U15565 ( .B1(n14693), .B2(n12379), .A(n14673), .ZN(n14994) );
  AND2_X1 U15566 ( .A1(n14700), .A2(n12380), .ZN(n12381) );
  NOR2_X1 U15567 ( .A1(n14679), .A2(n12381), .ZN(n15311) );
  INV_X1 U15568 ( .A(n15311), .ZN(n12382) );
  OAI22_X1 U15569 ( .A1(n14994), .A2(n18965), .B1(n12382), .B2(n18960), .ZN(
        n12383) );
  NOR2_X1 U15570 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12387), .ZN(n16447)
         );
  AOI211_X1 U15571 ( .C1(n15208), .C2(n12389), .A(n12388), .B(n19713), .ZN(
        n12399) );
  INV_X1 U15572 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19767) );
  OAI22_X1 U15573 ( .A1(n13882), .A2(n18941), .B1(n19767), .B2(n18923), .ZN(
        n12398) );
  OAI22_X1 U15574 ( .A1(n18961), .A2(n11898), .B1(n15206), .B2(n18955), .ZN(
        n12397) );
  NAND2_X1 U15575 ( .A1(n15042), .A2(n12391), .ZN(n12392) );
  NAND2_X1 U15576 ( .A1(n9648), .A2(n12392), .ZN(n15402) );
  AND2_X1 U15577 ( .A1(n15424), .A2(n12393), .ZN(n12394) );
  NOR2_X1 U15578 ( .A1(n15389), .A2(n12394), .ZN(n15399) );
  INV_X1 U15579 ( .A(n15399), .ZN(n12395) );
  OAI22_X1 U15580 ( .A1(n15402), .A2(n18965), .B1(n18960), .B2(n12395), .ZN(
        n12396) );
  OR4_X1 U15581 ( .A1(n12399), .A2(n12398), .A3(n12397), .A4(n12396), .ZN(
        P2_U2834) );
  AOI211_X1 U15582 ( .C1(n15188), .C2(n12401), .A(n12400), .B(n19713), .ZN(
        n12412) );
  NAND2_X1 U15583 ( .A1(n13904), .A2(n12402), .ZN(n12403) );
  AND2_X1 U15584 ( .A1(n13913), .A2(n12403), .ZN(n13908) );
  INV_X1 U15585 ( .A(n13908), .ZN(n13911) );
  OAI22_X1 U15586 ( .A1(n13911), .A2(n18941), .B1(n18961), .B2(n11903), .ZN(
        n12411) );
  OAI22_X1 U15587 ( .A1(n20877), .A2(n18955), .B1(n20860), .B2(n18923), .ZN(
        n12410) );
  NOR2_X1 U15588 ( .A1(n15027), .A2(n12404), .ZN(n12405) );
  OR2_X1 U15589 ( .A1(n15020), .A2(n12405), .ZN(n15379) );
  NAND2_X1 U15590 ( .A1(n15391), .A2(n12406), .ZN(n12407) );
  AND2_X1 U15591 ( .A1(n15098), .A2(n12407), .ZN(n15377) );
  INV_X1 U15592 ( .A(n15377), .ZN(n12408) );
  OAI22_X1 U15593 ( .A1(n15379), .A2(n18965), .B1(n18960), .B2(n12408), .ZN(
        n12409) );
  OR4_X1 U15594 ( .A1(n12412), .A2(n12411), .A3(n12410), .A4(n12409), .ZN(
        P2_U2832) );
  NOR3_X1 U15595 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16807) );
  NAND2_X1 U15596 ( .A1(n16807), .A2(n16801), .ZN(n16800) );
  NOR2_X1 U15597 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16800), .ZN(n16779) );
  INV_X1 U15598 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16775) );
  NAND2_X1 U15599 ( .A1(n16779), .A2(n16775), .ZN(n16772) );
  NOR2_X1 U15600 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16772), .ZN(n16752) );
  INV_X1 U15601 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16749) );
  NAND2_X1 U15602 ( .A1(n16752), .A2(n16749), .ZN(n16748) );
  INV_X1 U15603 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17049) );
  NAND2_X1 U15604 ( .A1(n16725), .A2(n17049), .ZN(n16722) );
  INV_X1 U15605 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17064) );
  NAND2_X1 U15606 ( .A1(n16704), .A2(n17064), .ZN(n16698) );
  INV_X1 U15607 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16676) );
  NAND2_X1 U15608 ( .A1(n16681), .A2(n16676), .ZN(n16668) );
  INV_X1 U15609 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17018) );
  NAND2_X1 U15610 ( .A1(n16656), .A2(n17018), .ZN(n16645) );
  INV_X1 U15611 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16623) );
  NAND2_X1 U15612 ( .A1(n16631), .A2(n16623), .ZN(n16622) );
  INV_X1 U15613 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16599) );
  NAND2_X1 U15614 ( .A1(n16608), .A2(n16599), .ZN(n16598) );
  INV_X1 U15615 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16936) );
  NAND2_X1 U15616 ( .A1(n16584), .A2(n16936), .ZN(n16578) );
  NOR2_X1 U15617 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16578), .ZN(n16563) );
  INV_X1 U15618 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16847) );
  NAND2_X1 U15619 ( .A1(n16563), .A2(n16847), .ZN(n16558) );
  NOR2_X1 U15620 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16558), .ZN(n16544) );
  INV_X1 U15621 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16536) );
  NAND2_X1 U15622 ( .A1(n16544), .A2(n16536), .ZN(n16535) );
  NOR2_X1 U15623 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16535), .ZN(n16529) );
  NAND2_X1 U15624 ( .A1(n18536), .A2(n18745), .ZN(n17301) );
  NAND2_X1 U15625 ( .A1(n18749), .A2(n18751), .ZN(n12413) );
  AOI211_X1 U15626 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16535), .A(n16529), .B(
        n16838), .ZN(n12433) );
  INV_X1 U15627 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n20831) );
  INV_X1 U15628 ( .A(n18751), .ZN(n18602) );
  AOI211_X1 U15629 ( .C1(n18750), .C2(n18748), .A(n18602), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18592) );
  INV_X1 U15630 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n20818) );
  INV_X1 U15631 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18664) );
  INV_X1 U15632 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18662) );
  INV_X1 U15633 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18647) );
  INV_X1 U15634 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18636) );
  NAND2_X1 U15635 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16812) );
  NOR2_X1 U15636 ( .A1(n18636), .A2(n16812), .ZN(n16792) );
  AND2_X1 U15637 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16792), .ZN(n16767) );
  NAND2_X1 U15638 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16767), .ZN(n16742) );
  INV_X1 U15639 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18644) );
  INV_X1 U15640 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18642) );
  NOR4_X1 U15641 ( .A1(n18647), .A2(n16742), .A3(n18644), .A4(n18642), .ZN(
        n16702) );
  INV_X1 U15642 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18650) );
  INV_X1 U15643 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18648) );
  NOR2_X1 U15644 ( .A1(n18650), .A2(n18648), .ZN(n16689) );
  NAND3_X1 U15645 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16702), .A3(n16689), 
        .ZN(n16663) );
  INV_X1 U15646 ( .A(n16663), .ZN(n16683) );
  NAND2_X1 U15647 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16683), .ZN(n16652) );
  NAND2_X1 U15648 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .ZN(n16618) );
  NOR2_X1 U15649 ( .A1(n16652), .A2(n16618), .ZN(n16655) );
  NAND2_X1 U15650 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16655), .ZN(n16627) );
  NOR3_X1 U15651 ( .A1(n18664), .A2(n18662), .A3(n16627), .ZN(n16591) );
  AND4_X1 U15652 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .A3(P3_REIP_REG_18__SCAN_IN), .A4(n16591), .ZN(n16572) );
  NAND3_X1 U15653 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(P3_REIP_REG_22__SCAN_IN), 
        .A3(n16572), .ZN(n16554) );
  NOR2_X1 U15654 ( .A1(n20818), .A2(n16554), .ZN(n16543) );
  AND2_X1 U15655 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16543), .ZN(n16537) );
  NAND2_X1 U15656 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16537), .ZN(n12415) );
  OR2_X1 U15657 ( .A1(n16831), .A2(n12415), .ZN(n16482) );
  NAND4_X1 U15658 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18762), .A3(n12414), 
        .A4(n18749), .ZN(n18608) );
  NOR2_X1 U15659 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n20828), .ZN(n18603) );
  INV_X1 U15660 ( .A(n18603), .ZN(n18472) );
  OR2_X1 U15661 ( .A1(n18605), .A2(n18472), .ZN(n18598) );
  INV_X1 U15662 ( .A(n16842), .ZN(n16826) );
  AOI221_X1 U15663 ( .B1(n20831), .B2(n16813), .C1(n12415), .C2(n16813), .A(
        n16826), .ZN(n16532) );
  AOI21_X1 U15664 ( .B1(n20831), .B2(n16482), .A(n16532), .ZN(n12432) );
  NOR2_X1 U15665 ( .A1(n16834), .A2(n17455), .ZN(n12419) );
  INV_X1 U15666 ( .A(n12419), .ZN(n12416) );
  NOR2_X1 U15667 ( .A1(n17456), .A2(n12416), .ZN(n17412) );
  INV_X1 U15668 ( .A(n16479), .ZN(n16480) );
  OAI21_X1 U15669 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17412), .A(
        n16480), .ZN(n17443) );
  INV_X1 U15670 ( .A(n17443), .ZN(n12427) );
  INV_X1 U15671 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12417) );
  NAND2_X1 U15672 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n12419), .ZN(
        n12418) );
  AOI21_X1 U15673 ( .B1(n12417), .B2(n12418), .A(n17412), .ZN(n17448) );
  OAI21_X1 U15674 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n12419), .A(
        n12418), .ZN(n17472) );
  INV_X1 U15675 ( .A(n17472), .ZN(n16547) );
  NOR2_X1 U15676 ( .A1(n16834), .A2(n17498), .ZN(n12423) );
  INV_X1 U15677 ( .A(n12423), .ZN(n12424) );
  NOR2_X1 U15678 ( .A1(n17499), .A2(n12424), .ZN(n12420) );
  INV_X1 U15679 ( .A(n12420), .ZN(n17447) );
  AOI21_X1 U15680 ( .B1(n9806), .B2(n17447), .A(n12419), .ZN(n17473) );
  INV_X1 U15681 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12421) );
  NAND2_X1 U15682 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n12423), .ZN(
        n12422) );
  AOI21_X1 U15683 ( .B1(n12421), .B2(n12422), .A(n12420), .ZN(n17491) );
  OAI21_X1 U15684 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n12423), .A(
        n12422), .ZN(n17516) );
  INV_X1 U15685 ( .A(n17516), .ZN(n16575) );
  AND2_X1 U15686 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17517), .ZN(
        n17488) );
  OAI21_X1 U15687 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17488), .A(
        n12424), .ZN(n12425) );
  INV_X1 U15688 ( .A(n12425), .ZN(n17519) );
  NOR2_X1 U15689 ( .A1(n16834), .A2(n17636), .ZN(n17612) );
  INV_X1 U15690 ( .A(n17612), .ZN(n16691) );
  NOR2_X1 U15691 ( .A1(n17614), .A2(n16691), .ZN(n16664) );
  NAND2_X1 U15692 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n16664), .ZN(
        n16650) );
  INV_X1 U15693 ( .A(n16650), .ZN(n17567) );
  NAND2_X1 U15694 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17567), .ZN(
        n16639) );
  NOR2_X1 U15695 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16639), .ZN(
        n16638) );
  NOR2_X1 U15696 ( .A1(n16573), .A2(n9794), .ZN(n16565) );
  NOR2_X1 U15697 ( .A1(n17491), .A2(n16565), .ZN(n16564) );
  NOR2_X1 U15698 ( .A1(n16564), .A2(n9794), .ZN(n16553) );
  NOR2_X1 U15699 ( .A1(n17473), .A2(n16553), .ZN(n16552) );
  NOR2_X1 U15700 ( .A1(n16552), .A2(n9794), .ZN(n16546) );
  NOR2_X1 U15701 ( .A1(n16547), .A2(n16546), .ZN(n16545) );
  AOI211_X1 U15702 ( .C1(n12427), .C2(n12426), .A(n16481), .B(n18608), .ZN(
        n12431) );
  INV_X1 U15703 ( .A(n12428), .ZN(n12429) );
  INV_X1 U15704 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n16894) );
  OAI22_X1 U15705 ( .A1(n9807), .A2(n16827), .B1(n16830), .B2(n16894), .ZN(
        n12430) );
  OR4_X1 U15706 ( .A1(n12433), .A2(n12432), .A3(n12431), .A4(n12430), .ZN(
        P3_U2645) );
  INV_X1 U15707 ( .A(n19050), .ZN(n12436) );
  NAND2_X1 U15708 ( .A1(n12436), .A2(n12435), .ZN(n18966) );
  INV_X1 U15709 ( .A(n18966), .ZN(n12439) );
  INV_X1 U15710 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n19874) );
  INV_X1 U15711 ( .A(n12447), .ZN(n12446) );
  AND2_X1 U15712 ( .A1(n19812), .A2(n12437), .ZN(n12441) );
  INV_X1 U15713 ( .A(n12441), .ZN(n12438) );
  OAI211_X1 U15714 ( .C1(n12439), .C2(n19874), .A(n12446), .B(n12438), .ZN(
        P2_U2814) );
  INV_X1 U15715 ( .A(n12440), .ZN(n12443) );
  OAI21_X1 U15716 ( .B1(n12441), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n19855), 
        .ZN(n12442) );
  OAI21_X1 U15717 ( .B1(n12443), .B2(n19855), .A(n12442), .ZN(P2_U3612) );
  NOR2_X1 U15718 ( .A1(n12626), .A2(n19878), .ZN(n12444) );
  NAND2_X1 U15719 ( .A1(n12625), .A2(n12763), .ZN(n12620) );
  NOR2_X1 U15720 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20586), .ZN(n12621) );
  AOI21_X1 U15721 ( .B1(n12620), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n12621), 
        .ZN(n12445) );
  NAND2_X1 U15722 ( .A1(n12704), .A2(n12445), .ZN(P1_U2801) );
  OAI21_X2 U15723 ( .B1(n12446), .B2(n19717), .A(n19051), .ZN(n12649) );
  INV_X1 U15724 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n12449) );
  INV_X1 U15725 ( .A(n19051), .ZN(n12494) );
  NAND3_X1 U15726 ( .A1(n12447), .A2(n14935), .A3(n19859), .ZN(n12501) );
  AOI22_X1 U15727 ( .A1(n15064), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n15061), .ZN(n19168) );
  NOR2_X1 U15728 ( .A1(n12501), .A2(n19168), .ZN(n12452) );
  AOI21_X1 U15729 ( .B1(P2_EAX_REG_1__SCAN_IN), .B2(n12494), .A(n12452), .ZN(
        n12448) );
  OAI21_X1 U15730 ( .B1(n12649), .B2(n12449), .A(n12448), .ZN(P2_U2968) );
  INV_X1 U15731 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n12451) );
  AOI22_X1 U15732 ( .A1(n15064), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n15061), .ZN(n19173) );
  NOR2_X1 U15733 ( .A1(n12501), .A2(n19173), .ZN(n12459) );
  AOI21_X1 U15734 ( .B1(P2_EAX_REG_3__SCAN_IN), .B2(n12494), .A(n12459), .ZN(
        n12450) );
  OAI21_X1 U15735 ( .B1(n12649), .B2(n12451), .A(n12450), .ZN(P2_U2970) );
  INV_X1 U15736 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n12454) );
  AOI21_X1 U15737 ( .B1(n12494), .B2(P2_EAX_REG_17__SCAN_IN), .A(n12452), .ZN(
        n12453) );
  OAI21_X1 U15738 ( .B1(n12649), .B2(n12454), .A(n12453), .ZN(P2_U2953) );
  INV_X1 U15739 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n12456) );
  INV_X1 U15740 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n20859) );
  INV_X1 U15741 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18108) );
  AOI22_X1 U15742 ( .A1(n15064), .A2(n20859), .B1(n18108), .B2(n15061), .ZN(
        n16152) );
  INV_X1 U15743 ( .A(n16152), .ZN(n13435) );
  NOR2_X1 U15744 ( .A1(n12501), .A2(n13435), .ZN(n12462) );
  AOI21_X1 U15745 ( .B1(P2_EAX_REG_2__SCAN_IN), .B2(n12494), .A(n12462), .ZN(
        n12455) );
  OAI21_X1 U15746 ( .B1(n12649), .B2(n12456), .A(n12455), .ZN(P2_U2969) );
  INV_X1 U15747 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n12458) );
  AOI22_X1 U15748 ( .A1(n15064), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n15061), .ZN(n19178) );
  NOR2_X1 U15749 ( .A1(n12501), .A2(n19178), .ZN(n12465) );
  AOI21_X1 U15750 ( .B1(P2_EAX_REG_5__SCAN_IN), .B2(n12494), .A(n12465), .ZN(
        n12457) );
  OAI21_X1 U15751 ( .B1(n12649), .B2(n12458), .A(n12457), .ZN(P2_U2972) );
  INV_X1 U15752 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n12461) );
  AOI21_X1 U15753 ( .B1(n12494), .B2(P2_EAX_REG_19__SCAN_IN), .A(n12459), .ZN(
        n12460) );
  OAI21_X1 U15754 ( .B1(n12649), .B2(n12461), .A(n12460), .ZN(P2_U2955) );
  INV_X1 U15755 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n12464) );
  AOI21_X1 U15756 ( .B1(P2_EAX_REG_18__SCAN_IN), .B2(n12494), .A(n12462), .ZN(
        n12463) );
  OAI21_X1 U15757 ( .B1(n12649), .B2(n12464), .A(n12463), .ZN(P2_U2954) );
  INV_X1 U15758 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n12467) );
  AOI21_X1 U15759 ( .B1(n12494), .B2(P2_EAX_REG_21__SCAN_IN), .A(n12465), .ZN(
        n12466) );
  OAI21_X1 U15760 ( .B1(n12649), .B2(n12467), .A(n12466), .ZN(P2_U2957) );
  INV_X1 U15761 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n12473) );
  INV_X1 U15762 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n12468) );
  OR2_X1 U15763 ( .A1(n15061), .A2(n12468), .ZN(n12470) );
  NAND2_X1 U15764 ( .A1(n15061), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12469) );
  AND2_X1 U15765 ( .A1(n12470), .A2(n12469), .ZN(n19000) );
  INV_X1 U15766 ( .A(n19000), .ZN(n12471) );
  NAND2_X1 U15767 ( .A1(n12674), .A2(n12471), .ZN(n12650) );
  NAND2_X1 U15768 ( .A1(n12494), .A2(P2_EAX_REG_11__SCAN_IN), .ZN(n12472) );
  OAI211_X1 U15769 ( .C1(n12649), .C2(n12473), .A(n12650), .B(n12472), .ZN(
        P2_U2978) );
  INV_X1 U15770 ( .A(P2_LWORD_REG_12__SCAN_IN), .ZN(n12479) );
  INV_X1 U15771 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n12474) );
  OR2_X1 U15772 ( .A1(n15061), .A2(n12474), .ZN(n12476) );
  NAND2_X1 U15773 ( .A1(n15061), .A2(BUF2_REG_12__SCAN_IN), .ZN(n12475) );
  AND2_X1 U15774 ( .A1(n12476), .A2(n12475), .ZN(n18998) );
  INV_X1 U15775 ( .A(n18998), .ZN(n12477) );
  NAND2_X1 U15776 ( .A1(n12674), .A2(n12477), .ZN(n12676) );
  NAND2_X1 U15777 ( .A1(n12494), .A2(P2_EAX_REG_12__SCAN_IN), .ZN(n12478) );
  OAI211_X1 U15778 ( .C1(n12649), .C2(n12479), .A(n12676), .B(n12478), .ZN(
        P2_U2979) );
  INV_X1 U15779 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n12482) );
  AOI22_X1 U15780 ( .A1(n15064), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n15061), .ZN(n19188) );
  INV_X1 U15781 ( .A(n19188), .ZN(n12480) );
  NAND2_X1 U15782 ( .A1(n12674), .A2(n12480), .ZN(n12664) );
  NAND2_X1 U15783 ( .A1(n12494), .A2(P2_EAX_REG_7__SCAN_IN), .ZN(n12481) );
  OAI211_X1 U15784 ( .C1(n12649), .C2(n12482), .A(n12664), .B(n12481), .ZN(
        P2_U2974) );
  INV_X1 U15785 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n12487) );
  OR2_X1 U15786 ( .A1(n15061), .A2(n16389), .ZN(n12484) );
  NAND2_X1 U15787 ( .A1(n15061), .A2(BUF2_REG_13__SCAN_IN), .ZN(n12483) );
  AND2_X1 U15788 ( .A1(n12484), .A2(n12483), .ZN(n18996) );
  INV_X1 U15789 ( .A(n18996), .ZN(n12485) );
  NAND2_X1 U15790 ( .A1(n12674), .A2(n12485), .ZN(n12656) );
  NAND2_X1 U15791 ( .A1(n12494), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n12486) );
  OAI211_X1 U15792 ( .C1(n12649), .C2(n12487), .A(n12656), .B(n12486), .ZN(
        P2_U2980) );
  INV_X1 U15793 ( .A(P2_LWORD_REG_9__SCAN_IN), .ZN(n12493) );
  INV_X1 U15794 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n12488) );
  OR2_X1 U15795 ( .A1(n15061), .A2(n12488), .ZN(n12490) );
  NAND2_X1 U15796 ( .A1(n15061), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12489) );
  AND2_X1 U15797 ( .A1(n12490), .A2(n12489), .ZN(n19005) );
  INV_X1 U15798 ( .A(n19005), .ZN(n12491) );
  NAND2_X1 U15799 ( .A1(n12674), .A2(n12491), .ZN(n12669) );
  NAND2_X1 U15800 ( .A1(n12494), .A2(P2_EAX_REG_9__SCAN_IN), .ZN(n12492) );
  OAI211_X1 U15801 ( .C1(n12649), .C2(n12493), .A(n12669), .B(n12492), .ZN(
        P2_U2976) );
  INV_X1 U15802 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n12496) );
  OAI22_X1 U15803 ( .A1(n15061), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n15064), .ZN(n19182) );
  INV_X1 U15804 ( .A(n19182), .ZN(n16141) );
  NAND2_X1 U15805 ( .A1(n12674), .A2(n16141), .ZN(n12666) );
  NAND2_X1 U15806 ( .A1(n12494), .A2(P2_EAX_REG_6__SCAN_IN), .ZN(n12495) );
  OAI211_X1 U15807 ( .C1(n12649), .C2(n12496), .A(n12666), .B(n12495), .ZN(
        P2_U2973) );
  INV_X1 U15808 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n12497) );
  INV_X1 U15809 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n19083) );
  INV_X1 U15810 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16414) );
  INV_X1 U15811 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18098) );
  AOI22_X1 U15812 ( .A1(n15064), .A2(n16414), .B1(n18098), .B2(n15061), .ZN(
        n18978) );
  INV_X1 U15813 ( .A(n18978), .ZN(n13238) );
  OAI222_X1 U15814 ( .A1(n12497), .A2(n12649), .B1(n19051), .B2(n19083), .C1(
        n13238), .C2(n12501), .ZN(P2_U2952) );
  INV_X1 U15815 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n12499) );
  INV_X1 U15816 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n12498) );
  OAI222_X1 U15817 ( .A1(n12499), .A2(n12649), .B1(n12501), .B2(n13238), .C1(
        n19051), .C2(n12498), .ZN(P2_U2967) );
  INV_X1 U15818 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n12502) );
  AOI22_X1 U15819 ( .A1(n15064), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n15061), .ZN(n18991) );
  INV_X1 U15820 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n12500) );
  OAI222_X1 U15821 ( .A1(n12502), .A2(n12649), .B1(n12501), .B2(n18991), .C1(
        n19051), .C2(n12500), .ZN(P2_U2982) );
  OR2_X1 U15822 ( .A1(n19050), .A2(n13312), .ZN(n12543) );
  NAND2_X1 U15823 ( .A1(n19860), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19864) );
  NAND2_X1 U15824 ( .A1(n19864), .A2(n14935), .ZN(n12503) );
  MUX2_X1 U15825 ( .A(n12503), .B(n12581), .S(n12504), .Z(n12513) );
  INV_X1 U15826 ( .A(n12504), .ZN(n12511) );
  OAI21_X1 U15827 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19839), .A(
        n12505), .ZN(n12582) );
  OAI21_X1 U15828 ( .B1(n12582), .B2(n12506), .A(n11776), .ZN(n12509) );
  INV_X1 U15829 ( .A(n12582), .ZN(n12553) );
  OAI211_X1 U15830 ( .C1(n14935), .C2(n12553), .A(n13344), .B(n12507), .ZN(
        n12508) );
  OAI211_X1 U15831 ( .C1(n12511), .C2(n12510), .A(n12509), .B(n12508), .ZN(
        n12512) );
  NAND2_X1 U15832 ( .A1(n12513), .A2(n12512), .ZN(n12514) );
  NAND2_X1 U15833 ( .A1(n12514), .A2(n12555), .ZN(n12517) );
  INV_X1 U15834 ( .A(n12555), .ZN(n12515) );
  NAND2_X1 U15835 ( .A1(n12515), .A2(n12581), .ZN(n12516) );
  NAND2_X1 U15836 ( .A1(n12517), .A2(n12516), .ZN(n12518) );
  NAND2_X1 U15837 ( .A1(n12518), .A2(n12522), .ZN(n12519) );
  NAND2_X1 U15838 ( .A1(n12519), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12521) );
  NAND2_X1 U15839 ( .A1(n11587), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12520) );
  NAND2_X1 U15840 ( .A1(n16269), .A2(n14935), .ZN(n19053) );
  NAND2_X1 U15841 ( .A1(n12525), .A2(n13436), .ZN(n12526) );
  NAND2_X1 U15842 ( .A1(n19050), .A2(n12526), .ZN(n12531) );
  NOR2_X1 U15843 ( .A1(n13345), .A2(n14935), .ZN(n12532) );
  OAI211_X1 U15844 ( .C1(n12532), .C2(n19860), .A(n11768), .B(n12772), .ZN(
        n12527) );
  NAND2_X1 U15845 ( .A1(n12527), .A2(n13436), .ZN(n12530) );
  NAND2_X1 U15846 ( .A1(n12528), .A2(n12772), .ZN(n12529) );
  NOR2_X1 U15847 ( .A1(n13344), .A2(n19865), .ZN(n12559) );
  NAND2_X1 U15848 ( .A1(n12529), .A2(n12559), .ZN(n13337) );
  NAND4_X1 U15849 ( .A1(n12524), .A2(n12531), .A3(n12530), .A4(n13337), .ZN(
        n12540) );
  INV_X1 U15850 ( .A(n12532), .ZN(n12533) );
  NOR2_X1 U15851 ( .A1(n12540), .A2(n12533), .ZN(n16274) );
  NAND2_X1 U15852 ( .A1(n16269), .A2(n16274), .ZN(n12535) );
  AND2_X1 U15853 ( .A1(n12440), .A2(n19859), .ZN(n16281) );
  NAND3_X1 U15854 ( .A1(n11807), .A2(n16271), .A3(n16281), .ZN(n12534) );
  NAND2_X1 U15855 ( .A1(n12535), .A2(n12534), .ZN(n12687) );
  INV_X1 U15856 ( .A(n12687), .ZN(n12542) );
  NAND2_X1 U15857 ( .A1(n12536), .A2(n12537), .ZN(n16272) );
  OR2_X1 U15858 ( .A1(n16269), .A2(n16272), .ZN(n12770) );
  OR2_X1 U15859 ( .A1(n11789), .A2(n13312), .ZN(n12538) );
  INV_X1 U15860 ( .A(n16271), .ZN(n16279) );
  NOR2_X1 U15861 ( .A1(n12538), .A2(n16279), .ZN(n12539) );
  NOR2_X1 U15862 ( .A1(n12540), .A2(n12539), .ZN(n13322) );
  AND2_X1 U15863 ( .A1(n12770), .A2(n13322), .ZN(n12541) );
  OAI211_X1 U15864 ( .C1(n12543), .C2(n19053), .A(n12542), .B(n12541), .ZN(
        n16285) );
  NAND2_X1 U15865 ( .A1(n16285), .A2(n19708), .ZN(n12545) );
  NAND2_X1 U15866 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19831) );
  NOR2_X1 U15867 ( .A1(n11587), .A2(n19831), .ZN(n16304) );
  AOI22_X1 U15868 ( .A1(n11587), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n16304), 
        .B2(P2_FLUSH_REG_SCAN_IN), .ZN(n12544) );
  NAND2_X1 U15869 ( .A1(n12545), .A2(n12544), .ZN(n15617) );
  NAND2_X1 U15870 ( .A1(n12546), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12547) );
  NAND2_X1 U15871 ( .A1(n12547), .A2(n16286), .ZN(n12565) );
  AND3_X1 U15872 ( .A1(n12549), .A2(n12548), .A3(n12565), .ZN(n16277) );
  NOR2_X1 U15873 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19710) );
  NAND3_X1 U15874 ( .A1(n15617), .A2(n16277), .A3(n19710), .ZN(n12550) );
  OAI21_X1 U15875 ( .B1(n15617), .B2(n16286), .A(n12550), .ZN(P2_U3595) );
  AND2_X1 U15876 ( .A1(n12554), .A2(n12553), .ZN(n12556) );
  OAI21_X1 U15877 ( .B1(n12557), .B2(n12556), .A(n12555), .ZN(n19841) );
  INV_X1 U15878 ( .A(n12559), .ZN(n12560) );
  OR2_X1 U15879 ( .A1(n16276), .A2(n12560), .ZN(n19842) );
  NOR2_X1 U15880 ( .A1(n19842), .A2(n19844), .ZN(n12561) );
  NAND2_X1 U15881 ( .A1(n19841), .A2(n12561), .ZN(n13321) );
  NOR2_X1 U15882 ( .A1(n16276), .A2(n12581), .ZN(n13327) );
  OAI21_X1 U15883 ( .B1(n12582), .B2(n12562), .A(n16271), .ZN(n12563) );
  INV_X1 U15884 ( .A(n12563), .ZN(n12566) );
  INV_X1 U15885 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12564) );
  OAI21_X1 U15886 ( .B1(n11963), .B2(n12565), .A(n12564), .ZN(n19830) );
  MUX2_X1 U15887 ( .A(n12566), .B(n19830), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n19848) );
  NAND2_X1 U15888 ( .A1(n13327), .A2(n19848), .ZN(n12567) );
  NAND2_X1 U15889 ( .A1(n13321), .A2(n12567), .ZN(n12568) );
  NAND2_X1 U15890 ( .A1(n12568), .A2(n19708), .ZN(n18776) );
  OR2_X1 U15891 ( .A1(n19812), .A2(n19710), .ZN(n19829) );
  NAND2_X1 U15892 ( .A1(n19829), .A2(n11587), .ZN(n12569) );
  AND2_X1 U15893 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19820) );
  INV_X1 U15894 ( .A(n12823), .ZN(n12571) );
  INV_X1 U15895 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n15620) );
  NAND2_X1 U15896 ( .A1(n15620), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12570) );
  NAND2_X1 U15897 ( .A1(n12571), .A2(n12570), .ZN(n12615) );
  OAI22_X1 U15898 ( .A1(n19129), .A2(n12904), .B1(n19736), .B2(n18921), .ZN(
        n12580) );
  OR2_X1 U15899 ( .A1(n12583), .A2(n14935), .ZN(n12614) );
  NAND2_X1 U15900 ( .A1(n12614), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12613) );
  INV_X1 U15901 ( .A(n12613), .ZN(n12572) );
  XOR2_X1 U15902 ( .A(n12583), .B(n12575), .Z(n12573) );
  NAND2_X1 U15903 ( .A1(n12572), .A2(n12573), .ZN(n12574) );
  XNOR2_X1 U15904 ( .A(n12573), .B(n12613), .ZN(n12598) );
  NAND2_X1 U15905 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n12598), .ZN(
        n12597) );
  NAND2_X1 U15906 ( .A1(n12574), .A2(n12597), .ZN(n13328) );
  XOR2_X1 U15907 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n13328), .Z(
        n12578) );
  OR2_X1 U15908 ( .A1(n14935), .A2(n12575), .ZN(n12576) );
  OR2_X1 U15909 ( .A1(n12583), .A2(n12576), .ZN(n13303) );
  XNOR2_X1 U15910 ( .A(n13302), .B(n13303), .ZN(n12577) );
  NAND2_X1 U15911 ( .A1(n12578), .A2(n12577), .ZN(n13330) );
  OAI21_X1 U15912 ( .B1(n12578), .B2(n12577), .A(n13330), .ZN(n19148) );
  NOR2_X1 U15913 ( .A1(n19148), .A2(n16194), .ZN(n12579) );
  AOI211_X1 U15914 ( .C1(n19118), .C2(n12903), .A(n12580), .B(n12579), .ZN(
        n12594) );
  MUX2_X1 U15915 ( .A(n12583), .B(n12582), .S(n12581), .Z(n12586) );
  INV_X1 U15916 ( .A(n12584), .ZN(n12585) );
  AOI21_X1 U15917 ( .B1(n12586), .B2(n13826), .A(n12585), .ZN(n13202) );
  NAND2_X1 U15918 ( .A1(n13202), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12612) );
  AND3_X1 U15919 ( .A1(n19177), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n12587) );
  OR2_X1 U15920 ( .A1(n12590), .A2(n12587), .ZN(n13127) );
  NOR2_X1 U15921 ( .A1(n12612), .A2(n13127), .ZN(n12588) );
  NAND2_X1 U15922 ( .A1(n12612), .A2(n13127), .ZN(n12601) );
  OAI21_X1 U15923 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12588), .A(
        n12601), .ZN(n12592) );
  OAI21_X1 U15924 ( .B1(n12590), .B2(n12589), .A(n13086), .ZN(n13308) );
  INV_X1 U15925 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13358) );
  XNOR2_X1 U15926 ( .A(n13308), .B(n13358), .ZN(n12591) );
  OR2_X1 U15927 ( .A1(n12592), .A2(n12591), .ZN(n19132) );
  OR2_X1 U15928 ( .A1(n18776), .A2(n11798), .ZN(n16192) );
  NAND2_X1 U15929 ( .A1(n12592), .A2(n12591), .ZN(n19130) );
  NAND3_X1 U15930 ( .A1(n19132), .A2(n19124), .A3(n19130), .ZN(n12593) );
  OAI211_X1 U15931 ( .C1(n13276), .C2(n16160), .A(n12594), .B(n12593), .ZN(
        P2_U3012) );
  XNOR2_X2 U15932 ( .A(n12595), .B(n12596), .ZN(n13267) );
  OAI21_X1 U15933 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12598), .A(
        n12597), .ZN(n19158) );
  OR2_X1 U15934 ( .A1(n18921), .A2(n19734), .ZN(n19164) );
  OAI21_X1 U15935 ( .B1(n19129), .B2(n13130), .A(n19164), .ZN(n12599) );
  INV_X1 U15936 ( .A(n12599), .ZN(n12600) );
  OAI21_X1 U15937 ( .B1(n19158), .B2(n16194), .A(n12600), .ZN(n12604) );
  OAI21_X1 U15938 ( .B1(n12612), .B2(n13127), .A(n12601), .ZN(n12602) );
  XNOR2_X1 U15939 ( .A(n12602), .B(n19150), .ZN(n19167) );
  NOR2_X1 U15940 ( .A1(n19167), .A2(n16192), .ZN(n12603) );
  AOI211_X1 U15941 ( .C1(n19118), .C2(n13130), .A(n12604), .B(n12603), .ZN(
        n12605) );
  OAI21_X1 U15942 ( .B1(n13267), .B2(n16160), .A(n12605), .ZN(P2_U3013) );
  INV_X1 U15943 ( .A(n12606), .ZN(n12609) );
  INV_X1 U15944 ( .A(n12607), .ZN(n12608) );
  NAND2_X1 U15945 ( .A1(n12609), .A2(n12608), .ZN(n12611) );
  INV_X1 U15946 ( .A(n13252), .ZN(n16249) );
  OAI21_X1 U15947 ( .B1(n13202), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12612), .ZN(n16247) );
  INV_X1 U15948 ( .A(n16247), .ZN(n12618) );
  OAI21_X1 U15949 ( .B1(n12614), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12613), .ZN(n16255) );
  INV_X1 U15950 ( .A(n19129), .ZN(n16184) );
  OAI21_X1 U15951 ( .B1(n16184), .B2(n12615), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12616) );
  INV_X2 U15952 ( .A(n18921), .ZN(n19119) );
  NAND2_X1 U15953 ( .A1(n19119), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n16253) );
  OAI211_X1 U15954 ( .C1(n16194), .C2(n16255), .A(n12616), .B(n16253), .ZN(
        n12617) );
  AOI21_X1 U15955 ( .B1(n19124), .B2(n12618), .A(n12617), .ZN(n12619) );
  OAI21_X1 U15956 ( .B1(n16249), .B2(n16160), .A(n12619), .ZN(P2_U3014) );
  OAI21_X1 U15957 ( .B1(n12621), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n20757), 
        .ZN(n12622) );
  OAI21_X1 U15958 ( .B1(n12623), .B2(n20757), .A(n12622), .ZN(P1_U3487) );
  OR2_X1 U15959 ( .A1(n12800), .A2(n12624), .ZN(n12629) );
  INV_X1 U15960 ( .A(n12625), .ZN(n12627) );
  NAND2_X1 U15961 ( .A1(n12627), .A2(n12626), .ZN(n12628) );
  NAND2_X1 U15962 ( .A1(n12629), .A2(n12628), .ZN(n19879) );
  NAND3_X1 U15963 ( .A1(n10261), .A2(n15849), .A3(n12817), .ZN(n12630) );
  AND2_X1 U15964 ( .A1(n12630), .A2(n20659), .ZN(n20761) );
  OR2_X1 U15965 ( .A1(n19879), .A2(n20761), .ZN(n15820) );
  AND2_X1 U15966 ( .A1(n15820), .A2(n12763), .ZN(n19886) );
  INV_X1 U15967 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n12648) );
  NAND2_X1 U15968 ( .A1(n12632), .A2(n12631), .ZN(n15816) );
  NAND4_X1 U15969 ( .A1(n12636), .A2(n12635), .A3(n12634), .A4(n12633), .ZN(
        n12637) );
  AND3_X1 U15970 ( .A1(n12949), .A2(n15816), .A3(n12637), .ZN(n12644) );
  NAND2_X1 U15971 ( .A1(n12800), .A2(n12638), .ZN(n12643) );
  INV_X1 U15972 ( .A(n12639), .ZN(n12641) );
  NAND2_X1 U15973 ( .A1(n12641), .A2(n12640), .ZN(n12642) );
  OAI211_X1 U15974 ( .C1(n12800), .C2(n12644), .A(n12643), .B(n12642), .ZN(
        n12645) );
  NAND2_X1 U15975 ( .A1(n12645), .A2(n20105), .ZN(n15817) );
  INV_X1 U15976 ( .A(n15817), .ZN(n12646) );
  NAND2_X1 U15977 ( .A1(n19886), .A2(n12646), .ZN(n12647) );
  OAI21_X1 U15978 ( .B1(n19886), .B2(n12648), .A(n12647), .ZN(P1_U3484) );
  INV_X1 U15979 ( .A(n12649), .ZN(n12681) );
  NAND2_X1 U15980 ( .A1(n12681), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n12651) );
  OAI211_X1 U15981 ( .C1(n19051), .C2(n19063), .A(n12651), .B(n12650), .ZN(
        P2_U2963) );
  INV_X1 U15982 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19098) );
  NAND2_X1 U15983 ( .A1(n12681), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n12652) );
  MUX2_X1 U15984 ( .A(BUF1_REG_8__SCAN_IN), .B(BUF2_REG_8__SCAN_IN), .S(n15061), .Z(n19009) );
  NAND2_X1 U15985 ( .A1(n12674), .A2(n19009), .ZN(n12660) );
  OAI211_X1 U15986 ( .C1(n19098), .C2(n19051), .A(n12652), .B(n12660), .ZN(
        P2_U2975) );
  INV_X1 U15987 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n19065) );
  NAND2_X1 U15988 ( .A1(n12681), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12655) );
  NAND2_X1 U15989 ( .A1(n15061), .A2(BUF2_REG_10__SCAN_IN), .ZN(n12654) );
  INV_X1 U15990 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16393) );
  OR2_X1 U15991 ( .A1(n15061), .A2(n16393), .ZN(n12653) );
  NAND2_X1 U15992 ( .A1(n12654), .A2(n12653), .ZN(n19002) );
  NAND2_X1 U15993 ( .A1(n12674), .A2(n19002), .ZN(n12662) );
  OAI211_X1 U15994 ( .C1(n19065), .C2(n19051), .A(n12655), .B(n12662), .ZN(
        P2_U2962) );
  INV_X1 U15995 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n19059) );
  NAND2_X1 U15996 ( .A1(n12681), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n12657) );
  OAI211_X1 U15997 ( .C1(n19051), .C2(n19059), .A(n12657), .B(n12656), .ZN(
        P2_U2965) );
  NAND2_X1 U15998 ( .A1(n12681), .A2(P2_UWORD_REG_4__SCAN_IN), .ZN(n12658) );
  OAI22_X1 U15999 ( .A1(n15061), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n15064), .ZN(n19032) );
  INV_X1 U16000 ( .A(n19032), .ZN(n16147) );
  NAND2_X1 U16001 ( .A1(n12674), .A2(n16147), .ZN(n12678) );
  OAI211_X1 U16002 ( .C1(n19051), .C2(n12659), .A(n12658), .B(n12678), .ZN(
        P2_U2956) );
  NAND2_X1 U16003 ( .A1(n12681), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n12661) );
  OAI211_X1 U16004 ( .C1(n15101), .C2(n19051), .A(n12661), .B(n12660), .ZN(
        P2_U2960) );
  INV_X1 U16005 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19094) );
  NAND2_X1 U16006 ( .A1(n12681), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n12663) );
  OAI211_X1 U16007 ( .C1(n19094), .C2(n19051), .A(n12663), .B(n12662), .ZN(
        P2_U2977) );
  NAND2_X1 U16008 ( .A1(n12681), .A2(P2_UWORD_REG_7__SCAN_IN), .ZN(n12665) );
  OAI211_X1 U16009 ( .C1(n19051), .C2(n19070), .A(n12665), .B(n12664), .ZN(
        P2_U2959) );
  INV_X1 U16010 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n12668) );
  NAND2_X1 U16011 ( .A1(n12681), .A2(P2_UWORD_REG_6__SCAN_IN), .ZN(n12667) );
  OAI211_X1 U16012 ( .C1(n19051), .C2(n12668), .A(n12667), .B(n12666), .ZN(
        P2_U2958) );
  INV_X1 U16013 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n19067) );
  NAND2_X1 U16014 ( .A1(n12681), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n12670) );
  OAI211_X1 U16015 ( .C1(n19051), .C2(n19067), .A(n12670), .B(n12669), .ZN(
        P2_U2961) );
  INV_X1 U16016 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19087) );
  NAND2_X1 U16017 ( .A1(n12681), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n12675) );
  NAND2_X1 U16018 ( .A1(n15061), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12673) );
  INV_X1 U16019 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n12671) );
  OR2_X1 U16020 ( .A1(n15061), .A2(n12671), .ZN(n12672) );
  NAND2_X1 U16021 ( .A1(n12673), .A2(n12672), .ZN(n18993) );
  NAND2_X1 U16022 ( .A1(n12674), .A2(n18993), .ZN(n12682) );
  OAI211_X1 U16023 ( .C1(n19087), .C2(n19051), .A(n12675), .B(n12682), .ZN(
        P2_U2981) );
  NAND2_X1 U16024 ( .A1(n12681), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n12677) );
  OAI211_X1 U16025 ( .C1(n19051), .C2(n19061), .A(n12677), .B(n12676), .ZN(
        P2_U2964) );
  INV_X1 U16026 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n12680) );
  NAND2_X1 U16027 ( .A1(n12681), .A2(P2_LWORD_REG_4__SCAN_IN), .ZN(n12679) );
  OAI211_X1 U16028 ( .C1(n12680), .C2(n19051), .A(n12679), .B(n12678), .ZN(
        P2_U2971) );
  INV_X1 U16029 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n19057) );
  NAND2_X1 U16030 ( .A1(n12681), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n12683) );
  OAI211_X1 U16031 ( .C1(n19057), .C2(n19051), .A(n12683), .B(n12682), .ZN(
        P2_U2966) );
  AND2_X1 U16032 ( .A1(n12685), .A2(n12684), .ZN(n12686) );
  AND2_X1 U16033 ( .A1(n12772), .A2(n19177), .ZN(n12689) );
  NAND2_X1 U16034 ( .A1(n19014), .A2(n12689), .ZN(n15127) );
  INV_X1 U16035 ( .A(n12690), .ZN(n12691) );
  NAND2_X1 U16036 ( .A1(n19014), .A2(n12691), .ZN(n15065) );
  NAND2_X1 U16037 ( .A1(n15127), .A2(n15065), .ZN(n19008) );
  INV_X1 U16038 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19416) );
  OAI21_X1 U16039 ( .B1(n19181), .B2(n11587), .A(n19416), .ZN(n12827) );
  AOI22_X1 U16040 ( .A1(n12827), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19812), .B2(n19839), .ZN(n12692) );
  NAND2_X1 U16041 ( .A1(n19865), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12694) );
  AND4_X1 U16042 ( .A1(n19181), .A2(n12694), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n19416), .ZN(n12695) );
  NOR2_X1 U16043 ( .A1(n12697), .A2(n12696), .ZN(n12698) );
  NOR2_X1 U16044 ( .A1(n12699), .A2(n12698), .ZN(n16245) );
  NAND2_X1 U16045 ( .A1(n13421), .A2(n16245), .ZN(n19042) );
  NAND2_X1 U16046 ( .A1(n19014), .A2(n12700), .ZN(n18984) );
  OAI211_X1 U16047 ( .C1(n13421), .C2(n16245), .A(n19042), .B(n19044), .ZN(
        n12702) );
  AND2_X1 U16048 ( .A1(n19014), .A2(n11773), .ZN(n19040) );
  AOI22_X1 U16049 ( .A1(n19040), .A2(n16245), .B1(n19039), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n12701) );
  OAI211_X1 U16050 ( .C1(n19048), .C2(n13238), .A(n12702), .B(n12701), .ZN(
        P2_U2919) );
  NAND2_X1 U16051 ( .A1(n12896), .A2(n12946), .ZN(n12845) );
  INV_X1 U16052 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20007) );
  INV_X2 U16053 ( .A(n12896), .ZN(n12890) );
  NAND2_X1 U16054 ( .A1(n12890), .A2(P1_LWORD_REG_1__SCAN_IN), .ZN(n12707) );
  NOR2_X2 U16055 ( .A1(n12704), .A2(n12703), .ZN(n12893) );
  NAND2_X1 U16056 ( .A1(n13389), .A2(DATAI_1_), .ZN(n12706) );
  NAND2_X1 U16057 ( .A1(n13387), .A2(BUF1_REG_1__SCAN_IN), .ZN(n12705) );
  AND2_X1 U16058 ( .A1(n12706), .A2(n12705), .ZN(n20082) );
  INV_X1 U16059 ( .A(n20082), .ZN(n14335) );
  NAND2_X1 U16060 ( .A1(n12893), .A2(n14335), .ZN(n12717) );
  OAI211_X1 U16061 ( .C1(n12845), .C2(n20007), .A(n12707), .B(n12717), .ZN(
        P1_U2953) );
  INV_X1 U16062 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20005) );
  NAND2_X1 U16063 ( .A1(n12890), .A2(P1_LWORD_REG_2__SCAN_IN), .ZN(n12710) );
  NAND2_X1 U16064 ( .A1(n13389), .A2(DATAI_2_), .ZN(n12709) );
  NAND2_X1 U16065 ( .A1(n13387), .A2(BUF1_REG_2__SCAN_IN), .ZN(n12708) );
  AND2_X1 U16066 ( .A1(n12709), .A2(n12708), .ZN(n13395) );
  INV_X1 U16067 ( .A(n13395), .ZN(n14330) );
  NAND2_X1 U16068 ( .A1(n12893), .A2(n14330), .ZN(n12725) );
  OAI211_X1 U16069 ( .C1(n12845), .C2(n20005), .A(n12710), .B(n12725), .ZN(
        P1_U2954) );
  INV_X1 U16070 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13017) );
  NAND2_X1 U16071 ( .A1(n12890), .A2(P1_UWORD_REG_3__SCAN_IN), .ZN(n12713) );
  NAND2_X1 U16072 ( .A1(n13389), .A2(DATAI_3_), .ZN(n12712) );
  NAND2_X1 U16073 ( .A1(n13387), .A2(BUF1_REG_3__SCAN_IN), .ZN(n12711) );
  AND2_X1 U16074 ( .A1(n12712), .A2(n12711), .ZN(n20088) );
  INV_X1 U16075 ( .A(n20088), .ZN(n14325) );
  NAND2_X1 U16076 ( .A1(n12893), .A2(n14325), .ZN(n12874) );
  OAI211_X1 U16077 ( .C1(n12845), .C2(n13017), .A(n12713), .B(n12874), .ZN(
        P1_U2940) );
  INV_X1 U16078 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13019) );
  NAND2_X1 U16079 ( .A1(n12890), .A2(P1_UWORD_REG_4__SCAN_IN), .ZN(n12716) );
  INV_X1 U16080 ( .A(DATAI_4_), .ZN(n12715) );
  NAND2_X1 U16081 ( .A1(n13387), .A2(BUF1_REG_4__SCAN_IN), .ZN(n12714) );
  OAI21_X1 U16082 ( .B1(n13387), .B2(n12715), .A(n12714), .ZN(n14320) );
  NAND2_X1 U16083 ( .A1(n12893), .A2(n14320), .ZN(n12877) );
  OAI211_X1 U16084 ( .C1(n12845), .C2(n13019), .A(n12716), .B(n12877), .ZN(
        P1_U2941) );
  INV_X1 U16085 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n12749) );
  NAND2_X1 U16086 ( .A1(n12890), .A2(P1_UWORD_REG_1__SCAN_IN), .ZN(n12718) );
  OAI211_X1 U16087 ( .C1(n12845), .C2(n12749), .A(n12718), .B(n12717), .ZN(
        P1_U2938) );
  INV_X1 U16088 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13025) );
  NAND2_X1 U16089 ( .A1(n12890), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n12721) );
  INV_X1 U16090 ( .A(DATAI_13_), .ZN(n12720) );
  NAND2_X1 U16091 ( .A1(n13387), .A2(BUF1_REG_13__SCAN_IN), .ZN(n12719) );
  OAI21_X1 U16092 ( .B1(n13387), .B2(n12720), .A(n12719), .ZN(n14269) );
  NAND2_X1 U16093 ( .A1(n12893), .A2(n14269), .ZN(n12865) );
  OAI211_X1 U16094 ( .C1(n12845), .C2(n13025), .A(n12721), .B(n12865), .ZN(
        P1_U2950) );
  INV_X1 U16095 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13027) );
  NAND2_X1 U16096 ( .A1(n12890), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n12724) );
  INV_X1 U16097 ( .A(DATAI_14_), .ZN(n12723) );
  NAND2_X1 U16098 ( .A1(n13387), .A2(BUF1_REG_14__SCAN_IN), .ZN(n12722) );
  OAI21_X1 U16099 ( .B1(n13387), .B2(n12723), .A(n12722), .ZN(n14264) );
  NAND2_X1 U16100 ( .A1(n12893), .A2(n14264), .ZN(n12861) );
  OAI211_X1 U16101 ( .C1(n12845), .C2(n13027), .A(n12724), .B(n12861), .ZN(
        P1_U2951) );
  INV_X1 U16102 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13029) );
  NAND2_X1 U16103 ( .A1(n12890), .A2(P1_UWORD_REG_2__SCAN_IN), .ZN(n12726) );
  OAI211_X1 U16104 ( .C1(n12845), .C2(n13029), .A(n12726), .B(n12725), .ZN(
        P1_U2939) );
  INV_X1 U16105 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n12752) );
  NAND2_X1 U16106 ( .A1(n12890), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n12729) );
  INV_X1 U16107 ( .A(DATAI_9_), .ZN(n12728) );
  NAND2_X1 U16108 ( .A1(n13387), .A2(BUF1_REG_9__SCAN_IN), .ZN(n12727) );
  OAI21_X1 U16109 ( .B1(n13387), .B2(n12728), .A(n12727), .ZN(n14293) );
  NAND2_X1 U16110 ( .A1(n12893), .A2(n14293), .ZN(n12887) );
  OAI211_X1 U16111 ( .C1(n12845), .C2(n12752), .A(n12729), .B(n12887), .ZN(
        P1_U2946) );
  INV_X1 U16112 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20012) );
  NAND2_X1 U16113 ( .A1(n12890), .A2(P1_LWORD_REG_0__SCAN_IN), .ZN(n12732) );
  NAND2_X1 U16114 ( .A1(n13389), .A2(DATAI_0_), .ZN(n12731) );
  NAND2_X1 U16115 ( .A1(n13387), .A2(BUF1_REG_0__SCAN_IN), .ZN(n12730) );
  AND2_X1 U16116 ( .A1(n12731), .A2(n12730), .ZN(n20076) );
  INV_X1 U16117 ( .A(n20076), .ZN(n14343) );
  NAND2_X1 U16118 ( .A1(n12893), .A2(n14343), .ZN(n12872) );
  OAI211_X1 U16119 ( .C1(n12845), .C2(n20012), .A(n12732), .B(n12872), .ZN(
        P1_U2952) );
  INV_X1 U16120 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13032) );
  NAND2_X1 U16121 ( .A1(n13389), .A2(DATAI_5_), .ZN(n12734) );
  NAND2_X1 U16122 ( .A1(n13387), .A2(BUF1_REG_5__SCAN_IN), .ZN(n12733) );
  AND2_X1 U16123 ( .A1(n12734), .A2(n12733), .ZN(n20094) );
  INV_X1 U16124 ( .A(n20094), .ZN(n14314) );
  NAND2_X1 U16125 ( .A1(n12893), .A2(n14314), .ZN(n12878) );
  NAND2_X1 U16126 ( .A1(n12890), .A2(P1_UWORD_REG_5__SCAN_IN), .ZN(n12735) );
  OAI211_X1 U16127 ( .C1(n12845), .C2(n13032), .A(n12878), .B(n12735), .ZN(
        P1_U2942) );
  OR2_X1 U16128 ( .A1(n12737), .A2(n12736), .ZN(n12738) );
  NAND2_X1 U16129 ( .A1(n12840), .A2(n12738), .ZN(n19970) );
  INV_X1 U16130 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19960) );
  NAND2_X1 U16131 ( .A1(n10704), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n14622) );
  OAI21_X1 U16132 ( .B1(n20024), .B2(n19960), .A(n14622), .ZN(n12739) );
  AOI21_X1 U16133 ( .B1(n15976), .B2(n19960), .A(n12739), .ZN(n12743) );
  OR2_X1 U16134 ( .A1(n12740), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14621) );
  NAND3_X1 U16135 ( .A1(n14621), .A2(n12741), .A3(n20019), .ZN(n12742) );
  OAI211_X1 U16136 ( .C1(n19970), .C2(n15947), .A(n12743), .B(n12742), .ZN(
        P1_U2998) );
  INV_X1 U16137 ( .A(n12744), .ZN(n15828) );
  INV_X1 U16138 ( .A(n15849), .ZN(n12745) );
  OAI211_X1 U16139 ( .C1(n12962), .C2(n15828), .A(n12745), .B(n12763), .ZN(
        n12746) );
  INV_X1 U16140 ( .A(n12746), .ZN(n12747) );
  NAND2_X1 U16141 ( .A1(n19979), .A2(n20074), .ZN(n13031) );
  NOR2_X1 U16142 ( .A1(n20652), .A2(n20648), .ZN(n16122) );
  NAND2_X1 U16143 ( .A1(n20649), .A2(n16122), .ZN(n20758) );
  INV_X2 U16144 ( .A(n20758), .ZN(n20009) );
  AOI22_X1 U16145 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n19999), .B1(n20009), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n12748) );
  OAI21_X1 U16146 ( .B1(n12749), .B2(n13031), .A(n12748), .ZN(P1_U2919) );
  INV_X1 U16147 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n12871) );
  AOI22_X1 U16148 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n19999), .B1(n20009), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n12750) );
  OAI21_X1 U16149 ( .B1(n12871), .B2(n13031), .A(n12750), .ZN(P1_U2914) );
  AOI22_X1 U16150 ( .A1(n20009), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n19999), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n12751) );
  OAI21_X1 U16151 ( .B1(n12752), .B2(n13031), .A(n12751), .ZN(P1_U2911) );
  INV_X1 U16152 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n12849) );
  AOI22_X1 U16153 ( .A1(n20009), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n19999), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12753) );
  OAI21_X1 U16154 ( .B1(n12849), .B2(n13031), .A(n12753), .ZN(P1_U2909) );
  INV_X1 U16155 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n12853) );
  AOI22_X1 U16156 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20009), .B1(n19999), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12754) );
  OAI21_X1 U16157 ( .B1(n12853), .B2(n13031), .A(n12754), .ZN(P1_U2908) );
  OAI21_X1 U16158 ( .B1(n12757), .B2(n12756), .A(n12755), .ZN(n13443) );
  INV_X1 U16159 ( .A(n12758), .ZN(n12761) );
  NOR2_X1 U16160 ( .A1(n12759), .A2(n12817), .ZN(n12760) );
  NAND2_X1 U16161 ( .A1(n12761), .A2(n12760), .ZN(n12762) );
  NOR2_X1 U16162 ( .A1(n12766), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12767) );
  OR2_X1 U16163 ( .A1(n12768), .A2(n12767), .ZN(n13463) );
  OAI222_X1 U16164 ( .A1(n13443), .A2(n14254), .B1(n12769), .B2(n14260), .C1(
        n13463), .C2(n14259), .ZN(P1_U2872) );
  INV_X1 U16165 ( .A(n13352), .ZN(n15590) );
  NAND2_X1 U16166 ( .A1(n12770), .A2(n15590), .ZN(n12771) );
  NAND2_X1 U16167 ( .A1(n14743), .A2(n12772), .ZN(n15060) );
  MUX2_X1 U16168 ( .A(n16249), .B(n13199), .S(n15055), .Z(n12773) );
  OAI21_X1 U16169 ( .B1(n19834), .B2(n15060), .A(n12773), .ZN(P2_U2887) );
  NAND2_X1 U16170 ( .A1(n12827), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12774) );
  NAND2_X1 U16171 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19839), .ZN(
        n19479) );
  NAND2_X1 U16172 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19828), .ZN(
        n19447) );
  NAND2_X1 U16173 ( .A1(n19479), .A2(n19447), .ZN(n13423) );
  NAND2_X1 U16174 ( .A1(n19812), .A2(n13423), .ZN(n19481) );
  NAND2_X1 U16175 ( .A1(n12774), .A2(n19481), .ZN(n12775) );
  INV_X1 U16176 ( .A(n12785), .ZN(n12777) );
  NAND2_X1 U16177 ( .A1(n12776), .A2(n19181), .ZN(n14885) );
  INV_X1 U16178 ( .A(n14885), .ZN(n14916) );
  NAND2_X1 U16179 ( .A1(n14916), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12787) );
  MUX2_X1 U16180 ( .A(n13267), .B(n11783), .S(n15055), .Z(n12778) );
  OAI21_X1 U16181 ( .B1(n19814), .B2(n15060), .A(n12778), .ZN(P2_U2886) );
  NAND2_X1 U16182 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19510) );
  NAND2_X1 U16183 ( .A1(n19510), .A2(n19819), .ZN(n12780) );
  NAND2_X1 U16184 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19641) );
  INV_X1 U16185 ( .A(n19641), .ZN(n12779) );
  AND2_X1 U16186 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12779), .ZN(
        n12824) );
  INV_X1 U16187 ( .A(n12824), .ZN(n12825) );
  AND2_X1 U16188 ( .A1(n12780), .A2(n12825), .ZN(n13226) );
  AOI22_X1 U16189 ( .A1(n12827), .A2(n16257), .B1(n19812), .B2(n13226), .ZN(
        n12781) );
  INV_X1 U16190 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15639) );
  NOR2_X1 U16191 ( .A1(n14885), .A2(n15639), .ZN(n12783) );
  NAND2_X1 U16192 ( .A1(n12786), .A2(n12785), .ZN(n12790) );
  INV_X1 U16193 ( .A(n12787), .ZN(n12788) );
  MUX2_X1 U16194 ( .A(n13276), .B(n11829), .S(n15055), .Z(n12791) );
  OAI21_X1 U16195 ( .B1(n19813), .B2(n15060), .A(n12791), .ZN(P2_U2885) );
  INV_X1 U16196 ( .A(n20181), .ZN(n20735) );
  NAND3_X1 U16197 ( .A1(n12792), .A2(n12948), .A3(n11561), .ZN(n14640) );
  INV_X1 U16198 ( .A(n14640), .ZN(n12793) );
  OAI22_X1 U16199 ( .A1(n20735), .A2(n12793), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14637), .ZN(n15804) );
  OAI22_X1 U16200 ( .A1(n20648), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14657), .ZN(n12794) );
  AOI21_X1 U16201 ( .B1(n15804), .B2(n19877), .A(n12794), .ZN(n12807) );
  OAI211_X1 U16202 ( .C1(n13456), .C2(n13396), .A(n12796), .B(n12795), .ZN(
        n12797) );
  INV_X1 U16203 ( .A(n12797), .ZN(n12802) );
  INV_X1 U16204 ( .A(n12962), .ZN(n14636) );
  AOI21_X1 U16205 ( .B1(n14636), .B2(n14262), .A(n12798), .ZN(n12799) );
  NAND2_X1 U16206 ( .A1(n12800), .A2(n12799), .ZN(n12801) );
  NAND4_X1 U16207 ( .A1(n12804), .A2(n12803), .A3(n12802), .A4(n12801), .ZN(
        n12976) );
  INV_X1 U16208 ( .A(n12976), .ZN(n15806) );
  NAND2_X1 U16209 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16122), .ZN(n16127) );
  INV_X1 U16210 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19885) );
  OAI22_X1 U16211 ( .A1(n15806), .A2(n19878), .B1(n16127), .B2(n19885), .ZN(
        n16112) );
  AOI21_X1 U16212 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20649), .A(n16112), 
        .ZN(n14647) );
  NOR2_X1 U16213 ( .A1(n14636), .A2(n12805), .ZN(n15803) );
  AOI22_X1 U16214 ( .A1(n15803), .A2(n19877), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14647), .ZN(n12806) );
  OAI21_X1 U16215 ( .B1(n12807), .B2(n14647), .A(n12806), .ZN(P1_U3474) );
  INV_X1 U16216 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n20750) );
  OAI21_X1 U16217 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n12809), .A(
        n12808), .ZN(n20031) );
  OAI22_X1 U16218 ( .A1(n20036), .A2(n20750), .B1(n16106), .B2(n20031), .ZN(
        n12816) );
  INV_X1 U16219 ( .A(n20056), .ZN(n16046) );
  INV_X1 U16220 ( .A(n12810), .ZN(n12811) );
  OAI21_X1 U16221 ( .B1(n16046), .B2(n12811), .A(n20055), .ZN(n14623) );
  INV_X1 U16222 ( .A(n14624), .ZN(n12813) );
  INV_X1 U16223 ( .A(n12812), .ZN(n14628) );
  OAI21_X1 U16224 ( .B1(n12813), .B2(n14628), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12814) );
  OAI211_X1 U16225 ( .C1(n20038), .C2(n13463), .A(n14623), .B(n12814), .ZN(
        n12815) );
  OR2_X1 U16226 ( .A1(n12816), .A2(n12815), .ZN(P1_U3031) );
  XNOR2_X1 U16227 ( .A(n19975), .B(n12817), .ZN(n14627) );
  AOI22_X1 U16228 ( .A1(n14223), .A2(n14627), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n14222), .ZN(n12818) );
  OAI21_X1 U16229 ( .B1(n19970), .B2(n14254), .A(n12818), .ZN(P1_U2871) );
  NAND2_X1 U16230 ( .A1(n15615), .A2(n12823), .ZN(n12829) );
  NAND2_X1 U16231 ( .A1(n12824), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19648) );
  NAND2_X1 U16232 ( .A1(n19811), .A2(n12825), .ZN(n12826) );
  AND3_X1 U16233 ( .A1(n19648), .A2(n19812), .A3(n12826), .ZN(n13234) );
  AOI21_X1 U16234 ( .B1(n12827), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n13234), .ZN(n12828) );
  NAND2_X1 U16235 ( .A1(n12829), .A2(n12828), .ZN(n12831) );
  NOR2_X1 U16236 ( .A1(n14885), .A2(n19176), .ZN(n12830) );
  NAND2_X1 U16237 ( .A1(n12831), .A2(n12830), .ZN(n13004) );
  OR2_X1 U16238 ( .A1(n12831), .A2(n12830), .ZN(n12832) );
  NAND2_X1 U16239 ( .A1(n12833), .A2(n9669), .ZN(n12835) );
  MUX2_X1 U16240 ( .A(n13249), .B(n12838), .S(n15055), .Z(n12839) );
  OAI21_X1 U16241 ( .B1(n19445), .B2(n15060), .A(n12839), .ZN(P2_U2884) );
  OAI21_X1 U16242 ( .B1(n10096), .B2(n11077), .A(n12841), .ZN(n14200) );
  OAI21_X1 U16243 ( .B1(n12843), .B2(n12842), .A(n13101), .ZN(n14193) );
  INV_X1 U16244 ( .A(n14193), .ZN(n20060) );
  AOI22_X1 U16245 ( .A1(n14223), .A2(n20060), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n14222), .ZN(n12844) );
  OAI21_X1 U16246 ( .B1(n14200), .B2(n14254), .A(n12844), .ZN(P1_U2870) );
  NAND2_X1 U16247 ( .A1(n12890), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n12848) );
  INV_X1 U16248 ( .A(DATAI_11_), .ZN(n12847) );
  NAND2_X1 U16249 ( .A1(n13387), .A2(BUF1_REG_11__SCAN_IN), .ZN(n12846) );
  OAI21_X1 U16250 ( .B1(n13387), .B2(n12847), .A(n12846), .ZN(n14280) );
  NAND2_X1 U16251 ( .A1(n12893), .A2(n14280), .ZN(n12892) );
  OAI211_X1 U16252 ( .C1(n12898), .C2(n12849), .A(n12848), .B(n12892), .ZN(
        P1_U2948) );
  NAND2_X1 U16253 ( .A1(n12890), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n12852) );
  INV_X1 U16254 ( .A(DATAI_12_), .ZN(n12851) );
  NAND2_X1 U16255 ( .A1(n13387), .A2(BUF1_REG_12__SCAN_IN), .ZN(n12850) );
  OAI21_X1 U16256 ( .B1(n13387), .B2(n12851), .A(n12850), .ZN(n14275) );
  NAND2_X1 U16257 ( .A1(n12893), .A2(n14275), .ZN(n12863) );
  OAI211_X1 U16258 ( .C1(n12898), .C2(n12853), .A(n12852), .B(n12863), .ZN(
        P1_U2949) );
  INV_X1 U16259 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13023) );
  NAND2_X1 U16260 ( .A1(n12890), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n12856) );
  INV_X1 U16261 ( .A(DATAI_10_), .ZN(n12855) );
  NAND2_X1 U16262 ( .A1(n13387), .A2(BUF1_REG_10__SCAN_IN), .ZN(n12854) );
  OAI21_X1 U16263 ( .B1(n13387), .B2(n12855), .A(n12854), .ZN(n14288) );
  NAND2_X1 U16264 ( .A1(n12893), .A2(n14288), .ZN(n12889) );
  OAI211_X1 U16265 ( .C1(n12898), .C2(n13023), .A(n12856), .B(n12889), .ZN(
        P1_U2947) );
  INV_X1 U16266 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13015) );
  NAND2_X1 U16267 ( .A1(n12890), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n12859) );
  INV_X1 U16268 ( .A(DATAI_8_), .ZN(n12858) );
  NAND2_X1 U16269 ( .A1(n13387), .A2(BUF1_REG_8__SCAN_IN), .ZN(n12857) );
  OAI21_X1 U16270 ( .B1(n13387), .B2(n12858), .A(n12857), .ZN(n14299) );
  NAND2_X1 U16271 ( .A1(n12893), .A2(n14299), .ZN(n12885) );
  OAI211_X1 U16272 ( .C1(n12898), .C2(n13015), .A(n12859), .B(n12885), .ZN(
        P1_U2945) );
  INV_X1 U16273 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n19981) );
  NAND2_X1 U16274 ( .A1(n12890), .A2(P1_LWORD_REG_14__SCAN_IN), .ZN(n12860) );
  OAI211_X1 U16275 ( .C1(n12898), .C2(n19981), .A(n12861), .B(n12860), .ZN(
        P1_U2966) );
  INV_X1 U16276 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n19985) );
  NAND2_X1 U16277 ( .A1(n12890), .A2(P1_LWORD_REG_12__SCAN_IN), .ZN(n12862) );
  OAI211_X1 U16278 ( .C1(n12898), .C2(n19985), .A(n12863), .B(n12862), .ZN(
        P1_U2964) );
  INV_X1 U16279 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n19983) );
  NAND2_X1 U16280 ( .A1(n12890), .A2(P1_LWORD_REG_13__SCAN_IN), .ZN(n12864) );
  OAI211_X1 U16281 ( .C1(n12898), .C2(n19983), .A(n12865), .B(n12864), .ZN(
        P1_U2965) );
  INV_X1 U16282 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13013) );
  NAND2_X1 U16283 ( .A1(n12890), .A2(P1_UWORD_REG_7__SCAN_IN), .ZN(n12868) );
  NAND2_X1 U16284 ( .A1(n13389), .A2(DATAI_7_), .ZN(n12867) );
  NAND2_X1 U16285 ( .A1(n13387), .A2(BUF1_REG_7__SCAN_IN), .ZN(n12866) );
  AND2_X1 U16286 ( .A1(n12867), .A2(n12866), .ZN(n20108) );
  INV_X1 U16287 ( .A(n20108), .ZN(n14304) );
  NAND2_X1 U16288 ( .A1(n12893), .A2(n14304), .ZN(n12882) );
  OAI211_X1 U16289 ( .C1(n12898), .C2(n13013), .A(n12868), .B(n12882), .ZN(
        P1_U2944) );
  NAND2_X1 U16290 ( .A1(n12890), .A2(P1_UWORD_REG_6__SCAN_IN), .ZN(n12870) );
  INV_X1 U16291 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16401) );
  NAND2_X1 U16292 ( .A1(n13387), .A2(n16401), .ZN(n12869) );
  OAI21_X1 U16293 ( .B1(n13387), .B2(DATAI_6_), .A(n12869), .ZN(n20100) );
  INV_X1 U16294 ( .A(n20100), .ZN(n14309) );
  NAND2_X1 U16295 ( .A1(n12893), .A2(n14309), .ZN(n12880) );
  OAI211_X1 U16296 ( .C1(n12898), .C2(n12871), .A(n12870), .B(n12880), .ZN(
        P1_U2943) );
  INV_X1 U16297 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13021) );
  NAND2_X1 U16298 ( .A1(n12890), .A2(P1_UWORD_REG_0__SCAN_IN), .ZN(n12873) );
  OAI211_X1 U16299 ( .C1(n12898), .C2(n13021), .A(n12873), .B(n12872), .ZN(
        P1_U2937) );
  INV_X1 U16300 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20003) );
  NAND2_X1 U16301 ( .A1(n12890), .A2(P1_LWORD_REG_3__SCAN_IN), .ZN(n12875) );
  OAI211_X1 U16302 ( .C1(n12898), .C2(n20003), .A(n12875), .B(n12874), .ZN(
        P1_U2955) );
  INV_X1 U16303 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20001) );
  NAND2_X1 U16304 ( .A1(n12890), .A2(P1_LWORD_REG_4__SCAN_IN), .ZN(n12876) );
  OAI211_X1 U16305 ( .C1(n12898), .C2(n20001), .A(n12877), .B(n12876), .ZN(
        P1_U2956) );
  NAND2_X1 U16306 ( .A1(n12890), .A2(P1_LWORD_REG_5__SCAN_IN), .ZN(n12879) );
  OAI211_X1 U16307 ( .C1(n12898), .C2(n11111), .A(n12879), .B(n12878), .ZN(
        P1_U2957) );
  INV_X1 U16308 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n19997) );
  NAND2_X1 U16309 ( .A1(n12890), .A2(P1_LWORD_REG_6__SCAN_IN), .ZN(n12881) );
  OAI211_X1 U16310 ( .C1(n12898), .C2(n19997), .A(n12881), .B(n12880), .ZN(
        P1_U2958) );
  INV_X1 U16311 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n19995) );
  NAND2_X1 U16312 ( .A1(n12890), .A2(P1_LWORD_REG_7__SCAN_IN), .ZN(n12883) );
  OAI211_X1 U16313 ( .C1(n12898), .C2(n19995), .A(n12883), .B(n12882), .ZN(
        P1_U2959) );
  INV_X1 U16314 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n19993) );
  NAND2_X1 U16315 ( .A1(n12890), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n12884) );
  OAI211_X1 U16316 ( .C1(n12898), .C2(n19993), .A(n12885), .B(n12884), .ZN(
        P1_U2960) );
  INV_X1 U16317 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n19991) );
  NAND2_X1 U16318 ( .A1(n12890), .A2(P1_LWORD_REG_9__SCAN_IN), .ZN(n12886) );
  OAI211_X1 U16319 ( .C1(n12898), .C2(n19991), .A(n12887), .B(n12886), .ZN(
        P1_U2961) );
  INV_X1 U16320 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n19989) );
  NAND2_X1 U16321 ( .A1(n12890), .A2(P1_LWORD_REG_10__SCAN_IN), .ZN(n12888) );
  OAI211_X1 U16322 ( .C1(n12898), .C2(n19989), .A(n12889), .B(n12888), .ZN(
        P1_U2962) );
  INV_X1 U16323 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n19987) );
  NAND2_X1 U16324 ( .A1(n12890), .A2(P1_LWORD_REG_11__SCAN_IN), .ZN(n12891) );
  OAI211_X1 U16325 ( .C1(n12898), .C2(n19987), .A(n12892), .B(n12891), .ZN(
        P1_U2963) );
  INV_X1 U16326 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n13808) );
  INV_X1 U16327 ( .A(n12893), .ZN(n12897) );
  INV_X1 U16328 ( .A(DATAI_15_), .ZN(n12895) );
  INV_X1 U16329 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n12894) );
  MUX2_X1 U16330 ( .A(n12895), .B(n12894), .S(n13387), .Z(n13807) );
  INV_X1 U16331 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n19978) );
  OAI222_X1 U16332 ( .A1(n12898), .A2(n13808), .B1(n12897), .B2(n13807), .C1(
        n12896), .C2(n19978), .ZN(P1_U2967) );
  NAND2_X1 U16333 ( .A1(n12899), .A2(n20105), .ZN(n12900) );
  OAI222_X1 U16334 ( .A1(n14285), .A2(n19970), .B1(n14353), .B2(n20007), .C1(
        n14352), .C2(n20082), .ZN(P1_U2903) );
  OAI222_X1 U16335 ( .A1(n14285), .A2(n13443), .B1(n14353), .B2(n20012), .C1(
        n14352), .C2(n20076), .ZN(P1_U2904) );
  OAI222_X1 U16336 ( .A1(n14285), .A2(n14200), .B1(n14353), .B2(n20005), .C1(
        n14352), .C2(n13395), .ZN(P1_U2902) );
  NAND2_X1 U16337 ( .A1(n12901), .A2(n13124), .ZN(n12902) );
  XNOR2_X1 U16338 ( .A(n12903), .B(n12902), .ZN(n12917) );
  NAND2_X1 U16339 ( .A1(n18898), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n12907) );
  NOR2_X1 U16340 ( .A1(n18955), .A2(n12904), .ZN(n12905) );
  AOI21_X1 U16341 ( .B1(n18963), .B2(P2_REIP_REG_2__SCAN_IN), .A(n12905), .ZN(
        n12906) );
  OAI211_X1 U16342 ( .C1(n18941), .C2(n13308), .A(n12907), .B(n12906), .ZN(
        n12908) );
  NAND2_X1 U16343 ( .A1(n12910), .A2(n12909), .ZN(n12913) );
  INV_X1 U16344 ( .A(n12911), .ZN(n12912) );
  NAND2_X1 U16345 ( .A1(n12913), .A2(n12912), .ZN(n19817) );
  NAND2_X1 U16346 ( .A1(n19817), .A2(n18907), .ZN(n12914) );
  OAI211_X1 U16347 ( .C1(n19813), .C2(n18966), .A(n12915), .B(n12914), .ZN(
        n12916) );
  AOI21_X1 U16348 ( .B1(n12917), .B2(n18951), .A(n12916), .ZN(n12918) );
  INV_X1 U16349 ( .A(n12918), .ZN(P2_U2853) );
  AND2_X1 U16350 ( .A1(n13570), .A2(n12919), .ZN(n12921) );
  OR2_X1 U16351 ( .A1(n12921), .A2(n12920), .ZN(n13700) );
  NAND2_X1 U16352 ( .A1(n12901), .A2(n12922), .ZN(n12923) );
  XNOR2_X1 U16353 ( .A(n16213), .B(n12923), .ZN(n12924) );
  NAND2_X1 U16354 ( .A1(n12924), .A2(n18951), .ZN(n12935) );
  OR2_X1 U16355 ( .A1(n12925), .A2(n13033), .ZN(n12926) );
  NAND2_X1 U16356 ( .A1(n12926), .A2(n13109), .ZN(n13108) );
  INV_X1 U16357 ( .A(n13108), .ZN(n16215) );
  XNOR2_X1 U16358 ( .A(n12928), .B(n12927), .ZN(n19013) );
  INV_X1 U16359 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19741) );
  OAI21_X1 U16360 ( .B1(n19741), .B2(n18923), .A(n18921), .ZN(n12931) );
  NOR2_X1 U16361 ( .A1(n18961), .A2(n12929), .ZN(n12930) );
  AOI211_X1 U16362 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n18957), .A(
        n12931), .B(n12930), .ZN(n12932) );
  OAI21_X1 U16363 ( .B1(n18960), .B2(n19013), .A(n12932), .ZN(n12933) );
  AOI21_X1 U16364 ( .B1(n18902), .B2(n16215), .A(n12933), .ZN(n12934) );
  OAI211_X1 U16365 ( .C1(n18941), .C2(n13700), .A(n12935), .B(n12934), .ZN(
        P2_U2849) );
  OAI21_X1 U16366 ( .B1(n12938), .B2(n12937), .A(n12936), .ZN(n20061) );
  INV_X1 U16367 ( .A(n14200), .ZN(n12941) );
  AOI22_X1 U16368 ( .A1(n20013), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n10704), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n12939) );
  OAI21_X1 U16369 ( .B1(n20023), .B2(n14190), .A(n12939), .ZN(n12940) );
  AOI21_X1 U16370 ( .B1(n12941), .B2(n14447), .A(n12940), .ZN(n12942) );
  OAI21_X1 U16371 ( .B1(n20030), .B2(n20061), .A(n12942), .ZN(P1_U2997) );
  NOR2_X1 U16372 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20648), .ZN(n12979) );
  INV_X1 U16373 ( .A(n12944), .ZN(n14197) );
  NAND4_X1 U16374 ( .A1(n12948), .A2(n12947), .A3(n12946), .A4(n12945), .ZN(
        n12967) );
  XNOR2_X1 U16375 ( .A(n14642), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14649) );
  NAND2_X1 U16376 ( .A1(n12950), .A2(n12949), .ZN(n12959) );
  NAND2_X1 U16377 ( .A1(n12959), .A2(n14649), .ZN(n12953) );
  XNOR2_X1 U16378 ( .A(n10080), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12951) );
  NAND2_X1 U16379 ( .A1(n12962), .A2(n12951), .ZN(n12952) );
  OAI211_X1 U16380 ( .C1(n12967), .C2(n14649), .A(n12953), .B(n12952), .ZN(
        n12954) );
  AOI21_X1 U16381 ( .B1(n14197), .B2(n14640), .A(n12954), .ZN(n14654) );
  INV_X1 U16382 ( .A(n14654), .ZN(n12955) );
  MUX2_X1 U16383 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n12955), .S(
        n12976), .Z(n15811) );
  AOI22_X1 U16384 ( .A1(n12979), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15811), .B2(n20648), .ZN(n12972) );
  NAND2_X1 U16385 ( .A1(n12956), .A2(n14640), .ZN(n12970) );
  AOI21_X1 U16386 ( .B1(n14642), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n9816), .ZN(n12957) );
  NOR2_X1 U16387 ( .A1(n12958), .A2(n12957), .ZN(n14658) );
  MUX2_X1 U16388 ( .A(n12964), .B(n9816), .S(n14642), .Z(n12960) );
  OAI21_X1 U16389 ( .B1(n12961), .B2(n12960), .A(n12959), .ZN(n12966) );
  MUX2_X1 U16390 ( .A(n12961), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n10080), .Z(n12963) );
  OAI21_X1 U16391 ( .B1(n12964), .B2(n12963), .A(n12962), .ZN(n12965) );
  OAI211_X1 U16392 ( .C1(n14658), .C2(n12967), .A(n12966), .B(n12965), .ZN(
        n12968) );
  INV_X1 U16393 ( .A(n12968), .ZN(n12969) );
  NAND2_X1 U16394 ( .A1(n12970), .A2(n12969), .ZN(n14656) );
  MUX2_X1 U16395 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14656), .S(
        n12976), .Z(n15802) );
  AOI22_X1 U16396 ( .A1(n12979), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n20648), .B2(n15802), .ZN(n12971) );
  NOR2_X1 U16397 ( .A1(n12972), .A2(n12971), .ZN(n15814) );
  INV_X1 U16398 ( .A(n14643), .ZN(n12973) );
  NAND2_X1 U16399 ( .A1(n15814), .A2(n12973), .ZN(n15832) );
  INV_X1 U16400 ( .A(n20218), .ZN(n20479) );
  OR2_X1 U16401 ( .A1(n12974), .A2(n20479), .ZN(n12975) );
  XNOR2_X1 U16402 ( .A(n12975), .B(n16116), .ZN(n19949) );
  OAI21_X1 U16403 ( .B1(n19949), .B2(n11561), .A(n12976), .ZN(n12978) );
  AOI21_X1 U16404 ( .B1(n15806), .B2(n16116), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n12977) );
  NAND2_X1 U16405 ( .A1(n12978), .A2(n12977), .ZN(n12981) );
  NAND2_X1 U16406 ( .A1(n12979), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12980) );
  NAND2_X1 U16407 ( .A1(n12981), .A2(n12980), .ZN(n15830) );
  NOR2_X1 U16408 ( .A1(n15830), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n12982) );
  AOI21_X1 U16409 ( .B1(n15832), .B2(n12982), .A(n16127), .ZN(n12983) );
  NOR2_X1 U16410 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20760) );
  OR2_X1 U16411 ( .A1(n12983), .A2(n20117), .ZN(n20740) );
  INV_X1 U16412 ( .A(n12988), .ZN(n12985) );
  NOR2_X1 U16413 ( .A1(n12984), .A2(n12985), .ZN(n20542) );
  INV_X1 U16414 ( .A(n12986), .ZN(n12996) );
  NAND2_X1 U16415 ( .A1(n20542), .A2(n12996), .ZN(n20511) );
  AOI211_X1 U16416 ( .C1(n20511), .C2(n20450), .A(P1_STATE2_REG_3__SCAN_IN), 
        .B(n12987), .ZN(n12993) );
  INV_X1 U16417 ( .A(n13379), .ZN(n12991) );
  NAND2_X1 U16418 ( .A1(n20738), .A2(n20515), .ZN(n20477) );
  NOR2_X1 U16419 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20648), .ZN(n20736) );
  INV_X1 U16420 ( .A(n20736), .ZN(n12998) );
  OR2_X1 U16421 ( .A1(n12984), .A2(n12988), .ZN(n20311) );
  AND2_X1 U16422 ( .A1(n20369), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12989) );
  NAND2_X1 U16423 ( .A1(n12986), .A2(n12989), .ZN(n14632) );
  NOR2_X1 U16424 ( .A1(n20311), .A2(n14632), .ZN(n20318) );
  AOI21_X1 U16425 ( .B1(n12956), .B2(n12998), .A(n20318), .ZN(n12990) );
  OAI21_X1 U16426 ( .B1(n12991), .B2(n20477), .A(n12990), .ZN(n12992) );
  OAI21_X1 U16427 ( .B1(n12993), .B2(n12992), .A(n20740), .ZN(n12994) );
  OAI21_X1 U16428 ( .B1(n20740), .B2(n20442), .A(n12994), .ZN(P1_U3475) );
  INV_X1 U16429 ( .A(n20740), .ZN(n20743) );
  OR2_X1 U16430 ( .A1(n12986), .A2(n20586), .ZN(n12995) );
  NAND2_X1 U16431 ( .A1(n12995), .A2(n20477), .ZN(n20590) );
  NAND2_X1 U16432 ( .A1(n12996), .A2(n20515), .ZN(n12999) );
  INV_X1 U16433 ( .A(n12997), .ZN(n20543) );
  AOI22_X1 U16434 ( .A1(n20590), .A2(n12999), .B1(n20543), .B2(n12998), .ZN(
        n13001) );
  NAND2_X1 U16435 ( .A1(n20743), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13000) );
  OAI21_X1 U16436 ( .B1(n20743), .B2(n13001), .A(n13000), .ZN(P1_U3477) );
  NAND2_X1 U16437 ( .A1(n13002), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13003) );
  NAND2_X2 U16438 ( .A1(n13006), .A2(n13005), .ZN(n13215) );
  INV_X1 U16439 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15646) );
  NOR2_X1 U16440 ( .A1(n14885), .A2(n15646), .ZN(n13052) );
  OR2_X1 U16441 ( .A1(n13188), .A2(n13052), .ZN(n13007) );
  NAND2_X1 U16442 ( .A1(n13188), .A2(n13052), .ZN(n13104) );
  NAND2_X1 U16443 ( .A1(n13007), .A2(n13104), .ZN(n19027) );
  OR2_X1 U16444 ( .A1(n13009), .A2(n13008), .ZN(n13010) );
  AND2_X1 U16445 ( .A1(n13010), .A2(n13034), .ZN(n19120) );
  INV_X1 U16446 ( .A(n19120), .ZN(n18964) );
  MUX2_X1 U16447 ( .A(n11848), .B(n18964), .S(n14743), .Z(n13011) );
  OAI21_X1 U16448 ( .B1(n19027), .B2(n15060), .A(n13011), .ZN(P2_U2883) );
  AOI22_X1 U16449 ( .A1(n20009), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20008), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13012) );
  OAI21_X1 U16450 ( .B1(n13013), .B2(n13031), .A(n13012), .ZN(P1_U2913) );
  AOI22_X1 U16451 ( .A1(n20009), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20008), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13014) );
  OAI21_X1 U16452 ( .B1(n13015), .B2(n13031), .A(n13014), .ZN(P1_U2912) );
  AOI22_X1 U16453 ( .A1(n20009), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20008), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13016) );
  OAI21_X1 U16454 ( .B1(n13017), .B2(n13031), .A(n13016), .ZN(P1_U2917) );
  AOI22_X1 U16455 ( .A1(n20009), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20008), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13018) );
  OAI21_X1 U16456 ( .B1(n13019), .B2(n13031), .A(n13018), .ZN(P1_U2916) );
  AOI22_X1 U16457 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20009), .B1(n20008), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13020) );
  OAI21_X1 U16458 ( .B1(n13021), .B2(n13031), .A(n13020), .ZN(P1_U2920) );
  AOI22_X1 U16459 ( .A1(n20009), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20008), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13022) );
  OAI21_X1 U16460 ( .B1(n13023), .B2(n13031), .A(n13022), .ZN(P1_U2910) );
  AOI22_X1 U16461 ( .A1(n20009), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20008), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13024) );
  OAI21_X1 U16462 ( .B1(n13025), .B2(n13031), .A(n13024), .ZN(P1_U2907) );
  AOI22_X1 U16463 ( .A1(n20009), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n20008), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13026) );
  OAI21_X1 U16464 ( .B1(n13027), .B2(n13031), .A(n13026), .ZN(P1_U2906) );
  AOI22_X1 U16465 ( .A1(n20009), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20008), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13028) );
  OAI21_X1 U16466 ( .B1(n13029), .B2(n13031), .A(n13028), .ZN(P1_U2918) );
  AOI22_X1 U16467 ( .A1(n20009), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20008), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13030) );
  OAI21_X1 U16468 ( .B1(n13032), .B2(n13031), .A(n13030), .ZN(P1_U2915) );
  XOR2_X1 U16469 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13104), .Z(n13038)
         );
  AOI21_X1 U16470 ( .B1(n13035), .B2(n13034), .A(n13033), .ZN(n18948) );
  NOR2_X1 U16471 ( .A1(n14743), .A2(n12306), .ZN(n13036) );
  AOI21_X1 U16472 ( .B1(n18948), .B2(n14743), .A(n13036), .ZN(n13037) );
  OAI21_X1 U16473 ( .B1(n13038), .B2(n15060), .A(n13037), .ZN(P2_U2882) );
  INV_X1 U16474 ( .A(n19817), .ZN(n19137) );
  INV_X1 U16475 ( .A(n19040), .ZN(n18983) );
  XNOR2_X1 U16476 ( .A(n19813), .B(n19817), .ZN(n13044) );
  XNOR2_X1 U16477 ( .A(n13040), .B(n13039), .ZN(n19826) );
  NOR2_X1 U16478 ( .A1(n19824), .A2(n19826), .ZN(n13041) );
  AOI21_X1 U16479 ( .B1(n19826), .B2(n19824), .A(n13041), .ZN(n19043) );
  NAND2_X1 U16480 ( .A1(n19043), .A2(n19042), .ZN(n19041) );
  INV_X1 U16481 ( .A(n13041), .ZN(n13042) );
  NAND2_X1 U16482 ( .A1(n19041), .A2(n13042), .ZN(n13043) );
  NAND2_X1 U16483 ( .A1(n13043), .A2(n13044), .ZN(n19016) );
  OAI21_X1 U16484 ( .B1(n13044), .B2(n13043), .A(n19016), .ZN(n13045) );
  NAND2_X1 U16485 ( .A1(n13045), .A2(n19044), .ZN(n13047) );
  AOI22_X1 U16486 ( .A1(n19008), .A2(n16152), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19039), .ZN(n13046) );
  OAI211_X1 U16487 ( .C1(n19137), .C2(n18983), .A(n13047), .B(n13046), .ZN(
        P2_U2917) );
  OR2_X1 U16488 ( .A1(n13048), .A2(n9701), .ZN(n13049) );
  NAND2_X1 U16489 ( .A1(n13049), .A2(n13063), .ZN(n15557) );
  AND2_X1 U16490 ( .A1(n13188), .A2(n13052), .ZN(n13050) );
  INV_X1 U16491 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19194) );
  NAND2_X1 U16492 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13103) );
  NOR2_X1 U16493 ( .A1(n19194), .A2(n13103), .ZN(n13051) );
  AND2_X1 U16494 ( .A1(n13050), .A2(n13051), .ZN(n13055) );
  AND2_X1 U16495 ( .A1(n13054), .A2(n13051), .ZN(n13053) );
  AND2_X1 U16496 ( .A1(n13053), .A2(n13052), .ZN(n13060) );
  NAND2_X1 U16497 ( .A1(n13188), .A2(n13060), .ZN(n13058) );
  OAI211_X1 U16498 ( .C1(n13055), .C2(n13054), .A(n13058), .B(n15047), .ZN(
        n13057) );
  NAND2_X1 U16499 ( .A1(n15050), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13056) );
  OAI211_X1 U16500 ( .C1(n15557), .C2(n15050), .A(n13057), .B(n13056), .ZN(
        P2_U2879) );
  INV_X1 U16501 ( .A(n13058), .ZN(n13062) );
  INV_X1 U16502 ( .A(n13059), .ZN(n13061) );
  NAND2_X1 U16503 ( .A1(n13188), .A2(n13074), .ZN(n13072) );
  OAI211_X1 U16504 ( .C1(n13062), .C2(n13061), .A(n15047), .B(n13072), .ZN(
        n13068) );
  NAND2_X1 U16505 ( .A1(n13064), .A2(n13063), .ZN(n13066) );
  INV_X1 U16506 ( .A(n13069), .ZN(n13065) );
  NAND2_X1 U16507 ( .A1(n13066), .A2(n13065), .ZN(n18935) );
  INV_X1 U16508 ( .A(n18935), .ZN(n13998) );
  NAND2_X1 U16509 ( .A1(n13998), .A2(n14743), .ZN(n13067) );
  OAI211_X1 U16510 ( .C1(n14743), .C2(n9880), .A(n13068), .B(n13067), .ZN(
        P2_U2878) );
  OR2_X1 U16511 ( .A1(n13070), .A2(n13069), .ZN(n13071) );
  AND2_X1 U16512 ( .A1(n13071), .A2(n13173), .ZN(n16201) );
  INV_X1 U16513 ( .A(n16201), .ZN(n18924) );
  INV_X1 U16514 ( .A(n13072), .ZN(n13077) );
  INV_X1 U16515 ( .A(n13073), .ZN(n13076) );
  AND2_X1 U16516 ( .A1(n13188), .A2(n13186), .ZN(n13191) );
  INV_X1 U16517 ( .A(n13191), .ZN(n13075) );
  OAI211_X1 U16518 ( .C1(n13077), .C2(n13076), .A(n13075), .B(n15047), .ZN(
        n13079) );
  NAND2_X1 U16519 ( .A1(n15050), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n13078) );
  OAI211_X1 U16520 ( .C1(n18924), .C2(n15055), .A(n13079), .B(n13078), .ZN(
        P2_U2877) );
  NOR2_X1 U16521 ( .A1(n9927), .A2(n13080), .ZN(n13081) );
  XNOR2_X1 U16522 ( .A(n13081), .B(n13369), .ZN(n13096) );
  NOR2_X1 U16523 ( .A1(n19445), .A2(n18966), .ZN(n13095) );
  OR2_X1 U16524 ( .A1(n13083), .A2(n13082), .ZN(n13084) );
  NAND2_X1 U16525 ( .A1(n13084), .A2(n13498), .ZN(n19018) );
  INV_X1 U16526 ( .A(n13480), .ZN(n13088) );
  NAND2_X1 U16527 ( .A1(n13086), .A2(n13085), .ZN(n13087) );
  NAND2_X1 U16528 ( .A1(n13088), .A2(n13087), .ZN(n13305) );
  INV_X1 U16529 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13371) );
  NOR2_X1 U16530 ( .A1(n18955), .A2(n13371), .ZN(n13089) );
  AOI21_X1 U16531 ( .B1(n18963), .B2(P2_REIP_REG_3__SCAN_IN), .A(n13089), .ZN(
        n13091) );
  NAND2_X1 U16532 ( .A1(n18898), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n13090) );
  OAI211_X1 U16533 ( .C1(n13305), .C2(n18941), .A(n13091), .B(n13090), .ZN(
        n13092) );
  AOI21_X1 U16534 ( .B1(n15615), .B2(n18902), .A(n13092), .ZN(n13093) );
  OAI21_X1 U16535 ( .B1(n19018), .B2(n18960), .A(n13093), .ZN(n13094) );
  AOI211_X1 U16536 ( .C1(n13096), .C2(n18951), .A(n13095), .B(n13094), .ZN(
        n13097) );
  INV_X1 U16537 ( .A(n13097), .ZN(P2_U2852) );
  OAI21_X1 U16538 ( .B1(n13099), .B2(n13098), .A(n13155), .ZN(n13515) );
  OAI222_X1 U16539 ( .A1(n14285), .A2(n13515), .B1(n14353), .B2(n20003), .C1(
        n14352), .C2(n20088), .ZN(P1_U2901) );
  AOI21_X1 U16540 ( .B1(n13101), .B2(n13100), .A(n13180), .ZN(n20046) );
  INV_X1 U16541 ( .A(n20046), .ZN(n13512) );
  INV_X1 U16542 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13102) );
  OAI222_X1 U16543 ( .A1(n13512), .A2(n14259), .B1(n13102), .B2(n14260), .C1(
        n13515), .C2(n14254), .ZN(P1_U2869) );
  NOR2_X1 U16544 ( .A1(n13104), .A2(n20797), .ZN(n13105) );
  OR2_X1 U16545 ( .A1(n13104), .A2(n13103), .ZN(n13137) );
  OAI211_X1 U16546 ( .C1(n13105), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n15047), .B(n13137), .ZN(n13107) );
  NAND2_X1 U16547 ( .A1(n15055), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n13106) );
  OAI211_X1 U16548 ( .C1(n13108), .C2(n15050), .A(n13107), .B(n13106), .ZN(
        P2_U2881) );
  AOI21_X1 U16549 ( .B1(n13110), .B2(n13109), .A(n9701), .ZN(n13111) );
  INV_X1 U16550 ( .A(n13111), .ZN(n15565) );
  NOR2_X1 U16551 ( .A1(n9927), .A2(n13112), .ZN(n13113) );
  XNOR2_X1 U16552 ( .A(n13113), .B(n15292), .ZN(n13114) );
  NAND2_X1 U16553 ( .A1(n13114), .A2(n18951), .ZN(n13123) );
  INV_X1 U16554 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19743) );
  INV_X1 U16555 ( .A(n13115), .ZN(n13116) );
  XNOR2_X1 U16556 ( .A(n12920), .B(n13116), .ZN(n13831) );
  AOI22_X1 U16557 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n18957), .B1(
        n18958), .B2(n13831), .ZN(n13117) );
  OAI211_X1 U16558 ( .C1(n19743), .C2(n18923), .A(n13117), .B(n18921), .ZN(
        n13121) );
  XNOR2_X1 U16559 ( .A(n13119), .B(n13118), .ZN(n19012) );
  NOR2_X1 U16560 ( .A1(n19012), .A2(n18960), .ZN(n13120) );
  AOI211_X1 U16561 ( .C1(P2_EBX_REG_7__SCAN_IN), .C2(n18898), .A(n13121), .B(
        n13120), .ZN(n13122) );
  OAI211_X1 U16562 ( .C1(n15565), .C2(n18965), .A(n13123), .B(n13122), .ZN(
        P2_U2848) );
  NAND2_X1 U16563 ( .A1(n18951), .A2(n9927), .ZN(n18914) );
  OAI211_X1 U16564 ( .C1(n13196), .C2(n13125), .A(n12901), .B(n13124), .ZN(
        n15585) );
  OAI22_X1 U16565 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18914), .B1(
        n15585), .B2(n19713), .ZN(n13126) );
  INV_X1 U16566 ( .A(n13126), .ZN(n13136) );
  NAND2_X1 U16567 ( .A1(n19826), .A2(n18907), .ZN(n13133) );
  INV_X1 U16568 ( .A(n13127), .ZN(n13128) );
  NAND2_X1 U16569 ( .A1(n18958), .A2(n13128), .ZN(n13129) );
  OAI21_X1 U16570 ( .B1(n13130), .B2(n18955), .A(n13129), .ZN(n13131) );
  AOI21_X1 U16571 ( .B1(n18963), .B2(P2_REIP_REG_1__SCAN_IN), .A(n13131), .ZN(
        n13132) );
  OAI211_X1 U16572 ( .C1(n11783), .C2(n18961), .A(n13133), .B(n13132), .ZN(
        n13134) );
  AOI21_X1 U16573 ( .B1(n19157), .B2(n18902), .A(n13134), .ZN(n13135) );
  OAI211_X1 U16574 ( .C1(n18966), .C2(n19814), .A(n13136), .B(n13135), .ZN(
        P2_U2854) );
  XOR2_X1 U16575 ( .A(n13137), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13139)
         );
  MUX2_X1 U16576 ( .A(n12308), .B(n15565), .S(n14743), .Z(n13138) );
  OAI21_X1 U16577 ( .B1(n13139), .B2(n15060), .A(n13138), .ZN(P2_U2880) );
  NAND2_X1 U16578 ( .A1(n13141), .A2(n13140), .ZN(n13142) );
  NAND2_X1 U16579 ( .A1(n13824), .A2(n13142), .ZN(n13823) );
  NAND2_X1 U16580 ( .A1(n12901), .A2(n13143), .ZN(n13144) );
  XNOR2_X1 U16581 ( .A(n16206), .B(n13144), .ZN(n13145) );
  NAND2_X1 U16582 ( .A1(n13145), .A2(n18951), .ZN(n13154) );
  INV_X1 U16583 ( .A(n15557), .ZN(n16207) );
  AOI21_X1 U16584 ( .B1(n13147), .B2(n13146), .A(n9682), .ZN(n19007) );
  INV_X1 U16585 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n19745) );
  OAI21_X1 U16586 ( .B1(n19745), .B2(n18923), .A(n18921), .ZN(n13149) );
  NOR2_X1 U16587 ( .A1(n18955), .A2(n16212), .ZN(n13148) );
  AOI211_X1 U16588 ( .C1(n18907), .C2(n19007), .A(n13149), .B(n13148), .ZN(
        n13150) );
  OAI21_X1 U16589 ( .B1(n18961), .B2(n13151), .A(n13150), .ZN(n13152) );
  AOI21_X1 U16590 ( .B1(n16207), .B2(n18902), .A(n13152), .ZN(n13153) );
  OAI211_X1 U16591 ( .C1(n18941), .C2(n13823), .A(n13154), .B(n13153), .ZN(
        P2_U2847) );
  XOR2_X1 U16592 ( .A(n13156), .B(n13155), .Z(n20018) );
  INV_X1 U16593 ( .A(n20018), .ZN(n13181) );
  AOI22_X1 U16594 ( .A1(n13772), .A2(n14320), .B1(P1_EAX_REG_4__SCAN_IN), .B2(
        n14342), .ZN(n13157) );
  OAI21_X1 U16595 ( .B1(n13181), .B2(n14285), .A(n13157), .ZN(P1_U2900) );
  OAI21_X1 U16596 ( .B1(n13160), .B2(n13159), .A(n13158), .ZN(n13161) );
  INV_X1 U16597 ( .A(n13161), .ZN(n20049) );
  NAND2_X1 U16598 ( .A1(n20049), .A2(n20019), .ZN(n13165) );
  INV_X1 U16599 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n13162) );
  NOR2_X1 U16600 ( .A1(n20036), .A2(n13162), .ZN(n20045) );
  NOR2_X1 U16601 ( .A1(n20023), .A2(n13508), .ZN(n13163) );
  AOI211_X1 U16602 ( .C1(n20013), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20045), .B(n13163), .ZN(n13164) );
  OAI211_X1 U16603 ( .C1(n15947), .C2(n13515), .A(n13165), .B(n13164), .ZN(
        P1_U2996) );
  OR2_X1 U16604 ( .A1(n13167), .A2(n13166), .ZN(n14255) );
  NAND2_X1 U16605 ( .A1(n13167), .A2(n13166), .ZN(n13168) );
  NAND2_X1 U16606 ( .A1(n14255), .A2(n13168), .ZN(n16003) );
  INV_X1 U16607 ( .A(n14258), .ZN(n13169) );
  AOI21_X1 U16608 ( .B1(n13170), .B2(n13178), .A(n13169), .ZN(n16103) );
  AOI22_X1 U16609 ( .A1(n16103), .A2(n14223), .B1(P1_EBX_REG_5__SCAN_IN), .B2(
        n14222), .ZN(n13171) );
  OAI21_X1 U16610 ( .B1(n16003), .B2(n14254), .A(n13171), .ZN(P1_U2867) );
  XNOR2_X1 U16611 ( .A(n13191), .B(n13190), .ZN(n13177) );
  NAND2_X1 U16612 ( .A1(n13173), .A2(n13172), .ZN(n13174) );
  AND2_X1 U16613 ( .A1(n13184), .A2(n13174), .ZN(n18903) );
  NOR2_X1 U16614 ( .A1(n14743), .A2(n11866), .ZN(n13175) );
  AOI21_X1 U16615 ( .B1(n18903), .B2(n14743), .A(n13175), .ZN(n13176) );
  OAI21_X1 U16616 ( .B1(n13177), .B2(n15060), .A(n13176), .ZN(P2_U2876) );
  OAI21_X1 U16617 ( .B1(n13180), .B2(n13179), .A(n13178), .ZN(n20037) );
  INV_X1 U16618 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13182) );
  OAI222_X1 U16619 ( .A1(n20037), .A2(n14259), .B1(n13182), .B2(n14260), .C1(
        n14254), .C2(n13181), .ZN(P1_U2868) );
  AND2_X1 U16620 ( .A1(n13184), .A2(n13183), .ZN(n13185) );
  NOR2_X1 U16621 ( .A1(n13220), .A2(n13185), .ZN(n16186) );
  INV_X1 U16622 ( .A(n16186), .ZN(n18893) );
  AND2_X1 U16623 ( .A1(n13189), .A2(n13190), .ZN(n13187) );
  AND2_X1 U16624 ( .A1(n13188), .A2(n13213), .ZN(n13217) );
  AOI21_X1 U16625 ( .B1(n13191), .B2(n13190), .A(n13189), .ZN(n13192) );
  OR3_X1 U16626 ( .A1(n13217), .A2(n13192), .A3(n15060), .ZN(n13194) );
  NAND2_X1 U16627 ( .A1(n15055), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13193) );
  OAI211_X1 U16628 ( .C1(n18893), .C2(n15050), .A(n13194), .B(n13193), .ZN(
        P2_U2875) );
  INV_X1 U16629 ( .A(n18914), .ZN(n13195) );
  OAI21_X1 U16630 ( .B1(n18957), .B2(n13195), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13204) );
  NOR2_X1 U16631 ( .A1(n9927), .A2(n19713), .ZN(n18831) );
  INV_X1 U16632 ( .A(n13196), .ZN(n15577) );
  AOI22_X1 U16633 ( .A1(n18963), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n18831), 
        .B2(n15577), .ZN(n13198) );
  NAND2_X1 U16634 ( .A1(n16245), .A2(n18907), .ZN(n13197) );
  OAI211_X1 U16635 ( .C1(n18961), .C2(n13199), .A(n13198), .B(n13197), .ZN(
        n13201) );
  NOR2_X1 U16636 ( .A1(n16249), .A2(n18965), .ZN(n13200) );
  AOI211_X1 U16637 ( .C1(n18958), .C2(n13202), .A(n13201), .B(n13200), .ZN(
        n13203) );
  OAI211_X1 U16638 ( .C1(n18966), .C2(n19834), .A(n13204), .B(n13203), .ZN(
        P2_U2855) );
  OR2_X1 U16639 ( .A1(n13207), .A2(n13206), .ZN(n13208) );
  AND2_X1 U16640 ( .A1(n13205), .A2(n13208), .ZN(n15992) );
  OR2_X1 U16641 ( .A1(n13210), .A2(n13209), .ZN(n13211) );
  AND2_X1 U16642 ( .A1(n13417), .A2(n13211), .ZN(n19932) );
  AOI22_X1 U16643 ( .A1(n19932), .A2(n14223), .B1(P1_EBX_REG_7__SCAN_IN), .B2(
        n14222), .ZN(n13212) );
  OAI21_X1 U16644 ( .B1(n19929), .B2(n14254), .A(n13212), .ZN(P1_U2865) );
  OAI222_X1 U16645 ( .A1(n14285), .A2(n19929), .B1(n14353), .B2(n19995), .C1(
        n14352), .C2(n20108), .ZN(P1_U2897) );
  INV_X1 U16646 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n18875) );
  OAI211_X1 U16647 ( .C1(n13217), .C2(n13216), .A(n13405), .B(n15047), .ZN(
        n13223) );
  OR2_X1 U16648 ( .A1(n13220), .A2(n13219), .ZN(n13221) );
  NAND2_X1 U16649 ( .A1(n13218), .A2(n13221), .ZN(n18881) );
  INV_X1 U16650 ( .A(n18881), .ZN(n15481) );
  NAND2_X1 U16651 ( .A1(n15481), .A2(n14743), .ZN(n13222) );
  OAI211_X1 U16652 ( .C1(n14743), .C2(n18875), .A(n13223), .B(n13222), .ZN(
        P2_U2874) );
  NOR3_X1 U16653 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19819), .A3(
        n19811), .ZN(n19573) );
  NAND2_X1 U16654 ( .A1(n19573), .A2(n19839), .ZN(n13241) );
  NAND2_X1 U16655 ( .A1(n13269), .A2(n16249), .ZN(n13260) );
  OAI21_X1 U16656 ( .B1(n13669), .B2(n19852), .A(n19416), .ZN(n13233) );
  OAI21_X1 U16657 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(
        P2_STATE2_REG_1__SCAN_IN), .A(n11587), .ZN(n19863) );
  INV_X1 U16658 ( .A(n19863), .ZN(n13225) );
  AOI21_X4 U16659 ( .B1(n19831), .B2(n13225), .A(n16297), .ZN(n19650) );
  INV_X1 U16660 ( .A(n13226), .ZN(n13227) );
  NOR2_X1 U16661 ( .A1(n13227), .A2(n13423), .ZN(n19307) );
  INV_X1 U16662 ( .A(n19597), .ZN(n13229) );
  INV_X1 U16663 ( .A(n19568), .ZN(n13228) );
  INV_X1 U16664 ( .A(n19565), .ZN(n13230) );
  AOI21_X1 U16665 ( .B1(n19591), .B2(n19552), .A(n15620), .ZN(n13231) );
  AOI21_X1 U16666 ( .B1(n19307), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n13231), .ZN(n13232) );
  AOI211_X1 U16667 ( .C1(n13241), .C2(n13233), .A(n19650), .B(n13232), .ZN(
        n19541) );
  INV_X1 U16668 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13244) );
  INV_X1 U16669 ( .A(n13234), .ZN(n13237) );
  INV_X1 U16670 ( .A(n19307), .ZN(n13236) );
  INV_X1 U16671 ( .A(n13241), .ZN(n19559) );
  OAI21_X1 U16672 ( .B1(n13669), .B2(n19559), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13235) );
  OAI21_X1 U16673 ( .B1(n13237), .B2(n13236), .A(n13235), .ZN(n19560) );
  NOR2_X2 U16674 ( .A1(n13238), .A2(n19650), .ZN(n19646) );
  NOR2_X2 U16675 ( .A1(n13344), .A2(n19186), .ZN(n19645) );
  INV_X1 U16676 ( .A(n19645), .ZN(n19200) );
  AOI22_X1 U16677 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19190), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19189), .ZN(n19578) );
  INV_X1 U16678 ( .A(n19552), .ZN(n19561) );
  AOI22_X1 U16679 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19190), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19189), .ZN(n19660) );
  AOI22_X1 U16680 ( .A1(n19593), .A2(n19657), .B1(n19561), .B2(n19575), .ZN(
        n13240) );
  OAI21_X1 U16681 ( .B1(n19200), .B2(n13241), .A(n13240), .ZN(n13242) );
  AOI21_X1 U16682 ( .B1(n19560), .B2(n19646), .A(n13242), .ZN(n13243) );
  OAI21_X1 U16683 ( .B1(n19541), .B2(n13244), .A(n13243), .ZN(P2_U3144) );
  NOR2_X1 U16684 ( .A1(n13260), .A2(n13267), .ZN(n13245) );
  AOI22_X1 U16685 ( .A1(n13545), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13669), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13258) );
  AND2_X1 U16686 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n13267), .ZN(
        n13246) );
  NAND2_X1 U16687 ( .A1(n13246), .A2(n13286), .ZN(n13257) );
  INV_X1 U16688 ( .A(n13271), .ZN(n13249) );
  INV_X1 U16689 ( .A(n12595), .ZN(n13247) );
  AND2_X1 U16690 ( .A1(n13247), .A2(n13252), .ZN(n13250) );
  INV_X1 U16691 ( .A(n13250), .ZN(n13248) );
  NAND2_X1 U16692 ( .A1(n13269), .A2(n13250), .ZN(n13263) );
  INV_X1 U16693 ( .A(n13263), .ZN(n13251) );
  AND2_X1 U16694 ( .A1(n13271), .A2(n13251), .ZN(n13296) );
  AND2_X1 U16695 ( .A1(n12595), .A2(n13252), .ZN(n13275) );
  INV_X1 U16696 ( .A(n13275), .ZN(n13253) );
  NOR2_X1 U16697 ( .A1(n13269), .A2(n13253), .ZN(n13254) );
  AOI22_X1 U16698 ( .A1(n13287), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n19453), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13255) );
  NOR2_X2 U16699 ( .A1(n13259), .A2(n13267), .ZN(n15651) );
  NAND2_X1 U16700 ( .A1(n13249), .A2(n13224), .ZN(n13261) );
  NOR2_X2 U16701 ( .A1(n13261), .A2(n19157), .ZN(n13544) );
  AOI22_X1 U16702 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n15651), .B1(
        n13544), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13280) );
  INV_X1 U16703 ( .A(n13261), .ZN(n13262) );
  NAND2_X1 U16704 ( .A1(n13262), .A2(n19157), .ZN(n13425) );
  NOR2_X2 U16705 ( .A1(n13271), .A2(n13263), .ZN(n19388) );
  AND2_X1 U16706 ( .A1(n13271), .A2(n13264), .ZN(n13291) );
  AOI22_X1 U16707 ( .A1(n19388), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13291), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13265) );
  OAI21_X1 U16708 ( .B1(n13425), .B2(n13266), .A(n13265), .ZN(n13274) );
  AND2_X1 U16709 ( .A1(n13269), .A2(n13275), .ZN(n13270) );
  AOI22_X1 U16710 ( .A1(n19422), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n19569), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13272) );
  INV_X1 U16711 ( .A(n13272), .ZN(n13273) );
  NOR2_X1 U16712 ( .A1(n13274), .A2(n13273), .ZN(n13279) );
  NOR2_X2 U16713 ( .A1(n13277), .A2(n13276), .ZN(n19335) );
  AOI22_X1 U16714 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19335), .B1(
        n19197), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13278) );
  NAND4_X1 U16715 ( .A1(n13281), .A2(n13280), .A3(n13279), .A4(n13278), .ZN(
        n13282) );
  NAND2_X1 U16716 ( .A1(n13282), .A2(n14935), .ZN(n13285) );
  INV_X1 U16717 ( .A(n10101), .ZN(n13283) );
  NAND2_X1 U16718 ( .A1(n13283), .A2(n11798), .ZN(n13284) );
  INV_X1 U16719 ( .A(n13425), .ZN(n13674) );
  NAND2_X1 U16720 ( .A1(n15629), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13289) );
  AOI22_X1 U16721 ( .A1(n19388), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13291), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13295) );
  NAND2_X1 U16722 ( .A1(n19335), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n13294) );
  NAND2_X1 U16723 ( .A1(n19197), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13293) );
  AOI22_X1 U16724 ( .A1(n19422), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n19569), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13292) );
  AOI21_X1 U16725 ( .B1(n19453), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A(
        n11798), .ZN(n13298) );
  AOI22_X1 U16726 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n13669), .B1(
        n13545), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13297) );
  AOI22_X1 U16727 ( .A1(n13544), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n15651), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13300) );
  NAND2_X1 U16728 ( .A1(n13303), .A2(n13302), .ZN(n13488) );
  NAND2_X1 U16729 ( .A1(n13484), .A2(n13905), .ZN(n13306) );
  NAND2_X1 U16730 ( .A1(n13306), .A2(n13305), .ZN(n13575) );
  NOR2_X1 U16731 ( .A1(n13575), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13476) );
  INV_X1 U16732 ( .A(n13476), .ZN(n13307) );
  NAND2_X1 U16733 ( .A1(n13575), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13477) );
  NAND2_X1 U16734 ( .A1(n13307), .A2(n13477), .ZN(n13311) );
  INV_X1 U16735 ( .A(n13308), .ZN(n13309) );
  NAND2_X1 U16736 ( .A1(n13309), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13310) );
  NAND2_X1 U16737 ( .A1(n19132), .A2(n13310), .ZN(n13579) );
  INV_X1 U16738 ( .A(n13579), .ZN(n13478) );
  XNOR2_X1 U16739 ( .A(n13311), .B(n13478), .ZN(n13377) );
  INV_X1 U16740 ( .A(n13312), .ZN(n16280) );
  NAND2_X1 U16741 ( .A1(n13316), .A2(n16280), .ZN(n13325) );
  AOI21_X1 U16742 ( .B1(n13313), .B2(n13344), .A(n13345), .ZN(n13314) );
  NAND2_X1 U16743 ( .A1(n19053), .A2(n13314), .ZN(n13324) );
  MUX2_X1 U16744 ( .A(n13316), .B(n13315), .S(n14935), .Z(n13317) );
  NAND3_X1 U16745 ( .A1(n13317), .A2(n16271), .A3(n19859), .ZN(n13320) );
  NAND2_X1 U16746 ( .A1(n14935), .A2(n19848), .ZN(n13318) );
  OR2_X1 U16747 ( .A1(n16276), .A2(n13318), .ZN(n13319) );
  AND4_X1 U16748 ( .A1(n13322), .A2(n13321), .A3(n13320), .A4(n13319), .ZN(
        n13323) );
  OAI211_X1 U16749 ( .C1(n19053), .C2(n13325), .A(n13324), .B(n13323), .ZN(
        n13326) );
  NAND2_X1 U16750 ( .A1(n13326), .A2(n19708), .ZN(n13357) );
  INV_X1 U16751 ( .A(n13327), .ZN(n19849) );
  NAND2_X1 U16752 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13328), .ZN(
        n13329) );
  NAND2_X1 U16753 ( .A1(n13330), .A2(n13329), .ZN(n13485) );
  INV_X1 U16754 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13363) );
  XNOR2_X1 U16755 ( .A(n13485), .B(n13363), .ZN(n13483) );
  XOR2_X1 U16756 ( .A(n13484), .B(n13483), .Z(n13374) );
  NAND2_X1 U16757 ( .A1(n11807), .A2(n14935), .ZN(n13331) );
  AND2_X1 U16758 ( .A1(n16272), .A2(n13331), .ZN(n13332) );
  NAND2_X1 U16759 ( .A1(n15587), .A2(n11798), .ZN(n13334) );
  AND2_X1 U16760 ( .A1(n15591), .A2(n13334), .ZN(n13335) );
  NAND2_X1 U16761 ( .A1(n13336), .A2(n14935), .ZN(n15572) );
  NAND2_X1 U16762 ( .A1(n15572), .A2(n13337), .ZN(n13338) );
  NAND2_X1 U16763 ( .A1(n13338), .A2(n11768), .ZN(n13351) );
  NAND2_X1 U16764 ( .A1(n13340), .A2(n13339), .ZN(n13341) );
  NAND2_X1 U16765 ( .A1(n13341), .A2(n12440), .ZN(n13343) );
  NAND2_X1 U16766 ( .A1(n13343), .A2(n13342), .ZN(n13348) );
  OAI22_X1 U16767 ( .A1(n12440), .A2(n13345), .B1(n13436), .B2(n13344), .ZN(
        n13346) );
  INV_X1 U16768 ( .A(n13346), .ZN(n13347) );
  AND3_X1 U16769 ( .A1(n13349), .A2(n13348), .A3(n13347), .ZN(n13350) );
  NAND2_X1 U16770 ( .A1(n13351), .A2(n13350), .ZN(n15614) );
  NOR2_X1 U16771 ( .A1(n15614), .A2(n13352), .ZN(n13353) );
  NOR2_X1 U16772 ( .A1(n13357), .A2(n13353), .ZN(n15466) );
  INV_X1 U16773 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19151) );
  NOR2_X1 U16774 ( .A1(n19151), .A2(n19150), .ZN(n19149) );
  INV_X1 U16775 ( .A(n19149), .ZN(n13354) );
  NAND2_X1 U16776 ( .A1(n15466), .A2(n13354), .ZN(n13355) );
  AND2_X1 U16777 ( .A1(n13357), .A2(n18921), .ZN(n19154) );
  INV_X1 U16778 ( .A(n19154), .ZN(n16250) );
  NAND2_X1 U16779 ( .A1(n13355), .A2(n16250), .ZN(n19142) );
  INV_X1 U16780 ( .A(n16274), .ZN(n13356) );
  NOR2_X1 U16781 ( .A1(n13357), .A2(n13356), .ZN(n19143) );
  NOR2_X1 U16782 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19149), .ZN(
        n19145) );
  AND2_X1 U16783 ( .A1(n19143), .A2(n19145), .ZN(n13359) );
  AND2_X1 U16784 ( .A1(n15466), .A2(n13358), .ZN(n19133) );
  INV_X1 U16785 ( .A(n13701), .ZN(n13958) );
  INV_X1 U16786 ( .A(n19145), .ZN(n13360) );
  NAND2_X1 U16787 ( .A1(n19143), .A2(n13360), .ZN(n13362) );
  AND2_X1 U16788 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19149), .ZN(
        n19144) );
  NAND2_X1 U16789 ( .A1(n15466), .A2(n19144), .ZN(n13361) );
  NAND2_X1 U16790 ( .A1(n13362), .A2(n13361), .ZN(n13954) );
  AOI22_X1 U16791 ( .A1(n13954), .A2(n13363), .B1(n19119), .B2(
        P2_REIP_REG_3__SCAN_IN), .ZN(n13364) );
  OAI21_X1 U16792 ( .B1(n13958), .B2(n13363), .A(n13364), .ZN(n13365) );
  AOI21_X1 U16793 ( .B1(n19156), .B2(n15615), .A(n13365), .ZN(n13366) );
  OAI21_X1 U16794 ( .B1(n19018), .B2(n19136), .A(n13366), .ZN(n13367) );
  AOI21_X1 U16795 ( .B1(n13374), .B2(n16228), .A(n13367), .ZN(n13368) );
  OAI21_X1 U16796 ( .B1(n13377), .B2(n19166), .A(n13368), .ZN(P2_U3043) );
  NOR2_X1 U16797 ( .A1(n16190), .A2(n13369), .ZN(n13373) );
  INV_X1 U16798 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n13370) );
  OAI22_X1 U16799 ( .A1(n19129), .A2(n13371), .B1(n13370), .B2(n18921), .ZN(
        n13372) );
  AOI211_X1 U16800 ( .C1(n15615), .C2(n19121), .A(n13373), .B(n13372), .ZN(
        n13376) );
  NAND2_X1 U16801 ( .A1(n13374), .A2(n19123), .ZN(n13375) );
  OAI211_X1 U16802 ( .C1(n13377), .C2(n16192), .A(n13376), .B(n13375), .ZN(
        P2_U3011) );
  INV_X1 U16803 ( .A(n12984), .ZN(n13378) );
  NAND2_X1 U16804 ( .A1(n20542), .A2(n20312), .ZN(n20629) );
  OAI21_X1 U16805 ( .B1(n20127), .B2(n20642), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n13380) );
  NAND2_X1 U16806 ( .A1(n13380), .A2(n20738), .ZN(n13386) );
  OR2_X1 U16807 ( .A1(n14197), .A2(n12956), .ZN(n20146) );
  NAND2_X1 U16808 ( .A1(n20184), .A2(n12997), .ZN(n13381) );
  NAND2_X1 U16809 ( .A1(n20340), .A2(n20399), .ZN(n20220) );
  NOR2_X1 U16810 ( .A1(n13382), .A2(n20652), .ZN(n20223) );
  INV_X1 U16811 ( .A(n20223), .ZN(n20405) );
  OAI22_X1 U16812 ( .A1(n13386), .A2(n13381), .B1(n20220), .B2(n20405), .ZN(
        n20110) );
  INV_X1 U16813 ( .A(n20110), .ZN(n13402) );
  INV_X1 U16814 ( .A(n20618), .ZN(n13394) );
  INV_X1 U16815 ( .A(n13381), .ZN(n13385) );
  NAND3_X1 U16816 ( .A1(n20442), .A2(n20395), .A3(n20475), .ZN(n20116) );
  NOR2_X1 U16817 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20116), .ZN(
        n13397) );
  INV_X1 U16818 ( .A(n13397), .ZN(n20106) );
  NAND2_X1 U16819 ( .A1(n13382), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20544) );
  NAND2_X1 U16820 ( .A1(n20117), .A2(n20544), .ZN(n20342) );
  AOI21_X1 U16821 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20106), .A(n20342), 
        .ZN(n13384) );
  NAND2_X1 U16822 ( .A1(n20220), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13383) );
  OAI211_X1 U16823 ( .C1(n13386), .C2(n13385), .A(n13384), .B(n13383), .ZN(
        n20073) );
  NOR2_X2 U16824 ( .A1(n15947), .A2(n13389), .ZN(n20109) );
  AOI22_X1 U16825 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20109), .B1(DATAI_28_), 
        .B2(n13388), .ZN(n20622) );
  INV_X1 U16826 ( .A(n20622), .ZN(n20565) );
  AOI22_X1 U16827 ( .A1(n20642), .A2(n20565), .B1(n13397), .B2(n20617), .ZN(
        n13391) );
  OAI21_X1 U16828 ( .B1(n20568), .B2(n20141), .A(n13391), .ZN(n13392) );
  AOI21_X1 U16829 ( .B1(n20073), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A(
        n13392), .ZN(n13393) );
  OAI21_X1 U16830 ( .B1(n13402), .B2(n13394), .A(n13393), .ZN(P1_U3037) );
  NOR2_X2 U16831 ( .A1(n13395), .A2(n20224), .ZN(n20606) );
  INV_X1 U16832 ( .A(n20606), .ZN(n13401) );
  AOI22_X1 U16833 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20109), .B1(DATAI_18_), 
        .B2(n13388), .ZN(n20560) );
  INV_X1 U16834 ( .A(n20610), .ZN(n20557) );
  AOI22_X1 U16835 ( .A1(n20642), .A2(n20557), .B1(n13397), .B2(n20605), .ZN(
        n13398) );
  OAI21_X1 U16836 ( .B1(n20560), .B2(n20141), .A(n13398), .ZN(n13399) );
  AOI21_X1 U16837 ( .B1(n20073), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n13399), .ZN(n13400) );
  OAI21_X1 U16838 ( .B1(n13402), .B2(n13401), .A(n13400), .ZN(P1_U3035) );
  NAND2_X1 U16839 ( .A1(n13218), .A2(n13403), .ZN(n13404) );
  AND2_X1 U16840 ( .A1(n13527), .A2(n13404), .ZN(n18870) );
  INV_X1 U16841 ( .A(n18870), .ZN(n13411) );
  INV_X1 U16842 ( .A(n13405), .ZN(n13408) );
  INV_X1 U16843 ( .A(n13406), .ZN(n13407) );
  OAI211_X1 U16844 ( .C1(n13408), .C2(n13407), .A(n15047), .B(n13529), .ZN(
        n13410) );
  NAND2_X1 U16845 ( .A1(n15050), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n13409) );
  OAI211_X1 U16846 ( .C1(n13411), .C2(n15055), .A(n13410), .B(n13409), .ZN(
        P2_U2873) );
  INV_X1 U16847 ( .A(n13412), .ZN(n13413) );
  AOI21_X1 U16848 ( .B1(n13414), .B2(n13205), .A(n13413), .ZN(n19919) );
  INV_X1 U16849 ( .A(n19919), .ZN(n13420) );
  AOI22_X1 U16850 ( .A1(n13772), .A2(n14299), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n14342), .ZN(n13415) );
  OAI21_X1 U16851 ( .B1(n13420), .B2(n14285), .A(n13415), .ZN(P1_U2896) );
  INV_X1 U16852 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13419) );
  NAND2_X1 U16853 ( .A1(n13417), .A2(n13416), .ZN(n13418) );
  NAND2_X1 U16854 ( .A1(n13470), .A2(n13418), .ZN(n19917) );
  OAI222_X1 U16855 ( .A1(n13420), .A2(n14254), .B1(n14260), .B2(n13419), .C1(
        n19917), .C2(n14259), .ZN(P1_U2864) );
  NAND2_X1 U16856 ( .A1(n19445), .A2(n13421), .ZN(n19386) );
  NOR2_X2 U16857 ( .A1(n19798), .A2(n19309), .ZN(n19411) );
  OAI21_X1 U16858 ( .B1(n19367), .B2(n19411), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13424) );
  NAND2_X1 U16859 ( .A1(n19811), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19387) );
  INV_X1 U16860 ( .A(n19387), .ZN(n13422) );
  NAND2_X1 U16861 ( .A1(n13423), .A2(n13422), .ZN(n13434) );
  NAND2_X1 U16862 ( .A1(n13424), .A2(n13434), .ZN(n13430) );
  NOR2_X1 U16863 ( .A1(n19479), .A2(n19387), .ZN(n19380) );
  INV_X1 U16864 ( .A(n19380), .ZN(n13426) );
  AND2_X1 U16865 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n13426), .ZN(n13427) );
  NAND2_X1 U16866 ( .A1(n13425), .A2(n13427), .ZN(n13432) );
  OAI211_X1 U16867 ( .C1(n19380), .C2(n19416), .A(n13432), .B(n19604), .ZN(
        n13428) );
  INV_X1 U16868 ( .A(n13428), .ZN(n13429) );
  INV_X1 U16869 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13439) );
  AOI22_X1 U16870 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19190), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19189), .ZN(n19547) );
  AOI22_X1 U16871 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19189), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19190), .ZN(n19672) );
  INV_X1 U16872 ( .A(n19672), .ZN(n19544) );
  AOI22_X1 U16873 ( .A1(n19411), .A2(n19669), .B1(n19367), .B2(n19544), .ZN(
        n13438) );
  INV_X1 U16874 ( .A(n13431), .ZN(n19389) );
  INV_X1 U16875 ( .A(n13432), .ZN(n13433) );
  AOI211_X2 U16876 ( .C1(n19852), .C2(n13434), .A(n19389), .B(n13433), .ZN(
        n19381) );
  NOR2_X2 U16877 ( .A1(n13435), .A2(n19650), .ZN(n19668) );
  NOR2_X2 U16878 ( .A1(n13436), .A2(n19186), .ZN(n19667) );
  AOI22_X1 U16879 ( .A1(n19381), .A2(n19668), .B1(n19667), .B2(n19380), .ZN(
        n13437) );
  OAI211_X1 U16880 ( .C1(n19371), .C2(n13439), .A(n13438), .B(n13437), .ZN(
        P2_U3098) );
  NOR2_X1 U16881 ( .A1(n20757), .A2(n13440), .ZN(n13455) );
  NAND2_X1 U16882 ( .A1(n20080), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13452) );
  AND2_X1 U16883 ( .A1(n20659), .A2(n20515), .ZN(n13441) );
  NOR2_X1 U16884 ( .A1(n13452), .A2(n13441), .ZN(n13442) );
  INV_X1 U16885 ( .A(n13443), .ZN(n20027) );
  NAND2_X1 U16886 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20760), .ZN(n16118) );
  NOR2_X1 U16887 ( .A1(n16118), .A2(n20649), .ZN(n13447) );
  NAND2_X1 U16888 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20649), .ZN(n13445) );
  OAI21_X1 U16889 ( .B1(n13445), .B2(n13444), .A(n20036), .ZN(n13446) );
  NOR2_X1 U16890 ( .A1(n13457), .A2(n20648), .ZN(n13449) );
  OR2_X1 U16891 ( .A1(n20757), .A2(n10261), .ZN(n13450) );
  INV_X1 U16892 ( .A(n19969), .ZN(n19955) );
  AND2_X1 U16893 ( .A1(n13451), .A2(n20515), .ZN(n15827) );
  NAND2_X1 U16894 ( .A1(n19924), .A2(n14187), .ZN(n15886) );
  AOI22_X1 U16895 ( .A1(n20027), .A2(n19955), .B1(P1_REIP_REG_0__SCAN_IN), 
        .B2(n15886), .ZN(n13462) );
  INV_X1 U16896 ( .A(n13452), .ZN(n13453) );
  NOR2_X1 U16897 ( .A1(n15827), .A2(n13453), .ZN(n13454) );
  NAND2_X1 U16898 ( .A1(n13455), .A2(n13454), .ZN(n15924) );
  OR2_X1 U16899 ( .A1(n20757), .A2(n13456), .ZN(n19965) );
  AND2_X1 U16900 ( .A1(n13457), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13458) );
  OAI21_X1 U16901 ( .B1(n19962), .B2(n19961), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13459) );
  OAI21_X1 U16902 ( .B1(n19965), .B2(n20735), .A(n13459), .ZN(n13460) );
  AOI21_X1 U16903 ( .B1(P1_EBX_REG_0__SCAN_IN), .B2(n19967), .A(n13460), .ZN(
        n13461) );
  OAI211_X1 U16904 ( .C1(n19976), .C2(n13463), .A(n13462), .B(n13461), .ZN(
        P1_U2840) );
  AND2_X1 U16905 ( .A1(n13412), .A2(n13464), .ZN(n13466) );
  OR2_X1 U16906 ( .A1(n13466), .A2(n13465), .ZN(n19901) );
  AOI22_X1 U16907 ( .A1(n13772), .A2(n14293), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14342), .ZN(n13467) );
  OAI21_X1 U16908 ( .B1(n19901), .B2(n14285), .A(n13467), .ZN(P1_U2895) );
  INV_X1 U16909 ( .A(n13521), .ZN(n13468) );
  AOI21_X1 U16910 ( .B1(n13470), .B2(n13469), .A(n13468), .ZN(n19903) );
  AOI22_X1 U16911 ( .A1(n19903), .A2(n14223), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n14222), .ZN(n13471) );
  OAI21_X1 U16912 ( .B1(n19901), .B2(n14254), .A(n13471), .ZN(P1_U2863) );
  INV_X1 U16913 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20672) );
  NAND4_X1 U16914 ( .A1(n19972), .A2(P1_REIP_REG_1__SCAN_IN), .A3(
        P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n19952) );
  NOR2_X1 U16915 ( .A1(n20672), .A2(n19952), .ZN(n19935) );
  INV_X1 U16916 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20674) );
  AND4_X1 U16917 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_4__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n13534)
         );
  OAI21_X1 U16918 ( .B1(n19924), .B2(n13534), .A(n14187), .ZN(n19953) );
  AOI21_X1 U16919 ( .B1(n19962), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n10704), .ZN(n13473) );
  AOI22_X1 U16920 ( .A1(n19967), .A2(P1_EBX_REG_5__SCAN_IN), .B1(n19948), .B2(
        n16103), .ZN(n13472) );
  OAI211_X1 U16921 ( .C1(n16008), .C2(n19950), .A(n13473), .B(n13472), .ZN(
        n13474) );
  AOI221_X1 U16922 ( .B1(n19935), .B2(n20674), .C1(n19953), .C2(
        P1_REIP_REG_5__SCAN_IN), .A(n13474), .ZN(n13475) );
  OAI21_X1 U16923 ( .B1(n19969), .B2(n16003), .A(n13475), .ZN(P1_U2835) );
  AOI21_X1 U16924 ( .B1(n13478), .B2(n13477), .A(n13476), .ZN(n13482) );
  XNOR2_X1 U16925 ( .A(n13480), .B(n13479), .ZN(n13577) );
  INV_X1 U16926 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13591) );
  XNOR2_X1 U16927 ( .A(n13577), .B(n13591), .ZN(n13481) );
  XNOR2_X1 U16928 ( .A(n13482), .B(n13481), .ZN(n19125) );
  INV_X1 U16929 ( .A(n19125), .ZN(n13505) );
  NAND2_X1 U16930 ( .A1(n13484), .A2(n13483), .ZN(n13487) );
  NAND2_X1 U16931 ( .A1(n13485), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13486) );
  NAND2_X1 U16932 ( .A1(n13487), .A2(n13486), .ZN(n13495) );
  INV_X1 U16933 ( .A(n13495), .ZN(n13493) );
  XNOR2_X1 U16934 ( .A(n13543), .B(n13491), .ZN(n13494) );
  INV_X1 U16935 ( .A(n13494), .ZN(n13492) );
  NAND2_X1 U16936 ( .A1(n13495), .A2(n13494), .ZN(n13584) );
  NAND2_X1 U16937 ( .A1(n13585), .A2(n13584), .ZN(n13496) );
  XNOR2_X1 U16938 ( .A(n13496), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19122) );
  NAND2_X1 U16939 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13954), .ZN(
        n13590) );
  OR2_X1 U16940 ( .A1(n19143), .A2(n15466), .ZN(n19153) );
  AOI21_X1 U16941 ( .B1(n13363), .B2(n19153), .A(n13701), .ZN(n13598) );
  NAND2_X1 U16942 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19119), .ZN(n13497) );
  OAI221_X1 U16943 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n13590), .C1(
        n13591), .C2(n13598), .A(n13497), .ZN(n13503) );
  NAND2_X1 U16944 ( .A1(n13499), .A2(n13498), .ZN(n13501) );
  INV_X1 U16945 ( .A(n13593), .ZN(n13500) );
  NAND2_X1 U16946 ( .A1(n13501), .A2(n13500), .ZN(n19025) );
  OAI22_X1 U16947 ( .A1(n18964), .A2(n16248), .B1(n19136), .B2(n19025), .ZN(
        n13502) );
  AOI211_X1 U16948 ( .C1(n19122), .C2(n16228), .A(n13503), .B(n13502), .ZN(
        n13504) );
  OAI21_X1 U16949 ( .B1(n13505), .B2(n19166), .A(n13504), .ZN(P2_U3042) );
  INV_X1 U16950 ( .A(n19965), .ZN(n14198) );
  OAI221_X1 U16951 ( .B1(n19924), .B2(P1_REIP_REG_1__SCAN_IN), .C1(n19924), 
        .C2(P1_REIP_REG_2__SCAN_IN), .A(n14187), .ZN(n13506) );
  AOI22_X1 U16952 ( .A1(n19962), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n13506), .ZN(n13507) );
  OAI21_X1 U16953 ( .B1(n19950), .B2(n13508), .A(n13507), .ZN(n13509) );
  AOI21_X1 U16954 ( .B1(n19967), .B2(P1_EBX_REG_3__SCAN_IN), .A(n13509), .ZN(
        n13511) );
  NAND4_X1 U16955 ( .A1(n19972), .A2(P1_REIP_REG_2__SCAN_IN), .A3(n13162), 
        .A4(P1_REIP_REG_1__SCAN_IN), .ZN(n13510) );
  OAI211_X1 U16956 ( .C1(n13512), .C2(n19976), .A(n13511), .B(n13510), .ZN(
        n13513) );
  AOI21_X1 U16957 ( .B1(n14198), .B2(n12956), .A(n13513), .ZN(n13514) );
  OAI21_X1 U16958 ( .B1(n13515), .B2(n19969), .A(n13514), .ZN(P1_U2837) );
  INV_X1 U16959 ( .A(n13516), .ZN(n13519) );
  INV_X1 U16960 ( .A(n13465), .ZN(n13518) );
  AOI21_X1 U16961 ( .B1(n13519), .B2(n13518), .A(n13517), .ZN(n14483) );
  INV_X1 U16962 ( .A(n14483), .ZN(n13541) );
  AND2_X1 U16963 ( .A1(n13521), .A2(n13520), .ZN(n13522) );
  OR2_X1 U16964 ( .A1(n13522), .A2(n13735), .ZN(n16069) );
  OAI22_X1 U16965 ( .A1(n16069), .A2(n14259), .B1(n20911), .B2(n14260), .ZN(
        n13523) );
  INV_X1 U16966 ( .A(n13523), .ZN(n13524) );
  OAI21_X1 U16967 ( .B1(n13541), .B2(n14254), .A(n13524), .ZN(P1_U2862) );
  AOI22_X1 U16968 ( .A1(n13772), .A2(n14288), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n14342), .ZN(n13525) );
  OAI21_X1 U16969 ( .B1(n13541), .B2(n14285), .A(n13525), .ZN(P1_U2894) );
  AND2_X1 U16970 ( .A1(n13527), .A2(n13526), .ZN(n13528) );
  NOR2_X1 U16971 ( .A1(n13628), .A2(n13528), .ZN(n18859) );
  NOR2_X1 U16972 ( .A1(n14743), .A2(n11879), .ZN(n13532) );
  AOI211_X1 U16973 ( .C1(n13530), .C2(n13529), .A(n15060), .B(n13625), .ZN(
        n13531) );
  AOI211_X1 U16974 ( .C1(n18859), .C2(n14743), .A(n13532), .B(n13531), .ZN(
        n13533) );
  INV_X1 U16975 ( .A(n13533), .ZN(P2_U2872) );
  INV_X1 U16976 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20678) );
  NAND3_X1 U16977 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .A3(n13534), .ZN(n19923) );
  NOR2_X1 U16978 ( .A1(n20678), .A2(n19923), .ZN(n19915) );
  NAND2_X1 U16979 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n19915), .ZN(n19913) );
  NAND2_X1 U16980 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n13758) );
  NOR2_X1 U16981 ( .A1(n19913), .A2(n13758), .ZN(n14044) );
  NAND2_X1 U16982 ( .A1(n14044), .A2(n14187), .ZN(n15887) );
  AND2_X1 U16983 ( .A1(n15886), .A2(n15887), .ZN(n15942) );
  NOR2_X1 U16984 ( .A1(n19924), .A2(n19913), .ZN(n19902) );
  NAND2_X1 U16985 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n19902), .ZN(n13536) );
  AOI22_X1 U16986 ( .A1(n19967), .A2(P1_EBX_REG_10__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19962), .ZN(n13535) );
  OAI21_X1 U16987 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(n13536), .A(n13535), 
        .ZN(n13537) );
  AOI211_X1 U16988 ( .C1(P1_REIP_REG_10__SCAN_IN), .C2(n15942), .A(n10704), 
        .B(n13537), .ZN(n13540) );
  OAI22_X1 U16989 ( .A1(n16069), .A2(n19976), .B1(n14481), .B2(n19950), .ZN(
        n13538) );
  INV_X1 U16990 ( .A(n13538), .ZN(n13539) );
  OAI211_X1 U16991 ( .C1(n13541), .C2(n19928), .A(n13540), .B(n13539), .ZN(
        P1_U2830) );
  INV_X1 U16992 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13549) );
  INV_X1 U16993 ( .A(n13544), .ZN(n13548) );
  AOI22_X1 U16994 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n13545), .B1(
        n19453), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13547) );
  AOI22_X1 U16995 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n13296), .B1(
        n13291), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13546) );
  OAI211_X1 U16996 ( .C1(n13549), .C2(n13548), .A(n13547), .B(n13546), .ZN(
        n13550) );
  INV_X1 U16997 ( .A(n13550), .ZN(n13562) );
  AOI22_X1 U16998 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19422), .B1(
        n13669), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13558) );
  INV_X1 U16999 ( .A(n13287), .ZN(n13553) );
  INV_X1 U17000 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13552) );
  INV_X1 U17001 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13551) );
  INV_X1 U17002 ( .A(n13554), .ZN(n13557) );
  NAND2_X1 U17003 ( .A1(n19335), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n13556) );
  AOI22_X1 U17004 ( .A1(n19388), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n19569), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13555) );
  AOI22_X1 U17005 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n15651), .B1(
        n15629), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13560) );
  AOI22_X1 U17006 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19197), .B1(
        n13674), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13559) );
  NAND4_X1 U17007 ( .A1(n13562), .A2(n13561), .A3(n13560), .A4(n13559), .ZN(
        n13565) );
  NAND2_X1 U17008 ( .A1(n13563), .A2(n11798), .ZN(n13564) );
  INV_X1 U17009 ( .A(n13566), .ZN(n13567) );
  NAND2_X1 U17010 ( .A1(n13568), .A2(n13567), .ZN(n13569) );
  OAI21_X1 U17011 ( .B1(n13572), .B2(n13571), .A(n13570), .ZN(n18942) );
  INV_X1 U17012 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13597) );
  NAND2_X1 U17013 ( .A1(n13577), .A2(n13591), .ZN(n13576) );
  OAI21_X1 U17014 ( .B1(n13579), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n13576), .ZN(n13573) );
  INV_X1 U17015 ( .A(n13573), .ZN(n13574) );
  NAND2_X1 U17016 ( .A1(n13575), .A2(n13574), .ZN(n13581) );
  AND2_X1 U17017 ( .A1(n13576), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13578) );
  INV_X1 U17018 ( .A(n13577), .ZN(n18959) );
  AOI22_X1 U17019 ( .A1(n13579), .A2(n13578), .B1(n18959), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13580) );
  NAND2_X1 U17020 ( .A1(n13581), .A2(n13580), .ZN(n13693) );
  XNOR2_X1 U17021 ( .A(n13694), .B(n13693), .ZN(n13603) );
  INV_X1 U17022 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n13582) );
  NOR2_X1 U17023 ( .A1(n18921), .A2(n13582), .ZN(n13592) );
  INV_X1 U17024 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18956) );
  OAI22_X1 U17025 ( .A1(n19129), .A2(n18956), .B1(n16190), .B2(n18947), .ZN(
        n13583) );
  AOI211_X1 U17026 ( .C1(n19121), .C2(n18948), .A(n13592), .B(n13583), .ZN(
        n13589) );
  AND2_X1 U17027 ( .A1(n13586), .A2(n13597), .ZN(n13658) );
  NOR2_X1 U17028 ( .A1(n13686), .A2(n13658), .ZN(n13587) );
  XNOR2_X1 U17029 ( .A(n13659), .B(n13587), .ZN(n13601) );
  NAND2_X1 U17030 ( .A1(n13601), .A2(n19123), .ZN(n13588) );
  OAI211_X1 U17031 ( .C1(n13603), .C2(n16192), .A(n13589), .B(n13588), .ZN(
        P2_U3009) );
  AOI221_X1 U17032 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n13597), .C2(n13591), .A(
        n13590), .ZN(n13600) );
  AOI21_X1 U17033 ( .B1(n19156), .B2(n18948), .A(n13592), .ZN(n13596) );
  XNOR2_X1 U17034 ( .A(n13594), .B(n13593), .ZN(n19023) );
  OR2_X1 U17035 ( .A1(n19136), .A2(n19023), .ZN(n13595) );
  OAI211_X1 U17036 ( .C1(n13598), .C2(n13597), .A(n13596), .B(n13595), .ZN(
        n13599) );
  AOI211_X1 U17037 ( .C1(n13601), .C2(n16228), .A(n13600), .B(n13599), .ZN(
        n13602) );
  OAI21_X1 U17038 ( .B1(n19166), .B2(n13603), .A(n13602), .ZN(P2_U3041) );
  XNOR2_X1 U17039 ( .A(n13604), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13605) );
  XNOR2_X1 U17040 ( .A(n13606), .B(n13605), .ZN(n16090) );
  INV_X1 U17041 ( .A(n16090), .ZN(n13610) );
  AOI22_X1 U17042 ( .A1(n20013), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n10704), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13607) );
  OAI21_X1 U17043 ( .B1(n20023), .B2(n19911), .A(n13607), .ZN(n13608) );
  AOI21_X1 U17044 ( .B1(n19919), .B2(n14447), .A(n13608), .ZN(n13609) );
  OAI21_X1 U17045 ( .B1(n13610), .B2(n20030), .A(n13609), .ZN(P1_U2991) );
  AOI22_X1 U17046 ( .A1(n12053), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12144), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13617) );
  NAND2_X1 U17047 ( .A1(n12004), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n13613) );
  NAND2_X1 U17048 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n13612) );
  NAND2_X1 U17049 ( .A1(n11963), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13611) );
  AND3_X1 U17050 ( .A1(n13613), .A2(n13612), .A3(n13611), .ZN(n13616) );
  AOI22_X1 U17051 ( .A1(n14862), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14861), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13615) );
  AOI22_X1 U17052 ( .A1(n12056), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12057), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13614) );
  NAND4_X1 U17053 ( .A1(n13617), .A2(n13616), .A3(n13615), .A4(n13614), .ZN(
        n13623) );
  AOI22_X1 U17054 ( .A1(n14867), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13621) );
  AOI22_X1 U17055 ( .A1(n12026), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12027), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13620) );
  AOI22_X1 U17056 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13619) );
  NAND2_X1 U17057 ( .A1(n14868), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n13618) );
  NAND4_X1 U17058 ( .A1(n13621), .A2(n13620), .A3(n13619), .A4(n13618), .ZN(
        n13622) );
  OR2_X1 U17059 ( .A1(n13623), .A2(n13622), .ZN(n13624) );
  NOR2_X1 U17060 ( .A1(n13625), .A2(n13624), .ZN(n13626) );
  OR2_X1 U17061 ( .A1(n13646), .A2(n13626), .ZN(n18985) );
  XOR2_X1 U17062 ( .A(n13628), .B(n13627), .Z(n18849) );
  INV_X1 U17063 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n13629) );
  NOR2_X1 U17064 ( .A1(n14743), .A2(n13629), .ZN(n13630) );
  AOI21_X1 U17065 ( .B1(n18849), .B2(n14743), .A(n13630), .ZN(n13631) );
  OAI21_X1 U17066 ( .B1(n18985), .B2(n15060), .A(n13631), .ZN(P2_U2871) );
  AOI22_X1 U17067 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n12144), .B1(
        n12053), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13638) );
  NAND2_X1 U17068 ( .A1(n12004), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13634) );
  NAND2_X1 U17069 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n13633) );
  NAND2_X1 U17070 ( .A1(n11963), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13632) );
  AND3_X1 U17071 ( .A1(n13634), .A2(n13633), .A3(n13632), .ZN(n13637) );
  AOI22_X1 U17072 ( .A1(n14862), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14861), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13636) );
  AOI22_X1 U17073 ( .A1(n12056), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12057), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13635) );
  NAND4_X1 U17074 ( .A1(n13638), .A2(n13637), .A3(n13636), .A4(n13635), .ZN(
        n13644) );
  AOI22_X1 U17075 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n14867), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13642) );
  AOI22_X1 U17076 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12026), .B1(
        n12027), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13641) );
  AOI22_X1 U17077 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12003), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13640) );
  NAND2_X1 U17078 ( .A1(n14868), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n13639) );
  NAND4_X1 U17079 ( .A1(n13642), .A2(n13641), .A3(n13640), .A4(n13639), .ZN(
        n13643) );
  OR2_X1 U17080 ( .A1(n13644), .A2(n13643), .ZN(n13645) );
  OAI21_X1 U17081 ( .B1(n13646), .B2(n13645), .A(n13726), .ZN(n15135) );
  NAND2_X1 U17082 ( .A1(n15050), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13651) );
  INV_X1 U17083 ( .A(n13711), .ZN(n13647) );
  AOI21_X1 U17084 ( .B1(n13649), .B2(n13648), .A(n13647), .ZN(n18838) );
  NAND2_X1 U17085 ( .A1(n18838), .A2(n14743), .ZN(n13650) );
  OAI211_X1 U17086 ( .C1(n15135), .C2(n15060), .A(n13651), .B(n13650), .ZN(
        P2_U2870) );
  XNOR2_X1 U17087 ( .A(n9611), .B(n16081), .ZN(n13652) );
  XNOR2_X1 U17088 ( .A(n13653), .B(n13652), .ZN(n16078) );
  NAND2_X1 U17089 ( .A1(n16078), .A2(n20019), .ZN(n13657) );
  INV_X1 U17090 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n13654) );
  OAI22_X1 U17091 ( .A1(n20024), .A2(n19906), .B1(n20036), .B2(n13654), .ZN(
        n13655) );
  AOI21_X1 U17092 ( .B1(n15976), .B2(n19900), .A(n13655), .ZN(n13656) );
  OAI211_X1 U17093 ( .C1(n15947), .C2(n19901), .A(n13657), .B(n13656), .ZN(
        P1_U2990) );
  NAND2_X1 U17094 ( .A1(n15651), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n13663) );
  AOI22_X1 U17095 ( .A1(n13660), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n19453), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13662) );
  AOI22_X1 U17096 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n13545), .B1(
        n19569), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13661) );
  AOI22_X1 U17097 ( .A1(n13287), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13291), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13673) );
  INV_X1 U17098 ( .A(n19422), .ZN(n13667) );
  INV_X1 U17099 ( .A(n19388), .ZN(n13665) );
  OAI22_X1 U17100 ( .A1(n13667), .A2(n13666), .B1(n13665), .B2(n13664), .ZN(
        n13668) );
  INV_X1 U17101 ( .A(n13668), .ZN(n13672) );
  NAND2_X1 U17102 ( .A1(n19335), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n13671) );
  AOI22_X1 U17103 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n13669), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13670) );
  AOI22_X1 U17104 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19197), .B1(
        n13674), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13676) );
  AOI22_X1 U17105 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n15629), .B1(
        n13544), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13675) );
  NAND4_X1 U17106 ( .A1(n13678), .A2(n13677), .A3(n13676), .A4(n13675), .ZN(
        n13681) );
  NAND2_X1 U17107 ( .A1(n13679), .A2(n11798), .ZN(n13680) );
  NAND2_X1 U17108 ( .A1(n13935), .A2(n13684), .ZN(n13691) );
  NAND2_X1 U17109 ( .A1(n13699), .A2(n13936), .ZN(n13688) );
  NAND2_X1 U17110 ( .A1(n13686), .A2(n13685), .ZN(n13687) );
  OAI21_X1 U17111 ( .B1(n13692), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n13940), .ZN(n16214) );
  NAND2_X1 U17112 ( .A1(n13695), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13696) );
  NAND2_X1 U17113 ( .A1(n13697), .A2(n13696), .ZN(n13820) );
  INV_X1 U17114 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13953) );
  XNOR2_X1 U17115 ( .A(n13821), .B(n13953), .ZN(n13819) );
  XOR2_X1 U17116 ( .A(n13820), .B(n13819), .Z(n16216) );
  NAND3_X1 U17117 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13952) );
  AOI21_X1 U17118 ( .B1(n13952), .B2(n19153), .A(n13701), .ZN(n13707) );
  INV_X1 U17119 ( .A(n13954), .ZN(n13702) );
  NOR3_X1 U17120 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13702), .A3(
        n13952), .ZN(n13703) );
  AOI21_X1 U17121 ( .B1(n19119), .B2(P2_REIP_REG_6__SCAN_IN), .A(n13703), .ZN(
        n13704) );
  OAI21_X1 U17122 ( .B1(n19136), .B2(n19013), .A(n13704), .ZN(n13705) );
  AOI21_X1 U17123 ( .B1(n19156), .B2(n16215), .A(n13705), .ZN(n13706) );
  OAI21_X1 U17124 ( .B1(n13707), .B2(n13953), .A(n13706), .ZN(n13708) );
  AOI21_X1 U17125 ( .B1(n16216), .B2(n19131), .A(n13708), .ZN(n13709) );
  OAI21_X1 U17126 ( .B1(n19159), .B2(n16214), .A(n13709), .ZN(P2_U3040) );
  NAND2_X1 U17127 ( .A1(n13711), .A2(n13710), .ZN(n13712) );
  NAND2_X1 U17128 ( .A1(n15056), .A2(n13712), .ZN(n18825) );
  AOI22_X1 U17129 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n12144), .B1(
        n12053), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13719) );
  NAND2_X1 U17130 ( .A1(n12004), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n13715) );
  NAND2_X1 U17131 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n13714) );
  NAND2_X1 U17132 ( .A1(n11963), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13713) );
  AND3_X1 U17133 ( .A1(n13715), .A2(n13714), .A3(n13713), .ZN(n13718) );
  AOI22_X1 U17134 ( .A1(n14862), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14861), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13717) );
  AOI22_X1 U17135 ( .A1(n12056), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12057), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13716) );
  NAND4_X1 U17136 ( .A1(n13719), .A2(n13718), .A3(n13717), .A4(n13716), .ZN(
        n13725) );
  AOI22_X1 U17137 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n14867), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13723) );
  AOI22_X1 U17138 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n12026), .B1(
        n12027), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13722) );
  AOI22_X1 U17139 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12003), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13721) );
  NAND2_X1 U17140 ( .A1(n14868), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n13720) );
  NAND4_X1 U17141 ( .A1(n13723), .A2(n13722), .A3(n13721), .A4(n13720), .ZN(
        n13724) );
  NOR2_X1 U17142 ( .A1(n13725), .A2(n13724), .ZN(n13729) );
  INV_X1 U17143 ( .A(n14830), .ZN(n15054) );
  AOI21_X1 U17144 ( .B1(n13729), .B2(n13726), .A(n15054), .ZN(n16153) );
  NAND2_X1 U17145 ( .A1(n16153), .A2(n15047), .ZN(n13731) );
  NAND2_X1 U17146 ( .A1(n15055), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n13730) );
  OAI211_X1 U17147 ( .C1(n18825), .C2(n15050), .A(n13731), .B(n13730), .ZN(
        P2_U2869) );
  OAI21_X1 U17148 ( .B1(n13517), .B2(n13733), .A(n13732), .ZN(n13750) );
  XNOR2_X1 U17149 ( .A(n13750), .B(n13748), .ZN(n15984) );
  INV_X1 U17150 ( .A(n15984), .ZN(n13737) );
  AOI22_X1 U17151 ( .A1(n13772), .A2(n14280), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n14342), .ZN(n13734) );
  OAI21_X1 U17152 ( .B1(n13737), .B2(n14285), .A(n13734), .ZN(P1_U2893) );
  INV_X1 U17153 ( .A(n13797), .ZN(n13753) );
  OAI21_X1 U17154 ( .B1(n13736), .B2(n13735), .A(n13753), .ZN(n15939) );
  INV_X1 U17155 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n13738) );
  OAI222_X1 U17156 ( .A1(n15939), .A2(n14259), .B1(n13738), .B2(n14260), .C1(
        n13737), .C2(n14254), .ZN(P1_U2861) );
  INV_X1 U17157 ( .A(n13740), .ZN(n13741) );
  AOI21_X1 U17158 ( .B1(n13742), .B2(n13739), .A(n13741), .ZN(n15928) );
  INV_X1 U17159 ( .A(n15928), .ZN(n13747) );
  AOI22_X1 U17160 ( .A1(n13772), .A2(n14264), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14342), .ZN(n13743) );
  OAI21_X1 U17161 ( .B1(n13747), .B2(n14285), .A(n13743), .ZN(P1_U2890) );
  INV_X1 U17162 ( .A(n13804), .ZN(n13744) );
  AOI21_X1 U17163 ( .B1(n13745), .B2(n13754), .A(n13744), .ZN(n15921) );
  AOI22_X1 U17164 ( .A1(n15921), .A2(n14223), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n14222), .ZN(n13746) );
  OAI21_X1 U17165 ( .B1(n13747), .B2(n14254), .A(n13746), .ZN(P1_U2858) );
  INV_X1 U17166 ( .A(n13748), .ZN(n13749) );
  OAI21_X1 U17167 ( .B1(n13750), .B2(n13749), .A(n13732), .ZN(n13767) );
  AND2_X1 U17168 ( .A1(n13767), .A2(n13768), .ZN(n13769) );
  OAI21_X1 U17169 ( .B1(n13769), .B2(n13751), .A(n13739), .ZN(n14478) );
  OAI21_X1 U17170 ( .B1(n13753), .B2(n13795), .A(n13752), .ZN(n13755) );
  NAND2_X1 U17171 ( .A1(n13755), .A2(n13754), .ZN(n13766) );
  INV_X1 U17172 ( .A(n13766), .ZN(n16036) );
  AOI22_X1 U17173 ( .A1(n16036), .A2(n19948), .B1(n19967), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n13756) );
  OAI211_X1 U17174 ( .C1(n19905), .C2(n13757), .A(n13756), .B(n20036), .ZN(
        n13762) );
  NAND2_X1 U17175 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14180) );
  INV_X1 U17176 ( .A(n15933), .ZN(n15945) );
  NOR2_X1 U17177 ( .A1(n14180), .A2(n15945), .ZN(n13760) );
  OAI21_X1 U17178 ( .B1(n14180), .B2(n15887), .A(n15886), .ZN(n15937) );
  INV_X1 U17179 ( .A(n15937), .ZN(n13759) );
  MUX2_X1 U17180 ( .A(n13760), .B(n13759), .S(P1_REIP_REG_13__SCAN_IN), .Z(
        n13761) );
  AOI211_X1 U17181 ( .C1(n14475), .C2(n19961), .A(n13762), .B(n13761), .ZN(
        n13763) );
  OAI21_X1 U17182 ( .B1(n14478), .B2(n19928), .A(n13763), .ZN(P1_U2827) );
  AOI22_X1 U17183 ( .A1(n13772), .A2(n14269), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n14342), .ZN(n13764) );
  OAI21_X1 U17184 ( .B1(n14478), .B2(n14285), .A(n13764), .ZN(P1_U2891) );
  INV_X1 U17185 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n13765) );
  OAI222_X1 U17186 ( .A1(n13766), .A2(n14259), .B1(n13765), .B2(n14260), .C1(
        n14478), .C2(n14254), .ZN(P1_U2859) );
  INV_X1 U17187 ( .A(n13767), .ZN(n13771) );
  INV_X1 U17188 ( .A(n13768), .ZN(n13770) );
  AOI21_X1 U17189 ( .B1(n13771), .B2(n13770), .A(n13769), .ZN(n15974) );
  INV_X1 U17190 ( .A(n15974), .ZN(n13799) );
  AOI22_X1 U17191 ( .A1(n13772), .A2(n14275), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n14342), .ZN(n13773) );
  OAI21_X1 U17192 ( .B1(n13799), .B2(n14285), .A(n13773), .ZN(P1_U2892) );
  INV_X1 U17193 ( .A(n13775), .ZN(n13776) );
  NAND2_X1 U17194 ( .A1(n13774), .A2(n13776), .ZN(n14456) );
  INV_X1 U17195 ( .A(n13777), .ZN(n13778) );
  AOI21_X1 U17196 ( .B1(n14456), .B2(n13779), .A(n13778), .ZN(n13781) );
  XNOR2_X1 U17197 ( .A(n9611), .B(n14610), .ZN(n13780) );
  XNOR2_X1 U17198 ( .A(n13781), .B(n13780), .ZN(n13794) );
  INV_X1 U17199 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n13782) );
  NOR2_X1 U17200 ( .A1(n20036), .A2(n13782), .ZN(n13789) );
  INV_X1 U17201 ( .A(n20066), .ZN(n16085) );
  OAI21_X1 U17202 ( .B1(n16085), .B2(n20054), .A(n20056), .ZN(n16053) );
  NAND2_X1 U17203 ( .A1(n16053), .A2(n14610), .ZN(n13785) );
  OAI21_X1 U17204 ( .B1(n20034), .B2(n13783), .A(n20033), .ZN(n13784) );
  AOI21_X1 U17205 ( .B1(n16046), .B2(n13786), .A(n13784), .ZN(n16037) );
  OAI22_X1 U17206 ( .A1(n13786), .A2(n13785), .B1(n16037), .B2(n14610), .ZN(
        n13787) );
  AOI211_X1 U17207 ( .C1(n20059), .C2(n15921), .A(n13789), .B(n13787), .ZN(
        n13788) );
  OAI21_X1 U17208 ( .B1(n13794), .B2(n16106), .A(n13788), .ZN(P1_U3017) );
  AOI21_X1 U17209 ( .B1(n20013), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n13789), .ZN(n13790) );
  OAI21_X1 U17210 ( .B1(n20023), .B2(n13791), .A(n13790), .ZN(n13792) );
  AOI21_X1 U17211 ( .B1(n15928), .B2(n14447), .A(n13792), .ZN(n13793) );
  OAI21_X1 U17212 ( .B1(n13794), .B2(n20030), .A(n13793), .ZN(P1_U2985) );
  INV_X1 U17213 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n13798) );
  INV_X1 U17214 ( .A(n13795), .ZN(n13796) );
  XNOR2_X1 U17215 ( .A(n13797), .B(n13796), .ZN(n16049) );
  OAI222_X1 U17216 ( .A1(n14254), .A2(n13799), .B1(n13798), .B2(n14260), .C1(
        n14259), .C2(n16049), .ZN(P1_U2860) );
  INV_X1 U17217 ( .A(n13800), .ZN(n13801) );
  AOI21_X1 U17218 ( .B1(n13802), .B2(n13740), .A(n13801), .ZN(n15967) );
  INV_X1 U17219 ( .A(n15967), .ZN(n13809) );
  AND2_X1 U17220 ( .A1(n13804), .A2(n13803), .ZN(n13805) );
  NOR2_X1 U17221 ( .A1(n9694), .A2(n13805), .ZN(n16031) );
  AOI22_X1 U17222 ( .A1(n16031), .A2(n14223), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n14222), .ZN(n13806) );
  OAI21_X1 U17223 ( .B1(n13809), .B2(n14254), .A(n13806), .ZN(P1_U2857) );
  OAI222_X1 U17224 ( .A1(n14285), .A2(n13809), .B1(n14353), .B2(n13808), .C1(
        n14352), .C2(n13807), .ZN(P1_U2889) );
  OR2_X1 U17225 ( .A1(n9610), .A2(n13810), .ZN(n18550) );
  INV_X1 U17226 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18540) );
  NAND3_X1 U17227 ( .A1(n16940), .A2(n18550), .A3(n18540), .ZN(n18090) );
  NOR2_X1 U17228 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18090), .ZN(n13811) );
  NAND3_X1 U17229 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18703)
         );
  OAI21_X1 U17230 ( .B1(n13811), .B2(n18703), .A(n18142), .ZN(n18096) );
  INV_X1 U17231 ( .A(n18096), .ZN(n13812) );
  INV_X1 U17232 ( .A(n17671), .ZN(n17726) );
  NOR2_X1 U17233 ( .A1(n18744), .A2(n17726), .ZN(n15756) );
  AOI21_X1 U17234 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n15756), .ZN(n15757) );
  NOR2_X1 U17235 ( .A1(n13812), .A2(n15757), .ZN(n13814) );
  NOR2_X1 U17236 ( .A1(n20828), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18141) );
  OR2_X1 U17237 ( .A1(n18141), .A2(n13812), .ZN(n15755) );
  OR2_X1 U17238 ( .A1(n18445), .A2(n15755), .ZN(n13813) );
  MUX2_X1 U17239 ( .A(n13814), .B(n13813), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  INV_X1 U17240 ( .A(n13815), .ZN(n13816) );
  NAND2_X1 U17241 ( .A1(n13816), .A2(n9658), .ZN(n13817) );
  NAND2_X1 U17242 ( .A1(n14704), .A2(n13698), .ZN(n13978) );
  NAND2_X1 U17243 ( .A1(n13821), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13822) );
  NOR2_X1 U17244 ( .A1(n13823), .A2(n13905), .ZN(n13829) );
  NAND2_X1 U17245 ( .A1(n13829), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15548) );
  AND2_X1 U17246 ( .A1(n19177), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n13825) );
  MUX2_X1 U17247 ( .A(n13826), .B(n13825), .S(n13824), .Z(n13827) );
  NOR2_X1 U17248 ( .A1(n13827), .A2(n13833), .ZN(n18929) );
  NAND2_X1 U17249 ( .A1(n18929), .A2(n13929), .ZN(n13828) );
  INV_X1 U17250 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n13994) );
  NAND2_X1 U17251 ( .A1(n13828), .A2(n13994), .ZN(n13990) );
  INV_X1 U17252 ( .A(n13829), .ZN(n13830) );
  INV_X1 U17253 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15555) );
  NAND2_X1 U17254 ( .A1(n13830), .A2(n15555), .ZN(n15547) );
  INV_X1 U17255 ( .A(n13831), .ZN(n13832) );
  INV_X1 U17256 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n13943) );
  NAND2_X1 U17257 ( .A1(n13832), .A2(n13943), .ZN(n15287) );
  AND2_X1 U17258 ( .A1(n15547), .A2(n15287), .ZN(n13988) );
  NAND2_X1 U17259 ( .A1(n13833), .A2(n18918), .ZN(n13837) );
  NOR2_X1 U17260 ( .A1(n13833), .A2(n18918), .ZN(n13834) );
  NAND2_X1 U17261 ( .A1(n13916), .A2(n13834), .ZN(n13835) );
  AND2_X1 U17262 ( .A1(n13917), .A2(n13835), .ZN(n13836) );
  NAND2_X1 U17263 ( .A1(n13837), .A2(n13836), .ZN(n18919) );
  OR2_X1 U17264 ( .A1(n18919), .A2(n13905), .ZN(n13838) );
  INV_X1 U17265 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15527) );
  NAND2_X1 U17266 ( .A1(n13838), .A2(n15527), .ZN(n15534) );
  OR2_X1 U17267 ( .A1(n13840), .A2(n10109), .ZN(n18905) );
  INV_X1 U17268 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13841) );
  OAI21_X1 U17269 ( .B1(n18905), .B2(n13905), .A(n13841), .ZN(n15513) );
  AND4_X1 U17270 ( .A1(n13990), .A2(n13988), .A3(n15534), .A4(n15513), .ZN(
        n13842) );
  AND2_X1 U17271 ( .A1(n13929), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13843) );
  NAND2_X1 U17272 ( .A1(n18929), .A2(n13843), .ZN(n13991) );
  OR3_X1 U17273 ( .A1(n18919), .A2(n13905), .A3(n15527), .ZN(n15533) );
  NAND2_X1 U17274 ( .A1(n13991), .A2(n15533), .ZN(n15511) );
  NAND2_X1 U17275 ( .A1(n13929), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13844) );
  NOR2_X1 U17276 ( .A1(n18905), .A2(n13844), .ZN(n15512) );
  NOR2_X1 U17277 ( .A1(n15511), .A2(n15512), .ZN(n13845) );
  NAND2_X1 U17278 ( .A1(n9878), .A2(n13847), .ZN(n13848) );
  NAND2_X1 U17279 ( .A1(n13853), .A2(n13848), .ZN(n18890) );
  OR2_X1 U17280 ( .A1(n18890), .A2(n13905), .ZN(n15492) );
  INV_X1 U17281 ( .A(n15491), .ZN(n13851) );
  INV_X1 U17282 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n13850) );
  NAND2_X1 U17283 ( .A1(n13853), .A2(n13852), .ZN(n13854) );
  AND2_X1 U17284 ( .A1(n13875), .A2(n13854), .ZN(n18874) );
  AOI21_X1 U17285 ( .B1(n18874), .B2(n13929), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15276) );
  INV_X1 U17286 ( .A(n15276), .ZN(n13855) );
  NAND2_X1 U17287 ( .A1(n13916), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n13857) );
  MUX2_X1 U17288 ( .A(n13857), .B(n19177), .S(n13856), .Z(n13859) );
  NAND2_X1 U17289 ( .A1(n13859), .A2(n13858), .ZN(n18802) );
  OAI21_X1 U17290 ( .B1(n18802), .B2(n13905), .A(n15419), .ZN(n15215) );
  XNOR2_X1 U17291 ( .A(n9649), .B(n12309), .ZN(n18811) );
  NAND2_X1 U17292 ( .A1(n18811), .A2(n13929), .ZN(n13885) );
  INV_X1 U17293 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15418) );
  NAND2_X1 U17294 ( .A1(n13885), .A2(n15418), .ZN(n15226) );
  NAND2_X1 U17295 ( .A1(n13872), .A2(n13861), .ZN(n13862) );
  NAND2_X1 U17296 ( .A1(n9649), .A2(n13862), .ZN(n18821) );
  INV_X1 U17297 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15447) );
  OAI21_X1 U17298 ( .B1(n18821), .B2(n13905), .A(n15447), .ZN(n15238) );
  AND2_X1 U17299 ( .A1(n15226), .A2(n15238), .ZN(n15212) );
  AND2_X1 U17300 ( .A1(n15215), .A2(n15212), .ZN(n15200) );
  AND2_X1 U17301 ( .A1(n19177), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n13863) );
  AOI21_X1 U17302 ( .B1(n13864), .B2(n13863), .A(n13918), .ZN(n13866) );
  AND2_X1 U17303 ( .A1(n13866), .A2(n13865), .ZN(n18845) );
  NAND2_X1 U17304 ( .A1(n18845), .A2(n13929), .ZN(n13867) );
  NAND2_X1 U17305 ( .A1(n13867), .A2(n15786), .ZN(n13868) );
  OR2_X1 U17306 ( .A1(n13870), .A2(n13869), .ZN(n13871) );
  NAND2_X1 U17307 ( .A1(n13872), .A2(n13871), .ZN(n18835) );
  INV_X1 U17308 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15461) );
  OAI21_X1 U17309 ( .B1(n18835), .B2(n13905), .A(n15461), .ZN(n15250) );
  INV_X1 U17310 ( .A(n13873), .ZN(n13874) );
  XNOR2_X1 U17311 ( .A(n13875), .B(n13874), .ZN(n18866) );
  NAND2_X1 U17312 ( .A1(n18866), .A2(n13929), .ZN(n13876) );
  INV_X1 U17313 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n13949) );
  NAND2_X1 U17314 ( .A1(n13876), .A2(n13949), .ZN(n16176) );
  INV_X1 U17315 ( .A(n13877), .ZN(n13878) );
  XNOR2_X1 U17316 ( .A(n13879), .B(n13878), .ZN(n18856) );
  NAND2_X1 U17317 ( .A1(n18856), .A2(n13929), .ZN(n13880) );
  INV_X1 U17318 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16224) );
  NAND2_X1 U17319 ( .A1(n13880), .A2(n16224), .ZN(n15263) );
  AND4_X1 U17320 ( .A1(n15197), .A2(n15250), .A3(n16176), .A4(n15263), .ZN(
        n13881) );
  OAI21_X1 U17321 ( .B1(n13882), .B2(n13905), .A(n15205), .ZN(n15202) );
  INV_X1 U17322 ( .A(n13882), .ZN(n13884) );
  AND2_X1 U17323 ( .A1(n13929), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13883) );
  NAND2_X1 U17324 ( .A1(n13884), .A2(n13883), .ZN(n15201) );
  INV_X1 U17325 ( .A(n13885), .ZN(n13886) );
  NAND2_X1 U17326 ( .A1(n13886), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15227) );
  INV_X1 U17327 ( .A(n18835), .ZN(n13888) );
  AND2_X1 U17328 ( .A1(n13929), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13887) );
  NAND2_X1 U17329 ( .A1(n13888), .A2(n13887), .ZN(n15249) );
  NAND2_X1 U17330 ( .A1(n15249), .A2(n15247), .ZN(n15198) );
  AND2_X1 U17331 ( .A1(n13929), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13889) );
  NAND2_X1 U17332 ( .A1(n18856), .A2(n13889), .ZN(n15262) );
  AND2_X1 U17333 ( .A1(n13929), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13890) );
  NAND2_X1 U17334 ( .A1(n18866), .A2(n13890), .ZN(n16175) );
  AND2_X1 U17335 ( .A1(n13929), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13891) );
  NAND2_X1 U17336 ( .A1(n18874), .A2(n13891), .ZN(n15274) );
  NAND3_X1 U17337 ( .A1(n15262), .A2(n16175), .A3(n15274), .ZN(n13892) );
  NOR2_X1 U17338 ( .A1(n15198), .A2(n13892), .ZN(n13895) );
  INV_X1 U17339 ( .A(n18821), .ZN(n13894) );
  AND2_X1 U17340 ( .A1(n13929), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13893) );
  NAND2_X1 U17341 ( .A1(n13894), .A2(n13893), .ZN(n15237) );
  AND3_X1 U17342 ( .A1(n15227), .A2(n13895), .A3(n15237), .ZN(n13898) );
  INV_X1 U17343 ( .A(n18802), .ZN(n13897) );
  AND2_X1 U17344 ( .A1(n13929), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13896) );
  NAND2_X1 U17345 ( .A1(n13897), .A2(n13896), .ZN(n15214) );
  INV_X1 U17346 ( .A(n13899), .ZN(n13900) );
  NAND2_X1 U17347 ( .A1(n13902), .A2(n9870), .ZN(n13903) );
  NAND2_X1 U17348 ( .A1(n13904), .A2(n13903), .ZN(n15797) );
  OR2_X1 U17349 ( .A1(n15797), .A2(n13905), .ZN(n13906) );
  NAND2_X1 U17350 ( .A1(n13929), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13907) );
  OR2_X1 U17351 ( .A1(n15797), .A2(n13907), .ZN(n15386) );
  NAND2_X1 U17352 ( .A1(n13908), .A2(n13929), .ZN(n13909) );
  XNOR2_X1 U17353 ( .A(n13909), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15189) );
  NOR3_X1 U17354 ( .A1(n13911), .A2(n13905), .A3(n13910), .ZN(n13912) );
  NAND2_X1 U17355 ( .A1(n13914), .A2(n13917), .ZN(n16129) );
  NOR2_X1 U17356 ( .A1(n13919), .A2(n15010), .ZN(n13915) );
  NAND2_X1 U17357 ( .A1(n13916), .A2(n13915), .ZN(n13921) );
  AOI21_X1 U17358 ( .B1(n13919), .B2(n15010), .A(n13918), .ZN(n13920) );
  AOI21_X1 U17359 ( .B1(n14737), .B2(n13929), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15167) );
  XNOR2_X1 U17360 ( .A(n13923), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15159) );
  NAND2_X1 U17361 ( .A1(n13922), .A2(n13698), .ZN(n13980) );
  INV_X1 U17362 ( .A(n13923), .ZN(n13925) );
  AND2_X1 U17363 ( .A1(n13929), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13924) );
  AND2_X1 U17364 ( .A1(n14737), .A2(n13924), .ZN(n15166) );
  AOI21_X1 U17365 ( .B1(n13925), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15166), .ZN(n13975) );
  XOR2_X1 U17366 ( .A(n13927), .B(n13926), .Z(n14688) );
  INV_X1 U17367 ( .A(n14688), .ZN(n13928) );
  INV_X1 U17368 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15298) );
  OAI21_X1 U17369 ( .B1(n13928), .B2(n13905), .A(n15298), .ZN(n15137) );
  NAND2_X1 U17370 ( .A1(n15138), .A2(n15137), .ZN(n14009) );
  NAND3_X1 U17371 ( .A1(n14688), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n13698), .ZN(n15136) );
  NAND2_X1 U17372 ( .A1(n14009), .A2(n15136), .ZN(n13934) );
  INV_X1 U17373 ( .A(n14007), .ZN(n13932) );
  NOR2_X1 U17374 ( .A1(n14008), .A2(n13932), .ZN(n13933) );
  XNOR2_X1 U17375 ( .A(n13934), .B(n13933), .ZN(n13974) );
  NAND2_X1 U17376 ( .A1(n13937), .A2(n13936), .ZN(n13938) );
  NAND2_X1 U17377 ( .A1(n13938), .A2(n13699), .ZN(n13939) );
  XNOR2_X1 U17378 ( .A(n13945), .B(n13929), .ZN(n13942) );
  INV_X1 U17379 ( .A(n13942), .ZN(n13944) );
  NAND2_X1 U17380 ( .A1(n13947), .A2(n13929), .ZN(n13946) );
  NAND3_X1 U17381 ( .A1(n13947), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n13929), .ZN(n13948) );
  NAND2_X1 U17382 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16233) );
  NOR2_X1 U17383 ( .A1(n13949), .A2(n16233), .ZN(n15460) );
  NAND2_X1 U17384 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15506) );
  NOR2_X1 U17385 ( .A1(n13994), .A2(n15506), .ZN(n15475) );
  NAND2_X1 U17386 ( .A1(n15460), .A2(n15475), .ZN(n15412) );
  AND2_X1 U17387 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15462) );
  NAND2_X1 U17388 ( .A1(n15462), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15417) );
  NOR2_X1 U17389 ( .A1(n15412), .A2(n15417), .ZN(n15414) );
  INV_X1 U17390 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15349) );
  INV_X1 U17391 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15336) );
  NOR2_X1 U17392 ( .A1(n18921), .A2(n13951), .ZN(n13969) );
  AOI21_X1 U17393 ( .B1(n15066), .B2(n19155), .A(n13969), .ZN(n13965) );
  AND2_X1 U17394 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15337) );
  NAND4_X1 U17395 ( .A1(n15414), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15403) );
  NOR2_X1 U17396 ( .A1(n15205), .A2(n15403), .ZN(n15373) );
  NAND3_X1 U17397 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n15373), .ZN(n13956) );
  NAND2_X1 U17398 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15553) );
  NOR2_X1 U17399 ( .A1(n13953), .A2(n13952), .ZN(n13957) );
  NAND2_X1 U17400 ( .A1(n13957), .A2(n13954), .ZN(n15564) );
  NOR2_X1 U17401 ( .A1(n15553), .A2(n15564), .ZN(n15459) );
  INV_X1 U17402 ( .A(n15459), .ZN(n15505) );
  NOR2_X1 U17403 ( .A1(n13956), .A2(n15505), .ZN(n15365) );
  AND2_X1 U17404 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n15365), .ZN(
        n13955) );
  NAND2_X1 U17405 ( .A1(n15337), .A2(n13955), .ZN(n15308) );
  NOR2_X1 U17406 ( .A1(n15313), .A2(n15323), .ZN(n15307) );
  NAND2_X1 U17407 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15307), .ZN(
        n14026) );
  NOR2_X1 U17408 ( .A1(n15308), .A2(n14026), .ZN(n13963) );
  NAND2_X1 U17409 ( .A1(n19153), .A2(n13956), .ZN(n13960) );
  INV_X1 U17410 ( .A(n15552), .ZN(n15507) );
  NAND2_X1 U17411 ( .A1(n13958), .A2(n13957), .ZN(n15551) );
  NOR2_X1 U17412 ( .A1(n15551), .A2(n15553), .ZN(n15508) );
  OR2_X1 U17413 ( .A1(n15507), .A2(n15508), .ZN(n13993) );
  AND2_X1 U17414 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n13993), .ZN(
        n13959) );
  NAND2_X1 U17415 ( .A1(n13960), .A2(n13959), .ZN(n15364) );
  NAND2_X1 U17416 ( .A1(n15364), .A2(n15552), .ZN(n15350) );
  OAI21_X1 U17417 ( .B1(n15349), .B2(n15336), .A(n15552), .ZN(n13961) );
  NAND2_X1 U17418 ( .A1(n15350), .A2(n13961), .ZN(n15329) );
  AND2_X1 U17419 ( .A1(n19153), .A2(n14026), .ZN(n13962) );
  OR3_X1 U17420 ( .A1(n15329), .A2(n13962), .A3(n9989), .ZN(n14025) );
  OAI21_X1 U17421 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n13963), .A(
        n14025), .ZN(n13964) );
  OAI211_X1 U17422 ( .C1(n14983), .C2(n16248), .A(n13965), .B(n13964), .ZN(
        n13966) );
  AOI21_X1 U17423 ( .B1(n13972), .B2(n16228), .A(n13966), .ZN(n13967) );
  OAI21_X1 U17424 ( .B1(n13974), .B2(n19166), .A(n13967), .ZN(P2_U3016) );
  NOR2_X1 U17425 ( .A1(n16190), .A2(n14662), .ZN(n13968) );
  AOI211_X1 U17426 ( .C1(n16184), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n13969), .B(n13968), .ZN(n13970) );
  OAI21_X1 U17427 ( .B1(n14983), .B2(n16160), .A(n13970), .ZN(n13971) );
  AOI21_X1 U17428 ( .B1(n13972), .B2(n19123), .A(n13971), .ZN(n13973) );
  OAI21_X1 U17429 ( .B1(n13974), .B2(n16192), .A(n13973), .ZN(P2_U2984) );
  NAND2_X1 U17430 ( .A1(n13976), .A2(n13975), .ZN(n13977) );
  INV_X1 U17431 ( .A(n13977), .ZN(n13979) );
  XNOR2_X1 U17432 ( .A(n13977), .B(n13978), .ZN(n15150) );
  NAND2_X1 U17433 ( .A1(n15150), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15321) );
  XNOR2_X1 U17434 ( .A(n13980), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13981) );
  INV_X1 U17435 ( .A(n14994), .ZN(n15318) );
  NOR2_X1 U17436 ( .A1(n18921), .A2(n19779), .ZN(n15310) );
  AOI21_X1 U17437 ( .B1(n16184), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15310), .ZN(n13982) );
  OAI21_X1 U17438 ( .B1(n16190), .B2(n13983), .A(n13982), .ZN(n13985) );
  OAI21_X1 U17439 ( .B1(n15148), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15141), .ZN(n15315) );
  NOR2_X1 U17440 ( .A1(n15315), .A2(n16194), .ZN(n13984) );
  OAI21_X1 U17441 ( .B1(n15320), .B2(n16192), .A(n13986), .ZN(P2_U2986) );
  AND2_X1 U17442 ( .A1(n13987), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15257) );
  INV_X1 U17443 ( .A(n15257), .ZN(n15525) );
  OAI21_X1 U17444 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n13987), .A(
        n15525), .ZN(n14006) );
  NAND2_X1 U17445 ( .A1(n13989), .A2(n13988), .ZN(n15510) );
  INV_X1 U17446 ( .A(n13990), .ZN(n15509) );
  INV_X1 U17447 ( .A(n13991), .ZN(n15535) );
  NOR2_X1 U17448 ( .A1(n15509), .A2(n15535), .ZN(n13992) );
  XNOR2_X1 U17449 ( .A(n15510), .B(n13992), .ZN(n14004) );
  INV_X1 U17450 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19747) );
  OAI22_X1 U17451 ( .A1(n18921), .A2(n19747), .B1(n13994), .B2(n13993), .ZN(
        n13997) );
  OAI21_X1 U17452 ( .B1(n13995), .B2(n9682), .A(n15530), .ZN(n19006) );
  NOR2_X1 U17453 ( .A1(n19136), .A2(n19006), .ZN(n13996) );
  AOI211_X1 U17454 ( .C1(n13998), .C2(n19156), .A(n13997), .B(n13996), .ZN(
        n13999) );
  OAI21_X1 U17455 ( .B1(n15505), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n13999), .ZN(n14000) );
  AOI21_X1 U17456 ( .B1(n14004), .B2(n19131), .A(n14000), .ZN(n14001) );
  OAI21_X1 U17457 ( .B1(n14006), .B2(n19159), .A(n14001), .ZN(P2_U3037) );
  INV_X1 U17458 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18940) );
  OAI22_X1 U17459 ( .A1(n19129), .A2(n18940), .B1(n16190), .B2(n18934), .ZN(
        n14003) );
  OAI22_X1 U17460 ( .A1(n18935), .A2(n16160), .B1(n18921), .B2(n19747), .ZN(
        n14002) );
  AOI211_X1 U17461 ( .C1(n14004), .C2(n19124), .A(n14003), .B(n14002), .ZN(
        n14005) );
  OAI21_X1 U17462 ( .B1(n14006), .B2(n16194), .A(n14005), .ZN(P2_U3005) );
  OAI211_X1 U17463 ( .C1(n14009), .C2(n14008), .A(n14007), .B(n15136), .ZN(
        n14015) );
  INV_X1 U17464 ( .A(n14718), .ZN(n14012) );
  NOR2_X1 U17465 ( .A1(n14010), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14011) );
  MUX2_X1 U17466 ( .A(n14012), .B(n14011), .S(n19177), .Z(n14669) );
  NAND2_X1 U17467 ( .A1(n14669), .A2(n13698), .ZN(n14013) );
  XNOR2_X1 U17468 ( .A(n14013), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14014) );
  XNOR2_X1 U17469 ( .A(n14015), .B(n14014), .ZN(n14042) );
  NAND2_X1 U17470 ( .A1(n15140), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14016) );
  XNOR2_X1 U17471 ( .A(n14016), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14040) );
  NAND2_X1 U17472 ( .A1(n11927), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14019) );
  AOI22_X1 U17473 ( .A1(n14017), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n14018) );
  OAI211_X1 U17474 ( .C1(n14020), .C2(n14742), .A(n14019), .B(n14018), .ZN(
        n14024) );
  NAND3_X1 U17475 ( .A1(n14025), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15552), .ZN(n14028) );
  NOR4_X1 U17476 ( .A1(n15308), .A2(n9989), .A3(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A4(n14026), .ZN(n14027) );
  INV_X1 U17477 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19786) );
  NOR2_X1 U17478 ( .A1(n18921), .A2(n19786), .ZN(n14037) );
  AND2_X1 U17479 ( .A1(n14028), .A2(n10117), .ZN(n14032) );
  AOI222_X1 U17480 ( .A1(n11995), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n12000), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n12279), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14029) );
  XNOR2_X1 U17481 ( .A(n14030), .B(n14029), .ZN(n18975) );
  OAI211_X1 U17482 ( .C1(n14739), .C2(n16248), .A(n14032), .B(n14031), .ZN(
        n14033) );
  AOI21_X1 U17483 ( .B1(n14040), .B2(n16228), .A(n14033), .ZN(n14034) );
  OAI21_X1 U17484 ( .B1(n14042), .B2(n19166), .A(n14034), .ZN(P2_U3015) );
  NOR2_X1 U17485 ( .A1(n16190), .A2(n14035), .ZN(n14036) );
  AOI211_X1 U17486 ( .C1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n16184), .A(
        n14037), .B(n14036), .ZN(n14038) );
  OAI21_X1 U17487 ( .B1(n14739), .B2(n16160), .A(n14038), .ZN(n14039) );
  AOI21_X1 U17488 ( .B1(n14040), .B2(n19123), .A(n14039), .ZN(n14041) );
  OAI21_X1 U17489 ( .B1(n14042), .B2(n16192), .A(n14041), .ZN(P2_U2983) );
  NAND2_X1 U17490 ( .A1(n14043), .A2(n19942), .ZN(n14056) );
  INV_X1 U17491 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20701) );
  INV_X1 U17492 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20693) );
  INV_X1 U17493 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20691) );
  NAND4_X1 U17494 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(P1_REIP_REG_12__SCAN_IN), .A4(P1_REIP_REG_11__SCAN_IN), .ZN(n14178) );
  NOR3_X1 U17495 ( .A1(n20693), .A2(n20691), .A3(n14178), .ZN(n15905) );
  NAND2_X1 U17496 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n15905), .ZN(n15888) );
  NAND2_X1 U17497 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n15891) );
  NOR2_X1 U17498 ( .A1(n15888), .A2(n15891), .ZN(n15875) );
  NAND3_X1 U17499 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n14044), .A3(n15875), 
        .ZN(n15861) );
  NOR2_X1 U17500 ( .A1(n20701), .A2(n15861), .ZN(n14164) );
  NAND2_X1 U17501 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n14164), .ZN(n14154) );
  INV_X1 U17502 ( .A(n14154), .ZN(n14045) );
  AND2_X1 U17503 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n14045), .ZN(n14122) );
  NAND2_X1 U17504 ( .A1(n14122), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14051) );
  AND2_X1 U17505 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n14052) );
  INV_X1 U17506 ( .A(n14052), .ZN(n14046) );
  NOR2_X1 U17507 ( .A1(n14051), .A2(n14046), .ZN(n14047) );
  AND2_X1 U17508 ( .A1(n14187), .A2(n14047), .ZN(n14097) );
  NAND3_X1 U17509 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .A3(P1_REIP_REG_27__SCAN_IN), .ZN(n14063) );
  INV_X1 U17510 ( .A(n14063), .ZN(n14048) );
  NAND3_X1 U17511 ( .A1(n14097), .A2(P1_REIP_REG_30__SCAN_IN), .A3(n14048), 
        .ZN(n14049) );
  AND2_X1 U17512 ( .A1(n15886), .A2(n14049), .ZN(n14064) );
  INV_X1 U17513 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14201) );
  INV_X1 U17514 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14050) );
  OAI22_X1 U17515 ( .A1(n15924), .A2(n14201), .B1(n14050), .B2(n19905), .ZN(
        n14054) );
  NOR2_X1 U17516 ( .A1(n19924), .A2(n14051), .ZN(n14123) );
  NAND2_X1 U17517 ( .A1(n14123), .A2(n14052), .ZN(n14102) );
  INV_X1 U17518 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n20720) );
  NOR4_X1 U17519 ( .A1(n14102), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14063), 
        .A4(n20720), .ZN(n14053) );
  AOI211_X1 U17520 ( .C1(n14064), .C2(P1_REIP_REG_31__SCAN_IN), .A(n14054), 
        .B(n14053), .ZN(n14055) );
  OAI211_X1 U17521 ( .C1(n14202), .C2(n19976), .A(n14056), .B(n14055), .ZN(
        P1_U2809) );
  INV_X1 U17522 ( .A(n14360), .ZN(n14268) );
  INV_X1 U17523 ( .A(n14058), .ZN(n14059) );
  AOI22_X1 U17524 ( .A1(n14070), .A2(n14060), .B1(n14059), .B2(n14091), .ZN(
        n14061) );
  XOR2_X1 U17525 ( .A(n14062), .B(n14061), .Z(n14492) );
  INV_X1 U17526 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14204) );
  NOR2_X1 U17527 ( .A1(n14102), .A2(n14063), .ZN(n14065) );
  OAI21_X1 U17528 ( .B1(n14065), .B2(P1_REIP_REG_30__SCAN_IN), .A(n14064), 
        .ZN(n14067) );
  AOI22_X1 U17529 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19962), .B1(
        n19961), .B2(n14357), .ZN(n14066) );
  OAI211_X1 U17530 ( .C1(n15924), .C2(n14204), .A(n14067), .B(n14066), .ZN(
        n14068) );
  AOI21_X1 U17531 ( .B1(n14492), .B2(n19948), .A(n14068), .ZN(n14069) );
  OAI21_X1 U17532 ( .B1(n14268), .B2(n19928), .A(n14069), .ZN(P1_U2810) );
  OAI21_X1 U17533 ( .B1(n14091), .B2(n14071), .A(n14070), .ZN(n14495) );
  NAND2_X1 U17534 ( .A1(n14367), .A2(n19942), .ZN(n14081) );
  INV_X1 U17535 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n20710) );
  INV_X1 U17536 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20712) );
  NOR2_X1 U17537 ( .A1(n20710), .A2(n20712), .ZN(n14075) );
  INV_X1 U17538 ( .A(n15886), .ZN(n14179) );
  AOI21_X1 U17539 ( .B1(n14097), .B2(n14075), .A(n14179), .ZN(n14090) );
  INV_X1 U17540 ( .A(n14365), .ZN(n14076) );
  AOI22_X1 U17541 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19962), .B1(
        n19961), .B2(n14076), .ZN(n14077) );
  OAI21_X1 U17542 ( .B1(n15924), .B2(n14205), .A(n14077), .ZN(n14079) );
  NOR4_X1 U17543 ( .A1(n14102), .A2(P1_REIP_REG_29__SCAN_IN), .A3(n20712), 
        .A4(n20710), .ZN(n14078) );
  AOI211_X1 U17544 ( .C1(n14090), .C2(P1_REIP_REG_29__SCAN_IN), .A(n14079), 
        .B(n14078), .ZN(n14080) );
  OAI211_X1 U17545 ( .C1(n19976), .C2(n14495), .A(n14081), .B(n14080), .ZN(
        P1_U2811) );
  OR2_X1 U17546 ( .A1(n14082), .A2(n14083), .ZN(n14085) );
  AOI22_X1 U17547 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19962), .B1(
        n19961), .B2(n14377), .ZN(n14086) );
  OAI21_X1 U17548 ( .B1(n15924), .B2(n14087), .A(n14086), .ZN(n14089) );
  NOR3_X1 U17549 ( .A1(n14102), .A2(P1_REIP_REG_28__SCAN_IN), .A3(n20712), 
        .ZN(n14088) );
  AOI211_X1 U17550 ( .C1(n14090), .C2(P1_REIP_REG_28__SCAN_IN), .A(n14089), 
        .B(n14088), .ZN(n14094) );
  AOI21_X1 U17551 ( .B1(n14092), .B2(n14103), .A(n14091), .ZN(n14512) );
  NAND2_X1 U17552 ( .A1(n14512), .A2(n19948), .ZN(n14093) );
  OAI211_X1 U17553 ( .C1(n14375), .C2(n19928), .A(n14094), .B(n14093), .ZN(
        P1_U2812) );
  AOI21_X1 U17554 ( .B1(n14096), .B2(n14109), .A(n14082), .ZN(n14384) );
  INV_X1 U17555 ( .A(n14384), .ZN(n14286) );
  INV_X1 U17556 ( .A(n14097), .ZN(n14098) );
  AND2_X1 U17557 ( .A1(n15886), .A2(n14098), .ZN(n14112) );
  OAI22_X1 U17558 ( .A1(n14099), .A2(n19905), .B1(n19950), .B2(n14382), .ZN(
        n14100) );
  AOI21_X1 U17559 ( .B1(n19967), .B2(P1_EBX_REG_27__SCAN_IN), .A(n14100), .ZN(
        n14101) );
  OAI21_X1 U17560 ( .B1(n14102), .B2(P1_REIP_REG_27__SCAN_IN), .A(n14101), 
        .ZN(n14106) );
  OAI21_X1 U17561 ( .B1(n9675), .B2(n14104), .A(n14103), .ZN(n14516) );
  NOR2_X1 U17562 ( .A1(n14516), .A2(n19976), .ZN(n14105) );
  AOI211_X1 U17563 ( .C1(P1_REIP_REG_27__SCAN_IN), .C2(n14112), .A(n14106), 
        .B(n14105), .ZN(n14107) );
  OAI21_X1 U17564 ( .B1(n14286), .B2(n19928), .A(n14107), .ZN(P1_U2813) );
  AOI21_X1 U17565 ( .B1(n14111), .B2(n14128), .A(n9675), .ZN(n14535) );
  AOI21_X1 U17566 ( .B1(n14123), .B2(P1_REIP_REG_25__SCAN_IN), .A(
        P1_REIP_REG_26__SCAN_IN), .ZN(n14116) );
  INV_X1 U17567 ( .A(n14112), .ZN(n14115) );
  AOI22_X1 U17568 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19962), .B1(
        n19961), .B2(n14393), .ZN(n14114) );
  NAND2_X1 U17569 ( .A1(n19967), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n14113) );
  OAI211_X1 U17570 ( .C1(n14116), .C2(n14115), .A(n14114), .B(n14113), .ZN(
        n14117) );
  AOI21_X1 U17571 ( .B1(n14535), .B2(n19948), .A(n14117), .ZN(n14118) );
  OAI21_X1 U17572 ( .B1(n14390), .B2(n19928), .A(n14118), .ZN(P1_U2814) );
  AOI21_X1 U17573 ( .B1(n14121), .B2(n14119), .A(n14120), .ZN(n14403) );
  INV_X1 U17574 ( .A(n14403), .ZN(n14211) );
  INV_X1 U17575 ( .A(n14122), .ZN(n14139) );
  INV_X1 U17576 ( .A(n14187), .ZN(n19959) );
  AOI21_X1 U17577 ( .B1(n19972), .B2(n14139), .A(n19959), .ZN(n14153) );
  OAI21_X1 U17578 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n19924), .A(n14153), 
        .ZN(n14132) );
  INV_X1 U17579 ( .A(n14123), .ZN(n14127) );
  OAI22_X1 U17580 ( .A1(n14124), .A2(n19905), .B1(n19950), .B2(n14401), .ZN(
        n14125) );
  AOI21_X1 U17581 ( .B1(n19967), .B2(P1_EBX_REG_25__SCAN_IN), .A(n14125), .ZN(
        n14126) );
  OAI21_X1 U17582 ( .B1(n14127), .B2(P1_REIP_REG_25__SCAN_IN), .A(n14126), 
        .ZN(n14131) );
  OAI21_X1 U17583 ( .B1(n14136), .B2(n14129), .A(n14128), .ZN(n14541) );
  NOR2_X1 U17584 ( .A1(n14541), .A2(n19976), .ZN(n14130) );
  AOI211_X1 U17585 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n14132), .A(n14131), 
        .B(n14130), .ZN(n14133) );
  OAI21_X1 U17586 ( .B1(n14211), .B2(n19928), .A(n14133), .ZN(P1_U2815) );
  OAI21_X1 U17587 ( .B1(n14151), .B2(n14135), .A(n14119), .ZN(n14411) );
  AOI21_X1 U17588 ( .B1(n14137), .B2(n14148), .A(n14136), .ZN(n14554) );
  INV_X1 U17589 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n14143) );
  INV_X1 U17590 ( .A(n14414), .ZN(n14138) );
  OAI22_X1 U17591 ( .A1(n14410), .A2(n19905), .B1(n19950), .B2(n14138), .ZN(
        n14141) );
  NOR3_X1 U17592 ( .A1(n19924), .A2(P1_REIP_REG_24__SCAN_IN), .A3(n14139), 
        .ZN(n14140) );
  AOI211_X1 U17593 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n19967), .A(n14141), .B(
        n14140), .ZN(n14142) );
  OAI21_X1 U17594 ( .B1(n14153), .B2(n14143), .A(n14142), .ZN(n14144) );
  AOI21_X1 U17595 ( .B1(n14554), .B2(n19948), .A(n14144), .ZN(n14145) );
  OAI21_X1 U17596 ( .B1(n14411), .B2(n19928), .A(n14145), .ZN(P1_U2816) );
  INV_X1 U17597 ( .A(n14165), .ZN(n14147) );
  OAI21_X1 U17598 ( .B1(n9646), .B2(n14147), .A(n14146), .ZN(n14149) );
  NAND2_X1 U17599 ( .A1(n14149), .A2(n14148), .ZN(n14557) );
  INV_X1 U17600 ( .A(n14150), .ZN(n14162) );
  AOI21_X1 U17601 ( .B1(n14152), .B2(n14162), .A(n14151), .ZN(n14421) );
  NAND2_X1 U17602 ( .A1(n14421), .A2(n19942), .ZN(n14160) );
  INV_X1 U17603 ( .A(n14153), .ZN(n14158) );
  INV_X1 U17604 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20908) );
  OAI21_X1 U17605 ( .B1(n19924), .B2(n14154), .A(n20908), .ZN(n14157) );
  INV_X1 U17606 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14213) );
  NOR2_X1 U17607 ( .A1(n15924), .A2(n14213), .ZN(n14156) );
  OAI22_X1 U17608 ( .A1(n11405), .A2(n19905), .B1(n19950), .B2(n14419), .ZN(
        n14155) );
  AOI211_X1 U17609 ( .C1(n14158), .C2(n14157), .A(n14156), .B(n14155), .ZN(
        n14159) );
  OAI211_X1 U17610 ( .C1(n14557), .C2(n19976), .A(n14160), .B(n14159), .ZN(
        P1_U2817) );
  AOI21_X1 U17611 ( .B1(n14163), .B2(n14161), .A(n14150), .ZN(n14430) );
  INV_X1 U17612 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20703) );
  NAND2_X1 U17613 ( .A1(n14164), .A2(n20703), .ZN(n14173) );
  XNOR2_X1 U17614 ( .A(n9646), .B(n14165), .ZN(n14577) );
  NAND2_X1 U17615 ( .A1(n14577), .A2(n19948), .ZN(n14172) );
  NAND2_X1 U17616 ( .A1(n19961), .A2(n14426), .ZN(n14169) );
  NAND2_X1 U17617 ( .A1(n19962), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14168) );
  NAND2_X1 U17618 ( .A1(n20701), .A2(n19972), .ZN(n15860) );
  INV_X1 U17619 ( .A(n15860), .ZN(n14166) );
  AOI21_X1 U17620 ( .B1(n15861), .B2(n19972), .A(n19959), .ZN(n15877) );
  INV_X1 U17621 ( .A(n15877), .ZN(n15867) );
  OAI21_X1 U17622 ( .B1(n14166), .B2(n15867), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14167) );
  NAND3_X1 U17623 ( .A1(n14169), .A2(n14168), .A3(n14167), .ZN(n14170) );
  AOI21_X1 U17624 ( .B1(n19967), .B2(P1_EBX_REG_22__SCAN_IN), .A(n14170), .ZN(
        n14171) );
  OAI211_X1 U17625 ( .C1(n19924), .C2(n14173), .A(n14172), .B(n14171), .ZN(
        n14174) );
  AOI21_X1 U17626 ( .B1(n14430), .B2(n19942), .A(n14174), .ZN(n14175) );
  INV_X1 U17627 ( .A(n14175), .ZN(P1_U2818) );
  AOI21_X1 U17628 ( .B1(n14177), .B2(n13800), .A(n14176), .ZN(n14341) );
  INV_X1 U17629 ( .A(n14341), .ZN(n14465) );
  OAI21_X1 U17630 ( .B1(n14178), .B2(n15887), .A(n15886), .ZN(n15932) );
  OAI21_X1 U17631 ( .B1(n14179), .B2(P1_REIP_REG_15__SCAN_IN), .A(n15932), 
        .ZN(n15915) );
  INV_X1 U17632 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20688) );
  NOR3_X1 U17633 ( .A1(n20688), .A2(n14180), .A3(n15945), .ZN(n15920) );
  NAND2_X1 U17634 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n15920), .ZN(n15914) );
  OAI21_X1 U17635 ( .B1(n20691), .B2(n15914), .A(n20693), .ZN(n14181) );
  OAI21_X1 U17636 ( .B1(n20693), .B2(n15915), .A(n14181), .ZN(n14186) );
  OAI21_X1 U17637 ( .B1(n9694), .B2(n14182), .A(n14248), .ZN(n14616) );
  AOI22_X1 U17638 ( .A1(P1_EBX_REG_16__SCAN_IN), .A2(n19967), .B1(n14462), 
        .B2(n19961), .ZN(n14183) );
  OAI21_X1 U17639 ( .B1(n19976), .B2(n14616), .A(n14183), .ZN(n14184) );
  AOI211_X1 U17640 ( .C1(n19962), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n14184), .B(n10704), .ZN(n14185) );
  OAI211_X1 U17641 ( .C1(n14465), .C2(n19928), .A(n14186), .B(n14185), .ZN(
        P1_U2824) );
  OAI21_X1 U17642 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19924), .A(n14187), .ZN(
        n14188) );
  AOI22_X1 U17643 ( .A1(n19962), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n14188), .ZN(n14189) );
  OAI21_X1 U17644 ( .B1(n19950), .B2(n14190), .A(n14189), .ZN(n14191) );
  AOI21_X1 U17645 ( .B1(n19967), .B2(P1_EBX_REG_2__SCAN_IN), .A(n14191), .ZN(
        n14192) );
  OAI21_X1 U17646 ( .B1(n19976), .B2(n14193), .A(n14192), .ZN(n14196) );
  NAND2_X1 U17647 ( .A1(n19972), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n14194) );
  NOR2_X1 U17648 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n14194), .ZN(n14195) );
  AOI211_X1 U17649 ( .C1(n14198), .C2(n14197), .A(n14196), .B(n14195), .ZN(
        n14199) );
  OAI21_X1 U17650 ( .B1(n19969), .B2(n14200), .A(n14199), .ZN(P1_U2838) );
  OAI22_X1 U17651 ( .A1(n14202), .A2(n14259), .B1(n14260), .B2(n14201), .ZN(
        P1_U2841) );
  INV_X1 U17652 ( .A(n14492), .ZN(n14203) );
  OAI222_X1 U17653 ( .A1(n14254), .A2(n14268), .B1(n14204), .B2(n14260), .C1(
        n14203), .C2(n14259), .ZN(P1_U2842) );
  INV_X1 U17654 ( .A(n14367), .ZN(n14206) );
  OAI222_X1 U17655 ( .A1(n14254), .A2(n14206), .B1(n14205), .B2(n14260), .C1(
        n14495), .C2(n14259), .ZN(P1_U2843) );
  AOI22_X1 U17656 ( .A1(n14512), .A2(n14223), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n14222), .ZN(n14207) );
  OAI21_X1 U17657 ( .B1(n14375), .B2(n14254), .A(n14207), .ZN(P1_U2844) );
  INV_X1 U17658 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14208) );
  OAI222_X1 U17659 ( .A1(n14254), .A2(n14286), .B1(n14208), .B2(n14260), .C1(
        n14516), .C2(n14259), .ZN(P1_U2845) );
  AOI22_X1 U17660 ( .A1(n14535), .A2(n14223), .B1(P1_EBX_REG_26__SCAN_IN), 
        .B2(n14222), .ZN(n14209) );
  OAI21_X1 U17661 ( .B1(n14390), .B2(n14254), .A(n14209), .ZN(P1_U2846) );
  INV_X1 U17662 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14210) );
  OAI222_X1 U17663 ( .A1(n14254), .A2(n14211), .B1(n14210), .B2(n14260), .C1(
        n14541), .C2(n14259), .ZN(P1_U2847) );
  AOI22_X1 U17664 ( .A1(n14554), .A2(n14223), .B1(P1_EBX_REG_24__SCAN_IN), 
        .B2(n14222), .ZN(n14212) );
  OAI21_X1 U17665 ( .B1(n14411), .B2(n14254), .A(n14212), .ZN(P1_U2848) );
  INV_X1 U17666 ( .A(n14421), .ZN(n14214) );
  OAI222_X1 U17667 ( .A1(n14214), .A2(n14254), .B1(n14213), .B2(n14260), .C1(
        n14557), .C2(n14259), .ZN(P1_U2849) );
  INV_X1 U17668 ( .A(n14430), .ZN(n14216) );
  AOI22_X1 U17669 ( .A1(n14577), .A2(n14223), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n14222), .ZN(n14215) );
  OAI21_X1 U17670 ( .B1(n14216), .B2(n14254), .A(n14215), .ZN(P1_U2850) );
  OR2_X1 U17671 ( .A1(n14217), .A2(n14218), .ZN(n14219) );
  AND2_X1 U17672 ( .A1(n14161), .A2(n14219), .ZN(n15870) );
  INV_X1 U17673 ( .A(n15870), .ZN(n14225) );
  NAND2_X1 U17674 ( .A1(n9680), .A2(n14220), .ZN(n14221) );
  NAND2_X1 U17675 ( .A1(n9646), .A2(n14221), .ZN(n15868) );
  INV_X1 U17676 ( .A(n15868), .ZN(n14584) );
  AOI22_X1 U17677 ( .A1(n14584), .A2(n14223), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n14222), .ZN(n14224) );
  OAI21_X1 U17678 ( .B1(n14225), .B2(n14254), .A(n14224), .ZN(P1_U2851) );
  NOR2_X1 U17679 ( .A1(n14226), .A2(n14227), .ZN(n14228) );
  OR2_X1 U17680 ( .A1(n14217), .A2(n14228), .ZN(n14319) );
  INV_X1 U17681 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14231) );
  OR2_X1 U17682 ( .A1(n14234), .A2(n14229), .ZN(n14230) );
  NAND2_X1 U17683 ( .A1(n9680), .A2(n14230), .ZN(n15876) );
  OAI222_X1 U17684 ( .A1(n14319), .A2(n14254), .B1(n14260), .B2(n14231), .C1(
        n15876), .C2(n14259), .ZN(P1_U2852) );
  NOR2_X1 U17685 ( .A1(n14243), .A2(n14232), .ZN(n14233) );
  OR2_X1 U17686 ( .A1(n14234), .A2(n14233), .ZN(n15896) );
  INV_X1 U17687 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14238) );
  AND2_X1 U17688 ( .A1(n14236), .A2(n14235), .ZN(n14237) );
  OR2_X1 U17689 ( .A1(n14237), .A2(n14226), .ZN(n15948) );
  OAI222_X1 U17690 ( .A1(n15896), .A2(n14259), .B1(n14238), .B2(n14260), .C1(
        n15948), .C2(n14254), .ZN(P1_U2853) );
  XOR2_X1 U17691 ( .A(n14241), .B(n14240), .Z(n15903) );
  INV_X1 U17692 ( .A(n15903), .ZN(n14334) );
  AND2_X1 U17693 ( .A1(n14250), .A2(n14242), .ZN(n14244) );
  OR2_X1 U17694 ( .A1(n14244), .A2(n14243), .ZN(n16010) );
  OAI22_X1 U17695 ( .A1(n16010), .A2(n14259), .B1(n15898), .B2(n14260), .ZN(
        n14245) );
  INV_X1 U17696 ( .A(n14245), .ZN(n14246) );
  OAI21_X1 U17697 ( .B1(n14334), .B2(n14254), .A(n14246), .ZN(P1_U2854) );
  NAND2_X1 U17698 ( .A1(n14248), .A2(n14247), .ZN(n14249) );
  AND2_X1 U17699 ( .A1(n14250), .A2(n14249), .ZN(n16021) );
  INV_X1 U17700 ( .A(n16021), .ZN(n14252) );
  INV_X1 U17701 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n15907) );
  OAI21_X1 U17702 ( .B1(n14176), .B2(n14251), .A(n14240), .ZN(n15909) );
  OAI222_X1 U17703 ( .A1(n14252), .A2(n14259), .B1(n14260), .B2(n15907), .C1(
        n15909), .C2(n14254), .ZN(P1_U2855) );
  INV_X1 U17704 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14253) );
  OAI222_X1 U17705 ( .A1(n14465), .A2(n14254), .B1(n14260), .B2(n14253), .C1(
        n14616), .C2(n14259), .ZN(P1_U2856) );
  XOR2_X1 U17706 ( .A(n14256), .B(n14255), .Z(n19943) );
  INV_X1 U17707 ( .A(n19943), .ZN(n14351) );
  INV_X1 U17708 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n14261) );
  XNOR2_X1 U17709 ( .A(n14258), .B(n14257), .ZN(n19940) );
  OAI222_X1 U17710 ( .A1(n14254), .A2(n14351), .B1(n14261), .B2(n14260), .C1(
        n14259), .C2(n19940), .ZN(P1_U2866) );
  INV_X1 U17711 ( .A(n14262), .ZN(n14263) );
  AOI22_X1 U17712 ( .A1(n14344), .A2(n14264), .B1(n14342), .B2(
        P1_EAX_REG_30__SCAN_IN), .ZN(n14265) );
  OAI21_X1 U17713 ( .B1(n16360), .B2(n14337), .A(n14265), .ZN(n14266) );
  AOI21_X1 U17714 ( .B1(n14345), .B2(DATAI_30_), .A(n14266), .ZN(n14267) );
  OAI21_X1 U17715 ( .B1(n14268), .B2(n14285), .A(n14267), .ZN(P1_U2874) );
  NAND2_X1 U17716 ( .A1(n14367), .A2(n14340), .ZN(n14273) );
  AOI22_X1 U17717 ( .A1(n14344), .A2(n14269), .B1(n14342), .B2(
        P1_EAX_REG_29__SCAN_IN), .ZN(n14272) );
  NAND2_X1 U17718 ( .A1(n14345), .A2(DATAI_29_), .ZN(n14271) );
  NAND2_X1 U17719 ( .A1(n14346), .A2(BUF1_REG_29__SCAN_IN), .ZN(n14270) );
  NAND4_X1 U17720 ( .A1(n14273), .A2(n14272), .A3(n14271), .A4(n14270), .ZN(
        P1_U2875) );
  INV_X1 U17721 ( .A(n14375), .ZN(n14274) );
  NAND2_X1 U17722 ( .A1(n14274), .A2(n14340), .ZN(n14279) );
  AOI22_X1 U17723 ( .A1(n14344), .A2(n14275), .B1(n14342), .B2(
        P1_EAX_REG_28__SCAN_IN), .ZN(n14278) );
  NAND2_X1 U17724 ( .A1(n14345), .A2(DATAI_28_), .ZN(n14277) );
  NAND2_X1 U17725 ( .A1(n14346), .A2(BUF1_REG_28__SCAN_IN), .ZN(n14276) );
  NAND4_X1 U17726 ( .A1(n14279), .A2(n14278), .A3(n14277), .A4(n14276), .ZN(
        P1_U2876) );
  INV_X1 U17727 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n14282) );
  AOI22_X1 U17728 ( .A1(n14344), .A2(n14280), .B1(n14342), .B2(
        P1_EAX_REG_27__SCAN_IN), .ZN(n14281) );
  OAI21_X1 U17729 ( .B1(n14282), .B2(n14337), .A(n14281), .ZN(n14283) );
  AOI21_X1 U17730 ( .B1(n14345), .B2(DATAI_27_), .A(n14283), .ZN(n14284) );
  OAI21_X1 U17731 ( .B1(n14286), .B2(n14285), .A(n14284), .ZN(P1_U2877) );
  INV_X1 U17732 ( .A(n14390), .ZN(n14287) );
  NAND2_X1 U17733 ( .A1(n14287), .A2(n14340), .ZN(n14292) );
  AOI22_X1 U17734 ( .A1(n14344), .A2(n14288), .B1(n14342), .B2(
        P1_EAX_REG_26__SCAN_IN), .ZN(n14291) );
  NAND2_X1 U17735 ( .A1(n14345), .A2(DATAI_26_), .ZN(n14290) );
  NAND2_X1 U17736 ( .A1(n14346), .A2(BUF1_REG_26__SCAN_IN), .ZN(n14289) );
  NAND4_X1 U17737 ( .A1(n14292), .A2(n14291), .A3(n14290), .A4(n14289), .ZN(
        P1_U2878) );
  NAND2_X1 U17738 ( .A1(n14403), .A2(n14340), .ZN(n14297) );
  AOI22_X1 U17739 ( .A1(n14344), .A2(n14293), .B1(n14342), .B2(
        P1_EAX_REG_25__SCAN_IN), .ZN(n14296) );
  NAND2_X1 U17740 ( .A1(n14345), .A2(DATAI_25_), .ZN(n14295) );
  NAND2_X1 U17741 ( .A1(n14346), .A2(BUF1_REG_25__SCAN_IN), .ZN(n14294) );
  NAND4_X1 U17742 ( .A1(n14297), .A2(n14296), .A3(n14295), .A4(n14294), .ZN(
        P1_U2879) );
  INV_X1 U17743 ( .A(n14411), .ZN(n14298) );
  NAND2_X1 U17744 ( .A1(n14298), .A2(n14340), .ZN(n14303) );
  AOI22_X1 U17745 ( .A1(n14344), .A2(n14299), .B1(n14342), .B2(
        P1_EAX_REG_24__SCAN_IN), .ZN(n14302) );
  NAND2_X1 U17746 ( .A1(n14345), .A2(DATAI_24_), .ZN(n14301) );
  NAND2_X1 U17747 ( .A1(n14346), .A2(BUF1_REG_24__SCAN_IN), .ZN(n14300) );
  NAND4_X1 U17748 ( .A1(n14303), .A2(n14302), .A3(n14301), .A4(n14300), .ZN(
        P1_U2880) );
  NAND2_X1 U17749 ( .A1(n14421), .A2(n14340), .ZN(n14308) );
  AOI22_X1 U17750 ( .A1(n14344), .A2(n14304), .B1(n14342), .B2(
        P1_EAX_REG_23__SCAN_IN), .ZN(n14307) );
  NAND2_X1 U17751 ( .A1(n14345), .A2(DATAI_23_), .ZN(n14306) );
  NAND2_X1 U17752 ( .A1(n14346), .A2(BUF1_REG_23__SCAN_IN), .ZN(n14305) );
  NAND4_X1 U17753 ( .A1(n14308), .A2(n14307), .A3(n14306), .A4(n14305), .ZN(
        P1_U2881) );
  NAND2_X1 U17754 ( .A1(n14430), .A2(n14340), .ZN(n14313) );
  AOI22_X1 U17755 ( .A1(n14344), .A2(n14309), .B1(n14342), .B2(
        P1_EAX_REG_22__SCAN_IN), .ZN(n14312) );
  NAND2_X1 U17756 ( .A1(n14345), .A2(DATAI_22_), .ZN(n14311) );
  NAND2_X1 U17757 ( .A1(n14346), .A2(BUF1_REG_22__SCAN_IN), .ZN(n14310) );
  NAND4_X1 U17758 ( .A1(n14313), .A2(n14312), .A3(n14311), .A4(n14310), .ZN(
        P1_U2882) );
  INV_X1 U17759 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16376) );
  NAND2_X1 U17760 ( .A1(n14345), .A2(DATAI_21_), .ZN(n14316) );
  AOI22_X1 U17761 ( .A1(n14344), .A2(n14314), .B1(n14342), .B2(
        P1_EAX_REG_21__SCAN_IN), .ZN(n14315) );
  OAI211_X1 U17762 ( .C1(n16376), .C2(n14337), .A(n14316), .B(n14315), .ZN(
        n14317) );
  AOI21_X1 U17763 ( .B1(n15870), .B2(n14340), .A(n14317), .ZN(n14318) );
  INV_X1 U17764 ( .A(n14318), .ZN(P1_U2883) );
  NAND2_X1 U17765 ( .A1(n15880), .A2(n14340), .ZN(n14324) );
  AOI22_X1 U17766 ( .A1(n14344), .A2(n14320), .B1(n14342), .B2(
        P1_EAX_REG_20__SCAN_IN), .ZN(n14323) );
  NAND2_X1 U17767 ( .A1(n14345), .A2(DATAI_20_), .ZN(n14322) );
  NAND2_X1 U17768 ( .A1(n14346), .A2(BUF1_REG_20__SCAN_IN), .ZN(n14321) );
  NAND4_X1 U17769 ( .A1(n14324), .A2(n14323), .A3(n14322), .A4(n14321), .ZN(
        P1_U2884) );
  INV_X1 U17770 ( .A(n15948), .ZN(n15893) );
  INV_X1 U17771 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16380) );
  NAND2_X1 U17772 ( .A1(n14345), .A2(DATAI_19_), .ZN(n14327) );
  AOI22_X1 U17773 ( .A1(n14344), .A2(n14325), .B1(n14342), .B2(
        P1_EAX_REG_19__SCAN_IN), .ZN(n14326) );
  OAI211_X1 U17774 ( .C1(n16380), .C2(n14337), .A(n14327), .B(n14326), .ZN(
        n14328) );
  AOI21_X1 U17775 ( .B1(n15893), .B2(n14340), .A(n14328), .ZN(n14329) );
  INV_X1 U17776 ( .A(n14329), .ZN(P1_U2885) );
  AOI22_X1 U17777 ( .A1(n14344), .A2(n14330), .B1(n14342), .B2(
        P1_EAX_REG_18__SCAN_IN), .ZN(n14331) );
  OAI21_X1 U17778 ( .B1(n14337), .B2(n16382), .A(n14331), .ZN(n14332) );
  AOI21_X1 U17779 ( .B1(n14345), .B2(DATAI_18_), .A(n14332), .ZN(n14333) );
  OAI21_X1 U17780 ( .B1(n14334), .B2(n14285), .A(n14333), .ZN(P1_U2886) );
  AOI22_X1 U17781 ( .A1(n14344), .A2(n14335), .B1(n14342), .B2(
        P1_EAX_REG_17__SCAN_IN), .ZN(n14336) );
  OAI21_X1 U17782 ( .B1(n15130), .B2(n14337), .A(n14336), .ZN(n14338) );
  AOI21_X1 U17783 ( .B1(n14345), .B2(DATAI_17_), .A(n14338), .ZN(n14339) );
  OAI21_X1 U17784 ( .B1(n15909), .B2(n14285), .A(n14339), .ZN(P1_U2887) );
  NAND2_X1 U17785 ( .A1(n14341), .A2(n14340), .ZN(n14350) );
  AOI22_X1 U17786 ( .A1(n14344), .A2(n14343), .B1(n14342), .B2(
        P1_EAX_REG_16__SCAN_IN), .ZN(n14349) );
  NAND2_X1 U17787 ( .A1(n14345), .A2(DATAI_16_), .ZN(n14348) );
  NAND2_X1 U17788 ( .A1(n14346), .A2(BUF1_REG_16__SCAN_IN), .ZN(n14347) );
  NAND4_X1 U17789 ( .A1(n14350), .A2(n14349), .A3(n14348), .A4(n14347), .ZN(
        P1_U2888) );
  OAI222_X1 U17790 ( .A1(n14352), .A2(n20100), .B1(n14353), .B2(n19997), .C1(
        n14285), .C2(n14351), .ZN(P1_U2898) );
  OAI222_X1 U17791 ( .A1(n14285), .A2(n16003), .B1(n14353), .B2(n11111), .C1(
        n14352), .C2(n20094), .ZN(P1_U2899) );
  NAND2_X1 U17792 ( .A1(n14355), .A2(n14354), .ZN(n14356) );
  XNOR2_X1 U17793 ( .A(n14356), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14494) );
  NAND2_X1 U17794 ( .A1(n15976), .A2(n14357), .ZN(n14358) );
  NAND2_X1 U17795 ( .A1(n10704), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14486) );
  OAI211_X1 U17796 ( .C1(n20024), .C2(n20880), .A(n14358), .B(n14486), .ZN(
        n14359) );
  AOI21_X1 U17797 ( .B1(n14360), .B2(n14447), .A(n14359), .ZN(n14361) );
  OAI21_X1 U17798 ( .B1(n14494), .B2(n20030), .A(n14361), .ZN(P1_U2969) );
  XNOR2_X1 U17799 ( .A(n9611), .B(n14499), .ZN(n14362) );
  XNOR2_X1 U17800 ( .A(n14363), .B(n14362), .ZN(n14504) );
  NAND2_X1 U17801 ( .A1(n10704), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14498) );
  NAND2_X1 U17802 ( .A1(n20013), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14364) );
  OAI211_X1 U17803 ( .C1(n20023), .C2(n14365), .A(n14498), .B(n14364), .ZN(
        n14366) );
  AOI21_X1 U17804 ( .B1(n14367), .B2(n14447), .A(n14366), .ZN(n14368) );
  OAI21_X1 U17805 ( .B1(n14504), .B2(n20030), .A(n14368), .ZN(P1_U2970) );
  NAND2_X1 U17806 ( .A1(n9611), .A2(n14528), .ZN(n14386) );
  NAND2_X1 U17807 ( .A1(n14417), .A2(n14386), .ZN(n14372) );
  OAI21_X1 U17808 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n14369), .A(
        n14372), .ZN(n14371) );
  MUX2_X1 U17809 ( .A(n14520), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n15980), .Z(n14370) );
  OAI211_X1 U17810 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n14372), .A(
        n14371), .B(n14370), .ZN(n14374) );
  XNOR2_X1 U17811 ( .A(n14374), .B(n14373), .ZN(n14515) );
  NAND2_X1 U17812 ( .A1(n10704), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14505) );
  OAI21_X1 U17813 ( .B1(n20024), .B2(n20810), .A(n14505), .ZN(n14376) );
  MUX2_X1 U17814 ( .A(n14379), .B(n14378), .S(n15980), .Z(n14380) );
  XNOR2_X1 U17815 ( .A(n14380), .B(n14520), .ZN(n14525) );
  NOR2_X1 U17816 ( .A1(n20036), .A2(n20712), .ZN(n14517) );
  AOI21_X1 U17817 ( .B1(n20013), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14517), .ZN(n14381) );
  OAI21_X1 U17818 ( .B1(n20023), .B2(n14382), .A(n14381), .ZN(n14383) );
  AOI21_X1 U17819 ( .B1(n14384), .B2(n14447), .A(n14383), .ZN(n14385) );
  OAI21_X1 U17820 ( .B1(n20030), .B2(n14525), .A(n14385), .ZN(P1_U2972) );
  OAI211_X1 U17821 ( .C1(n14437), .C2(n14417), .A(n14387), .B(n14386), .ZN(
        n14388) );
  XNOR2_X1 U17822 ( .A(n14388), .B(n14529), .ZN(n14537) );
  NAND2_X1 U17823 ( .A1(n10704), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14532) );
  OAI21_X1 U17824 ( .B1(n20024), .B2(n14389), .A(n14532), .ZN(n14392) );
  NOR2_X1 U17825 ( .A1(n14390), .A2(n15947), .ZN(n14391) );
  OAI21_X1 U17826 ( .B1(n20030), .B2(n14537), .A(n14394), .ZN(P1_U2973) );
  OR3_X1 U17827 ( .A1(n14417), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14397) );
  NAND2_X1 U17828 ( .A1(n14395), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14406) );
  OR2_X1 U17829 ( .A1(n14406), .A2(n14408), .ZN(n14396) );
  MUX2_X1 U17830 ( .A(n14397), .B(n14396), .S(n15980), .Z(n14399) );
  XNOR2_X1 U17831 ( .A(n14399), .B(n14398), .ZN(n14545) );
  INV_X1 U17832 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20707) );
  NOR2_X1 U17833 ( .A1(n20036), .A2(n20707), .ZN(n14539) );
  AOI21_X1 U17834 ( .B1(n20013), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n14539), .ZN(n14400) );
  OAI21_X1 U17835 ( .B1(n20023), .B2(n14401), .A(n14400), .ZN(n14402) );
  AOI21_X1 U17836 ( .B1(n14403), .B2(n14447), .A(n14402), .ZN(n14404) );
  OAI21_X1 U17837 ( .B1(n20030), .B2(n14545), .A(n14404), .ZN(P1_U2974) );
  INV_X1 U17838 ( .A(n14417), .ZN(n14405) );
  NAND2_X1 U17839 ( .A1(n14405), .A2(n14406), .ZN(n14407) );
  MUX2_X1 U17840 ( .A(n14407), .B(n14406), .S(n15980), .Z(n14409) );
  XNOR2_X1 U17841 ( .A(n14409), .B(n14408), .ZN(n14556) );
  NAND2_X1 U17842 ( .A1(n10704), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14546) );
  OAI21_X1 U17843 ( .B1(n20024), .B2(n14410), .A(n14546), .ZN(n14413) );
  NOR2_X1 U17844 ( .A1(n14411), .A2(n15947), .ZN(n14412) );
  AOI211_X1 U17845 ( .C1(n15976), .C2(n14414), .A(n14413), .B(n14412), .ZN(
        n14415) );
  OAI21_X1 U17846 ( .B1(n20030), .B2(n14556), .A(n14415), .ZN(P1_U2975) );
  XNOR2_X1 U17847 ( .A(n9611), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14416) );
  XNOR2_X1 U17848 ( .A(n14417), .B(n14416), .ZN(n14566) );
  NOR2_X1 U17849 ( .A1(n20036), .A2(n20908), .ZN(n14558) );
  AOI21_X1 U17850 ( .B1(n20013), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n14558), .ZN(n14418) );
  OAI21_X1 U17851 ( .B1(n20023), .B2(n14419), .A(n14418), .ZN(n14420) );
  AOI21_X1 U17852 ( .B1(n14421), .B2(n14447), .A(n14420), .ZN(n14422) );
  OAI21_X1 U17853 ( .B1(n14566), .B2(n20030), .A(n14422), .ZN(P1_U2976) );
  NAND2_X1 U17854 ( .A1(n14424), .A2(n14423), .ZN(n14425) );
  XNOR2_X1 U17855 ( .A(n14425), .B(n14572), .ZN(n14579) );
  INV_X1 U17856 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14428) );
  NAND2_X1 U17857 ( .A1(n15976), .A2(n14426), .ZN(n14427) );
  NAND2_X1 U17858 ( .A1(n10704), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n14573) );
  OAI211_X1 U17859 ( .C1(n20024), .C2(n14428), .A(n14427), .B(n14573), .ZN(
        n14429) );
  AOI21_X1 U17860 ( .B1(n14430), .B2(n14447), .A(n14429), .ZN(n14431) );
  OAI21_X1 U17861 ( .B1(n20030), .B2(n14579), .A(n14431), .ZN(P1_U2977) );
  OR2_X1 U17862 ( .A1(n15980), .A2(n16014), .ZN(n14433) );
  AND2_X1 U17863 ( .A1(n14432), .A2(n14433), .ZN(n14599) );
  NOR2_X1 U17864 ( .A1(n9611), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14597) );
  INV_X1 U17865 ( .A(n14432), .ZN(n14434) );
  AND2_X1 U17866 ( .A1(n15980), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14596) );
  AOI22_X1 U17867 ( .A1(n14599), .A2(n14597), .B1(n14434), .B2(n14596), .ZN(
        n14444) );
  NOR2_X1 U17868 ( .A1(n14444), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14443) );
  INV_X1 U17869 ( .A(n14596), .ZN(n14435) );
  NOR3_X1 U17870 ( .A1(n14432), .A2(n14589), .A3(n14435), .ZN(n14436) );
  AOI21_X1 U17871 ( .B1(n14443), .B2(n14437), .A(n14436), .ZN(n14439) );
  XNOR2_X1 U17872 ( .A(n14439), .B(n14438), .ZN(n14587) );
  NAND2_X1 U17873 ( .A1(n10704), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14580) );
  NAND2_X1 U17874 ( .A1(n20013), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14440) );
  OAI211_X1 U17875 ( .C1(n20023), .C2(n15862), .A(n14580), .B(n14440), .ZN(
        n14441) );
  AOI21_X1 U17876 ( .B1(n15870), .B2(n14447), .A(n14441), .ZN(n14442) );
  OAI21_X1 U17877 ( .B1(n14587), .B2(n20030), .A(n14442), .ZN(P1_U2978) );
  AOI21_X1 U17878 ( .B1(n14444), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n14443), .ZN(n14595) );
  NAND2_X1 U17879 ( .A1(n15976), .A2(n15874), .ZN(n14445) );
  NAND2_X1 U17880 ( .A1(n10704), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n14588) );
  OAI211_X1 U17881 ( .C1(n20024), .C2(n15883), .A(n14445), .B(n14588), .ZN(
        n14446) );
  AOI21_X1 U17882 ( .B1(n15880), .B2(n14447), .A(n14446), .ZN(n14448) );
  OAI21_X1 U17883 ( .B1(n14595), .B2(n20030), .A(n14448), .ZN(P1_U2979) );
  OAI21_X1 U17884 ( .B1(n14450), .B2(n14449), .A(n14432), .ZN(n16011) );
  INV_X1 U17885 ( .A(n14451), .ZN(n15897) );
  AOI22_X1 U17886 ( .A1(n20013), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n10704), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14452) );
  OAI21_X1 U17887 ( .B1(n15897), .B2(n20023), .A(n14452), .ZN(n14453) );
  AOI21_X1 U17888 ( .B1(n15903), .B2(n14447), .A(n14453), .ZN(n14454) );
  OAI21_X1 U17889 ( .B1(n20030), .B2(n16011), .A(n14454), .ZN(P1_U2981) );
  AOI21_X1 U17890 ( .B1(n14456), .B2(n9679), .A(n14455), .ZN(n15965) );
  NAND2_X1 U17891 ( .A1(n15965), .A2(n15963), .ZN(n15954) );
  AOI21_X1 U17892 ( .B1(n15954), .B2(n15962), .A(n14457), .ZN(n14459) );
  INV_X1 U17893 ( .A(n14457), .ZN(n14458) );
  OAI22_X1 U17894 ( .A1(n14459), .A2(n15953), .B1(n14458), .B2(n15954), .ZN(
        n14619) );
  NAND2_X1 U17895 ( .A1(n14619), .A2(n20019), .ZN(n14464) );
  NAND2_X1 U17896 ( .A1(n10704), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n14615) );
  OAI21_X1 U17897 ( .B1(n20024), .B2(n14460), .A(n14615), .ZN(n14461) );
  AOI21_X1 U17898 ( .B1(n14462), .B2(n15976), .A(n14461), .ZN(n14463) );
  OAI211_X1 U17899 ( .C1(n15947), .C2(n14465), .A(n14464), .B(n14463), .ZN(
        P1_U2983) );
  INV_X1 U17900 ( .A(n13774), .ZN(n14469) );
  INV_X1 U17901 ( .A(n14466), .ZN(n14467) );
  AOI21_X1 U17902 ( .B1(n14469), .B2(n14468), .A(n14467), .ZN(n15972) );
  AND2_X1 U17903 ( .A1(n14470), .A2(n14471), .ZN(n15971) );
  NAND2_X1 U17904 ( .A1(n15972), .A2(n15971), .ZN(n15970) );
  NAND2_X1 U17905 ( .A1(n15970), .A2(n14471), .ZN(n14472) );
  XOR2_X1 U17906 ( .A(n14473), .B(n14472), .Z(n16039) );
  NAND2_X1 U17907 ( .A1(n16039), .A2(n20019), .ZN(n14477) );
  NAND2_X1 U17908 ( .A1(n10704), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n16034) );
  OAI21_X1 U17909 ( .B1(n20024), .B2(n13757), .A(n16034), .ZN(n14474) );
  AOI21_X1 U17910 ( .B1(n15976), .B2(n14475), .A(n14474), .ZN(n14476) );
  OAI211_X1 U17911 ( .C1(n15947), .C2(n14478), .A(n14477), .B(n14476), .ZN(
        P1_U2986) );
  INV_X1 U17912 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16074) );
  MUX2_X1 U17913 ( .A(n15979), .B(n13774), .S(n15980), .Z(n14479) );
  XOR2_X1 U17914 ( .A(n16074), .B(n14479), .Z(n16072) );
  INV_X1 U17915 ( .A(n16072), .ZN(n14485) );
  AOI22_X1 U17916 ( .A1(n20013), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n10704), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14480) );
  OAI21_X1 U17917 ( .B1(n20023), .B2(n14481), .A(n14480), .ZN(n14482) );
  AOI21_X1 U17918 ( .B1(n14483), .B2(n14447), .A(n14482), .ZN(n14484) );
  OAI21_X1 U17919 ( .B1(n14485), .B2(n20030), .A(n14484), .ZN(P1_U2989) );
  INV_X1 U17920 ( .A(n14486), .ZN(n14491) );
  AOI21_X1 U17921 ( .B1(n14489), .B2(n14488), .A(n14487), .ZN(n14490) );
  AOI211_X1 U17922 ( .C1(n14492), .C2(n20059), .A(n14491), .B(n14490), .ZN(
        n14493) );
  OAI21_X1 U17923 ( .B1(n14494), .B2(n16106), .A(n14493), .ZN(P1_U3001) );
  INV_X1 U17924 ( .A(n14495), .ZN(n14502) );
  INV_X1 U17925 ( .A(n14496), .ZN(n14500) );
  NAND3_X1 U17926 ( .A1(n14518), .A2(n14507), .A3(n14499), .ZN(n14497) );
  OAI211_X1 U17927 ( .C1(n14500), .C2(n14499), .A(n14498), .B(n14497), .ZN(
        n14501) );
  AOI21_X1 U17928 ( .B1(n14502), .B2(n20059), .A(n14501), .ZN(n14503) );
  OAI21_X1 U17929 ( .B1(n14504), .B2(n16106), .A(n14503), .ZN(P1_U3002) );
  INV_X1 U17930 ( .A(n14521), .ZN(n14511) );
  INV_X1 U17931 ( .A(n14505), .ZN(n14510) );
  NOR3_X1 U17932 ( .A1(n14508), .A2(n14507), .A3(n14506), .ZN(n14509) );
  AOI211_X1 U17933 ( .C1(n14511), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14510), .B(n14509), .ZN(n14514) );
  NAND2_X1 U17934 ( .A1(n14512), .A2(n20059), .ZN(n14513) );
  OAI211_X1 U17935 ( .C1(n14515), .C2(n16106), .A(n14514), .B(n14513), .ZN(
        P1_U3003) );
  INV_X1 U17936 ( .A(n14516), .ZN(n14523) );
  AOI21_X1 U17937 ( .B1(n14518), .B2(n14520), .A(n14517), .ZN(n14519) );
  OAI21_X1 U17938 ( .B1(n14521), .B2(n14520), .A(n14519), .ZN(n14522) );
  AOI21_X1 U17939 ( .B1(n14523), .B2(n20059), .A(n14522), .ZN(n14524) );
  OAI21_X1 U17940 ( .B1(n14525), .B2(n16106), .A(n14524), .ZN(P1_U3004) );
  INV_X1 U17941 ( .A(n14526), .ZN(n14548) );
  NOR3_X1 U17942 ( .A1(n14527), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n14548), .ZN(n14538) );
  OAI21_X1 U17943 ( .B1(n14540), .B2(n14538), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14533) );
  INV_X1 U17944 ( .A(n14527), .ZN(n14559) );
  INV_X1 U17945 ( .A(n14528), .ZN(n14530) );
  NAND3_X1 U17946 ( .A1(n14559), .A2(n14530), .A3(n14529), .ZN(n14531) );
  NAND3_X1 U17947 ( .A1(n14533), .A2(n14532), .A3(n14531), .ZN(n14534) );
  AOI21_X1 U17948 ( .B1(n14535), .B2(n20059), .A(n14534), .ZN(n14536) );
  OAI21_X1 U17949 ( .B1(n14537), .B2(n16106), .A(n14536), .ZN(P1_U3005) );
  AOI211_X1 U17950 ( .C1(n14540), .C2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n14539), .B(n14538), .ZN(n14544) );
  INV_X1 U17951 ( .A(n14541), .ZN(n14542) );
  NAND2_X1 U17952 ( .A1(n14542), .A2(n20059), .ZN(n14543) );
  OAI211_X1 U17953 ( .C1(n14545), .C2(n16106), .A(n14544), .B(n14543), .ZN(
        P1_U3006) );
  INV_X1 U17954 ( .A(n14546), .ZN(n14553) );
  INV_X1 U17955 ( .A(n14547), .ZN(n14549) );
  OAI21_X1 U17956 ( .B1(n14549), .B2(n16046), .A(n14548), .ZN(n14551) );
  AOI21_X1 U17957 ( .B1(n14559), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14550) );
  AOI21_X1 U17958 ( .B1(n14562), .B2(n14551), .A(n14550), .ZN(n14552) );
  AOI211_X1 U17959 ( .C1(n14554), .C2(n20059), .A(n14553), .B(n14552), .ZN(
        n14555) );
  OAI21_X1 U17960 ( .B1(n14556), .B2(n16106), .A(n14555), .ZN(P1_U3007) );
  INV_X1 U17961 ( .A(n14557), .ZN(n14564) );
  AOI21_X1 U17962 ( .B1(n14559), .B2(n14561), .A(n14558), .ZN(n14560) );
  OAI21_X1 U17963 ( .B1(n14562), .B2(n14561), .A(n14560), .ZN(n14563) );
  AOI21_X1 U17964 ( .B1(n14564), .B2(n20059), .A(n14563), .ZN(n14565) );
  OAI21_X1 U17965 ( .B1(n14566), .B2(n16106), .A(n14565), .ZN(P1_U3008) );
  INV_X1 U17966 ( .A(n14567), .ZN(n14569) );
  AOI22_X1 U17967 ( .A1(n20066), .A2(n14569), .B1(n16046), .B2(n14568), .ZN(
        n16042) );
  OR2_X1 U17968 ( .A1(n16042), .A2(n14570), .ZN(n14605) );
  NAND2_X1 U17969 ( .A1(n10042), .A2(n14572), .ZN(n14575) );
  NOR4_X1 U17970 ( .A1(n14605), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n14600), .A4(n14589), .ZN(n14581) );
  OAI21_X1 U17971 ( .B1(n14581), .B2(n14583), .A(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14574) );
  OAI211_X1 U17972 ( .C1(n14605), .C2(n14575), .A(n14574), .B(n14573), .ZN(
        n14576) );
  AOI21_X1 U17973 ( .B1(n14577), .B2(n20059), .A(n14576), .ZN(n14578) );
  OAI21_X1 U17974 ( .B1(n14579), .B2(n16106), .A(n14578), .ZN(P1_U3009) );
  INV_X1 U17975 ( .A(n14580), .ZN(n14582) );
  AOI211_X1 U17976 ( .C1(n14583), .C2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n14582), .B(n14581), .ZN(n14586) );
  NAND2_X1 U17977 ( .A1(n14584), .A2(n20059), .ZN(n14585) );
  OAI211_X1 U17978 ( .C1(n14587), .C2(n16106), .A(n14586), .B(n14585), .ZN(
        P1_U3010) );
  NOR2_X1 U17979 ( .A1(n15876), .A2(n20038), .ZN(n14593) );
  NOR3_X1 U17980 ( .A1(n14605), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n14600), .ZN(n14592) );
  INV_X1 U17981 ( .A(n14588), .ZN(n14591) );
  AOI211_X1 U17982 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n14602), .A(
        n14589), .B(n14601), .ZN(n14590) );
  NOR4_X1 U17983 ( .A1(n14593), .A2(n14592), .A3(n14591), .A4(n14590), .ZN(
        n14594) );
  OAI21_X1 U17984 ( .B1(n14595), .B2(n16106), .A(n14594), .ZN(P1_U3011) );
  NOR2_X1 U17985 ( .A1(n14597), .A2(n14596), .ZN(n14598) );
  XNOR2_X1 U17986 ( .A(n14599), .B(n14598), .ZN(n15946) );
  NOR2_X1 U17987 ( .A1(n14601), .A2(n14600), .ZN(n14604) );
  INV_X1 U17988 ( .A(n14602), .ZN(n14603) );
  AOI22_X1 U17989 ( .A1(n14604), .A2(n14603), .B1(n10704), .B2(
        P1_REIP_REG_19__SCAN_IN), .ZN(n14607) );
  OR2_X1 U17990 ( .A1(n14605), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14606) );
  OAI211_X1 U17991 ( .C1(n15896), .C2(n20038), .A(n14607), .B(n14606), .ZN(
        n14608) );
  INV_X1 U17992 ( .A(n14608), .ZN(n14609) );
  OAI21_X1 U17993 ( .B1(n15946), .B2(n16106), .A(n14609), .ZN(P1_U3012) );
  INV_X1 U17994 ( .A(n16013), .ZN(n16020) );
  NOR2_X1 U17995 ( .A1(n16020), .A2(n14610), .ZN(n14612) );
  INV_X1 U17996 ( .A(n14612), .ZN(n16028) );
  NOR2_X1 U17997 ( .A1(n10501), .A2(n16028), .ZN(n14614) );
  OAI21_X1 U17998 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16009), .A(
        n16037), .ZN(n14611) );
  AOI21_X1 U17999 ( .B1(n14612), .B2(n10501), .A(n14611), .ZN(n16027) );
  INV_X1 U18000 ( .A(n16027), .ZN(n14613) );
  MUX2_X1 U18001 ( .A(n14614), .B(n14613), .S(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .Z(n14618) );
  OAI21_X1 U18002 ( .B1(n14616), .B2(n20038), .A(n14615), .ZN(n14617) );
  AOI211_X1 U18003 ( .C1(n14619), .C2(n20063), .A(n14618), .B(n14617), .ZN(
        n14620) );
  INV_X1 U18004 ( .A(n14620), .ZN(P1_U3015) );
  NAND3_X1 U18005 ( .A1(n14621), .A2(n12741), .A3(n20063), .ZN(n14631) );
  INV_X1 U18006 ( .A(n14622), .ZN(n14626) );
  AOI21_X1 U18007 ( .B1(n14624), .B2(n14623), .A(n14641), .ZN(n14625) );
  AOI211_X1 U18008 ( .C1(n20059), .C2(n14627), .A(n14626), .B(n14625), .ZN(
        n14630) );
  OAI211_X1 U18009 ( .C1(n14628), .C2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n16086), .B(n14641), .ZN(n14629) );
  NAND3_X1 U18010 ( .A1(n14631), .A2(n14630), .A3(n14629), .ZN(P1_U3030) );
  INV_X1 U18011 ( .A(n20590), .ZN(n14633) );
  MUX2_X1 U18012 ( .A(n14633), .B(n14632), .S(n12984), .Z(n14634) );
  OAI21_X1 U18013 ( .B1(n20736), .B2(n12944), .A(n14634), .ZN(n14635) );
  MUX2_X1 U18014 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n14635), .S(
        n20740), .Z(P1_U3476) );
  NOR2_X1 U18015 ( .A1(n14636), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14639) );
  NOR3_X1 U18016 ( .A1(n14637), .A2(n14642), .A3(n14643), .ZN(n14638) );
  AOI211_X1 U18017 ( .C1(n20543), .C2(n14640), .A(n14639), .B(n14638), .ZN(
        n15805) );
  INV_X1 U18018 ( .A(n19877), .ZN(n14659) );
  AOI22_X1 U18019 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n14641), .B2(n10512), .ZN(
        n14652) );
  INV_X1 U18020 ( .A(n14652), .ZN(n14645) );
  NOR2_X1 U18021 ( .A1(n20648), .A2(n20055), .ZN(n14651) );
  NOR3_X1 U18022 ( .A1(n14643), .A2(n14642), .A3(n14657), .ZN(n14644) );
  AOI21_X1 U18023 ( .B1(n14645), .B2(n14651), .A(n14644), .ZN(n14646) );
  OAI21_X1 U18024 ( .B1(n15805), .B2(n14659), .A(n14646), .ZN(n14648) );
  INV_X1 U18025 ( .A(n14647), .ZN(n16117) );
  MUX2_X1 U18026 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14648), .S(
        n16117), .Z(P1_U3473) );
  INV_X1 U18027 ( .A(n14649), .ZN(n14650) );
  INV_X1 U18028 ( .A(n14657), .ZN(n15836) );
  AOI22_X1 U18029 ( .A1(n14652), .A2(n14651), .B1(n14650), .B2(n15836), .ZN(
        n14653) );
  OAI21_X1 U18030 ( .B1(n14654), .B2(n14659), .A(n14653), .ZN(n14655) );
  MUX2_X1 U18031 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14655), .S(
        n16117), .Z(P1_U3472) );
  INV_X1 U18032 ( .A(n14656), .ZN(n14660) );
  OAI22_X1 U18033 ( .A1(n14660), .A2(n14659), .B1(n14658), .B2(n14657), .ZN(
        n14661) );
  MUX2_X1 U18034 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14661), .S(
        n16117), .Z(P1_U3469) );
  NAND4_X1 U18035 ( .A1(n14676), .A2(n18951), .A3(n12901), .A4(n14662), .ZN(
        n14671) );
  INV_X1 U18036 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14663) );
  OAI22_X1 U18037 ( .A1(n14664), .A2(n14742), .B1(n14663), .B2(n18955), .ZN(
        n14665) );
  AOI21_X1 U18038 ( .B1(P2_REIP_REG_31__SCAN_IN), .B2(n18963), .A(n14665), 
        .ZN(n14666) );
  OAI21_X1 U18039 ( .B1(n14667), .B2(n18960), .A(n14666), .ZN(n14668) );
  AOI21_X1 U18040 ( .B1(n14669), .B2(n18958), .A(n14668), .ZN(n14670) );
  OAI211_X1 U18041 ( .C1(n14739), .C2(n18965), .A(n14671), .B(n14670), .ZN(
        P2_U2824) );
  NAND2_X1 U18042 ( .A1(n14673), .A2(n14672), .ZN(n14674) );
  NAND2_X1 U18043 ( .A1(n14675), .A2(n14674), .ZN(n15303) );
  AOI21_X1 U18044 ( .B1(n14677), .B2(n15144), .A(n14676), .ZN(n14678) );
  NAND2_X1 U18045 ( .A1(n14678), .A2(n18951), .ZN(n14690) );
  INV_X1 U18046 ( .A(n14679), .ZN(n14682) );
  INV_X1 U18047 ( .A(n14680), .ZN(n14681) );
  NAND2_X1 U18048 ( .A1(n14682), .A2(n14681), .ZN(n14683) );
  AOI22_X1 U18049 ( .A1(n18963), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18957), .ZN(n14686) );
  NAND2_X1 U18050 ( .A1(n18898), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14685) );
  OAI211_X1 U18051 ( .C1(n15301), .C2(n18960), .A(n14686), .B(n14685), .ZN(
        n14687) );
  AOI21_X1 U18052 ( .B1(n14688), .B2(n18958), .A(n14687), .ZN(n14689) );
  OAI211_X1 U18053 ( .C1(n15303), .C2(n18965), .A(n14690), .B(n14689), .ZN(
        P2_U2826) );
  NOR2_X1 U18054 ( .A1(n14708), .A2(n14691), .ZN(n14692) );
  OR2_X1 U18055 ( .A1(n14693), .A2(n14692), .ZN(n15331) );
  AOI211_X1 U18056 ( .C1(n15154), .C2(n14695), .A(n14694), .B(n19713), .ZN(
        n14696) );
  INV_X1 U18057 ( .A(n14696), .ZN(n14706) );
  NAND2_X1 U18058 ( .A1(n14697), .A2(n14698), .ZN(n14699) );
  NAND2_X1 U18059 ( .A1(n14700), .A2(n14699), .ZN(n15327) );
  AOI22_X1 U18060 ( .A1(P2_REIP_REG_27__SCAN_IN), .A2(n18963), .B1(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n18957), .ZN(n14702) );
  NAND2_X1 U18061 ( .A1(n18898), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14701) );
  OAI211_X1 U18062 ( .C1(n15327), .C2(n18960), .A(n14702), .B(n14701), .ZN(
        n14703) );
  AOI21_X1 U18063 ( .B1(n14704), .B2(n18958), .A(n14703), .ZN(n14705) );
  OAI211_X1 U18064 ( .C1(n15331), .C2(n18965), .A(n14706), .B(n14705), .ZN(
        P2_U2828) );
  AND2_X1 U18065 ( .A1(n14727), .A2(n14707), .ZN(n14709) );
  OR2_X1 U18066 ( .A1(n14709), .A2(n14708), .ZN(n15344) );
  OR2_X1 U18067 ( .A1(n14724), .A2(n14710), .ZN(n14711) );
  NAND2_X1 U18068 ( .A1(n14697), .A2(n14711), .ZN(n15340) );
  INV_X1 U18069 ( .A(n15340), .ZN(n14722) );
  NOR2_X1 U18070 ( .A1(n9940), .A2(n18955), .ZN(n14715) );
  AOI211_X1 U18071 ( .C1(n10103), .C2(n14713), .A(n19713), .B(n14712), .ZN(
        n14714) );
  AOI211_X1 U18072 ( .C1(n18963), .C2(P2_REIP_REG_26__SCAN_IN), .A(n14715), 
        .B(n14714), .ZN(n14716) );
  OAI21_X1 U18073 ( .B1(n18961), .B2(n14717), .A(n14716), .ZN(n14721) );
  AOI211_X1 U18074 ( .C1(P2_EBX_REG_26__SCAN_IN), .C2(n14719), .A(n18941), .B(
        n14718), .ZN(n14720) );
  AOI211_X1 U18075 ( .C1(n14722), .C2(n18907), .A(n14721), .B(n14720), .ZN(
        n14723) );
  OAI21_X1 U18076 ( .B1(n15344), .B2(n18965), .A(n14723), .ZN(P2_U2829) );
  INV_X1 U18077 ( .A(n14724), .ZN(n14725) );
  OAI21_X1 U18078 ( .B1(n15100), .B2(n14726), .A(n14725), .ZN(n15353) );
  INV_X1 U18079 ( .A(n14727), .ZN(n14728) );
  AOI21_X1 U18080 ( .B1(n14729), .B2(n15018), .A(n14728), .ZN(n15356) );
  NAND2_X1 U18081 ( .A1(n15356), .A2(n18902), .ZN(n14732) );
  INV_X1 U18082 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19774) );
  OAI22_X1 U18083 ( .A1(n18923), .A2(n19774), .B1(n15172), .B2(n18955), .ZN(
        n14730) );
  AOI21_X1 U18084 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n18898), .A(n14730), .ZN(
        n14731) );
  OAI211_X1 U18085 ( .C1(n15353), .C2(n18960), .A(n14732), .B(n14731), .ZN(
        n14736) );
  AOI211_X1 U18086 ( .C1(n14734), .C2(n15170), .A(n19713), .B(n14733), .ZN(
        n14735) );
  AOI211_X1 U18087 ( .C1(n18958), .C2(n14737), .A(n14736), .B(n14735), .ZN(
        n14738) );
  INV_X1 U18088 ( .A(n14738), .ZN(P2_U2830) );
  INV_X1 U18089 ( .A(n14739), .ZN(n14740) );
  NAND2_X1 U18090 ( .A1(n14740), .A2(n14743), .ZN(n14741) );
  OAI21_X1 U18091 ( .B1(n14743), .B2(n14742), .A(n14741), .ZN(P2_U2856) );
  AOI22_X1 U18092 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n11963), .B1(
        n11964), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14745) );
  NAND2_X1 U18093 ( .A1(n14861), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n14744) );
  AND2_X1 U18094 ( .A1(n14745), .A2(n14744), .ZN(n14749) );
  AOI22_X1 U18095 ( .A1(n14862), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14748) );
  AOI22_X1 U18096 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12057), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14747) );
  AOI22_X1 U18097 ( .A1(n12056), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14746) );
  NAND4_X1 U18098 ( .A1(n14749), .A2(n14748), .A3(n14747), .A4(n14746), .ZN(
        n14755) );
  AOI22_X1 U18099 ( .A1(n12053), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14867), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14753) );
  AOI22_X1 U18100 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n12026), .B1(
        n12027), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14752) );
  AOI22_X1 U18101 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12003), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14751) );
  NAND2_X1 U18102 ( .A1(n14868), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n14750) );
  NAND4_X1 U18103 ( .A1(n14753), .A2(n14752), .A3(n14751), .A4(n14750), .ZN(
        n14754) );
  OR2_X1 U18104 ( .A1(n14755), .A2(n14754), .ZN(n14877) );
  AOI22_X1 U18105 ( .A1(n14787), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14966), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14764) );
  NAND2_X1 U18106 ( .A1(n14756), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n14760) );
  OR2_X1 U18107 ( .A1(n14758), .A2(n14757), .ZN(n14973) );
  NAND2_X1 U18108 ( .A1(n14967), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14759) );
  AND3_X1 U18109 ( .A1(n14760), .A2(n14973), .A3(n14759), .ZN(n14763) );
  AOI22_X1 U18110 ( .A1(n14968), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14972), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14762) );
  AOI22_X1 U18111 ( .A1(n14903), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11946), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14761) );
  NAND4_X1 U18112 ( .A1(n14764), .A2(n14763), .A3(n14762), .A4(n14761), .ZN(
        n14772) );
  AOI22_X1 U18113 ( .A1(n14787), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14971), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14770) );
  NAND2_X1 U18114 ( .A1(n14966), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n14766) );
  INV_X1 U18115 ( .A(n14973), .ZN(n14938) );
  NAND2_X1 U18116 ( .A1(n14967), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n14765) );
  AND3_X1 U18117 ( .A1(n14766), .A2(n14938), .A3(n14765), .ZN(n14769) );
  AOI22_X1 U18118 ( .A1(n14968), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14972), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14768) );
  AOI22_X1 U18119 ( .A1(n14903), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11946), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14767) );
  NAND4_X1 U18120 ( .A1(n14770), .A2(n14769), .A3(n14768), .A4(n14767), .ZN(
        n14771) );
  AND2_X1 U18121 ( .A1(n14772), .A2(n14771), .ZN(n14888) );
  AND2_X1 U18122 ( .A1(n14877), .A2(n14888), .ZN(n14876) );
  INV_X1 U18123 ( .A(n14876), .ZN(n14886) );
  AOI22_X1 U18124 ( .A1(n14787), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14966), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14778) );
  AOI22_X1 U18125 ( .A1(n14968), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14972), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14777) );
  AOI22_X1 U18126 ( .A1(n14971), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14903), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14776) );
  NAND2_X1 U18127 ( .A1(n14967), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n14774) );
  NAND2_X1 U18128 ( .A1(n11946), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n14773) );
  AND3_X1 U18129 ( .A1(n14774), .A2(n14973), .A3(n14773), .ZN(n14775) );
  NAND4_X1 U18130 ( .A1(n14778), .A2(n14777), .A3(n14776), .A4(n14775), .ZN(
        n14786) );
  AOI22_X1 U18131 ( .A1(n14787), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14966), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14784) );
  AOI22_X1 U18132 ( .A1(n14968), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14972), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14783) );
  AOI22_X1 U18133 ( .A1(n14971), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14903), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14782) );
  NAND2_X1 U18134 ( .A1(n14967), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n14780) );
  NAND2_X1 U18135 ( .A1(n11946), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n14779) );
  AND3_X1 U18136 ( .A1(n14780), .A2(n14938), .A3(n14779), .ZN(n14781) );
  NAND4_X1 U18137 ( .A1(n14784), .A2(n14783), .A3(n14782), .A4(n14781), .ZN(
        n14785) );
  NAND2_X1 U18138 ( .A1(n14786), .A2(n14785), .ZN(n14887) );
  NOR2_X1 U18139 ( .A1(n14886), .A2(n14887), .ZN(n14890) );
  AOI22_X1 U18140 ( .A1(n14787), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14966), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14793) );
  AOI22_X1 U18141 ( .A1(n14968), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14972), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14792) );
  AOI22_X1 U18142 ( .A1(n14756), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14903), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14791) );
  NAND2_X1 U18143 ( .A1(n14967), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14789) );
  NAND2_X1 U18144 ( .A1(n11946), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n14788) );
  AND3_X1 U18145 ( .A1(n14789), .A2(n14973), .A3(n14788), .ZN(n14790) );
  NAND4_X1 U18146 ( .A1(n14793), .A2(n14792), .A3(n14791), .A4(n14790), .ZN(
        n14801) );
  AOI22_X1 U18147 ( .A1(n14787), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14966), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14799) );
  AOI22_X1 U18148 ( .A1(n14968), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14972), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14798) );
  AOI22_X1 U18149 ( .A1(n14971), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14903), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14797) );
  NAND2_X1 U18150 ( .A1(n14967), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n14795) );
  NAND2_X1 U18151 ( .A1(n11946), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n14794) );
  AND3_X1 U18152 ( .A1(n14795), .A2(n14938), .A3(n14794), .ZN(n14796) );
  NAND4_X1 U18153 ( .A1(n14799), .A2(n14798), .A3(n14797), .A4(n14796), .ZN(
        n14800) );
  AND2_X1 U18154 ( .A1(n14801), .A2(n14800), .ZN(n14891) );
  NAND2_X1 U18155 ( .A1(n14890), .A2(n14891), .ZN(n14889) );
  AOI22_X1 U18156 ( .A1(n14787), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14966), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14807) );
  AOI22_X1 U18157 ( .A1(n14968), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14972), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14806) );
  AOI22_X1 U18158 ( .A1(n14756), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14903), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14805) );
  NAND2_X1 U18159 ( .A1(n14967), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n14803) );
  NAND2_X1 U18160 ( .A1(n11946), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n14802) );
  AND3_X1 U18161 ( .A1(n14803), .A2(n14973), .A3(n14802), .ZN(n14804) );
  NAND4_X1 U18162 ( .A1(n14807), .A2(n14806), .A3(n14805), .A4(n14804), .ZN(
        n14815) );
  AOI22_X1 U18163 ( .A1(n14787), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14966), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14813) );
  AOI22_X1 U18164 ( .A1(n14968), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14972), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14812) );
  AOI22_X1 U18165 ( .A1(n14971), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14903), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14811) );
  NAND2_X1 U18166 ( .A1(n14967), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n14809) );
  NAND2_X1 U18167 ( .A1(n11946), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n14808) );
  AND3_X1 U18168 ( .A1(n14809), .A2(n14938), .A3(n14808), .ZN(n14810) );
  NAND4_X1 U18169 ( .A1(n14813), .A2(n14812), .A3(n14811), .A4(n14810), .ZN(
        n14814) );
  NAND2_X1 U18170 ( .A1(n14815), .A2(n14814), .ZN(n14897) );
  AOI21_X1 U18171 ( .B1(n14889), .B2(n14897), .A(n14885), .ZN(n14816) );
  OR2_X1 U18172 ( .A1(n14889), .A2(n14897), .ZN(n14900) );
  AOI22_X1 U18173 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n12144), .B1(
        n12053), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14823) );
  NAND2_X1 U18174 ( .A1(n12004), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n14819) );
  NAND2_X1 U18175 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n14818) );
  NAND2_X1 U18176 ( .A1(n11963), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n14817) );
  AND3_X1 U18177 ( .A1(n14819), .A2(n14818), .A3(n14817), .ZN(n14822) );
  AOI22_X1 U18178 ( .A1(n14862), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14861), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14821) );
  AOI22_X1 U18179 ( .A1(n12056), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12057), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14820) );
  NAND4_X1 U18180 ( .A1(n14823), .A2(n14822), .A3(n14821), .A4(n14820), .ZN(
        n14829) );
  AOI22_X1 U18181 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n14867), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14827) );
  AOI22_X1 U18182 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n12026), .B1(
        n12027), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14826) );
  AOI22_X1 U18183 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12003), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14825) );
  NAND2_X1 U18184 ( .A1(n14868), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n14824) );
  NAND4_X1 U18185 ( .A1(n14827), .A2(n14826), .A3(n14825), .A4(n14824), .ZN(
        n14828) );
  NOR2_X1 U18186 ( .A1(n14829), .A2(n14828), .ZN(n15051) );
  NOR2_X2 U18187 ( .A1(n14830), .A2(n15051), .ZN(n15043) );
  AOI22_X1 U18188 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12053), .B1(
        n12144), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14837) );
  NAND2_X1 U18189 ( .A1(n12004), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n14833) );
  NAND2_X1 U18190 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n14832) );
  NAND2_X1 U18191 ( .A1(n11963), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14831) );
  AND3_X1 U18192 ( .A1(n14833), .A2(n14832), .A3(n14831), .ZN(n14836) );
  AOI22_X1 U18193 ( .A1(n14862), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n14861), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14835) );
  AOI22_X1 U18194 ( .A1(n12056), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12057), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14834) );
  NAND4_X1 U18195 ( .A1(n14837), .A2(n14836), .A3(n14835), .A4(n14834), .ZN(
        n14843) );
  AOI22_X1 U18196 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n14867), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14841) );
  AOI22_X1 U18197 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n12026), .B1(
        n12027), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14840) );
  AOI22_X1 U18198 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12003), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14839) );
  NAND2_X1 U18199 ( .A1(n14868), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n14838) );
  NAND4_X1 U18200 ( .A1(n14841), .A2(n14840), .A3(n14839), .A4(n14838), .ZN(
        n14842) );
  NOR2_X1 U18201 ( .A1(n14843), .A2(n14842), .ZN(n15044) );
  AOI22_X1 U18202 ( .A1(n12053), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12144), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14851) );
  NAND2_X1 U18203 ( .A1(n12004), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n14847) );
  NAND2_X1 U18204 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n14846) );
  NAND2_X1 U18205 ( .A1(n11963), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n14845) );
  AND3_X1 U18206 ( .A1(n14847), .A2(n14846), .A3(n14845), .ZN(n14850) );
  AOI22_X1 U18207 ( .A1(n14862), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14861), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14849) );
  AOI22_X1 U18208 ( .A1(n12056), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12057), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14848) );
  NAND4_X1 U18209 ( .A1(n14851), .A2(n14850), .A3(n14849), .A4(n14848), .ZN(
        n14857) );
  AOI22_X1 U18210 ( .A1(n14867), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14855) );
  AOI22_X1 U18211 ( .A1(n12026), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12027), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14854) );
  AOI22_X1 U18212 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14853) );
  NAND2_X1 U18213 ( .A1(n14868), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n14852) );
  NAND4_X1 U18214 ( .A1(n14855), .A2(n14854), .A3(n14853), .A4(n14852), .ZN(
        n14856) );
  OR2_X1 U18215 ( .A1(n14857), .A2(n14856), .ZN(n15036) );
  AOI22_X1 U18216 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n12144), .B1(
        n12053), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14866) );
  NAND2_X1 U18217 ( .A1(n12004), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n14860) );
  NAND2_X1 U18218 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n14859) );
  NAND2_X1 U18219 ( .A1(n11963), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n14858) );
  AND3_X1 U18220 ( .A1(n14860), .A2(n14859), .A3(n14858), .ZN(n14865) );
  AOI22_X1 U18221 ( .A1(n14862), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14861), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14864) );
  AOI22_X1 U18222 ( .A1(n12056), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12057), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14863) );
  NAND4_X1 U18223 ( .A1(n14866), .A2(n14865), .A3(n14864), .A4(n14863), .ZN(
        n14874) );
  AOI22_X1 U18224 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n11980), .B1(
        n14867), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14872) );
  AOI22_X1 U18225 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n12026), .B1(
        n12027), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14871) );
  AOI22_X1 U18226 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12003), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14870) );
  NAND2_X1 U18227 ( .A1(n14868), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n14869) );
  NAND4_X1 U18228 ( .A1(n14872), .A2(n14871), .A3(n14870), .A4(n14869), .ZN(
        n14873) );
  NOR2_X1 U18229 ( .A1(n14874), .A2(n14873), .ZN(n15032) );
  NAND2_X1 U18230 ( .A1(n14876), .A2(n14935), .ZN(n14881) );
  INV_X1 U18231 ( .A(n14877), .ZN(n14879) );
  NAND2_X1 U18232 ( .A1(n19865), .A2(n14888), .ZN(n14878) );
  NAND2_X1 U18233 ( .A1(n14879), .A2(n14878), .ZN(n14880) );
  XNOR2_X2 U18234 ( .A(n15031), .B(n9709), .ZN(n15025) );
  INV_X1 U18235 ( .A(n14888), .ZN(n14882) );
  NOR2_X1 U18236 ( .A1(n14935), .A2(n14882), .ZN(n15024) );
  AOI211_X1 U18237 ( .C1(n14887), .C2(n14886), .A(n14885), .B(n14890), .ZN(
        n15015) );
  NOR2_X1 U18238 ( .A1(n19865), .A2(n14887), .ZN(n15017) );
  OAI211_X1 U18239 ( .C1(n14890), .C2(n14891), .A(n14889), .B(n14916), .ZN(
        n14894) );
  INV_X1 U18240 ( .A(n14891), .ZN(n14892) );
  NOR2_X1 U18241 ( .A1(n14935), .A2(n14892), .ZN(n15008) );
  INV_X1 U18242 ( .A(n14897), .ZN(n14898) );
  NAND2_X1 U18243 ( .A1(n11798), .A2(n14898), .ZN(n15003) );
  AOI21_X2 U18244 ( .B1(n9700), .B2(n14899), .A(n15002), .ZN(n14919) );
  INV_X1 U18245 ( .A(n14900), .ZN(n14917) );
  AOI22_X1 U18246 ( .A1(n14787), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14966), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14907) );
  NAND2_X1 U18247 ( .A1(n14971), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n14902) );
  NAND2_X1 U18248 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n14901) );
  AND3_X1 U18249 ( .A1(n14902), .A2(n14938), .A3(n14901), .ZN(n14906) );
  AOI22_X1 U18250 ( .A1(n14967), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14972), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14905) );
  AOI22_X1 U18251 ( .A1(n14903), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11946), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14904) );
  NAND4_X1 U18252 ( .A1(n14907), .A2(n14906), .A3(n14905), .A4(n14904), .ZN(
        n14915) );
  AOI22_X1 U18253 ( .A1(n14787), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14966), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14913) );
  AOI22_X1 U18254 ( .A1(n14968), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14967), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14912) );
  AOI22_X1 U18255 ( .A1(n14971), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14903), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14911) );
  NAND2_X1 U18256 ( .A1(n11946), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n14909) );
  NAND2_X1 U18257 ( .A1(n14972), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n14908) );
  AND3_X1 U18258 ( .A1(n14909), .A2(n14908), .A3(n14973), .ZN(n14910) );
  NAND4_X1 U18259 ( .A1(n14913), .A2(n14912), .A3(n14911), .A4(n14910), .ZN(
        n14914) );
  AND2_X1 U18260 ( .A1(n14915), .A2(n14914), .ZN(n14920) );
  NAND2_X1 U18261 ( .A1(n14917), .A2(n14920), .ZN(n14991) );
  OAI211_X1 U18262 ( .C1(n14917), .C2(n14920), .A(n14916), .B(n14991), .ZN(
        n14918) );
  NAND2_X1 U18263 ( .A1(n11798), .A2(n14920), .ZN(n14998) );
  AOI22_X1 U18264 ( .A1(n14787), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14966), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14926) );
  AOI22_X1 U18265 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14972), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14925) );
  AOI22_X1 U18266 ( .A1(n14756), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14903), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14924) );
  NAND2_X1 U18267 ( .A1(n14967), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n14922) );
  NAND2_X1 U18268 ( .A1(n11946), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n14921) );
  AND3_X1 U18269 ( .A1(n14922), .A2(n14973), .A3(n14921), .ZN(n14923) );
  NAND4_X1 U18270 ( .A1(n14926), .A2(n14925), .A3(n14924), .A4(n14923), .ZN(
        n14934) );
  AOI22_X1 U18271 ( .A1(n14787), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14966), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14932) );
  AOI22_X1 U18272 ( .A1(n14968), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14972), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14931) );
  AOI22_X1 U18273 ( .A1(n14971), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14903), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14930) );
  NAND2_X1 U18274 ( .A1(n14967), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n14928) );
  NAND2_X1 U18275 ( .A1(n11946), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n14927) );
  AND3_X1 U18276 ( .A1(n14928), .A2(n14938), .A3(n14927), .ZN(n14929) );
  NAND4_X1 U18277 ( .A1(n14932), .A2(n14931), .A3(n14930), .A4(n14929), .ZN(
        n14933) );
  AND2_X1 U18278 ( .A1(n14934), .A2(n14933), .ZN(n14992) );
  INV_X1 U18279 ( .A(n14991), .ZN(n14937) );
  AND2_X1 U18280 ( .A1(n14935), .A2(n14992), .ZN(n14936) );
  AND2_X1 U18281 ( .A1(n14937), .A2(n14936), .ZN(n14956) );
  INV_X1 U18282 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14940) );
  NAND2_X1 U18283 ( .A1(n14971), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n14939) );
  OAI211_X1 U18284 ( .C1(n14941), .C2(n14940), .A(n14939), .B(n14938), .ZN(
        n14942) );
  INV_X1 U18285 ( .A(n14942), .ZN(n14946) );
  AOI22_X1 U18286 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14967), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14945) );
  AOI22_X1 U18287 ( .A1(n14787), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11946), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14944) );
  AOI22_X1 U18288 ( .A1(n14966), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14903), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14943) );
  NAND4_X1 U18289 ( .A1(n14946), .A2(n14945), .A3(n14944), .A4(n14943), .ZN(
        n14954) );
  AOI22_X1 U18290 ( .A1(n14787), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14966), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14952) );
  AOI22_X1 U18291 ( .A1(n14967), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14972), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14951) );
  AOI22_X1 U18292 ( .A1(n14756), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14903), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14950) );
  NAND2_X1 U18293 ( .A1(n14968), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n14948) );
  NAND2_X1 U18294 ( .A1(n11946), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n14947) );
  AND3_X1 U18295 ( .A1(n14948), .A2(n14973), .A3(n14947), .ZN(n14949) );
  NAND4_X1 U18296 ( .A1(n14952), .A2(n14951), .A3(n14950), .A4(n14949), .ZN(
        n14953) );
  AND2_X1 U18297 ( .A1(n14954), .A2(n14953), .ZN(n14955) );
  NAND2_X1 U18298 ( .A1(n14956), .A2(n14955), .ZN(n14957) );
  OAI21_X1 U18299 ( .B1(n14956), .B2(n14955), .A(n14957), .ZN(n14987) );
  INV_X1 U18300 ( .A(n14957), .ZN(n14958) );
  AOI22_X1 U18301 ( .A1(n14787), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14971), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14961) );
  AOI22_X1 U18302 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14972), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14960) );
  NAND2_X1 U18303 ( .A1(n14961), .A2(n14960), .ZN(n14980) );
  INV_X1 U18304 ( .A(n11946), .ZN(n14965) );
  INV_X1 U18305 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14964) );
  AOI22_X1 U18306 ( .A1(n14966), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14903), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14963) );
  AOI21_X1 U18307 ( .B1(n14967), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n14973), .ZN(n14962) );
  OAI211_X1 U18308 ( .C1(n14965), .C2(n14964), .A(n14963), .B(n14962), .ZN(
        n14979) );
  AOI22_X1 U18309 ( .A1(n14787), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14966), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14970) );
  AOI22_X1 U18310 ( .A1(n14968), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14967), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14969) );
  NAND2_X1 U18311 ( .A1(n14970), .A2(n14969), .ZN(n14978) );
  AOI22_X1 U18312 ( .A1(n14971), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14903), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14976) );
  NAND2_X1 U18313 ( .A1(n14972), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n14975) );
  NAND2_X1 U18314 ( .A1(n11946), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n14974) );
  NAND4_X1 U18315 ( .A1(n14976), .A2(n14975), .A3(n14974), .A4(n14973), .ZN(
        n14977) );
  OAI22_X1 U18316 ( .A1(n14980), .A2(n14979), .B1(n14978), .B2(n14977), .ZN(
        n14981) );
  XNOR2_X1 U18317 ( .A(n14982), .B(n14981), .ZN(n15069) );
  NOR2_X1 U18318 ( .A1(n14983), .A2(n15055), .ZN(n14984) );
  AOI21_X1 U18319 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n15050), .A(n14984), .ZN(
        n14985) );
  OAI21_X1 U18320 ( .B1(n15069), .B2(n15060), .A(n14985), .ZN(P2_U2857) );
  INV_X1 U18321 ( .A(n14986), .ZN(n15071) );
  NAND2_X1 U18322 ( .A1(n14988), .A2(n14987), .ZN(n15070) );
  NAND3_X1 U18323 ( .A1(n15071), .A2(n15047), .A3(n15070), .ZN(n14990) );
  NAND2_X1 U18324 ( .A1(n15050), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14989) );
  OAI211_X1 U18325 ( .C1(n15055), .C2(n15303), .A(n14990), .B(n14989), .ZN(
        P2_U2858) );
  NAND2_X1 U18326 ( .A1(n9600), .A2(n14991), .ZN(n14993) );
  XNOR2_X1 U18327 ( .A(n14993), .B(n14992), .ZN(n15080) );
  NOR2_X1 U18328 ( .A1(n14994), .A2(n15055), .ZN(n14995) );
  AOI21_X1 U18329 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n15050), .A(n14995), .ZN(
        n14996) );
  OAI21_X1 U18330 ( .B1(n15080), .B2(n15060), .A(n14996), .ZN(P2_U2859) );
  AOI21_X1 U18331 ( .B1(n14999), .B2(n14998), .A(n14997), .ZN(n15081) );
  NAND2_X1 U18332 ( .A1(n15081), .A2(n15047), .ZN(n15001) );
  NAND2_X1 U18333 ( .A1(n15055), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15000) );
  OAI211_X1 U18334 ( .C1(n15055), .C2(n15331), .A(n15001), .B(n15000), .ZN(
        P2_U2860) );
  AOI21_X1 U18335 ( .B1(n15004), .B2(n15003), .A(n15002), .ZN(n15090) );
  NAND2_X1 U18336 ( .A1(n15090), .A2(n15047), .ZN(n15006) );
  NAND2_X1 U18337 ( .A1(n15050), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15005) );
  OAI211_X1 U18338 ( .C1(n15344), .C2(n15050), .A(n15006), .B(n15005), .ZN(
        P2_U2861) );
  OAI21_X1 U18339 ( .B1(n15009), .B2(n15008), .A(n15007), .ZN(n15096) );
  NOR2_X1 U18340 ( .A1(n14743), .A2(n15010), .ZN(n15011) );
  AOI21_X1 U18341 ( .B1(n15356), .B2(n14743), .A(n15011), .ZN(n15012) );
  OAI21_X1 U18342 ( .B1(n15096), .B2(n15060), .A(n15012), .ZN(P2_U2862) );
  OAI21_X1 U18343 ( .B1(n15015), .B2(n15014), .A(n15013), .ZN(n15016) );
  XOR2_X1 U18344 ( .A(n15017), .B(n15016), .Z(n15106) );
  OAI21_X1 U18345 ( .B1(n15020), .B2(n15019), .A(n15018), .ZN(n15368) );
  NOR2_X1 U18346 ( .A1(n15368), .A2(n15055), .ZN(n15021) );
  AOI21_X1 U18347 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n15055), .A(n15021), .ZN(
        n15022) );
  OAI21_X1 U18348 ( .B1(n15106), .B2(n15060), .A(n15022), .ZN(P2_U2863) );
  OAI21_X1 U18349 ( .B1(n15025), .B2(n15024), .A(n15023), .ZN(n15112) );
  MUX2_X1 U18350 ( .A(n15379), .B(n11903), .S(n15055), .Z(n15026) );
  OAI21_X1 U18351 ( .B1(n15112), .B2(n15060), .A(n15026), .ZN(P2_U2864) );
  INV_X1 U18352 ( .A(n15027), .ZN(n15030) );
  NAND2_X1 U18353 ( .A1(n9648), .A2(n15028), .ZN(n15029) );
  NAND2_X1 U18354 ( .A1(n15030), .A2(n15029), .ZN(n16159) );
  AOI21_X1 U18355 ( .B1(n15032), .B2(n15035), .A(n14883), .ZN(n16143) );
  NAND2_X1 U18356 ( .A1(n16143), .A2(n15047), .ZN(n15034) );
  NAND2_X1 U18357 ( .A1(n15055), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n15033) );
  OAI211_X1 U18358 ( .C1(n16159), .C2(n15055), .A(n15034), .B(n15033), .ZN(
        P2_U2865) );
  OAI21_X1 U18359 ( .B1(n15046), .B2(n15036), .A(n15035), .ZN(n15117) );
  NOR2_X1 U18360 ( .A1(n15402), .A2(n15055), .ZN(n15037) );
  AOI21_X1 U18361 ( .B1(P2_EBX_REG_21__SCAN_IN), .B2(n15055), .A(n15037), .ZN(
        n15038) );
  OAI21_X1 U18362 ( .B1(n15117), .B2(n15060), .A(n15038), .ZN(P2_U2866) );
  OR2_X1 U18363 ( .A1(n15039), .A2(n15040), .ZN(n15041) );
  NAND2_X1 U18364 ( .A1(n15042), .A2(n15041), .ZN(n18797) );
  AND2_X1 U18365 ( .A1(n15052), .A2(n15044), .ZN(n15045) );
  NOR2_X1 U18366 ( .A1(n15046), .A2(n15045), .ZN(n16148) );
  NAND2_X1 U18367 ( .A1(n16148), .A2(n15047), .ZN(n15049) );
  NAND2_X1 U18368 ( .A1(n15050), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n15048) );
  OAI211_X1 U18369 ( .C1(n18797), .C2(n15050), .A(n15049), .B(n15048), .ZN(
        P2_U2867) );
  INV_X1 U18370 ( .A(n15051), .ZN(n15053) );
  OAI21_X1 U18371 ( .B1(n15054), .B2(n15053), .A(n15052), .ZN(n15124) );
  NAND2_X1 U18372 ( .A1(n15055), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n15059) );
  AOI21_X1 U18373 ( .B1(n15057), .B2(n15056), .A(n15039), .ZN(n18808) );
  NAND2_X1 U18374 ( .A1(n18808), .A2(n14743), .ZN(n15058) );
  OAI211_X1 U18375 ( .C1(n15124), .C2(n15060), .A(n15059), .B(n15058), .ZN(
        P2_U2868) );
  NOR2_X2 U18376 ( .A1(n15065), .A2(n15061), .ZN(n18981) );
  INV_X1 U18377 ( .A(n18993), .ZN(n15062) );
  OAI22_X1 U18378 ( .A1(n15127), .A2(n15062), .B1(n19014), .B2(n19057), .ZN(
        n15063) );
  AOI21_X1 U18379 ( .B1(n18981), .B2(BUF1_REG_30__SCAN_IN), .A(n15063), .ZN(
        n15068) );
  NOR2_X2 U18380 ( .A1(n15065), .A2(n15064), .ZN(n18980) );
  AOI22_X1 U18381 ( .A1(n15066), .A2(n19040), .B1(n18980), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n15067) );
  OAI211_X1 U18382 ( .C1(n15069), .C2(n18984), .A(n15068), .B(n15067), .ZN(
        P2_U2889) );
  NAND3_X1 U18383 ( .A1(n15071), .A2(n19044), .A3(n15070), .ZN(n15076) );
  INV_X1 U18384 ( .A(n15301), .ZN(n15073) );
  OAI22_X1 U18385 ( .A1(n15127), .A2(n18996), .B1(n19014), .B2(n19059), .ZN(
        n15072) );
  AOI21_X1 U18386 ( .B1(n15073), .B2(n19040), .A(n15072), .ZN(n15075) );
  AOI22_X1 U18387 ( .A1(n18981), .A2(BUF1_REG_29__SCAN_IN), .B1(n18980), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n15074) );
  NAND3_X1 U18388 ( .A1(n15076), .A2(n15075), .A3(n15074), .ZN(P2_U2890) );
  OAI22_X1 U18389 ( .A1(n15127), .A2(n18998), .B1(n19014), .B2(n19061), .ZN(
        n15077) );
  AOI21_X1 U18390 ( .B1(n15311), .B2(n19040), .A(n15077), .ZN(n15079) );
  AOI22_X1 U18391 ( .A1(n18981), .A2(BUF1_REG_28__SCAN_IN), .B1(n18980), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n15078) );
  OAI211_X1 U18392 ( .C1(n15080), .C2(n18984), .A(n15079), .B(n15078), .ZN(
        P2_U2891) );
  INV_X1 U18393 ( .A(n15081), .ZN(n15086) );
  INV_X1 U18394 ( .A(n15327), .ZN(n15083) );
  OAI22_X1 U18395 ( .A1(n15127), .A2(n19000), .B1(n19014), .B2(n19063), .ZN(
        n15082) );
  AOI21_X1 U18396 ( .B1(n15083), .B2(n19040), .A(n15082), .ZN(n15085) );
  AOI22_X1 U18397 ( .A1(n18981), .A2(BUF1_REG_27__SCAN_IN), .B1(n18980), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n15084) );
  OAI211_X1 U18398 ( .C1(n15086), .C2(n18984), .A(n15085), .B(n15084), .ZN(
        P2_U2892) );
  AOI22_X1 U18399 ( .A1(n18981), .A2(BUF1_REG_26__SCAN_IN), .B1(n18980), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n15088) );
  INV_X1 U18400 ( .A(n15127), .ZN(n18979) );
  AOI22_X1 U18401 ( .A1(n18979), .A2(n19002), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n19039), .ZN(n15087) );
  OAI211_X1 U18402 ( .C1(n18983), .C2(n15340), .A(n15088), .B(n15087), .ZN(
        n15089) );
  AOI21_X1 U18403 ( .B1(n15090), .B2(n19044), .A(n15089), .ZN(n15091) );
  INV_X1 U18404 ( .A(n15091), .ZN(P2_U2893) );
  INV_X1 U18405 ( .A(n15353), .ZN(n15093) );
  OAI22_X1 U18406 ( .A1(n15127), .A2(n19005), .B1(n19014), .B2(n19067), .ZN(
        n15092) );
  AOI21_X1 U18407 ( .B1(n15093), .B2(n19040), .A(n15092), .ZN(n15095) );
  AOI22_X1 U18408 ( .A1(n18981), .A2(BUF1_REG_25__SCAN_IN), .B1(n18980), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n15094) );
  OAI211_X1 U18409 ( .C1(n15096), .C2(n18984), .A(n15095), .B(n15094), .ZN(
        P2_U2894) );
  AND2_X1 U18410 ( .A1(n15098), .A2(n15097), .ZN(n15099) );
  NOR2_X1 U18411 ( .A1(n15100), .A2(n15099), .ZN(n16131) );
  INV_X1 U18412 ( .A(n19009), .ZN(n15102) );
  OAI22_X1 U18413 ( .A1(n15127), .A2(n15102), .B1(n19014), .B2(n15101), .ZN(
        n15103) );
  AOI21_X1 U18414 ( .B1(n19040), .B2(n16131), .A(n15103), .ZN(n15105) );
  AOI22_X1 U18415 ( .A1(n18981), .A2(BUF1_REG_24__SCAN_IN), .B1(n18980), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n15104) );
  OAI211_X1 U18416 ( .C1(n15106), .C2(n18984), .A(n15105), .B(n15104), .ZN(
        P2_U2895) );
  OAI22_X1 U18417 ( .A1(n15127), .A2(n19188), .B1(n19014), .B2(n19070), .ZN(
        n15110) );
  INV_X1 U18418 ( .A(n18981), .ZN(n15131) );
  INV_X1 U18419 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n15108) );
  INV_X1 U18420 ( .A(n18980), .ZN(n15129) );
  INV_X1 U18421 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n15107) );
  OAI22_X1 U18422 ( .A1(n15131), .A2(n15108), .B1(n15129), .B2(n15107), .ZN(
        n15109) );
  AOI211_X1 U18423 ( .C1(n19040), .C2(n15377), .A(n15110), .B(n15109), .ZN(
        n15111) );
  OAI21_X1 U18424 ( .B1(n15112), .B2(n18984), .A(n15111), .ZN(P2_U2896) );
  OAI22_X1 U18425 ( .A1(n15127), .A2(n19178), .B1(n19014), .B2(n19073), .ZN(
        n15115) );
  INV_X1 U18426 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n15113) );
  OAI22_X1 U18427 ( .A1(n15131), .A2(n16376), .B1(n15129), .B2(n15113), .ZN(
        n15114) );
  AOI211_X1 U18428 ( .C1(n19040), .C2(n15399), .A(n15115), .B(n15114), .ZN(
        n15116) );
  OAI21_X1 U18429 ( .B1(n15117), .B2(n18984), .A(n15116), .ZN(P2_U2898) );
  OR2_X1 U18430 ( .A1(n15118), .A2(n15448), .ZN(n15119) );
  NAND2_X1 U18431 ( .A1(n15422), .A2(n15119), .ZN(n15437) );
  INV_X1 U18432 ( .A(n15437), .ZN(n18807) );
  INV_X1 U18433 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n19076) );
  OAI22_X1 U18434 ( .A1(n15127), .A2(n19173), .B1(n19014), .B2(n19076), .ZN(
        n15122) );
  INV_X1 U18435 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n15120) );
  OAI22_X1 U18436 ( .A1(n15131), .A2(n16380), .B1(n15129), .B2(n15120), .ZN(
        n15121) );
  AOI211_X1 U18437 ( .C1(n19040), .C2(n18807), .A(n15122), .B(n15121), .ZN(
        n15123) );
  OAI21_X1 U18438 ( .B1(n15124), .B2(n18984), .A(n15123), .ZN(P2_U2900) );
  NAND2_X1 U18439 ( .A1(n15780), .A2(n15125), .ZN(n15126) );
  NAND2_X1 U18440 ( .A1(n15450), .A2(n15126), .ZN(n15458) );
  INV_X1 U18441 ( .A(n15458), .ZN(n18837) );
  INV_X1 U18442 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n19080) );
  OAI22_X1 U18443 ( .A1(n15127), .A2(n19168), .B1(n19014), .B2(n19080), .ZN(
        n15133) );
  INV_X1 U18444 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n15130) );
  INV_X1 U18445 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n15128) );
  OAI22_X1 U18446 ( .A1(n15131), .A2(n15130), .B1(n15129), .B2(n15128), .ZN(
        n15132) );
  AOI211_X1 U18447 ( .C1(n19040), .C2(n18837), .A(n15133), .B(n15132), .ZN(
        n15134) );
  OAI21_X1 U18448 ( .B1(n15135), .B2(n18984), .A(n15134), .ZN(P2_U2902) );
  NAND2_X1 U18449 ( .A1(n15137), .A2(n15136), .ZN(n15139) );
  XOR2_X1 U18450 ( .A(n15139), .B(n15138), .Z(n15306) );
  AOI21_X1 U18451 ( .B1(n15298), .B2(n15141), .A(n15140), .ZN(n15304) );
  INV_X1 U18452 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19782) );
  OR2_X1 U18453 ( .A1(n18921), .A2(n19782), .ZN(n15300) );
  OAI21_X1 U18454 ( .B1(n19129), .B2(n15142), .A(n15300), .ZN(n15143) );
  AOI21_X1 U18455 ( .B1(n19118), .B2(n15144), .A(n15143), .ZN(n15145) );
  OAI21_X1 U18456 ( .B1(n15303), .B2(n16160), .A(n15145), .ZN(n15146) );
  AOI21_X1 U18457 ( .B1(n15304), .B2(n19123), .A(n15146), .ZN(n15147) );
  OAI21_X1 U18458 ( .B1(n15306), .B2(n16192), .A(n15147), .ZN(P2_U2985) );
  INV_X1 U18459 ( .A(n15148), .ZN(n15149) );
  OAI21_X1 U18460 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15160), .A(
        n15149), .ZN(n15335) );
  OR2_X1 U18461 ( .A1(n15150), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15322) );
  NAND3_X1 U18462 ( .A1(n15322), .A2(n15321), .A3(n19124), .ZN(n15156) );
  INV_X1 U18463 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19778) );
  OR2_X1 U18464 ( .A1(n18921), .A2(n19778), .ZN(n15326) );
  OAI21_X1 U18465 ( .B1(n19129), .B2(n15151), .A(n15326), .ZN(n15153) );
  NOR2_X1 U18466 ( .A1(n15331), .A2(n16160), .ZN(n15152) );
  AOI211_X1 U18467 ( .C1(n19118), .C2(n15154), .A(n15153), .B(n15152), .ZN(
        n15155) );
  OAI211_X1 U18468 ( .C1(n16194), .C2(n15335), .A(n15156), .B(n15155), .ZN(
        P2_U2987) );
  NOR2_X1 U18469 ( .A1(n15157), .A2(n15166), .ZN(n15158) );
  XOR2_X1 U18470 ( .A(n15159), .B(n15158), .Z(n15348) );
  AOI21_X1 U18471 ( .B1(n15336), .B2(n15358), .A(n15160), .ZN(n15346) );
  INV_X1 U18472 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n15161) );
  OR2_X1 U18473 ( .A1(n18921), .A2(n15161), .ZN(n15339) );
  OAI21_X1 U18474 ( .B1(n19129), .B2(n9940), .A(n15339), .ZN(n15162) );
  AOI21_X1 U18475 ( .B1(n19118), .B2(n10103), .A(n15162), .ZN(n15163) );
  OAI21_X1 U18476 ( .B1(n15344), .B2(n16160), .A(n15163), .ZN(n15164) );
  AOI21_X1 U18477 ( .B1(n15346), .B2(n19123), .A(n15164), .ZN(n15165) );
  OAI21_X1 U18478 ( .B1(n15348), .B2(n16192), .A(n15165), .ZN(P2_U2988) );
  NOR2_X1 U18479 ( .A1(n15167), .A2(n15166), .ZN(n15169) );
  XOR2_X1 U18480 ( .A(n15169), .B(n15168), .Z(n15361) );
  NAND2_X1 U18481 ( .A1(n19118), .A2(n15170), .ZN(n15171) );
  NAND2_X1 U18482 ( .A1(n19119), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15352) );
  OAI211_X1 U18483 ( .C1(n19129), .C2(n15172), .A(n15171), .B(n15352), .ZN(
        n15173) );
  AOI21_X1 U18484 ( .B1(n15356), .B2(n19121), .A(n15173), .ZN(n15175) );
  NAND2_X1 U18485 ( .A1(n15180), .A2(n15349), .ZN(n15357) );
  NAND3_X1 U18486 ( .A1(n15358), .A2(n19123), .A3(n15357), .ZN(n15174) );
  OAI211_X1 U18487 ( .C1(n15361), .C2(n16192), .A(n15175), .B(n15174), .ZN(
        P2_U2989) );
  XNOR2_X1 U18488 ( .A(n15177), .B(n15176), .ZN(n15372) );
  INV_X1 U18489 ( .A(n15368), .ZN(n16132) );
  INV_X1 U18490 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19772) );
  NOR2_X1 U18491 ( .A1(n18921), .A2(n19772), .ZN(n15363) );
  AOI21_X1 U18492 ( .B1(n16184), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15363), .ZN(n15178) );
  OAI21_X1 U18493 ( .B1(n16190), .B2(n15179), .A(n15178), .ZN(n15182) );
  OAI21_X1 U18494 ( .B1(n15184), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15180), .ZN(n15362) );
  NOR2_X1 U18495 ( .A1(n15362), .A2(n16194), .ZN(n15181) );
  AOI211_X1 U18496 ( .C1(n19121), .C2(n16132), .A(n15182), .B(n15181), .ZN(
        n15183) );
  OAI21_X1 U18497 ( .B1(n15372), .B2(n16192), .A(n15183), .ZN(P2_U2990) );
  INV_X1 U18498 ( .A(n15184), .ZN(n15185) );
  OAI21_X1 U18499 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n16157), .A(
        n15185), .ZN(n15384) );
  NAND2_X1 U18500 ( .A1(n19119), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n15374) );
  OAI21_X1 U18501 ( .B1(n19129), .B2(n20877), .A(n15374), .ZN(n15187) );
  NOR2_X1 U18502 ( .A1(n15379), .A2(n16160), .ZN(n15186) );
  AOI211_X1 U18503 ( .C1(n19118), .C2(n15188), .A(n15187), .B(n15186), .ZN(
        n15192) );
  XOR2_X1 U18504 ( .A(n15190), .B(n15189), .Z(n15381) );
  NAND2_X1 U18505 ( .A1(n15381), .A2(n19124), .ZN(n15191) );
  OAI211_X1 U18506 ( .C1(n15384), .C2(n16194), .A(n15192), .B(n15191), .ZN(
        P2_U2991) );
  NAND2_X1 U18507 ( .A1(n15193), .A2(n15274), .ZN(n16178) );
  INV_X1 U18508 ( .A(n16178), .ZN(n15195) );
  INV_X1 U18509 ( .A(n16176), .ZN(n15194) );
  OAI21_X2 U18510 ( .B1(n15195), .B2(n15194), .A(n16175), .ZN(n15264) );
  INV_X1 U18511 ( .A(n15262), .ZN(n15196) );
  NOR2_X2 U18512 ( .A1(n15782), .A2(n15783), .ZN(n15781) );
  OAI21_X1 U18513 ( .B1(n15781), .B2(n15198), .A(n15250), .ZN(n15240) );
  AND2_X1 U18514 ( .A1(n15240), .A2(n15237), .ZN(n15229) );
  NAND2_X1 U18515 ( .A1(n15229), .A2(n15227), .ZN(n15213) );
  INV_X1 U18516 ( .A(n15214), .ZN(n15199) );
  AOI21_X1 U18517 ( .B1(n15213), .B2(n15200), .A(n15199), .ZN(n15204) );
  NAND2_X1 U18518 ( .A1(n15202), .A2(n15201), .ZN(n15203) );
  XNOR2_X1 U18519 ( .A(n15204), .B(n15203), .ZN(n15410) );
  AOI21_X1 U18520 ( .B1(n15205), .B2(n15219), .A(n9650), .ZN(n15407) );
  NAND2_X1 U18521 ( .A1(n19119), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15401) );
  OAI21_X1 U18522 ( .B1(n19129), .B2(n15206), .A(n15401), .ZN(n15207) );
  AOI21_X1 U18523 ( .B1(n19118), .B2(n15208), .A(n15207), .ZN(n15209) );
  OAI21_X1 U18524 ( .B1(n15402), .B2(n16160), .A(n15209), .ZN(n15210) );
  AOI21_X1 U18525 ( .B1(n15407), .B2(n19123), .A(n15210), .ZN(n15211) );
  OAI21_X1 U18526 ( .B1(n15410), .B2(n16192), .A(n15211), .ZN(P2_U2993) );
  NAND2_X1 U18527 ( .A1(n15213), .A2(n15212), .ZN(n15217) );
  NAND2_X1 U18528 ( .A1(n15215), .A2(n15214), .ZN(n15216) );
  XNOR2_X1 U18529 ( .A(n15217), .B(n15216), .ZN(n15433) );
  INV_X1 U18530 ( .A(n15219), .ZN(n15220) );
  AOI21_X1 U18531 ( .B1(n15419), .B2(n15218), .A(n15220), .ZN(n15431) );
  NOR2_X1 U18532 ( .A1(n18797), .A2(n16160), .ZN(n15224) );
  NAND2_X1 U18533 ( .A1(n19119), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n15425) );
  NAND2_X1 U18534 ( .A1(n16184), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15221) );
  OAI211_X1 U18535 ( .C1(n16190), .C2(n15222), .A(n15425), .B(n15221), .ZN(
        n15223) );
  AOI211_X1 U18536 ( .C1(n15431), .C2(n19123), .A(n15224), .B(n15223), .ZN(
        n15225) );
  OAI21_X1 U18537 ( .B1(n15433), .B2(n16192), .A(n15225), .ZN(P2_U2994) );
  NAND2_X1 U18538 ( .A1(n15227), .A2(n15226), .ZN(n15231) );
  INV_X1 U18539 ( .A(n15238), .ZN(n15228) );
  NOR2_X1 U18540 ( .A1(n15229), .A2(n15228), .ZN(n15230) );
  XOR2_X1 U18541 ( .A(n15231), .B(n15230), .Z(n15444) );
  NAND2_X1 U18542 ( .A1(n18810), .A2(n19118), .ZN(n15232) );
  NAND2_X1 U18543 ( .A1(n19119), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15435) );
  OAI211_X1 U18544 ( .C1(n19129), .C2(n15233), .A(n15232), .B(n15435), .ZN(
        n15234) );
  AOI21_X1 U18545 ( .B1(n18808), .B2(n19121), .A(n15234), .ZN(n15236) );
  NAND2_X1 U18546 ( .A1(n9811), .A2(n15418), .ZN(n15441) );
  NAND3_X1 U18547 ( .A1(n15441), .A2(n19123), .A3(n15218), .ZN(n15235) );
  OAI211_X1 U18548 ( .C1(n15444), .C2(n16192), .A(n15236), .B(n15235), .ZN(
        P2_U2995) );
  NAND2_X1 U18549 ( .A1(n15238), .A2(n15237), .ZN(n15239) );
  XNOR2_X1 U18550 ( .A(n15240), .B(n15239), .ZN(n15456) );
  INV_X1 U18551 ( .A(n15241), .ZN(n15259) );
  AOI21_X1 U18552 ( .B1(n15447), .B2(n15259), .A(n15242), .ZN(n15454) );
  NOR2_X1 U18553 ( .A1(n18825), .A2(n16160), .ZN(n15245) );
  AOI22_X1 U18554 ( .A1(n16184), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n19119), .ZN(n15243) );
  OAI21_X1 U18555 ( .B1(n18818), .B2(n16190), .A(n15243), .ZN(n15244) );
  AOI211_X1 U18556 ( .C1(n15454), .C2(n19123), .A(n15245), .B(n15244), .ZN(
        n15246) );
  OAI21_X1 U18557 ( .B1(n15456), .B2(n16192), .A(n15246), .ZN(P2_U2996) );
  INV_X1 U18558 ( .A(n15247), .ZN(n15248) );
  NOR2_X1 U18559 ( .A1(n15781), .A2(n15248), .ZN(n15252) );
  NAND2_X1 U18560 ( .A1(n15250), .A2(n15249), .ZN(n15251) );
  XNOR2_X1 U18561 ( .A(n15252), .B(n15251), .ZN(n15474) );
  NOR2_X1 U18562 ( .A1(n18841), .A2(n16190), .ZN(n15255) );
  INV_X1 U18563 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15253) );
  NAND2_X1 U18564 ( .A1(n19119), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15457) );
  OAI21_X1 U18565 ( .B1(n19129), .B2(n15253), .A(n15457), .ZN(n15254) );
  AOI211_X1 U18566 ( .C1(n18838), .C2(n19121), .A(n15255), .B(n15254), .ZN(
        n15261) );
  INV_X1 U18567 ( .A(n15506), .ZN(n15256) );
  INV_X1 U18568 ( .A(n15462), .ZN(n15258) );
  NOR2_X1 U18569 ( .A1(n16179), .A2(n15258), .ZN(n16168) );
  OAI211_X1 U18570 ( .C1(n16168), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n19123), .B(n15259), .ZN(n15260) );
  OAI211_X1 U18571 ( .C1(n15474), .C2(n16192), .A(n15261), .B(n15260), .ZN(
        P2_U2997) );
  NAND2_X1 U18572 ( .A1(n15263), .A2(n15262), .ZN(n15265) );
  XOR2_X1 U18573 ( .A(n15265), .B(n15264), .Z(n16231) );
  NOR2_X1 U18574 ( .A1(n16224), .A2(n16179), .ZN(n16170) );
  AOI21_X1 U18575 ( .B1(n16224), .B2(n16179), .A(n16170), .ZN(n16227) );
  INV_X1 U18576 ( .A(n16227), .ZN(n15267) );
  INV_X1 U18577 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n15266) );
  OAI22_X1 U18578 ( .A1(n16194), .A2(n15267), .B1(n15266), .B2(n18921), .ZN(
        n15270) );
  INV_X1 U18579 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15268) );
  OAI22_X1 U18580 ( .A1(n19129), .A2(n15268), .B1(n16190), .B2(n18854), .ZN(
        n15269) );
  AOI211_X1 U18581 ( .C1(n19121), .C2(n18859), .A(n15270), .B(n15269), .ZN(
        n15271) );
  OAI21_X1 U18582 ( .B1(n16231), .B2(n16192), .A(n15271), .ZN(P2_U2999) );
  NAND2_X1 U18583 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15488), .ZN(
        n15489) );
  INV_X1 U18584 ( .A(n15488), .ZN(n15517) );
  NOR2_X1 U18585 ( .A1(n16233), .A2(n15517), .ZN(n16180) );
  AOI21_X1 U18586 ( .B1(n20796), .B2(n15489), .A(n16180), .ZN(n15272) );
  INV_X1 U18587 ( .A(n15272), .ZN(n15487) );
  INV_X1 U18588 ( .A(n15274), .ZN(n15275) );
  NOR2_X1 U18589 ( .A1(n15276), .A2(n15275), .ZN(n15277) );
  XNOR2_X1 U18590 ( .A(n15273), .B(n15277), .ZN(n15485) );
  OAI22_X1 U18591 ( .A1(n19129), .A2(n18886), .B1(n16190), .B2(n15278), .ZN(
        n15280) );
  NAND2_X1 U18592 ( .A1(n19119), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n15479) );
  OAI21_X1 U18593 ( .B1(n18881), .B2(n16160), .A(n15479), .ZN(n15279) );
  AOI211_X1 U18594 ( .C1(n15485), .C2(n19124), .A(n15280), .B(n15279), .ZN(
        n15281) );
  OAI21_X1 U18595 ( .B1(n15487), .B2(n16194), .A(n15281), .ZN(P2_U3001) );
  INV_X1 U18596 ( .A(n15282), .ZN(n15284) );
  NOR2_X1 U18597 ( .A1(n15284), .A2(n15283), .ZN(n15285) );
  XNOR2_X1 U18598 ( .A(n15286), .B(n15285), .ZN(n15570) );
  INV_X1 U18599 ( .A(n15546), .ZN(n15291) );
  INV_X1 U18600 ( .A(n15287), .ZN(n15545) );
  OAI21_X1 U18601 ( .B1(n15289), .B2(n15545), .A(n15288), .ZN(n15290) );
  OAI21_X1 U18602 ( .B1(n15291), .B2(n15545), .A(n15290), .ZN(n15568) );
  INV_X1 U18603 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15293) );
  OAI22_X1 U18604 ( .A1(n19129), .A2(n15293), .B1(n16190), .B2(n15292), .ZN(
        n15295) );
  OAI22_X1 U18605 ( .A1(n15565), .A2(n16160), .B1(n18921), .B2(n19743), .ZN(
        n15294) );
  AOI211_X1 U18606 ( .C1(n15568), .C2(n19124), .A(n15295), .B(n15294), .ZN(
        n15296) );
  OAI21_X1 U18607 ( .B1(n15570), .B2(n16194), .A(n15296), .ZN(P2_U3007) );
  NOR2_X1 U18608 ( .A1(n15308), .A2(n15307), .ZN(n15297) );
  NOR2_X1 U18609 ( .A1(n15329), .A2(n15297), .ZN(n15314) );
  INV_X1 U18610 ( .A(n15314), .ZN(n15302) );
  INV_X1 U18611 ( .A(n15308), .ZN(n15324) );
  NAND3_X1 U18612 ( .A1(n15324), .A2(n15307), .A3(n15298), .ZN(n15299) );
  OAI21_X1 U18613 ( .B1(n15306), .B2(n19166), .A(n15305), .ZN(P2_U3017) );
  NOR3_X1 U18614 ( .A1(n15308), .A2(n15307), .A3(n15323), .ZN(n15309) );
  AOI211_X1 U18615 ( .C1(n15311), .C2(n19155), .A(n15310), .B(n15309), .ZN(
        n15312) );
  OAI21_X1 U18616 ( .B1(n15314), .B2(n15313), .A(n15312), .ZN(n15317) );
  NOR2_X1 U18617 ( .A1(n15315), .A2(n19159), .ZN(n15316) );
  NAND3_X1 U18618 ( .A1(n15322), .A2(n15321), .A3(n19131), .ZN(n15334) );
  NAND2_X1 U18619 ( .A1(n15324), .A2(n15323), .ZN(n15325) );
  OAI211_X1 U18620 ( .C1(n15327), .C2(n19136), .A(n15326), .B(n15325), .ZN(
        n15328) );
  AOI21_X1 U18621 ( .B1(n15329), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15328), .ZN(n15330) );
  OAI21_X1 U18622 ( .B1(n15331), .B2(n16248), .A(n15330), .ZN(n15332) );
  INV_X1 U18623 ( .A(n15332), .ZN(n15333) );
  OAI211_X1 U18624 ( .C1(n15335), .C2(n19159), .A(n15334), .B(n15333), .ZN(
        P2_U3019) );
  NAND3_X1 U18625 ( .A1(n15349), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15365), .ZN(n15351) );
  NAND2_X1 U18626 ( .A1(n15350), .A2(n15351), .ZN(n15342) );
  NAND3_X1 U18627 ( .A1(n15337), .A2(n15336), .A3(n15365), .ZN(n15338) );
  OAI211_X1 U18628 ( .C1(n15340), .C2(n19136), .A(n15339), .B(n15338), .ZN(
        n15341) );
  AOI21_X1 U18629 ( .B1(n15342), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15341), .ZN(n15343) );
  OAI21_X1 U18630 ( .B1(n15344), .B2(n16248), .A(n15343), .ZN(n15345) );
  AOI21_X1 U18631 ( .B1(n15346), .B2(n16228), .A(n15345), .ZN(n15347) );
  OAI21_X1 U18632 ( .B1(n15348), .B2(n19166), .A(n15347), .ZN(P2_U3020) );
  NOR2_X1 U18633 ( .A1(n15350), .A2(n15349), .ZN(n15355) );
  OAI211_X1 U18634 ( .C1(n15353), .C2(n19136), .A(n15352), .B(n15351), .ZN(
        n15354) );
  AOI211_X1 U18635 ( .C1(n15356), .C2(n19156), .A(n15355), .B(n15354), .ZN(
        n15360) );
  NAND3_X1 U18636 ( .A1(n15358), .A2(n16228), .A3(n15357), .ZN(n15359) );
  OAI211_X1 U18637 ( .C1(n15361), .C2(n19166), .A(n15360), .B(n15359), .ZN(
        P2_U3021) );
  INV_X1 U18638 ( .A(n15362), .ZN(n15370) );
  AOI21_X1 U18639 ( .B1(n19155), .B2(n16131), .A(n15363), .ZN(n15367) );
  OAI21_X1 U18640 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15365), .A(
        n15364), .ZN(n15366) );
  OAI211_X1 U18641 ( .C1(n15368), .C2(n16248), .A(n15367), .B(n15366), .ZN(
        n15369) );
  AOI21_X1 U18642 ( .B1(n15370), .B2(n16228), .A(n15369), .ZN(n15371) );
  OAI21_X1 U18643 ( .B1(n15372), .B2(n19166), .A(n15371), .ZN(P2_U3022) );
  AOI21_X1 U18644 ( .B1(n15508), .B2(n15373), .A(n15507), .ZN(n15406) );
  NAND2_X1 U18645 ( .A1(n15373), .A2(n15459), .ZN(n15393) );
  XNOR2_X1 U18646 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15375) );
  OAI21_X1 U18647 ( .B1(n15393), .B2(n15375), .A(n15374), .ZN(n15376) );
  AOI21_X1 U18648 ( .B1(n19155), .B2(n15377), .A(n15376), .ZN(n15378) );
  OAI21_X1 U18649 ( .B1(n15379), .B2(n16248), .A(n15378), .ZN(n15380) );
  AOI21_X1 U18650 ( .B1(n15406), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15380), .ZN(n15383) );
  NAND2_X1 U18651 ( .A1(n15381), .A2(n19131), .ZN(n15382) );
  OAI211_X1 U18652 ( .C1(n15384), .C2(n19159), .A(n15383), .B(n15382), .ZN(
        P2_U3023) );
  NAND2_X1 U18653 ( .A1(n9685), .A2(n15386), .ZN(n15387) );
  XNOR2_X1 U18654 ( .A(n15385), .B(n15387), .ZN(n16161) );
  NOR2_X1 U18655 ( .A1(n9650), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16158) );
  OR3_X1 U18656 ( .A1(n16158), .A2(n16157), .A3(n19159), .ZN(n15398) );
  OR2_X1 U18657 ( .A1(n15389), .A2(n15388), .ZN(n15390) );
  AND2_X1 U18658 ( .A1(n15391), .A2(n15390), .ZN(n16142) );
  NAND2_X1 U18659 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19119), .ZN(n15392) );
  OAI21_X1 U18660 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15393), .A(
        n15392), .ZN(n15394) );
  AOI21_X1 U18661 ( .B1(n19155), .B2(n16142), .A(n15394), .ZN(n15395) );
  OAI21_X1 U18662 ( .B1(n16159), .B2(n16248), .A(n15395), .ZN(n15396) );
  AOI21_X1 U18663 ( .B1(n15406), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15396), .ZN(n15397) );
  OAI211_X1 U18664 ( .C1(n16161), .C2(n19166), .A(n15398), .B(n15397), .ZN(
        P2_U3024) );
  NAND2_X1 U18665 ( .A1(n19155), .A2(n15399), .ZN(n15400) );
  OAI211_X1 U18666 ( .C1(n15402), .C2(n16248), .A(n15401), .B(n15400), .ZN(
        n15405) );
  NOR3_X1 U18667 ( .A1(n15505), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15403), .ZN(n15404) );
  AOI211_X1 U18668 ( .C1(n15406), .C2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15405), .B(n15404), .ZN(n15409) );
  NAND2_X1 U18669 ( .A1(n15407), .A2(n16228), .ZN(n15408) );
  OAI211_X1 U18670 ( .C1(n15410), .C2(n19166), .A(n15409), .B(n15408), .ZN(
        P2_U3025) );
  INV_X1 U18671 ( .A(n15508), .ZN(n15411) );
  OR2_X1 U18672 ( .A1(n15412), .A2(n15411), .ZN(n15413) );
  NAND2_X1 U18673 ( .A1(n15552), .A2(n15413), .ZN(n16223) );
  INV_X1 U18674 ( .A(n16223), .ZN(n15416) );
  NAND2_X1 U18675 ( .A1(n15459), .A2(n15414), .ZN(n15446) );
  NOR2_X1 U18676 ( .A1(n15446), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15415) );
  AOI211_X1 U18677 ( .C1(n15417), .C2(n19153), .A(n15416), .B(n15415), .ZN(
        n15445) );
  NOR2_X1 U18678 ( .A1(n15446), .A2(n15447), .ZN(n15420) );
  NAND2_X1 U18679 ( .A1(n15420), .A2(n15418), .ZN(n15434) );
  AOI21_X1 U18680 ( .B1(n15445), .B2(n15434), .A(n15419), .ZN(n15430) );
  NAND3_X1 U18681 ( .A1(n15420), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n15419), .ZN(n15428) );
  NAND2_X1 U18682 ( .A1(n15422), .A2(n15421), .ZN(n15423) );
  AND2_X1 U18683 ( .A1(n15424), .A2(n15423), .ZN(n18795) );
  INV_X1 U18684 ( .A(n15425), .ZN(n15426) );
  AOI21_X1 U18685 ( .B1(n19155), .B2(n18795), .A(n15426), .ZN(n15427) );
  OAI211_X1 U18686 ( .C1(n18797), .C2(n16248), .A(n15428), .B(n15427), .ZN(
        n15429) );
  AOI211_X1 U18687 ( .C1(n15431), .C2(n16228), .A(n15430), .B(n15429), .ZN(
        n15432) );
  OAI21_X1 U18688 ( .B1(n15433), .B2(n19166), .A(n15432), .ZN(P2_U3026) );
  INV_X1 U18689 ( .A(n15445), .ZN(n15440) );
  INV_X1 U18690 ( .A(n15434), .ZN(n15439) );
  NAND2_X1 U18691 ( .A1(n18808), .A2(n19156), .ZN(n15436) );
  OAI211_X1 U18692 ( .C1(n19136), .C2(n15437), .A(n15436), .B(n15435), .ZN(
        n15438) );
  AOI211_X1 U18693 ( .C1(n15440), .C2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15439), .B(n15438), .ZN(n15443) );
  NAND3_X1 U18694 ( .A1(n15441), .A2(n16228), .A3(n15218), .ZN(n15442) );
  OAI211_X1 U18695 ( .C1(n15444), .C2(n19166), .A(n15443), .B(n15442), .ZN(
        P2_U3027) );
  AOI21_X1 U18696 ( .B1(n15447), .B2(n15446), .A(n15445), .ZN(n15453) );
  AOI21_X1 U18697 ( .B1(n15450), .B2(n15449), .A(n15448), .ZN(n18823) );
  AOI22_X1 U18698 ( .A1(n19155), .A2(n18823), .B1(n19119), .B2(
        P2_REIP_REG_18__SCAN_IN), .ZN(n15451) );
  OAI21_X1 U18699 ( .B1(n18825), .B2(n16248), .A(n15451), .ZN(n15452) );
  AOI211_X1 U18700 ( .C1(n15454), .C2(n16228), .A(n15453), .B(n15452), .ZN(
        n15455) );
  OAI21_X1 U18701 ( .B1(n15456), .B2(n19166), .A(n15455), .ZN(P2_U3028) );
  OAI21_X1 U18702 ( .B1(n19136), .B2(n15458), .A(n15457), .ZN(n15464) );
  NAND2_X1 U18703 ( .A1(n15475), .A2(n15459), .ZN(n16232) );
  INV_X1 U18704 ( .A(n16232), .ZN(n15498) );
  NAND2_X1 U18705 ( .A1(n15460), .A2(n15498), .ZN(n16225) );
  OAI21_X1 U18706 ( .B1(n16179), .B2(n19159), .A(n16225), .ZN(n15785) );
  AND3_X1 U18707 ( .A1(n15785), .A2(n15462), .A3(n15461), .ZN(n15463) );
  AOI211_X1 U18708 ( .C1(n18838), .C2(n19156), .A(n15464), .B(n15463), .ZN(
        n15473) );
  NOR2_X1 U18709 ( .A1(n19143), .A2(n16228), .ZN(n15465) );
  OR2_X1 U18710 ( .A1(n16168), .A2(n15465), .ZN(n15469) );
  NAND2_X1 U18711 ( .A1(n15466), .A2(n16224), .ZN(n15467) );
  AND2_X1 U18712 ( .A1(n16223), .A2(n15467), .ZN(n15468) );
  NAND2_X1 U18713 ( .A1(n15469), .A2(n15468), .ZN(n15784) );
  INV_X1 U18714 ( .A(n19153), .ZN(n15470) );
  NOR2_X1 U18715 ( .A1(n15470), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15471) );
  OAI21_X1 U18716 ( .B1(n15784), .B2(n15471), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15472) );
  OAI211_X1 U18717 ( .C1(n15474), .C2(n19166), .A(n15473), .B(n15472), .ZN(
        P2_U3029) );
  AOI21_X1 U18718 ( .B1(n15475), .B2(n15508), .A(n15507), .ZN(n15497) );
  AOI21_X1 U18719 ( .B1(n15498), .B2(n16233), .A(n15497), .ZN(n16234) );
  AOI21_X1 U18720 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15498), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15483) );
  OAI21_X1 U18721 ( .B1(n15478), .B2(n15477), .A(n15476), .ZN(n18997) );
  OAI21_X1 U18722 ( .B1(n19136), .B2(n18997), .A(n15479), .ZN(n15480) );
  AOI21_X1 U18723 ( .B1(n15481), .B2(n19156), .A(n15480), .ZN(n15482) );
  OAI21_X1 U18724 ( .B1(n16234), .B2(n15483), .A(n15482), .ZN(n15484) );
  AOI21_X1 U18725 ( .B1(n15485), .B2(n19131), .A(n15484), .ZN(n15486) );
  OAI21_X1 U18726 ( .B1(n15487), .B2(n19159), .A(n15486), .ZN(P2_U3033) );
  OR2_X1 U18727 ( .A1(n15488), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15490) );
  INV_X1 U18728 ( .A(n16185), .ZN(n15503) );
  XNOR2_X1 U18729 ( .A(n15492), .B(n13850), .ZN(n15493) );
  XNOR2_X1 U18730 ( .A(n15491), .B(n15493), .ZN(n16187) );
  XNOR2_X1 U18731 ( .A(n15494), .B(n15495), .ZN(n18999) );
  INV_X1 U18732 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19752) );
  NOR2_X1 U18733 ( .A1(n19752), .A2(n18921), .ZN(n15496) );
  AOI221_X1 U18734 ( .B1(n15498), .B2(n13850), .C1(n15497), .C2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n15496), .ZN(n15500) );
  NAND2_X1 U18735 ( .A1(n16186), .A2(n19156), .ZN(n15499) );
  OAI211_X1 U18736 ( .C1(n18999), .C2(n19136), .A(n15500), .B(n15499), .ZN(
        n15501) );
  AOI21_X1 U18737 ( .B1(n16187), .B2(n19131), .A(n15501), .ZN(n15502) );
  OAI21_X1 U18738 ( .B1(n15503), .B2(n19159), .A(n15502), .ZN(P2_U3034) );
  OAI21_X1 U18739 ( .B1(n9714), .B2(n15504), .A(n15494), .ZN(n19001) );
  NOR2_X1 U18740 ( .A1(n13994), .A2(n15505), .ZN(n15528) );
  OAI211_X1 U18741 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n15528), .B(n15506), .ZN(
        n15523) );
  INV_X1 U18742 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n15520) );
  AOI21_X1 U18743 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15508), .A(
        n15507), .ZN(n15529) );
  NOR2_X1 U18744 ( .A1(n15510), .A2(n15509), .ZN(n15536) );
  AOI21_X1 U18745 ( .B1(n15536), .B2(n15534), .A(n15511), .ZN(n15516) );
  INV_X1 U18746 ( .A(n15512), .ZN(n15514) );
  NAND2_X1 U18747 ( .A1(n15514), .A2(n15513), .ZN(n15515) );
  XNOR2_X1 U18748 ( .A(n15516), .B(n15515), .ZN(n16193) );
  NOR2_X1 U18749 ( .A1(n15525), .A2(n15527), .ZN(n15524) );
  OAI21_X1 U18750 ( .B1(n15524), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15517), .ZN(n16195) );
  OAI22_X1 U18751 ( .A1(n16193), .A2(n19166), .B1(n19159), .B2(n16195), .ZN(
        n15518) );
  AOI21_X1 U18752 ( .B1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15529), .A(
        n15518), .ZN(n15519) );
  OAI21_X1 U18753 ( .B1(n18921), .B2(n15520), .A(n15519), .ZN(n15521) );
  AOI21_X1 U18754 ( .B1(n19156), .B2(n18903), .A(n15521), .ZN(n15522) );
  OAI211_X1 U18755 ( .C1(n19001), .C2(n19136), .A(n15523), .B(n15522), .ZN(
        P2_U3035) );
  AOI21_X1 U18756 ( .B1(n15527), .B2(n15525), .A(n15524), .ZN(n16200) );
  NAND2_X1 U18757 ( .A1(n16200), .A2(n16228), .ZN(n15542) );
  INV_X1 U18758 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19749) );
  NOR2_X1 U18759 ( .A1(n19749), .A2(n18921), .ZN(n15526) );
  AOI221_X1 U18760 ( .B1(n15529), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), 
        .C1(n15528), .C2(n15527), .A(n15526), .ZN(n15541) );
  XNOR2_X1 U18761 ( .A(n15531), .B(n15530), .ZN(n19004) );
  INV_X1 U18762 ( .A(n19004), .ZN(n15532) );
  AOI22_X1 U18763 ( .A1(n19156), .A2(n16201), .B1(n19155), .B2(n15532), .ZN(
        n15540) );
  NAND2_X1 U18764 ( .A1(n15534), .A2(n15533), .ZN(n15538) );
  NOR2_X1 U18765 ( .A1(n15536), .A2(n15535), .ZN(n15537) );
  XOR2_X1 U18766 ( .A(n15538), .B(n15537), .Z(n16202) );
  NAND2_X1 U18767 ( .A1(n16202), .A2(n19131), .ZN(n15539) );
  NAND4_X1 U18768 ( .A1(n15542), .A2(n15541), .A3(n15540), .A4(n15539), .ZN(
        P2_U3036) );
  XOR2_X1 U18769 ( .A(n15544), .B(n15543), .Z(n16209) );
  INV_X1 U18770 ( .A(n16209), .ZN(n15561) );
  NOR2_X1 U18771 ( .A1(n15546), .A2(n15545), .ZN(n15550) );
  NAND2_X1 U18772 ( .A1(n15548), .A2(n15547), .ZN(n15549) );
  XNOR2_X1 U18773 ( .A(n15550), .B(n15549), .ZN(n16208) );
  NAND2_X1 U18774 ( .A1(n15552), .A2(n15551), .ZN(n15563) );
  OAI21_X1 U18775 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n15553), .ZN(n15554) );
  OAI22_X1 U18776 ( .A1(n15555), .A2(n15563), .B1(n15564), .B2(n15554), .ZN(
        n15559) );
  AOI22_X1 U18777 ( .A1(n19155), .A2(n19007), .B1(n19119), .B2(
        P2_REIP_REG_8__SCAN_IN), .ZN(n15556) );
  OAI21_X1 U18778 ( .B1(n16248), .B2(n15557), .A(n15556), .ZN(n15558) );
  AOI211_X1 U18779 ( .C1(n16208), .C2(n19131), .A(n15559), .B(n15558), .ZN(
        n15560) );
  OAI21_X1 U18780 ( .B1(n15561), .B2(n19159), .A(n15560), .ZN(P2_U3038) );
  NAND2_X1 U18781 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19119), .ZN(n15562) );
  OAI221_X1 U18782 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n15564), .C1(
        n13943), .C2(n15563), .A(n15562), .ZN(n15567) );
  OAI22_X1 U18783 ( .A1(n19012), .A2(n19136), .B1(n16248), .B2(n15565), .ZN(
        n15566) );
  AOI211_X1 U18784 ( .C1(n15568), .C2(n19131), .A(n15567), .B(n15566), .ZN(
        n15569) );
  OAI21_X1 U18785 ( .B1(n15570), .B2(n19159), .A(n15569), .ZN(P2_U3039) );
  INV_X1 U18786 ( .A(n15614), .ZN(n15576) );
  INV_X1 U18787 ( .A(n15587), .ZN(n15608) );
  INV_X1 U18788 ( .A(n12536), .ZN(n15571) );
  NAND2_X1 U18789 ( .A1(n15572), .A2(n15571), .ZN(n15581) );
  INV_X1 U18790 ( .A(n15581), .ZN(n15574) );
  MUX2_X1 U18791 ( .A(n15608), .B(n15574), .S(n15573), .Z(n15575) );
  OAI21_X1 U18792 ( .B1(n16249), .B2(n15576), .A(n15575), .ZN(n16261) );
  AOI22_X1 U18793 ( .A1(n9927), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n15577), .B2(n12901), .ZN(n15584) );
  AOI22_X1 U18794 ( .A1(n16261), .A2(n19710), .B1(P2_STATE2_REG_1__SCAN_IN), 
        .B2(n15584), .ZN(n15578) );
  OAI21_X1 U18795 ( .B1(n15579), .B2(n15616), .A(n15578), .ZN(n15580) );
  MUX2_X1 U18796 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n15580), .S(
        n15617), .Z(P2_U3601) );
  INV_X1 U18797 ( .A(n19710), .ZN(n19799) );
  OAI21_X1 U18798 ( .B1(n11937), .B2(n11936), .A(n15581), .ZN(n15582) );
  OAI21_X1 U18799 ( .B1(n15608), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n15582), .ZN(n15583) );
  AOI21_X1 U18800 ( .B1(n19157), .B2(n15614), .A(n15583), .ZN(n16265) );
  OR2_X1 U18801 ( .A1(n15584), .A2(n12437), .ZN(n15599) );
  OAI21_X1 U18802 ( .B1(n12901), .B2(n19150), .A(n15585), .ZN(n15598) );
  OAI222_X1 U18803 ( .A1(n19814), .A2(n15616), .B1(n19799), .B2(n16265), .C1(
        n15599), .C2(n15598), .ZN(n15586) );
  MUX2_X1 U18804 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15586), .S(
        n15617), .Z(P2_U3600) );
  NOR2_X1 U18805 ( .A1(n16257), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15596) );
  INV_X1 U18806 ( .A(n12546), .ZN(n15607) );
  NAND2_X1 U18807 ( .A1(n15587), .A2(n15607), .ZN(n15604) );
  INV_X1 U18808 ( .A(n16272), .ZN(n15588) );
  OR2_X1 U18809 ( .A1(n16274), .A2(n15588), .ZN(n15605) );
  INV_X1 U18810 ( .A(n11947), .ZN(n15589) );
  NAND2_X1 U18811 ( .A1(n15589), .A2(n11737), .ZN(n15606) );
  NAND2_X1 U18812 ( .A1(n11670), .A2(n15606), .ZN(n15592) );
  NAND2_X1 U18813 ( .A1(n15605), .A2(n15592), .ZN(n15595) );
  NAND2_X1 U18814 ( .A1(n15591), .A2(n15590), .ZN(n15602) );
  INV_X1 U18815 ( .A(n15592), .ZN(n15593) );
  NAND2_X1 U18816 ( .A1(n15602), .A2(n15593), .ZN(n15594) );
  OAI211_X1 U18817 ( .C1(n15596), .C2(n15604), .A(n15595), .B(n15594), .ZN(
        n15597) );
  INV_X1 U18818 ( .A(n15598), .ZN(n15600) );
  OAI222_X1 U18819 ( .A1(n19813), .A2(n15616), .B1(n16259), .B2(n19799), .C1(
        n15600), .C2(n15599), .ZN(n15601) );
  MUX2_X1 U18820 ( .A(n16257), .B(n15601), .S(n15617), .Z(P2_U3599) );
  NAND2_X1 U18821 ( .A1(n15602), .A2(n9604), .ZN(n15603) );
  NAND3_X1 U18822 ( .A1(n15604), .A2(n15603), .A3(n15606), .ZN(n15612) );
  INV_X1 U18823 ( .A(n15605), .ZN(n15610) );
  INV_X1 U18824 ( .A(n15606), .ZN(n15609) );
  OAI22_X1 U18825 ( .A1(n15610), .A2(n15609), .B1(n15608), .B2(n15607), .ZN(
        n15611) );
  MUX2_X1 U18826 ( .A(n15612), .B(n15611), .S(n11637), .Z(n15613) );
  AOI211_X1 U18827 ( .C1(n15615), .C2(n15614), .A(n11980), .B(n15613), .ZN(
        n16256) );
  OAI22_X1 U18828 ( .A1(n19445), .A2(n15616), .B1(n16256), .B2(n19799), .ZN(
        n15618) );
  MUX2_X1 U18829 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15618), .S(
        n15617), .Z(P2_U3596) );
  NAND2_X1 U18830 ( .A1(n19812), .A2(n15642), .ZN(n15619) );
  NAND2_X1 U18831 ( .A1(n19812), .A2(n15620), .ZN(n19800) );
  INV_X1 U18832 ( .A(n15632), .ZN(n15622) );
  NOR2_X1 U18833 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19278) );
  NAND2_X1 U18834 ( .A1(n19278), .A2(n19828), .ZN(n19206) );
  NOR2_X1 U18835 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19206), .ZN(
        n19187) );
  INV_X1 U18836 ( .A(n19187), .ZN(n15641) );
  AND2_X1 U18837 ( .A1(n19648), .A2(n15641), .ZN(n15631) );
  NAND2_X1 U18838 ( .A1(n15622), .A2(n15631), .ZN(n15626) );
  NAND2_X1 U18839 ( .A1(n15629), .A2(n19416), .ZN(n15624) );
  NOR2_X1 U18840 ( .A1(n19812), .A2(n19187), .ZN(n15623) );
  AOI21_X1 U18841 ( .B1(n15624), .B2(n15623), .A(n19650), .ZN(n15625) );
  INV_X1 U18842 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15635) );
  INV_X1 U18843 ( .A(n19702), .ZN(n15627) );
  OAI22_X1 U18844 ( .A1(n19660), .A2(n15627), .B1(n19200), .B2(n15641), .ZN(
        n15628) );
  AOI21_X1 U18845 ( .B1(n19246), .B2(n19657), .A(n15628), .ZN(n15634) );
  OAI21_X1 U18846 ( .B1(n15629), .B2(n19187), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15630) );
  NAND2_X1 U18847 ( .A1(n19191), .A2(n19646), .ZN(n15633) );
  OAI211_X1 U18848 ( .C1(n19195), .C2(n15635), .A(n15634), .B(n15633), .ZN(
        P2_U3048) );
  INV_X1 U18849 ( .A(n19667), .ZN(n19217) );
  OAI22_X1 U18850 ( .A1(n19547), .A2(n15642), .B1(n19217), .B2(n15641), .ZN(
        n15636) );
  AOI21_X1 U18851 ( .B1(n19702), .B2(n19544), .A(n15636), .ZN(n15638) );
  NAND2_X1 U18852 ( .A1(n19191), .A2(n19668), .ZN(n15637) );
  OAI211_X1 U18853 ( .C1(n19195), .C2(n15639), .A(n15638), .B(n15637), .ZN(
        P2_U3050) );
  AOI22_X1 U18854 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19189), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19190), .ZN(n19684) );
  INV_X1 U18855 ( .A(n19684), .ZN(n19621) );
  AOI22_X1 U18856 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19190), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19189), .ZN(n19624) );
  NAND2_X1 U18857 ( .A1(n15640), .A2(n19172), .ZN(n19260) );
  OAI22_X1 U18858 ( .A1(n19624), .A2(n15642), .B1(n15641), .B2(n19260), .ZN(
        n15643) );
  AOI21_X1 U18859 ( .B1(n19702), .B2(n19621), .A(n15643), .ZN(n15645) );
  NOR2_X2 U18860 ( .A1(n19032), .A2(n19650), .ZN(n19680) );
  NAND2_X1 U18861 ( .A1(n19191), .A2(n19680), .ZN(n15644) );
  OAI211_X1 U18862 ( .C1(n19195), .C2(n15646), .A(n15645), .B(n15644), .ZN(
        P2_U3052) );
  INV_X1 U18863 ( .A(n19278), .ZN(n19277) );
  NOR2_X1 U18864 ( .A1(n19479), .A2(n19277), .ZN(n19270) );
  AOI21_X1 U18865 ( .B1(n15651), .B2(n19416), .A(n19270), .ZN(n15649) );
  NOR2_X1 U18866 ( .A1(n19481), .A2(n19277), .ZN(n15652) );
  AOI221_X1 U18867 ( .B1(n19272), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19302), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n15652), .ZN(n15648) );
  MUX2_X1 U18868 ( .A(n15649), .B(n15648), .S(n19812), .Z(n15650) );
  INV_X1 U18869 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15657) );
  AOI22_X1 U18870 ( .A1(n19302), .A2(n19657), .B1(n19272), .B2(n19575), .ZN(
        n15656) );
  OAI21_X1 U18871 ( .B1(n15651), .B2(n19270), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15654) );
  INV_X1 U18872 ( .A(n15652), .ZN(n15653) );
  NAND2_X1 U18873 ( .A1(n15654), .A2(n15653), .ZN(n19271) );
  AOI22_X1 U18874 ( .A1(n19271), .A2(n19646), .B1(n19645), .B2(n19270), .ZN(
        n15655) );
  OAI211_X1 U18875 ( .C1(n19276), .C2(n15657), .A(n15656), .B(n15655), .ZN(
        P2_U3064) );
  NAND3_X1 U18876 ( .A1(n18136), .A2(n18119), .A3(n15658), .ZN(n15659) );
  INV_X1 U18877 ( .A(n17145), .ZN(n17142) );
  INV_X2 U18878 ( .A(n17146), .ZN(n17141) );
  AOI22_X1 U18879 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17053), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15664) );
  AOI22_X1 U18880 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15747), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15663) );
  AOI22_X1 U18881 ( .A1(n17072), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15741), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15662) );
  AOI22_X1 U18882 ( .A1(n16928), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15742), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15661) );
  NAND4_X1 U18883 ( .A1(n15664), .A2(n15663), .A3(n15662), .A4(n15661), .ZN(
        n15670) );
  AOI22_X1 U18884 ( .A1(n17088), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15668) );
  AOI22_X1 U18885 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15667) );
  AOI22_X1 U18886 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15666) );
  AOI22_X1 U18887 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15665) );
  NAND4_X1 U18888 ( .A1(n15668), .A2(n15667), .A3(n15666), .A4(n15665), .ZN(
        n15669) );
  NOR2_X1 U18889 ( .A1(n15670), .A2(n15669), .ZN(n16886) );
  AOI22_X1 U18890 ( .A1(n15741), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15674) );
  AOI22_X1 U18891 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15673) );
  AOI22_X1 U18892 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15672) );
  AOI22_X1 U18893 ( .A1(n17067), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15671) );
  NAND4_X1 U18894 ( .A1(n15674), .A2(n15673), .A3(n15672), .A4(n15671), .ZN(
        n15680) );
  AOI22_X1 U18895 ( .A1(n15747), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15678) );
  AOI22_X1 U18896 ( .A1(n17072), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17088), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15677) );
  AOI22_X1 U18897 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17053), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15676) );
  AOI22_X1 U18898 ( .A1(n16928), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15675) );
  NAND4_X1 U18899 ( .A1(n15678), .A2(n15677), .A3(n15676), .A4(n15675), .ZN(
        n15679) );
  NOR2_X1 U18900 ( .A1(n15680), .A2(n15679), .ZN(n16896) );
  AOI22_X1 U18901 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15684) );
  AOI22_X1 U18902 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15683) );
  AOI22_X1 U18903 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15682) );
  AOI22_X1 U18904 ( .A1(n17067), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15681) );
  NAND4_X1 U18905 ( .A1(n15684), .A2(n15683), .A3(n15682), .A4(n15681), .ZN(
        n15690) );
  AOI22_X1 U18906 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15688) );
  AOI22_X1 U18907 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15741), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15687) );
  AOI22_X1 U18908 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15747), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15686) );
  AOI22_X1 U18909 ( .A1(n17072), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17088), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15685) );
  NAND4_X1 U18910 ( .A1(n15688), .A2(n15687), .A3(n15686), .A4(n15685), .ZN(
        n15689) );
  NOR2_X1 U18911 ( .A1(n15690), .A2(n15689), .ZN(n16907) );
  AOI22_X1 U18912 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15694) );
  AOI22_X1 U18913 ( .A1(n17088), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15693) );
  AOI22_X1 U18914 ( .A1(n17072), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15741), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15692) );
  AOI22_X1 U18915 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15742), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15691) );
  NAND4_X1 U18916 ( .A1(n15694), .A2(n15693), .A3(n15692), .A4(n15691), .ZN(
        n15700) );
  AOI22_X1 U18917 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15698) );
  AOI22_X1 U18918 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15697) );
  AOI22_X1 U18919 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15696) );
  AOI22_X1 U18920 ( .A1(n16928), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n15747), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15695) );
  NAND4_X1 U18921 ( .A1(n15698), .A2(n15697), .A3(n15696), .A4(n15695), .ZN(
        n15699) );
  NOR2_X1 U18922 ( .A1(n15700), .A2(n15699), .ZN(n16906) );
  NOR2_X1 U18923 ( .A1(n16907), .A2(n16906), .ZN(n16902) );
  AOI22_X1 U18924 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17109), .B1(
        n17081), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15710) );
  AOI22_X1 U18925 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17105), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n17088), .ZN(n15709) );
  AOI22_X1 U18926 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17106), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17104), .ZN(n15701) );
  OAI21_X1 U18927 ( .B1(n18107), .B2(n15722), .A(n15701), .ZN(n15707) );
  AOI22_X1 U18928 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17090), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15705) );
  AOI22_X1 U18929 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n9618), .ZN(n15704) );
  AOI22_X1 U18930 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n15747), .ZN(n15703) );
  AOI22_X1 U18931 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n15742), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15702) );
  NAND4_X1 U18932 ( .A1(n15705), .A2(n15704), .A3(n15703), .A4(n15702), .ZN(
        n15706) );
  AOI211_X1 U18933 ( .C1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .C2(n17089), .A(
        n15707), .B(n15706), .ZN(n15708) );
  NAND3_X1 U18934 ( .A1(n15710), .A2(n15709), .A3(n15708), .ZN(n16901) );
  NAND2_X1 U18935 ( .A1(n16902), .A2(n16901), .ZN(n16900) );
  NOR2_X1 U18936 ( .A1(n16896), .A2(n16900), .ZN(n16892) );
  AOI22_X1 U18937 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15720) );
  AOI22_X1 U18938 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15719) );
  AOI22_X1 U18939 ( .A1(n17072), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15711) );
  OAI21_X1 U18940 ( .B1(n16910), .B2(n20794), .A(n15711), .ZN(n15717) );
  AOI22_X1 U18941 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9616), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15715) );
  AOI22_X1 U18942 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15714) );
  AOI22_X1 U18943 ( .A1(n17067), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15713) );
  AOI22_X1 U18944 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17088), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15712) );
  NAND4_X1 U18945 ( .A1(n15715), .A2(n15714), .A3(n15713), .A4(n15712), .ZN(
        n15716) );
  AOI211_X1 U18946 ( .C1(n17117), .C2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A(
        n15717), .B(n15716), .ZN(n15718) );
  NAND3_X1 U18947 ( .A1(n15720), .A2(n15719), .A3(n15718), .ZN(n16891) );
  NAND2_X1 U18948 ( .A1(n16892), .A2(n16891), .ZN(n16890) );
  NOR2_X1 U18949 ( .A1(n16886), .A2(n16890), .ZN(n16885) );
  AOI22_X1 U18950 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15731) );
  AOI22_X1 U18951 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15730) );
  AOI22_X1 U18952 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17088), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15721) );
  OAI21_X1 U18953 ( .B1(n15722), .B2(n20890), .A(n15721), .ZN(n15728) );
  AOI22_X1 U18954 ( .A1(n17107), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9618), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15726) );
  AOI22_X1 U18955 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15725) );
  AOI22_X1 U18956 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15742), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15724) );
  AOI22_X1 U18957 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17090), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15723) );
  NAND4_X1 U18958 ( .A1(n15726), .A2(n15725), .A3(n15724), .A4(n15723), .ZN(
        n15727) );
  AOI211_X1 U18959 ( .C1(n17101), .C2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n15728), .B(n15727), .ZN(n15729) );
  NAND3_X1 U18960 ( .A1(n15731), .A2(n15730), .A3(n15729), .ZN(n15732) );
  NAND2_X1 U18961 ( .A1(n16885), .A2(n15732), .ZN(n16880) );
  OAI21_X1 U18962 ( .B1(n16885), .B2(n15732), .A(n16880), .ZN(n17168) );
  AND2_X1 U18963 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16878) );
  NAND2_X1 U18964 ( .A1(n18136), .A2(n17142), .ZN(n17148) );
  INV_X1 U18965 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n16848) );
  INV_X1 U18966 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n15735) );
  NAND3_X1 U18967 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17134) );
  INV_X1 U18968 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n15734) );
  NAND2_X1 U18969 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .ZN(n17048) );
  NAND4_X1 U18970 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .A4(P3_EBX_REG_4__SCAN_IN), .ZN(n15733) );
  NOR4_X1 U18971 ( .A1(n17064), .A2(n15734), .A3(n17048), .A4(n15733), .ZN(
        n17035) );
  NAND3_X1 U18972 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17136), .A3(n17035), 
        .ZN(n15739) );
  NAND2_X1 U18973 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17005), .ZN(n16979) );
  NAND2_X1 U18974 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16966), .ZN(n16935) );
  NOR2_X1 U18975 ( .A1(n17240), .A2(n16935), .ZN(n16937) );
  NAND2_X1 U18976 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16937), .ZN(n16923) );
  NAND2_X1 U18977 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n16905), .ZN(n16899) );
  NOR2_X1 U18978 ( .A1(n16894), .A2(n16536), .ZN(n16895) );
  NAND2_X1 U18979 ( .A1(n16904), .A2(n16895), .ZN(n15736) );
  NAND2_X1 U18980 ( .A1(n17141), .A2(n15736), .ZN(n16893) );
  OAI21_X1 U18981 ( .B1(n16878), .B2(n17148), .A(n16893), .ZN(n16882) );
  INV_X1 U18982 ( .A(n15736), .ZN(n16887) );
  INV_X1 U18983 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16889) );
  NOR2_X1 U18984 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16889), .ZN(n15737) );
  AOI22_X1 U18985 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16882), .B1(n16887), 
        .B2(n15737), .ZN(n15738) );
  OAI21_X1 U18986 ( .B1(n17141), .B2(n17168), .A(n15738), .ZN(P3_U2675) );
  INV_X1 U18987 ( .A(n15739), .ZN(n15740) );
  OAI21_X1 U18988 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n15740), .A(n17141), .ZN(
        n15754) );
  AOI22_X1 U18989 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15746) );
  AOI22_X1 U18990 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15745) );
  AOI22_X1 U18991 ( .A1(n17072), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15741), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15744) );
  AOI22_X1 U18992 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15742), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15743) );
  NAND4_X1 U18993 ( .A1(n15746), .A2(n15745), .A3(n15744), .A4(n15743), .ZN(
        n15753) );
  AOI22_X1 U18994 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15747), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15751) );
  AOI22_X1 U18995 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17088), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15750) );
  AOI22_X1 U18996 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15749) );
  AOI22_X1 U18997 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9618), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15748) );
  NAND4_X1 U18998 ( .A1(n15751), .A2(n15750), .A3(n15749), .A4(n15748), .ZN(
        n15752) );
  NOR2_X1 U18999 ( .A1(n15753), .A2(n15752), .ZN(n17249) );
  OAI22_X1 U19000 ( .A1(n17032), .A2(n15754), .B1(n17249), .B2(n17141), .ZN(
        P3_U2690) );
  NAND2_X1 U19001 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18280) );
  AOI221_X1 U19002 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18280), .C1(n15756), 
        .C2(n18280), .A(n15755), .ZN(n18095) );
  NOR2_X1 U19003 ( .A1(n15757), .A2(n18575), .ZN(n15758) );
  OAI21_X1 U19004 ( .B1(n15758), .B2(n18445), .A(n18096), .ZN(n18093) );
  AOI22_X1 U19005 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18095), .B1(
        n18093), .B2(n18580), .ZN(P3_U2865) );
  NOR2_X1 U19006 ( .A1(n15759), .A2(n18748), .ZN(n17302) );
  OAI211_X1 U19007 ( .C1(n17302), .C2(n15854), .A(n18536), .B(n18751), .ZN(
        n15760) );
  OAI211_X1 U19008 ( .C1(n15763), .C2(n15762), .A(n15761), .B(n15760), .ZN(
        n18567) );
  NOR2_X1 U19009 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n20828), .ZN(n18100) );
  INV_X1 U19010 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18091) );
  NOR2_X1 U19011 ( .A1(n18091), .A2(n18703), .ZN(n15764) );
  AOI211_X1 U19012 ( .C1(n18745), .C2(n18567), .A(n18100), .B(n15764), .ZN(
        n18730) );
  INV_X1 U19013 ( .A(n18730), .ZN(n18728) );
  AOI21_X1 U19014 ( .B1(n18550), .B2(n18540), .A(n15765), .ZN(n18590) );
  NAND3_X1 U19015 ( .A1(n18728), .A2(n18763), .A3(n18590), .ZN(n15766) );
  OAI21_X1 U19016 ( .B1(n18728), .B2(n18540), .A(n15766), .ZN(P3_U3284) );
  NAND2_X1 U19017 ( .A1(n17564), .A2(n10849), .ZN(n16343) );
  OAI221_X1 U19018 ( .B1(n16345), .B2(n16340), .C1(n16345), .C2(n10849), .A(
        n16343), .ZN(n15767) );
  XNOR2_X1 U19019 ( .A(n16320), .B(n15767), .ZN(n16322) );
  NOR2_X1 U19020 ( .A1(n17964), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16347) );
  OAI21_X1 U19021 ( .B1(n10849), .B2(n16347), .A(n18076), .ZN(n15771) );
  NAND2_X1 U19022 ( .A1(n15768), .A2(n18071), .ZN(n18068) );
  NOR2_X1 U19023 ( .A1(n16339), .A2(n18068), .ZN(n17916) );
  INV_X1 U19024 ( .A(n16318), .ZN(n17780) );
  OAI21_X1 U19025 ( .B1(n16319), .B2(n18079), .A(n15769), .ZN(n15770) );
  AOI21_X1 U19026 ( .B1(n17916), .B2(n16311), .A(n15770), .ZN(n15845) );
  NAND2_X1 U19027 ( .A1(n15771), .A2(n15845), .ZN(n15772) );
  AOI22_X1 U19028 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15772), .B1(
        n9612), .B2(P3_REIP_REG_29__SCAN_IN), .ZN(n15776) );
  INV_X1 U19029 ( .A(n16321), .ZN(n16317) );
  INV_X1 U19030 ( .A(n17995), .ZN(n17953) );
  AOI22_X1 U19031 ( .A1(n18530), .A2(n16318), .B1(n17778), .B2(n17953), .ZN(
        n15774) );
  AOI21_X1 U19032 ( .B1(n15774), .B2(n15773), .A(n18086), .ZN(n15847) );
  NAND3_X1 U19033 ( .A1(n16317), .A2(n15847), .A3(n16320), .ZN(n15775) );
  OAI211_X1 U19034 ( .C1(n16322), .C2(n17998), .A(n15776), .B(n15775), .ZN(
        P3_U2833) );
  OR2_X1 U19035 ( .A1(n15778), .A2(n15777), .ZN(n15779) );
  NAND2_X1 U19036 ( .A1(n15780), .A2(n15779), .ZN(n18982) );
  INV_X1 U19037 ( .A(n18982), .ZN(n18848) );
  AOI22_X1 U19038 ( .A1(n18849), .A2(n19156), .B1(n19155), .B2(n18848), .ZN(
        n15789) );
  AOI21_X1 U19039 ( .B1(n15783), .B2(n15782), .A(n15781), .ZN(n16167) );
  AOI22_X1 U19040 ( .A1(n16167), .A2(n19131), .B1(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15784), .ZN(n15788) );
  NAND3_X1 U19041 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n15786), .A3(
        n15785), .ZN(n15787) );
  NAND2_X1 U19042 ( .A1(P2_REIP_REG_16__SCAN_IN), .A2(n19119), .ZN(n16172) );
  NAND4_X1 U19043 ( .A1(n15789), .A2(n15788), .A3(n15787), .A4(n16172), .ZN(
        P2_U3030) );
  INV_X1 U19044 ( .A(n16142), .ZN(n15790) );
  OAI22_X1 U19045 ( .A1(n16159), .A2(n18965), .B1(n18960), .B2(n15790), .ZN(
        n15791) );
  INV_X1 U19046 ( .A(n15791), .ZN(n15801) );
  AOI211_X1 U19047 ( .C1(n15794), .C2(n15792), .A(n15793), .B(n19713), .ZN(
        n15799) );
  INV_X1 U19048 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15795) );
  OAI222_X1 U19049 ( .A1(n18941), .A2(n15797), .B1(n15796), .B2(n18961), .C1(
        n15795), .C2(n18955), .ZN(n15798) );
  AOI211_X1 U19050 ( .C1(n18963), .C2(P2_REIP_REG_22__SCAN_IN), .A(n15799), 
        .B(n15798), .ZN(n15800) );
  NAND2_X1 U19051 ( .A1(n15801), .A2(n15800), .ZN(P2_U2833) );
  INV_X1 U19052 ( .A(n15802), .ZN(n15813) );
  NOR3_X1 U19053 ( .A1(n15804), .A2(n15803), .A3(n20742), .ZN(n15809) );
  AOI211_X1 U19054 ( .C1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n15809), .A(
        n15806), .B(n15805), .ZN(n15807) );
  INV_X1 U19055 ( .A(n15807), .ZN(n15808) );
  OAI21_X1 U19056 ( .B1(n15809), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15808), .ZN(n15810) );
  AOI222_X1 U19057 ( .A1(n15811), .A2(n20395), .B1(n15811), .B2(n15810), .C1(
        n20395), .C2(n15810), .ZN(n15812) );
  AOI222_X1 U19058 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15813), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15812), .C1(n15813), 
        .C2(n15812), .ZN(n15815) );
  AOI211_X1 U19059 ( .C1(n15815), .C2(n20072), .A(n15814), .B(n15830), .ZN(
        n15823) );
  NOR2_X1 U19060 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(P1_MORE_REG_SCAN_IN), .ZN(
        n15819) );
  AND2_X1 U19061 ( .A1(n15816), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n15818) );
  OAI211_X1 U19062 ( .C1(n15820), .C2(n15819), .A(n15818), .B(n15817), .ZN(
        n15821) );
  INV_X1 U19063 ( .A(n15821), .ZN(n15822) );
  AND2_X1 U19064 ( .A1(n15823), .A2(n15822), .ZN(n15829) );
  INV_X1 U19065 ( .A(n15824), .ZN(n15825) );
  AOI21_X1 U19066 ( .B1(n20759), .B2(n15825), .A(n15834), .ZN(n15826) );
  AOI21_X1 U19067 ( .B1(n15828), .B2(n15827), .A(n15826), .ZN(n16124) );
  OAI21_X1 U19068 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(n15829), .A(n16124), 
        .ZN(n16119) );
  INV_X1 U19069 ( .A(n15829), .ZN(n15835) );
  INV_X1 U19070 ( .A(n15830), .ZN(n15831) );
  NAND3_X1 U19071 ( .A1(n15832), .A2(n15831), .A3(n16122), .ZN(n20734) );
  OAI211_X1 U19072 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20659), .A(n20734), 
        .B(n16118), .ZN(n15833) );
  AOI211_X1 U19073 ( .C1(n15835), .C2(n15834), .A(n15833), .B(n20649), .ZN(
        n15839) );
  NAND2_X1 U19074 ( .A1(n20760), .A2(n15836), .ZN(n15837) );
  AOI21_X1 U19075 ( .B1(n15837), .B2(n16119), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n15838) );
  AOI21_X1 U19076 ( .B1(n16119), .B2(n15839), .A(n15838), .ZN(P1_U3161) );
  NAND2_X1 U19077 ( .A1(n15840), .A2(n9771), .ZN(n15841) );
  XNOR2_X1 U19078 ( .A(n15841), .B(n15843), .ZN(n16316) );
  NOR2_X1 U19079 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15842), .ZN(
        n16312) );
  AOI21_X1 U19080 ( .B1(n15845), .B2(n15844), .A(n15843), .ZN(n15846) );
  AOI21_X1 U19081 ( .B1(n16312), .B2(n15847), .A(n15846), .ZN(n15848) );
  NAND2_X1 U19082 ( .A1(n9612), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16307) );
  OAI211_X1 U19083 ( .C1(n17998), .C2(n16316), .A(n15848), .B(n16307), .ZN(
        P3_U2832) );
  INV_X1 U19084 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20658) );
  INV_X1 U19085 ( .A(HOLD), .ZN(n20668) );
  NOR2_X1 U19086 ( .A1(n20658), .A2(n20668), .ZN(n20655) );
  AOI22_X1 U19087 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n15850) );
  NAND2_X1 U19088 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20759), .ZN(n20662) );
  OAI211_X1 U19089 ( .C1(n20655), .C2(n15850), .A(n15849), .B(n20662), .ZN(
        P1_U3195) );
  AND2_X1 U19090 ( .A1(n19999), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR2_X1 U19091 ( .A1(n19717), .A2(n11587), .ZN(n19709) );
  NAND2_X1 U19092 ( .A1(n19709), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n15852) );
  AOI21_X1 U19093 ( .B1(n19820), .B2(n11587), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15851) );
  AOI21_X1 U19094 ( .B1(n15852), .B2(n15851), .A(n16304), .ZN(P2_U3178) );
  INV_X1 U19095 ( .A(n19848), .ZN(n15853) );
  AOI221_X1 U19096 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16304), .C1(n15853), .C2(
        n16304), .A(n19604), .ZN(n19837) );
  INV_X1 U19097 ( .A(n19837), .ZN(n19838) );
  NOR2_X1 U19098 ( .A1(n16292), .A2(n19838), .ZN(P2_U3047) );
  NAND3_X1 U19099 ( .A1(n15854), .A2(n18536), .A3(n18751), .ZN(n15857) );
  NAND3_X1 U19100 ( .A1(n18101), .A2(n18750), .A3(n15855), .ZN(n15856) );
  NAND2_X1 U19101 ( .A1(n18136), .A2(n17151), .ZN(n17198) );
  INV_X1 U19102 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17375) );
  NAND2_X1 U19103 ( .A1(n15858), .A2(n17151), .ZN(n20931) );
  INV_X1 U19104 ( .A(n20931), .ZN(n17295) );
  AOI22_X1 U19105 ( .A1(n17295), .A2(BUF2_REG_0__SCAN_IN), .B1(n17271), .B2(
        n17763), .ZN(n15859) );
  OAI221_X1 U19106 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17198), .C1(n17375), 
        .C2(n17151), .A(n15859), .ZN(P3_U2735) );
  OAI22_X1 U19107 ( .A1(n15862), .A2(n19950), .B1(n15861), .B2(n15860), .ZN(
        n15863) );
  INV_X1 U19108 ( .A(n15863), .ZN(n15873) );
  INV_X1 U19109 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15865) );
  OAI22_X1 U19110 ( .A1(n15924), .A2(n15865), .B1(n19905), .B2(n15864), .ZN(
        n15866) );
  AOI21_X1 U19111 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n15867), .A(n15866), 
        .ZN(n15872) );
  NOR2_X1 U19112 ( .A1(n15868), .A2(n19976), .ZN(n15869) );
  AOI21_X1 U19113 ( .B1(n15870), .B2(n19942), .A(n15869), .ZN(n15871) );
  NAND3_X1 U19114 ( .A1(n15873), .A2(n15872), .A3(n15871), .ZN(P1_U2819) );
  AOI22_X1 U19115 ( .A1(n19967), .A2(P1_EBX_REG_20__SCAN_IN), .B1(n15874), 
        .B2(n19961), .ZN(n15882) );
  AOI21_X1 U19116 ( .B1(n15875), .B2(n15933), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n15878) );
  OAI22_X1 U19117 ( .A1(n15878), .A2(n15877), .B1(n19976), .B2(n15876), .ZN(
        n15879) );
  AOI21_X1 U19118 ( .B1(n15880), .B2(n19942), .A(n15879), .ZN(n15881) );
  OAI211_X1 U19119 ( .C1(n15883), .C2(n19905), .A(n15882), .B(n15881), .ZN(
        P1_U2820) );
  INV_X1 U19120 ( .A(n15952), .ZN(n15884) );
  AOI21_X1 U19121 ( .B1(n19961), .B2(n15884), .A(n10704), .ZN(n15885) );
  OAI21_X1 U19122 ( .B1(n11318), .B2(n19905), .A(n15885), .ZN(n15890) );
  OAI21_X1 U19123 ( .B1(n15888), .B2(n15887), .A(n15886), .ZN(n15912) );
  INV_X1 U19124 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20698) );
  NOR2_X1 U19125 ( .A1(n15912), .A2(n20698), .ZN(n15889) );
  AOI211_X1 U19126 ( .C1(P1_EBX_REG_19__SCAN_IN), .C2(n19967), .A(n15890), .B(
        n15889), .ZN(n15895) );
  INV_X1 U19127 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20696) );
  NAND3_X1 U19128 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n15905), .A3(n15933), 
        .ZN(n15901) );
  AOI21_X1 U19129 ( .B1(n20698), .B2(n20696), .A(n15901), .ZN(n15892) );
  AOI22_X1 U19130 ( .A1(n15893), .A2(n19942), .B1(n15892), .B2(n15891), .ZN(
        n15894) );
  OAI211_X1 U19131 ( .C1(n19976), .C2(n15896), .A(n15895), .B(n15894), .ZN(
        P1_U2821) );
  OAI22_X1 U19132 ( .A1(n15924), .A2(n15898), .B1(n15897), .B2(n19950), .ZN(
        n15899) );
  AOI211_X1 U19133 ( .C1(n19962), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n10704), .B(n15899), .ZN(n15900) );
  OAI221_X1 U19134 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n15901), .C1(n20696), 
        .C2(n15912), .A(n15900), .ZN(n15902) );
  AOI21_X1 U19135 ( .B1(n15903), .B2(n19942), .A(n15902), .ZN(n15904) );
  OAI21_X1 U19136 ( .B1(n19976), .B2(n16010), .A(n15904), .ZN(P1_U2822) );
  AOI21_X1 U19137 ( .B1(n15905), .B2(n15933), .A(P1_REIP_REG_17__SCAN_IN), 
        .ZN(n15913) );
  OAI22_X1 U19138 ( .A1(n15924), .A2(n15907), .B1(n15906), .B2(n19905), .ZN(
        n15908) );
  AOI211_X1 U19139 ( .C1(n19961), .C2(n15958), .A(n10704), .B(n15908), .ZN(
        n15911) );
  INV_X1 U19140 ( .A(n15909), .ZN(n15959) );
  AOI22_X1 U19141 ( .A1(n15959), .A2(n19942), .B1(n19948), .B2(n16021), .ZN(
        n15910) );
  OAI211_X1 U19142 ( .C1(n15913), .C2(n15912), .A(n15911), .B(n15910), .ZN(
        P1_U2823) );
  AOI22_X1 U19143 ( .A1(n15966), .A2(n19961), .B1(n19948), .B2(n16031), .ZN(
        n15919) );
  AOI22_X1 U19144 ( .A1(n19967), .A2(P1_EBX_REG_15__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n19962), .ZN(n15918) );
  NAND2_X1 U19145 ( .A1(n20691), .A2(n15914), .ZN(n15916) );
  AOI22_X1 U19146 ( .A1(n15967), .A2(n19942), .B1(n15916), .B2(n15915), .ZN(
        n15917) );
  NAND4_X1 U19147 ( .A1(n15919), .A2(n15918), .A3(n15917), .A4(n20036), .ZN(
        P1_U2825) );
  NOR2_X1 U19148 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n15920), .ZN(n15931) );
  AOI22_X1 U19149 ( .A1(n15922), .A2(n19961), .B1(n19948), .B2(n15921), .ZN(
        n15930) );
  NOR2_X1 U19150 ( .A1(n15924), .A2(n15923), .ZN(n15927) );
  OAI21_X1 U19151 ( .B1(n19905), .B2(n15925), .A(n20036), .ZN(n15926) );
  AOI211_X1 U19152 ( .C1(n15928), .C2(n19942), .A(n15927), .B(n15926), .ZN(
        n15929) );
  OAI211_X1 U19153 ( .C1(n15932), .C2(n15931), .A(n15930), .B(n15929), .ZN(
        P1_U2826) );
  AOI21_X1 U19154 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n15933), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n15938) );
  AOI22_X1 U19155 ( .A1(n19967), .A2(P1_EBX_REG_12__SCAN_IN), .B1(n15975), 
        .B2(n19961), .ZN(n15936) );
  OAI22_X1 U19156 ( .A1(n20864), .A2(n19905), .B1(n19976), .B2(n16049), .ZN(
        n15934) );
  AOI211_X1 U19157 ( .C1(n15974), .C2(n19942), .A(n10704), .B(n15934), .ZN(
        n15935) );
  OAI211_X1 U19158 ( .C1(n15938), .C2(n15937), .A(n15936), .B(n15935), .ZN(
        P1_U2828) );
  INV_X1 U19159 ( .A(n15939), .ZN(n16059) );
  AOI22_X1 U19160 ( .A1(n16059), .A2(n19948), .B1(n19967), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n15940) );
  OAI21_X1 U19161 ( .B1(n15987), .B2(n19950), .A(n15940), .ZN(n15941) );
  AOI211_X1 U19162 ( .C1(n19962), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n10704), .B(n15941), .ZN(n15944) );
  AOI22_X1 U19163 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n15942), .B1(n19942), 
        .B2(n15984), .ZN(n15943) );
  OAI211_X1 U19164 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n15945), .A(n15944), 
        .B(n15943), .ZN(P1_U2829) );
  AOI22_X1 U19165 ( .A1(n20013), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n10704), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15951) );
  OAI22_X1 U19166 ( .A1(n15948), .A2(n15947), .B1(n20030), .B2(n15946), .ZN(
        n15949) );
  INV_X1 U19167 ( .A(n15949), .ZN(n15950) );
  OAI211_X1 U19168 ( .C1(n20023), .C2(n15952), .A(n15951), .B(n15950), .ZN(
        P1_U2980) );
  NAND2_X1 U19169 ( .A1(n15953), .A2(n15956), .ZN(n15955) );
  MUX2_X1 U19170 ( .A(n15956), .B(n15955), .S(n15954), .Z(n15957) );
  XNOR2_X1 U19171 ( .A(n15957), .B(n16018), .ZN(n16026) );
  AOI22_X1 U19172 ( .A1(n20013), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n10704), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n15961) );
  AOI22_X1 U19173 ( .A1(n15959), .A2(n14447), .B1(n15958), .B2(n15976), .ZN(
        n15960) );
  OAI211_X1 U19174 ( .C1(n20030), .C2(n16026), .A(n15961), .B(n15960), .ZN(
        P1_U2982) );
  NAND2_X1 U19175 ( .A1(n15963), .A2(n15962), .ZN(n15964) );
  XNOR2_X1 U19176 ( .A(n15965), .B(n15964), .ZN(n16033) );
  AOI22_X1 U19177 ( .A1(n20013), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n10704), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15969) );
  AOI22_X1 U19178 ( .A1(n15967), .A2(n14447), .B1(n15966), .B2(n15976), .ZN(
        n15968) );
  OAI211_X1 U19179 ( .C1(n16033), .C2(n20030), .A(n15969), .B(n15968), .ZN(
        P1_U2984) );
  OAI21_X1 U19180 ( .B1(n15972), .B2(n15971), .A(n15970), .ZN(n15973) );
  INV_X1 U19181 ( .A(n15973), .ZN(n16058) );
  AOI22_X1 U19182 ( .A1(n20013), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n10704), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15978) );
  AOI22_X1 U19183 ( .A1(n15976), .A2(n15975), .B1(n14447), .B2(n15974), .ZN(
        n15977) );
  OAI211_X1 U19184 ( .C1(n16058), .C2(n20030), .A(n15978), .B(n15977), .ZN(
        P1_U2987) );
  AOI22_X1 U19185 ( .A1(n20013), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n10704), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15986) );
  NOR2_X1 U19186 ( .A1(n15979), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15982) );
  NOR2_X1 U19187 ( .A1(n13774), .A2(n16074), .ZN(n15981) );
  MUX2_X1 U19188 ( .A(n15982), .B(n15981), .S(n15980), .Z(n15983) );
  INV_X1 U19189 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n20815) );
  XNOR2_X1 U19190 ( .A(n15983), .B(n20815), .ZN(n16061) );
  AOI22_X1 U19191 ( .A1(n20019), .A2(n16061), .B1(n14447), .B2(n15984), .ZN(
        n15985) );
  OAI211_X1 U19192 ( .C1(n20023), .C2(n15987), .A(n15986), .B(n15985), .ZN(
        P1_U2988) );
  AOI22_X1 U19193 ( .A1(n20013), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n10704), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15994) );
  NAND2_X1 U19194 ( .A1(n15989), .A2(n15988), .ZN(n15990) );
  XNOR2_X1 U19195 ( .A(n15991), .B(n15990), .ZN(n16092) );
  AOI22_X1 U19196 ( .A1(n16092), .A2(n20019), .B1(n14447), .B2(n15992), .ZN(
        n15993) );
  OAI211_X1 U19197 ( .C1(n20023), .C2(n19927), .A(n15994), .B(n15993), .ZN(
        P1_U2992) );
  AOI22_X1 U19198 ( .A1(n20013), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n10704), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15999) );
  XNOR2_X1 U19199 ( .A(n15995), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15996) );
  XNOR2_X1 U19200 ( .A(n15997), .B(n15996), .ZN(n16099) );
  AOI22_X1 U19201 ( .A1(n16099), .A2(n20019), .B1(n14447), .B2(n19943), .ZN(
        n15998) );
  OAI211_X1 U19202 ( .C1(n20023), .C2(n19937), .A(n15999), .B(n15998), .ZN(
        P1_U2993) );
  AOI22_X1 U19203 ( .A1(n20013), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n10704), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n16007) );
  OAI21_X1 U19204 ( .B1(n16002), .B2(n16001), .A(n16000), .ZN(n16107) );
  INV_X1 U19205 ( .A(n16107), .ZN(n16005) );
  INV_X1 U19206 ( .A(n16003), .ZN(n16004) );
  AOI22_X1 U19207 ( .A1(n16005), .A2(n20019), .B1(n14447), .B2(n16004), .ZN(
        n16006) );
  OAI211_X1 U19208 ( .C1(n20023), .C2(n16008), .A(n16007), .B(n16006), .ZN(
        P1_U2994) );
  OAI21_X1 U19209 ( .B1(n16009), .B2(n16015), .A(n16037), .ZN(n16022) );
  OAI22_X1 U19210 ( .A1(n16011), .A2(n16106), .B1(n20038), .B2(n16010), .ZN(
        n16012) );
  AOI21_X1 U19211 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n16022), .A(
        n16012), .ZN(n16017) );
  NAND3_X1 U19212 ( .A1(n16015), .A2(n16014), .A3(n16013), .ZN(n16016) );
  OAI211_X1 U19213 ( .C1(n20696), .C2(n20036), .A(n16017), .B(n16016), .ZN(
        P1_U3013) );
  NAND3_X1 U19214 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16019) );
  OAI21_X1 U19215 ( .B1(n16020), .B2(n16019), .A(n16018), .ZN(n16023) );
  AOI22_X1 U19216 ( .A1(n16023), .A2(n16022), .B1(n20059), .B2(n16021), .ZN(
        n16025) );
  NAND2_X1 U19217 ( .A1(n10704), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16024) );
  OAI211_X1 U19218 ( .C1(n16026), .C2(n16106), .A(n16025), .B(n16024), .ZN(
        P1_U3014) );
  NOR2_X1 U19219 ( .A1(n20036), .A2(n20691), .ZN(n16030) );
  AOI21_X1 U19220 ( .B1(n10501), .B2(n16028), .A(n16027), .ZN(n16029) );
  AOI211_X1 U19221 ( .C1(n16031), .C2(n20059), .A(n16030), .B(n16029), .ZN(
        n16032) );
  OAI21_X1 U19222 ( .B1(n16033), .B2(n16106), .A(n16032), .ZN(P1_U3016) );
  INV_X1 U19223 ( .A(n16034), .ZN(n16035) );
  AOI21_X1 U19224 ( .B1(n16036), .B2(n20059), .A(n16035), .ZN(n16041) );
  INV_X1 U19225 ( .A(n16037), .ZN(n16038) );
  AOI22_X1 U19226 ( .A1(n16039), .A2(n20063), .B1(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16038), .ZN(n16040) );
  OAI211_X1 U19227 ( .C1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n16042), .A(
        n16041), .B(n16040), .ZN(P1_U3018) );
  AOI21_X1 U19228 ( .B1(n16043), .B2(n16065), .A(n20034), .ZN(n16045) );
  OAI21_X1 U19229 ( .B1(n16044), .B2(n20056), .A(n20033), .ZN(n16083) );
  AOI211_X1 U19230 ( .C1(n16046), .C2(n16055), .A(n16045), .B(n16083), .ZN(
        n16064) );
  NOR2_X1 U19231 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16047), .ZN(
        n16060) );
  NAND2_X1 U19232 ( .A1(n16060), .A2(n20066), .ZN(n16048) );
  AOI21_X1 U19233 ( .B1(n16064), .B2(n16048), .A(n10499), .ZN(n16051) );
  INV_X1 U19234 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20686) );
  OAI22_X1 U19235 ( .A1(n16049), .A2(n20038), .B1(n20686), .B2(n20036), .ZN(
        n16050) );
  NOR2_X1 U19236 ( .A1(n16051), .A2(n16050), .ZN(n16057) );
  INV_X1 U19237 ( .A(n16052), .ZN(n20032) );
  NAND2_X1 U19238 ( .A1(n20032), .A2(n16053), .ZN(n20047) );
  INV_X1 U19239 ( .A(n16087), .ZN(n16102) );
  OR3_X1 U19240 ( .A1(n16055), .A2(n16102), .A3(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16056) );
  OAI211_X1 U19241 ( .C1(n16058), .C2(n16106), .A(n16057), .B(n16056), .ZN(
        P1_U3019) );
  AOI22_X1 U19242 ( .A1(n16059), .A2(n20059), .B1(n10704), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n16063) );
  AOI22_X1 U19243 ( .A1(n20063), .A2(n16061), .B1(n16087), .B2(n16060), .ZN(
        n16062) );
  OAI211_X1 U19244 ( .C1(n16064), .C2(n20815), .A(n16063), .B(n16062), .ZN(
        P1_U3020) );
  OAI21_X1 U19245 ( .B1(n16065), .B2(n20034), .A(n16068), .ZN(n16067) );
  OAI21_X1 U19246 ( .B1(n16083), .B2(n16067), .A(n16066), .ZN(n16080) );
  NAND2_X1 U19247 ( .A1(n16068), .A2(n16087), .ZN(n16076) );
  AOI221_X1 U19248 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n16074), .C2(n16081), .A(
        n16076), .ZN(n16071) );
  INV_X1 U19249 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20683) );
  OAI22_X1 U19250 ( .A1(n16069), .A2(n20038), .B1(n20683), .B2(n20036), .ZN(
        n16070) );
  AOI211_X1 U19251 ( .C1(n16072), .C2(n20063), .A(n16071), .B(n16070), .ZN(
        n16073) );
  OAI21_X1 U19252 ( .B1(n16074), .B2(n16080), .A(n16073), .ZN(P1_U3021) );
  AOI22_X1 U19253 ( .A1(n19903), .A2(n20059), .B1(n10704), .B2(
        P1_REIP_REG_9__SCAN_IN), .ZN(n16075) );
  OAI21_X1 U19254 ( .B1(n16076), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16075), .ZN(n16077) );
  AOI21_X1 U19255 ( .B1(n16078), .B2(n20063), .A(n16077), .ZN(n16079) );
  OAI21_X1 U19256 ( .B1(n16081), .B2(n16080), .A(n16079), .ZN(P1_U3022) );
  NAND2_X1 U19257 ( .A1(n20039), .A2(n16104), .ZN(n16111) );
  INV_X1 U19258 ( .A(n20034), .ZN(n20035) );
  INV_X1 U19259 ( .A(n20039), .ZN(n16082) );
  OR2_X1 U19260 ( .A1(n16082), .A2(n20054), .ZN(n16084) );
  AOI21_X1 U19261 ( .B1(n20035), .B2(n16084), .A(n16083), .ZN(n16105) );
  OAI21_X1 U19262 ( .B1(n16085), .B2(n16111), .A(n16105), .ZN(n16098) );
  AOI21_X1 U19263 ( .B1(n10606), .B2(n16086), .A(n16098), .ZN(n16094) );
  NAND2_X1 U19264 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16087), .ZN(
        n16096) );
  AOI221_X1 U19265 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n20843), .C2(n16095), .A(
        n16096), .ZN(n16089) );
  INV_X1 U19266 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20679) );
  OAI22_X1 U19267 ( .A1(n19917), .A2(n20038), .B1(n20679), .B2(n20036), .ZN(
        n16088) );
  AOI211_X1 U19268 ( .C1(n16090), .C2(n20063), .A(n16089), .B(n16088), .ZN(
        n16091) );
  OAI21_X1 U19269 ( .B1(n16094), .B2(n20843), .A(n16091), .ZN(P1_U3023) );
  AOI222_X1 U19270 ( .A1(n16092), .A2(n20063), .B1(n20059), .B2(n19932), .C1(
        P1_REIP_REG_7__SCAN_IN), .C2(n10704), .ZN(n16093) );
  OAI221_X1 U19271 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16096), .C1(
        n16095), .C2(n16094), .A(n16093), .ZN(P1_U3024) );
  INV_X1 U19272 ( .A(n19940), .ZN(n16097) );
  AOI22_X1 U19273 ( .A1(n20059), .A2(n16097), .B1(n10704), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n16101) );
  AOI22_X1 U19274 ( .A1(n16099), .A2(n20063), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16098), .ZN(n16100) );
  OAI211_X1 U19275 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16102), .A(
        n16101), .B(n16100), .ZN(P1_U3025) );
  AOI22_X1 U19276 ( .A1(n16103), .A2(n20059), .B1(n10704), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n16110) );
  OAI22_X1 U19277 ( .A1(n16107), .A2(n16106), .B1(n16105), .B2(n16104), .ZN(
        n16108) );
  INV_X1 U19278 ( .A(n16108), .ZN(n16109) );
  OAI211_X1 U19279 ( .C1(n20047), .C2(n16111), .A(n16110), .B(n16109), .ZN(
        P1_U3026) );
  INV_X1 U19280 ( .A(n19949), .ZN(n16114) );
  NAND4_X1 U19281 ( .A1(n16114), .A2(n19877), .A3(n16113), .A4(n16112), .ZN(
        n16115) );
  OAI21_X1 U19282 ( .B1(n16117), .B2(n16116), .A(n16115), .ZN(P1_U3468) );
  INV_X1 U19283 ( .A(n16118), .ZN(n16126) );
  AND2_X1 U19284 ( .A1(n16119), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n16128) );
  NAND4_X1 U19285 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20652), .A4(n20659), .ZN(n16120) );
  NAND2_X1 U19286 ( .A1(n16121), .A2(n16120), .ZN(n20650) );
  NOR2_X1 U19287 ( .A1(n16122), .A2(n20650), .ZN(n16123) );
  OAI22_X1 U19288 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n16128), .B1(n16124), 
        .B2(n16123), .ZN(n16125) );
  AOI211_X1 U19289 ( .C1(n20760), .C2(n20759), .A(n16126), .B(n16125), .ZN(
        P1_U3162) );
  INV_X1 U19290 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20481) );
  OAI21_X1 U19291 ( .B1(n16128), .B2(n20481), .A(n16127), .ZN(P1_U3466) );
  OAI22_X1 U19292 ( .A1(n16129), .A2(n18941), .B1(n19772), .B2(n18923), .ZN(
        n16130) );
  INV_X1 U19293 ( .A(n16130), .ZN(n16140) );
  AOI22_X1 U19294 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18957), .B1(
        P2_EBX_REG_24__SCAN_IN), .B2(n18898), .ZN(n16139) );
  AOI22_X1 U19295 ( .A1(n16132), .A2(n18902), .B1(n18907), .B2(n16131), .ZN(
        n16138) );
  AOI21_X1 U19296 ( .B1(n16135), .B2(n16134), .A(n16133), .ZN(n16136) );
  NAND2_X1 U19297 ( .A1(n18951), .A2(n16136), .ZN(n16137) );
  NAND4_X1 U19298 ( .A1(n16140), .A2(n16139), .A3(n16138), .A4(n16137), .ZN(
        P2_U2831) );
  AOI22_X1 U19299 ( .A1(n18979), .A2(n16141), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n19039), .ZN(n16146) );
  AOI22_X1 U19300 ( .A1(n18981), .A2(BUF1_REG_22__SCAN_IN), .B1(n18980), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n16145) );
  AOI22_X1 U19301 ( .A1(n16143), .A2(n19044), .B1(n19040), .B2(n16142), .ZN(
        n16144) );
  NAND3_X1 U19302 ( .A1(n16146), .A2(n16145), .A3(n16144), .ZN(P2_U2897) );
  AOI22_X1 U19303 ( .A1(n18979), .A2(n16147), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n19039), .ZN(n16151) );
  AOI22_X1 U19304 ( .A1(n18981), .A2(BUF1_REG_20__SCAN_IN), .B1(n18980), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16150) );
  AOI22_X1 U19305 ( .A1(n16148), .A2(n19044), .B1(n19040), .B2(n18795), .ZN(
        n16149) );
  NAND3_X1 U19306 ( .A1(n16151), .A2(n16150), .A3(n16149), .ZN(P2_U2899) );
  AOI22_X1 U19307 ( .A1(n18979), .A2(n16152), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n19039), .ZN(n16156) );
  AOI22_X1 U19308 ( .A1(n18981), .A2(BUF1_REG_18__SCAN_IN), .B1(n18980), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n16155) );
  AOI22_X1 U19309 ( .A1(n16153), .A2(n19044), .B1(n19040), .B2(n18823), .ZN(
        n16154) );
  NAND3_X1 U19310 ( .A1(n16156), .A2(n16155), .A3(n16154), .ZN(P2_U2901) );
  AOI22_X1 U19311 ( .A1(n16184), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19119), .ZN(n16165) );
  NOR3_X1 U19312 ( .A1(n16158), .A2(n16157), .A3(n16194), .ZN(n16163) );
  OAI22_X1 U19313 ( .A1(n16161), .A2(n16192), .B1(n16160), .B2(n16159), .ZN(
        n16162) );
  NOR2_X1 U19314 ( .A1(n16163), .A2(n16162), .ZN(n16164) );
  OAI211_X1 U19315 ( .C1(n16190), .C2(n16166), .A(n16165), .B(n16164), .ZN(
        P2_U2992) );
  AOI22_X1 U19316 ( .A1(n16184), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n19118), .B2(n18844), .ZN(n16174) );
  AOI22_X1 U19317 ( .A1(n16167), .A2(n19124), .B1(n19121), .B2(n18849), .ZN(
        n16173) );
  INV_X1 U19318 ( .A(n16168), .ZN(n16169) );
  OAI211_X1 U19319 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n16170), .A(
        n16169), .B(n19123), .ZN(n16171) );
  NAND4_X1 U19320 ( .A1(n16174), .A2(n16173), .A3(n16172), .A4(n16171), .ZN(
        P2_U2998) );
  AOI22_X1 U19321 ( .A1(n16184), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19119), .ZN(n16183) );
  NAND2_X1 U19322 ( .A1(n16176), .A2(n16175), .ZN(n16177) );
  XNOR2_X1 U19323 ( .A(n16178), .B(n16177), .ZN(n16241) );
  OAI21_X1 U19324 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16180), .A(
        n16179), .ZN(n16244) );
  INV_X1 U19325 ( .A(n16244), .ZN(n16181) );
  AOI222_X1 U19326 ( .A1(n16241), .A2(n19124), .B1(n19121), .B2(n18870), .C1(
        n16181), .C2(n19123), .ZN(n16182) );
  OAI211_X1 U19327 ( .C1(n16190), .C2(n18865), .A(n16183), .B(n16182), .ZN(
        P2_U3000) );
  AOI22_X1 U19328 ( .A1(n16184), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19119), .ZN(n16189) );
  AOI222_X1 U19329 ( .A1(n16187), .A2(n19124), .B1(n19121), .B2(n16186), .C1(
        n19123), .C2(n16185), .ZN(n16188) );
  OAI211_X1 U19330 ( .C1(n16190), .C2(n18888), .A(n16189), .B(n16188), .ZN(
        P2_U3002) );
  AOI22_X1 U19331 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19119), .B1(n19118), 
        .B2(n16191), .ZN(n16198) );
  OAI22_X1 U19332 ( .A1(n16195), .A2(n16194), .B1(n16193), .B2(n16192), .ZN(
        n16196) );
  AOI21_X1 U19333 ( .B1(n19121), .B2(n18903), .A(n16196), .ZN(n16197) );
  OAI211_X1 U19334 ( .C1(n19129), .C2(n16199), .A(n16198), .B(n16197), .ZN(
        P2_U3003) );
  AOI22_X1 U19335 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19119), .B1(n19118), 
        .B2(n18916), .ZN(n16204) );
  AOI222_X1 U19336 ( .A1(n16202), .A2(n19124), .B1(n19121), .B2(n16201), .C1(
        n19123), .C2(n16200), .ZN(n16203) );
  OAI211_X1 U19337 ( .C1(n19129), .C2(n16205), .A(n16204), .B(n16203), .ZN(
        P2_U3004) );
  AOI22_X1 U19338 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19119), .B1(n19118), 
        .B2(n16206), .ZN(n16211) );
  AOI222_X1 U19339 ( .A1(n16209), .A2(n19123), .B1(n16208), .B2(n19124), .C1(
        n19121), .C2(n16207), .ZN(n16210) );
  OAI211_X1 U19340 ( .C1(n19129), .C2(n16212), .A(n16211), .B(n16210), .ZN(
        P2_U3006) );
  AOI22_X1 U19341 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n19119), .B1(n19118), 
        .B2(n16213), .ZN(n16219) );
  INV_X1 U19342 ( .A(n16214), .ZN(n16217) );
  AOI222_X1 U19343 ( .A1(n19123), .A2(n16217), .B1(n16216), .B2(n19124), .C1(
        n19121), .C2(n16215), .ZN(n16218) );
  OAI211_X1 U19344 ( .C1(n19129), .C2(n20876), .A(n16219), .B(n16218), .ZN(
        P2_U3008) );
  INV_X1 U19345 ( .A(n16237), .ZN(n16220) );
  XNOR2_X1 U19346 ( .A(n16221), .B(n16220), .ZN(n18990) );
  NAND2_X1 U19347 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19119), .ZN(n16222) );
  OAI221_X1 U19348 ( .B1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16225), 
        .C1(n16224), .C2(n16223), .A(n16222), .ZN(n16226) );
  AOI21_X1 U19349 ( .B1(n19155), .B2(n18990), .A(n16226), .ZN(n16230) );
  AOI22_X1 U19350 ( .A1(n18859), .A2(n19156), .B1(n16228), .B2(n16227), .ZN(
        n16229) );
  OAI211_X1 U19351 ( .C1(n16231), .C2(n19166), .A(n16230), .B(n16229), .ZN(
        P2_U3031) );
  NOR2_X1 U19352 ( .A1(n16233), .A2(n16232), .ZN(n16236) );
  INV_X1 U19353 ( .A(n16234), .ZN(n16235) );
  MUX2_X1 U19354 ( .A(n16236), .B(n16235), .S(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n16240) );
  AOI21_X1 U19355 ( .B1(n16238), .B2(n15476), .A(n16237), .ZN(n18869) );
  INV_X1 U19356 ( .A(n18869), .ZN(n18995) );
  INV_X1 U19357 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19756) );
  OAI22_X1 U19358 ( .A1(n19136), .A2(n18995), .B1(n19756), .B2(n18921), .ZN(
        n16239) );
  NOR2_X1 U19359 ( .A1(n16240), .A2(n16239), .ZN(n16243) );
  AOI22_X1 U19360 ( .A1(n16241), .A2(n19131), .B1(n19156), .B2(n18870), .ZN(
        n16242) );
  OAI211_X1 U19361 ( .C1(n19159), .C2(n16244), .A(n16243), .B(n16242), .ZN(
        P2_U3032) );
  INV_X1 U19362 ( .A(n16245), .ZN(n16246) );
  OAI22_X1 U19363 ( .A1(n19166), .A2(n16247), .B1(n19136), .B2(n16246), .ZN(
        n16252) );
  OAI22_X1 U19364 ( .A1(n16250), .A2(n19151), .B1(n16249), .B2(n16248), .ZN(
        n16251) );
  AOI211_X1 U19365 ( .C1(n19151), .C2(n19153), .A(n16252), .B(n16251), .ZN(
        n16254) );
  OAI211_X1 U19366 ( .C1(n19159), .C2(n16255), .A(n16254), .B(n16253), .ZN(
        P2_U3046) );
  MUX2_X1 U19367 ( .A(n11637), .B(n16256), .S(n16285), .Z(n16288) );
  NOR2_X1 U19368 ( .A1(n16285), .A2(n16257), .ZN(n16258) );
  AOI21_X1 U19369 ( .B1(n16259), .B2(n16285), .A(n16258), .ZN(n16284) );
  OAI21_X1 U19370 ( .B1(n16284), .B2(n19819), .A(n19811), .ZN(n16260) );
  OAI21_X1 U19371 ( .B1(n16288), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n16260), .ZN(n16267) );
  INV_X1 U19372 ( .A(n16285), .ZN(n16264) );
  INV_X1 U19373 ( .A(n16265), .ZN(n16262) );
  AOI211_X1 U19374 ( .C1(n16262), .C2(n19828), .A(n19839), .B(n16261), .ZN(
        n16263) );
  AOI211_X1 U19375 ( .C1(n16265), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n16264), .B(n16263), .ZN(n16266) );
  AOI22_X1 U19376 ( .A1(n16267), .A2(n16266), .B1(n16284), .B2(n19278), .ZN(
        n16268) );
  OAI21_X1 U19377 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16288), .A(
        n16268), .ZN(n16291) );
  INV_X1 U19378 ( .A(n16269), .ZN(n16275) );
  OAI22_X1 U19379 ( .A1(n16275), .A2(n16272), .B1(n16270), .B2(n16271), .ZN(
        n16273) );
  AOI21_X1 U19380 ( .B1(n16275), .B2(n16274), .A(n16273), .ZN(n19847) );
  INV_X1 U19381 ( .A(n16276), .ZN(n16278) );
  AOI21_X1 U19382 ( .B1(n16278), .B2(n19860), .A(n16277), .ZN(n16283) );
  NOR4_X1 U19383 ( .A1(n16270), .A2(n16281), .A3(n16280), .A4(n16279), .ZN(
        n18775) );
  OAI21_X1 U19384 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n18775), .ZN(n16282) );
  NAND3_X1 U19385 ( .A1(n19847), .A2(n16283), .A3(n16282), .ZN(n16290) );
  INV_X1 U19386 ( .A(n16284), .ZN(n16287) );
  OAI22_X1 U19387 ( .A1(n16288), .A2(n16287), .B1(n16286), .B2(n16285), .ZN(
        n16289) );
  AOI211_X1 U19388 ( .C1(n16292), .C2(n16291), .A(n16290), .B(n16289), .ZN(
        n16303) );
  NOR2_X1 U19389 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n11587), .ZN(n19711) );
  AOI21_X1 U19390 ( .B1(n19717), .B2(n19711), .A(n16293), .ZN(n16302) );
  AOI211_X1 U19391 ( .C1(n16295), .C2(n16294), .A(n19853), .B(n19852), .ZN(
        n16298) );
  OAI221_X1 U19392 ( .B1(n12437), .B2(n11587), .C1(n16303), .C2(n11587), .A(
        n16298), .ZN(n16296) );
  INV_X1 U19393 ( .A(n16296), .ZN(n19715) );
  NOR2_X1 U19394 ( .A1(n19715), .A2(n11587), .ZN(n16306) );
  OAI21_X1 U19395 ( .B1(n16297), .B2(n16306), .A(n19863), .ZN(n16300) );
  NAND3_X1 U19396 ( .A1(n19717), .A2(n16298), .A3(n11587), .ZN(n16299) );
  AOI22_X1 U19397 ( .A1(n19848), .A2(n16304), .B1(n16300), .B2(n16299), .ZN(
        n16301) );
  OAI211_X1 U19398 ( .C1(n16303), .C2(n19049), .A(n16302), .B(n16301), .ZN(
        P2_U3176) );
  INV_X1 U19399 ( .A(n16304), .ZN(n16305) );
  OAI21_X1 U19400 ( .B1(n16306), .B2(n19416), .A(n16305), .ZN(P2_U3593) );
  XOR2_X1 U19401 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n16327), .Z(
        n16494) );
  INV_X1 U19402 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16499) );
  OAI221_X1 U19403 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16309), .C1(
        n16499), .C2(n16308), .A(n16307), .ZN(n16310) );
  AOI21_X1 U19404 ( .B1(n17532), .B2(n16494), .A(n16310), .ZN(n16315) );
  NAND2_X1 U19405 ( .A1(n17603), .A2(n16311), .ZN(n16323) );
  OAI21_X1 U19406 ( .B1(n16319), .B2(n17768), .A(n16323), .ZN(n16313) );
  NAND2_X1 U19407 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17497), .ZN(
        n17481) );
  AOI22_X1 U19408 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16313), .B1(
        n16312), .B2(n17436), .ZN(n16314) );
  OAI211_X1 U19409 ( .C1(n17678), .C2(n16316), .A(n16315), .B(n16314), .ZN(
        P3_U2800) );
  NAND2_X1 U19410 ( .A1(n16318), .A2(n16317), .ZN(n16348) );
  AOI211_X1 U19411 ( .C1(n16320), .C2(n16348), .A(n16319), .B(n17768), .ZN(
        n16326) );
  NOR2_X1 U19412 ( .A1(n16321), .A2(n17424), .ZN(n16350) );
  NOR2_X1 U19413 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16350), .ZN(
        n16324) );
  OAI22_X1 U19414 ( .A1(n16324), .A2(n16323), .B1(n17678), .B2(n16322), .ZN(
        n16325) );
  NOR2_X1 U19415 ( .A1(n16326), .A2(n16325), .ZN(n16334) );
  INV_X1 U19416 ( .A(n18069), .ZN(n17985) );
  NAND2_X1 U19417 ( .A1(n17985), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16333) );
  INV_X1 U19418 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16511) );
  AOI21_X1 U19419 ( .B1(n16511), .B2(n16477), .A(n16327), .ZN(n16505) );
  OAI21_X1 U19420 ( .B1(n16328), .B2(n17532), .A(n16505), .ZN(n16332) );
  OAI221_X1 U19421 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18478), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n16330), .A(n16329), .ZN(
        n16331) );
  NAND4_X1 U19422 ( .A1(n16334), .A2(n16333), .A3(n16332), .A4(n16331), .ZN(
        P3_U2801) );
  NAND2_X1 U19423 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n10849), .ZN(
        n17428) );
  INV_X1 U19424 ( .A(n17775), .ZN(n16337) );
  INV_X1 U19425 ( .A(n17954), .ZN(n17643) );
  AOI22_X1 U19426 ( .A1(n18530), .A2(n17643), .B1(n17644), .B2(n17953), .ZN(
        n17938) );
  INV_X1 U19427 ( .A(n17904), .ZN(n16335) );
  INV_X1 U19428 ( .A(n17991), .ZN(n18052) );
  AOI22_X1 U19429 ( .A1(n18566), .A2(n16335), .B1(n18052), .B2(n17921), .ZN(
        n17937) );
  AOI21_X1 U19430 ( .B1(n17938), .B2(n17937), .A(n17552), .ZN(n17839) );
  NAND2_X1 U19431 ( .A1(n16336), .A2(n17839), .ZN(n17819) );
  NOR2_X1 U19432 ( .A1(n18086), .A2(n17819), .ZN(n17807) );
  NAND2_X1 U19433 ( .A1(n16337), .A2(n17807), .ZN(n17769) );
  OAI21_X1 U19434 ( .B1(n10849), .B2(n17564), .A(n16343), .ZN(n16338) );
  INV_X1 U19435 ( .A(n16338), .ZN(n17415) );
  NAND3_X1 U19436 ( .A1(n16340), .A2(n17415), .A3(n16339), .ZN(n16341) );
  OAI21_X1 U19437 ( .B1(n16343), .B2(n16342), .A(n16341), .ZN(n16344) );
  AOI22_X1 U19438 ( .A1(n9612), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n18085), 
        .B2(n16344), .ZN(n16354) );
  NOR2_X1 U19439 ( .A1(n17416), .A2(n17415), .ZN(n17414) );
  NOR4_X1 U19440 ( .A1(n16345), .A2(n17278), .A3(n17414), .A4(n18534), .ZN(
        n16352) );
  AOI211_X1 U19441 ( .C1(n18530), .C2(n16348), .A(n16347), .B(n16346), .ZN(
        n16349) );
  OAI21_X1 U19442 ( .B1(n16350), .B2(n17995), .A(n16349), .ZN(n16351) );
  OAI211_X1 U19443 ( .C1(n16352), .C2(n16351), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18069), .ZN(n16353) );
  OAI211_X1 U19444 ( .C1(n17428), .C2(n17769), .A(n16354), .B(n16353), .ZN(
        P3_U2834) );
  NOR3_X1 U19445 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16356) );
  NOR4_X1 U19446 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16355) );
  NAND4_X1 U19447 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16356), .A3(n16355), .A4(
        U215), .ZN(U213) );
  INV_X1 U19448 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16449) );
  INV_X2 U19449 ( .A(U214), .ZN(n16411) );
  INV_X1 U19450 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16450) );
  OAI222_X1 U19451 ( .A1(U212), .A2(n16449), .B1(n16413), .B2(n16358), .C1(
        U214), .C2(n16450), .ZN(U216) );
  INV_X1 U19452 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16360) );
  AOI22_X1 U19453 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16399), .ZN(n16359) );
  OAI21_X1 U19454 ( .B1(n16360), .B2(n16413), .A(n16359), .ZN(U217) );
  INV_X1 U19455 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16362) );
  AOI22_X1 U19456 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16399), .ZN(n16361) );
  OAI21_X1 U19457 ( .B1(n16362), .B2(n16413), .A(n16361), .ZN(U218) );
  INV_X1 U19458 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16364) );
  AOI22_X1 U19459 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16399), .ZN(n16363) );
  OAI21_X1 U19460 ( .B1(n16364), .B2(n16413), .A(n16363), .ZN(U219) );
  AOI22_X1 U19461 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16399), .ZN(n16365) );
  OAI21_X1 U19462 ( .B1(n14282), .B2(n16413), .A(n16365), .ZN(U220) );
  INV_X1 U19463 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16367) );
  AOI22_X1 U19464 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16399), .ZN(n16366) );
  OAI21_X1 U19465 ( .B1(n16367), .B2(n16413), .A(n16366), .ZN(U221) );
  INV_X1 U19466 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16369) );
  AOI22_X1 U19467 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16399), .ZN(n16368) );
  OAI21_X1 U19468 ( .B1(n16369), .B2(n16413), .A(n16368), .ZN(U222) );
  INV_X1 U19469 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16371) );
  AOI22_X1 U19470 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16399), .ZN(n16370) );
  OAI21_X1 U19471 ( .B1(n16371), .B2(n16413), .A(n16370), .ZN(U223) );
  AOI22_X1 U19472 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16399), .ZN(n16372) );
  OAI21_X1 U19473 ( .B1(n15108), .B2(n16413), .A(n16372), .ZN(U224) );
  INV_X1 U19474 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16374) );
  AOI22_X1 U19475 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16399), .ZN(n16373) );
  OAI21_X1 U19476 ( .B1(n16374), .B2(n16413), .A(n16373), .ZN(U225) );
  AOI22_X1 U19477 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16399), .ZN(n16375) );
  OAI21_X1 U19478 ( .B1(n16376), .B2(n16413), .A(n16375), .ZN(U226) );
  INV_X1 U19479 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16378) );
  AOI22_X1 U19480 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16399), .ZN(n16377) );
  OAI21_X1 U19481 ( .B1(n16378), .B2(n16413), .A(n16377), .ZN(U227) );
  AOI22_X1 U19482 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16399), .ZN(n16379) );
  OAI21_X1 U19483 ( .B1(n16380), .B2(n16413), .A(n16379), .ZN(U228) );
  INV_X1 U19484 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16382) );
  AOI22_X1 U19485 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16399), .ZN(n16381) );
  OAI21_X1 U19486 ( .B1(n16382), .B2(n16413), .A(n16381), .ZN(U229) );
  AOI22_X1 U19487 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16399), .ZN(n16383) );
  OAI21_X1 U19488 ( .B1(n15130), .B2(n16413), .A(n16383), .ZN(U230) );
  INV_X1 U19489 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16385) );
  AOI22_X1 U19490 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16399), .ZN(n16384) );
  OAI21_X1 U19491 ( .B1(n16385), .B2(n16413), .A(n16384), .ZN(U231) );
  AOI22_X1 U19492 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16399), .ZN(n16386) );
  OAI21_X1 U19493 ( .B1(n12894), .B2(n16413), .A(n16386), .ZN(U232) );
  AOI22_X1 U19494 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16399), .ZN(n16387) );
  OAI21_X1 U19495 ( .B1(n12671), .B2(n16413), .A(n16387), .ZN(U233) );
  INV_X1 U19496 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16389) );
  AOI22_X1 U19497 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16399), .ZN(n16388) );
  OAI21_X1 U19498 ( .B1(n16389), .B2(n16413), .A(n16388), .ZN(U234) );
  AOI22_X1 U19499 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16399), .ZN(n16390) );
  OAI21_X1 U19500 ( .B1(n12474), .B2(n16413), .A(n16390), .ZN(U235) );
  AOI22_X1 U19501 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16399), .ZN(n16391) );
  OAI21_X1 U19502 ( .B1(n12468), .B2(n16413), .A(n16391), .ZN(U236) );
  AOI22_X1 U19503 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16399), .ZN(n16392) );
  OAI21_X1 U19504 ( .B1(n16393), .B2(n16413), .A(n16392), .ZN(U237) );
  AOI22_X1 U19505 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16399), .ZN(n16394) );
  OAI21_X1 U19506 ( .B1(n12488), .B2(n16413), .A(n16394), .ZN(U238) );
  INV_X1 U19507 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16396) );
  AOI22_X1 U19508 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16399), .ZN(n16395) );
  OAI21_X1 U19509 ( .B1(n16396), .B2(n16413), .A(n16395), .ZN(U239) );
  INV_X1 U19510 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16398) );
  AOI22_X1 U19511 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16399), .ZN(n16397) );
  OAI21_X1 U19512 ( .B1(n16398), .B2(n16413), .A(n16397), .ZN(U240) );
  AOI22_X1 U19513 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16399), .ZN(n16400) );
  OAI21_X1 U19514 ( .B1(n16401), .B2(n16413), .A(n16400), .ZN(U241) );
  INV_X1 U19515 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16403) );
  AOI22_X1 U19516 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16399), .ZN(n16402) );
  OAI21_X1 U19517 ( .B1(n16403), .B2(n16413), .A(n16402), .ZN(U242) );
  INV_X1 U19518 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16405) );
  AOI22_X1 U19519 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16399), .ZN(n16404) );
  OAI21_X1 U19520 ( .B1(n16405), .B2(n16413), .A(n16404), .ZN(U243) );
  INV_X1 U19521 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16407) );
  AOI22_X1 U19522 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16399), .ZN(n16406) );
  OAI21_X1 U19523 ( .B1(n16407), .B2(n16413), .A(n16406), .ZN(U244) );
  AOI22_X1 U19524 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16399), .ZN(n16408) );
  OAI21_X1 U19525 ( .B1(n20859), .B2(n16413), .A(n16408), .ZN(U245) );
  INV_X1 U19526 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16410) );
  AOI22_X1 U19527 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16399), .ZN(n16409) );
  OAI21_X1 U19528 ( .B1(n16410), .B2(n16413), .A(n16409), .ZN(U246) );
  AOI22_X1 U19529 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16411), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16399), .ZN(n16412) );
  OAI21_X1 U19530 ( .B1(n16414), .B2(n16413), .A(n16412), .ZN(U247) );
  INV_X1 U19531 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16415) );
  AOI22_X1 U19532 ( .A1(n16445), .A2(n16415), .B1(n18098), .B2(U215), .ZN(U251) );
  OAI22_X1 U19533 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16445), .ZN(n16416) );
  INV_X1 U19534 ( .A(n16416), .ZN(U252) );
  INV_X1 U19535 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16417) );
  AOI22_X1 U19536 ( .A1(n16445), .A2(n16417), .B1(n18108), .B2(U215), .ZN(U253) );
  INV_X1 U19537 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16418) );
  INV_X1 U19538 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18113) );
  AOI22_X1 U19539 ( .A1(n16445), .A2(n16418), .B1(n18113), .B2(U215), .ZN(U254) );
  INV_X1 U19540 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16419) );
  INV_X1 U19541 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18118) );
  AOI22_X1 U19542 ( .A1(n16445), .A2(n16419), .B1(n18118), .B2(U215), .ZN(U255) );
  INV_X1 U19543 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16420) );
  INV_X1 U19544 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18123) );
  AOI22_X1 U19545 ( .A1(n16447), .A2(n16420), .B1(n18123), .B2(U215), .ZN(U256) );
  INV_X1 U19546 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16421) );
  INV_X1 U19547 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n20932) );
  AOI22_X1 U19548 ( .A1(n16445), .A2(n16421), .B1(n20932), .B2(U215), .ZN(U257) );
  INV_X1 U19549 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16422) );
  INV_X1 U19550 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18131) );
  AOI22_X1 U19551 ( .A1(n16445), .A2(n16422), .B1(n18131), .B2(U215), .ZN(U258) );
  INV_X1 U19552 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16423) );
  INV_X1 U19553 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17276) );
  AOI22_X1 U19554 ( .A1(n16447), .A2(n16423), .B1(n17276), .B2(U215), .ZN(U259) );
  INV_X1 U19555 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16424) );
  INV_X1 U19556 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17269) );
  AOI22_X1 U19557 ( .A1(n16445), .A2(n16424), .B1(n17269), .B2(U215), .ZN(U260) );
  INV_X1 U19558 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16425) );
  INV_X1 U19559 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17265) );
  AOI22_X1 U19560 ( .A1(n16447), .A2(n16425), .B1(n17265), .B2(U215), .ZN(U261) );
  OAI22_X1 U19561 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16445), .ZN(n16426) );
  INV_X1 U19562 ( .A(n16426), .ZN(U262) );
  INV_X1 U19563 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16427) );
  INV_X1 U19564 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17257) );
  AOI22_X1 U19565 ( .A1(n16445), .A2(n16427), .B1(n17257), .B2(U215), .ZN(U263) );
  INV_X1 U19566 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16428) );
  INV_X1 U19567 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17252) );
  AOI22_X1 U19568 ( .A1(n16445), .A2(n16428), .B1(n17252), .B2(U215), .ZN(U264) );
  OAI22_X1 U19569 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16447), .ZN(n16429) );
  INV_X1 U19570 ( .A(n16429), .ZN(U265) );
  OAI22_X1 U19571 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16447), .ZN(n16430) );
  INV_X1 U19572 ( .A(n16430), .ZN(U266) );
  OAI22_X1 U19573 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16447), .ZN(n16431) );
  INV_X1 U19574 ( .A(n16431), .ZN(U267) );
  INV_X1 U19575 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n16432) );
  AOI22_X1 U19576 ( .A1(n16445), .A2(n16432), .B1(n15128), .B2(U215), .ZN(U268) );
  OAI22_X1 U19577 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16447), .ZN(n16433) );
  INV_X1 U19578 ( .A(n16433), .ZN(U269) );
  OAI22_X1 U19579 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16447), .ZN(n16434) );
  INV_X1 U19580 ( .A(n16434), .ZN(U270) );
  OAI22_X1 U19581 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16447), .ZN(n16435) );
  INV_X1 U19582 ( .A(n16435), .ZN(U271) );
  INV_X1 U19583 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n16436) );
  AOI22_X1 U19584 ( .A1(n16445), .A2(n16436), .B1(n15113), .B2(U215), .ZN(U272) );
  OAI22_X1 U19585 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16445), .ZN(n16437) );
  INV_X1 U19586 ( .A(n16437), .ZN(U273) );
  OAI22_X1 U19587 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16445), .ZN(n16438) );
  INV_X1 U19588 ( .A(n16438), .ZN(U274) );
  OAI22_X1 U19589 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16445), .ZN(n16439) );
  INV_X1 U19590 ( .A(n16439), .ZN(U275) );
  OAI22_X1 U19591 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16445), .ZN(n16440) );
  INV_X1 U19592 ( .A(n16440), .ZN(U276) );
  OAI22_X1 U19593 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16445), .ZN(n16441) );
  INV_X1 U19594 ( .A(n16441), .ZN(U277) );
  OAI22_X1 U19595 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16445), .ZN(n16442) );
  INV_X1 U19596 ( .A(n16442), .ZN(U278) );
  OAI22_X1 U19597 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16445), .ZN(n16443) );
  INV_X1 U19598 ( .A(n16443), .ZN(U279) );
  OAI22_X1 U19599 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16445), .ZN(n16444) );
  INV_X1 U19600 ( .A(n16444), .ZN(U280) );
  OAI22_X1 U19601 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16445), .ZN(n16446) );
  INV_X1 U19602 ( .A(n16446), .ZN(U281) );
  INV_X1 U19603 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18133) );
  AOI22_X1 U19604 ( .A1(n16447), .A2(n16449), .B1(n18133), .B2(U215), .ZN(U282) );
  INV_X1 U19605 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16448) );
  AOI222_X1 U19606 ( .A1(n16450), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16449), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16448), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16451) );
  INV_X1 U19607 ( .A(n16453), .ZN(n16452) );
  INV_X1 U19608 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18651) );
  INV_X1 U19609 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19750) );
  AOI22_X1 U19610 ( .A1(n16452), .A2(n18651), .B1(n19750), .B2(n16453), .ZN(
        U347) );
  INV_X1 U19611 ( .A(n16453), .ZN(n16454) );
  INV_X1 U19612 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18649) );
  INV_X1 U19613 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19748) );
  AOI22_X1 U19614 ( .A1(n16454), .A2(n18649), .B1(n19748), .B2(n16453), .ZN(
        U348) );
  INV_X1 U19615 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18646) );
  INV_X1 U19616 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19746) );
  AOI22_X1 U19617 ( .A1(n16452), .A2(n18646), .B1(n19746), .B2(n16453), .ZN(
        U349) );
  INV_X1 U19618 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18645) );
  INV_X1 U19619 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19744) );
  AOI22_X1 U19620 ( .A1(n16452), .A2(n18645), .B1(n19744), .B2(n16453), .ZN(
        U350) );
  INV_X1 U19621 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18643) );
  INV_X1 U19622 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19742) );
  AOI22_X1 U19623 ( .A1(n16452), .A2(n18643), .B1(n19742), .B2(n16453), .ZN(
        U351) );
  INV_X1 U19624 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18640) );
  INV_X1 U19625 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19740) );
  AOI22_X1 U19626 ( .A1(n16452), .A2(n18640), .B1(n19740), .B2(n16453), .ZN(
        U352) );
  INV_X1 U19627 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18639) );
  INV_X1 U19628 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19739) );
  AOI22_X1 U19629 ( .A1(n16454), .A2(n18639), .B1(n19739), .B2(n16453), .ZN(
        U353) );
  INV_X1 U19630 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18637) );
  AOI22_X1 U19631 ( .A1(n16452), .A2(n18637), .B1(n19738), .B2(n16453), .ZN(
        U354) );
  INV_X1 U19632 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18689) );
  INV_X1 U19633 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19785) );
  AOI22_X1 U19634 ( .A1(n16452), .A2(n18689), .B1(n19785), .B2(n16453), .ZN(
        U355) );
  INV_X1 U19635 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18686) );
  INV_X1 U19636 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19783) );
  AOI22_X1 U19637 ( .A1(n16452), .A2(n18686), .B1(n19783), .B2(n16453), .ZN(
        U356) );
  INV_X1 U19638 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18683) );
  INV_X1 U19639 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19781) );
  AOI22_X1 U19640 ( .A1(n16452), .A2(n18683), .B1(n19781), .B2(n16453), .ZN(
        U357) );
  INV_X1 U19641 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18682) );
  INV_X1 U19642 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19777) );
  AOI22_X1 U19643 ( .A1(n16452), .A2(n18682), .B1(n19777), .B2(n16453), .ZN(
        U358) );
  INV_X1 U19644 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18681) );
  INV_X1 U19645 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19776) );
  AOI22_X1 U19646 ( .A1(n16452), .A2(n18681), .B1(n19776), .B2(n16453), .ZN(
        U359) );
  INV_X1 U19647 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18680) );
  INV_X1 U19648 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19775) );
  AOI22_X1 U19649 ( .A1(n16452), .A2(n18680), .B1(n19775), .B2(n16453), .ZN(
        U360) );
  INV_X1 U19650 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18678) );
  INV_X1 U19651 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19773) );
  AOI22_X1 U19652 ( .A1(n16452), .A2(n18678), .B1(n19773), .B2(n16453), .ZN(
        U361) );
  INV_X1 U19653 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18676) );
  INV_X1 U19654 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19771) );
  AOI22_X1 U19655 ( .A1(n16452), .A2(n18676), .B1(n19771), .B2(n16453), .ZN(
        U362) );
  INV_X1 U19656 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18675) );
  INV_X1 U19657 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19770) );
  AOI22_X1 U19658 ( .A1(n16452), .A2(n18675), .B1(n19770), .B2(n16453), .ZN(
        U363) );
  INV_X1 U19659 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18672) );
  INV_X1 U19660 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19768) );
  AOI22_X1 U19661 ( .A1(n16452), .A2(n18672), .B1(n19768), .B2(n16453), .ZN(
        U364) );
  INV_X1 U19662 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18635) );
  INV_X1 U19663 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19737) );
  AOI22_X1 U19664 ( .A1(n16452), .A2(n18635), .B1(n19737), .B2(n16453), .ZN(
        U365) );
  INV_X1 U19665 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18670) );
  INV_X1 U19666 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20892) );
  AOI22_X1 U19667 ( .A1(n16452), .A2(n18670), .B1(n20892), .B2(n16453), .ZN(
        U366) );
  INV_X1 U19668 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18669) );
  INV_X1 U19669 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19765) );
  AOI22_X1 U19670 ( .A1(n16452), .A2(n18669), .B1(n19765), .B2(n16453), .ZN(
        U367) );
  INV_X1 U19671 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18667) );
  INV_X1 U19672 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19763) );
  AOI22_X1 U19673 ( .A1(n16452), .A2(n18667), .B1(n19763), .B2(n16453), .ZN(
        U368) );
  INV_X1 U19674 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18665) );
  INV_X1 U19675 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19761) );
  AOI22_X1 U19676 ( .A1(n16452), .A2(n18665), .B1(n19761), .B2(n16453), .ZN(
        U369) );
  INV_X1 U19677 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18663) );
  INV_X1 U19678 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19759) );
  AOI22_X1 U19679 ( .A1(n16452), .A2(n18663), .B1(n19759), .B2(n16453), .ZN(
        U370) );
  INV_X1 U19680 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18661) );
  INV_X1 U19681 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19758) );
  AOI22_X1 U19682 ( .A1(n16454), .A2(n18661), .B1(n19758), .B2(n16453), .ZN(
        U371) );
  INV_X1 U19683 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18659) );
  INV_X1 U19684 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19757) );
  AOI22_X1 U19685 ( .A1(n16454), .A2(n18659), .B1(n19757), .B2(n16453), .ZN(
        U372) );
  INV_X1 U19686 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18657) );
  INV_X1 U19687 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19755) );
  AOI22_X1 U19688 ( .A1(n16454), .A2(n18657), .B1(n19755), .B2(n16453), .ZN(
        U373) );
  INV_X1 U19689 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18654) );
  INV_X1 U19690 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19753) );
  AOI22_X1 U19691 ( .A1(n16454), .A2(n18654), .B1(n19753), .B2(n16453), .ZN(
        U374) );
  INV_X1 U19692 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18653) );
  INV_X1 U19693 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19751) );
  AOI22_X1 U19694 ( .A1(n16454), .A2(n18653), .B1(n19751), .B2(n16453), .ZN(
        U375) );
  INV_X1 U19695 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18632) );
  INV_X1 U19696 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19735) );
  AOI22_X1 U19697 ( .A1(n16454), .A2(n18632), .B1(n19735), .B2(n16453), .ZN(
        U376) );
  INV_X1 U19698 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16455) );
  NOR2_X1 U19699 ( .A1(n18618), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18620) );
  OAI22_X1 U19700 ( .A1(n18629), .A2(n18620), .B1(n18618), .B2(
        P3_STATE_REG_0__SCAN_IN), .ZN(n18614) );
  INV_X1 U19701 ( .A(n18614), .ZN(n18702) );
  INV_X1 U19702 ( .A(n18702), .ZN(n18615) );
  OAI21_X1 U19703 ( .B1(n18629), .B2(n16455), .A(n18615), .ZN(P3_U2633) );
  NOR3_X1 U19704 ( .A1(n16462), .A2(n16461), .A3(n18600), .ZN(n17304) );
  INV_X1 U19705 ( .A(P3_CODEFETCH_REG_SCAN_IN), .ZN(n16457) );
  OAI22_X1 U19706 ( .A1(n17304), .A2(n16457), .B1(n18605), .B2(n16456), .ZN(
        P3_U2634) );
  INV_X1 U19707 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18631) );
  AOI21_X1 U19708 ( .B1(n18629), .B2(n18631), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16458) );
  AOI22_X1 U19709 ( .A1(n18761), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16458), 
        .B2(n18759), .ZN(P3_U2635) );
  NOR2_X1 U19710 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18616) );
  OAI21_X1 U19711 ( .B1(n18616), .B2(BS16), .A(n18702), .ZN(n18700) );
  OAI21_X1 U19712 ( .B1(n18702), .B2(n18749), .A(n18700), .ZN(P3_U2636) );
  INV_X1 U19713 ( .A(n16459), .ZN(n16460) );
  NOR3_X1 U19714 ( .A1(n16462), .A2(n16461), .A3(n16460), .ZN(n18537) );
  NOR2_X1 U19715 ( .A1(n18537), .A2(n18600), .ZN(n18741) );
  OAI21_X1 U19716 ( .B1(n18741), .B2(n18091), .A(n16463), .ZN(P3_U2637) );
  NOR4_X1 U19717 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n16467) );
  NOR4_X1 U19718 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16466) );
  NOR4_X1 U19719 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16465) );
  NOR4_X1 U19720 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n16464) );
  NAND4_X1 U19721 ( .A1(n16467), .A2(n16466), .A3(n16465), .A4(n16464), .ZN(
        n16473) );
  NOR4_X1 U19722 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n16471) );
  AOI211_X1 U19723 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_28__SCAN_IN), .B(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16470) );
  NOR4_X1 U19724 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16469) );
  NOR4_X1 U19725 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16468) );
  NAND4_X1 U19726 ( .A1(n16471), .A2(n16470), .A3(n16469), .A4(n16468), .ZN(
        n16472) );
  NOR2_X1 U19727 ( .A1(n16473), .A2(n16472), .ZN(n18739) );
  INV_X1 U19728 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18696) );
  NOR3_X1 U19729 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16475) );
  OAI21_X1 U19730 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16475), .A(n18739), .ZN(
        n16474) );
  OAI21_X1 U19731 ( .B1(n18739), .B2(n18696), .A(n16474), .ZN(P3_U2638) );
  INV_X1 U19732 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18693) );
  NOR2_X1 U19733 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18733) );
  OAI21_X1 U19734 ( .B1(n16475), .B2(n18733), .A(n18739), .ZN(n16476) );
  OAI21_X1 U19735 ( .B1(n18739), .B2(n18693), .A(n16476), .ZN(P3_U2639) );
  NAND2_X1 U19736 ( .A1(n16529), .A2(n16889), .ZN(n16528) );
  NOR2_X1 U19737 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16528), .ZN(n16512) );
  INV_X1 U19738 ( .A(n16512), .ZN(n16502) );
  NOR2_X1 U19739 ( .A1(n16838), .A2(n16492), .ZN(n16495) );
  INV_X1 U19740 ( .A(n16495), .ZN(n16491) );
  INV_X1 U19741 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n20847) );
  NOR2_X1 U19742 ( .A1(n16480), .A2(n20847), .ZN(n16478) );
  OAI21_X1 U19743 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16478), .A(
        n16477), .ZN(n17421) );
  INV_X1 U19744 ( .A(n17421), .ZN(n16515) );
  OAI22_X1 U19745 ( .A1(n16480), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B1(
        n20847), .B2(n16479), .ZN(n17430) );
  NOR2_X1 U19746 ( .A1(n16481), .A2(n9794), .ZN(n16524) );
  NOR2_X1 U19747 ( .A1(n17430), .A2(n16524), .ZN(n16523) );
  NOR2_X1 U19748 ( .A1(n16523), .A2(n9794), .ZN(n16514) );
  NOR2_X1 U19749 ( .A1(n16515), .A2(n16514), .ZN(n16513) );
  NOR2_X1 U19750 ( .A1(n16513), .A2(n9794), .ZN(n16504) );
  NOR2_X1 U19751 ( .A1(n16505), .A2(n16504), .ZN(n16503) );
  INV_X1 U19752 ( .A(n18608), .ZN(n16820) );
  NAND2_X1 U19753 ( .A1(n9795), .A2(n16820), .ZN(n16828) );
  NOR3_X1 U19754 ( .A1(n16494), .A2(n16493), .A3(n16828), .ZN(n16486) );
  NOR2_X1 U19755 ( .A1(n20831), .A2(n16482), .ZN(n16519) );
  NAND4_X1 U19756 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16519), .ZN(n16487) );
  NAND2_X1 U19757 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n18688), .ZN(n16483) );
  OAI22_X1 U19758 ( .A1(n16484), .A2(n16827), .B1(n16487), .B2(n16483), .ZN(
        n16485) );
  AOI211_X1 U19759 ( .C1(n16818), .C2(P3_EBX_REG_31__SCAN_IN), .A(n16486), .B(
        n16485), .ZN(n16490) );
  NOR2_X1 U19760 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16487), .ZN(n16496) );
  NOR2_X1 U19761 ( .A1(n16826), .A2(n16813), .ZN(n16653) );
  INV_X1 U19762 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18684) );
  INV_X1 U19763 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18685) );
  INV_X1 U19764 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n20825) );
  NOR3_X1 U19765 ( .A1(n18684), .A2(n18685), .A3(n20825), .ZN(n16488) );
  OAI21_X1 U19766 ( .B1(n16653), .B2(n16488), .A(n16532), .ZN(n16508) );
  OAI21_X1 U19767 ( .B1(n16496), .B2(n16508), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n16489) );
  OAI211_X1 U19768 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16491), .A(n16490), .B(
        n16489), .ZN(P3_U2640) );
  NAND2_X1 U19769 ( .A1(n16840), .A2(n16492), .ZN(n16501) );
  AOI21_X1 U19770 ( .B1(P3_REIP_REG_30__SCAN_IN), .B2(n16508), .A(n16496), 
        .ZN(n16497) );
  OAI211_X1 U19771 ( .C1(n16827), .C2(n16499), .A(n16498), .B(n16497), .ZN(
        P3_U2641) );
  NOR3_X1 U19772 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n18684), .A3(n20825), 
        .ZN(n16500) );
  AOI22_X1 U19773 ( .A1(n16841), .A2(P3_EBX_REG_29__SCAN_IN), .B1(n16519), 
        .B2(n16500), .ZN(n16510) );
  AOI21_X1 U19774 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16502), .A(n16501), .ZN(
        n16507) );
  AOI211_X1 U19775 ( .C1(n16505), .C2(n16504), .A(n16503), .B(n18608), .ZN(
        n16506) );
  AOI211_X1 U19776 ( .C1(P3_REIP_REG_29__SCAN_IN), .C2(n16508), .A(n16507), 
        .B(n16506), .ZN(n16509) );
  OAI211_X1 U19777 ( .C1(n16511), .C2(n16827), .A(n16510), .B(n16509), .ZN(
        P3_U2642) );
  AOI22_X1 U19778 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16791), .B1(
        n16841), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16522) );
  AOI211_X1 U19779 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16528), .A(n16512), .B(
        n16838), .ZN(n16518) );
  NAND2_X1 U19780 ( .A1(n16519), .A2(n20825), .ZN(n16525) );
  AOI21_X1 U19781 ( .B1(n16532), .B2(n16525), .A(n18684), .ZN(n16517) );
  AOI211_X1 U19782 ( .C1(n16515), .C2(n16514), .A(n16513), .B(n18608), .ZN(
        n16516) );
  NOR3_X1 U19783 ( .A1(n16518), .A2(n16517), .A3(n16516), .ZN(n16521) );
  NAND3_X1 U19784 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16519), .A3(n18684), 
        .ZN(n16520) );
  NAND3_X1 U19785 ( .A1(n16522), .A2(n16521), .A3(n16520), .ZN(P3_U2643) );
  AOI211_X1 U19786 ( .C1(n17430), .C2(n16524), .A(n16523), .B(n18608), .ZN(
        n16527) );
  OAI21_X1 U19787 ( .B1(n16827), .B2(n20847), .A(n16525), .ZN(n16526) );
  AOI211_X1 U19788 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n16841), .A(n16527), .B(
        n16526), .ZN(n16531) );
  OAI211_X1 U19789 ( .C1(n16529), .C2(n16889), .A(n16840), .B(n16528), .ZN(
        n16530) );
  OAI211_X1 U19790 ( .C1(n16532), .C2(n20825), .A(n16531), .B(n16530), .ZN(
        P3_U2644) );
  AOI22_X1 U19791 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n16791), .B1(
        n16818), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n16541) );
  NOR2_X1 U19792 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16831), .ZN(n16542) );
  INV_X1 U19793 ( .A(n16554), .ZN(n16562) );
  OAI221_X1 U19794 ( .B1(n16831), .B2(P3_REIP_REG_23__SCAN_IN), .C1(n16831), 
        .C2(n16562), .A(n16842), .ZN(n16557) );
  AOI211_X1 U19795 ( .C1(n17448), .C2(n16533), .A(n9690), .B(n18608), .ZN(
        n16534) );
  AOI221_X1 U19796 ( .B1(n16542), .B2(P3_REIP_REG_25__SCAN_IN), .C1(n16557), 
        .C2(P3_REIP_REG_25__SCAN_IN), .A(n16534), .ZN(n16540) );
  OAI211_X1 U19797 ( .C1(n16544), .C2(n16536), .A(n16840), .B(n16535), .ZN(
        n16539) );
  INV_X1 U19798 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18679) );
  NAND3_X1 U19799 ( .A1(n16813), .A2(n16537), .A3(n18679), .ZN(n16538) );
  NAND4_X1 U19800 ( .A1(n16541), .A2(n16540), .A3(n16539), .A4(n16538), .ZN(
        P3_U2646) );
  INV_X1 U19801 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17462) );
  AOI22_X1 U19802 ( .A1(n16841), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16543), 
        .B2(n16542), .ZN(n16551) );
  AOI211_X1 U19803 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16558), .A(n16544), .B(
        n16838), .ZN(n16549) );
  AOI211_X1 U19804 ( .C1(n16547), .C2(n16546), .A(n16545), .B(n18608), .ZN(
        n16548) );
  AOI211_X1 U19805 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16557), .A(n16549), 
        .B(n16548), .ZN(n16550) );
  OAI211_X1 U19806 ( .C1(n17462), .C2(n16827), .A(n16551), .B(n16550), .ZN(
        P3_U2647) );
  AOI22_X1 U19807 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n16791), .B1(
        n16841), .B2(P3_EBX_REG_23__SCAN_IN), .ZN(n16561) );
  AOI211_X1 U19808 ( .C1(n17473), .C2(n16553), .A(n16552), .B(n18608), .ZN(
        n16556) );
  NOR3_X1 U19809 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16831), .A3(n16554), 
        .ZN(n16555) );
  AOI211_X1 U19810 ( .C1(n16557), .C2(P3_REIP_REG_23__SCAN_IN), .A(n16556), 
        .B(n16555), .ZN(n16560) );
  OAI211_X1 U19811 ( .C1(n16563), .C2(n16847), .A(n16840), .B(n16558), .ZN(
        n16559) );
  NAND3_X1 U19812 ( .A1(n16561), .A2(n16560), .A3(n16559), .ZN(P3_U2648) );
  AOI22_X1 U19813 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n16791), .B1(
        n16841), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n16571) );
  AOI21_X1 U19814 ( .B1(n16562), .B2(n16842), .A(n16653), .ZN(n16569) );
  INV_X1 U19815 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18673) );
  NAND2_X1 U19816 ( .A1(n16813), .A2(n16572), .ZN(n16581) );
  INV_X1 U19817 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18674) );
  OAI21_X1 U19818 ( .B1(n18673), .B2(n16581), .A(n18674), .ZN(n16568) );
  AOI211_X1 U19819 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16578), .A(n16563), .B(
        n16838), .ZN(n16567) );
  AOI211_X1 U19820 ( .C1(n17491), .C2(n16565), .A(n16564), .B(n18608), .ZN(
        n16566) );
  AOI211_X1 U19821 ( .C1(n16569), .C2(n16568), .A(n16567), .B(n16566), .ZN(
        n16570) );
  NAND2_X1 U19822 ( .A1(n16571), .A2(n16570), .ZN(P3_U2649) );
  OAI21_X1 U19823 ( .B1(n16572), .B2(n16831), .A(n16842), .ZN(n16588) );
  AOI211_X1 U19824 ( .C1(n16575), .C2(n16574), .A(n16573), .B(n18608), .ZN(
        n16577) );
  INV_X1 U19825 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17505) );
  OAI22_X1 U19826 ( .A1(n17505), .A2(n16827), .B1(n16830), .B2(n16936), .ZN(
        n16576) );
  AOI211_X1 U19827 ( .C1(n16588), .C2(P3_REIP_REG_21__SCAN_IN), .A(n16577), 
        .B(n16576), .ZN(n16580) );
  OAI211_X1 U19828 ( .C1(n16584), .C2(n16936), .A(n16840), .B(n16578), .ZN(
        n16579) );
  OAI211_X1 U19829 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n16581), .A(n16580), 
        .B(n16579), .ZN(P3_U2650) );
  AOI22_X1 U19830 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n16791), .B1(
        n16841), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n16590) );
  NAND2_X1 U19831 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n16601) );
  NAND2_X1 U19832 ( .A1(n16813), .A2(n16591), .ZN(n16600) );
  INV_X1 U19833 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18671) );
  OAI21_X1 U19834 ( .B1(n16601), .B2(n16600), .A(n18671), .ZN(n16587) );
  AOI211_X1 U19835 ( .C1(n17519), .C2(n16583), .A(n16582), .B(n18608), .ZN(
        n16586) );
  AOI211_X1 U19836 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16598), .A(n16584), .B(
        n16838), .ZN(n16585) );
  AOI211_X1 U19837 ( .C1(n16588), .C2(n16587), .A(n16586), .B(n16585), .ZN(
        n16589) );
  NAND2_X1 U19838 ( .A1(n16590), .A2(n16589), .ZN(P3_U2651) );
  OAI21_X1 U19839 ( .B1(n16591), .B2(n16831), .A(n16842), .ZN(n16619) );
  INV_X1 U19840 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16595) );
  NOR2_X1 U19841 ( .A1(n16834), .A2(n17533), .ZN(n17530) );
  NAND2_X1 U19842 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17530), .ZN(
        n16592) );
  AOI21_X1 U19843 ( .B1(n16595), .B2(n16592), .A(n17488), .ZN(n17531) );
  OAI21_X1 U19844 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17530), .A(
        n16592), .ZN(n17545) );
  INV_X1 U19845 ( .A(n17545), .ZN(n16607) );
  AOI21_X1 U19846 ( .B1(n17530), .B2(n16638), .A(n9794), .ZN(n16606) );
  NOR2_X1 U19847 ( .A1(n16607), .A2(n16606), .ZN(n16605) );
  NOR2_X1 U19848 ( .A1(n16605), .A2(n9794), .ZN(n16594) );
  OAI21_X1 U19849 ( .B1(n17531), .B2(n16594), .A(n16820), .ZN(n16593) );
  AOI21_X1 U19850 ( .B1(n17531), .B2(n16594), .A(n16593), .ZN(n16597) );
  OAI22_X1 U19851 ( .A1(n16595), .A2(n16827), .B1(n16830), .B2(n16599), .ZN(
        n16596) );
  AOI211_X1 U19852 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(n16619), .A(n16597), 
        .B(n16596), .ZN(n16604) );
  OAI211_X1 U19853 ( .C1(n16608), .C2(n16599), .A(n16840), .B(n16598), .ZN(
        n16603) );
  INV_X1 U19854 ( .A(n16600), .ZN(n16612) );
  OAI211_X1 U19855 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(P3_REIP_REG_18__SCAN_IN), .A(n16612), .B(n16601), .ZN(n16602) );
  NAND4_X1 U19856 ( .A1(n16604), .A2(n18069), .A3(n16603), .A4(n16602), .ZN(
        P3_U2652) );
  AOI211_X1 U19857 ( .C1(n16607), .C2(n16606), .A(n16605), .B(n18608), .ZN(
        n16610) );
  AOI211_X1 U19858 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16622), .A(n16608), .B(
        n16838), .ZN(n16609) );
  AOI211_X1 U19859 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16841), .A(n16610), .B(
        n16609), .ZN(n16614) );
  INV_X1 U19860 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18666) );
  INV_X1 U19861 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17548) );
  OAI21_X1 U19862 ( .B1(n17548), .B2(n16827), .A(n18069), .ZN(n16611) );
  AOI221_X1 U19863 ( .B1(n16612), .B2(n18666), .C1(n16619), .C2(
        P3_REIP_REG_18__SCAN_IN), .A(n16611), .ZN(n16613) );
  NAND2_X1 U19864 ( .A1(n16614), .A2(n16613), .ZN(P3_U2653) );
  AOI22_X1 U19865 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16791), .B1(
        n16841), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n16626) );
  INV_X1 U19866 ( .A(n16639), .ZN(n16616) );
  NAND2_X1 U19867 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16616), .ZN(
        n16615) );
  AOI21_X1 U19868 ( .B1(n9798), .B2(n16615), .A(n17530), .ZN(n17558) );
  OAI21_X1 U19869 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16616), .A(
        n16615), .ZN(n17572) );
  AOI21_X1 U19870 ( .B1(n16638), .B2(n17572), .A(n9794), .ZN(n16617) );
  XOR2_X1 U19871 ( .A(n17558), .B(n16617), .Z(n16621) );
  NOR3_X1 U19872 ( .A1(n16831), .A2(n16652), .A3(n16618), .ZN(n16643) );
  NAND2_X1 U19873 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16643), .ZN(n16637) );
  OAI21_X1 U19874 ( .B1(n18662), .B2(n16637), .A(n18664), .ZN(n16620) );
  AOI22_X1 U19875 ( .A1(n16820), .A2(n16621), .B1(n16620), .B2(n16619), .ZN(
        n16625) );
  OAI211_X1 U19876 ( .C1(n16631), .C2(n16623), .A(n16840), .B(n16622), .ZN(
        n16624) );
  NAND4_X1 U19877 ( .A1(n16626), .A2(n16625), .A3(n18069), .A4(n16624), .ZN(
        P3_U2654) );
  AOI21_X1 U19878 ( .B1(n16813), .B2(n16627), .A(n16826), .ZN(n16641) );
  INV_X1 U19879 ( .A(n17572), .ZN(n16630) );
  NOR2_X1 U19880 ( .A1(n16638), .A2(n9794), .ZN(n16629) );
  INV_X1 U19881 ( .A(n16629), .ZN(n16628) );
  AOI221_X1 U19882 ( .B1(n16630), .B2(n16629), .C1(n17572), .C2(n16628), .A(
        n18608), .ZN(n16635) );
  AOI211_X1 U19883 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16645), .A(n16631), .B(
        n16838), .ZN(n16634) );
  AOI22_X1 U19884 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16791), .B1(
        n16841), .B2(P3_EBX_REG_16__SCAN_IN), .ZN(n16632) );
  INV_X1 U19885 ( .A(n16632), .ZN(n16633) );
  NOR4_X1 U19886 ( .A1(n17985), .A2(n16635), .A3(n16634), .A4(n16633), .ZN(
        n16636) );
  OAI221_X1 U19887 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(n16637), .C1(n18662), 
        .C2(n16641), .A(n16636), .ZN(P3_U2655) );
  AOI22_X1 U19888 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n16791), .B1(
        n16841), .B2(P3_EBX_REG_15__SCAN_IN), .ZN(n16649) );
  NOR2_X1 U19889 ( .A1(n16638), .A2(n16828), .ZN(n16640) );
  OAI21_X1 U19890 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17567), .A(
        n16639), .ZN(n17577) );
  AOI21_X1 U19891 ( .B1(n16640), .B2(n17577), .A(n9612), .ZN(n16648) );
  INV_X1 U19892 ( .A(n16641), .ZN(n16644) );
  NAND2_X1 U19893 ( .A1(n16820), .A2(n9794), .ZN(n16824) );
  INV_X1 U19894 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16829) );
  OAI21_X1 U19895 ( .B1(n9794), .B2(n16829), .A(n16820), .ZN(n16761) );
  AOI211_X1 U19896 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n16824), .A(
        n16761), .B(n17577), .ZN(n16642) );
  AOI221_X1 U19897 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16644), .C1(n16643), 
        .C2(n16644), .A(n16642), .ZN(n16647) );
  OAI211_X1 U19898 ( .C1(n16656), .C2(n17018), .A(n16840), .B(n16645), .ZN(
        n16646) );
  NAND4_X1 U19899 ( .A1(n16649), .A2(n16648), .A3(n16647), .A4(n16646), .ZN(
        P3_U2656) );
  OAI21_X1 U19900 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16664), .A(
        n16650), .ZN(n17593) );
  NOR2_X1 U19901 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16834), .ZN(
        n16821) );
  NAND2_X1 U19902 ( .A1(n17592), .A2(n16821), .ZN(n16667) );
  NAND2_X1 U19903 ( .A1(n9795), .A2(n16667), .ZN(n16651) );
  XNOR2_X1 U19904 ( .A(n17593), .B(n16651), .ZN(n16661) );
  AOI21_X1 U19905 ( .B1(n16841), .B2(P3_EBX_REG_14__SCAN_IN), .A(n9612), .ZN(
        n16660) );
  NOR2_X1 U19906 ( .A1(n16831), .A2(n16652), .ZN(n16662) );
  INV_X1 U19907 ( .A(n16653), .ZN(n16839) );
  AOI22_X1 U19908 ( .A1(n16662), .A2(P3_REIP_REG_13__SCAN_IN), .B1(
        P3_REIP_REG_14__SCAN_IN), .B2(n16839), .ZN(n16654) );
  AOI21_X1 U19909 ( .B1(n16655), .B2(n16842), .A(n16654), .ZN(n16658) );
  AOI211_X1 U19910 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16668), .A(n16656), .B(
        n16838), .ZN(n16657) );
  AOI211_X1 U19911 ( .C1(n16791), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16658), .B(n16657), .ZN(n16659) );
  OAI211_X1 U19912 ( .C1(n18608), .C2(n16661), .A(n16660), .B(n16659), .ZN(
        P3_U2657) );
  INV_X1 U19913 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18656) );
  AOI22_X1 U19914 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n16791), .B1(
        n16662), .B2(n18656), .ZN(n16675) );
  AOI21_X1 U19915 ( .B1(n16813), .B2(n16663), .A(n16826), .ZN(n16696) );
  OAI21_X1 U19916 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n16831), .A(n16696), 
        .ZN(n16673) );
  INV_X1 U19917 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17625) );
  NOR2_X1 U19918 ( .A1(n17625), .A2(n16691), .ZN(n16666) );
  INV_X1 U19919 ( .A(n16666), .ZN(n16677) );
  INV_X1 U19920 ( .A(n16664), .ZN(n16665) );
  OAI21_X1 U19921 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16666), .A(
        n16665), .ZN(n17616) );
  AOI211_X1 U19922 ( .C1(n16677), .C2(n16824), .A(n16761), .B(n17616), .ZN(
        n16672) );
  NAND2_X1 U19923 ( .A1(n17616), .A2(n16667), .ZN(n16670) );
  OAI211_X1 U19924 ( .C1(n16681), .C2(n16676), .A(n16840), .B(n16668), .ZN(
        n16669) );
  OAI211_X1 U19925 ( .C1(n16828), .C2(n16670), .A(n18069), .B(n16669), .ZN(
        n16671) );
  AOI211_X1 U19926 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16673), .A(n16672), 
        .B(n16671), .ZN(n16674) );
  OAI211_X1 U19927 ( .C1(n16830), .C2(n16676), .A(n16675), .B(n16674), .ZN(
        P3_U2658) );
  OAI21_X1 U19928 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17612), .A(
        n16677), .ZN(n17621) );
  NAND2_X1 U19929 ( .A1(n17672), .A2(n16821), .ZN(n16741) );
  INV_X1 U19930 ( .A(n16741), .ZN(n16692) );
  AOI21_X1 U19931 ( .B1(n16679), .B2(n16692), .A(n16678), .ZN(n16680) );
  XOR2_X1 U19932 ( .A(n17621), .B(n16680), .Z(n16688) );
  AOI211_X1 U19933 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16698), .A(n16681), .B(
        n16838), .ZN(n16686) );
  INV_X1 U19934 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18655) );
  NOR2_X1 U19935 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16831), .ZN(n16682) );
  AOI22_X1 U19936 ( .A1(n16841), .A2(P3_EBX_REG_12__SCAN_IN), .B1(n16683), 
        .B2(n16682), .ZN(n16684) );
  OAI211_X1 U19937 ( .C1(n16696), .C2(n18655), .A(n16684), .B(n18069), .ZN(
        n16685) );
  AOI211_X1 U19938 ( .C1(n16791), .C2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16686), .B(n16685), .ZN(n16687) );
  OAI21_X1 U19939 ( .B1(n18608), .B2(n16688), .A(n16687), .ZN(P3_U2659) );
  AND2_X1 U19940 ( .A1(n16813), .A2(n16702), .ZN(n16711) );
  AOI21_X1 U19941 ( .B1(n16689), .B2(n16711), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16695) );
  NAND2_X1 U19942 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17672), .ZN(
        n16739) );
  NOR2_X1 U19943 ( .A1(n16690), .A2(n16739), .ZN(n16707) );
  OAI21_X1 U19944 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16707), .A(
        n16691), .ZN(n17639) );
  AOI21_X1 U19945 ( .B1(n16693), .B2(n16692), .A(n9794), .ZN(n16710) );
  XOR2_X1 U19946 ( .A(n17639), .B(n16710), .Z(n16694) );
  OAI22_X1 U19947 ( .A1(n16696), .A2(n16695), .B1(n18608), .B2(n16694), .ZN(
        n16697) );
  AOI211_X1 U19948 ( .C1(n16818), .C2(P3_EBX_REG_11__SCAN_IN), .A(n9612), .B(
        n16697), .ZN(n16700) );
  OAI211_X1 U19949 ( .C1(n16704), .C2(n17064), .A(n16840), .B(n16698), .ZN(
        n16699) );
  OAI211_X1 U19950 ( .C1(n16827), .C2(n16701), .A(n16700), .B(n16699), .ZN(
        P3_U2660) );
  AOI22_X1 U19951 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16791), .B1(
        n16841), .B2(P3_EBX_REG_10__SCAN_IN), .ZN(n16715) );
  OAI21_X1 U19952 ( .B1(n16831), .B2(n16702), .A(n16842), .ZN(n16727) );
  INV_X1 U19953 ( .A(n16727), .ZN(n16703) );
  NAND2_X1 U19954 ( .A1(n16711), .A2(n18648), .ZN(n16719) );
  NAND2_X1 U19955 ( .A1(n16703), .A2(n16719), .ZN(n16706) );
  AOI211_X1 U19956 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16722), .A(n16704), .B(
        n16838), .ZN(n16705) );
  AOI211_X1 U19957 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(n16706), .A(n9612), .B(
        n16705), .ZN(n16714) );
  NOR2_X1 U19958 ( .A1(n17680), .A2(n16739), .ZN(n16729) );
  NAND2_X1 U19959 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16729), .ZN(
        n16716) );
  AOI21_X1 U19960 ( .B1(n16708), .B2(n16716), .A(n16707), .ZN(n17654) );
  INV_X1 U19961 ( .A(n16824), .ZN(n16733) );
  OR2_X1 U19962 ( .A1(n17680), .A2(n16741), .ZN(n16717) );
  AOI221_X1 U19963 ( .B1(n17662), .B2(n17654), .C1(n16717), .C2(n17654), .A(
        n18608), .ZN(n16709) );
  OAI22_X1 U19964 ( .A1(n17654), .A2(n16710), .B1(n16733), .B2(n16709), .ZN(
        n16713) );
  NAND3_X1 U19965 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16711), .A3(n18650), 
        .ZN(n16712) );
  NAND4_X1 U19966 ( .A1(n16715), .A2(n16714), .A3(n16713), .A4(n16712), .ZN(
        P3_U2661) );
  OAI21_X1 U19967 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16729), .A(
        n16716), .ZN(n17659) );
  NAND2_X1 U19968 ( .A1(n9795), .A2(n16717), .ZN(n16731) );
  OAI21_X1 U19969 ( .B1(n17659), .B2(n16731), .A(n16820), .ZN(n16718) );
  AOI21_X1 U19970 ( .B1(n17659), .B2(n16731), .A(n16718), .ZN(n16721) );
  OAI211_X1 U19971 ( .C1(n16830), .C2(n17049), .A(n18069), .B(n16719), .ZN(
        n16720) );
  AOI211_X1 U19972 ( .C1(P3_REIP_REG_9__SCAN_IN), .C2(n16727), .A(n16721), .B(
        n16720), .ZN(n16724) );
  OAI211_X1 U19973 ( .C1(n16725), .C2(n17049), .A(n16840), .B(n16722), .ZN(
        n16723) );
  OAI211_X1 U19974 ( .C1(n16827), .C2(n17662), .A(n16724), .B(n16723), .ZN(
        P3_U2662) );
  AOI22_X1 U19975 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16791), .B1(
        n16841), .B2(P3_EBX_REG_8__SCAN_IN), .ZN(n16738) );
  AOI211_X1 U19976 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16748), .A(n16725), .B(
        n16838), .ZN(n16726) );
  AOI211_X1 U19977 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n16727), .A(n9612), .B(
        n16726), .ZN(n16737) );
  NOR2_X1 U19978 ( .A1(n16831), .A2(n16742), .ZN(n16728) );
  NAND4_X1 U19979 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .A3(n16728), .A4(n18647), .ZN(n16736) );
  INV_X1 U19980 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16730) );
  NAND3_X1 U19981 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17672), .A3(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16740) );
  AOI21_X1 U19982 ( .B1(n16730), .B2(n16740), .A(n16729), .ZN(n17673) );
  INV_X1 U19983 ( .A(n16731), .ZN(n16734) );
  INV_X1 U19984 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17687) );
  AOI221_X1 U19985 ( .B1(n17687), .B2(n17673), .C1(n16741), .C2(n17673), .A(
        n18608), .ZN(n16732) );
  OAI22_X1 U19986 ( .A1(n17673), .A2(n16734), .B1(n16733), .B2(n16732), .ZN(
        n16735) );
  NAND4_X1 U19987 ( .A1(n16738), .A2(n16737), .A3(n16736), .A4(n16735), .ZN(
        P3_U2663) );
  INV_X1 U19988 ( .A(n16739), .ZN(n16753) );
  OAI21_X1 U19989 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16753), .A(
        n16740), .ZN(n17697) );
  NAND2_X1 U19990 ( .A1(n9795), .A2(n16741), .ZN(n16755) );
  XOR2_X1 U19991 ( .A(n17697), .B(n16755), .Z(n16747) );
  INV_X1 U19992 ( .A(n16742), .ZN(n16743) );
  NOR2_X1 U19993 ( .A1(n16743), .A2(n16831), .ZN(n16766) );
  NOR2_X1 U19994 ( .A1(n16826), .A2(n16766), .ZN(n16769) );
  NAND3_X1 U19995 ( .A1(n16743), .A2(n16813), .A3(n18642), .ZN(n16757) );
  AOI21_X1 U19996 ( .B1(n16769), .B2(n16757), .A(n18644), .ZN(n16746) );
  NAND4_X1 U19997 ( .A1(n16743), .A2(n16813), .A3(P3_REIP_REG_6__SCAN_IN), 
        .A4(n18644), .ZN(n16744) );
  OAI211_X1 U19998 ( .C1(n16830), .C2(n16749), .A(n18069), .B(n16744), .ZN(
        n16745) );
  AOI211_X1 U19999 ( .C1(n16820), .C2(n16747), .A(n16746), .B(n16745), .ZN(
        n16751) );
  OAI211_X1 U20000 ( .C1(n16752), .C2(n16749), .A(n16840), .B(n16748), .ZN(
        n16750) );
  OAI211_X1 U20001 ( .C1(n16827), .C2(n17687), .A(n16751), .B(n16750), .ZN(
        P3_U2664) );
  AOI211_X1 U20002 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16772), .A(n16752), .B(
        n16838), .ZN(n16760) );
  NOR2_X1 U20003 ( .A1(n16834), .A2(n17700), .ZN(n16764) );
  INV_X1 U20004 ( .A(n16764), .ZN(n16754) );
  AOI21_X1 U20005 ( .B1(n17707), .B2(n16754), .A(n16753), .ZN(n17704) );
  NOR3_X1 U20006 ( .A1(n17704), .A2(n18608), .A3(n16755), .ZN(n16756) );
  NOR2_X1 U20007 ( .A1(n16756), .A2(n9612), .ZN(n16758) );
  OAI211_X1 U20008 ( .C1(n16769), .C2(n18642), .A(n16758), .B(n16757), .ZN(
        n16759) );
  AOI211_X1 U20009 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16818), .A(n16760), .B(
        n16759), .ZN(n16763) );
  INV_X1 U20010 ( .A(n16761), .ZN(n16833) );
  OAI211_X1 U20011 ( .C1(n16764), .C2(n9794), .A(n17704), .B(n16833), .ZN(
        n16762) );
  OAI211_X1 U20012 ( .C1(n16827), .C2(n17707), .A(n16763), .B(n16762), .ZN(
        P3_U2665) );
  INV_X1 U20013 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16765) );
  NAND2_X1 U20014 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17708), .ZN(
        n16780) );
  AOI21_X1 U20015 ( .B1(n16765), .B2(n16780), .A(n16764), .ZN(n17713) );
  OAI21_X1 U20016 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16780), .A(
        n9795), .ZN(n16785) );
  XNOR2_X1 U20017 ( .A(n17713), .B(n16785), .ZN(n16771) );
  INV_X1 U20018 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18641) );
  AOI22_X1 U20019 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n16791), .B1(
        n16767), .B2(n16766), .ZN(n16768) );
  OAI211_X1 U20020 ( .C1(n16769), .C2(n18641), .A(n16768), .B(n18069), .ZN(
        n16770) );
  AOI21_X1 U20021 ( .B1(n16820), .B2(n16771), .A(n16770), .ZN(n16774) );
  OAI211_X1 U20022 ( .C1(n16779), .C2(n16775), .A(n16840), .B(n16772), .ZN(
        n16773) );
  OAI211_X1 U20023 ( .C1(n16775), .C2(n16830), .A(n16774), .B(n16773), .ZN(
        P3_U2666) );
  NOR2_X1 U20024 ( .A1(n16776), .A2(n18743), .ZN(n18767) );
  INV_X1 U20025 ( .A(n18767), .ZN(n16777) );
  AOI21_X1 U20026 ( .B1(n9645), .B2(n18540), .A(n16777), .ZN(n16778) );
  AOI211_X1 U20027 ( .C1(n16841), .C2(P3_EBX_REG_4__SCAN_IN), .A(n9612), .B(
        n16778), .ZN(n16790) );
  AOI211_X1 U20028 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16800), .A(n16779), .B(
        n16838), .ZN(n16783) );
  NAND2_X1 U20029 ( .A1(n16813), .A2(n16792), .ZN(n16781) );
  NOR2_X1 U20030 ( .A1(n16834), .A2(n17725), .ZN(n16795) );
  OAI21_X1 U20031 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16795), .A(
        n16780), .ZN(n17728) );
  OAI22_X1 U20032 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16781), .B1(n16824), 
        .B2(n17728), .ZN(n16782) );
  AOI211_X1 U20033 ( .C1(n16791), .C2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n16783), .B(n16782), .ZN(n16789) );
  INV_X1 U20034 ( .A(n17728), .ZN(n16786) );
  INV_X1 U20035 ( .A(n16821), .ZN(n16784) );
  OR2_X1 U20036 ( .A1(n17725), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17732) );
  OAI22_X1 U20037 ( .A1(n16786), .A2(n16785), .B1(n16784), .B2(n17732), .ZN(
        n16787) );
  OAI21_X1 U20038 ( .B1(n16792), .B2(n16831), .A(n16842), .ZN(n16798) );
  AOI22_X1 U20039 ( .A1(n16820), .A2(n16787), .B1(P3_REIP_REG_4__SCAN_IN), 
        .B2(n16798), .ZN(n16788) );
  NAND3_X1 U20040 ( .A1(n16790), .A2(n16789), .A3(n16788), .ZN(P3_U2667) );
  AOI22_X1 U20041 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n16791), .B1(
        n16841), .B2(P3_EBX_REG_3__SCAN_IN), .ZN(n16805) );
  INV_X1 U20042 ( .A(n16812), .ZN(n16794) );
  NOR2_X1 U20043 ( .A1(n16792), .A2(n16831), .ZN(n16793) );
  NOR3_X1 U20044 ( .A1(n9610), .A2(n20898), .A3(n18717), .ZN(n16809) );
  INV_X1 U20045 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18554) );
  OAI21_X1 U20046 ( .B1(n16809), .B2(n18554), .A(n9599), .ZN(n18705) );
  AOI22_X1 U20047 ( .A1(n16794), .A2(n16793), .B1(n18767), .B2(n18705), .ZN(
        n16804) );
  INV_X1 U20048 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16796) );
  NAND2_X1 U20049 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16806) );
  AOI21_X1 U20050 ( .B1(n16796), .B2(n16806), .A(n16795), .ZN(n17739) );
  AOI21_X1 U20051 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n16821), .A(
        n9794), .ZN(n16819) );
  XOR2_X1 U20052 ( .A(n17739), .B(n16819), .Z(n16799) );
  AOI22_X1 U20053 ( .A1(n16820), .A2(n16799), .B1(P3_REIP_REG_3__SCAN_IN), 
        .B2(n16798), .ZN(n16803) );
  OAI211_X1 U20054 ( .C1(n16807), .C2(n16801), .A(n16840), .B(n16800), .ZN(
        n16802) );
  NAND4_X1 U20055 ( .A1(n16805), .A2(n16804), .A3(n16803), .A4(n16802), .ZN(
        P3_U2668) );
  OAI21_X1 U20056 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16806), .ZN(n17749) );
  OR2_X1 U20057 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), .ZN(
        n16808) );
  AOI211_X1 U20058 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16808), .A(n16807), .B(
        n16838), .ZN(n16817) );
  INV_X1 U20059 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17752) );
  NAND2_X1 U20060 ( .A1(n18717), .A2(n18560), .ZN(n18556) );
  INV_X1 U20061 ( .A(n16809), .ZN(n16810) );
  NAND2_X1 U20062 ( .A1(n18556), .A2(n16810), .ZN(n18711) );
  INV_X1 U20063 ( .A(n18711), .ZN(n16811) );
  AOI22_X1 U20064 ( .A1(n16826), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n16811), 
        .B2(n18767), .ZN(n16815) );
  OAI211_X1 U20065 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16813), .B(n16812), .ZN(n16814) );
  OAI211_X1 U20066 ( .C1(n16827), .C2(n17752), .A(n16815), .B(n16814), .ZN(
        n16816) );
  AOI211_X1 U20067 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16818), .A(n16817), .B(
        n16816), .ZN(n16823) );
  OAI211_X1 U20068 ( .C1(n16821), .C2(n17749), .A(n16820), .B(n16819), .ZN(
        n16822) );
  OAI211_X1 U20069 ( .C1(n16824), .C2(n17749), .A(n16823), .B(n16822), .ZN(
        P3_U2669) );
  NAND2_X1 U20070 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17137) );
  OAI21_X1 U20071 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17137), .ZN(n17144) );
  NAND2_X1 U20072 ( .A1(n18560), .A2(n16825), .ZN(n18572) );
  INV_X1 U20073 ( .A(n18572), .ZN(n18721) );
  AOI22_X1 U20074 ( .A1(n16826), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n18721), 
        .B2(n18767), .ZN(n16837) );
  OAI21_X1 U20075 ( .B1(n16829), .B2(n16828), .A(n16827), .ZN(n16835) );
  INV_X1 U20076 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17143) );
  OAI22_X1 U20077 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16831), .B1(n16830), 
        .B2(n17143), .ZN(n16832) );
  AOI221_X1 U20078 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16835), .C1(
        n16834), .C2(n16833), .A(n16832), .ZN(n16836) );
  OAI211_X1 U20079 ( .C1(n16838), .C2(n17144), .A(n16837), .B(n16836), .ZN(
        P3_U2670) );
  AOI22_X1 U20080 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n16839), .B1(n18767), 
        .B2(n20898), .ZN(n16845) );
  OAI21_X1 U20081 ( .B1(n16841), .B2(n16840), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n16844) );
  NAND3_X1 U20082 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18713), .A3(
        n16842), .ZN(n16843) );
  NAND3_X1 U20083 ( .A1(n16845), .A2(n16844), .A3(n16843), .ZN(P3_U2671) );
  INV_X1 U20084 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16853) );
  NAND3_X1 U20085 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n16878), .ZN(n16846) );
  NOR4_X1 U20086 ( .A1(n16848), .A2(n16847), .A3(n16935), .A4(n16846), .ZN(
        n16849) );
  NAND3_X1 U20087 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16895), .A3(n16849), 
        .ZN(n16852) );
  NOR2_X1 U20088 ( .A1(n16853), .A2(n16852), .ZN(n16877) );
  NAND2_X1 U20089 ( .A1(n17141), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16851) );
  NAND2_X1 U20090 ( .A1(n16877), .A2(n18136), .ZN(n16850) );
  OAI22_X1 U20091 ( .A1(n16877), .A2(n16851), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16850), .ZN(P3_U2672) );
  NAND2_X1 U20092 ( .A1(n16853), .A2(n16852), .ZN(n16854) );
  NAND2_X1 U20093 ( .A1(n16854), .A2(n17141), .ZN(n16876) );
  AOI22_X1 U20094 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17081), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16858) );
  AOI22_X1 U20095 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16857) );
  AOI22_X1 U20096 ( .A1(n17067), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16856) );
  AOI22_X1 U20097 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n15741), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16855) );
  NAND4_X1 U20098 ( .A1(n16858), .A2(n16857), .A3(n16856), .A4(n16855), .ZN(
        n16864) );
  AOI22_X1 U20099 ( .A1(n17107), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16862) );
  AOI22_X1 U20100 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17053), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16861) );
  AOI22_X1 U20101 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16860) );
  AOI22_X1 U20102 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16859) );
  NAND4_X1 U20103 ( .A1(n16862), .A2(n16861), .A3(n16860), .A4(n16859), .ZN(
        n16863) );
  NOR2_X1 U20104 ( .A1(n16864), .A2(n16863), .ZN(n16881) );
  NOR2_X1 U20105 ( .A1(n16881), .A2(n16880), .ZN(n16879) );
  AOI22_X1 U20106 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16868) );
  AOI22_X1 U20107 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16867) );
  AOI22_X1 U20108 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16866) );
  AOI22_X1 U20109 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16865) );
  NAND4_X1 U20110 ( .A1(n16868), .A2(n16867), .A3(n16866), .A4(n16865), .ZN(
        n16874) );
  AOI22_X1 U20111 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15741), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16872) );
  AOI22_X1 U20112 ( .A1(n17107), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17081), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16871) );
  AOI22_X1 U20113 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16870) );
  AOI22_X1 U20114 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16869) );
  NAND4_X1 U20115 ( .A1(n16872), .A2(n16871), .A3(n16870), .A4(n16869), .ZN(
        n16873) );
  NOR2_X1 U20116 ( .A1(n16874), .A2(n16873), .ZN(n16875) );
  XOR2_X1 U20117 ( .A(n16879), .B(n16875), .Z(n17158) );
  OAI22_X1 U20118 ( .A1(n16877), .A2(n16876), .B1(n17158), .B2(n17141), .ZN(
        P3_U2673) );
  NAND2_X1 U20119 ( .A1(n16887), .A2(n16878), .ZN(n16884) );
  AOI21_X1 U20120 ( .B1(n16881), .B2(n16880), .A(n16879), .ZN(n17160) );
  AOI22_X1 U20121 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16882), .B1(n17160), 
        .B2(n17146), .ZN(n16883) );
  OAI21_X1 U20122 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16884), .A(n16883), .ZN(
        P3_U2674) );
  AOI21_X1 U20123 ( .B1(n16886), .B2(n16890), .A(n16885), .ZN(n17170) );
  AOI22_X1 U20124 ( .A1(n17170), .A2(n17146), .B1(n16887), .B2(n16889), .ZN(
        n16888) );
  OAI21_X1 U20125 ( .B1(n16889), .B2(n16893), .A(n16888), .ZN(P3_U2676) );
  OAI21_X1 U20126 ( .B1(n16892), .B2(n16891), .A(n16890), .ZN(n17178) );
  NAND2_X1 U20127 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n16904), .ZN(n16897) );
  OAI222_X1 U20128 ( .A1(n17178), .A2(n17141), .B1(n16897), .B2(n16895), .C1(
        n16894), .C2(n16893), .ZN(P3_U2677) );
  XNOR2_X1 U20129 ( .A(n16896), .B(n16900), .ZN(n17184) );
  OAI211_X1 U20130 ( .C1(n16904), .C2(P3_EBX_REG_25__SCAN_IN), .A(n17141), .B(
        n16897), .ZN(n16898) );
  OAI21_X1 U20131 ( .B1(n17184), .B2(n17141), .A(n16898), .ZN(P3_U2678) );
  INV_X1 U20132 ( .A(n16899), .ZN(n16909) );
  AOI21_X1 U20133 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17141), .A(n16909), .ZN(
        n16903) );
  OAI21_X1 U20134 ( .B1(n16902), .B2(n16901), .A(n16900), .ZN(n17189) );
  OAI22_X1 U20135 ( .A1(n16904), .A2(n16903), .B1(n17141), .B2(n17189), .ZN(
        P3_U2679) );
  AOI21_X1 U20136 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17141), .A(n16905), .ZN(
        n16908) );
  XNOR2_X1 U20137 ( .A(n16907), .B(n16906), .ZN(n17194) );
  OAI22_X1 U20138 ( .A1(n16909), .A2(n16908), .B1(n17141), .B2(n17194), .ZN(
        P3_U2680) );
  AOI22_X1 U20139 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16920) );
  AOI22_X1 U20140 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n15741), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16919) );
  INV_X1 U20141 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18130) );
  AOI22_X1 U20142 ( .A1(n17104), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9618), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16911) );
  OAI21_X1 U20143 ( .B1(n16940), .B2(n18130), .A(n16911), .ZN(n16917) );
  AOI22_X1 U20144 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16915) );
  AOI22_X1 U20145 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16914) );
  AOI22_X1 U20146 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16913) );
  AOI22_X1 U20147 ( .A1(n17067), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16912) );
  NAND4_X1 U20148 ( .A1(n16915), .A2(n16914), .A3(n16913), .A4(n16912), .ZN(
        n16916) );
  AOI211_X1 U20149 ( .C1(n17087), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n16917), .B(n16916), .ZN(n16918) );
  NAND3_X1 U20150 ( .A1(n16920), .A2(n16919), .A3(n16918), .ZN(n17195) );
  INV_X1 U20151 ( .A(n17195), .ZN(n16922) );
  NAND3_X1 U20152 ( .A1(n16923), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17141), 
        .ZN(n16921) );
  OAI221_X1 U20153 ( .B1(n16923), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17141), 
        .C2(n16922), .A(n16921), .ZN(P3_U2681) );
  AOI22_X1 U20154 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9616), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16927) );
  AOI22_X1 U20155 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9618), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16926) );
  AOI22_X1 U20156 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16925) );
  AOI22_X1 U20157 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17087), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16924) );
  NAND4_X1 U20158 ( .A1(n16927), .A2(n16926), .A3(n16925), .A4(n16924), .ZN(
        n16934) );
  AOI22_X1 U20159 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16932) );
  AOI22_X1 U20160 ( .A1(n17088), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16931) );
  AOI22_X1 U20161 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16930) );
  AOI22_X1 U20162 ( .A1(n17106), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16929) );
  NAND4_X1 U20163 ( .A1(n16932), .A2(n16931), .A3(n16930), .A4(n16929), .ZN(
        n16933) );
  NOR2_X1 U20164 ( .A1(n16934), .A2(n16933), .ZN(n17205) );
  AND2_X1 U20165 ( .A1(n17141), .A2(n16935), .ZN(n16950) );
  AOI22_X1 U20166 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16950), .B1(n16937), 
        .B2(n16936), .ZN(n16938) );
  OAI21_X1 U20167 ( .B1(n17205), .B2(n17141), .A(n16938), .ZN(P3_U2682) );
  AOI22_X1 U20168 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16949) );
  AOI22_X1 U20169 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17087), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16948) );
  AOI22_X1 U20170 ( .A1(n17067), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16939) );
  OAI21_X1 U20171 ( .B1(n16940), .B2(n18122), .A(n16939), .ZN(n16946) );
  AOI22_X1 U20172 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16944) );
  AOI22_X1 U20173 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16943) );
  AOI22_X1 U20174 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17081), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16942) );
  AOI22_X1 U20175 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n15741), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16941) );
  NAND4_X1 U20176 ( .A1(n16944), .A2(n16943), .A3(n16942), .A4(n16941), .ZN(
        n16945) );
  AOI211_X1 U20177 ( .C1(n17105), .C2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n16946), .B(n16945), .ZN(n16947) );
  NAND3_X1 U20178 ( .A1(n16949), .A2(n16948), .A3(n16947), .ZN(n17208) );
  INV_X1 U20179 ( .A(n17208), .ZN(n16952) );
  OAI21_X1 U20180 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16966), .A(n16950), .ZN(
        n16951) );
  OAI21_X1 U20181 ( .B1(n16952), .B2(n17141), .A(n16951), .ZN(P3_U2683) );
  INV_X1 U20182 ( .A(n16977), .ZN(n16953) );
  OAI21_X1 U20183 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n16953), .A(n17141), .ZN(
        n16965) );
  AOI22_X1 U20184 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9618), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16958) );
  AOI22_X1 U20185 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16957) );
  AOI22_X1 U20186 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16956) );
  AOI22_X1 U20187 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16955) );
  NAND4_X1 U20188 ( .A1(n16958), .A2(n16957), .A3(n16956), .A4(n16955), .ZN(
        n16964) );
  AOI22_X1 U20189 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17087), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16962) );
  AOI22_X1 U20190 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17081), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16961) );
  AOI22_X1 U20191 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n16960) );
  AOI22_X1 U20192 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9616), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16959) );
  NAND4_X1 U20193 ( .A1(n16962), .A2(n16961), .A3(n16960), .A4(n16959), .ZN(
        n16963) );
  NOR2_X1 U20194 ( .A1(n16964), .A2(n16963), .ZN(n17218) );
  OAI22_X1 U20195 ( .A1(n16966), .A2(n16965), .B1(n17218), .B2(n17141), .ZN(
        P3_U2684) );
  AOI22_X1 U20196 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n16970) );
  AOI22_X1 U20197 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n15741), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16969) );
  AOI22_X1 U20198 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16968) );
  AOI22_X1 U20199 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16967) );
  NAND4_X1 U20200 ( .A1(n16970), .A2(n16969), .A3(n16968), .A4(n16967), .ZN(
        n16976) );
  AOI22_X1 U20201 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n16974) );
  AOI22_X1 U20202 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n16973) );
  AOI22_X1 U20203 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9618), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16972) );
  AOI22_X1 U20204 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17087), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16971) );
  NAND4_X1 U20205 ( .A1(n16974), .A2(n16973), .A3(n16972), .A4(n16971), .ZN(
        n16975) );
  NOR2_X1 U20206 ( .A1(n16976), .A2(n16975), .ZN(n17223) );
  OAI21_X1 U20207 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n16992), .A(n16977), .ZN(
        n16978) );
  AOI22_X1 U20208 ( .A1(n17146), .A2(n17223), .B1(n16978), .B2(n17141), .ZN(
        P3_U2685) );
  INV_X1 U20209 ( .A(n16979), .ZN(n16980) );
  OAI21_X1 U20210 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n16980), .A(n17141), .ZN(
        n16991) );
  AOI22_X1 U20211 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n17105), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n17089), .ZN(n16984) );
  AOI22_X1 U20212 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17053), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n9614), .ZN(n16983) );
  AOI22_X1 U20213 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17104), .ZN(n16982) );
  AOI22_X1 U20214 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17067), .ZN(n16981) );
  NAND4_X1 U20215 ( .A1(n16984), .A2(n16983), .A3(n16982), .A4(n16981), .ZN(
        n16990) );
  AOI22_X1 U20216 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n17106), .ZN(n16988) );
  AOI22_X1 U20217 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17108), .B1(
        n15741), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16987) );
  AOI22_X1 U20218 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17088), .B1(
        n17090), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n16986) );
  AOI22_X1 U20219 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17087), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n16985) );
  NAND4_X1 U20220 ( .A1(n16988), .A2(n16987), .A3(n16986), .A4(n16985), .ZN(
        n16989) );
  NOR2_X1 U20221 ( .A1(n16990), .A2(n16989), .ZN(n17228) );
  OAI22_X1 U20222 ( .A1(n16992), .A2(n16991), .B1(n17228), .B2(n17141), .ZN(
        P3_U2686) );
  AOI22_X1 U20223 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n16996) );
  AOI22_X1 U20224 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17053), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16995) );
  AOI22_X1 U20225 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n16994) );
  AOI22_X1 U20226 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16993) );
  NAND4_X1 U20227 ( .A1(n16996), .A2(n16995), .A3(n16994), .A4(n16993), .ZN(
        n17002) );
  AOI22_X1 U20228 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9616), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17000) );
  AOI22_X1 U20229 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n16999) );
  AOI22_X1 U20230 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17087), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n16998) );
  AOI22_X1 U20231 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16997) );
  NAND4_X1 U20232 ( .A1(n17000), .A2(n16999), .A3(n16998), .A4(n16997), .ZN(
        n17001) );
  NOR2_X1 U20233 ( .A1(n17002), .A2(n17001), .ZN(n17235) );
  OAI22_X1 U20234 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17240), .B1(n17146), 
        .B2(n17005), .ZN(n17003) );
  OAI21_X1 U20235 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17005), .A(n17003), .ZN(
        n17004) );
  OAI21_X1 U20236 ( .B1(n17235), .B2(n17141), .A(n17004), .ZN(P3_U2687) );
  OR2_X1 U20237 ( .A1(n17146), .A2(n17005), .ZN(n17019) );
  AOI22_X1 U20238 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17016) );
  AOI22_X1 U20239 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n15741), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17015) );
  AOI22_X1 U20240 ( .A1(n17106), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17006) );
  OAI21_X1 U20241 ( .B1(n17007), .B2(n20912), .A(n17006), .ZN(n17013) );
  AOI22_X1 U20242 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17011) );
  AOI22_X1 U20243 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17087), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17010) );
  AOI22_X1 U20244 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17009) );
  AOI22_X1 U20245 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17008) );
  NAND4_X1 U20246 ( .A1(n17011), .A2(n17010), .A3(n17009), .A4(n17008), .ZN(
        n17012) );
  AOI211_X1 U20247 ( .C1(n17117), .C2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n17013), .B(n17012), .ZN(n17014) );
  NAND3_X1 U20248 ( .A1(n17016), .A2(n17015), .A3(n17014), .ZN(n17237) );
  NAND2_X1 U20249 ( .A1(n17146), .A2(n17237), .ZN(n17017) );
  OAI221_X1 U20250 ( .B1(n17019), .B2(n17018), .C1(n17019), .C2(n17031), .A(
        n17017), .ZN(P3_U2688) );
  AOI22_X1 U20251 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17087), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17030) );
  AOI22_X1 U20252 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17029) );
  AOI22_X1 U20253 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17020) );
  OAI21_X1 U20254 ( .B1(n17103), .B2(n18130), .A(n17020), .ZN(n17027) );
  AOI22_X1 U20255 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9616), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17025) );
  AOI22_X1 U20256 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17090), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17024) );
  AOI22_X1 U20257 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17023) );
  AOI22_X1 U20258 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17081), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17022) );
  NAND4_X1 U20259 ( .A1(n17025), .A2(n17024), .A3(n17023), .A4(n17022), .ZN(
        n17026) );
  AOI211_X1 U20260 ( .C1(n17106), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n17027), .B(n17026), .ZN(n17028) );
  NAND3_X1 U20261 ( .A1(n17030), .A2(n17029), .A3(n17028), .ZN(n17244) );
  INV_X1 U20262 ( .A(n17244), .ZN(n17034) );
  OAI21_X1 U20263 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17032), .A(n17031), .ZN(
        n17033) );
  AOI22_X1 U20264 ( .A1(n17146), .A2(n17034), .B1(n17033), .B2(n17141), .ZN(
        P3_U2689) );
  NAND3_X1 U20265 ( .A1(n18136), .A2(n17136), .A3(n17035), .ZN(n17047) );
  AOI22_X1 U20266 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17039) );
  AOI22_X1 U20267 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17053), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17038) );
  AOI22_X1 U20268 ( .A1(n17106), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17037) );
  AOI22_X1 U20269 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17036) );
  NAND4_X1 U20270 ( .A1(n17039), .A2(n17038), .A3(n17037), .A4(n17036), .ZN(
        n17045) );
  AOI22_X1 U20271 ( .A1(n17107), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17088), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17043) );
  AOI22_X1 U20272 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17042) );
  AOI22_X1 U20273 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17081), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17041) );
  AOI22_X1 U20274 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9616), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17040) );
  NAND4_X1 U20275 ( .A1(n17043), .A2(n17042), .A3(n17041), .A4(n17040), .ZN(
        n17044) );
  NOR2_X1 U20276 ( .A1(n17045), .A2(n17044), .ZN(n17254) );
  NAND3_X1 U20277 ( .A1(n17047), .A2(P3_EBX_REG_12__SCAN_IN), .A3(n17141), 
        .ZN(n17046) );
  OAI221_X1 U20278 ( .B1(n17047), .B2(P3_EBX_REG_12__SCAN_IN), .C1(n17141), 
        .C2(n17254), .A(n17046), .ZN(P3_U2691) );
  NAND2_X1 U20279 ( .A1(n17141), .A2(n17047), .ZN(n17065) );
  NAND3_X1 U20280 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(P3_EBX_REG_4__SCAN_IN), 
        .A3(n17136), .ZN(n17126) );
  NOR2_X1 U20281 ( .A1(n17048), .A2(n17126), .ZN(n17125) );
  NAND2_X1 U20282 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17125), .ZN(n17121) );
  NOR2_X1 U20283 ( .A1(n17049), .A2(n17121), .ZN(n17099) );
  NAND2_X1 U20284 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17099), .ZN(n17079) );
  AOI22_X1 U20285 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17062) );
  AOI22_X1 U20286 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17061) );
  AOI22_X1 U20287 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17051) );
  OAI21_X1 U20288 ( .B1(n17052), .B2(n20794), .A(n17051), .ZN(n17059) );
  AOI22_X1 U20289 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n15741), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17057) );
  AOI22_X1 U20290 ( .A1(n17107), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17056) );
  AOI22_X1 U20291 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17053), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17055) );
  AOI22_X1 U20292 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17054) );
  NAND4_X1 U20293 ( .A1(n17057), .A2(n17056), .A3(n17055), .A4(n17054), .ZN(
        n17058) );
  AOI211_X1 U20294 ( .C1(n17082), .C2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A(
        n17059), .B(n17058), .ZN(n17060) );
  NAND3_X1 U20295 ( .A1(n17062), .A2(n17061), .A3(n17060), .ZN(n17258) );
  NAND2_X1 U20296 ( .A1(n17146), .A2(n17258), .ZN(n17063) );
  OAI221_X1 U20297 ( .B1(n17065), .B2(n17064), .C1(n17065), .C2(n17079), .A(
        n17063), .ZN(P3_U2692) );
  AOI22_X1 U20298 ( .A1(n17107), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17081), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17071) );
  AOI22_X1 U20299 ( .A1(n17106), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9616), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17070) );
  AOI22_X1 U20300 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17069) );
  AOI22_X1 U20301 ( .A1(n17067), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17068) );
  NAND4_X1 U20302 ( .A1(n17071), .A2(n17070), .A3(n17069), .A4(n17068), .ZN(
        n17078) );
  AOI22_X1 U20303 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9618), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17076) );
  AOI22_X1 U20304 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17110), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17075) );
  AOI22_X1 U20305 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17088), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17074) );
  AOI22_X1 U20306 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17072), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17073) );
  NAND4_X1 U20307 ( .A1(n17076), .A2(n17075), .A3(n17074), .A4(n17073), .ZN(
        n17077) );
  NOR2_X1 U20308 ( .A1(n17078), .A2(n17077), .ZN(n17262) );
  OAI21_X1 U20309 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17099), .A(n17079), .ZN(
        n17080) );
  AOI22_X1 U20310 ( .A1(n17146), .A2(n17262), .B1(n17080), .B2(n17141), .ZN(
        P3_U2693) );
  AOI22_X1 U20311 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17081), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17086) );
  AOI22_X1 U20312 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17085) );
  AOI22_X1 U20313 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n9614), .ZN(n17084) );
  AOI22_X1 U20314 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17104), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n17067), .ZN(n17083) );
  NAND4_X1 U20315 ( .A1(n17086), .A2(n17085), .A3(n17084), .A4(n17083), .ZN(
        n17096) );
  AOI22_X1 U20316 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17087), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17094) );
  AOI22_X1 U20317 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17089), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17088), .ZN(n17093) );
  AOI22_X1 U20318 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17090), .ZN(n17092) );
  AOI22_X1 U20319 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9616), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17091) );
  NAND4_X1 U20320 ( .A1(n17094), .A2(n17093), .A3(n17092), .A4(n17091), .ZN(
        n17095) );
  NOR2_X1 U20321 ( .A1(n17096), .A2(n17095), .ZN(n17266) );
  INV_X1 U20322 ( .A(n17121), .ZN(n17097) );
  OAI21_X1 U20323 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17097), .A(n17141), .ZN(
        n17098) );
  OAI22_X1 U20324 ( .A1(n17266), .A2(n17141), .B1(n17099), .B2(n17098), .ZN(
        P3_U2694) );
  AOI22_X1 U20325 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n15741), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17120) );
  AOI22_X1 U20326 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17100), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17119) );
  AOI22_X1 U20327 ( .A1(n17072), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17081), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17102) );
  OAI21_X1 U20328 ( .B1(n17103), .B2(n18104), .A(n17102), .ZN(n17116) );
  AOI22_X1 U20329 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17114) );
  AOI22_X1 U20330 ( .A1(n17107), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17106), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17113) );
  AOI22_X1 U20331 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17112) );
  AOI22_X1 U20332 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17111) );
  NAND4_X1 U20333 ( .A1(n17114), .A2(n17113), .A3(n17112), .A4(n17111), .ZN(
        n17115) );
  AOI211_X1 U20334 ( .C1(n17117), .C2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n17116), .B(n17115), .ZN(n17118) );
  NAND3_X1 U20335 ( .A1(n17120), .A2(n17119), .A3(n17118), .ZN(n17270) );
  INV_X1 U20336 ( .A(n17270), .ZN(n17123) );
  OAI21_X1 U20337 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17125), .A(n17121), .ZN(
        n17122) );
  AOI22_X1 U20338 ( .A1(n17146), .A2(n17123), .B1(n17122), .B2(n17141), .ZN(
        P3_U2695) );
  NOR2_X1 U20339 ( .A1(n17240), .A2(n17126), .ZN(n17127) );
  AOI22_X1 U20340 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17141), .B1(
        P3_EBX_REG_6__SCAN_IN), .B2(n17127), .ZN(n17124) );
  INV_X1 U20341 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18140) );
  OAI22_X1 U20342 ( .A1(n17125), .A2(n17124), .B1(n18140), .B2(n17141), .ZN(
        P3_U2696) );
  INV_X1 U20343 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17129) );
  NAND2_X1 U20344 ( .A1(n17141), .A2(n17126), .ZN(n17130) );
  AOI22_X1 U20345 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n17146), .B1(
        n17127), .B2(n17129), .ZN(n17128) );
  OAI21_X1 U20346 ( .B1(n17129), .B2(n17130), .A(n17128), .ZN(P3_U2697) );
  AOI21_X1 U20347 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17136), .A(
        P3_EBX_REG_5__SCAN_IN), .ZN(n17131) );
  OAI22_X1 U20348 ( .A1(n17131), .A2(n17130), .B1(n20890), .B2(n17141), .ZN(
        P3_U2698) );
  NAND2_X1 U20349 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17136), .ZN(n17132) );
  OAI21_X1 U20350 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17136), .A(n17132), .ZN(
        n17133) );
  AOI22_X1 U20351 ( .A1(n17146), .A2(n18122), .B1(n17133), .B2(n17141), .ZN(
        P3_U2699) );
  NOR2_X1 U20352 ( .A1(n17134), .A2(n17148), .ZN(n17139) );
  AOI21_X1 U20353 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17141), .A(n17139), .ZN(
        n17135) );
  INV_X1 U20354 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18117) );
  OAI22_X1 U20355 ( .A1(n17136), .A2(n17135), .B1(n18117), .B2(n17141), .ZN(
        P3_U2700) );
  INV_X1 U20356 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18112) );
  INV_X1 U20357 ( .A(n17137), .ZN(n17138) );
  AOI221_X1 U20358 ( .B1(n17138), .B2(n17142), .C1(n17240), .C2(n17142), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17140) );
  AOI211_X1 U20359 ( .C1(n17146), .C2(n18112), .A(n17140), .B(n17139), .ZN(
        P3_U2701) );
  OAI222_X1 U20360 ( .A1(n17144), .A2(n17148), .B1(n17143), .B2(n17142), .C1(
        n18107), .C2(n17141), .ZN(P3_U2702) );
  AOI22_X1 U20361 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17146), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17145), .ZN(n17147) );
  OAI21_X1 U20362 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17148), .A(n17147), .ZN(
        P3_U2703) );
  INV_X1 U20363 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17371) );
  INV_X1 U20364 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17367) );
  INV_X1 U20365 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17363) );
  INV_X1 U20366 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17357) );
  INV_X1 U20367 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17411) );
  INV_X1 U20368 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17377) );
  INV_X1 U20369 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17383) );
  NAND4_X1 U20370 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .A3(P3_EAX_REG_2__SCAN_IN), .A4(P3_EAX_REG_5__SCAN_IN), .ZN(n17149) );
  NOR3_X1 U20371 ( .A1(n17377), .A2(n17383), .A3(n17149), .ZN(n17277) );
  NAND2_X1 U20372 ( .A1(n17277), .A2(P3_EAX_REG_7__SCAN_IN), .ZN(n17241) );
  NAND3_X1 U20373 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .A3(P3_EAX_REG_8__SCAN_IN), .ZN(n17242) );
  NAND2_X1 U20374 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .ZN(n17243) );
  NOR2_X1 U20375 ( .A1(n17242), .A2(n17243), .ZN(n17150) );
  NAND4_X1 U20376 ( .A1(n17272), .A2(P3_EAX_REG_14__SCAN_IN), .A3(
        P3_EAX_REG_11__SCAN_IN), .A4(n17150), .ZN(n17236) );
  INV_X1 U20377 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17353) );
  INV_X1 U20378 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17351) );
  NOR2_X1 U20379 ( .A1(n17353), .A2(n17351), .ZN(n17197) );
  NAND4_X1 U20380 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_17__SCAN_IN), .A4(n17197), .ZN(n17203) );
  NAND2_X1 U20381 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17191), .ZN(n17190) );
  NAND2_X1 U20382 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17179), .ZN(n17175) );
  NAND2_X1 U20383 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17174), .ZN(n17165) );
  NAND2_X1 U20384 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17164), .ZN(n17155) );
  NAND3_X1 U20385 ( .A1(n20926), .A2(P3_EAX_REG_31__SCAN_IN), .A3(n17155), 
        .ZN(n17153) );
  NOR2_X2 U20386 ( .A1(n18127), .A2(n17297), .ZN(n17229) );
  NAND2_X1 U20387 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17229), .ZN(n17152) );
  OAI211_X1 U20388 ( .C1(P3_EAX_REG_31__SCAN_IN), .C2(n17155), .A(n17153), .B(
        n17152), .ZN(P3_U2704) );
  NOR2_X2 U20389 ( .A1(n17154), .A2(n17297), .ZN(n17230) );
  AOI22_X1 U20390 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17230), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17229), .ZN(n17157) );
  OAI211_X1 U20391 ( .C1(n17164), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17297), .B(
        n17155), .ZN(n17156) );
  OAI211_X1 U20392 ( .C1(n17158), .C2(n20928), .A(n17157), .B(n17156), .ZN(
        P3_U2705) );
  INV_X1 U20393 ( .A(n17165), .ZN(n17159) );
  AOI21_X1 U20394 ( .B1(P3_EAX_REG_29__SCAN_IN), .B2(n20926), .A(n17159), .ZN(
        n17163) );
  AOI22_X1 U20395 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17230), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17229), .ZN(n17162) );
  NAND2_X1 U20396 ( .A1(n17271), .A2(n17160), .ZN(n17161) );
  OAI211_X1 U20397 ( .C1(n17164), .C2(n17163), .A(n17162), .B(n17161), .ZN(
        P3_U2706) );
  AOI22_X1 U20398 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17230), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17229), .ZN(n17167) );
  OAI211_X1 U20399 ( .C1(n17174), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17297), .B(
        n17165), .ZN(n17166) );
  OAI211_X1 U20400 ( .C1(n17168), .C2(n20928), .A(n17167), .B(n17166), .ZN(
        P3_U2707) );
  INV_X1 U20401 ( .A(n17175), .ZN(n17169) );
  AOI21_X1 U20402 ( .B1(P3_EAX_REG_27__SCAN_IN), .B2(n20926), .A(n17169), .ZN(
        n17173) );
  AOI22_X1 U20403 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17230), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17229), .ZN(n17172) );
  NAND2_X1 U20404 ( .A1(n17271), .A2(n17170), .ZN(n17171) );
  OAI211_X1 U20405 ( .C1(n17174), .C2(n17173), .A(n17172), .B(n17171), .ZN(
        P3_U2708) );
  AOI22_X1 U20406 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17230), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17229), .ZN(n17177) );
  OAI211_X1 U20407 ( .C1(n17179), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17297), .B(
        n17175), .ZN(n17176) );
  OAI211_X1 U20408 ( .C1(n17178), .C2(n20928), .A(n17177), .B(n17176), .ZN(
        P3_U2709) );
  AOI22_X1 U20409 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17230), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17229), .ZN(n17183) );
  INV_X1 U20410 ( .A(n17185), .ZN(n17181) );
  INV_X1 U20411 ( .A(n17179), .ZN(n17180) );
  OAI211_X1 U20412 ( .C1(n17181), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17297), .B(
        n17180), .ZN(n17182) );
  OAI211_X1 U20413 ( .C1(n17184), .C2(n20928), .A(n17183), .B(n17182), .ZN(
        P3_U2710) );
  AOI22_X1 U20414 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17230), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17229), .ZN(n17188) );
  OAI211_X1 U20415 ( .C1(n17186), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17297), .B(
        n17185), .ZN(n17187) );
  OAI211_X1 U20416 ( .C1(n17189), .C2(n20928), .A(n17188), .B(n17187), .ZN(
        P3_U2711) );
  AOI22_X1 U20417 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17230), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17229), .ZN(n17193) );
  OAI211_X1 U20418 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17191), .A(n20926), .B(
        n17190), .ZN(n17192) );
  OAI211_X1 U20419 ( .C1(n17194), .C2(n20928), .A(n17193), .B(n17192), .ZN(
        P3_U2712) );
  NOR2_X1 U20420 ( .A1(n17240), .A2(n17231), .ZN(n17225) );
  NAND2_X1 U20421 ( .A1(n17225), .A2(n17357), .ZN(n17202) );
  AOI22_X1 U20422 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17229), .B1(n17271), .B2(
        n17195), .ZN(n17201) );
  INV_X1 U20423 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17349) );
  INV_X1 U20424 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17347) );
  NOR2_X1 U20425 ( .A1(n17349), .A2(n17347), .ZN(n17196) );
  NAND2_X1 U20426 ( .A1(n17196), .A2(n17225), .ZN(n17219) );
  INV_X1 U20427 ( .A(n17219), .ZN(n17215) );
  NAND2_X1 U20428 ( .A1(n17197), .A2(n17215), .ZN(n17209) );
  NAND2_X1 U20429 ( .A1(n20926), .A2(n17209), .ZN(n17212) );
  OAI21_X1 U20430 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17198), .A(n17212), .ZN(
        n17199) );
  AOI22_X1 U20431 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17230), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17199), .ZN(n17200) );
  OAI211_X1 U20432 ( .C1(n17203), .C2(n17202), .A(n17201), .B(n17200), .ZN(
        P3_U2713) );
  INV_X1 U20433 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17355) );
  INV_X1 U20434 ( .A(n17229), .ZN(n17204) );
  OAI22_X1 U20435 ( .A1(n17205), .A2(n20928), .B1(n15113), .B2(n17204), .ZN(
        n17206) );
  AOI21_X1 U20436 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17230), .A(n17206), .ZN(
        n17207) );
  OAI221_X1 U20437 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17209), .C1(n17355), 
        .C2(n17212), .A(n17207), .ZN(P3_U2714) );
  AOI22_X1 U20438 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17230), .B1(n17271), .B2(
        n17208), .ZN(n17211) );
  NOR2_X1 U20439 ( .A1(n17351), .A2(n17219), .ZN(n17213) );
  AOI22_X1 U20440 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17229), .B1(n17213), .B2(
        n17209), .ZN(n17210) );
  OAI211_X1 U20441 ( .C1(n17353), .C2(n17212), .A(n17211), .B(n17210), .ZN(
        P3_U2715) );
  AOI22_X1 U20442 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17230), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17229), .ZN(n17217) );
  INV_X1 U20443 ( .A(n17213), .ZN(n17214) );
  OAI211_X1 U20444 ( .C1(n17215), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17297), .B(
        n17214), .ZN(n17216) );
  OAI211_X1 U20445 ( .C1(n17218), .C2(n20928), .A(n17217), .B(n17216), .ZN(
        P3_U2716) );
  AOI22_X1 U20446 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17230), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17229), .ZN(n17222) );
  NAND2_X1 U20447 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17225), .ZN(n17224) );
  INV_X1 U20448 ( .A(n17224), .ZN(n17220) );
  OAI211_X1 U20449 ( .C1(n17220), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17297), .B(
        n17219), .ZN(n17221) );
  OAI211_X1 U20450 ( .C1(n17223), .C2(n20928), .A(n17222), .B(n17221), .ZN(
        P3_U2717) );
  AOI22_X1 U20451 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17230), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17229), .ZN(n17227) );
  OAI211_X1 U20452 ( .C1(n17225), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17297), .B(
        n17224), .ZN(n17226) );
  OAI211_X1 U20453 ( .C1(n17228), .C2(n20928), .A(n17227), .B(n17226), .ZN(
        P3_U2718) );
  AOI22_X1 U20454 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17230), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17229), .ZN(n17234) );
  OAI211_X1 U20455 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17232), .A(n20926), .B(
        n17231), .ZN(n17233) );
  OAI211_X1 U20456 ( .C1(n17235), .C2(n20928), .A(n17234), .B(n17233), .ZN(
        P3_U2719) );
  OR2_X1 U20457 ( .A1(n17240), .A2(n17236), .ZN(n17239) );
  NAND2_X1 U20458 ( .A1(n20926), .A2(n17236), .ZN(n17246) );
  AOI22_X1 U20459 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17295), .B1(n17271), .B2(
        n17237), .ZN(n17238) );
  OAI221_X1 U20460 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(n17239), .C1(n17411), 
        .C2(n17246), .A(n17238), .ZN(P3_U2720) );
  INV_X1 U20461 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17397) );
  NOR2_X1 U20462 ( .A1(n17240), .A2(n17296), .ZN(n17294) );
  INV_X1 U20463 ( .A(n17294), .ZN(n17281) );
  INV_X1 U20464 ( .A(n17279), .ZN(n17261) );
  NOR2_X1 U20465 ( .A1(n17397), .A2(n17260), .ZN(n17253) );
  INV_X1 U20466 ( .A(n17253), .ZN(n17248) );
  NOR2_X1 U20467 ( .A1(n17243), .A2(n17248), .ZN(n17250) );
  INV_X1 U20468 ( .A(n17250), .ZN(n17247) );
  INV_X1 U20469 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17406) );
  AOI22_X1 U20470 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17295), .B1(n17271), .B2(
        n17244), .ZN(n17245) );
  OAI221_X1 U20471 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n17247), .C1(n17406), 
        .C2(n17246), .A(n17245), .ZN(P3_U2721) );
  INV_X1 U20472 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17400) );
  NOR2_X1 U20473 ( .A1(n17400), .A2(n17248), .ZN(n17256) );
  AOI21_X1 U20474 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n20926), .A(n17256), .ZN(
        n17251) );
  OAI222_X1 U20475 ( .A1(n20931), .A2(n17252), .B1(n17251), .B2(n17250), .C1(
        n20928), .C2(n17249), .ZN(P3_U2722) );
  AOI21_X1 U20476 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n20926), .A(n17253), .ZN(
        n17255) );
  OAI222_X1 U20477 ( .A1(n20931), .A2(n17257), .B1(n17256), .B2(n17255), .C1(
        n20928), .C2(n17254), .ZN(P3_U2723) );
  NAND2_X1 U20478 ( .A1(n20926), .A2(n17260), .ZN(n17264) );
  AOI22_X1 U20479 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17295), .B1(n17271), .B2(
        n17258), .ZN(n17259) );
  OAI221_X1 U20480 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17260), .C1(n17397), 
        .C2(n17264), .A(n17259), .ZN(P3_U2724) );
  INV_X1 U20481 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17393) );
  INV_X1 U20482 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17391) );
  NOR3_X1 U20483 ( .A1(n17393), .A2(n17391), .A3(n17261), .ZN(n17268) );
  NOR2_X1 U20484 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17268), .ZN(n17263) );
  OAI222_X1 U20485 ( .A1(n20931), .A2(n17265), .B1(n17264), .B2(n17263), .C1(
        n20928), .C2(n17262), .ZN(P3_U2725) );
  AOI22_X1 U20486 ( .A1(n17279), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n17297), .ZN(n17267) );
  OAI222_X1 U20487 ( .A1(n20931), .A2(n17269), .B1(n17268), .B2(n17267), .C1(
        n20928), .C2(n17266), .ZN(P3_U2726) );
  AOI22_X1 U20488 ( .A1(n17271), .A2(n17270), .B1(n17279), .B2(n17391), .ZN(
        n17275) );
  INV_X1 U20489 ( .A(n17272), .ZN(n17273) );
  NAND3_X1 U20490 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n20926), .A3(n17273), .ZN(
        n17274) );
  OAI211_X1 U20491 ( .C1(n20931), .C2(n17276), .A(n17275), .B(n17274), .ZN(
        P3_U2727) );
  AND2_X1 U20492 ( .A1(n17277), .A2(n17294), .ZN(n20930) );
  AOI21_X1 U20493 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n20926), .A(n20930), .ZN(
        n17280) );
  OAI222_X1 U20494 ( .A1(n20931), .A2(n18131), .B1(n17280), .B2(n17279), .C1(
        n20928), .C2(n17278), .ZN(P3_U2728) );
  INV_X1 U20495 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17385) );
  INV_X1 U20496 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17379) );
  NOR3_X1 U20497 ( .A1(n17377), .A2(n17379), .A3(n17281), .ZN(n17293) );
  AND2_X1 U20498 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17293), .ZN(n17290) );
  NAND2_X1 U20499 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17290), .ZN(n17282) );
  NOR2_X1 U20500 ( .A1(n17385), .A2(n17282), .ZN(n20925) );
  INV_X1 U20501 ( .A(n17282), .ZN(n17287) );
  AOI21_X1 U20502 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n20926), .A(n17287), .ZN(
        n17284) );
  OAI222_X1 U20503 ( .A1(n18123), .A2(n20931), .B1(n20925), .B2(n17284), .C1(
        n20928), .C2(n17283), .ZN(P3_U2730) );
  AOI21_X1 U20504 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n20926), .A(n17290), .ZN(
        n17286) );
  OAI222_X1 U20505 ( .A1(n18118), .A2(n20931), .B1(n17287), .B2(n17286), .C1(
        n20928), .C2(n17285), .ZN(P3_U2731) );
  AOI21_X1 U20506 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n20926), .A(n17293), .ZN(
        n17289) );
  OAI222_X1 U20507 ( .A1(n18113), .A2(n20931), .B1(n17290), .B2(n17289), .C1(
        n20928), .C2(n17288), .ZN(P3_U2732) );
  AOI22_X1 U20508 ( .A1(n17294), .A2(P3_EAX_REG_1__SCAN_IN), .B1(
        P3_EAX_REG_2__SCAN_IN), .B2(n17297), .ZN(n17292) );
  OAI222_X1 U20509 ( .A1(n18108), .A2(n20931), .B1(n17293), .B2(n17292), .C1(
        n20928), .C2(n17291), .ZN(P3_U2733) );
  AOI22_X1 U20510 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17295), .B1(n17294), .B2(
        n17377), .ZN(n17299) );
  NAND3_X1 U20511 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17297), .A3(n17296), .ZN(
        n17298) );
  OAI211_X1 U20512 ( .C1(n17300), .C2(n20928), .A(n17299), .B(n17298), .ZN(
        P3_U2734) );
  INV_X1 U20513 ( .A(n17610), .ZN(n18613) );
  INV_X1 U20514 ( .A(n17301), .ZN(n17343) );
  AND2_X1 U20515 ( .A1(n17317), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20516 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17373) );
  INV_X1 U20517 ( .A(n18748), .ZN(n17305) );
  NAND3_X1 U20518 ( .A1(n17306), .A2(n17305), .A3(n17304), .ZN(n17323) );
  AOI22_X1 U20519 ( .A1(n18747), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17317), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17307) );
  OAI21_X1 U20520 ( .B1(n17373), .B2(n17323), .A(n17307), .ZN(P3_U2737) );
  AOI22_X1 U20521 ( .A1(n18747), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17317), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17308) );
  OAI21_X1 U20522 ( .B1(n17371), .B2(n17323), .A(n17308), .ZN(P3_U2738) );
  INV_X1 U20523 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17369) );
  AOI22_X1 U20524 ( .A1(n18747), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17317), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17309) );
  OAI21_X1 U20525 ( .B1(n17369), .B2(n17323), .A(n17309), .ZN(P3_U2739) );
  AOI22_X1 U20526 ( .A1(n18747), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17310) );
  OAI21_X1 U20527 ( .B1(n17367), .B2(n17323), .A(n17310), .ZN(P3_U2740) );
  INV_X1 U20528 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17365) );
  AOI22_X1 U20529 ( .A1(n18747), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17317), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17311) );
  OAI21_X1 U20530 ( .B1(n17365), .B2(n17323), .A(n17311), .ZN(P3_U2741) );
  AOI22_X1 U20531 ( .A1(n18747), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17317), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17312) );
  OAI21_X1 U20532 ( .B1(n17363), .B2(n17323), .A(n17312), .ZN(P3_U2742) );
  INV_X1 U20533 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17361) );
  AOI22_X1 U20534 ( .A1(n18747), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17317), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17313) );
  OAI21_X1 U20535 ( .B1(n17361), .B2(n17323), .A(n17313), .ZN(P3_U2743) );
  INV_X1 U20536 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17359) );
  AOI22_X1 U20537 ( .A1(n17340), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17317), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17314) );
  OAI21_X1 U20538 ( .B1(n17359), .B2(n17323), .A(n17314), .ZN(P3_U2744) );
  AOI22_X1 U20539 ( .A1(n17340), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17317), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17315) );
  OAI21_X1 U20540 ( .B1(n17357), .B2(n17323), .A(n17315), .ZN(P3_U2745) );
  AOI22_X1 U20541 ( .A1(n17340), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17317), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17316) );
  OAI21_X1 U20542 ( .B1(n17355), .B2(n17323), .A(n17316), .ZN(P3_U2746) );
  AOI22_X1 U20543 ( .A1(n17340), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17317), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17318) );
  OAI21_X1 U20544 ( .B1(n17353), .B2(n17323), .A(n17318), .ZN(P3_U2747) );
  AOI22_X1 U20545 ( .A1(n17340), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(
        P3_DATAO_REG_19__SCAN_IN), .B2(n17339), .ZN(n17319) );
  OAI21_X1 U20546 ( .B1(n17351), .B2(n17323), .A(n17319), .ZN(P3_U2748) );
  AOI22_X1 U20547 ( .A1(n17340), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17320) );
  OAI21_X1 U20548 ( .B1(n17349), .B2(n17323), .A(n17320), .ZN(P3_U2749) );
  AOI22_X1 U20549 ( .A1(n17340), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17321) );
  OAI21_X1 U20550 ( .B1(n17347), .B2(n17323), .A(n17321), .ZN(P3_U2750) );
  INV_X1 U20551 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17345) );
  AOI22_X1 U20552 ( .A1(n17340), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17322) );
  OAI21_X1 U20553 ( .B1(n17345), .B2(n17323), .A(n17322), .ZN(P3_U2751) );
  AOI22_X1 U20554 ( .A1(n17340), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17324) );
  OAI21_X1 U20555 ( .B1(n17411), .B2(n17342), .A(n17324), .ZN(P3_U2752) );
  AOI22_X1 U20556 ( .A1(n17340), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17325) );
  OAI21_X1 U20557 ( .B1(n17406), .B2(n17342), .A(n17325), .ZN(P3_U2753) );
  INV_X1 U20558 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17402) );
  AOI22_X1 U20559 ( .A1(n17340), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17326) );
  OAI21_X1 U20560 ( .B1(n17402), .B2(n17342), .A(n17326), .ZN(P3_U2754) );
  AOI22_X1 U20561 ( .A1(n17340), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17327) );
  OAI21_X1 U20562 ( .B1(n17400), .B2(n17342), .A(n17327), .ZN(P3_U2755) );
  AOI22_X1 U20563 ( .A1(n17340), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17328) );
  OAI21_X1 U20564 ( .B1(n17397), .B2(n17342), .A(n17328), .ZN(P3_U2756) );
  INV_X1 U20565 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17395) );
  AOI22_X1 U20566 ( .A1(n17340), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17329) );
  OAI21_X1 U20567 ( .B1(n17395), .B2(n17342), .A(n17329), .ZN(P3_U2757) );
  AOI22_X1 U20568 ( .A1(n17340), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(
        P3_DATAO_REG_9__SCAN_IN), .B2(n17339), .ZN(n17330) );
  OAI21_X1 U20569 ( .B1(n17393), .B2(n17342), .A(n17330), .ZN(P3_U2758) );
  AOI22_X1 U20570 ( .A1(n17340), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17331) );
  OAI21_X1 U20571 ( .B1(n17391), .B2(n17342), .A(n17331), .ZN(P3_U2759) );
  INV_X1 U20572 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17389) );
  AOI22_X1 U20573 ( .A1(n17340), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17332) );
  OAI21_X1 U20574 ( .B1(n17389), .B2(n17342), .A(n17332), .ZN(P3_U2760) );
  INV_X1 U20575 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17387) );
  AOI22_X1 U20576 ( .A1(n17340), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17333) );
  OAI21_X1 U20577 ( .B1(n17387), .B2(n17342), .A(n17333), .ZN(P3_U2761) );
  AOI22_X1 U20578 ( .A1(n17340), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17334) );
  OAI21_X1 U20579 ( .B1(n17385), .B2(n17342), .A(n17334), .ZN(P3_U2762) );
  AOI22_X1 U20580 ( .A1(n17340), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17335) );
  OAI21_X1 U20581 ( .B1(n17383), .B2(n17342), .A(n17335), .ZN(P3_U2763) );
  INV_X1 U20582 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17381) );
  AOI22_X1 U20583 ( .A1(n17340), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17336) );
  OAI21_X1 U20584 ( .B1(n17381), .B2(n17342), .A(n17336), .ZN(P3_U2764) );
  AOI22_X1 U20585 ( .A1(n17340), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17337) );
  OAI21_X1 U20586 ( .B1(n17379), .B2(n17342), .A(n17337), .ZN(P3_U2765) );
  AOI22_X1 U20587 ( .A1(n17340), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17338) );
  OAI21_X1 U20588 ( .B1(n17377), .B2(n17342), .A(n17338), .ZN(P3_U2766) );
  AOI22_X1 U20589 ( .A1(n17340), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17339), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17341) );
  OAI21_X1 U20590 ( .B1(n17375), .B2(n17342), .A(n17341), .ZN(P3_U2767) );
  NAND3_X1 U20591 ( .A1(n18750), .A2(n18593), .A3(n17343), .ZN(n17410) );
  OAI211_X1 U20592 ( .C1(n18750), .C2(n18751), .A(n18593), .B(n17343), .ZN(
        n17398) );
  AOI22_X1 U20593 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17403), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17407), .ZN(n17344) );
  OAI21_X1 U20594 ( .B1(n17345), .B2(n17405), .A(n17344), .ZN(P3_U2768) );
  AOI22_X1 U20595 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17403), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17407), .ZN(n17346) );
  OAI21_X1 U20596 ( .B1(n17347), .B2(n17405), .A(n17346), .ZN(P3_U2769) );
  AOI22_X1 U20597 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17403), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17407), .ZN(n17348) );
  OAI21_X1 U20598 ( .B1(n17349), .B2(n17405), .A(n17348), .ZN(P3_U2770) );
  AOI22_X1 U20599 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17403), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17407), .ZN(n17350) );
  OAI21_X1 U20600 ( .B1(n17351), .B2(n17405), .A(n17350), .ZN(P3_U2771) );
  AOI22_X1 U20601 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17408), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17407), .ZN(n17352) );
  OAI21_X1 U20602 ( .B1(n17353), .B2(n17405), .A(n17352), .ZN(P3_U2772) );
  AOI22_X1 U20603 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17408), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17407), .ZN(n17354) );
  OAI21_X1 U20604 ( .B1(n17355), .B2(n17405), .A(n17354), .ZN(P3_U2773) );
  AOI22_X1 U20605 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17408), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17407), .ZN(n17356) );
  OAI21_X1 U20606 ( .B1(n17357), .B2(n17405), .A(n17356), .ZN(P3_U2774) );
  AOI22_X1 U20607 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17408), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17407), .ZN(n17358) );
  OAI21_X1 U20608 ( .B1(n17359), .B2(n17405), .A(n17358), .ZN(P3_U2775) );
  AOI22_X1 U20609 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17408), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17407), .ZN(n17360) );
  OAI21_X1 U20610 ( .B1(n17361), .B2(n17405), .A(n17360), .ZN(P3_U2776) );
  AOI22_X1 U20611 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17408), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17407), .ZN(n17362) );
  OAI21_X1 U20612 ( .B1(n17363), .B2(n17405), .A(n17362), .ZN(P3_U2777) );
  AOI22_X1 U20613 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17408), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17407), .ZN(n17364) );
  OAI21_X1 U20614 ( .B1(n17365), .B2(n17405), .A(n17364), .ZN(P3_U2778) );
  AOI22_X1 U20615 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17408), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17407), .ZN(n17366) );
  OAI21_X1 U20616 ( .B1(n17367), .B2(n17405), .A(n17366), .ZN(P3_U2779) );
  AOI22_X1 U20617 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17403), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17407), .ZN(n17368) );
  OAI21_X1 U20618 ( .B1(n17369), .B2(n17410), .A(n17368), .ZN(P3_U2780) );
  AOI22_X1 U20619 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17403), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17407), .ZN(n17370) );
  OAI21_X1 U20620 ( .B1(n17371), .B2(n17410), .A(n17370), .ZN(P3_U2781) );
  AOI22_X1 U20621 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17403), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17407), .ZN(n17372) );
  OAI21_X1 U20622 ( .B1(n17373), .B2(n17410), .A(n17372), .ZN(P3_U2782) );
  AOI22_X1 U20623 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17403), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17407), .ZN(n17374) );
  OAI21_X1 U20624 ( .B1(n17375), .B2(n17410), .A(n17374), .ZN(P3_U2783) );
  AOI22_X1 U20625 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17403), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17407), .ZN(n17376) );
  OAI21_X1 U20626 ( .B1(n17377), .B2(n17410), .A(n17376), .ZN(P3_U2784) );
  AOI22_X1 U20627 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17403), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17407), .ZN(n17378) );
  OAI21_X1 U20628 ( .B1(n17379), .B2(n17410), .A(n17378), .ZN(P3_U2785) );
  AOI22_X1 U20629 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17403), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17398), .ZN(n17380) );
  OAI21_X1 U20630 ( .B1(n17381), .B2(n17410), .A(n17380), .ZN(P3_U2786) );
  AOI22_X1 U20631 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17403), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17398), .ZN(n17382) );
  OAI21_X1 U20632 ( .B1(n17383), .B2(n17410), .A(n17382), .ZN(P3_U2787) );
  AOI22_X1 U20633 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17403), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17398), .ZN(n17384) );
  OAI21_X1 U20634 ( .B1(n17385), .B2(n17410), .A(n17384), .ZN(P3_U2788) );
  AOI22_X1 U20635 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17403), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17398), .ZN(n17386) );
  OAI21_X1 U20636 ( .B1(n17387), .B2(n17410), .A(n17386), .ZN(P3_U2789) );
  AOI22_X1 U20637 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17403), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17398), .ZN(n17388) );
  OAI21_X1 U20638 ( .B1(n17389), .B2(n17410), .A(n17388), .ZN(P3_U2790) );
  AOI22_X1 U20639 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17403), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17398), .ZN(n17390) );
  OAI21_X1 U20640 ( .B1(n17391), .B2(n17405), .A(n17390), .ZN(P3_U2791) );
  AOI22_X1 U20641 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17403), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17398), .ZN(n17392) );
  OAI21_X1 U20642 ( .B1(n17393), .B2(n17410), .A(n17392), .ZN(P3_U2792) );
  AOI22_X1 U20643 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17408), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17398), .ZN(n17394) );
  OAI21_X1 U20644 ( .B1(n17395), .B2(n17410), .A(n17394), .ZN(P3_U2793) );
  AOI22_X1 U20645 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17403), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17398), .ZN(n17396) );
  OAI21_X1 U20646 ( .B1(n17397), .B2(n17410), .A(n17396), .ZN(P3_U2794) );
  AOI22_X1 U20647 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17403), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17398), .ZN(n17399) );
  OAI21_X1 U20648 ( .B1(n17400), .B2(n17410), .A(n17399), .ZN(P3_U2795) );
  AOI22_X1 U20649 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17408), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17407), .ZN(n17401) );
  OAI21_X1 U20650 ( .B1(n17402), .B2(n17410), .A(n17401), .ZN(P3_U2796) );
  AOI22_X1 U20651 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17403), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17407), .ZN(n17404) );
  OAI21_X1 U20652 ( .B1(n17406), .B2(n17405), .A(n17404), .ZN(P3_U2797) );
  AOI22_X1 U20653 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17408), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17407), .ZN(n17409) );
  OAI21_X1 U20654 ( .B1(n17411), .B2(n17410), .A(n17409), .ZN(P3_U2798) );
  INV_X1 U20655 ( .A(n17436), .ZN(n17427) );
  OAI21_X1 U20656 ( .B1(n17412), .B2(n18613), .A(n17764), .ZN(n17413) );
  AOI21_X1 U20657 ( .B1(n17726), .B2(n17417), .A(n17413), .ZN(n17442) );
  OAI21_X1 U20658 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17490), .A(
        n17442), .ZN(n17433) );
  AOI211_X1 U20659 ( .C1(n17416), .C2(n17415), .A(n17414), .B(n17678), .ZN(
        n17423) );
  NAND2_X1 U20660 ( .A1(n17985), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17420) );
  NOR2_X1 U20661 ( .A1(n17613), .A2(n17417), .ZN(n17434) );
  OAI211_X1 U20662 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17434), .B(n17418), .ZN(n17419) );
  OAI211_X1 U20663 ( .C1(n17622), .C2(n17421), .A(n17420), .B(n17419), .ZN(
        n17422) );
  AOI211_X1 U20664 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17433), .A(
        n17423), .B(n17422), .ZN(n17426) );
  NAND2_X1 U20665 ( .A1(n17768), .A2(n12354), .ZN(n17521) );
  AOI22_X1 U20666 ( .A1(n17755), .A2(n17780), .B1(n17603), .B2(n17424), .ZN(
        n17444) );
  NAND2_X1 U20667 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17444), .ZN(
        n17435) );
  NAND3_X1 U20668 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17521), .A3(
        n17435), .ZN(n17425) );
  OAI211_X1 U20669 ( .C1(n17428), .C2(n17427), .A(n17426), .B(n17425), .ZN(
        P3_U2802) );
  AOI21_X1 U20670 ( .B1(n17677), .B2(n17429), .A(n9666), .ZN(n17785) );
  INV_X1 U20671 ( .A(n17430), .ZN(n17431) );
  OAI22_X1 U20672 ( .A1(n18069), .A2(n20825), .B1(n17622), .B2(n17431), .ZN(
        n17432) );
  AOI221_X1 U20673 ( .B1(n17434), .B2(n20847), .C1(n17433), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17432), .ZN(n17438) );
  OAI21_X1 U20674 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17436), .A(
        n17435), .ZN(n17437) );
  OAI211_X1 U20675 ( .C1(n17785), .C2(n17678), .A(n17438), .B(n17437), .ZN(
        P3_U2803) );
  AOI21_X1 U20676 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17440), .A(
        n17439), .ZN(n17792) );
  NOR2_X1 U20677 ( .A1(n17532), .A2(n12345), .ZN(n17518) );
  AOI21_X1 U20678 ( .B1(n9719), .B2(n18478), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17441) );
  OAI22_X1 U20679 ( .A1(n17518), .A2(n17443), .B1(n17442), .B2(n17441), .ZN(
        n17446) );
  INV_X1 U20680 ( .A(n17444), .ZN(n17445) );
  INV_X1 U20681 ( .A(n17764), .ZN(n17724) );
  AND2_X1 U20682 ( .A1(n17455), .A2(n18478), .ZN(n17484) );
  AOI211_X1 U20683 ( .C1(n17610), .C2(n17447), .A(n17724), .B(n17484), .ZN(
        n17476) );
  OAI21_X1 U20684 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17490), .A(
        n17476), .ZN(n17461) );
  AOI22_X1 U20685 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17461), .B1(
        n17532), .B2(n17448), .ZN(n17459) );
  XNOR2_X1 U20686 ( .A(n17449), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17803) );
  XNOR2_X1 U20687 ( .A(n17450), .B(n17797), .ZN(n17805) );
  OAI21_X1 U20688 ( .B1(n17677), .B2(n17452), .A(n17451), .ZN(n17453) );
  XNOR2_X1 U20689 ( .A(n17453), .B(n17797), .ZN(n17801) );
  OAI22_X1 U20690 ( .A1(n17768), .A2(n17805), .B1(n17678), .B2(n17801), .ZN(
        n17454) );
  AOI21_X1 U20691 ( .B1(n17603), .B2(n17803), .A(n17454), .ZN(n17458) );
  NAND2_X1 U20692 ( .A1(n17985), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17799) );
  NOR2_X1 U20693 ( .A1(n17613), .A2(n17455), .ZN(n17463) );
  OAI211_X1 U20694 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17463), .B(n17456), .ZN(n17457) );
  NAND4_X1 U20695 ( .A1(n17459), .A2(n17458), .A3(n17799), .A4(n17457), .ZN(
        P3_U2805) );
  INV_X1 U20696 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18677) );
  NOR2_X1 U20697 ( .A1(n18069), .A2(n18677), .ZN(n17460) );
  AOI221_X1 U20698 ( .B1(n17463), .B2(n17462), .C1(n17461), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17460), .ZN(n17471) );
  INV_X1 U20699 ( .A(n17481), .ZN(n17469) );
  NOR2_X1 U20700 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17818), .ZN(
        n17806) );
  INV_X1 U20701 ( .A(n17811), .ZN(n17464) );
  AOI22_X1 U20702 ( .A1(n17755), .A2(n17464), .B1(n17603), .B2(n17808), .ZN(
        n17487) );
  AOI21_X1 U20703 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17466), .A(
        n17465), .ZN(n17817) );
  OAI22_X1 U20704 ( .A1(n17487), .A2(n17467), .B1(n17817), .B2(n17678), .ZN(
        n17468) );
  AOI21_X1 U20705 ( .B1(n17469), .B2(n17806), .A(n17468), .ZN(n17470) );
  OAI211_X1 U20706 ( .C1(n17622), .C2(n17472), .A(n17471), .B(n17470), .ZN(
        P3_U2806) );
  NAND2_X1 U20707 ( .A1(n17985), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17475) );
  OAI21_X1 U20708 ( .B1(n17532), .B2(n12345), .A(n17473), .ZN(n17474) );
  OAI211_X1 U20709 ( .C1(n17476), .C2(n9806), .A(n17475), .B(n17474), .ZN(
        n17483) );
  AOI22_X1 U20710 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17677), .B1(
        n17478), .B2(n17494), .ZN(n17479) );
  NAND2_X1 U20711 ( .A1(n17477), .A2(n17479), .ZN(n17480) );
  XNOR2_X1 U20712 ( .A(n17480), .B(n17818), .ZN(n17823) );
  OAI22_X1 U20713 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17481), .B1(
        n17823), .B2(n17678), .ZN(n17482) );
  AOI211_X1 U20714 ( .C1(n17485), .C2(n17484), .A(n17483), .B(n17482), .ZN(
        n17486) );
  OAI21_X1 U20715 ( .B1(n17487), .B2(n17818), .A(n17486), .ZN(P3_U2807) );
  OAI21_X1 U20716 ( .B1(n17488), .B2(n18613), .A(n17764), .ZN(n17489) );
  AOI21_X1 U20717 ( .B1(n17726), .B2(n17498), .A(n17489), .ZN(n17527) );
  OAI21_X1 U20718 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17490), .A(
        n17527), .ZN(n17504) );
  AOI22_X1 U20719 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17504), .B1(
        n17532), .B2(n17491), .ZN(n17502) );
  NAND2_X1 U20720 ( .A1(n17755), .A2(n17891), .ZN(n17589) );
  OAI21_X1 U20721 ( .B1(n17824), .B2(n12354), .A(n17589), .ZN(n17550) );
  AOI21_X1 U20722 ( .B1(n17827), .B2(n17521), .A(n17550), .ZN(n17512) );
  INV_X1 U20723 ( .A(n17492), .ZN(n17565) );
  AOI221_X1 U20724 ( .B1(n17565), .B2(n17494), .C1(n17827), .C2(n17494), .A(
        n17493), .ZN(n17495) );
  XNOR2_X1 U20725 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17495), .ZN(
        n17838) );
  OAI22_X1 U20726 ( .A1(n17512), .A2(n17833), .B1(n17678), .B2(n17838), .ZN(
        n17496) );
  AOI21_X1 U20727 ( .B1(n17497), .B2(n17833), .A(n17496), .ZN(n17501) );
  NAND2_X1 U20728 ( .A1(n17985), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17836) );
  NOR2_X1 U20729 ( .A1(n17613), .A2(n17498), .ZN(n17506) );
  OAI211_X1 U20730 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17506), .B(n17499), .ZN(n17500) );
  NAND4_X1 U20731 ( .A1(n17502), .A2(n17501), .A3(n17836), .A4(n17500), .ZN(
        P3_U2808) );
  NOR2_X1 U20732 ( .A1(n18069), .A2(n18673), .ZN(n17503) );
  AOI221_X1 U20733 ( .B1(n17506), .B2(n17505), .C1(n17504), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17503), .ZN(n17515) );
  INV_X1 U20734 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n20862) );
  NOR3_X1 U20735 ( .A1(n20862), .A2(n17677), .A3(n17507), .ZN(n17528) );
  INV_X1 U20736 ( .A(n17508), .ZN(n17544) );
  AOI22_X1 U20737 ( .A1(n17844), .A2(n17528), .B1(n17544), .B2(n17509), .ZN(
        n17510) );
  XNOR2_X1 U20738 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17510), .ZN(
        n17840) );
  NAND2_X1 U20739 ( .A1(n17844), .A2(n17511), .ZN(n17848) );
  NAND2_X1 U20740 ( .A1(n17551), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17842) );
  OAI22_X1 U20741 ( .A1(n17512), .A2(n17511), .B1(n17848), .B2(n17541), .ZN(
        n17513) );
  AOI21_X1 U20742 ( .B1(n17666), .B2(n17840), .A(n17513), .ZN(n17514) );
  OAI211_X1 U20743 ( .C1(n17622), .C2(n17516), .A(n17515), .B(n17514), .ZN(
        P3_U2809) );
  AOI21_X1 U20744 ( .B1(n17517), .B2(n18478), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17526) );
  AOI22_X1 U20745 ( .A1(n9612), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n17519), 
        .B2(n17738), .ZN(n17525) );
  OAI221_X1 U20746 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17542), 
        .C1(n17540), .C2(n17528), .A(n17477), .ZN(n17520) );
  XNOR2_X1 U20747 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17520), .ZN(
        n17849) );
  NAND3_X1 U20748 ( .A1(n17551), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17851) );
  AOI21_X1 U20749 ( .B1(n17521), .B2(n17851), .A(n17550), .ZN(n17539) );
  NAND2_X1 U20750 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17522), .ZN(
        n17857) );
  OAI22_X1 U20751 ( .A1(n17539), .A2(n17522), .B1(n17857), .B2(n17541), .ZN(
        n17523) );
  AOI21_X1 U20752 ( .B1(n17666), .B2(n17849), .A(n17523), .ZN(n17524) );
  OAI211_X1 U20753 ( .C1(n17527), .C2(n17526), .A(n17525), .B(n17524), .ZN(
        P3_U2810) );
  AOI21_X1 U20754 ( .B1(n17542), .B2(n17544), .A(n17528), .ZN(n17529) );
  XNOR2_X1 U20755 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n17529), .ZN(
        n17858) );
  AOI21_X1 U20756 ( .B1(n17726), .B2(n17533), .A(n17724), .ZN(n17555) );
  OAI21_X1 U20757 ( .B1(n17530), .B2(n18613), .A(n17555), .ZN(n17547) );
  AOI22_X1 U20758 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17547), .B1(
        n17532), .B2(n17531), .ZN(n17536) );
  NAND2_X1 U20759 ( .A1(n17985), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17860) );
  NOR2_X1 U20760 ( .A1(n17613), .A2(n17533), .ZN(n17549) );
  OAI211_X1 U20761 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17549), .B(n17534), .ZN(n17535) );
  NAND3_X1 U20762 ( .A1(n17536), .A2(n17860), .A3(n17535), .ZN(n17537) );
  AOI21_X1 U20763 ( .B1(n17666), .B2(n17858), .A(n17537), .ZN(n17538) );
  OAI221_X1 U20764 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17541), 
        .C1(n17540), .C2(n17539), .A(n17538), .ZN(P3_U2811) );
  AOI21_X1 U20765 ( .B1(n17564), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17542), .ZN(n17543) );
  XNOR2_X1 U20766 ( .A(n17544), .B(n17543), .ZN(n17872) );
  NAND2_X1 U20767 ( .A1(n17985), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n17870) );
  OAI21_X1 U20768 ( .B1(n17622), .B2(n17545), .A(n17870), .ZN(n17546) );
  AOI221_X1 U20769 ( .B1(n17549), .B2(n17548), .C1(n17547), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17546), .ZN(n17554) );
  INV_X1 U20770 ( .A(n17550), .ZN(n17575) );
  OAI21_X1 U20771 ( .B1(n17551), .B2(n17576), .A(n17575), .ZN(n17561) );
  NOR2_X1 U20772 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17552), .ZN(
        n17868) );
  AOI22_X1 U20773 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17561), .B1(
        n17868), .B2(n17642), .ZN(n17553) );
  OAI211_X1 U20774 ( .C1(n17678), .C2(n17872), .A(n17554), .B(n17553), .ZN(
        P3_U2812) );
  NAND2_X1 U20775 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n20867), .ZN(
        n17879) );
  AOI21_X1 U20776 ( .B1(n9724), .B2(n18478), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17556) );
  NAND2_X1 U20777 ( .A1(n17985), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n17877) );
  OAI21_X1 U20778 ( .B1(n17556), .B2(n17555), .A(n17877), .ZN(n17557) );
  AOI21_X1 U20779 ( .B1(n17558), .B2(n17738), .A(n17557), .ZN(n17563) );
  OAI21_X1 U20780 ( .B1(n17560), .B2(n20867), .A(n17559), .ZN(n17876) );
  AOI22_X1 U20781 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17561), .B1(
        n17666), .B2(n17876), .ZN(n17562) );
  OAI211_X1 U20782 ( .C1(n17576), .C2(n17879), .A(n17563), .B(n17562), .ZN(
        P3_U2813) );
  NAND2_X1 U20783 ( .A1(n17564), .A2(n17644), .ZN(n17664) );
  INV_X1 U20784 ( .A(n17664), .ZN(n17633) );
  AOI22_X1 U20785 ( .A1(n17677), .A2(n17565), .B1(n17633), .B2(n17873), .ZN(
        n17566) );
  XNOR2_X1 U20786 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17566), .ZN(
        n17885) );
  AOI21_X1 U20787 ( .B1(n17726), .B2(n17568), .A(n17724), .ZN(n17595) );
  OAI21_X1 U20788 ( .B1(n17567), .B2(n18613), .A(n17595), .ZN(n17579) );
  AOI22_X1 U20789 ( .A1(n9612), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17579), .ZN(n17571) );
  NOR2_X1 U20790 ( .A1(n17613), .A2(n17568), .ZN(n17581) );
  OAI211_X1 U20791 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17581), .B(n17569), .ZN(n17570) );
  OAI211_X1 U20792 ( .C1(n17622), .C2(n17572), .A(n17571), .B(n17570), .ZN(
        n17573) );
  AOI21_X1 U20793 ( .B1(n17666), .B2(n17885), .A(n17573), .ZN(n17574) );
  OAI221_X1 U20794 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17576), 
        .C1(n20793), .C2(n17575), .A(n17574), .ZN(P3_U2814) );
  NOR2_X1 U20795 ( .A1(n17598), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17890) );
  INV_X1 U20796 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17580) );
  NAND2_X1 U20797 ( .A1(n17985), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n17899) );
  OAI21_X1 U20798 ( .B1(n17622), .B2(n17577), .A(n17899), .ZN(n17578) );
  AOI221_X1 U20799 ( .B1(n17581), .B2(n17580), .C1(n17579), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17578), .ZN(n17588) );
  NOR3_X1 U20800 ( .A1(n17602), .A2(n17936), .A3(n17909), .ZN(n17582) );
  AOI21_X1 U20801 ( .B1(n17607), .B2(n17582), .A(n17590), .ZN(n17583) );
  AOI221_X1 U20802 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17939), 
        .C1(n17677), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17583), .ZN(
        n17584) );
  XNOR2_X1 U20803 ( .A(n17584), .B(n10835), .ZN(n17898) );
  NOR2_X1 U20804 ( .A1(n17824), .A2(n12354), .ZN(n17586) );
  NAND2_X1 U20805 ( .A1(n10835), .A2(n17585), .ZN(n17895) );
  AOI22_X1 U20806 ( .A1(n17666), .A2(n17898), .B1(n17586), .B2(n17895), .ZN(
        n17587) );
  OAI211_X1 U20807 ( .C1(n17890), .C2(n17589), .A(n17588), .B(n17587), .ZN(
        P3_U2815) );
  AOI22_X1 U20808 ( .A1(n17633), .A2(n17907), .B1(n17590), .B2(n17939), .ZN(
        n17591) );
  XNOR2_X1 U20809 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17591), .ZN(
        n17917) );
  INV_X1 U20810 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18658) );
  NOR2_X1 U20811 ( .A1(n18069), .A2(n18658), .ZN(n17597) );
  AOI21_X1 U20812 ( .B1(n17592), .B2(n18478), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17594) );
  OAI22_X1 U20813 ( .A1(n17595), .A2(n17594), .B1(n17518), .B2(n17593), .ZN(
        n17596) );
  AOI211_X1 U20814 ( .C1(n17666), .C2(n17917), .A(n17597), .B(n17596), .ZN(
        n17605) );
  AOI21_X1 U20815 ( .B1(n17602), .B2(n17599), .A(n17598), .ZN(n17914) );
  AOI21_X1 U20816 ( .B1(n17602), .B2(n17601), .A(n17600), .ZN(n17915) );
  AOI22_X1 U20817 ( .A1(n17755), .A2(n17914), .B1(n17603), .B2(n17915), .ZN(
        n17604) );
  NAND2_X1 U20818 ( .A1(n17605), .A2(n17604), .ZN(P3_U2816) );
  AOI22_X1 U20819 ( .A1(n17607), .A2(n17942), .B1(n17939), .B2(n17677), .ZN(
        n17608) );
  AOI21_X1 U20820 ( .B1(n17677), .B2(n17606), .A(n17608), .ZN(n17609) );
  XNOR2_X1 U20821 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17609), .ZN(
        n17935) );
  AOI21_X1 U20822 ( .B1(n17726), .B2(n17636), .A(n17610), .ZN(n17611) );
  OAI21_X1 U20823 ( .B1(n17612), .B2(n17611), .A(n17764), .ZN(n17624) );
  NOR2_X1 U20824 ( .A1(n17613), .A2(n17636), .ZN(n17626) );
  OAI211_X1 U20825 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17626), .B(n17614), .ZN(n17615) );
  NAND2_X1 U20826 ( .A1(n17985), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17933) );
  OAI211_X1 U20827 ( .C1(n17622), .C2(n17616), .A(n17615), .B(n17933), .ZN(
        n17617) );
  AOI21_X1 U20828 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17624), .A(
        n17617), .ZN(n17620) );
  OAI22_X1 U20829 ( .A1(n17928), .A2(n17768), .B1(n17618), .B2(n12354), .ZN(
        n17628) );
  NOR2_X1 U20830 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17905), .ZN(
        n17931) );
  AOI22_X1 U20831 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17628), .B1(
        n17931), .B2(n17642), .ZN(n17619) );
  OAI211_X1 U20832 ( .C1(n17678), .C2(n17935), .A(n17620), .B(n17619), .ZN(
        P3_U2817) );
  NAND2_X1 U20833 ( .A1(n17985), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n17947) );
  OAI21_X1 U20834 ( .B1(n17622), .B2(n17621), .A(n17947), .ZN(n17623) );
  AOI221_X1 U20835 ( .B1(n17626), .B2(n17625), .C1(n17624), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n17623), .ZN(n17631) );
  OAI21_X1 U20836 ( .B1(n17936), .B2(n17664), .A(n17606), .ZN(n17627) );
  XNOR2_X1 U20837 ( .A(n17627), .B(n17939), .ZN(n17946) );
  AOI22_X1 U20838 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17628), .B1(
        n17666), .B2(n17946), .ZN(n17630) );
  INV_X1 U20839 ( .A(n17642), .ZN(n17670) );
  OR3_X1 U20840 ( .A1(n17936), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n17670), .ZN(n17629) );
  NAND3_X1 U20841 ( .A1(n17631), .A2(n17630), .A3(n17629), .ZN(P3_U2818) );
  AOI21_X1 U20842 ( .B1(n17633), .B2(n17922), .A(n17632), .ZN(n17635) );
  XNOR2_X1 U20843 ( .A(n17635), .B(n17634), .ZN(n17963) );
  NOR2_X1 U20844 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17958), .ZN(
        n17950) );
  INV_X1 U20845 ( .A(n17636), .ZN(n17638) );
  INV_X1 U20846 ( .A(n17672), .ZN(n17685) );
  NOR3_X1 U20847 ( .A1(n17685), .A2(n17680), .A3(n18134), .ZN(n17661) );
  NAND3_X1 U20848 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A3(n17661), .ZN(n17650) );
  NAND2_X1 U20849 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n17758), .ZN(
        n17637) );
  AOI22_X1 U20850 ( .A1(n17638), .A2(n18478), .B1(n17650), .B2(n17637), .ZN(
        n17641) );
  INV_X1 U20851 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18652) );
  OAI22_X1 U20852 ( .A1(n17518), .A2(n17639), .B1(n18069), .B2(n18652), .ZN(
        n17640) );
  AOI211_X1 U20853 ( .C1(n17950), .C2(n17642), .A(n17641), .B(n17640), .ZN(
        n17646) );
  NOR2_X1 U20854 ( .A1(n17922), .A2(n17670), .ZN(n17656) );
  OAI22_X1 U20855 ( .A1(n17644), .A2(n12354), .B1(n17768), .B2(n17643), .ZN(
        n17667) );
  OAI21_X1 U20856 ( .B1(n17656), .B2(n17667), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17645) );
  OAI211_X1 U20857 ( .C1(n17963), .C2(n17678), .A(n17646), .B(n17645), .ZN(
        P3_U2819) );
  OAI221_X1 U20858 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17647), .C1(
        n10834), .C2(n17664), .A(n10833), .ZN(n17649) );
  NAND4_X1 U20859 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n10832), .A3(
        n10834), .A4(n17677), .ZN(n17648) );
  OAI211_X1 U20860 ( .C1(n17664), .C2(n17958), .A(n17649), .B(n17648), .ZN(
        n17973) );
  INV_X1 U20861 ( .A(n17650), .ZN(n17652) );
  AOI22_X1 U20862 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17661), .B1(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17758), .ZN(n17651) );
  NAND2_X1 U20863 ( .A1(n17985), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n17971) );
  OAI21_X1 U20864 ( .B1(n17652), .B2(n17651), .A(n17971), .ZN(n17653) );
  AOI21_X1 U20865 ( .B1(n17654), .B2(n17738), .A(n17653), .ZN(n17658) );
  AOI22_X1 U20866 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17667), .B1(
        n17656), .B2(n17655), .ZN(n17657) );
  OAI211_X1 U20867 ( .C1(n17678), .C2(n17973), .A(n17658), .B(n17657), .ZN(
        P3_U2820) );
  NOR2_X1 U20868 ( .A1(n17662), .A2(n17661), .ZN(n17663) );
  OAI22_X1 U20869 ( .A1(n17518), .A2(n17659), .B1(n18069), .B2(n18648), .ZN(
        n17660) );
  AOI221_X1 U20870 ( .B1(n17758), .B2(n17663), .C1(n17662), .C2(n17661), .A(
        n17660), .ZN(n17669) );
  NAND2_X1 U20871 ( .A1(n17664), .A2(n17647), .ZN(n17665) );
  XNOR2_X1 U20872 ( .A(n17665), .B(n10834), .ZN(n17981) );
  AOI22_X1 U20873 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17667), .B1(
        n17666), .B2(n17981), .ZN(n17668) );
  OAI211_X1 U20874 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n17670), .A(
        n17669), .B(n17668), .ZN(P3_U2821) );
  OAI21_X1 U20875 ( .B1(n17672), .B2(n17671), .A(n17764), .ZN(n17686) );
  AOI22_X1 U20876 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17686), .B1(
        n17673), .B2(n17738), .ZN(n17684) );
  AOI21_X1 U20877 ( .B1(n17675), .B2(n18004), .A(n17674), .ZN(n17996) );
  AOI21_X1 U20878 ( .B1(n17677), .B2(n17994), .A(n17676), .ZN(n17999) );
  OAI22_X1 U20879 ( .A1(n17999), .A2(n17678), .B1(n12354), .B2(n17994), .ZN(
        n17679) );
  AOI21_X1 U20880 ( .B1(n17755), .B2(n17996), .A(n17679), .ZN(n17683) );
  NAND2_X1 U20881 ( .A1(n17985), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18002) );
  NOR2_X1 U20882 ( .A1(n17685), .A2(n17687), .ZN(n17681) );
  OAI211_X1 U20883 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17681), .A(
        n18478), .B(n17680), .ZN(n17682) );
  NAND4_X1 U20884 ( .A1(n17684), .A2(n17683), .A3(n18002), .A4(n17682), .ZN(
        P3_U2822) );
  NOR2_X1 U20885 ( .A1(n17685), .A2(n18134), .ZN(n17688) );
  NOR2_X1 U20886 ( .A1(n18069), .A2(n18644), .ZN(n18006) );
  AOI221_X1 U20887 ( .B1(n17688), .B2(n17687), .C1(n17686), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18006), .ZN(n17696) );
  NAND2_X1 U20888 ( .A1(n17690), .A2(n17689), .ZN(n17691) );
  XNOR2_X1 U20889 ( .A(n17691), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18008) );
  AOI21_X1 U20890 ( .B1(n17694), .B2(n17693), .A(n17692), .ZN(n18007) );
  AOI22_X1 U20891 ( .A1(n17755), .A2(n18008), .B1(n17759), .B2(n18007), .ZN(
        n17695) );
  OAI211_X1 U20892 ( .C1(n17518), .C2(n17697), .A(n17696), .B(n17695), .ZN(
        P3_U2823) );
  OAI21_X1 U20893 ( .B1(n18134), .B2(n17700), .A(n17758), .ZN(n17716) );
  AOI21_X1 U20894 ( .B1(n9707), .B2(n17699), .A(n17698), .ZN(n18021) );
  NOR2_X1 U20895 ( .A1(n18069), .A2(n18642), .ZN(n18018) );
  NOR3_X1 U20896 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17700), .A3(
        n18134), .ZN(n17701) );
  AOI211_X1 U20897 ( .C1(n17759), .C2(n18021), .A(n18018), .B(n17701), .ZN(
        n17706) );
  AOI21_X1 U20898 ( .B1(n17703), .B2(n18019), .A(n17702), .ZN(n18022) );
  AOI22_X1 U20899 ( .A1(n17755), .A2(n18022), .B1(n17704), .B2(n17738), .ZN(
        n17705) );
  OAI211_X1 U20900 ( .C1(n17707), .C2(n17716), .A(n17706), .B(n17705), .ZN(
        P3_U2824) );
  AOI21_X1 U20901 ( .B1(n17708), .B2(n17764), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17717) );
  AOI21_X1 U20902 ( .B1(n18016), .B2(n17710), .A(n17709), .ZN(n18027) );
  AOI22_X1 U20903 ( .A1(n17755), .A2(n18027), .B1(n17985), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17715) );
  AOI21_X1 U20904 ( .B1(n18016), .B2(n17712), .A(n17711), .ZN(n18026) );
  AOI22_X1 U20905 ( .A1(n17759), .A2(n18026), .B1(n17713), .B2(n17738), .ZN(
        n17714) );
  OAI211_X1 U20906 ( .C1(n17717), .C2(n17716), .A(n17715), .B(n17714), .ZN(
        P3_U2825) );
  AOI21_X1 U20907 ( .B1(n17720), .B2(n17719), .A(n17718), .ZN(n18038) );
  AOI22_X1 U20908 ( .A1(n17755), .A2(n18038), .B1(n9612), .B2(
        P3_REIP_REG_4__SCAN_IN), .ZN(n17731) );
  AOI21_X1 U20909 ( .B1(n17723), .B2(n17722), .A(n17721), .ZN(n18036) );
  AOI21_X1 U20910 ( .B1(n17726), .B2(n17725), .A(n17724), .ZN(n17742) );
  OAI22_X1 U20911 ( .A1(n17518), .A2(n17728), .B1(n17727), .B2(n17742), .ZN(
        n17729) );
  AOI21_X1 U20912 ( .B1(n17759), .B2(n18036), .A(n17729), .ZN(n17730) );
  OAI211_X1 U20913 ( .C1(n18134), .C2(n17732), .A(n17731), .B(n17730), .ZN(
        P3_U2826) );
  AOI21_X1 U20914 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17764), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17743) );
  AOI21_X1 U20915 ( .B1(n17735), .B2(n17734), .A(n17733), .ZN(n18044) );
  AOI22_X1 U20916 ( .A1(n17755), .A2(n18044), .B1(n9612), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n17741) );
  AOI21_X1 U20917 ( .B1(n18031), .B2(n17737), .A(n17736), .ZN(n18043) );
  AOI22_X1 U20918 ( .A1(n17759), .A2(n18043), .B1(n17739), .B2(n17738), .ZN(
        n17740) );
  OAI211_X1 U20919 ( .C1(n17743), .C2(n17742), .A(n17741), .B(n17740), .ZN(
        P3_U2827) );
  AOI21_X1 U20920 ( .B1(n17746), .B2(n17745), .A(n17744), .ZN(n18063) );
  INV_X1 U20921 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18634) );
  NOR2_X1 U20922 ( .A1(n18069), .A2(n18634), .ZN(n18050) );
  XNOR2_X1 U20923 ( .A(n17748), .B(n17747), .ZN(n18067) );
  OAI22_X1 U20924 ( .A1(n17518), .A2(n17749), .B1(n17767), .B2(n18067), .ZN(
        n17750) );
  AOI211_X1 U20925 ( .C1(n17755), .C2(n18063), .A(n18050), .B(n17750), .ZN(
        n17751) );
  OAI221_X1 U20926 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18134), .C1(
        n17752), .C2(n17764), .A(n17751), .ZN(P3_U2828) );
  NOR2_X1 U20927 ( .A1(n17763), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17753) );
  XOR2_X1 U20928 ( .A(n17753), .B(n17757), .Z(n18080) );
  INV_X1 U20929 ( .A(n18080), .ZN(n17754) );
  AOI22_X1 U20930 ( .A1(n17755), .A2(n17754), .B1(n9612), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17761) );
  AOI21_X1 U20931 ( .B1(n17757), .B2(n17762), .A(n17756), .ZN(n18075) );
  AOI22_X1 U20932 ( .A1(n17759), .A2(n18075), .B1(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17758), .ZN(n17760) );
  OAI211_X1 U20933 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n17518), .A(
        n17761), .B(n17760), .ZN(P3_U2829) );
  OAI21_X1 U20934 ( .B1(n17763), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17762), .ZN(n18082) );
  INV_X1 U20935 ( .A(n18082), .ZN(n18084) );
  NAND3_X1 U20936 ( .A1(n18710), .A2(n18613), .A3(n17764), .ZN(n17765) );
  AOI22_X1 U20937 ( .A1(n9612), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17765), .ZN(n17766) );
  OAI221_X1 U20938 ( .B1(n18084), .B2(n17768), .C1(n18082), .C2(n17767), .A(
        n17766), .ZN(P3_U2830) );
  INV_X1 U20939 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17770) );
  OAI21_X1 U20940 ( .B1(n18086), .B2(n17770), .A(n17769), .ZN(n17782) );
  INV_X1 U20941 ( .A(n18559), .ZN(n18570) );
  AOI21_X1 U20942 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n17771), .A(
        n18552), .ZN(n17830) );
  OAI22_X1 U20943 ( .A1(n18570), .A2(n17771), .B1(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17988), .ZN(n17772) );
  NOR2_X1 U20944 ( .A1(n17830), .A2(n17772), .ZN(n17810) );
  OAI211_X1 U20945 ( .C1(n17988), .C2(n17773), .A(n17810), .B(n17812), .ZN(
        n17793) );
  AOI22_X1 U20946 ( .A1(n18559), .A2(n17797), .B1(n18568), .B2(n17774), .ZN(
        n17777) );
  NAND2_X1 U20947 ( .A1(n18566), .A2(n17775), .ZN(n17776) );
  OAI211_X1 U20948 ( .C1(n17778), .C2(n17995), .A(n17777), .B(n17776), .ZN(
        n17779) );
  AOI211_X1 U20949 ( .C1(n18530), .C2(n17780), .A(n17793), .B(n17779), .ZN(
        n17788) );
  OAI211_X1 U20950 ( .C1(n18570), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n17788), .ZN(n17781) );
  AOI22_X1 U20951 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18051), .B1(
        n17782), .B2(n17781), .ZN(n17784) );
  NAND2_X1 U20952 ( .A1(n9612), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17783) );
  OAI211_X1 U20953 ( .C1(n17785), .C2(n17998), .A(n17784), .B(n17783), .ZN(
        P3_U2835) );
  AOI22_X1 U20954 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18071), .B1(
        n17786), .B2(n17807), .ZN(n17787) );
  AOI21_X1 U20955 ( .B1(n17788), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n17787), .ZN(n17789) );
  AOI21_X1 U20956 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n18051), .A(
        n17789), .ZN(n17791) );
  NAND2_X1 U20957 ( .A1(n9612), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17790) );
  OAI211_X1 U20958 ( .C1(n17792), .C2(n17998), .A(n17791), .B(n17790), .ZN(
        P3_U2836) );
  AOI211_X1 U20959 ( .C1(n18566), .C2(n17794), .A(n17797), .B(n17793), .ZN(
        n17795) );
  AOI211_X1 U20960 ( .C1(n17797), .C2(n17796), .A(n17795), .B(n18086), .ZN(
        n17798) );
  AOI21_X1 U20961 ( .B1(n18051), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17798), .ZN(n17800) );
  OAI211_X1 U20962 ( .C1(n17801), .C2(n17998), .A(n17800), .B(n17799), .ZN(
        n17802) );
  AOI21_X1 U20963 ( .B1(n17916), .B2(n17803), .A(n17802), .ZN(n17804) );
  OAI21_X1 U20964 ( .B1(n18079), .B2(n17805), .A(n17804), .ZN(P3_U2837) );
  AOI22_X1 U20965 ( .A1(n9612), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n17807), 
        .B2(n17806), .ZN(n17816) );
  INV_X1 U20966 ( .A(n18530), .ZN(n17927) );
  AOI21_X1 U20967 ( .B1(n17953), .B2(n17808), .A(n18051), .ZN(n17809) );
  OAI211_X1 U20968 ( .C1(n17811), .C2(n17927), .A(n17810), .B(n17809), .ZN(
        n17814) );
  NOR2_X1 U20969 ( .A1(n17818), .A2(n17814), .ZN(n17813) );
  AOI21_X1 U20970 ( .B1(n17813), .B2(n17812), .A(n9612), .ZN(n17821) );
  OAI211_X1 U20971 ( .C1(n17883), .C2(n17814), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17821), .ZN(n17815) );
  OAI211_X1 U20972 ( .C1(n17817), .C2(n17998), .A(n17816), .B(n17815), .ZN(
        P3_U2838) );
  OAI21_X1 U20973 ( .B1(n18051), .B2(n17819), .A(n17818), .ZN(n17820) );
  AOI22_X1 U20974 ( .A1(n9612), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n17821), 
        .B2(n17820), .ZN(n17822) );
  OAI21_X1 U20975 ( .B1(n17998), .B2(n17823), .A(n17822), .ZN(P3_U2839) );
  INV_X1 U20976 ( .A(n17839), .ZN(n17832) );
  OAI21_X1 U20977 ( .B1(n17844), .B2(n18035), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17829) );
  NOR2_X1 U20978 ( .A1(n17824), .A2(n17995), .ZN(n17894) );
  AOI21_X1 U20979 ( .B1(n18530), .B2(n17891), .A(n17894), .ZN(n17841) );
  NAND2_X1 U20980 ( .A1(n17927), .A2(n17995), .ZN(n17957) );
  NOR2_X1 U20981 ( .A1(n18570), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17826) );
  OAI21_X1 U20982 ( .B1(n17863), .B2(n17851), .A(n18559), .ZN(n17825) );
  OAI221_X1 U20983 ( .B1(n18035), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), 
        .C1(n18035), .C2(n17864), .A(n17825), .ZN(n17850) );
  AOI211_X1 U20984 ( .C1(n17827), .C2(n17957), .A(n17826), .B(n17850), .ZN(
        n17843) );
  OAI211_X1 U20985 ( .C1(n17964), .C2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n17841), .B(n17843), .ZN(n17828) );
  NOR3_X1 U20986 ( .A1(n17830), .A2(n17829), .A3(n17828), .ZN(n17831) );
  AOI221_X1 U20987 ( .B1(n17834), .B2(n17833), .C1(n17832), .C2(n17833), .A(
        n17831), .ZN(n17835) );
  AOI22_X1 U20988 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18051), .B1(
        n18071), .B2(n17835), .ZN(n17837) );
  OAI211_X1 U20989 ( .C1(n17838), .C2(n17998), .A(n17837), .B(n17836), .ZN(
        P3_U2840) );
  NAND3_X1 U20990 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18071), .A3(
        n17839), .ZN(n17862) );
  AOI22_X1 U20991 ( .A1(n9612), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n17982), 
        .B2(n17840), .ZN(n17847) );
  NAND2_X1 U20992 ( .A1(n18071), .A2(n17841), .ZN(n17884) );
  NOR2_X1 U20993 ( .A1(n18566), .A2(n18568), .ZN(n17903) );
  NAND2_X1 U20994 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17921), .ZN(
        n17974) );
  INV_X1 U20995 ( .A(n17974), .ZN(n17951) );
  NAND2_X1 U20996 ( .A1(n17873), .A2(n17951), .ZN(n17880) );
  OAI21_X1 U20997 ( .B1(n17842), .B2(n17880), .A(n18568), .ZN(n17852) );
  OAI211_X1 U20998 ( .C1(n17903), .C2(n17844), .A(n17852), .B(n17843), .ZN(
        n17845) );
  OAI211_X1 U20999 ( .C1(n17884), .C2(n17845), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18069), .ZN(n17846) );
  OAI211_X1 U21000 ( .C1(n17848), .C2(n17862), .A(n17847), .B(n17846), .ZN(
        P3_U2841) );
  AOI22_X1 U21001 ( .A1(n9612), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n17982), 
        .B2(n17849), .ZN(n17856) );
  AOI211_X1 U21002 ( .C1(n17851), .C2(n17957), .A(n17884), .B(n17850), .ZN(
        n17853) );
  AOI21_X1 U21003 ( .B1(n17853), .B2(n17852), .A(n9612), .ZN(n17859) );
  NOR3_X1 U21004 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17903), .A3(
        n18762), .ZN(n17854) );
  OAI21_X1 U21005 ( .B1(n17859), .B2(n17854), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17855) );
  OAI211_X1 U21006 ( .C1(n17857), .C2(n17862), .A(n17856), .B(n17855), .ZN(
        P3_U2842) );
  AOI22_X1 U21007 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17859), .B1(
        n17982), .B2(n17858), .ZN(n17861) );
  OAI211_X1 U21008 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17862), .A(
        n17861), .B(n17860), .ZN(P3_U2843) );
  NOR3_X1 U21009 ( .A1(n18054), .A2(n17863), .A3(n20793), .ZN(n17865) );
  OAI22_X1 U21010 ( .A1(n17988), .A2(n17865), .B1(n17864), .B2(n18035), .ZN(
        n17866) );
  AOI211_X1 U21011 ( .C1(n17867), .C2(n17957), .A(n17884), .B(n17866), .ZN(
        n17874) );
  AOI221_X1 U21012 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17874), 
        .C1(n17988), .C2(n17874), .A(n9612), .ZN(n17869) );
  AOI22_X1 U21013 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17869), .B1(
        n17980), .B2(n17868), .ZN(n17871) );
  OAI211_X1 U21014 ( .C1(n17998), .C2(n17872), .A(n17871), .B(n17870), .ZN(
        P3_U2844) );
  NAND2_X1 U21015 ( .A1(n17873), .A2(n17980), .ZN(n17888) );
  NOR3_X1 U21016 ( .A1(n9612), .A2(n17874), .A3(n20867), .ZN(n17875) );
  AOI21_X1 U21017 ( .B1(n17982), .B2(n17876), .A(n17875), .ZN(n17878) );
  OAI211_X1 U21018 ( .C1(n17888), .C2(n17879), .A(n17878), .B(n17877), .ZN(
        P3_U2845) );
  INV_X1 U21019 ( .A(n17889), .ZN(n17882) );
  NOR2_X1 U21020 ( .A1(n18570), .A2(n17921), .ZN(n17966) );
  AOI211_X1 U21021 ( .C1(n17880), .C2(n18568), .A(n10835), .B(n17966), .ZN(
        n17881) );
  NAND2_X1 U21022 ( .A1(n18566), .A2(n17904), .ZN(n17976) );
  OAI211_X1 U21023 ( .C1(n17964), .C2(n17882), .A(n17881), .B(n17976), .ZN(
        n17896) );
  OAI221_X1 U21024 ( .B1(n17884), .B2(n17883), .C1(n17884), .C2(n17896), .A(
        n18069), .ZN(n17887) );
  AOI22_X1 U21025 ( .A1(n9612), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n17982), 
        .B2(n17885), .ZN(n17886) );
  OAI221_X1 U21026 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17888), 
        .C1(n20793), .C2(n17887), .A(n17886), .ZN(P3_U2846) );
  OAI21_X1 U21027 ( .B1(n17889), .B2(n17937), .A(n10835), .ZN(n17897) );
  INV_X1 U21028 ( .A(n17890), .ZN(n17893) );
  AND2_X1 U21029 ( .A1(n17891), .A2(n18530), .ZN(n17892) );
  AOI222_X1 U21030 ( .A1(n17897), .A2(n17896), .B1(n17895), .B2(n17894), .C1(
        n17893), .C2(n17892), .ZN(n17901) );
  AOI22_X1 U21031 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18051), .B1(
        n17982), .B2(n17898), .ZN(n17900) );
  OAI211_X1 U21032 ( .C1(n17901), .C2(n18086), .A(n17900), .B(n17899), .ZN(
        P3_U2847) );
  INV_X1 U21033 ( .A(n17907), .ZN(n17902) );
  NOR2_X1 U21034 ( .A1(n17902), .A2(n17937), .ZN(n17912) );
  INV_X1 U21035 ( .A(n17903), .ZN(n18070) );
  AOI21_X1 U21036 ( .B1(n17942), .B2(n17951), .A(n18552), .ZN(n17929) );
  OAI21_X1 U21037 ( .B1(n17905), .B2(n17904), .A(n18566), .ZN(n17906) );
  OAI221_X1 U21038 ( .B1(n18570), .B2(n17907), .C1(n18570), .C2(n17921), .A(
        n17906), .ZN(n17908) );
  AOI211_X1 U21039 ( .C1(n17909), .C2(n18070), .A(n17929), .B(n17908), .ZN(
        n17910) );
  INV_X1 U21040 ( .A(n17910), .ZN(n17911) );
  MUX2_X1 U21041 ( .A(n17912), .B(n17911), .S(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n17913) );
  AOI21_X1 U21042 ( .B1(n18530), .B2(n17914), .A(n17913), .ZN(n17920) );
  AOI22_X1 U21043 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18051), .B1(
        n17985), .B2(P3_REIP_REG_14__SCAN_IN), .ZN(n17919) );
  AOI22_X1 U21044 ( .A1(n17982), .A2(n17917), .B1(n17916), .B2(n17915), .ZN(
        n17918) );
  OAI211_X1 U21045 ( .C1(n17920), .C2(n18086), .A(n17919), .B(n17918), .ZN(
        P3_U2848) );
  NOR2_X1 U21046 ( .A1(n18570), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17940) );
  AOI21_X1 U21047 ( .B1(n17922), .B2(n17921), .A(n18570), .ZN(n17923) );
  AOI21_X1 U21048 ( .B1(n17936), .B2(n18566), .A(n17923), .ZN(n17924) );
  INV_X1 U21049 ( .A(n17924), .ZN(n17960) );
  AOI21_X1 U21050 ( .B1(n17953), .B2(n17925), .A(n17960), .ZN(n17926) );
  OAI211_X1 U21051 ( .C1(n17928), .C2(n17927), .A(n17926), .B(n17976), .ZN(
        n17943) );
  NOR4_X1 U21052 ( .A1(n17940), .A2(n17929), .A3(n18086), .A4(n17943), .ZN(
        n17930) );
  AOI22_X1 U21053 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17932), .B1(
        n17980), .B2(n17931), .ZN(n17934) );
  OAI211_X1 U21054 ( .C1(n17935), .C2(n17998), .A(n17934), .B(n17933), .ZN(
        P3_U2849) );
  AOI21_X1 U21055 ( .B1(n17938), .B2(n17937), .A(n17936), .ZN(n17945) );
  NOR3_X1 U21056 ( .A1(n17940), .A2(n17939), .A3(n18568), .ZN(n17941) );
  AOI21_X1 U21057 ( .B1(n17951), .B2(n17942), .A(n17941), .ZN(n17944) );
  OAI22_X1 U21058 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17945), .B1(
        n17944), .B2(n17943), .ZN(n17949) );
  AOI22_X1 U21059 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18051), .B1(
        n17982), .B2(n17946), .ZN(n17948) );
  OAI211_X1 U21060 ( .C1(n18086), .C2(n17949), .A(n17948), .B(n17947), .ZN(
        P3_U2850) );
  AOI22_X1 U21061 ( .A1(n9612), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n17980), 
        .B2(n17950), .ZN(n17962) );
  AOI21_X1 U21062 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17951), .A(
        n18552), .ZN(n17956) );
  AOI22_X1 U21063 ( .A1(n18530), .A2(n17954), .B1(n17953), .B2(n17952), .ZN(
        n17977) );
  NAND3_X1 U21064 ( .A1(n18071), .A2(n17977), .A3(n17976), .ZN(n17955) );
  AOI211_X1 U21065 ( .C1(n17958), .C2(n17957), .A(n17956), .B(n17955), .ZN(
        n17968) );
  OAI21_X1 U21066 ( .B1(n18552), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17968), .ZN(n17959) );
  OAI211_X1 U21067 ( .C1(n17960), .C2(n17959), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18069), .ZN(n17961) );
  OAI211_X1 U21068 ( .C1(n17963), .C2(n17998), .A(n17962), .B(n17961), .ZN(
        P3_U2851) );
  INV_X1 U21069 ( .A(n17964), .ZN(n17965) );
  OAI21_X1 U21070 ( .B1(n17966), .B2(n10834), .A(n17965), .ZN(n17967) );
  AOI21_X1 U21071 ( .B1(n17968), .B2(n17967), .A(n9612), .ZN(n17970) );
  NOR2_X1 U21072 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n10834), .ZN(
        n17969) );
  AOI22_X1 U21073 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17970), .B1(
        n17980), .B2(n17969), .ZN(n17972) );
  OAI211_X1 U21074 ( .C1(n17998), .C2(n17973), .A(n17972), .B(n17971), .ZN(
        P3_U2852) );
  OAI211_X1 U21075 ( .C1(n18004), .C2(n18568), .A(n18053), .B(n17974), .ZN(
        n17975) );
  NAND4_X1 U21076 ( .A1(n17977), .A2(n18072), .A3(n17976), .A4(n17975), .ZN(
        n17979) );
  OAI221_X1 U21077 ( .B1(n17979), .B2(n18559), .C1(n17979), .C2(n17978), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17984) );
  AOI22_X1 U21078 ( .A1(n17982), .A2(n17981), .B1(n17980), .B2(n10834), .ZN(
        n17983) );
  OAI221_X1 U21079 ( .B1(n17985), .B2(n17984), .C1(n18069), .C2(n18648), .A(
        n17983), .ZN(P3_U2853) );
  OAI22_X1 U21080 ( .A1(n17988), .A2(n17987), .B1(n17986), .B2(n18035), .ZN(
        n17989) );
  NOR2_X1 U21081 ( .A1(n18054), .A2(n17989), .ZN(n18017) );
  OAI211_X1 U21082 ( .C1(n17990), .C2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n18017), .ZN(n18010) );
  AOI21_X1 U21083 ( .B1(n18076), .B2(n18010), .A(n18051), .ZN(n18005) );
  OAI22_X1 U21084 ( .A1(n18035), .A2(n18058), .B1(n17991), .B2(n18032), .ZN(
        n18046) );
  INV_X1 U21085 ( .A(n18046), .ZN(n18015) );
  NOR2_X1 U21086 ( .A1(n18015), .A2(n17992), .ZN(n18009) );
  NAND4_X1 U21087 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n18009), .A4(n18004), .ZN(
        n17993) );
  OAI21_X1 U21088 ( .B1(n17995), .B2(n17994), .A(n17993), .ZN(n18001) );
  INV_X1 U21089 ( .A(n17996), .ZN(n17997) );
  OAI22_X1 U21090 ( .A1(n17999), .A2(n17998), .B1(n18079), .B2(n17997), .ZN(
        n18000) );
  AOI21_X1 U21091 ( .B1(n18071), .B2(n18001), .A(n18000), .ZN(n18003) );
  OAI211_X1 U21092 ( .C1(n18005), .C2(n18004), .A(n18003), .B(n18002), .ZN(
        P3_U2854) );
  AOI21_X1 U21093 ( .B1(n18051), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18006), .ZN(n18014) );
  AOI22_X1 U21094 ( .A1(n18083), .A2(n18008), .B1(n18085), .B2(n18007), .ZN(
        n18013) );
  AND2_X1 U21095 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18009), .ZN(
        n18011) );
  OAI211_X1 U21096 ( .C1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n18011), .A(
        n18071), .B(n18010), .ZN(n18012) );
  NAND3_X1 U21097 ( .A1(n18014), .A2(n18013), .A3(n18012), .ZN(P3_U2855) );
  NOR3_X1 U21098 ( .A1(n18015), .A2(n18086), .A3(n18031), .ZN(n18037) );
  NAND2_X1 U21099 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18037), .ZN(
        n18030) );
  NOR2_X1 U21100 ( .A1(n18016), .A2(n18030), .ZN(n18020) );
  OAI21_X1 U21101 ( .B1(n18017), .B2(n18086), .A(n18072), .ZN(n18025) );
  AOI221_X1 U21102 ( .B1(n18020), .B2(n18019), .C1(n18025), .C2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(n18018), .ZN(n18024) );
  AOI22_X1 U21103 ( .A1(n18083), .A2(n18022), .B1(n18085), .B2(n18021), .ZN(
        n18023) );
  NAND2_X1 U21104 ( .A1(n18024), .A2(n18023), .ZN(P3_U2856) );
  AOI22_X1 U21105 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18025), .B1(
        n9612), .B2(P3_REIP_REG_5__SCAN_IN), .ZN(n18029) );
  AOI22_X1 U21106 ( .A1(n18083), .A2(n18027), .B1(n18085), .B2(n18026), .ZN(
        n18028) );
  OAI211_X1 U21107 ( .C1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n18030), .A(
        n18029), .B(n18028), .ZN(P3_U2857) );
  INV_X1 U21108 ( .A(n18058), .ZN(n18034) );
  AOI211_X1 U21109 ( .C1(n18053), .C2(n18032), .A(n18054), .B(n18031), .ZN(
        n18033) );
  OAI21_X1 U21110 ( .B1(n18035), .B2(n18034), .A(n18033), .ZN(n18045) );
  AOI21_X1 U21111 ( .B1(n18076), .B2(n18045), .A(n18051), .ZN(n18042) );
  AOI22_X1 U21112 ( .A1(n9612), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18085), .B2(
        n18036), .ZN(n18040) );
  AOI22_X1 U21113 ( .A1(n18038), .A2(n18083), .B1(n18037), .B2(n18041), .ZN(
        n18039) );
  OAI211_X1 U21114 ( .C1(n18042), .C2(n18041), .A(n18040), .B(n18039), .ZN(
        P3_U2858) );
  AOI22_X1 U21115 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18051), .B1(
        n9612), .B2(P3_REIP_REG_3__SCAN_IN), .ZN(n18049) );
  AOI22_X1 U21116 ( .A1(n18083), .A2(n18044), .B1(n18085), .B2(n18043), .ZN(
        n18048) );
  OAI211_X1 U21117 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n18046), .A(
        n18071), .B(n18045), .ZN(n18047) );
  NAND3_X1 U21118 ( .A1(n18049), .A2(n18048), .A3(n18047), .ZN(P3_U2859) );
  AOI21_X1 U21119 ( .B1(n18051), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n18050), .ZN(n18066) );
  NAND2_X1 U21120 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18052), .ZN(
        n18062) );
  NOR2_X1 U21121 ( .A1(n18727), .A2(n18709), .ZN(n18057) );
  OAI21_X1 U21122 ( .B1(n18709), .B2(n18054), .A(n18053), .ZN(n18055) );
  INV_X1 U21123 ( .A(n18055), .ZN(n18056) );
  AOI21_X1 U21124 ( .B1(n18057), .B2(n18566), .A(n18056), .ZN(n18060) );
  NAND2_X1 U21125 ( .A1(n18566), .A2(n18058), .ZN(n18059) );
  OAI221_X1 U21126 ( .B1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n18062), .C1(
        n18061), .C2(n18060), .A(n18059), .ZN(n18064) );
  AOI22_X1 U21127 ( .A1(n18071), .A2(n18064), .B1(n18083), .B2(n18063), .ZN(
        n18065) );
  OAI211_X1 U21128 ( .C1(n18068), .C2(n18067), .A(n18066), .B(n18065), .ZN(
        P3_U2860) );
  INV_X1 U21129 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18633) );
  NOR2_X1 U21130 ( .A1(n18069), .A2(n18633), .ZN(n18074) );
  NAND3_X1 U21131 ( .A1(n18071), .A2(n18727), .A3(n18070), .ZN(n18088) );
  AOI21_X1 U21132 ( .B1(n18072), .B2(n18088), .A(n18709), .ZN(n18073) );
  AOI211_X1 U21133 ( .C1(n18075), .C2(n18085), .A(n18074), .B(n18073), .ZN(
        n18078) );
  OAI211_X1 U21134 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18559), .A(
        n18076), .B(n18709), .ZN(n18077) );
  OAI211_X1 U21135 ( .C1(n18080), .C2(n18079), .A(n18078), .B(n18077), .ZN(
        P3_U2861) );
  AND2_X1 U21136 ( .A1(n9612), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18081) );
  AOI221_X1 U21137 ( .B1(n18085), .B2(n18084), .C1(n18083), .C2(n18082), .A(
        n18081), .ZN(n18089) );
  OAI211_X1 U21138 ( .C1(n18559), .C2(n18086), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n18069), .ZN(n18087) );
  NAND3_X1 U21139 ( .A1(n18089), .A2(n18088), .A3(n18087), .ZN(P3_U2862) );
  AOI211_X1 U21140 ( .C1(n18091), .C2(n18090), .A(n18762), .B(n18710), .ZN(
        n18595) );
  OAI21_X1 U21141 ( .B1(n18595), .B2(n18141), .A(n18096), .ZN(n18092) );
  OAI221_X1 U21142 ( .B1(n18392), .B2(n18744), .C1(n18392), .C2(n18096), .A(
        n18092), .ZN(P3_U2863) );
  INV_X1 U21143 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18583) );
  NOR2_X1 U21144 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18580), .ZN(
        n18281) );
  INV_X1 U21145 ( .A(n18281), .ZN(n18279) );
  NOR2_X1 U21146 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18583), .ZN(
        n18371) );
  NAND2_X1 U21147 ( .A1(n18445), .A2(n18371), .ZN(n18395) );
  AND2_X1 U21148 ( .A1(n18279), .A2(n18395), .ZN(n18094) );
  OAI22_X1 U21149 ( .A1(n18095), .A2(n18583), .B1(n18094), .B2(n18093), .ZN(
        P3_U2866) );
  NOR2_X1 U21150 ( .A1(n18584), .A2(n18096), .ZN(P3_U2867) );
  NOR2_X1 U21151 ( .A1(n18583), .A2(n18280), .ZN(n18476) );
  NAND2_X1 U21152 ( .A1(n18392), .A2(n18476), .ZN(n18470) );
  INV_X1 U21153 ( .A(n18470), .ZN(n18448) );
  NOR2_X1 U21154 ( .A1(n18580), .A2(n18583), .ZN(n18419) );
  NAND2_X1 U21155 ( .A1(n18419), .A2(n18575), .ZN(n18417) );
  NOR2_X2 U21156 ( .A1(n18392), .A2(n18417), .ZN(n18524) );
  NOR2_X1 U21157 ( .A1(n18448), .A2(n18524), .ZN(n18441) );
  NAND2_X1 U21158 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18574) );
  INV_X1 U21159 ( .A(n18419), .ZN(n18097) );
  NOR2_X2 U21160 ( .A1(n18574), .A2(n18097), .ZN(n18471) );
  NAND2_X1 U21161 ( .A1(n18575), .A2(n18392), .ZN(n18576) );
  NAND2_X1 U21162 ( .A1(n18580), .A2(n18583), .ZN(n18168) );
  NOR2_X1 U21163 ( .A1(n18576), .A2(n18168), .ZN(n18184) );
  CLKBUF_X1 U21164 ( .A(n18184), .Z(n18209) );
  NOR2_X1 U21165 ( .A1(n18471), .A2(n18209), .ZN(n18170) );
  OAI21_X1 U21166 ( .B1(n18392), .B2(n20828), .A(n18396), .ZN(n18347) );
  OAI22_X1 U21167 ( .A1(n18441), .A2(n18134), .B1(n18170), .B2(n18347), .ZN(
        n18139) );
  AND2_X1 U21168 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18478), .ZN(n18479) );
  NOR2_X2 U21169 ( .A1(n18142), .A2(n18098), .ZN(n18473) );
  NOR2_X1 U21170 ( .A1(n18603), .A2(n18170), .ZN(n18132) );
  AOI22_X1 U21171 ( .A1(n18524), .A2(n18479), .B1(n18473), .B2(n18132), .ZN(
        n18103) );
  NAND2_X1 U21172 ( .A1(n18478), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18452) );
  INV_X1 U21173 ( .A(n18452), .ZN(n18474) );
  NAND2_X1 U21174 ( .A1(n18100), .A2(n18099), .ZN(n18135) );
  NOR2_X1 U21175 ( .A1(n18101), .A2(n18135), .ZN(n18447) );
  AOI22_X1 U21176 ( .A1(n18474), .A2(n18448), .B1(n18209), .B2(n18447), .ZN(
        n18102) );
  OAI211_X1 U21177 ( .C1(n18104), .C2(n18139), .A(n18103), .B(n18102), .ZN(
        P3_U2868) );
  NOR2_X2 U21178 ( .A1(n18134), .A2(n15128), .ZN(n18485) );
  AND2_X1 U21179 ( .A1(n18396), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18483) );
  AOI22_X1 U21180 ( .A1(n18448), .A2(n18485), .B1(n18132), .B2(n18483), .ZN(
        n18106) );
  AND2_X1 U21181 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18478), .ZN(n18484) );
  NOR2_X1 U21182 ( .A1(n18750), .A2(n18135), .ZN(n18145) );
  AOI22_X1 U21183 ( .A1(n18524), .A2(n18484), .B1(n18209), .B2(n18145), .ZN(
        n18105) );
  OAI211_X1 U21184 ( .C1(n18107), .C2(n18139), .A(n18106), .B(n18105), .ZN(
        P3_U2869) );
  AND2_X1 U21185 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18478), .ZN(n18489) );
  NOR2_X2 U21186 ( .A1(n18142), .A2(n18108), .ZN(n18490) );
  AOI22_X1 U21187 ( .A1(n18524), .A2(n18489), .B1(n18132), .B2(n18490), .ZN(
        n18111) );
  AND2_X1 U21188 ( .A1(n18478), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18491) );
  NOR2_X1 U21189 ( .A1(n18109), .A2(n18135), .ZN(n18148) );
  AOI22_X1 U21190 ( .A1(n18448), .A2(n18491), .B1(n18184), .B2(n18148), .ZN(
        n18110) );
  OAI211_X1 U21191 ( .C1(n18112), .C2(n18139), .A(n18111), .B(n18110), .ZN(
        P3_U2870) );
  AND2_X1 U21192 ( .A1(n18478), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18496) );
  NOR2_X2 U21193 ( .A1(n18142), .A2(n18113), .ZN(n18495) );
  AOI22_X1 U21194 ( .A1(n18448), .A2(n18496), .B1(n18132), .B2(n18495), .ZN(
        n18116) );
  AND2_X1 U21195 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18478), .ZN(n18497) );
  NOR2_X1 U21196 ( .A1(n18114), .A2(n18135), .ZN(n18151) );
  AOI22_X1 U21197 ( .A1(n18524), .A2(n18497), .B1(n18184), .B2(n18151), .ZN(
        n18115) );
  OAI211_X1 U21198 ( .C1(n18117), .C2(n18139), .A(n18116), .B(n18115), .ZN(
        P3_U2871) );
  AND2_X1 U21199 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18478), .ZN(n18502) );
  NOR2_X2 U21200 ( .A1(n18142), .A2(n18118), .ZN(n18501) );
  AOI22_X1 U21201 ( .A1(n18524), .A2(n18502), .B1(n18132), .B2(n18501), .ZN(
        n18121) );
  AND2_X1 U21202 ( .A1(n18478), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18503) );
  NOR2_X1 U21203 ( .A1(n18119), .A2(n18135), .ZN(n18154) );
  AOI22_X1 U21204 ( .A1(n18448), .A2(n18503), .B1(n18184), .B2(n18154), .ZN(
        n18120) );
  OAI211_X1 U21205 ( .C1(n18122), .C2(n18139), .A(n18121), .B(n18120), .ZN(
        P3_U2872) );
  NOR2_X2 U21206 ( .A1(n18134), .A2(n15113), .ZN(n18509) );
  NOR2_X2 U21207 ( .A1(n18142), .A2(n18123), .ZN(n18507) );
  AOI22_X1 U21208 ( .A1(n18448), .A2(n18509), .B1(n18132), .B2(n18507), .ZN(
        n18126) );
  AND2_X1 U21209 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18478), .ZN(n18508) );
  NOR2_X1 U21210 ( .A1(n18124), .A2(n18135), .ZN(n18157) );
  AOI22_X1 U21211 ( .A1(n18524), .A2(n18508), .B1(n18184), .B2(n18157), .ZN(
        n18125) );
  OAI211_X1 U21212 ( .C1(n20890), .C2(n18139), .A(n18126), .B(n18125), .ZN(
        P3_U2873) );
  AND2_X1 U21213 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18478), .ZN(n18515) );
  NOR2_X2 U21214 ( .A1(n18142), .A2(n20932), .ZN(n18513) );
  AOI22_X1 U21215 ( .A1(n18524), .A2(n18515), .B1(n18132), .B2(n18513), .ZN(
        n18129) );
  AND2_X1 U21216 ( .A1(n18478), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18514) );
  NOR2_X1 U21217 ( .A1(n18127), .A2(n18135), .ZN(n18160) );
  AOI22_X1 U21218 ( .A1(n18448), .A2(n18514), .B1(n18184), .B2(n18160), .ZN(
        n18128) );
  OAI211_X1 U21219 ( .C1(n18130), .C2(n18139), .A(n18129), .B(n18128), .ZN(
        P3_U2874) );
  AND2_X1 U21220 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18478), .ZN(n18523) );
  NOR2_X2 U21221 ( .A1(n18131), .A2(n18142), .ZN(n18520) );
  AOI22_X1 U21222 ( .A1(n18448), .A2(n18523), .B1(n18132), .B2(n18520), .ZN(
        n18138) );
  NOR2_X2 U21223 ( .A1(n18134), .A2(n18133), .ZN(n18522) );
  NOR2_X1 U21224 ( .A1(n18136), .A2(n18135), .ZN(n18163) );
  AOI22_X1 U21225 ( .A1(n18524), .A2(n18522), .B1(n18184), .B2(n18163), .ZN(
        n18137) );
  OAI211_X1 U21226 ( .C1(n18140), .C2(n18139), .A(n18138), .B(n18137), .ZN(
        P3_U2875) );
  INV_X1 U21227 ( .A(n18447), .ZN(n18482) );
  INV_X1 U21228 ( .A(n18168), .ZN(n18193) );
  NOR2_X1 U21229 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18392), .ZN(
        n18325) );
  NAND2_X1 U21230 ( .A1(n18193), .A2(n18325), .ZN(n18169) );
  NAND2_X1 U21231 ( .A1(n18575), .A2(n18472), .ZN(n18326) );
  NOR2_X1 U21232 ( .A1(n18168), .A2(n18326), .ZN(n18164) );
  AOI22_X1 U21233 ( .A1(n18474), .A2(n18471), .B1(n18473), .B2(n18164), .ZN(
        n18144) );
  NOR2_X1 U21234 ( .A1(n18142), .A2(n18141), .ZN(n18475) );
  INV_X1 U21235 ( .A(n18475), .ZN(n18192) );
  NOR2_X1 U21236 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18192), .ZN(
        n18418) );
  AOI22_X1 U21237 ( .A1(n18478), .A2(n18476), .B1(n18193), .B2(n18418), .ZN(
        n18165) );
  AOI22_X1 U21238 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18165), .B1(
        n18448), .B2(n18479), .ZN(n18143) );
  OAI211_X1 U21239 ( .C1(n18482), .C2(n18169), .A(n18144), .B(n18143), .ZN(
        P3_U2876) );
  INV_X1 U21240 ( .A(n18145), .ZN(n18488) );
  AOI22_X1 U21241 ( .A1(n18448), .A2(n18484), .B1(n18483), .B2(n18164), .ZN(
        n18147) );
  AOI22_X1 U21242 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18165), .B1(
        n18471), .B2(n18485), .ZN(n18146) );
  OAI211_X1 U21243 ( .C1(n18488), .C2(n18169), .A(n18147), .B(n18146), .ZN(
        P3_U2877) );
  INV_X1 U21244 ( .A(n18148), .ZN(n18494) );
  AOI22_X1 U21245 ( .A1(n18471), .A2(n18491), .B1(n18490), .B2(n18164), .ZN(
        n18150) );
  AOI22_X1 U21246 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18165), .B1(
        n18448), .B2(n18489), .ZN(n18149) );
  OAI211_X1 U21247 ( .C1(n18494), .C2(n18169), .A(n18150), .B(n18149), .ZN(
        P3_U2878) );
  INV_X1 U21248 ( .A(n18151), .ZN(n18500) );
  AOI22_X1 U21249 ( .A1(n18448), .A2(n18497), .B1(n18495), .B2(n18164), .ZN(
        n18153) );
  AOI22_X1 U21250 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18165), .B1(
        n18471), .B2(n18496), .ZN(n18152) );
  OAI211_X1 U21251 ( .C1(n18500), .C2(n18169), .A(n18153), .B(n18152), .ZN(
        P3_U2879) );
  INV_X1 U21252 ( .A(n18154), .ZN(n18506) );
  AOI22_X1 U21253 ( .A1(n18471), .A2(n18503), .B1(n18501), .B2(n18164), .ZN(
        n18156) );
  AOI22_X1 U21254 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18165), .B1(
        n18448), .B2(n18502), .ZN(n18155) );
  OAI211_X1 U21255 ( .C1(n18506), .C2(n18169), .A(n18156), .B(n18155), .ZN(
        P3_U2880) );
  INV_X1 U21256 ( .A(n18157), .ZN(n18512) );
  AOI22_X1 U21257 ( .A1(n18471), .A2(n18509), .B1(n18507), .B2(n18164), .ZN(
        n18159) );
  AOI22_X1 U21258 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18165), .B1(
        n18448), .B2(n18508), .ZN(n18158) );
  OAI211_X1 U21259 ( .C1(n18512), .C2(n18169), .A(n18159), .B(n18158), .ZN(
        P3_U2881) );
  INV_X1 U21260 ( .A(n18160), .ZN(n18518) );
  AOI22_X1 U21261 ( .A1(n18448), .A2(n18515), .B1(n18513), .B2(n18164), .ZN(
        n18162) );
  AOI22_X1 U21262 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18165), .B1(
        n18471), .B2(n18514), .ZN(n18161) );
  OAI211_X1 U21263 ( .C1(n18518), .C2(n18169), .A(n18162), .B(n18161), .ZN(
        P3_U2882) );
  AOI22_X1 U21264 ( .A1(n18448), .A2(n18522), .B1(n18520), .B2(n18164), .ZN(
        n18167) );
  AOI22_X1 U21265 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18165), .B1(
        n18471), .B2(n18523), .ZN(n18166) );
  OAI211_X1 U21266 ( .C1(n18528), .C2(n18169), .A(n18167), .B(n18166), .ZN(
        P3_U2883) );
  NOR2_X1 U21267 ( .A1(n18575), .A2(n18168), .ZN(n18236) );
  NAND2_X1 U21268 ( .A1(n18236), .A2(n18392), .ZN(n18191) );
  INV_X1 U21269 ( .A(n18169), .ZN(n18231) );
  INV_X1 U21270 ( .A(n18191), .ZN(n18252) );
  NOR2_X1 U21271 ( .A1(n18231), .A2(n18252), .ZN(n18214) );
  INV_X1 U21272 ( .A(n18445), .ZN(n18348) );
  AOI221_X1 U21273 ( .B1(n18214), .B2(n18348), .C1(n18214), .C2(n18170), .A(
        n18347), .ZN(n18171) );
  INV_X1 U21274 ( .A(n18171), .ZN(n18188) );
  NOR2_X1 U21275 ( .A1(n18603), .A2(n18214), .ZN(n18187) );
  AOI22_X1 U21276 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18188), .B1(
        n18473), .B2(n18187), .ZN(n18173) );
  AOI22_X1 U21277 ( .A1(n18474), .A2(n18209), .B1(n18471), .B2(n18479), .ZN(
        n18172) );
  OAI211_X1 U21278 ( .C1(n18482), .C2(n18191), .A(n18173), .B(n18172), .ZN(
        P3_U2884) );
  AOI22_X1 U21279 ( .A1(n18471), .A2(n18484), .B1(n18483), .B2(n18187), .ZN(
        n18175) );
  AOI22_X1 U21280 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18188), .B1(
        n18184), .B2(n18485), .ZN(n18174) );
  OAI211_X1 U21281 ( .C1(n18488), .C2(n18191), .A(n18175), .B(n18174), .ZN(
        P3_U2885) );
  AOI22_X1 U21282 ( .A1(n18471), .A2(n18489), .B1(n18490), .B2(n18187), .ZN(
        n18177) );
  AOI22_X1 U21283 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18188), .B1(
        n18184), .B2(n18491), .ZN(n18176) );
  OAI211_X1 U21284 ( .C1(n18494), .C2(n18191), .A(n18177), .B(n18176), .ZN(
        P3_U2886) );
  AOI22_X1 U21285 ( .A1(n18471), .A2(n18497), .B1(n18495), .B2(n18187), .ZN(
        n18179) );
  AOI22_X1 U21286 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18188), .B1(
        n18184), .B2(n18496), .ZN(n18178) );
  OAI211_X1 U21287 ( .C1(n18500), .C2(n18191), .A(n18179), .B(n18178), .ZN(
        P3_U2887) );
  AOI22_X1 U21288 ( .A1(n18471), .A2(n18502), .B1(n18501), .B2(n18187), .ZN(
        n18181) );
  AOI22_X1 U21289 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18188), .B1(
        n18184), .B2(n18503), .ZN(n18180) );
  OAI211_X1 U21290 ( .C1(n18506), .C2(n18191), .A(n18181), .B(n18180), .ZN(
        P3_U2888) );
  AOI22_X1 U21291 ( .A1(n18209), .A2(n18509), .B1(n18507), .B2(n18187), .ZN(
        n18183) );
  AOI22_X1 U21292 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18188), .B1(
        n18471), .B2(n18508), .ZN(n18182) );
  OAI211_X1 U21293 ( .C1(n18512), .C2(n18191), .A(n18183), .B(n18182), .ZN(
        P3_U2889) );
  AOI22_X1 U21294 ( .A1(n18471), .A2(n18515), .B1(n18513), .B2(n18187), .ZN(
        n18186) );
  AOI22_X1 U21295 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18188), .B1(
        n18184), .B2(n18514), .ZN(n18185) );
  OAI211_X1 U21296 ( .C1(n18518), .C2(n18191), .A(n18186), .B(n18185), .ZN(
        P3_U2890) );
  AOI22_X1 U21297 ( .A1(n18209), .A2(n18523), .B1(n18520), .B2(n18187), .ZN(
        n18190) );
  AOI22_X1 U21298 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18188), .B1(
        n18471), .B2(n18522), .ZN(n18189) );
  OAI211_X1 U21299 ( .C1(n18528), .C2(n18191), .A(n18190), .B(n18189), .ZN(
        P3_U2891) );
  NAND2_X1 U21300 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18236), .ZN(
        n18213) );
  AND2_X1 U21301 ( .A1(n18472), .A2(n18236), .ZN(n18208) );
  AOI22_X1 U21302 ( .A1(n18209), .A2(n18479), .B1(n18473), .B2(n18208), .ZN(
        n18195) );
  AOI21_X1 U21303 ( .B1(n18575), .B2(n18348), .A(n18192), .ZN(n18282) );
  NAND2_X1 U21304 ( .A1(n18193), .A2(n18282), .ZN(n18210) );
  AOI22_X1 U21305 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18210), .B1(
        n18474), .B2(n18231), .ZN(n18194) );
  OAI211_X1 U21306 ( .C1(n18482), .C2(n18213), .A(n18195), .B(n18194), .ZN(
        P3_U2892) );
  AOI22_X1 U21307 ( .A1(n18209), .A2(n18484), .B1(n18483), .B2(n18208), .ZN(
        n18197) );
  AOI22_X1 U21308 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18210), .B1(
        n18485), .B2(n18231), .ZN(n18196) );
  OAI211_X1 U21309 ( .C1(n18488), .C2(n18213), .A(n18197), .B(n18196), .ZN(
        P3_U2893) );
  AOI22_X1 U21310 ( .A1(n18209), .A2(n18489), .B1(n18490), .B2(n18208), .ZN(
        n18199) );
  AOI22_X1 U21311 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18210), .B1(
        n18491), .B2(n18231), .ZN(n18198) );
  OAI211_X1 U21312 ( .C1(n18494), .C2(n18213), .A(n18199), .B(n18198), .ZN(
        P3_U2894) );
  AOI22_X1 U21313 ( .A1(n18209), .A2(n18497), .B1(n18495), .B2(n18208), .ZN(
        n18201) );
  AOI22_X1 U21314 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18210), .B1(
        n18496), .B2(n18231), .ZN(n18200) );
  OAI211_X1 U21315 ( .C1(n18500), .C2(n18213), .A(n18201), .B(n18200), .ZN(
        P3_U2895) );
  AOI22_X1 U21316 ( .A1(n18209), .A2(n18502), .B1(n18501), .B2(n18208), .ZN(
        n18203) );
  AOI22_X1 U21317 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18210), .B1(
        n18503), .B2(n18231), .ZN(n18202) );
  OAI211_X1 U21318 ( .C1(n18506), .C2(n18213), .A(n18203), .B(n18202), .ZN(
        P3_U2896) );
  AOI22_X1 U21319 ( .A1(n18509), .A2(n18231), .B1(n18507), .B2(n18208), .ZN(
        n18205) );
  AOI22_X1 U21320 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18210), .B1(
        n18209), .B2(n18508), .ZN(n18204) );
  OAI211_X1 U21321 ( .C1(n18512), .C2(n18213), .A(n18205), .B(n18204), .ZN(
        P3_U2897) );
  AOI22_X1 U21322 ( .A1(n18514), .A2(n18231), .B1(n18513), .B2(n18208), .ZN(
        n18207) );
  AOI22_X1 U21323 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18210), .B1(
        n18209), .B2(n18515), .ZN(n18206) );
  OAI211_X1 U21324 ( .C1(n18518), .C2(n18213), .A(n18207), .B(n18206), .ZN(
        P3_U2898) );
  AOI22_X1 U21325 ( .A1(n18209), .A2(n18522), .B1(n18520), .B2(n18208), .ZN(
        n18212) );
  AOI22_X1 U21326 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18210), .B1(
        n18523), .B2(n18231), .ZN(n18211) );
  OAI211_X1 U21327 ( .C1(n18528), .C2(n18213), .A(n18212), .B(n18211), .ZN(
        P3_U2899) );
  INV_X1 U21328 ( .A(n18576), .ZN(n18394) );
  NAND2_X1 U21329 ( .A1(n18394), .A2(n18281), .ZN(n18235) );
  INV_X1 U21330 ( .A(n18213), .ZN(n18274) );
  INV_X1 U21331 ( .A(n18235), .ZN(n18298) );
  NOR2_X1 U21332 ( .A1(n18274), .A2(n18298), .ZN(n18257) );
  NOR2_X1 U21333 ( .A1(n18603), .A2(n18257), .ZN(n18230) );
  AOI22_X1 U21334 ( .A1(n18474), .A2(n18252), .B1(n18473), .B2(n18230), .ZN(
        n18217) );
  OAI21_X1 U21335 ( .B1(n18214), .B2(n18348), .A(n18257), .ZN(n18215) );
  OAI211_X1 U21336 ( .C1(n18298), .C2(n20828), .A(n18396), .B(n18215), .ZN(
        n18232) );
  AOI22_X1 U21337 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18232), .B1(
        n18479), .B2(n18231), .ZN(n18216) );
  OAI211_X1 U21338 ( .C1(n18482), .C2(n18235), .A(n18217), .B(n18216), .ZN(
        P3_U2900) );
  AOI22_X1 U21339 ( .A1(n18485), .A2(n18252), .B1(n18483), .B2(n18230), .ZN(
        n18219) );
  AOI22_X1 U21340 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18232), .B1(
        n18484), .B2(n18231), .ZN(n18218) );
  OAI211_X1 U21341 ( .C1(n18488), .C2(n18235), .A(n18219), .B(n18218), .ZN(
        P3_U2901) );
  AOI22_X1 U21342 ( .A1(n18490), .A2(n18230), .B1(n18489), .B2(n18231), .ZN(
        n18221) );
  AOI22_X1 U21343 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18232), .B1(
        n18491), .B2(n18252), .ZN(n18220) );
  OAI211_X1 U21344 ( .C1(n18494), .C2(n18235), .A(n18221), .B(n18220), .ZN(
        P3_U2902) );
  AOI22_X1 U21345 ( .A1(n18496), .A2(n18252), .B1(n18495), .B2(n18230), .ZN(
        n18223) );
  AOI22_X1 U21346 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18232), .B1(
        n18497), .B2(n18231), .ZN(n18222) );
  OAI211_X1 U21347 ( .C1(n18500), .C2(n18235), .A(n18223), .B(n18222), .ZN(
        P3_U2903) );
  AOI22_X1 U21348 ( .A1(n18502), .A2(n18231), .B1(n18501), .B2(n18230), .ZN(
        n18225) );
  AOI22_X1 U21349 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18232), .B1(
        n18503), .B2(n18252), .ZN(n18224) );
  OAI211_X1 U21350 ( .C1(n18506), .C2(n18235), .A(n18225), .B(n18224), .ZN(
        P3_U2904) );
  AOI22_X1 U21351 ( .A1(n18509), .A2(n18252), .B1(n18507), .B2(n18230), .ZN(
        n18227) );
  AOI22_X1 U21352 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18232), .B1(
        n18508), .B2(n18231), .ZN(n18226) );
  OAI211_X1 U21353 ( .C1(n18512), .C2(n18235), .A(n18227), .B(n18226), .ZN(
        P3_U2905) );
  AOI22_X1 U21354 ( .A1(n18515), .A2(n18231), .B1(n18513), .B2(n18230), .ZN(
        n18229) );
  AOI22_X1 U21355 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18232), .B1(
        n18514), .B2(n18252), .ZN(n18228) );
  OAI211_X1 U21356 ( .C1(n18518), .C2(n18235), .A(n18229), .B(n18228), .ZN(
        P3_U2906) );
  AOI22_X1 U21357 ( .A1(n18522), .A2(n18231), .B1(n18520), .B2(n18230), .ZN(
        n18234) );
  AOI22_X1 U21358 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18232), .B1(
        n18523), .B2(n18252), .ZN(n18233) );
  OAI211_X1 U21359 ( .C1(n18528), .C2(n18235), .A(n18234), .B(n18233), .ZN(
        P3_U2907) );
  NAND2_X1 U21360 ( .A1(n18325), .A2(n18281), .ZN(n18256) );
  NOR2_X1 U21361 ( .A1(n18326), .A2(n18279), .ZN(n18251) );
  AOI22_X1 U21362 ( .A1(n18474), .A2(n18274), .B1(n18473), .B2(n18251), .ZN(
        n18238) );
  AOI22_X1 U21363 ( .A1(n18478), .A2(n18236), .B1(n18418), .B2(n18281), .ZN(
        n18253) );
  AOI22_X1 U21364 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18253), .B1(
        n18479), .B2(n18252), .ZN(n18237) );
  OAI211_X1 U21365 ( .C1(n18482), .C2(n18256), .A(n18238), .B(n18237), .ZN(
        P3_U2908) );
  AOI22_X1 U21366 ( .A1(n18484), .A2(n18252), .B1(n18483), .B2(n18251), .ZN(
        n18240) );
  AOI22_X1 U21367 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18253), .B1(
        n18485), .B2(n18274), .ZN(n18239) );
  OAI211_X1 U21368 ( .C1(n18488), .C2(n18256), .A(n18240), .B(n18239), .ZN(
        P3_U2909) );
  AOI22_X1 U21369 ( .A1(n18490), .A2(n18251), .B1(n18489), .B2(n18252), .ZN(
        n18242) );
  AOI22_X1 U21370 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18253), .B1(
        n18491), .B2(n18274), .ZN(n18241) );
  OAI211_X1 U21371 ( .C1(n18494), .C2(n18256), .A(n18242), .B(n18241), .ZN(
        P3_U2910) );
  AOI22_X1 U21372 ( .A1(n18496), .A2(n18274), .B1(n18495), .B2(n18251), .ZN(
        n18244) );
  AOI22_X1 U21373 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18253), .B1(
        n18497), .B2(n18252), .ZN(n18243) );
  OAI211_X1 U21374 ( .C1(n18500), .C2(n18256), .A(n18244), .B(n18243), .ZN(
        P3_U2911) );
  AOI22_X1 U21375 ( .A1(n18503), .A2(n18274), .B1(n18501), .B2(n18251), .ZN(
        n18246) );
  AOI22_X1 U21376 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18253), .B1(
        n18502), .B2(n18252), .ZN(n18245) );
  OAI211_X1 U21377 ( .C1(n18506), .C2(n18256), .A(n18246), .B(n18245), .ZN(
        P3_U2912) );
  AOI22_X1 U21378 ( .A1(n18509), .A2(n18274), .B1(n18507), .B2(n18251), .ZN(
        n18248) );
  AOI22_X1 U21379 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18253), .B1(
        n18508), .B2(n18252), .ZN(n18247) );
  OAI211_X1 U21380 ( .C1(n18512), .C2(n18256), .A(n18248), .B(n18247), .ZN(
        P3_U2913) );
  AOI22_X1 U21381 ( .A1(n18514), .A2(n18274), .B1(n18513), .B2(n18251), .ZN(
        n18250) );
  AOI22_X1 U21382 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18253), .B1(
        n18515), .B2(n18252), .ZN(n18249) );
  OAI211_X1 U21383 ( .C1(n18518), .C2(n18256), .A(n18250), .B(n18249), .ZN(
        P3_U2914) );
  AOI22_X1 U21384 ( .A1(n18522), .A2(n18252), .B1(n18520), .B2(n18251), .ZN(
        n18255) );
  AOI22_X1 U21385 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18253), .B1(
        n18523), .B2(n18274), .ZN(n18254) );
  OAI211_X1 U21386 ( .C1(n18528), .C2(n18256), .A(n18255), .B(n18254), .ZN(
        P3_U2915) );
  INV_X1 U21387 ( .A(n18343), .ZN(n18278) );
  INV_X1 U21388 ( .A(n18256), .ZN(n18320) );
  NOR2_X1 U21389 ( .A1(n18320), .A2(n18343), .ZN(n18303) );
  NOR2_X1 U21390 ( .A1(n18603), .A2(n18303), .ZN(n18273) );
  AOI22_X1 U21391 ( .A1(n18474), .A2(n18298), .B1(n18473), .B2(n18273), .ZN(
        n18260) );
  OAI21_X1 U21392 ( .B1(n18257), .B2(n18348), .A(n18303), .ZN(n18258) );
  OAI211_X1 U21393 ( .C1(n18343), .C2(n20828), .A(n18396), .B(n18258), .ZN(
        n18275) );
  AOI22_X1 U21394 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18275), .B1(
        n18479), .B2(n18274), .ZN(n18259) );
  OAI211_X1 U21395 ( .C1(n18482), .C2(n18278), .A(n18260), .B(n18259), .ZN(
        P3_U2916) );
  AOI22_X1 U21396 ( .A1(n18485), .A2(n18298), .B1(n18483), .B2(n18273), .ZN(
        n18262) );
  AOI22_X1 U21397 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18275), .B1(
        n18484), .B2(n18274), .ZN(n18261) );
  OAI211_X1 U21398 ( .C1(n18488), .C2(n18278), .A(n18262), .B(n18261), .ZN(
        P3_U2917) );
  AOI22_X1 U21399 ( .A1(n18490), .A2(n18273), .B1(n18489), .B2(n18274), .ZN(
        n18264) );
  AOI22_X1 U21400 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18275), .B1(
        n18491), .B2(n18298), .ZN(n18263) );
  OAI211_X1 U21401 ( .C1(n18494), .C2(n18278), .A(n18264), .B(n18263), .ZN(
        P3_U2918) );
  AOI22_X1 U21402 ( .A1(n18497), .A2(n18274), .B1(n18495), .B2(n18273), .ZN(
        n18266) );
  AOI22_X1 U21403 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18275), .B1(
        n18496), .B2(n18298), .ZN(n18265) );
  OAI211_X1 U21404 ( .C1(n18500), .C2(n18278), .A(n18266), .B(n18265), .ZN(
        P3_U2919) );
  AOI22_X1 U21405 ( .A1(n18502), .A2(n18274), .B1(n18501), .B2(n18273), .ZN(
        n18268) );
  AOI22_X1 U21406 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18275), .B1(
        n18503), .B2(n18298), .ZN(n18267) );
  OAI211_X1 U21407 ( .C1(n18506), .C2(n18278), .A(n18268), .B(n18267), .ZN(
        P3_U2920) );
  AOI22_X1 U21408 ( .A1(n18508), .A2(n18274), .B1(n18507), .B2(n18273), .ZN(
        n18270) );
  AOI22_X1 U21409 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18275), .B1(
        n18509), .B2(n18298), .ZN(n18269) );
  OAI211_X1 U21410 ( .C1(n18512), .C2(n18278), .A(n18270), .B(n18269), .ZN(
        P3_U2921) );
  AOI22_X1 U21411 ( .A1(n18515), .A2(n18274), .B1(n18513), .B2(n18273), .ZN(
        n18272) );
  AOI22_X1 U21412 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18275), .B1(
        n18514), .B2(n18298), .ZN(n18271) );
  OAI211_X1 U21413 ( .C1(n18518), .C2(n18278), .A(n18272), .B(n18271), .ZN(
        P3_U2922) );
  AOI22_X1 U21414 ( .A1(n18523), .A2(n18298), .B1(n18520), .B2(n18273), .ZN(
        n18277) );
  AOI22_X1 U21415 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18275), .B1(
        n18522), .B2(n18274), .ZN(n18276) );
  OAI211_X1 U21416 ( .C1(n18528), .C2(n18278), .A(n18277), .B(n18276), .ZN(
        P3_U2923) );
  NOR2_X2 U21417 ( .A1(n18574), .A2(n18279), .ZN(n18366) );
  INV_X1 U21418 ( .A(n18366), .ZN(n18302) );
  NOR2_X1 U21419 ( .A1(n18280), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18327) );
  AND2_X1 U21420 ( .A1(n18472), .A2(n18327), .ZN(n18297) );
  AOI22_X1 U21421 ( .A1(n18479), .A2(n18298), .B1(n18473), .B2(n18297), .ZN(
        n18284) );
  NAND2_X1 U21422 ( .A1(n18282), .A2(n18281), .ZN(n18299) );
  AOI22_X1 U21423 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18299), .B1(
        n18474), .B2(n18320), .ZN(n18283) );
  OAI211_X1 U21424 ( .C1(n18482), .C2(n18302), .A(n18284), .B(n18283), .ZN(
        P3_U2924) );
  AOI22_X1 U21425 ( .A1(n18484), .A2(n18298), .B1(n18483), .B2(n18297), .ZN(
        n18286) );
  AOI22_X1 U21426 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18299), .B1(
        n18485), .B2(n18320), .ZN(n18285) );
  OAI211_X1 U21427 ( .C1(n18488), .C2(n18302), .A(n18286), .B(n18285), .ZN(
        P3_U2925) );
  AOI22_X1 U21428 ( .A1(n18490), .A2(n18297), .B1(n18489), .B2(n18298), .ZN(
        n18288) );
  AOI22_X1 U21429 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18299), .B1(
        n18491), .B2(n18320), .ZN(n18287) );
  OAI211_X1 U21430 ( .C1(n18494), .C2(n18302), .A(n18288), .B(n18287), .ZN(
        P3_U2926) );
  AOI22_X1 U21431 ( .A1(n18496), .A2(n18320), .B1(n18495), .B2(n18297), .ZN(
        n18290) );
  AOI22_X1 U21432 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18299), .B1(
        n18497), .B2(n18298), .ZN(n18289) );
  OAI211_X1 U21433 ( .C1(n18500), .C2(n18302), .A(n18290), .B(n18289), .ZN(
        P3_U2927) );
  AOI22_X1 U21434 ( .A1(n18503), .A2(n18320), .B1(n18501), .B2(n18297), .ZN(
        n18292) );
  AOI22_X1 U21435 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18299), .B1(
        n18502), .B2(n18298), .ZN(n18291) );
  OAI211_X1 U21436 ( .C1(n18506), .C2(n18302), .A(n18292), .B(n18291), .ZN(
        P3_U2928) );
  AOI22_X1 U21437 ( .A1(n18508), .A2(n18298), .B1(n18507), .B2(n18297), .ZN(
        n18294) );
  AOI22_X1 U21438 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18299), .B1(
        n18509), .B2(n18320), .ZN(n18293) );
  OAI211_X1 U21439 ( .C1(n18512), .C2(n18302), .A(n18294), .B(n18293), .ZN(
        P3_U2929) );
  AOI22_X1 U21440 ( .A1(n18514), .A2(n18320), .B1(n18513), .B2(n18297), .ZN(
        n18296) );
  AOI22_X1 U21441 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18299), .B1(
        n18515), .B2(n18298), .ZN(n18295) );
  OAI211_X1 U21442 ( .C1(n18518), .C2(n18302), .A(n18296), .B(n18295), .ZN(
        P3_U2930) );
  AOI22_X1 U21443 ( .A1(n18523), .A2(n18320), .B1(n18520), .B2(n18297), .ZN(
        n18301) );
  AOI22_X1 U21444 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18299), .B1(
        n18522), .B2(n18298), .ZN(n18300) );
  OAI211_X1 U21445 ( .C1(n18528), .C2(n18302), .A(n18301), .B(n18300), .ZN(
        P3_U2931) );
  NAND2_X1 U21446 ( .A1(n18394), .A2(n18371), .ZN(n18324) );
  INV_X1 U21447 ( .A(n18324), .ZN(n18388) );
  NOR2_X1 U21448 ( .A1(n18366), .A2(n18388), .ZN(n18349) );
  NOR2_X1 U21449 ( .A1(n18603), .A2(n18349), .ZN(n18319) );
  AOI22_X1 U21450 ( .A1(n18474), .A2(n18343), .B1(n18473), .B2(n18319), .ZN(
        n18306) );
  OAI21_X1 U21451 ( .B1(n18303), .B2(n18348), .A(n18349), .ZN(n18304) );
  OAI211_X1 U21452 ( .C1(n18388), .C2(n20828), .A(n18396), .B(n18304), .ZN(
        n18321) );
  AOI22_X1 U21453 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18321), .B1(
        n18479), .B2(n18320), .ZN(n18305) );
  OAI211_X1 U21454 ( .C1(n18482), .C2(n18324), .A(n18306), .B(n18305), .ZN(
        P3_U2932) );
  AOI22_X1 U21455 ( .A1(n18485), .A2(n18343), .B1(n18483), .B2(n18319), .ZN(
        n18308) );
  AOI22_X1 U21456 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18321), .B1(
        n18484), .B2(n18320), .ZN(n18307) );
  OAI211_X1 U21457 ( .C1(n18488), .C2(n18324), .A(n18308), .B(n18307), .ZN(
        P3_U2933) );
  AOI22_X1 U21458 ( .A1(n18490), .A2(n18319), .B1(n18489), .B2(n18320), .ZN(
        n18310) );
  AOI22_X1 U21459 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18321), .B1(
        n18491), .B2(n18343), .ZN(n18309) );
  OAI211_X1 U21460 ( .C1(n18494), .C2(n18324), .A(n18310), .B(n18309), .ZN(
        P3_U2934) );
  AOI22_X1 U21461 ( .A1(n18497), .A2(n18320), .B1(n18495), .B2(n18319), .ZN(
        n18312) );
  AOI22_X1 U21462 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18321), .B1(
        n18496), .B2(n18343), .ZN(n18311) );
  OAI211_X1 U21463 ( .C1(n18500), .C2(n18324), .A(n18312), .B(n18311), .ZN(
        P3_U2935) );
  AOI22_X1 U21464 ( .A1(n18502), .A2(n18320), .B1(n18501), .B2(n18319), .ZN(
        n18314) );
  AOI22_X1 U21465 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18321), .B1(
        n18503), .B2(n18343), .ZN(n18313) );
  OAI211_X1 U21466 ( .C1(n18506), .C2(n18324), .A(n18314), .B(n18313), .ZN(
        P3_U2936) );
  AOI22_X1 U21467 ( .A1(n18509), .A2(n18343), .B1(n18507), .B2(n18319), .ZN(
        n18316) );
  AOI22_X1 U21468 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18321), .B1(
        n18508), .B2(n18320), .ZN(n18315) );
  OAI211_X1 U21469 ( .C1(n18512), .C2(n18324), .A(n18316), .B(n18315), .ZN(
        P3_U2937) );
  AOI22_X1 U21470 ( .A1(n18515), .A2(n18320), .B1(n18513), .B2(n18319), .ZN(
        n18318) );
  AOI22_X1 U21471 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18321), .B1(
        n18514), .B2(n18343), .ZN(n18317) );
  OAI211_X1 U21472 ( .C1(n18518), .C2(n18324), .A(n18318), .B(n18317), .ZN(
        P3_U2938) );
  AOI22_X1 U21473 ( .A1(n18523), .A2(n18343), .B1(n18520), .B2(n18319), .ZN(
        n18323) );
  AOI22_X1 U21474 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18321), .B1(
        n18522), .B2(n18320), .ZN(n18322) );
  OAI211_X1 U21475 ( .C1(n18528), .C2(n18324), .A(n18323), .B(n18322), .ZN(
        P3_U2939) );
  NAND2_X1 U21476 ( .A1(n18325), .A2(n18371), .ZN(n18372) );
  INV_X1 U21477 ( .A(n18371), .ZN(n18370) );
  NOR2_X1 U21478 ( .A1(n18326), .A2(n18370), .ZN(n18342) );
  AOI22_X1 U21479 ( .A1(n18479), .A2(n18343), .B1(n18473), .B2(n18342), .ZN(
        n18329) );
  AOI22_X1 U21480 ( .A1(n18478), .A2(n18327), .B1(n18418), .B2(n18371), .ZN(
        n18344) );
  AOI22_X1 U21481 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18344), .B1(
        n18474), .B2(n18366), .ZN(n18328) );
  OAI211_X1 U21482 ( .C1(n18482), .C2(n18372), .A(n18329), .B(n18328), .ZN(
        P3_U2940) );
  AOI22_X1 U21483 ( .A1(n18485), .A2(n18366), .B1(n18483), .B2(n18342), .ZN(
        n18331) );
  AOI22_X1 U21484 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18344), .B1(
        n18484), .B2(n18343), .ZN(n18330) );
  OAI211_X1 U21485 ( .C1(n18488), .C2(n18372), .A(n18331), .B(n18330), .ZN(
        P3_U2941) );
  AOI22_X1 U21486 ( .A1(n18491), .A2(n18366), .B1(n18490), .B2(n18342), .ZN(
        n18333) );
  AOI22_X1 U21487 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18344), .B1(
        n18489), .B2(n18343), .ZN(n18332) );
  OAI211_X1 U21488 ( .C1(n18494), .C2(n18372), .A(n18333), .B(n18332), .ZN(
        P3_U2942) );
  AOI22_X1 U21489 ( .A1(n18497), .A2(n18343), .B1(n18495), .B2(n18342), .ZN(
        n18335) );
  AOI22_X1 U21490 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18344), .B1(
        n18496), .B2(n18366), .ZN(n18334) );
  OAI211_X1 U21491 ( .C1(n18500), .C2(n18372), .A(n18335), .B(n18334), .ZN(
        P3_U2943) );
  AOI22_X1 U21492 ( .A1(n18502), .A2(n18343), .B1(n18501), .B2(n18342), .ZN(
        n18337) );
  AOI22_X1 U21493 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18344), .B1(
        n18503), .B2(n18366), .ZN(n18336) );
  OAI211_X1 U21494 ( .C1(n18506), .C2(n18372), .A(n18337), .B(n18336), .ZN(
        P3_U2944) );
  AOI22_X1 U21495 ( .A1(n18508), .A2(n18343), .B1(n18507), .B2(n18342), .ZN(
        n18339) );
  AOI22_X1 U21496 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18344), .B1(
        n18509), .B2(n18366), .ZN(n18338) );
  OAI211_X1 U21497 ( .C1(n18512), .C2(n18372), .A(n18339), .B(n18338), .ZN(
        P3_U2945) );
  AOI22_X1 U21498 ( .A1(n18514), .A2(n18366), .B1(n18513), .B2(n18342), .ZN(
        n18341) );
  AOI22_X1 U21499 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18344), .B1(
        n18515), .B2(n18343), .ZN(n18340) );
  OAI211_X1 U21500 ( .C1(n18518), .C2(n18372), .A(n18341), .B(n18340), .ZN(
        P3_U2946) );
  AOI22_X1 U21501 ( .A1(n18523), .A2(n18366), .B1(n18520), .B2(n18342), .ZN(
        n18346) );
  AOI22_X1 U21502 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18344), .B1(
        n18522), .B2(n18343), .ZN(n18345) );
  OAI211_X1 U21503 ( .C1(n18528), .C2(n18372), .A(n18346), .B(n18345), .ZN(
        P3_U2947) );
  NOR2_X1 U21504 ( .A1(n18575), .A2(n18370), .ZN(n18420) );
  NAND2_X1 U21505 ( .A1(n18420), .A2(n18392), .ZN(n18393) );
  AOI21_X1 U21506 ( .B1(n18372), .B2(n18393), .A(n18603), .ZN(n18365) );
  AOI22_X1 U21507 ( .A1(n18479), .A2(n18366), .B1(n18473), .B2(n18365), .ZN(
        n18352) );
  INV_X1 U21508 ( .A(n18347), .ZN(n18443) );
  OAI211_X1 U21509 ( .C1(n18349), .C2(n18348), .A(n18372), .B(n18393), .ZN(
        n18350) );
  NAND2_X1 U21510 ( .A1(n18443), .A2(n18350), .ZN(n18367) );
  AOI22_X1 U21511 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18367), .B1(
        n18474), .B2(n18388), .ZN(n18351) );
  OAI211_X1 U21512 ( .C1(n18482), .C2(n18393), .A(n18352), .B(n18351), .ZN(
        P3_U2948) );
  AOI22_X1 U21513 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18367), .B1(
        n18483), .B2(n18365), .ZN(n18354) );
  AOI22_X1 U21514 ( .A1(n18484), .A2(n18366), .B1(n18485), .B2(n18388), .ZN(
        n18353) );
  OAI211_X1 U21515 ( .C1(n18488), .C2(n18393), .A(n18354), .B(n18353), .ZN(
        P3_U2949) );
  AOI22_X1 U21516 ( .A1(n18490), .A2(n18365), .B1(n18489), .B2(n18366), .ZN(
        n18356) );
  AOI22_X1 U21517 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18367), .B1(
        n18491), .B2(n18388), .ZN(n18355) );
  OAI211_X1 U21518 ( .C1(n18494), .C2(n18393), .A(n18356), .B(n18355), .ZN(
        P3_U2950) );
  AOI22_X1 U21519 ( .A1(n18497), .A2(n18366), .B1(n18495), .B2(n18365), .ZN(
        n18358) );
  AOI22_X1 U21520 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18367), .B1(
        n18496), .B2(n18388), .ZN(n18357) );
  OAI211_X1 U21521 ( .C1(n18500), .C2(n18393), .A(n18358), .B(n18357), .ZN(
        P3_U2951) );
  AOI22_X1 U21522 ( .A1(n18502), .A2(n18366), .B1(n18501), .B2(n18365), .ZN(
        n18360) );
  AOI22_X1 U21523 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18367), .B1(
        n18503), .B2(n18388), .ZN(n18359) );
  OAI211_X1 U21524 ( .C1(n18506), .C2(n18393), .A(n18360), .B(n18359), .ZN(
        P3_U2952) );
  AOI22_X1 U21525 ( .A1(n18508), .A2(n18366), .B1(n18507), .B2(n18365), .ZN(
        n18362) );
  AOI22_X1 U21526 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18367), .B1(
        n18509), .B2(n18388), .ZN(n18361) );
  OAI211_X1 U21527 ( .C1(n18512), .C2(n18393), .A(n18362), .B(n18361), .ZN(
        P3_U2953) );
  AOI22_X1 U21528 ( .A1(n18514), .A2(n18388), .B1(n18513), .B2(n18365), .ZN(
        n18364) );
  AOI22_X1 U21529 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18367), .B1(
        n18515), .B2(n18366), .ZN(n18363) );
  OAI211_X1 U21530 ( .C1(n18518), .C2(n18393), .A(n18364), .B(n18363), .ZN(
        P3_U2954) );
  AOI22_X1 U21531 ( .A1(n18523), .A2(n18388), .B1(n18520), .B2(n18365), .ZN(
        n18369) );
  AOI22_X1 U21532 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18367), .B1(
        n18522), .B2(n18366), .ZN(n18368) );
  OAI211_X1 U21533 ( .C1(n18528), .C2(n18393), .A(n18369), .B(n18368), .ZN(
        P3_U2955) );
  NOR2_X2 U21534 ( .A1(n18574), .A2(n18370), .ZN(n18466) );
  INV_X1 U21535 ( .A(n18466), .ZN(n18442) );
  AND2_X1 U21536 ( .A1(n18472), .A2(n18420), .ZN(n18387) );
  AOI22_X1 U21537 ( .A1(n18479), .A2(n18388), .B1(n18473), .B2(n18387), .ZN(
        n18374) );
  AOI22_X1 U21538 ( .A1(n18478), .A2(n18371), .B1(n18475), .B2(n18420), .ZN(
        n18389) );
  INV_X1 U21539 ( .A(n18372), .ZN(n18413) );
  AOI22_X1 U21540 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18389), .B1(
        n18474), .B2(n18413), .ZN(n18373) );
  OAI211_X1 U21541 ( .C1(n18482), .C2(n18442), .A(n18374), .B(n18373), .ZN(
        P3_U2956) );
  AOI22_X1 U21542 ( .A1(n18485), .A2(n18413), .B1(n18483), .B2(n18387), .ZN(
        n18376) );
  AOI22_X1 U21543 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18389), .B1(
        n18484), .B2(n18388), .ZN(n18375) );
  OAI211_X1 U21544 ( .C1(n18488), .C2(n18442), .A(n18376), .B(n18375), .ZN(
        P3_U2957) );
  AOI22_X1 U21545 ( .A1(n18491), .A2(n18413), .B1(n18490), .B2(n18387), .ZN(
        n18378) );
  AOI22_X1 U21546 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18389), .B1(
        n18489), .B2(n18388), .ZN(n18377) );
  OAI211_X1 U21547 ( .C1(n18494), .C2(n18442), .A(n18378), .B(n18377), .ZN(
        P3_U2958) );
  AOI22_X1 U21548 ( .A1(n18497), .A2(n18388), .B1(n18495), .B2(n18387), .ZN(
        n18380) );
  AOI22_X1 U21549 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18389), .B1(
        n18496), .B2(n18413), .ZN(n18379) );
  OAI211_X1 U21550 ( .C1(n18500), .C2(n18442), .A(n18380), .B(n18379), .ZN(
        P3_U2959) );
  AOI22_X1 U21551 ( .A1(n18502), .A2(n18388), .B1(n18501), .B2(n18387), .ZN(
        n18382) );
  AOI22_X1 U21552 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18389), .B1(
        n18503), .B2(n18413), .ZN(n18381) );
  OAI211_X1 U21553 ( .C1(n18506), .C2(n18442), .A(n18382), .B(n18381), .ZN(
        P3_U2960) );
  AOI22_X1 U21554 ( .A1(n18509), .A2(n18413), .B1(n18507), .B2(n18387), .ZN(
        n18384) );
  AOI22_X1 U21555 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18389), .B1(
        n18508), .B2(n18388), .ZN(n18383) );
  OAI211_X1 U21556 ( .C1(n18512), .C2(n18442), .A(n18384), .B(n18383), .ZN(
        P3_U2961) );
  AOI22_X1 U21557 ( .A1(n18515), .A2(n18388), .B1(n18513), .B2(n18387), .ZN(
        n18386) );
  AOI22_X1 U21558 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18389), .B1(
        n18514), .B2(n18413), .ZN(n18385) );
  OAI211_X1 U21559 ( .C1(n18518), .C2(n18442), .A(n18386), .B(n18385), .ZN(
        P3_U2962) );
  AOI22_X1 U21560 ( .A1(n18523), .A2(n18413), .B1(n18520), .B2(n18387), .ZN(
        n18391) );
  AOI22_X1 U21561 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18389), .B1(
        n18522), .B2(n18388), .ZN(n18390) );
  OAI211_X1 U21562 ( .C1(n18528), .C2(n18442), .A(n18391), .B(n18390), .ZN(
        P3_U2963) );
  INV_X1 U21563 ( .A(n18417), .ZN(n18477) );
  NAND2_X1 U21564 ( .A1(n18477), .A2(n18392), .ZN(n18451) );
  INV_X1 U21565 ( .A(n18393), .ZN(n18436) );
  AOI21_X1 U21566 ( .B1(n18442), .B2(n18451), .A(n18603), .ZN(n18412) );
  AOI22_X1 U21567 ( .A1(n18474), .A2(n18436), .B1(n18473), .B2(n18412), .ZN(
        n18399) );
  INV_X1 U21568 ( .A(n18451), .ZN(n18521) );
  AOI211_X1 U21569 ( .C1(n18442), .C2(n18395), .A(P3_STATE2_REG_3__SCAN_IN), 
        .B(n18394), .ZN(n18397) );
  OAI21_X1 U21570 ( .B1(n18521), .B2(n18397), .A(n18396), .ZN(n18414) );
  AOI22_X1 U21571 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18414), .B1(
        n18479), .B2(n18413), .ZN(n18398) );
  OAI211_X1 U21572 ( .C1(n18482), .C2(n18451), .A(n18399), .B(n18398), .ZN(
        P3_U2964) );
  AOI22_X1 U21573 ( .A1(n18485), .A2(n18436), .B1(n18483), .B2(n18412), .ZN(
        n18401) );
  AOI22_X1 U21574 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18414), .B1(
        n18484), .B2(n18413), .ZN(n18400) );
  OAI211_X1 U21575 ( .C1(n18488), .C2(n18451), .A(n18401), .B(n18400), .ZN(
        P3_U2965) );
  AOI22_X1 U21576 ( .A1(n18490), .A2(n18412), .B1(n18489), .B2(n18413), .ZN(
        n18403) );
  AOI22_X1 U21577 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18414), .B1(
        n18491), .B2(n18436), .ZN(n18402) );
  OAI211_X1 U21578 ( .C1(n18494), .C2(n18451), .A(n18403), .B(n18402), .ZN(
        P3_U2966) );
  AOI22_X1 U21579 ( .A1(n18496), .A2(n18436), .B1(n18495), .B2(n18412), .ZN(
        n18405) );
  AOI22_X1 U21580 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18414), .B1(
        n18497), .B2(n18413), .ZN(n18404) );
  OAI211_X1 U21581 ( .C1(n18500), .C2(n18451), .A(n18405), .B(n18404), .ZN(
        P3_U2967) );
  AOI22_X1 U21582 ( .A1(n18502), .A2(n18413), .B1(n18501), .B2(n18412), .ZN(
        n18407) );
  AOI22_X1 U21583 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18414), .B1(
        n18503), .B2(n18436), .ZN(n18406) );
  OAI211_X1 U21584 ( .C1(n18506), .C2(n18451), .A(n18407), .B(n18406), .ZN(
        P3_U2968) );
  AOI22_X1 U21585 ( .A1(n18508), .A2(n18413), .B1(n18507), .B2(n18412), .ZN(
        n18409) );
  AOI22_X1 U21586 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18414), .B1(
        n18509), .B2(n18436), .ZN(n18408) );
  OAI211_X1 U21587 ( .C1(n18512), .C2(n18451), .A(n18409), .B(n18408), .ZN(
        P3_U2969) );
  AOI22_X1 U21588 ( .A1(n18515), .A2(n18413), .B1(n18513), .B2(n18412), .ZN(
        n18411) );
  AOI22_X1 U21589 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18414), .B1(
        n18514), .B2(n18436), .ZN(n18410) );
  OAI211_X1 U21590 ( .C1(n18518), .C2(n18451), .A(n18411), .B(n18410), .ZN(
        P3_U2970) );
  AOI22_X1 U21591 ( .A1(n18522), .A2(n18413), .B1(n18520), .B2(n18412), .ZN(
        n18416) );
  AOI22_X1 U21592 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18414), .B1(
        n18523), .B2(n18436), .ZN(n18415) );
  OAI211_X1 U21593 ( .C1(n18528), .C2(n18451), .A(n18416), .B(n18415), .ZN(
        P3_U2971) );
  NOR2_X1 U21594 ( .A1(n18603), .A2(n18417), .ZN(n18435) );
  AOI22_X1 U21595 ( .A1(n18479), .A2(n18436), .B1(n18473), .B2(n18435), .ZN(
        n18422) );
  AOI22_X1 U21596 ( .A1(n18478), .A2(n18420), .B1(n18419), .B2(n18418), .ZN(
        n18437) );
  AOI22_X1 U21597 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18437), .B1(
        n18524), .B2(n18447), .ZN(n18421) );
  OAI211_X1 U21598 ( .C1(n18452), .C2(n18442), .A(n18422), .B(n18421), .ZN(
        P3_U2972) );
  INV_X1 U21599 ( .A(n18524), .ZN(n18440) );
  AOI22_X1 U21600 ( .A1(n18485), .A2(n18466), .B1(n18483), .B2(n18435), .ZN(
        n18424) );
  AOI22_X1 U21601 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18437), .B1(
        n18484), .B2(n18436), .ZN(n18423) );
  OAI211_X1 U21602 ( .C1(n18440), .C2(n18488), .A(n18424), .B(n18423), .ZN(
        P3_U2973) );
  AOI22_X1 U21603 ( .A1(n18491), .A2(n18466), .B1(n18490), .B2(n18435), .ZN(
        n18426) );
  AOI22_X1 U21604 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18437), .B1(
        n18489), .B2(n18436), .ZN(n18425) );
  OAI211_X1 U21605 ( .C1(n18440), .C2(n18494), .A(n18426), .B(n18425), .ZN(
        P3_U2974) );
  AOI22_X1 U21606 ( .A1(n18496), .A2(n18466), .B1(n18495), .B2(n18435), .ZN(
        n18428) );
  AOI22_X1 U21607 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18437), .B1(
        n18497), .B2(n18436), .ZN(n18427) );
  OAI211_X1 U21608 ( .C1(n18440), .C2(n18500), .A(n18428), .B(n18427), .ZN(
        P3_U2975) );
  AOI22_X1 U21609 ( .A1(n18503), .A2(n18466), .B1(n18501), .B2(n18435), .ZN(
        n18430) );
  AOI22_X1 U21610 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18437), .B1(
        n18502), .B2(n18436), .ZN(n18429) );
  OAI211_X1 U21611 ( .C1(n18440), .C2(n18506), .A(n18430), .B(n18429), .ZN(
        P3_U2976) );
  AOI22_X1 U21612 ( .A1(n18508), .A2(n18436), .B1(n18507), .B2(n18435), .ZN(
        n18432) );
  AOI22_X1 U21613 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18437), .B1(
        n18509), .B2(n18466), .ZN(n18431) );
  OAI211_X1 U21614 ( .C1(n18440), .C2(n18512), .A(n18432), .B(n18431), .ZN(
        P3_U2977) );
  AOI22_X1 U21615 ( .A1(n18515), .A2(n18436), .B1(n18513), .B2(n18435), .ZN(
        n18434) );
  AOI22_X1 U21616 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18437), .B1(
        n18514), .B2(n18466), .ZN(n18433) );
  OAI211_X1 U21617 ( .C1(n18440), .C2(n18518), .A(n18434), .B(n18433), .ZN(
        P3_U2978) );
  AOI22_X1 U21618 ( .A1(n18522), .A2(n18436), .B1(n18520), .B2(n18435), .ZN(
        n18439) );
  AOI22_X1 U21619 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18437), .B1(
        n18523), .B2(n18466), .ZN(n18438) );
  OAI211_X1 U21620 ( .C1(n18440), .C2(n18528), .A(n18439), .B(n18438), .ZN(
        P3_U2979) );
  NOR2_X1 U21621 ( .A1(n18603), .A2(n18441), .ZN(n18465) );
  AOI22_X1 U21622 ( .A1(n18479), .A2(n18466), .B1(n18473), .B2(n18465), .ZN(
        n18450) );
  INV_X1 U21623 ( .A(n18441), .ZN(n18446) );
  NAND2_X1 U21624 ( .A1(n18442), .A2(n18451), .ZN(n18444) );
  OAI221_X1 U21625 ( .B1(n18446), .B2(n18445), .C1(n18446), .C2(n18444), .A(
        n18443), .ZN(n18467) );
  AOI22_X1 U21626 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18467), .B1(
        n18448), .B2(n18447), .ZN(n18449) );
  OAI211_X1 U21627 ( .C1(n18452), .C2(n18451), .A(n18450), .B(n18449), .ZN(
        P3_U2980) );
  AOI22_X1 U21628 ( .A1(n18484), .A2(n18466), .B1(n18483), .B2(n18465), .ZN(
        n18454) );
  AOI22_X1 U21629 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18467), .B1(
        n18485), .B2(n18521), .ZN(n18453) );
  OAI211_X1 U21630 ( .C1(n18470), .C2(n18488), .A(n18454), .B(n18453), .ZN(
        P3_U2981) );
  AOI22_X1 U21631 ( .A1(n18491), .A2(n18521), .B1(n18490), .B2(n18465), .ZN(
        n18456) );
  AOI22_X1 U21632 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18467), .B1(
        n18489), .B2(n18466), .ZN(n18455) );
  OAI211_X1 U21633 ( .C1(n18470), .C2(n18494), .A(n18456), .B(n18455), .ZN(
        P3_U2982) );
  AOI22_X1 U21634 ( .A1(n18496), .A2(n18521), .B1(n18495), .B2(n18465), .ZN(
        n18458) );
  AOI22_X1 U21635 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18467), .B1(
        n18497), .B2(n18466), .ZN(n18457) );
  OAI211_X1 U21636 ( .C1(n18470), .C2(n18500), .A(n18458), .B(n18457), .ZN(
        P3_U2983) );
  AOI22_X1 U21637 ( .A1(n18502), .A2(n18466), .B1(n18501), .B2(n18465), .ZN(
        n18460) );
  AOI22_X1 U21638 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18467), .B1(
        n18503), .B2(n18521), .ZN(n18459) );
  OAI211_X1 U21639 ( .C1(n18470), .C2(n18506), .A(n18460), .B(n18459), .ZN(
        P3_U2984) );
  AOI22_X1 U21640 ( .A1(n18508), .A2(n18466), .B1(n18507), .B2(n18465), .ZN(
        n18462) );
  AOI22_X1 U21641 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18467), .B1(
        n18509), .B2(n18521), .ZN(n18461) );
  OAI211_X1 U21642 ( .C1(n18470), .C2(n18512), .A(n18462), .B(n18461), .ZN(
        P3_U2985) );
  AOI22_X1 U21643 ( .A1(n18515), .A2(n18466), .B1(n18513), .B2(n18465), .ZN(
        n18464) );
  AOI22_X1 U21644 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18467), .B1(
        n18514), .B2(n18521), .ZN(n18463) );
  OAI211_X1 U21645 ( .C1(n18470), .C2(n18518), .A(n18464), .B(n18463), .ZN(
        P3_U2986) );
  AOI22_X1 U21646 ( .A1(n18522), .A2(n18466), .B1(n18520), .B2(n18465), .ZN(
        n18469) );
  AOI22_X1 U21647 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18467), .B1(
        n18523), .B2(n18521), .ZN(n18468) );
  OAI211_X1 U21648 ( .C1(n18470), .C2(n18528), .A(n18469), .B(n18468), .ZN(
        P3_U2987) );
  INV_X1 U21649 ( .A(n18471), .ZN(n18529) );
  AND2_X1 U21650 ( .A1(n18472), .A2(n18476), .ZN(n18519) );
  AOI22_X1 U21651 ( .A1(n18474), .A2(n18524), .B1(n18473), .B2(n18519), .ZN(
        n18481) );
  AOI22_X1 U21652 ( .A1(n18478), .A2(n18477), .B1(n18476), .B2(n18475), .ZN(
        n18525) );
  AOI22_X1 U21653 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18525), .B1(
        n18479), .B2(n18521), .ZN(n18480) );
  OAI211_X1 U21654 ( .C1(n18529), .C2(n18482), .A(n18481), .B(n18480), .ZN(
        P3_U2988) );
  AOI22_X1 U21655 ( .A1(n18484), .A2(n18521), .B1(n18483), .B2(n18519), .ZN(
        n18487) );
  AOI22_X1 U21656 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18525), .B1(
        n18524), .B2(n18485), .ZN(n18486) );
  OAI211_X1 U21657 ( .C1(n18529), .C2(n18488), .A(n18487), .B(n18486), .ZN(
        P3_U2989) );
  AOI22_X1 U21658 ( .A1(n18490), .A2(n18519), .B1(n18489), .B2(n18521), .ZN(
        n18493) );
  AOI22_X1 U21659 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18525), .B1(
        n18524), .B2(n18491), .ZN(n18492) );
  OAI211_X1 U21660 ( .C1(n18529), .C2(n18494), .A(n18493), .B(n18492), .ZN(
        P3_U2990) );
  AOI22_X1 U21661 ( .A1(n18524), .A2(n18496), .B1(n18495), .B2(n18519), .ZN(
        n18499) );
  AOI22_X1 U21662 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18525), .B1(
        n18497), .B2(n18521), .ZN(n18498) );
  OAI211_X1 U21663 ( .C1(n18529), .C2(n18500), .A(n18499), .B(n18498), .ZN(
        P3_U2991) );
  AOI22_X1 U21664 ( .A1(n18502), .A2(n18521), .B1(n18501), .B2(n18519), .ZN(
        n18505) );
  AOI22_X1 U21665 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18525), .B1(
        n18524), .B2(n18503), .ZN(n18504) );
  OAI211_X1 U21666 ( .C1(n18529), .C2(n18506), .A(n18505), .B(n18504), .ZN(
        P3_U2992) );
  AOI22_X1 U21667 ( .A1(n18508), .A2(n18521), .B1(n18507), .B2(n18519), .ZN(
        n18511) );
  AOI22_X1 U21668 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18525), .B1(
        n18524), .B2(n18509), .ZN(n18510) );
  OAI211_X1 U21669 ( .C1(n18529), .C2(n18512), .A(n18511), .B(n18510), .ZN(
        P3_U2993) );
  AOI22_X1 U21670 ( .A1(n18524), .A2(n18514), .B1(n18513), .B2(n18519), .ZN(
        n18517) );
  AOI22_X1 U21671 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18525), .B1(
        n18515), .B2(n18521), .ZN(n18516) );
  OAI211_X1 U21672 ( .C1(n18529), .C2(n18518), .A(n18517), .B(n18516), .ZN(
        P3_U2994) );
  AOI22_X1 U21673 ( .A1(n18522), .A2(n18521), .B1(n18520), .B2(n18519), .ZN(
        n18527) );
  AOI22_X1 U21674 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18525), .B1(
        n18524), .B2(n18523), .ZN(n18526) );
  OAI211_X1 U21675 ( .C1(n18529), .C2(n18528), .A(n18527), .B(n18526), .ZN(
        P3_U2995) );
  NOR2_X1 U21676 ( .A1(n18566), .A2(n18530), .ZN(n18532) );
  OAI222_X1 U21677 ( .A1(n18536), .A2(n18535), .B1(n18534), .B2(n18533), .C1(
        n18532), .C2(n18531), .ZN(n18742) );
  OAI21_X1 U21678 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18537), .ZN(n18538) );
  OAI211_X1 U21679 ( .C1(n18540), .C2(n18567), .A(n18539), .B(n18538), .ZN(
        n18589) );
  INV_X1 U21680 ( .A(n18567), .ZN(n18578) );
  AOI22_X1 U21681 ( .A1(n18544), .A2(n18543), .B1(n18542), .B2(n18541), .ZN(
        n18545) );
  INV_X1 U21682 ( .A(n18545), .ZN(n18547) );
  NOR2_X1 U21683 ( .A1(n18546), .A2(n18547), .ZN(n18563) );
  INV_X1 U21684 ( .A(n18563), .ZN(n18551) );
  OR3_X1 U21685 ( .A1(n18554), .A2(n18548), .A3(n18547), .ZN(n18549) );
  AOI22_X1 U21686 ( .A1(n20898), .A2(n18551), .B1(n18550), .B2(n18549), .ZN(
        n18557) );
  NOR2_X1 U21687 ( .A1(n9610), .A2(n18717), .ZN(n18553) );
  OAI21_X1 U21688 ( .B1(n18552), .B2(n20898), .A(n18570), .ZN(n18558) );
  AOI22_X1 U21689 ( .A1(n18566), .A2(n18556), .B1(n18553), .B2(n18558), .ZN(
        n18555) );
  AOI22_X1 U21690 ( .A1(n18557), .A2(n18556), .B1(n18555), .B2(n18554), .ZN(
        n18706) );
  AOI22_X1 U21691 ( .A1(n18578), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n18706), .B2(n18567), .ZN(n18587) );
  INV_X1 U21692 ( .A(n18558), .ZN(n18571) );
  NOR3_X1 U21693 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18571), .A3(
        n9610), .ZN(n18565) );
  NAND2_X1 U21694 ( .A1(n9610), .A2(n18559), .ZN(n18562) );
  INV_X1 U21695 ( .A(n18560), .ZN(n18561) );
  AOI211_X1 U21696 ( .C1(n18563), .C2(n18562), .A(n18561), .B(n18717), .ZN(
        n18564) );
  AOI211_X1 U21697 ( .C1(n18566), .C2(n18711), .A(n18565), .B(n18564), .ZN(
        n18714) );
  AOI22_X1 U21698 ( .A1(n18578), .A2(n18717), .B1(n18714), .B2(n18567), .ZN(
        n18582) );
  NOR2_X1 U21699 ( .A1(n18569), .A2(n18568), .ZN(n18573) );
  AOI22_X1 U21700 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18570), .B1(
        n18573), .B2(n20898), .ZN(n18726) );
  OAI22_X1 U21701 ( .A1(n18573), .A2(n18572), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18571), .ZN(n18722) );
  AOI222_X1 U21702 ( .A1(n18726), .A2(n18722), .B1(n18726), .B2(n18575), .C1(
        n18722), .C2(n18574), .ZN(n18577) );
  OAI21_X1 U21703 ( .B1(n18578), .B2(n18577), .A(n18576), .ZN(n18581) );
  AND2_X1 U21704 ( .A1(n18582), .A2(n18581), .ZN(n18579) );
  OAI221_X1 U21705 ( .B1(n18582), .B2(n18581), .C1(n18580), .C2(n18579), .A(
        n18584), .ZN(n18586) );
  AOI21_X1 U21706 ( .B1(n18584), .B2(n18583), .A(n18582), .ZN(n18585) );
  AOI222_X1 U21707 ( .A1(n18587), .A2(n18586), .B1(n18587), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18586), .C2(n18585), .ZN(
        n18588) );
  NOR4_X1 U21708 ( .A1(n18590), .A2(n18742), .A3(n18589), .A4(n18588), .ZN(
        n18601) );
  AOI22_X1 U21709 ( .A1(n18725), .A2(n18754), .B1(n18602), .B2(n18747), .ZN(
        n18591) );
  INV_X1 U21710 ( .A(n18591), .ZN(n18597) );
  NAND3_X1 U21711 ( .A1(n18750), .A2(n18593), .A3(n18592), .ZN(n18594) );
  NAND3_X1 U21712 ( .A1(n18601), .A2(n18745), .A3(n18594), .ZN(n18704) );
  OAI21_X1 U21713 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18751), .A(n18704), 
        .ZN(n18604) );
  NOR2_X1 U21714 ( .A1(n18595), .A2(n18604), .ZN(n18596) );
  MUX2_X1 U21715 ( .A(n18597), .B(n18596), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18599) );
  OAI211_X1 U21716 ( .C1(n18601), .C2(n18600), .A(n18599), .B(n18598), .ZN(
        P3_U2996) );
  NAND2_X1 U21717 ( .A1(n18602), .A2(n18747), .ZN(n18607) );
  NAND4_X1 U21718 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n18602), .A4(n18762), .ZN(n18610) );
  OR3_X1 U21719 ( .A1(n18605), .A2(n18604), .A3(n18603), .ZN(n18606) );
  NAND4_X1 U21720 ( .A1(n18608), .A2(n18607), .A3(n18610), .A4(n18606), .ZN(
        P3_U2997) );
  OAI21_X1 U21721 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18609), .ZN(n18612) );
  INV_X1 U21722 ( .A(n18610), .ZN(n18611) );
  AOI21_X1 U21723 ( .B1(n18613), .B2(n18612), .A(n18611), .ZN(P3_U2998) );
  AND2_X1 U21724 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18614), .ZN(
        P3_U2999) );
  AND2_X1 U21725 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18614), .ZN(
        P3_U3000) );
  AND2_X1 U21726 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18614), .ZN(
        P3_U3001) );
  INV_X1 U21727 ( .A(P3_DATAWIDTH_REG_28__SCAN_IN), .ZN(n20800) );
  NOR2_X1 U21728 ( .A1(n20800), .A2(n18702), .ZN(P3_U3002) );
  AND2_X1 U21729 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18614), .ZN(
        P3_U3003) );
  AND2_X1 U21730 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18614), .ZN(
        P3_U3004) );
  AND2_X1 U21731 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18614), .ZN(
        P3_U3005) );
  AND2_X1 U21732 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18614), .ZN(
        P3_U3006) );
  AND2_X1 U21733 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18614), .ZN(
        P3_U3007) );
  AND2_X1 U21734 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18614), .ZN(
        P3_U3008) );
  AND2_X1 U21735 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18614), .ZN(
        P3_U3009) );
  AND2_X1 U21736 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18615), .ZN(
        P3_U3010) );
  AND2_X1 U21737 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18615), .ZN(
        P3_U3011) );
  AND2_X1 U21738 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18615), .ZN(
        P3_U3012) );
  AND2_X1 U21739 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18615), .ZN(
        P3_U3013) );
  AND2_X1 U21740 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18615), .ZN(
        P3_U3014) );
  AND2_X1 U21741 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18615), .ZN(
        P3_U3015) );
  AND2_X1 U21742 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18615), .ZN(
        P3_U3016) );
  AND2_X1 U21743 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18615), .ZN(
        P3_U3017) );
  AND2_X1 U21744 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18615), .ZN(
        P3_U3018) );
  AND2_X1 U21745 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18615), .ZN(
        P3_U3019) );
  AND2_X1 U21746 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18615), .ZN(
        P3_U3020) );
  AND2_X1 U21747 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18615), .ZN(P3_U3021) );
  AND2_X1 U21748 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18615), .ZN(P3_U3022) );
  AND2_X1 U21749 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18615), .ZN(P3_U3023) );
  AND2_X1 U21750 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18615), .ZN(P3_U3024) );
  AND2_X1 U21751 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18615), .ZN(P3_U3025) );
  AND2_X1 U21752 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18615), .ZN(P3_U3026) );
  AND2_X1 U21753 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18615), .ZN(P3_U3027) );
  AND2_X1 U21754 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18615), .ZN(P3_U3028) );
  NOR2_X1 U21755 ( .A1(n18751), .A2(n18618), .ZN(n18623) );
  OAI21_X1 U21756 ( .B1(n18616), .B2(n20668), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18617) );
  AOI22_X1 U21757 ( .A1(n18623), .A2(n18631), .B1(n18759), .B2(n18617), .ZN(
        n18619) );
  NAND3_X1 U21758 ( .A1(NA), .A2(n18629), .A3(n18618), .ZN(n18624) );
  OAI211_X1 U21759 ( .C1(P3_STATE_REG_0__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18619), .B(n18624), .ZN(P3_U3029) );
  NOR2_X1 U21760 ( .A1(n18631), .A2(n20668), .ZN(n18627) );
  INV_X1 U21761 ( .A(n18627), .ZN(n18621) );
  AOI22_X1 U21762 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(n18621), .B1(HOLD), 
        .B2(n18620), .ZN(n18622) );
  INV_X1 U21763 ( .A(n18623), .ZN(n18625) );
  OAI211_X1 U21764 ( .C1(n18622), .C2(n18629), .A(n18625), .B(n18748), .ZN(
        P3_U3030) );
  AOI21_X1 U21765 ( .B1(n18629), .B2(n18624), .A(n18623), .ZN(n18630) );
  OAI22_X1 U21766 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18625), .ZN(n18626) );
  OAI22_X1 U21767 ( .A1(n18627), .A2(n18626), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18628) );
  OAI22_X1 U21768 ( .A1(n18630), .A2(n18631), .B1(n18629), .B2(n18628), .ZN(
        P3_U3031) );
  OAI222_X1 U21769 ( .A1(n18633), .A2(n18691), .B1(n18632), .B2(n18697), .C1(
        n18634), .C2(n18687), .ZN(P3_U3032) );
  OAI222_X1 U21770 ( .A1(n18687), .A2(n18636), .B1(n18635), .B2(n18697), .C1(
        n18634), .C2(n18691), .ZN(P3_U3033) );
  INV_X1 U21771 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18638) );
  OAI222_X1 U21772 ( .A1(n18687), .A2(n18638), .B1(n18637), .B2(n18697), .C1(
        n18636), .C2(n18691), .ZN(P3_U3034) );
  OAI222_X1 U21773 ( .A1(n18687), .A2(n18641), .B1(n18639), .B2(n18697), .C1(
        n18638), .C2(n18691), .ZN(P3_U3035) );
  OAI222_X1 U21774 ( .A1(n18641), .A2(n18691), .B1(n18640), .B2(n18697), .C1(
        n18642), .C2(n18687), .ZN(P3_U3036) );
  OAI222_X1 U21775 ( .A1(n18687), .A2(n18644), .B1(n18643), .B2(n18697), .C1(
        n18642), .C2(n18691), .ZN(P3_U3037) );
  OAI222_X1 U21776 ( .A1(n18687), .A2(n18647), .B1(n18645), .B2(n18697), .C1(
        n18644), .C2(n18691), .ZN(P3_U3038) );
  OAI222_X1 U21777 ( .A1(n18647), .A2(n18691), .B1(n18646), .B2(n18697), .C1(
        n18648), .C2(n18687), .ZN(P3_U3039) );
  OAI222_X1 U21778 ( .A1(n18687), .A2(n18650), .B1(n18649), .B2(n18697), .C1(
        n18648), .C2(n18691), .ZN(P3_U3040) );
  OAI222_X1 U21779 ( .A1(n18687), .A2(n18652), .B1(n18651), .B2(n18697), .C1(
        n18650), .C2(n18691), .ZN(P3_U3041) );
  OAI222_X1 U21780 ( .A1(n18687), .A2(n18655), .B1(n18653), .B2(n18697), .C1(
        n18652), .C2(n18691), .ZN(P3_U3042) );
  OAI222_X1 U21781 ( .A1(n18655), .A2(n18691), .B1(n18654), .B2(n18697), .C1(
        n18656), .C2(n18687), .ZN(P3_U3043) );
  OAI222_X1 U21782 ( .A1(n18687), .A2(n18658), .B1(n18657), .B2(n18697), .C1(
        n18656), .C2(n18691), .ZN(P3_U3044) );
  INV_X1 U21783 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18660) );
  OAI222_X1 U21784 ( .A1(n18687), .A2(n18660), .B1(n18659), .B2(n18761), .C1(
        n18658), .C2(n18691), .ZN(P3_U3045) );
  OAI222_X1 U21785 ( .A1(n18687), .A2(n18662), .B1(n18661), .B2(n18761), .C1(
        n18660), .C2(n18691), .ZN(P3_U3046) );
  OAI222_X1 U21786 ( .A1(n18687), .A2(n18664), .B1(n18663), .B2(n18761), .C1(
        n18662), .C2(n18691), .ZN(P3_U3047) );
  OAI222_X1 U21787 ( .A1(n18687), .A2(n18666), .B1(n18665), .B2(n18761), .C1(
        n18664), .C2(n18691), .ZN(P3_U3048) );
  INV_X1 U21788 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18668) );
  OAI222_X1 U21789 ( .A1(n18687), .A2(n18668), .B1(n18667), .B2(n18761), .C1(
        n18666), .C2(n18691), .ZN(P3_U3049) );
  OAI222_X1 U21790 ( .A1(n18687), .A2(n18671), .B1(n18669), .B2(n18761), .C1(
        n18668), .C2(n18691), .ZN(P3_U3050) );
  OAI222_X1 U21791 ( .A1(n18671), .A2(n18691), .B1(n18670), .B2(n18761), .C1(
        n18673), .C2(n18687), .ZN(P3_U3051) );
  OAI222_X1 U21792 ( .A1(n18673), .A2(n18691), .B1(n18672), .B2(n18761), .C1(
        n18674), .C2(n18687), .ZN(P3_U3052) );
  OAI222_X1 U21793 ( .A1(n18687), .A2(n20818), .B1(n18675), .B2(n18761), .C1(
        n18674), .C2(n18691), .ZN(P3_U3053) );
  OAI222_X1 U21794 ( .A1(n20818), .A2(n18691), .B1(n18676), .B2(n18761), .C1(
        n18677), .C2(n18687), .ZN(P3_U3054) );
  OAI222_X1 U21795 ( .A1(n18687), .A2(n18679), .B1(n18678), .B2(n18761), .C1(
        n18677), .C2(n18691), .ZN(P3_U3055) );
  OAI222_X1 U21796 ( .A1(n18687), .A2(n20831), .B1(n18680), .B2(n18697), .C1(
        n18679), .C2(n18691), .ZN(P3_U3056) );
  OAI222_X1 U21797 ( .A1(n18687), .A2(n20825), .B1(n18681), .B2(n18697), .C1(
        n20831), .C2(n18691), .ZN(P3_U3057) );
  OAI222_X1 U21798 ( .A1(n18687), .A2(n18684), .B1(n18682), .B2(n18697), .C1(
        n20825), .C2(n18691), .ZN(P3_U3058) );
  OAI222_X1 U21799 ( .A1(n18684), .A2(n18691), .B1(n18683), .B2(n18697), .C1(
        n18685), .C2(n18687), .ZN(P3_U3059) );
  INV_X1 U21800 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18690) );
  OAI222_X1 U21801 ( .A1(n18687), .A2(n18690), .B1(n18686), .B2(n18697), .C1(
        n18685), .C2(n18691), .ZN(P3_U3060) );
  OAI222_X1 U21802 ( .A1(n18691), .A2(n18690), .B1(n18689), .B2(n18697), .C1(
        n18688), .C2(n18687), .ZN(P3_U3061) );
  INV_X1 U21803 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18692) );
  AOI22_X1 U21804 ( .A1(n18761), .A2(n18693), .B1(n18692), .B2(n18759), .ZN(
        P3_U3274) );
  INV_X1 U21805 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18734) );
  INV_X1 U21806 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18694) );
  AOI22_X1 U21807 ( .A1(n18761), .A2(n18734), .B1(n18694), .B2(n18759), .ZN(
        P3_U3275) );
  INV_X1 U21808 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18695) );
  AOI22_X1 U21809 ( .A1(n18697), .A2(n18696), .B1(n18695), .B2(n18759), .ZN(
        P3_U3276) );
  INV_X1 U21810 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18737) );
  INV_X1 U21811 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18698) );
  AOI22_X1 U21812 ( .A1(n18761), .A2(n18737), .B1(n18698), .B2(n18759), .ZN(
        P3_U3277) );
  OAI21_X1 U21813 ( .B1(n18702), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18700), 
        .ZN(n18699) );
  INV_X1 U21814 ( .A(n18699), .ZN(P3_U3280) );
  INV_X1 U21815 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18701) );
  OAI21_X1 U21816 ( .B1(n18702), .B2(n18701), .A(n18700), .ZN(P3_U3281) );
  OAI221_X1 U21817 ( .B1(n20828), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n20828), 
        .C2(n18704), .A(n18703), .ZN(P3_U3282) );
  AOI22_X1 U21818 ( .A1(n18763), .A2(n18706), .B1(n18725), .B2(n18705), .ZN(
        n18707) );
  AOI22_X1 U21819 ( .A1(n18730), .A2(n18554), .B1(n18707), .B2(n18728), .ZN(
        P3_U3285) );
  AOI22_X1 U21820 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n18709), .B2(n18708), .ZN(
        n18718) );
  NOR2_X1 U21821 ( .A1(n18710), .A2(n18727), .ZN(n18719) );
  INV_X1 U21822 ( .A(n18725), .ZN(n18712) );
  OAI22_X1 U21823 ( .A1(n18714), .A2(n18713), .B1(n18712), .B2(n18711), .ZN(
        n18715) );
  AOI21_X1 U21824 ( .B1(n18718), .B2(n18719), .A(n18715), .ZN(n18716) );
  AOI22_X1 U21825 ( .A1(n18730), .A2(n18717), .B1(n18716), .B2(n18728), .ZN(
        P3_U3288) );
  INV_X1 U21826 ( .A(n18718), .ZN(n18720) );
  AOI222_X1 U21827 ( .A1(n18722), .A2(n18763), .B1(n18725), .B2(n18721), .C1(
        n18720), .C2(n18719), .ZN(n18723) );
  AOI22_X1 U21828 ( .A1(n18730), .A2(n9610), .B1(n18723), .B2(n18728), .ZN(
        P3_U3289) );
  AOI222_X1 U21829 ( .A1(n18727), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18763), 
        .B2(n18726), .C1(n20898), .C2(n18725), .ZN(n18729) );
  AOI22_X1 U21830 ( .A1(n18730), .A2(n9743), .B1(n18729), .B2(n18728), .ZN(
        P3_U3290) );
  INV_X1 U21831 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18732) );
  NOR3_X1 U21832 ( .A1(n18732), .A2(P3_REIP_REG_0__SCAN_IN), .A3(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18731) );
  AOI221_X1 U21833 ( .B1(n18733), .B2(n18732), .C1(P3_REIP_REG_1__SCAN_IN), 
        .C2(P3_REIP_REG_0__SCAN_IN), .A(n18731), .ZN(n18735) );
  INV_X1 U21834 ( .A(n18739), .ZN(n18736) );
  AOI22_X1 U21835 ( .A1(n18739), .A2(n18735), .B1(n18734), .B2(n18736), .ZN(
        P3_U3292) );
  NOR2_X1 U21836 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n18738) );
  AOI22_X1 U21837 ( .A1(n18739), .A2(n18738), .B1(n18737), .B2(n18736), .ZN(
        P3_U3293) );
  INV_X1 U21838 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18740) );
  AOI22_X1 U21839 ( .A1(n18761), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18740), 
        .B2(n18759), .ZN(P3_U3294) );
  MUX2_X1 U21840 ( .A(P3_MORE_REG_SCAN_IN), .B(n18742), .S(n18741), .Z(
        P3_U3295) );
  OAI21_X1 U21841 ( .B1(n18745), .B2(n18744), .A(n18743), .ZN(n18746) );
  AOI21_X1 U21842 ( .B1(n18747), .B2(n18751), .A(n18746), .ZN(n18758) );
  AOI21_X1 U21843 ( .B1(n18750), .B2(n18749), .A(n18748), .ZN(n18752) );
  OAI211_X1 U21844 ( .C1(n18753), .C2(n18752), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18751), .ZN(n18755) );
  AOI21_X1 U21845 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18755), .A(n18754), 
        .ZN(n18757) );
  NAND2_X1 U21846 ( .A1(n18758), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18756) );
  OAI21_X1 U21847 ( .B1(n18758), .B2(n18757), .A(n18756), .ZN(P3_U3296) );
  INV_X1 U21848 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18768) );
  INV_X1 U21849 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18760) );
  AOI22_X1 U21850 ( .A1(n18761), .A2(n18768), .B1(n18760), .B2(n18759), .ZN(
        P3_U3297) );
  AOI21_X1 U21851 ( .B1(n18763), .B2(n18762), .A(n18765), .ZN(n18769) );
  INV_X1 U21852 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18766) );
  AOI22_X1 U21853 ( .A1(n18769), .A2(n18766), .B1(n18765), .B2(n18764), .ZN(
        P3_U3298) );
  AOI21_X1 U21854 ( .B1(n18769), .B2(n18768), .A(n18767), .ZN(P3_U3299) );
  INV_X1 U21855 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18771) );
  INV_X1 U21856 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19733) );
  NAND2_X1 U21857 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19733), .ZN(n19723) );
  INV_X1 U21858 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n18770) );
  NAND2_X1 U21859 ( .A1(n19721), .A2(n18770), .ZN(n19722) );
  OAI21_X1 U21860 ( .B1(n19721), .B2(n19723), .A(n19722), .ZN(n19797) );
  INV_X1 U21861 ( .A(n19797), .ZN(n19716) );
  OAI21_X1 U21862 ( .B1(n19721), .B2(n18771), .A(n19716), .ZN(P2_U2815) );
  AOI22_X1 U21863 ( .A1(n19855), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n19710), 
        .B2(n19711), .ZN(n18772) );
  INV_X1 U21864 ( .A(n18772), .ZN(P2_U2816) );
  AOI22_X1 U21865 ( .A1(P2_D_C_N_REG_SCAN_IN), .A2(n19872), .B1(n18774), .B2(
        n19721), .ZN(n18773) );
  OAI21_X1 U21866 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n19872), .A(n18773), 
        .ZN(P2_U2817) );
  OAI21_X1 U21867 ( .B1(n18774), .B2(BS16), .A(n19797), .ZN(n19795) );
  OAI21_X1 U21868 ( .B1(n19797), .B2(n15620), .A(n19795), .ZN(P2_U2818) );
  NOR2_X1 U21869 ( .A1(n18775), .A2(n19049), .ZN(n19850) );
  OAI21_X1 U21870 ( .B1(n19850), .B2(n12564), .A(n18776), .ZN(P2_U2819) );
  NOR4_X1 U21871 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18780) );
  NOR4_X1 U21872 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n18779) );
  NOR4_X1 U21873 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18778) );
  NOR4_X1 U21874 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18777) );
  NAND4_X1 U21875 ( .A1(n18780), .A2(n18779), .A3(n18778), .A4(n18777), .ZN(
        n18786) );
  NOR4_X1 U21876 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18784) );
  AOI211_X1 U21877 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_10__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18783) );
  NOR4_X1 U21878 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n18782) );
  NOR4_X1 U21879 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n18781) );
  NAND4_X1 U21880 ( .A1(n18784), .A2(n18783), .A3(n18782), .A4(n18781), .ZN(
        n18785) );
  NOR2_X1 U21881 ( .A1(n18786), .A2(n18785), .ZN(n18794) );
  INV_X1 U21882 ( .A(n18794), .ZN(n18793) );
  NOR2_X1 U21883 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18793), .ZN(n18787) );
  INV_X1 U21884 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19793) );
  AOI22_X1 U21885 ( .A1(n18787), .A2(n18788), .B1(n18793), .B2(n19793), .ZN(
        P2_U2820) );
  OR3_X1 U21886 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18792) );
  INV_X1 U21887 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19791) );
  AOI22_X1 U21888 ( .A1(n18787), .A2(n18792), .B1(n18793), .B2(n19791), .ZN(
        P2_U2821) );
  INV_X1 U21889 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19796) );
  NAND2_X1 U21890 ( .A1(n18787), .A2(n19796), .ZN(n18791) );
  OAI21_X1 U21891 ( .B1(n19734), .B2(n18788), .A(n18794), .ZN(n18789) );
  OAI21_X1 U21892 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18794), .A(n18789), 
        .ZN(n18790) );
  OAI221_X1 U21893 ( .B1(n18791), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18791), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18790), .ZN(P2_U2822) );
  INV_X1 U21894 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19789) );
  OAI221_X1 U21895 ( .B1(n18794), .B2(n19789), .C1(n18793), .C2(n18792), .A(
        n18791), .ZN(P2_U2823) );
  INV_X1 U21896 ( .A(n18795), .ZN(n18796) );
  OAI22_X1 U21897 ( .A1(n18797), .A2(n18965), .B1(n18960), .B2(n18796), .ZN(
        n18798) );
  INV_X1 U21898 ( .A(n18798), .ZN(n18806) );
  AOI211_X1 U21899 ( .C1(n18800), .C2(n9708), .A(n18799), .B(n19713), .ZN(
        n18804) );
  AOI22_X1 U21900 ( .A1(n18898), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n18963), .ZN(n18801) );
  OAI21_X1 U21901 ( .B1(n18802), .B2(n18941), .A(n18801), .ZN(n18803) );
  AOI211_X1 U21902 ( .C1(n18957), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n18804), .B(n18803), .ZN(n18805) );
  NAND2_X1 U21903 ( .A1(n18806), .A2(n18805), .ZN(P2_U2835) );
  AOI22_X1 U21904 ( .A1(n18808), .A2(n18902), .B1(n18907), .B2(n18807), .ZN(
        n18816) );
  AOI211_X1 U21905 ( .C1(n18810), .C2(n18809), .A(n9718), .B(n19713), .ZN(
        n18814) );
  INV_X1 U21906 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19764) );
  AOI22_X1 U21907 ( .A1(n18811), .A2(n18958), .B1(P2_EBX_REG_19__SCAN_IN), 
        .B2(n18898), .ZN(n18812) );
  OAI211_X1 U21908 ( .C1(n19764), .C2(n18923), .A(n18812), .B(n18921), .ZN(
        n18813) );
  AOI211_X1 U21909 ( .C1(n18957), .C2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n18814), .B(n18813), .ZN(n18815) );
  NAND2_X1 U21910 ( .A1(n18816), .A2(n18815), .ZN(P2_U2836) );
  XNOR2_X1 U21911 ( .A(n18818), .B(n18817), .ZN(n18829) );
  OAI222_X1 U21912 ( .A1(n18941), .A2(n18821), .B1(n18820), .B2(n18961), .C1(
        n18819), .C2(n18955), .ZN(n18822) );
  AOI211_X1 U21913 ( .C1(P2_REIP_REG_18__SCAN_IN), .C2(n18963), .A(n19119), 
        .B(n18822), .ZN(n18828) );
  INV_X1 U21914 ( .A(n18823), .ZN(n18824) );
  OAI22_X1 U21915 ( .A1(n18825), .A2(n18965), .B1(n18960), .B2(n18824), .ZN(
        n18826) );
  INV_X1 U21916 ( .A(n18826), .ZN(n18827) );
  OAI211_X1 U21917 ( .C1(n19713), .C2(n18829), .A(n18828), .B(n18827), .ZN(
        P2_U2837) );
  AOI22_X1 U21918 ( .A1(n18898), .A2(P2_EBX_REG_17__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n18957), .ZN(n18834) );
  OAI211_X1 U21919 ( .C1(n18832), .C2(n18841), .A(n18831), .B(n18830), .ZN(
        n18833) );
  OAI211_X1 U21920 ( .C1(n18835), .C2(n18941), .A(n18834), .B(n18833), .ZN(
        n18836) );
  AOI211_X1 U21921 ( .C1(P2_REIP_REG_17__SCAN_IN), .C2(n18963), .A(n19119), 
        .B(n18836), .ZN(n18840) );
  AOI22_X1 U21922 ( .A1(n18838), .A2(n18902), .B1(n18907), .B2(n18837), .ZN(
        n18839) );
  OAI211_X1 U21923 ( .C1(n18841), .C2(n18914), .A(n18840), .B(n18839), .ZN(
        P2_U2838) );
  NAND2_X1 U21924 ( .A1(n12901), .A2(n18842), .ZN(n18843) );
  XOR2_X1 U21925 ( .A(n18844), .B(n18843), .Z(n18852) );
  AOI222_X1 U21926 ( .A1(n18898), .A2(P2_EBX_REG_16__SCAN_IN), .B1(n18845), 
        .B2(n18958), .C1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n18957), .ZN(
        n18846) );
  INV_X1 U21927 ( .A(n18846), .ZN(n18847) );
  AOI211_X1 U21928 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n18963), .A(n19119), 
        .B(n18847), .ZN(n18851) );
  AOI22_X1 U21929 ( .A1(n18849), .A2(n18902), .B1(n18907), .B2(n18848), .ZN(
        n18850) );
  OAI211_X1 U21930 ( .C1(n19713), .C2(n18852), .A(n18851), .B(n18850), .ZN(
        P2_U2839) );
  NOR2_X1 U21931 ( .A1(n9927), .A2(n18853), .ZN(n18855) );
  XOR2_X1 U21932 ( .A(n18855), .B(n18854), .Z(n18862) );
  AOI22_X1 U21933 ( .A1(n18856), .A2(n18958), .B1(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18957), .ZN(n18857) );
  OAI21_X1 U21934 ( .B1(n18961), .B2(n11879), .A(n18857), .ZN(n18858) );
  AOI211_X1 U21935 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n18963), .A(n19119), 
        .B(n18858), .ZN(n18861) );
  AOI22_X1 U21936 ( .A1(n18859), .A2(n18902), .B1(n18907), .B2(n18990), .ZN(
        n18860) );
  OAI211_X1 U21937 ( .C1(n19713), .C2(n18862), .A(n18861), .B(n18860), .ZN(
        P2_U2840) );
  NAND2_X1 U21938 ( .A1(n12901), .A2(n18863), .ZN(n18864) );
  XNOR2_X1 U21939 ( .A(n18865), .B(n18864), .ZN(n18873) );
  AOI22_X1 U21940 ( .A1(n18866), .A2(n18958), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n18957), .ZN(n18867) );
  OAI211_X1 U21941 ( .C1(n19756), .C2(n18923), .A(n18867), .B(n18921), .ZN(
        n18868) );
  AOI21_X1 U21942 ( .B1(P2_EBX_REG_14__SCAN_IN), .B2(n18898), .A(n18868), .ZN(
        n18872) );
  AOI22_X1 U21943 ( .A1(n18870), .A2(n18902), .B1(n18907), .B2(n18869), .ZN(
        n18871) );
  OAI211_X1 U21944 ( .C1(n19713), .C2(n18873), .A(n18872), .B(n18871), .ZN(
        P2_U2841) );
  INV_X1 U21945 ( .A(n18874), .ZN(n18876) );
  OAI22_X1 U21946 ( .A1(n18876), .A2(n18941), .B1(n18961), .B2(n18875), .ZN(
        n18877) );
  AOI211_X1 U21947 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n18963), .A(n19119), 
        .B(n18877), .ZN(n18885) );
  NOR2_X1 U21948 ( .A1(n9927), .A2(n18878), .ZN(n18879) );
  XOR2_X1 U21949 ( .A(n18880), .B(n18879), .Z(n18883) );
  OAI22_X1 U21950 ( .A1(n18881), .A2(n18965), .B1(n18960), .B2(n18997), .ZN(
        n18882) );
  AOI21_X1 U21951 ( .B1(n18883), .B2(n18951), .A(n18882), .ZN(n18884) );
  OAI211_X1 U21952 ( .C1(n18886), .C2(n18955), .A(n18885), .B(n18884), .ZN(
        P2_U2842) );
  AND2_X1 U21953 ( .A1(n12901), .A2(n18887), .ZN(n18909) );
  XOR2_X1 U21954 ( .A(n18909), .B(n18888), .Z(n18897) );
  OAI22_X1 U21955 ( .A1(n18890), .A2(n18941), .B1(n18961), .B2(n18889), .ZN(
        n18891) );
  INV_X1 U21956 ( .A(n18891), .ZN(n18892) );
  OAI211_X1 U21957 ( .C1(n19752), .C2(n18923), .A(n18892), .B(n18921), .ZN(
        n18895) );
  OAI22_X1 U21958 ( .A1(n18999), .A2(n18960), .B1(n18965), .B2(n18893), .ZN(
        n18894) );
  AOI211_X1 U21959 ( .C1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n18957), .A(
        n18895), .B(n18894), .ZN(n18896) );
  OAI21_X1 U21960 ( .B1(n18897), .B2(n19713), .A(n18896), .ZN(P2_U2843) );
  INV_X1 U21961 ( .A(n19001), .ZN(n18908) );
  NAND2_X1 U21962 ( .A1(n18963), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n18900) );
  AOI22_X1 U21963 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n18957), .B1(
        P2_EBX_REG_11__SCAN_IN), .B2(n18898), .ZN(n18899) );
  NAND3_X1 U21964 ( .A1(n18900), .A2(n18899), .A3(n18921), .ZN(n18901) );
  AOI21_X1 U21965 ( .B1(n18903), .B2(n18902), .A(n18901), .ZN(n18904) );
  OAI21_X1 U21966 ( .B1(n18905), .B2(n18941), .A(n18904), .ZN(n18906) );
  AOI21_X1 U21967 ( .B1(n18908), .B2(n18907), .A(n18906), .ZN(n18912) );
  OAI211_X1 U21968 ( .C1(n18910), .C2(n18913), .A(n18951), .B(n18909), .ZN(
        n18911) );
  OAI211_X1 U21969 ( .C1(n18914), .C2(n18913), .A(n18912), .B(n18911), .ZN(
        P2_U2844) );
  NAND2_X1 U21970 ( .A1(n12901), .A2(n18915), .ZN(n18917) );
  XOR2_X1 U21971 ( .A(n18917), .B(n18916), .Z(n18928) );
  OAI22_X1 U21972 ( .A1(n18919), .A2(n18941), .B1(n18961), .B2(n18918), .ZN(
        n18920) );
  INV_X1 U21973 ( .A(n18920), .ZN(n18922) );
  OAI211_X1 U21974 ( .C1(n19749), .C2(n18923), .A(n18922), .B(n18921), .ZN(
        n18926) );
  OAI22_X1 U21975 ( .A1(n18924), .A2(n18965), .B1(n18960), .B2(n19004), .ZN(
        n18925) );
  AOI211_X1 U21976 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n18957), .A(
        n18926), .B(n18925), .ZN(n18927) );
  OAI21_X1 U21977 ( .B1(n18928), .B2(n19713), .A(n18927), .ZN(P2_U2845) );
  INV_X1 U21978 ( .A(n18929), .ZN(n18930) );
  OAI22_X1 U21979 ( .A1(n18930), .A2(n18941), .B1(n18961), .B2(n9880), .ZN(
        n18931) );
  AOI211_X1 U21980 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n18963), .A(n19119), .B(
        n18931), .ZN(n18939) );
  NOR2_X1 U21981 ( .A1(n9927), .A2(n18932), .ZN(n18933) );
  XNOR2_X1 U21982 ( .A(n18934), .B(n18933), .ZN(n18937) );
  OAI22_X1 U21983 ( .A1(n18935), .A2(n18965), .B1(n18960), .B2(n19006), .ZN(
        n18936) );
  AOI21_X1 U21984 ( .B1(n18937), .B2(n18951), .A(n18936), .ZN(n18938) );
  OAI211_X1 U21985 ( .C1(n18940), .C2(n18955), .A(n18939), .B(n18938), .ZN(
        P2_U2846) );
  OAI22_X1 U21986 ( .A1(n18942), .A2(n18941), .B1(n18961), .B2(n12306), .ZN(
        n18943) );
  AOI211_X1 U21987 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n18963), .A(n19119), .B(
        n18943), .ZN(n18954) );
  NOR2_X1 U21988 ( .A1(n9927), .A2(n18944), .ZN(n18946) );
  XNOR2_X1 U21989 ( .A(n18947), .B(n18946), .ZN(n18952) );
  INV_X1 U21990 ( .A(n18948), .ZN(n18949) );
  OAI22_X1 U21991 ( .A1(n18949), .A2(n18965), .B1(n19023), .B2(n18960), .ZN(
        n18950) );
  AOI21_X1 U21992 ( .B1(n18952), .B2(n18951), .A(n18950), .ZN(n18953) );
  OAI211_X1 U21993 ( .C1(n18956), .C2(n18955), .A(n18954), .B(n18953), .ZN(
        P2_U2850) );
  AOI22_X1 U21994 ( .A1(n18959), .A2(n18958), .B1(n18957), .B2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18974) );
  OAI22_X1 U21995 ( .A1(n18961), .A2(n11848), .B1(n19025), .B2(n18960), .ZN(
        n18962) );
  AOI211_X1 U21996 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n18963), .A(n19119), .B(
        n18962), .ZN(n18973) );
  OAI22_X1 U21997 ( .A1(n19027), .A2(n18966), .B1(n18965), .B2(n18964), .ZN(
        n18967) );
  INV_X1 U21998 ( .A(n18967), .ZN(n18972) );
  AND2_X1 U21999 ( .A1(n12901), .A2(n18968), .ZN(n18970) );
  AOI21_X1 U22000 ( .B1(n19117), .B2(n18970), .A(n19713), .ZN(n18969) );
  OAI21_X1 U22001 ( .B1(n19117), .B2(n18970), .A(n18969), .ZN(n18971) );
  NAND4_X1 U22002 ( .A1(n18974), .A2(n18973), .A3(n18972), .A4(n18971), .ZN(
        P2_U2851) );
  AOI22_X1 U22003 ( .A1(n18975), .A2(n19040), .B1(n18980), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n18977) );
  AOI22_X1 U22004 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19039), .B1(n18981), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n18976) );
  NAND2_X1 U22005 ( .A1(n18977), .A2(n18976), .ZN(P2_U2888) );
  AOI22_X1 U22006 ( .A1(n18979), .A2(n18978), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n19039), .ZN(n18989) );
  AOI22_X1 U22007 ( .A1(n18981), .A2(BUF1_REG_16__SCAN_IN), .B1(n18980), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n18988) );
  OAI22_X1 U22008 ( .A1(n18985), .A2(n18984), .B1(n18983), .B2(n18982), .ZN(
        n18986) );
  INV_X1 U22009 ( .A(n18986), .ZN(n18987) );
  NAND3_X1 U22010 ( .A1(n18989), .A2(n18988), .A3(n18987), .ZN(P2_U2903) );
  INV_X1 U22011 ( .A(n18990), .ZN(n18992) );
  OAI222_X1 U22012 ( .A1(n18992), .A2(n19024), .B1(n12500), .B2(n19014), .C1(
        n18991), .C2(n19048), .ZN(P2_U2904) );
  AOI22_X1 U22013 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19039), .B1(n18993), 
        .B2(n19008), .ZN(n18994) );
  OAI21_X1 U22014 ( .B1(n19024), .B2(n18995), .A(n18994), .ZN(P2_U2905) );
  INV_X1 U22015 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19089) );
  OAI222_X1 U22016 ( .A1(n18997), .A2(n19024), .B1(n19089), .B2(n19014), .C1(
        n19048), .C2(n18996), .ZN(P2_U2906) );
  INV_X1 U22017 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n20850) );
  OAI222_X1 U22018 ( .A1(n18999), .A2(n19024), .B1(n20850), .B2(n19014), .C1(
        n19048), .C2(n18998), .ZN(P2_U2907) );
  INV_X1 U22019 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19092) );
  OAI222_X1 U22020 ( .A1(n19001), .A2(n19024), .B1(n19092), .B2(n19014), .C1(
        n19048), .C2(n19000), .ZN(P2_U2908) );
  AOI22_X1 U22021 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19039), .B1(n19002), 
        .B2(n19008), .ZN(n19003) );
  OAI21_X1 U22022 ( .B1(n19024), .B2(n19004), .A(n19003), .ZN(P2_U2909) );
  INV_X1 U22023 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19096) );
  OAI222_X1 U22024 ( .A1(n19006), .A2(n19024), .B1(n19096), .B2(n19014), .C1(
        n19048), .C2(n19005), .ZN(P2_U2910) );
  INV_X1 U22025 ( .A(n19007), .ZN(n19011) );
  AOI22_X1 U22026 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n19039), .B1(n19009), .B2(
        n19008), .ZN(n19010) );
  OAI21_X1 U22027 ( .B1(n19024), .B2(n19011), .A(n19010), .ZN(P2_U2911) );
  INV_X1 U22028 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19100) );
  OAI222_X1 U22029 ( .A1(n19012), .A2(n19024), .B1(n19100), .B2(n19014), .C1(
        n19048), .C2(n19188), .ZN(P2_U2912) );
  INV_X1 U22030 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19102) );
  OAI222_X1 U22031 ( .A1(n19013), .A2(n19024), .B1(n19102), .B2(n19014), .C1(
        n19048), .C2(n19182), .ZN(P2_U2913) );
  INV_X1 U22032 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19104) );
  OAI22_X1 U22033 ( .A1(n19104), .A2(n19014), .B1(n19178), .B2(n19048), .ZN(
        n19015) );
  INV_X1 U22034 ( .A(n19015), .ZN(n19022) );
  INV_X1 U22035 ( .A(n19018), .ZN(n19804) );
  INV_X1 U22036 ( .A(n19445), .ZN(n19803) );
  INV_X1 U22037 ( .A(n19813), .ZN(n19017) );
  OAI21_X1 U22038 ( .B1(n19017), .B2(n19817), .A(n19016), .ZN(n19034) );
  XOR2_X1 U22039 ( .A(n19018), .B(n19445), .Z(n19035) );
  NAND2_X1 U22040 ( .A1(n19034), .A2(n19035), .ZN(n19033) );
  OAI21_X1 U22041 ( .B1(n19804), .B2(n19803), .A(n19033), .ZN(n19019) );
  NAND2_X1 U22042 ( .A1(n19019), .A2(n19025), .ZN(n19028) );
  INV_X1 U22043 ( .A(n19027), .ZN(n19020) );
  NAND3_X1 U22044 ( .A1(n19028), .A2(n19020), .A3(n19044), .ZN(n19021) );
  OAI211_X1 U22045 ( .C1(n19024), .C2(n19023), .A(n19022), .B(n19021), .ZN(
        P2_U2914) );
  INV_X1 U22046 ( .A(n19025), .ZN(n19026) );
  AOI22_X1 U22047 ( .A1(n19040), .A2(n19026), .B1(n19039), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n19031) );
  XNOR2_X1 U22048 ( .A(n19028), .B(n19027), .ZN(n19029) );
  NAND2_X1 U22049 ( .A1(n19029), .A2(n19044), .ZN(n19030) );
  OAI211_X1 U22050 ( .C1(n19032), .C2(n19048), .A(n19031), .B(n19030), .ZN(
        P2_U2915) );
  AOI22_X1 U22051 ( .A1(n19804), .A2(n19040), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19039), .ZN(n19038) );
  OAI21_X1 U22052 ( .B1(n19035), .B2(n19034), .A(n19033), .ZN(n19036) );
  NAND2_X1 U22053 ( .A1(n19036), .A2(n19044), .ZN(n19037) );
  OAI211_X1 U22054 ( .C1(n19173), .C2(n19048), .A(n19038), .B(n19037), .ZN(
        P2_U2916) );
  AOI22_X1 U22055 ( .A1(n19040), .A2(n19826), .B1(n19039), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19047) );
  OAI21_X1 U22056 ( .B1(n19043), .B2(n19042), .A(n19041), .ZN(n19045) );
  NAND2_X1 U22057 ( .A1(n19045), .A2(n19044), .ZN(n19046) );
  OAI211_X1 U22058 ( .C1(n19168), .C2(n19048), .A(n19047), .B(n19046), .ZN(
        P2_U2918) );
  OR2_X1 U22059 ( .A1(n19050), .A2(n19049), .ZN(n19052) );
  OAI21_X1 U22060 ( .B1(n19053), .B2(n19052), .A(n19051), .ZN(n19054) );
  AND2_X1 U22061 ( .A1(n19054), .A2(n19866), .ZN(n19084) );
  NOR2_X1 U22062 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19831), .ZN(n19106) );
  AND2_X1 U22063 ( .A1(n19114), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NAND2_X1 U22064 ( .A1(n19084), .A2(n19055), .ZN(n19082) );
  AOI22_X1 U22065 ( .A1(n19858), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19111), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n19056) );
  OAI21_X1 U22066 ( .B1(n19057), .B2(n19082), .A(n19056), .ZN(P2_U2921) );
  AOI22_X1 U22067 ( .A1(n19858), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19111), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n19058) );
  OAI21_X1 U22068 ( .B1(n19059), .B2(n19082), .A(n19058), .ZN(P2_U2922) );
  AOI22_X1 U22069 ( .A1(n19858), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19111), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n19060) );
  OAI21_X1 U22070 ( .B1(n19061), .B2(n19082), .A(n19060), .ZN(P2_U2923) );
  AOI22_X1 U22071 ( .A1(n19858), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19114), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n19062) );
  OAI21_X1 U22072 ( .B1(n19063), .B2(n19082), .A(n19062), .ZN(P2_U2924) );
  AOI22_X1 U22073 ( .A1(n19858), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19111), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n19064) );
  OAI21_X1 U22074 ( .B1(n19065), .B2(n19082), .A(n19064), .ZN(P2_U2925) );
  AOI22_X1 U22075 ( .A1(n19858), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19114), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n19066) );
  OAI21_X1 U22076 ( .B1(n19067), .B2(n19082), .A(n19066), .ZN(P2_U2926) );
  AOI22_X1 U22077 ( .A1(n19858), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19111), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n19068) );
  OAI21_X1 U22078 ( .B1(n15101), .B2(n19082), .A(n19068), .ZN(P2_U2927) );
  AOI22_X1 U22079 ( .A1(n19858), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19111), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n19069) );
  OAI21_X1 U22080 ( .B1(n19070), .B2(n19082), .A(n19069), .ZN(P2_U2928) );
  AOI22_X1 U22081 ( .A1(n19858), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19111), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n19071) );
  OAI21_X1 U22082 ( .B1(n12668), .B2(n19082), .A(n19071), .ZN(P2_U2929) );
  AOI22_X1 U22083 ( .A1(n19858), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19111), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n19072) );
  OAI21_X1 U22084 ( .B1(n19073), .B2(n19082), .A(n19072), .ZN(P2_U2930) );
  AOI22_X1 U22085 ( .A1(n19858), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19111), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n19074) );
  OAI21_X1 U22086 ( .B1(n12659), .B2(n19082), .A(n19074), .ZN(P2_U2931) );
  AOI22_X1 U22087 ( .A1(n19858), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19111), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n19075) );
  OAI21_X1 U22088 ( .B1(n19076), .B2(n19082), .A(n19075), .ZN(P2_U2932) );
  INV_X1 U22089 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n19078) );
  AOI22_X1 U22090 ( .A1(n19858), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19111), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n19077) );
  OAI21_X1 U22091 ( .B1(n19078), .B2(n19082), .A(n19077), .ZN(P2_U2933) );
  AOI22_X1 U22092 ( .A1(n19858), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19111), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n19079) );
  OAI21_X1 U22093 ( .B1(n19080), .B2(n19082), .A(n19079), .ZN(P2_U2934) );
  AOI22_X1 U22094 ( .A1(n19858), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19111), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n19081) );
  OAI21_X1 U22095 ( .B1(n19083), .B2(n19082), .A(n19081), .ZN(P2_U2935) );
  AOI22_X1 U22096 ( .A1(n19858), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19111), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19085) );
  OAI21_X1 U22097 ( .B1(n12500), .B2(n19116), .A(n19085), .ZN(P2_U2936) );
  AOI22_X1 U22098 ( .A1(n19858), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19111), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19086) );
  OAI21_X1 U22099 ( .B1(n19087), .B2(n19116), .A(n19086), .ZN(P2_U2937) );
  AOI22_X1 U22100 ( .A1(n19858), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19111), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19088) );
  OAI21_X1 U22101 ( .B1(n19089), .B2(n19116), .A(n19088), .ZN(P2_U2938) );
  AOI22_X1 U22102 ( .A1(n19106), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19111), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19090) );
  OAI21_X1 U22103 ( .B1(n20850), .B2(n19116), .A(n19090), .ZN(P2_U2939) );
  AOI22_X1 U22104 ( .A1(n19106), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19114), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19091) );
  OAI21_X1 U22105 ( .B1(n19092), .B2(n19116), .A(n19091), .ZN(P2_U2940) );
  AOI22_X1 U22106 ( .A1(n19106), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19114), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19093) );
  OAI21_X1 U22107 ( .B1(n19094), .B2(n19116), .A(n19093), .ZN(P2_U2941) );
  AOI22_X1 U22108 ( .A1(n19106), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19114), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19095) );
  OAI21_X1 U22109 ( .B1(n19096), .B2(n19116), .A(n19095), .ZN(P2_U2942) );
  AOI22_X1 U22110 ( .A1(n19106), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19114), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19097) );
  OAI21_X1 U22111 ( .B1(n19098), .B2(n19116), .A(n19097), .ZN(P2_U2943) );
  AOI22_X1 U22112 ( .A1(n19106), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19114), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19099) );
  OAI21_X1 U22113 ( .B1(n19100), .B2(n19116), .A(n19099), .ZN(P2_U2944) );
  AOI22_X1 U22114 ( .A1(n19106), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19114), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19101) );
  OAI21_X1 U22115 ( .B1(n19102), .B2(n19116), .A(n19101), .ZN(P2_U2945) );
  AOI22_X1 U22116 ( .A1(n19106), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19114), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19103) );
  OAI21_X1 U22117 ( .B1(n19104), .B2(n19116), .A(n19103), .ZN(P2_U2946) );
  AOI22_X1 U22118 ( .A1(n19106), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19111), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19105) );
  OAI21_X1 U22119 ( .B1(n12680), .B2(n19116), .A(n19105), .ZN(P2_U2947) );
  INV_X1 U22120 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19108) );
  AOI22_X1 U22121 ( .A1(n19106), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19111), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19107) );
  OAI21_X1 U22122 ( .B1(n19108), .B2(n19116), .A(n19107), .ZN(P2_U2948) );
  INV_X1 U22123 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19110) );
  AOI22_X1 U22124 ( .A1(n19858), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19111), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19109) );
  OAI21_X1 U22125 ( .B1(n19110), .B2(n19116), .A(n19109), .ZN(P2_U2949) );
  INV_X1 U22126 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19113) );
  AOI22_X1 U22127 ( .A1(n19858), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19111), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19112) );
  OAI21_X1 U22128 ( .B1(n19113), .B2(n19116), .A(n19112), .ZN(P2_U2950) );
  AOI22_X1 U22129 ( .A1(P2_LWORD_REG_0__SCAN_IN), .A2(n19858), .B1(n19114), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19115) );
  OAI21_X1 U22130 ( .B1(n12498), .B2(n19116), .A(n19115), .ZN(P2_U2951) );
  AOI22_X1 U22131 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19119), .B1(n19118), 
        .B2(n19117), .ZN(n19127) );
  AOI222_X1 U22132 ( .A1(n19125), .A2(n19124), .B1(n19123), .B2(n19122), .C1(
        n19121), .C2(n19120), .ZN(n19126) );
  OAI211_X1 U22133 ( .C1(n19129), .C2(n19128), .A(n19127), .B(n19126), .ZN(
        P2_U3010) );
  NAND3_X1 U22134 ( .A1(n19132), .A2(n19131), .A3(n19130), .ZN(n19135) );
  NAND2_X1 U22135 ( .A1(n19133), .A2(n19149), .ZN(n19134) );
  OAI211_X1 U22136 ( .C1(n19736), .C2(n18921), .A(n19135), .B(n19134), .ZN(
        n19139) );
  NOR2_X1 U22137 ( .A1(n19137), .A2(n19136), .ZN(n19138) );
  INV_X1 U22138 ( .A(n19140), .ZN(n19141) );
  AOI21_X1 U22139 ( .B1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n19142), .A(
        n19141), .ZN(n19147) );
  OAI21_X1 U22140 ( .B1(n19145), .B2(n19144), .A(n19143), .ZN(n19146) );
  OAI211_X1 U22141 ( .C1(n19148), .C2(n19159), .A(n19147), .B(n19146), .ZN(
        P2_U3044) );
  AOI21_X1 U22142 ( .B1(n19151), .B2(n19150), .A(n19149), .ZN(n19152) );
  NAND2_X1 U22143 ( .A1(n19153), .A2(n19152), .ZN(n19163) );
  AOI22_X1 U22144 ( .A1(n19155), .A2(n19826), .B1(n19154), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19162) );
  NAND2_X1 U22145 ( .A1(n19157), .A2(n19156), .ZN(n19161) );
  OR2_X1 U22146 ( .A1(n19159), .A2(n19158), .ZN(n19160) );
  AND4_X1 U22147 ( .A1(n19163), .A2(n19162), .A3(n19161), .A4(n19160), .ZN(
        n19165) );
  OAI211_X1 U22148 ( .C1(n19167), .C2(n19166), .A(n19165), .B(n19164), .ZN(
        P2_U3045) );
  INV_X1 U22149 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19171) );
  AOI22_X1 U22150 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19190), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19189), .ZN(n19666) );
  AOI22_X1 U22151 ( .A1(n19611), .A2(n19702), .B1(n19187), .B2(n19661), .ZN(
        n19170) );
  NOR2_X2 U22152 ( .A1(n19168), .A2(n19650), .ZN(n19662) );
  AOI22_X1 U22153 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19190), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19189), .ZN(n19614) );
  AOI22_X1 U22154 ( .A1(n19662), .A2(n19191), .B1(n19246), .B2(n19663), .ZN(
        n19169) );
  OAI211_X1 U22155 ( .C1(n19195), .C2(n19171), .A(n19170), .B(n19169), .ZN(
        P2_U3049) );
  AOI22_X1 U22156 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19189), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19190), .ZN(n19678) );
  INV_X1 U22157 ( .A(n19678), .ZN(n19617) );
  AND2_X1 U22158 ( .A1(n11768), .A2(n19172), .ZN(n19673) );
  AOI22_X1 U22159 ( .A1(n19617), .A2(n19702), .B1(n19187), .B2(n19673), .ZN(
        n19175) );
  NOR2_X2 U22160 ( .A1(n19173), .A2(n19650), .ZN(n19674) );
  AOI22_X1 U22161 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19190), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19189), .ZN(n19620) );
  AOI22_X1 U22162 ( .A1(n19674), .A2(n19191), .B1(n19246), .B2(n19675), .ZN(
        n19174) );
  OAI211_X1 U22163 ( .C1(n19195), .C2(n19176), .A(n19175), .B(n19174), .ZN(
        P2_U3051) );
  INV_X1 U22164 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20797) );
  AOI22_X1 U22165 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19189), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19190), .ZN(n19690) );
  NOR2_X2 U22166 ( .A1(n19177), .A2(n19186), .ZN(n19685) );
  AOI22_X1 U22167 ( .A1(n19625), .A2(n19702), .B1(n19187), .B2(n19685), .ZN(
        n19180) );
  NOR2_X2 U22168 ( .A1(n19178), .A2(n19650), .ZN(n19686) );
  AOI22_X1 U22169 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19190), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19189), .ZN(n19628) );
  AOI22_X1 U22170 ( .A1(n19686), .A2(n19191), .B1(n19246), .B2(n19687), .ZN(
        n19179) );
  OAI211_X1 U22171 ( .C1(n19195), .C2(n20797), .A(n19180), .B(n19179), .ZN(
        P2_U3053) );
  AOI22_X1 U22172 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19190), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19189), .ZN(n19696) );
  INV_X1 U22173 ( .A(n19696), .ZN(n19555) );
  NOR2_X2 U22174 ( .A1(n19181), .A2(n19186), .ZN(n19691) );
  AOI22_X1 U22175 ( .A1(n19555), .A2(n19702), .B1(n19187), .B2(n19691), .ZN(
        n19184) );
  NOR2_X2 U22176 ( .A1(n19182), .A2(n19650), .ZN(n19692) );
  AOI22_X1 U22177 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19190), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19189), .ZN(n19558) );
  AOI22_X1 U22178 ( .A1(n19692), .A2(n19191), .B1(n19246), .B2(n19693), .ZN(
        n19183) );
  OAI211_X1 U22179 ( .C1(n19195), .C2(n19185), .A(n19184), .B(n19183), .ZN(
        P2_U3054) );
  AOI22_X1 U22180 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19190), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19189), .ZN(n19707) );
  NOR2_X2 U22181 ( .A1(n11773), .A2(n19186), .ZN(n19697) );
  AOI22_X1 U22182 ( .A1(n19635), .A2(n19702), .B1(n19187), .B2(n19697), .ZN(
        n19193) );
  NOR2_X2 U22183 ( .A1(n19188), .A2(n19650), .ZN(n19699) );
  AOI22_X1 U22184 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19190), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19189), .ZN(n19640) );
  INV_X1 U22185 ( .A(n19640), .ZN(n19701) );
  AOI22_X1 U22186 ( .A1(n19699), .A2(n19191), .B1(n19246), .B2(n19701), .ZN(
        n19192) );
  OAI211_X1 U22187 ( .C1(n19195), .C2(n19194), .A(n19193), .B(n19192), .ZN(
        P2_U3055) );
  NOR2_X1 U22188 ( .A1(n19447), .A2(n19277), .ZN(n19209) );
  INV_X1 U22189 ( .A(n19209), .ZN(n19241) );
  NAND2_X1 U22190 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19241), .ZN(n19196) );
  NOR2_X1 U22191 ( .A1(n19197), .A2(n19196), .ZN(n19205) );
  INV_X1 U22192 ( .A(n19206), .ZN(n19198) );
  NOR2_X1 U22193 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19198), .ZN(n19199) );
  INV_X1 U22194 ( .A(n19646), .ZN(n19201) );
  OAI22_X1 U22195 ( .A1(n19244), .A2(n19201), .B1(n19200), .B2(n19241), .ZN(
        n19202) );
  INV_X1 U22196 ( .A(n19202), .ZN(n19211) );
  NAND2_X1 U22197 ( .A1(n19445), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19391) );
  INV_X1 U22198 ( .A(n19391), .ZN(n19204) );
  INV_X1 U22199 ( .A(n19452), .ZN(n19203) );
  NAND2_X1 U22200 ( .A1(n19204), .A2(n19203), .ZN(n19207) );
  AOI21_X1 U22201 ( .B1(n19207), .B2(n19206), .A(n19205), .ZN(n19208) );
  OAI211_X1 U22202 ( .C1(n19209), .C2(n19416), .A(n19208), .B(n19604), .ZN(
        n19247) );
  AOI22_X1 U22203 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19247), .B1(
        n19246), .B2(n19575), .ZN(n19210) );
  OAI211_X1 U22204 ( .C1(n19578), .C2(n19250), .A(n19211), .B(n19210), .ZN(
        P2_U3056) );
  INV_X1 U22205 ( .A(n19662), .ZN(n19213) );
  INV_X1 U22206 ( .A(n19661), .ZN(n19212) );
  OAI22_X1 U22207 ( .A1(n19244), .A2(n19213), .B1(n19212), .B2(n19241), .ZN(
        n19214) );
  INV_X1 U22208 ( .A(n19214), .ZN(n19216) );
  AOI22_X1 U22209 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19247), .B1(
        n19246), .B2(n19611), .ZN(n19215) );
  OAI211_X1 U22210 ( .C1(n19614), .C2(n19250), .A(n19216), .B(n19215), .ZN(
        P2_U3057) );
  INV_X1 U22211 ( .A(n19668), .ZN(n19218) );
  OAI22_X1 U22212 ( .A1(n19244), .A2(n19218), .B1(n19217), .B2(n19241), .ZN(
        n19219) );
  INV_X1 U22213 ( .A(n19219), .ZN(n19221) );
  AOI22_X1 U22214 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19247), .B1(
        n19246), .B2(n19544), .ZN(n19220) );
  OAI211_X1 U22215 ( .C1(n19547), .C2(n19250), .A(n19221), .B(n19220), .ZN(
        P2_U3058) );
  INV_X1 U22216 ( .A(n19674), .ZN(n19223) );
  INV_X1 U22217 ( .A(n19673), .ZN(n19222) );
  OAI22_X1 U22218 ( .A1(n19244), .A2(n19223), .B1(n19222), .B2(n19241), .ZN(
        n19224) );
  INV_X1 U22219 ( .A(n19224), .ZN(n19226) );
  AOI22_X1 U22220 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19247), .B1(
        n19246), .B2(n19617), .ZN(n19225) );
  OAI211_X1 U22221 ( .C1(n19620), .C2(n19250), .A(n19226), .B(n19225), .ZN(
        P2_U3059) );
  INV_X1 U22222 ( .A(n19680), .ZN(n19227) );
  OAI22_X1 U22223 ( .A1(n19244), .A2(n19227), .B1(n19260), .B2(n19241), .ZN(
        n19228) );
  INV_X1 U22224 ( .A(n19228), .ZN(n19230) );
  AOI22_X1 U22225 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19247), .B1(
        n19246), .B2(n19621), .ZN(n19229) );
  OAI211_X1 U22226 ( .C1(n19624), .C2(n19250), .A(n19230), .B(n19229), .ZN(
        P2_U3060) );
  INV_X1 U22227 ( .A(n19686), .ZN(n19232) );
  INV_X1 U22228 ( .A(n19685), .ZN(n19231) );
  OAI22_X1 U22229 ( .A1(n19244), .A2(n19232), .B1(n19231), .B2(n19241), .ZN(
        n19233) );
  INV_X1 U22230 ( .A(n19233), .ZN(n19235) );
  AOI22_X1 U22231 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19247), .B1(
        n19246), .B2(n19625), .ZN(n19234) );
  OAI211_X1 U22232 ( .C1(n19628), .C2(n19250), .A(n19235), .B(n19234), .ZN(
        P2_U3061) );
  INV_X1 U22233 ( .A(n19692), .ZN(n19237) );
  INV_X1 U22234 ( .A(n19691), .ZN(n19236) );
  OAI22_X1 U22235 ( .A1(n19244), .A2(n19237), .B1(n19236), .B2(n19241), .ZN(
        n19238) );
  INV_X1 U22236 ( .A(n19238), .ZN(n19240) );
  AOI22_X1 U22237 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19247), .B1(
        n19246), .B2(n19555), .ZN(n19239) );
  OAI211_X1 U22238 ( .C1(n19558), .C2(n19250), .A(n19240), .B(n19239), .ZN(
        P2_U3062) );
  INV_X1 U22239 ( .A(n19699), .ZN(n19243) );
  INV_X1 U22240 ( .A(n19697), .ZN(n19242) );
  OAI22_X1 U22241 ( .A1(n19244), .A2(n19243), .B1(n19242), .B2(n19241), .ZN(
        n19245) );
  INV_X1 U22242 ( .A(n19245), .ZN(n19249) );
  AOI22_X1 U22243 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19247), .B1(
        n19246), .B2(n19635), .ZN(n19248) );
  OAI211_X1 U22244 ( .C1(n19640), .C2(n19250), .A(n19249), .B(n19248), .ZN(
        P2_U3063) );
  INV_X1 U22245 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n19253) );
  AOI22_X1 U22246 ( .A1(n19271), .A2(n19662), .B1(n19270), .B2(n19661), .ZN(
        n19252) );
  AOI22_X1 U22247 ( .A1(n19302), .A2(n19663), .B1(n19272), .B2(n19611), .ZN(
        n19251) );
  OAI211_X1 U22248 ( .C1(n19276), .C2(n19253), .A(n19252), .B(n19251), .ZN(
        P2_U3065) );
  INV_X1 U22249 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n19256) );
  AOI22_X1 U22250 ( .A1(n19271), .A2(n19668), .B1(n19270), .B2(n19667), .ZN(
        n19255) );
  AOI22_X1 U22251 ( .A1(n19302), .A2(n19669), .B1(n19272), .B2(n19544), .ZN(
        n19254) );
  OAI211_X1 U22252 ( .C1(n19276), .C2(n19256), .A(n19255), .B(n19254), .ZN(
        P2_U3066) );
  INV_X1 U22253 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n19259) );
  AOI22_X1 U22254 ( .A1(n19271), .A2(n19674), .B1(n19270), .B2(n19673), .ZN(
        n19258) );
  AOI22_X1 U22255 ( .A1(n19302), .A2(n19675), .B1(n19272), .B2(n19617), .ZN(
        n19257) );
  OAI211_X1 U22256 ( .C1(n19276), .C2(n19259), .A(n19258), .B(n19257), .ZN(
        P2_U3067) );
  INV_X1 U22257 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n19263) );
  AOI22_X1 U22258 ( .A1(n19271), .A2(n19680), .B1(n19270), .B2(n19679), .ZN(
        n19262) );
  AOI22_X1 U22259 ( .A1(n19302), .A2(n19681), .B1(n19272), .B2(n19621), .ZN(
        n19261) );
  OAI211_X1 U22260 ( .C1(n19276), .C2(n19263), .A(n19262), .B(n19261), .ZN(
        P2_U3068) );
  INV_X1 U22261 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n19266) );
  AOI22_X1 U22262 ( .A1(n19271), .A2(n19686), .B1(n19270), .B2(n19685), .ZN(
        n19265) );
  AOI22_X1 U22263 ( .A1(n19302), .A2(n19687), .B1(n19272), .B2(n19625), .ZN(
        n19264) );
  OAI211_X1 U22264 ( .C1(n19276), .C2(n19266), .A(n19265), .B(n19264), .ZN(
        P2_U3069) );
  INV_X1 U22265 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n19269) );
  AOI22_X1 U22266 ( .A1(n19271), .A2(n19692), .B1(n19270), .B2(n19691), .ZN(
        n19268) );
  AOI22_X1 U22267 ( .A1(n19302), .A2(n19693), .B1(n19272), .B2(n19555), .ZN(
        n19267) );
  OAI211_X1 U22268 ( .C1(n19276), .C2(n19269), .A(n19268), .B(n19267), .ZN(
        P2_U3070) );
  INV_X1 U22269 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n19275) );
  AOI22_X1 U22270 ( .A1(n19271), .A2(n19699), .B1(n19270), .B2(n19697), .ZN(
        n19274) );
  AOI22_X1 U22271 ( .A1(n19302), .A2(n19701), .B1(n19272), .B2(n19635), .ZN(
        n19273) );
  OAI211_X1 U22272 ( .C1(n19276), .C2(n19275), .A(n19274), .B(n19273), .ZN(
        P2_U3071) );
  NOR2_X1 U22273 ( .A1(n19510), .A2(n19277), .ZN(n19301) );
  AOI22_X1 U22274 ( .A1(n19575), .A2(n19302), .B1(n19645), .B2(n19301), .ZN(
        n19287) );
  OAI21_X1 U22275 ( .B1(n19391), .B2(n19516), .A(n19812), .ZN(n19285) );
  NAND2_X1 U22276 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19278), .ZN(
        n19284) );
  INV_X1 U22277 ( .A(n19284), .ZN(n19282) );
  OAI21_X1 U22278 ( .B1(n13660), .B2(n19852), .A(n19416), .ZN(n19280) );
  INV_X1 U22279 ( .A(n19301), .ZN(n19279) );
  NAND2_X1 U22280 ( .A1(n19280), .A2(n19279), .ZN(n19281) );
  OAI211_X1 U22281 ( .C1(n19285), .C2(n19282), .A(n19604), .B(n19281), .ZN(
        n19304) );
  OAI21_X1 U22282 ( .B1(n13660), .B2(n19301), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19283) );
  OAI21_X1 U22283 ( .B1(n19285), .B2(n19284), .A(n19283), .ZN(n19303) );
  AOI22_X1 U22284 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19304), .B1(
        n19646), .B2(n19303), .ZN(n19286) );
  OAI211_X1 U22285 ( .C1(n19578), .C2(n19334), .A(n19287), .B(n19286), .ZN(
        P2_U3072) );
  AOI22_X1 U22286 ( .A1(n19663), .A2(n19324), .B1(n19301), .B2(n19661), .ZN(
        n19289) );
  AOI22_X1 U22287 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19304), .B1(
        n19662), .B2(n19303), .ZN(n19288) );
  OAI211_X1 U22288 ( .C1(n19666), .C2(n19298), .A(n19289), .B(n19288), .ZN(
        P2_U3073) );
  AOI22_X1 U22289 ( .A1(n19669), .A2(n19324), .B1(n19667), .B2(n19301), .ZN(
        n19291) );
  AOI22_X1 U22290 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19304), .B1(
        n19668), .B2(n19303), .ZN(n19290) );
  OAI211_X1 U22291 ( .C1(n19672), .C2(n19298), .A(n19291), .B(n19290), .ZN(
        P2_U3074) );
  AOI22_X1 U22292 ( .A1(n19675), .A2(n19324), .B1(n19301), .B2(n19673), .ZN(
        n19293) );
  AOI22_X1 U22293 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19304), .B1(
        n19674), .B2(n19303), .ZN(n19292) );
  OAI211_X1 U22294 ( .C1(n19678), .C2(n19298), .A(n19293), .B(n19292), .ZN(
        P2_U3075) );
  AOI22_X1 U22295 ( .A1(n19681), .A2(n19324), .B1(n19679), .B2(n19301), .ZN(
        n19295) );
  AOI22_X1 U22296 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19304), .B1(
        n19680), .B2(n19303), .ZN(n19294) );
  OAI211_X1 U22297 ( .C1(n19684), .C2(n19298), .A(n19295), .B(n19294), .ZN(
        P2_U3076) );
  AOI22_X1 U22298 ( .A1(n19687), .A2(n19324), .B1(n19301), .B2(n19685), .ZN(
        n19297) );
  AOI22_X1 U22299 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19304), .B1(
        n19686), .B2(n19303), .ZN(n19296) );
  OAI211_X1 U22300 ( .C1(n19690), .C2(n19298), .A(n19297), .B(n19296), .ZN(
        P2_U3077) );
  AOI22_X1 U22301 ( .A1(n19555), .A2(n19302), .B1(n19301), .B2(n19691), .ZN(
        n19300) );
  AOI22_X1 U22302 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19304), .B1(
        n19692), .B2(n19303), .ZN(n19299) );
  OAI211_X1 U22303 ( .C1(n19558), .C2(n19334), .A(n19300), .B(n19299), .ZN(
        P2_U3078) );
  AOI22_X1 U22304 ( .A1(n19635), .A2(n19302), .B1(n19301), .B2(n19697), .ZN(
        n19306) );
  AOI22_X1 U22305 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19304), .B1(
        n19699), .B2(n19303), .ZN(n19305) );
  OAI211_X1 U22306 ( .C1(n19640), .C2(n19334), .A(n19306), .B(n19305), .ZN(
        P2_U3079) );
  NAND2_X1 U22307 ( .A1(n19307), .A2(n19811), .ZN(n19312) );
  INV_X1 U22308 ( .A(n19812), .ZN(n19807) );
  NOR2_X1 U22309 ( .A1(n19387), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19339) );
  INV_X1 U22310 ( .A(n19339), .ZN(n19341) );
  NOR2_X1 U22311 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19341), .ZN(
        n19329) );
  OAI21_X1 U22312 ( .B1(n13544), .B2(n19329), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19308) );
  OAI21_X1 U22313 ( .B1(n19312), .B2(n19807), .A(n19308), .ZN(n19330) );
  AOI22_X1 U22314 ( .A1(n19330), .A2(n19646), .B1(n19645), .B2(n19329), .ZN(
        n19315) );
  OAI21_X1 U22315 ( .B1(n19324), .B2(n19349), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19311) );
  AOI211_X1 U22316 ( .C1(n13544), .C2(n19416), .A(n19329), .B(n19812), .ZN(
        n19310) );
  AOI211_X1 U22317 ( .C1(n19312), .C2(n19311), .A(n19650), .B(n19310), .ZN(
        n19313) );
  AOI22_X1 U22318 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19331), .B1(
        n19349), .B2(n19657), .ZN(n19314) );
  OAI211_X1 U22319 ( .C1(n19660), .C2(n19334), .A(n19315), .B(n19314), .ZN(
        P2_U3080) );
  AOI22_X1 U22320 ( .A1(n19330), .A2(n19662), .B1(n19661), .B2(n19329), .ZN(
        n19317) );
  AOI22_X1 U22321 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19331), .B1(
        n19324), .B2(n19611), .ZN(n19316) );
  OAI211_X1 U22322 ( .C1(n19614), .C2(n19363), .A(n19317), .B(n19316), .ZN(
        P2_U3081) );
  AOI22_X1 U22323 ( .A1(n19330), .A2(n19668), .B1(n19667), .B2(n19329), .ZN(
        n19319) );
  AOI22_X1 U22324 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19331), .B1(
        n19349), .B2(n19669), .ZN(n19318) );
  OAI211_X1 U22325 ( .C1(n19672), .C2(n19334), .A(n19319), .B(n19318), .ZN(
        P2_U3082) );
  AOI22_X1 U22326 ( .A1(n19330), .A2(n19674), .B1(n19673), .B2(n19329), .ZN(
        n19321) );
  AOI22_X1 U22327 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19331), .B1(
        n19324), .B2(n19617), .ZN(n19320) );
  OAI211_X1 U22328 ( .C1(n19620), .C2(n19363), .A(n19321), .B(n19320), .ZN(
        P2_U3083) );
  AOI22_X1 U22329 ( .A1(n19330), .A2(n19680), .B1(n19679), .B2(n19329), .ZN(
        n19323) );
  AOI22_X1 U22330 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19331), .B1(
        n19324), .B2(n19621), .ZN(n19322) );
  OAI211_X1 U22331 ( .C1(n19624), .C2(n19363), .A(n19323), .B(n19322), .ZN(
        P2_U3084) );
  AOI22_X1 U22332 ( .A1(n19330), .A2(n19686), .B1(n19685), .B2(n19329), .ZN(
        n19326) );
  AOI22_X1 U22333 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19331), .B1(
        n19324), .B2(n19625), .ZN(n19325) );
  OAI211_X1 U22334 ( .C1(n19628), .C2(n19363), .A(n19326), .B(n19325), .ZN(
        P2_U3085) );
  AOI22_X1 U22335 ( .A1(n19330), .A2(n19692), .B1(n19691), .B2(n19329), .ZN(
        n19328) );
  AOI22_X1 U22336 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19331), .B1(
        n19349), .B2(n19693), .ZN(n19327) );
  OAI211_X1 U22337 ( .C1(n19696), .C2(n19334), .A(n19328), .B(n19327), .ZN(
        P2_U3086) );
  AOI22_X1 U22338 ( .A1(n19330), .A2(n19699), .B1(n19697), .B2(n19329), .ZN(
        n19333) );
  AOI22_X1 U22339 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19331), .B1(
        n19349), .B2(n19701), .ZN(n19332) );
  OAI211_X1 U22340 ( .C1(n19707), .C2(n19334), .A(n19333), .B(n19332), .ZN(
        P2_U3087) );
  NOR2_X1 U22341 ( .A1(n19447), .A2(n19387), .ZN(n19358) );
  AOI22_X1 U22342 ( .A1(n19575), .A2(n19349), .B1(n19645), .B2(n19358), .ZN(
        n19344) );
  OAI21_X1 U22343 ( .B1(n19391), .B2(n19568), .A(n19812), .ZN(n19342) );
  INV_X1 U22344 ( .A(n19335), .ZN(n19337) );
  INV_X1 U22345 ( .A(n19358), .ZN(n19336) );
  OAI211_X1 U22346 ( .C1(n19337), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19336), 
        .B(n19807), .ZN(n19338) );
  OAI211_X1 U22347 ( .C1(n19342), .C2(n19339), .A(n19604), .B(n19338), .ZN(
        n19360) );
  OAI21_X1 U22348 ( .B1(n19335), .B2(n19358), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19340) );
  OAI21_X1 U22349 ( .B1(n19342), .B2(n19341), .A(n19340), .ZN(n19359) );
  AOI22_X1 U22350 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19360), .B1(
        n19646), .B2(n19359), .ZN(n19343) );
  OAI211_X1 U22351 ( .C1(n19578), .C2(n19385), .A(n19344), .B(n19343), .ZN(
        P2_U3088) );
  AOI22_X1 U22352 ( .A1(n19611), .A2(n19349), .B1(n19358), .B2(n19661), .ZN(
        n19346) );
  AOI22_X1 U22353 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19360), .B1(
        n19662), .B2(n19359), .ZN(n19345) );
  OAI211_X1 U22354 ( .C1(n19614), .C2(n19385), .A(n19346), .B(n19345), .ZN(
        P2_U3089) );
  AOI22_X1 U22355 ( .A1(n19544), .A2(n19349), .B1(n19667), .B2(n19358), .ZN(
        n19348) );
  AOI22_X1 U22356 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19360), .B1(
        n19668), .B2(n19359), .ZN(n19347) );
  OAI211_X1 U22357 ( .C1(n19547), .C2(n19385), .A(n19348), .B(n19347), .ZN(
        P2_U3090) );
  AOI22_X1 U22358 ( .A1(n19617), .A2(n19349), .B1(n19358), .B2(n19673), .ZN(
        n19351) );
  AOI22_X1 U22359 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19360), .B1(
        n19674), .B2(n19359), .ZN(n19350) );
  OAI211_X1 U22360 ( .C1(n19620), .C2(n19385), .A(n19351), .B(n19350), .ZN(
        P2_U3091) );
  AOI22_X1 U22361 ( .A1(n19681), .A2(n19367), .B1(n19679), .B2(n19358), .ZN(
        n19353) );
  AOI22_X1 U22362 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19360), .B1(
        n19680), .B2(n19359), .ZN(n19352) );
  OAI211_X1 U22363 ( .C1(n19684), .C2(n19363), .A(n19353), .B(n19352), .ZN(
        P2_U3092) );
  AOI22_X1 U22364 ( .A1(n19687), .A2(n19367), .B1(n19358), .B2(n19685), .ZN(
        n19355) );
  AOI22_X1 U22365 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19360), .B1(
        n19686), .B2(n19359), .ZN(n19354) );
  OAI211_X1 U22366 ( .C1(n19690), .C2(n19363), .A(n19355), .B(n19354), .ZN(
        P2_U3093) );
  AOI22_X1 U22367 ( .A1(n19693), .A2(n19367), .B1(n19691), .B2(n19358), .ZN(
        n19357) );
  AOI22_X1 U22368 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19360), .B1(
        n19692), .B2(n19359), .ZN(n19356) );
  OAI211_X1 U22369 ( .C1(n19696), .C2(n19363), .A(n19357), .B(n19356), .ZN(
        P2_U3094) );
  AOI22_X1 U22370 ( .A1(n19701), .A2(n19367), .B1(n19358), .B2(n19697), .ZN(
        n19362) );
  AOI22_X1 U22371 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19360), .B1(
        n19699), .B2(n19359), .ZN(n19361) );
  OAI211_X1 U22372 ( .C1(n19707), .C2(n19363), .A(n19362), .B(n19361), .ZN(
        P2_U3095) );
  INV_X1 U22373 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n19366) );
  AOI22_X1 U22374 ( .A1(n19381), .A2(n19646), .B1(n19645), .B2(n19380), .ZN(
        n19365) );
  AOI22_X1 U22375 ( .A1(n19411), .A2(n19657), .B1(n19367), .B2(n19575), .ZN(
        n19364) );
  OAI211_X1 U22376 ( .C1(n19371), .C2(n19366), .A(n19365), .B(n19364), .ZN(
        P2_U3096) );
  INV_X1 U22377 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n19370) );
  AOI22_X1 U22378 ( .A1(n19381), .A2(n19662), .B1(n19380), .B2(n19661), .ZN(
        n19369) );
  AOI22_X1 U22379 ( .A1(n19411), .A2(n19663), .B1(n19367), .B2(n19611), .ZN(
        n19368) );
  OAI211_X1 U22380 ( .C1(n19371), .C2(n19370), .A(n19369), .B(n19368), .ZN(
        P2_U3097) );
  AOI22_X1 U22381 ( .A1(n19381), .A2(n19674), .B1(n19380), .B2(n19673), .ZN(
        n19373) );
  AOI22_X1 U22382 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19382), .B1(
        n19411), .B2(n19675), .ZN(n19372) );
  OAI211_X1 U22383 ( .C1(n19678), .C2(n19385), .A(n19373), .B(n19372), .ZN(
        P2_U3099) );
  AOI22_X1 U22384 ( .A1(n19381), .A2(n19680), .B1(n19380), .B2(n19679), .ZN(
        n19375) );
  AOI22_X1 U22385 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19382), .B1(
        n19411), .B2(n19681), .ZN(n19374) );
  OAI211_X1 U22386 ( .C1(n19684), .C2(n19385), .A(n19375), .B(n19374), .ZN(
        P2_U3100) );
  AOI22_X1 U22387 ( .A1(n19381), .A2(n19686), .B1(n19380), .B2(n19685), .ZN(
        n19377) );
  AOI22_X1 U22388 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19382), .B1(
        n19411), .B2(n19687), .ZN(n19376) );
  OAI211_X1 U22389 ( .C1(n19690), .C2(n19385), .A(n19377), .B(n19376), .ZN(
        P2_U3101) );
  AOI22_X1 U22390 ( .A1(n19381), .A2(n19692), .B1(n19380), .B2(n19691), .ZN(
        n19379) );
  AOI22_X1 U22391 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19382), .B1(
        n19411), .B2(n19693), .ZN(n19378) );
  OAI211_X1 U22392 ( .C1(n19696), .C2(n19385), .A(n19379), .B(n19378), .ZN(
        P2_U3102) );
  AOI22_X1 U22393 ( .A1(n19381), .A2(n19699), .B1(n19380), .B2(n19697), .ZN(
        n19384) );
  AOI22_X1 U22394 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19382), .B1(
        n19411), .B2(n19701), .ZN(n19383) );
  OAI211_X1 U22395 ( .C1(n19707), .C2(n19385), .A(n19384), .B(n19383), .ZN(
        P2_U3103) );
  NOR2_X1 U22396 ( .A1(n19641), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19394) );
  INV_X1 U22397 ( .A(n19394), .ZN(n19390) );
  NOR2_X1 U22398 ( .A1(n19510), .A2(n19387), .ZN(n19421) );
  NOR3_X1 U22399 ( .A1(n19388), .A2(n19421), .A3(n19852), .ZN(n19392) );
  AOI211_X2 U22400 ( .C1(n19390), .C2(n19852), .A(n19389), .B(n19392), .ZN(
        n19410) );
  AOI22_X1 U22401 ( .A1(n19410), .A2(n19646), .B1(n19645), .B2(n19421), .ZN(
        n19397) );
  OR2_X1 U22402 ( .A1(n19391), .A2(n19798), .ZN(n19808) );
  INV_X1 U22403 ( .A(n19808), .ZN(n19395) );
  INV_X1 U22404 ( .A(n19421), .ZN(n19418) );
  AOI211_X1 U22405 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19418), .A(n19650), 
        .B(n19392), .ZN(n19393) );
  OAI21_X1 U22406 ( .B1(n19395), .B2(n19394), .A(n19393), .ZN(n19412) );
  AOI22_X1 U22407 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19412), .B1(
        n19411), .B2(n19575), .ZN(n19396) );
  OAI211_X1 U22408 ( .C1(n19578), .C2(n19444), .A(n19397), .B(n19396), .ZN(
        P2_U3104) );
  AOI22_X1 U22409 ( .A1(n19410), .A2(n19662), .B1(n19421), .B2(n19661), .ZN(
        n19399) );
  AOI22_X1 U22410 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19412), .B1(
        n19411), .B2(n19611), .ZN(n19398) );
  OAI211_X1 U22411 ( .C1(n19614), .C2(n19444), .A(n19399), .B(n19398), .ZN(
        P2_U3105) );
  AOI22_X1 U22412 ( .A1(n19410), .A2(n19668), .B1(n19667), .B2(n19421), .ZN(
        n19401) );
  AOI22_X1 U22413 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19412), .B1(
        n19411), .B2(n19544), .ZN(n19400) );
  OAI211_X1 U22414 ( .C1(n19547), .C2(n19444), .A(n19401), .B(n19400), .ZN(
        P2_U3106) );
  AOI22_X1 U22415 ( .A1(n19410), .A2(n19674), .B1(n19421), .B2(n19673), .ZN(
        n19403) );
  AOI22_X1 U22416 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19412), .B1(
        n19411), .B2(n19617), .ZN(n19402) );
  OAI211_X1 U22417 ( .C1(n19620), .C2(n19444), .A(n19403), .B(n19402), .ZN(
        P2_U3107) );
  AOI22_X1 U22418 ( .A1(n19410), .A2(n19680), .B1(n19679), .B2(n19421), .ZN(
        n19405) );
  AOI22_X1 U22419 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19412), .B1(
        n19411), .B2(n19621), .ZN(n19404) );
  OAI211_X1 U22420 ( .C1(n19624), .C2(n19444), .A(n19405), .B(n19404), .ZN(
        P2_U3108) );
  AOI22_X1 U22421 ( .A1(n19410), .A2(n19686), .B1(n19421), .B2(n19685), .ZN(
        n19407) );
  AOI22_X1 U22422 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19412), .B1(
        n19411), .B2(n19625), .ZN(n19406) );
  OAI211_X1 U22423 ( .C1(n19628), .C2(n19444), .A(n19407), .B(n19406), .ZN(
        P2_U3109) );
  AOI22_X1 U22424 ( .A1(n19410), .A2(n19692), .B1(n19421), .B2(n19691), .ZN(
        n19409) );
  AOI22_X1 U22425 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19412), .B1(
        n19411), .B2(n19555), .ZN(n19408) );
  OAI211_X1 U22426 ( .C1(n19558), .C2(n19444), .A(n19409), .B(n19408), .ZN(
        P2_U3110) );
  AOI22_X1 U22427 ( .A1(n19410), .A2(n19699), .B1(n19421), .B2(n19697), .ZN(
        n19414) );
  AOI22_X1 U22428 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19412), .B1(
        n19411), .B2(n19635), .ZN(n19413) );
  OAI211_X1 U22429 ( .C1(n19640), .C2(n19444), .A(n19414), .B(n19413), .ZN(
        P2_U3111) );
  NOR2_X1 U22430 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19811), .ZN(
        n19512) );
  NAND2_X1 U22431 ( .A1(n19512), .A2(n19828), .ZN(n19455) );
  NOR2_X1 U22432 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19455), .ZN(
        n19439) );
  AOI22_X1 U22433 ( .A1(n19657), .A2(n19474), .B1(n19645), .B2(n19439), .ZN(
        n19426) );
  AOI21_X1 U22434 ( .B1(n19473), .B2(n19444), .A(n15620), .ZN(n19415) );
  NOR2_X1 U22435 ( .A1(n19415), .A2(n19807), .ZN(n19420) );
  OAI21_X1 U22436 ( .B1(n19422), .B2(n19852), .A(n19416), .ZN(n19417) );
  AOI21_X1 U22437 ( .B1(n19420), .B2(n19418), .A(n19417), .ZN(n19419) );
  OAI21_X1 U22438 ( .B1(n19421), .B2(n19439), .A(n19420), .ZN(n19424) );
  OAI21_X1 U22439 ( .B1(n19422), .B2(n19439), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19423) );
  AOI22_X1 U22440 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19441), .B1(
        n19646), .B2(n19440), .ZN(n19425) );
  OAI211_X1 U22441 ( .C1(n19660), .C2(n19444), .A(n19426), .B(n19425), .ZN(
        P2_U3112) );
  AOI22_X1 U22442 ( .A1(n19663), .A2(n19474), .B1(n19439), .B2(n19661), .ZN(
        n19428) );
  AOI22_X1 U22443 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19441), .B1(
        n19662), .B2(n19440), .ZN(n19427) );
  OAI211_X1 U22444 ( .C1(n19666), .C2(n19444), .A(n19428), .B(n19427), .ZN(
        P2_U3113) );
  AOI22_X1 U22445 ( .A1(n19669), .A2(n19474), .B1(n19667), .B2(n19439), .ZN(
        n19430) );
  AOI22_X1 U22446 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19441), .B1(
        n19668), .B2(n19440), .ZN(n19429) );
  OAI211_X1 U22447 ( .C1(n19672), .C2(n19444), .A(n19430), .B(n19429), .ZN(
        P2_U3114) );
  AOI22_X1 U22448 ( .A1(n19675), .A2(n19474), .B1(n19673), .B2(n19439), .ZN(
        n19432) );
  AOI22_X1 U22449 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19441), .B1(
        n19674), .B2(n19440), .ZN(n19431) );
  OAI211_X1 U22450 ( .C1(n19678), .C2(n19444), .A(n19432), .B(n19431), .ZN(
        P2_U3115) );
  AOI22_X1 U22451 ( .A1(n19681), .A2(n19474), .B1(n19679), .B2(n19439), .ZN(
        n19434) );
  AOI22_X1 U22452 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19441), .B1(
        n19680), .B2(n19440), .ZN(n19433) );
  OAI211_X1 U22453 ( .C1(n19684), .C2(n19444), .A(n19434), .B(n19433), .ZN(
        P2_U3116) );
  AOI22_X1 U22454 ( .A1(n19687), .A2(n19474), .B1(n19439), .B2(n19685), .ZN(
        n19436) );
  AOI22_X1 U22455 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19441), .B1(
        n19686), .B2(n19440), .ZN(n19435) );
  OAI211_X1 U22456 ( .C1(n19690), .C2(n19444), .A(n19436), .B(n19435), .ZN(
        P2_U3117) );
  AOI22_X1 U22457 ( .A1(n19693), .A2(n19474), .B1(n19691), .B2(n19439), .ZN(
        n19438) );
  AOI22_X1 U22458 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19441), .B1(
        n19692), .B2(n19440), .ZN(n19437) );
  OAI211_X1 U22459 ( .C1(n19696), .C2(n19444), .A(n19438), .B(n19437), .ZN(
        P2_U3118) );
  AOI22_X1 U22460 ( .A1(n19701), .A2(n19474), .B1(n19697), .B2(n19439), .ZN(
        n19443) );
  AOI22_X1 U22461 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19441), .B1(
        n19699), .B2(n19440), .ZN(n19442) );
  OAI211_X1 U22462 ( .C1(n19707), .C2(n19444), .A(n19443), .B(n19442), .ZN(
        P2_U3119) );
  OR2_X1 U22463 ( .A1(n19445), .A2(n15620), .ZN(n19647) );
  OAI21_X1 U22464 ( .B1(n19647), .B2(n19452), .A(n19812), .ZN(n19456) );
  INV_X1 U22465 ( .A(n19455), .ZN(n19446) );
  OR2_X1 U22466 ( .A1(n19456), .A2(n19446), .ZN(n19451) );
  INV_X1 U22467 ( .A(n19512), .ZN(n19515) );
  NOR2_X1 U22468 ( .A1(n19447), .A2(n19515), .ZN(n19483) );
  NOR2_X1 U22469 ( .A1(n19812), .A2(n19483), .ZN(n19449) );
  NAND2_X1 U22470 ( .A1(n19453), .A2(n19416), .ZN(n19448) );
  AOI21_X1 U22471 ( .B1(n19449), .B2(n19448), .A(n19650), .ZN(n19450) );
  INV_X1 U22472 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n19459) );
  AOI22_X1 U22473 ( .A1(n19657), .A2(n19482), .B1(n19645), .B2(n19483), .ZN(
        n19458) );
  OAI21_X1 U22474 ( .B1(n19453), .B2(n19483), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19454) );
  OAI21_X1 U22475 ( .B1(n19456), .B2(n19455), .A(n19454), .ZN(n19475) );
  AOI22_X1 U22476 ( .A1(n19646), .A2(n19475), .B1(n19474), .B2(n19575), .ZN(
        n19457) );
  OAI211_X1 U22477 ( .C1(n19460), .C2(n19459), .A(n19458), .B(n19457), .ZN(
        P2_U3120) );
  AOI22_X1 U22478 ( .A1(n19611), .A2(n19474), .B1(n19661), .B2(n19483), .ZN(
        n19462) );
  AOI22_X1 U22479 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19476), .B1(
        n19662), .B2(n19475), .ZN(n19461) );
  OAI211_X1 U22480 ( .C1(n19614), .C2(n19509), .A(n19462), .B(n19461), .ZN(
        P2_U3121) );
  AOI22_X1 U22481 ( .A1(n19669), .A2(n19482), .B1(n19667), .B2(n19483), .ZN(
        n19464) );
  AOI22_X1 U22482 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19476), .B1(
        n19668), .B2(n19475), .ZN(n19463) );
  OAI211_X1 U22483 ( .C1(n19672), .C2(n19473), .A(n19464), .B(n19463), .ZN(
        P2_U3122) );
  AOI22_X1 U22484 ( .A1(n19675), .A2(n19482), .B1(n19673), .B2(n19483), .ZN(
        n19466) );
  AOI22_X1 U22485 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19476), .B1(
        n19674), .B2(n19475), .ZN(n19465) );
  OAI211_X1 U22486 ( .C1(n19678), .C2(n19473), .A(n19466), .B(n19465), .ZN(
        P2_U3123) );
  AOI22_X1 U22487 ( .A1(n19681), .A2(n19482), .B1(n19679), .B2(n19483), .ZN(
        n19468) );
  AOI22_X1 U22488 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19476), .B1(
        n19680), .B2(n19475), .ZN(n19467) );
  OAI211_X1 U22489 ( .C1(n19684), .C2(n19473), .A(n19468), .B(n19467), .ZN(
        P2_U3124) );
  AOI22_X1 U22490 ( .A1(n19687), .A2(n19482), .B1(n19685), .B2(n19483), .ZN(
        n19470) );
  AOI22_X1 U22491 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19476), .B1(
        n19686), .B2(n19475), .ZN(n19469) );
  OAI211_X1 U22492 ( .C1(n19690), .C2(n19473), .A(n19470), .B(n19469), .ZN(
        P2_U3125) );
  AOI22_X1 U22493 ( .A1(n19693), .A2(n19482), .B1(n19691), .B2(n19483), .ZN(
        n19472) );
  AOI22_X1 U22494 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19476), .B1(
        n19692), .B2(n19475), .ZN(n19471) );
  OAI211_X1 U22495 ( .C1(n19696), .C2(n19473), .A(n19472), .B(n19471), .ZN(
        P2_U3126) );
  AOI22_X1 U22496 ( .A1(n19635), .A2(n19474), .B1(n19697), .B2(n19483), .ZN(
        n19478) );
  AOI22_X1 U22497 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19476), .B1(
        n19699), .B2(n19475), .ZN(n19477) );
  OAI211_X1 U22498 ( .C1(n19640), .C2(n19509), .A(n19478), .B(n19477), .ZN(
        P2_U3127) );
  NOR2_X1 U22499 ( .A1(n19479), .A2(n19515), .ZN(n19504) );
  OAI21_X1 U22500 ( .B1(n13287), .B2(n19504), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19480) );
  OAI21_X1 U22501 ( .B1(n19515), .B2(n19481), .A(n19480), .ZN(n19505) );
  AOI22_X1 U22502 ( .A1(n19505), .A2(n19646), .B1(n19645), .B2(n19504), .ZN(
        n19491) );
  OAI21_X1 U22503 ( .B1(n19537), .B2(n19482), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19485) );
  INV_X1 U22504 ( .A(n19483), .ZN(n19484) );
  AOI21_X1 U22505 ( .B1(n19485), .B2(n19484), .A(n19807), .ZN(n19489) );
  NAND3_X1 U22506 ( .A1(n13287), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19416), 
        .ZN(n19487) );
  INV_X1 U22507 ( .A(n19504), .ZN(n19486) );
  NAND2_X1 U22508 ( .A1(n19487), .A2(n19486), .ZN(n19488) );
  AOI22_X1 U22509 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19506), .B1(
        n19537), .B2(n19657), .ZN(n19490) );
  OAI211_X1 U22510 ( .C1(n19660), .C2(n19509), .A(n19491), .B(n19490), .ZN(
        P2_U3128) );
  AOI22_X1 U22511 ( .A1(n19505), .A2(n19662), .B1(n19661), .B2(n19504), .ZN(
        n19493) );
  AOI22_X1 U22512 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19506), .B1(
        n19537), .B2(n19663), .ZN(n19492) );
  OAI211_X1 U22513 ( .C1(n19666), .C2(n19509), .A(n19493), .B(n19492), .ZN(
        P2_U3129) );
  AOI22_X1 U22514 ( .A1(n19505), .A2(n19668), .B1(n19667), .B2(n19504), .ZN(
        n19495) );
  AOI22_X1 U22515 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19506), .B1(
        n19537), .B2(n19669), .ZN(n19494) );
  OAI211_X1 U22516 ( .C1(n19672), .C2(n19509), .A(n19495), .B(n19494), .ZN(
        P2_U3130) );
  AOI22_X1 U22517 ( .A1(n19505), .A2(n19674), .B1(n19673), .B2(n19504), .ZN(
        n19497) );
  AOI22_X1 U22518 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19506), .B1(
        n19537), .B2(n19675), .ZN(n19496) );
  OAI211_X1 U22519 ( .C1(n19678), .C2(n19509), .A(n19497), .B(n19496), .ZN(
        P2_U3131) );
  AOI22_X1 U22520 ( .A1(n19505), .A2(n19680), .B1(n19679), .B2(n19504), .ZN(
        n19499) );
  AOI22_X1 U22521 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19506), .B1(
        n19537), .B2(n19681), .ZN(n19498) );
  OAI211_X1 U22522 ( .C1(n19684), .C2(n19509), .A(n19499), .B(n19498), .ZN(
        P2_U3132) );
  AOI22_X1 U22523 ( .A1(n19505), .A2(n19686), .B1(n19685), .B2(n19504), .ZN(
        n19501) );
  AOI22_X1 U22524 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19506), .B1(
        n19537), .B2(n19687), .ZN(n19500) );
  OAI211_X1 U22525 ( .C1(n19690), .C2(n19509), .A(n19501), .B(n19500), .ZN(
        P2_U3133) );
  AOI22_X1 U22526 ( .A1(n19505), .A2(n19692), .B1(n19691), .B2(n19504), .ZN(
        n19503) );
  AOI22_X1 U22527 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19506), .B1(
        n19537), .B2(n19693), .ZN(n19502) );
  OAI211_X1 U22528 ( .C1(n19696), .C2(n19509), .A(n19503), .B(n19502), .ZN(
        P2_U3134) );
  AOI22_X1 U22529 ( .A1(n19505), .A2(n19699), .B1(n19697), .B2(n19504), .ZN(
        n19508) );
  AOI22_X1 U22530 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19506), .B1(
        n19537), .B2(n19701), .ZN(n19507) );
  OAI211_X1 U22531 ( .C1(n19707), .C2(n19509), .A(n19508), .B(n19507), .ZN(
        P2_U3135) );
  NAND2_X1 U22532 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19512), .ZN(
        n19514) );
  INV_X1 U22533 ( .A(n19510), .ZN(n19511) );
  NAND2_X1 U22534 ( .A1(n19512), .A2(n19511), .ZN(n19517) );
  INV_X1 U22535 ( .A(n19517), .ZN(n19535) );
  OAI21_X1 U22536 ( .B1(n13291), .B2(n19535), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19513) );
  OAI21_X1 U22537 ( .B1(n19514), .B2(n19807), .A(n19513), .ZN(n19536) );
  AOI22_X1 U22538 ( .A1(n19536), .A2(n19646), .B1(n19645), .B2(n19535), .ZN(
        n19522) );
  OAI22_X1 U22539 ( .A1(n19647), .A2(n19516), .B1(n19828), .B2(n19515), .ZN(
        n19520) );
  INV_X1 U22540 ( .A(n13291), .ZN(n19518) );
  OAI211_X1 U22541 ( .C1(n19518), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19517), 
        .B(n19807), .ZN(n19519) );
  NAND3_X1 U22542 ( .A1(n19520), .A2(n19604), .A3(n19519), .ZN(n19538) );
  AOI22_X1 U22543 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19538), .B1(
        n19537), .B2(n19575), .ZN(n19521) );
  OAI211_X1 U22544 ( .C1(n19578), .C2(n19552), .A(n19522), .B(n19521), .ZN(
        P2_U3136) );
  AOI22_X1 U22545 ( .A1(n19536), .A2(n19662), .B1(n19661), .B2(n19535), .ZN(
        n19524) );
  AOI22_X1 U22546 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19538), .B1(
        n19537), .B2(n19611), .ZN(n19523) );
  OAI211_X1 U22547 ( .C1(n19614), .C2(n19552), .A(n19524), .B(n19523), .ZN(
        P2_U3137) );
  AOI22_X1 U22548 ( .A1(n19536), .A2(n19668), .B1(n19667), .B2(n19535), .ZN(
        n19526) );
  AOI22_X1 U22549 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19538), .B1(
        n19537), .B2(n19544), .ZN(n19525) );
  OAI211_X1 U22550 ( .C1(n19547), .C2(n19552), .A(n19526), .B(n19525), .ZN(
        P2_U3138) );
  AOI22_X1 U22551 ( .A1(n19536), .A2(n19674), .B1(n19673), .B2(n19535), .ZN(
        n19528) );
  AOI22_X1 U22552 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19538), .B1(
        n19537), .B2(n19617), .ZN(n19527) );
  OAI211_X1 U22553 ( .C1(n19620), .C2(n19552), .A(n19528), .B(n19527), .ZN(
        P2_U3139) );
  AOI22_X1 U22554 ( .A1(n19536), .A2(n19680), .B1(n19679), .B2(n19535), .ZN(
        n19530) );
  AOI22_X1 U22555 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19538), .B1(
        n19537), .B2(n19621), .ZN(n19529) );
  OAI211_X1 U22556 ( .C1(n19624), .C2(n19552), .A(n19530), .B(n19529), .ZN(
        P2_U3140) );
  AOI22_X1 U22557 ( .A1(n19536), .A2(n19686), .B1(n19685), .B2(n19535), .ZN(
        n19532) );
  AOI22_X1 U22558 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19538), .B1(
        n19537), .B2(n19625), .ZN(n19531) );
  OAI211_X1 U22559 ( .C1(n19628), .C2(n19552), .A(n19532), .B(n19531), .ZN(
        P2_U3141) );
  AOI22_X1 U22560 ( .A1(n19536), .A2(n19692), .B1(n19691), .B2(n19535), .ZN(
        n19534) );
  AOI22_X1 U22561 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19538), .B1(
        n19537), .B2(n19555), .ZN(n19533) );
  OAI211_X1 U22562 ( .C1(n19558), .C2(n19552), .A(n19534), .B(n19533), .ZN(
        P2_U3142) );
  AOI22_X1 U22563 ( .A1(n19536), .A2(n19699), .B1(n19697), .B2(n19535), .ZN(
        n19540) );
  AOI22_X1 U22564 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19538), .B1(
        n19537), .B2(n19635), .ZN(n19539) );
  OAI211_X1 U22565 ( .C1(n19640), .C2(n19552), .A(n19540), .B(n19539), .ZN(
        P2_U3143) );
  AOI22_X1 U22566 ( .A1(n19560), .A2(n19662), .B1(n19661), .B2(n19559), .ZN(
        n19543) );
  AOI22_X1 U22567 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19562), .B1(
        n19593), .B2(n19663), .ZN(n19542) );
  OAI211_X1 U22568 ( .C1(n19666), .C2(n19552), .A(n19543), .B(n19542), .ZN(
        P2_U3145) );
  AOI22_X1 U22569 ( .A1(n19560), .A2(n19668), .B1(n19667), .B2(n19559), .ZN(
        n19546) );
  AOI22_X1 U22570 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19562), .B1(
        n19561), .B2(n19544), .ZN(n19545) );
  OAI211_X1 U22571 ( .C1(n19547), .C2(n19591), .A(n19546), .B(n19545), .ZN(
        P2_U3146) );
  AOI22_X1 U22572 ( .A1(n19560), .A2(n19674), .B1(n19673), .B2(n19559), .ZN(
        n19549) );
  AOI22_X1 U22573 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19562), .B1(
        n19593), .B2(n19675), .ZN(n19548) );
  OAI211_X1 U22574 ( .C1(n19678), .C2(n19552), .A(n19549), .B(n19548), .ZN(
        P2_U3147) );
  AOI22_X1 U22575 ( .A1(n19560), .A2(n19680), .B1(n19679), .B2(n19559), .ZN(
        n19551) );
  AOI22_X1 U22576 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19562), .B1(
        n19593), .B2(n19681), .ZN(n19550) );
  OAI211_X1 U22577 ( .C1(n19684), .C2(n19552), .A(n19551), .B(n19550), .ZN(
        P2_U3148) );
  AOI22_X1 U22578 ( .A1(n19560), .A2(n19686), .B1(n19685), .B2(n19559), .ZN(
        n19554) );
  AOI22_X1 U22579 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19562), .B1(
        n19561), .B2(n19625), .ZN(n19553) );
  OAI211_X1 U22580 ( .C1(n19628), .C2(n19591), .A(n19554), .B(n19553), .ZN(
        P2_U3149) );
  AOI22_X1 U22581 ( .A1(n19560), .A2(n19692), .B1(n19691), .B2(n19559), .ZN(
        n19557) );
  AOI22_X1 U22582 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19562), .B1(
        n19561), .B2(n19555), .ZN(n19556) );
  OAI211_X1 U22583 ( .C1(n19558), .C2(n19591), .A(n19557), .B(n19556), .ZN(
        P2_U3150) );
  AOI22_X1 U22584 ( .A1(n19560), .A2(n19699), .B1(n19697), .B2(n19559), .ZN(
        n19564) );
  AOI22_X1 U22585 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19562), .B1(
        n19561), .B2(n19635), .ZN(n19563) );
  OAI211_X1 U22586 ( .C1(n19640), .C2(n19591), .A(n19564), .B(n19563), .ZN(
        P2_U3151) );
  INV_X1 U22587 ( .A(n19573), .ZN(n19567) );
  NOR2_X1 U22588 ( .A1(n19839), .A2(n19567), .ZN(n19600) );
  OAI21_X1 U22589 ( .B1(n19569), .B2(n19600), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19566) );
  OAI21_X1 U22590 ( .B1(n19567), .B2(n19807), .A(n19566), .ZN(n19592) );
  AOI22_X1 U22591 ( .A1(n19592), .A2(n19646), .B1(n19645), .B2(n19600), .ZN(
        n19577) );
  NOR2_X1 U22592 ( .A1(n19647), .A2(n19568), .ZN(n19574) );
  INV_X1 U22593 ( .A(n19569), .ZN(n19571) );
  INV_X1 U22594 ( .A(n19600), .ZN(n19570) );
  OAI211_X1 U22595 ( .C1(n19571), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19570), 
        .B(n19807), .ZN(n19572) );
  OAI211_X1 U22596 ( .C1(n19574), .C2(n19573), .A(n19604), .B(n19572), .ZN(
        n19594) );
  AOI22_X1 U22597 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19594), .B1(
        n19593), .B2(n19575), .ZN(n19576) );
  OAI211_X1 U22598 ( .C1(n19578), .C2(n19632), .A(n19577), .B(n19576), .ZN(
        P2_U3152) );
  AOI22_X1 U22599 ( .A1(n19592), .A2(n19662), .B1(n19661), .B2(n19600), .ZN(
        n19580) );
  AOI22_X1 U22600 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19594), .B1(
        n19634), .B2(n19663), .ZN(n19579) );
  OAI211_X1 U22601 ( .C1(n19666), .C2(n19591), .A(n19580), .B(n19579), .ZN(
        P2_U3153) );
  AOI22_X1 U22602 ( .A1(n19592), .A2(n19668), .B1(n19667), .B2(n19600), .ZN(
        n19582) );
  AOI22_X1 U22603 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19594), .B1(
        n19634), .B2(n19669), .ZN(n19581) );
  OAI211_X1 U22604 ( .C1(n19672), .C2(n19591), .A(n19582), .B(n19581), .ZN(
        P2_U3154) );
  AOI22_X1 U22605 ( .A1(n19592), .A2(n19674), .B1(n19673), .B2(n19600), .ZN(
        n19584) );
  AOI22_X1 U22606 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19594), .B1(
        n19634), .B2(n19675), .ZN(n19583) );
  OAI211_X1 U22607 ( .C1(n19678), .C2(n19591), .A(n19584), .B(n19583), .ZN(
        P2_U3155) );
  AOI22_X1 U22608 ( .A1(n19592), .A2(n19680), .B1(n19679), .B2(n19600), .ZN(
        n19586) );
  AOI22_X1 U22609 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19594), .B1(
        n19593), .B2(n19621), .ZN(n19585) );
  OAI211_X1 U22610 ( .C1(n19624), .C2(n19632), .A(n19586), .B(n19585), .ZN(
        P2_U3156) );
  AOI22_X1 U22611 ( .A1(n19592), .A2(n19686), .B1(n19685), .B2(n19600), .ZN(
        n19588) );
  AOI22_X1 U22612 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19594), .B1(
        n19593), .B2(n19625), .ZN(n19587) );
  OAI211_X1 U22613 ( .C1(n19628), .C2(n19632), .A(n19588), .B(n19587), .ZN(
        P2_U3157) );
  AOI22_X1 U22614 ( .A1(n19592), .A2(n19692), .B1(n19691), .B2(n19600), .ZN(
        n19590) );
  AOI22_X1 U22615 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19594), .B1(
        n19634), .B2(n19693), .ZN(n19589) );
  OAI211_X1 U22616 ( .C1(n19696), .C2(n19591), .A(n19590), .B(n19589), .ZN(
        P2_U3158) );
  AOI22_X1 U22617 ( .A1(n19592), .A2(n19699), .B1(n19697), .B2(n19600), .ZN(
        n19596) );
  AOI22_X1 U22618 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19594), .B1(
        n19593), .B2(n19635), .ZN(n19595) );
  OAI211_X1 U22619 ( .C1(n19640), .C2(n19632), .A(n19596), .B(n19595), .ZN(
        P2_U3159) );
  NOR3_X2 U22620 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19811), .A3(
        n19641), .ZN(n19633) );
  AOI22_X1 U22621 ( .A1(n19657), .A2(n19629), .B1(n19645), .B2(n19633), .ZN(
        n19610) );
  NOR3_X1 U22622 ( .A1(n19634), .A2(n19629), .A3(n19807), .ZN(n19599) );
  INV_X1 U22623 ( .A(n19800), .ZN(n19598) );
  NOR2_X1 U22624 ( .A1(n19599), .A2(n19598), .ZN(n19608) );
  NOR2_X1 U22625 ( .A1(n19633), .A2(n19600), .ZN(n19607) );
  INV_X1 U22626 ( .A(n19607), .ZN(n19605) );
  INV_X1 U22627 ( .A(n13545), .ZN(n19602) );
  INV_X1 U22628 ( .A(n19633), .ZN(n19601) );
  OAI211_X1 U22629 ( .C1(n19602), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19601), 
        .B(n19807), .ZN(n19603) );
  OAI211_X1 U22630 ( .C1(n19608), .C2(n19605), .A(n19604), .B(n19603), .ZN(
        n19637) );
  OAI21_X1 U22631 ( .B1(n13545), .B2(n19633), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19606) );
  AOI22_X1 U22632 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19637), .B1(
        n19646), .B2(n19636), .ZN(n19609) );
  OAI211_X1 U22633 ( .C1(n19660), .C2(n19632), .A(n19610), .B(n19609), .ZN(
        P2_U3160) );
  AOI22_X1 U22634 ( .A1(n19611), .A2(n19634), .B1(n19633), .B2(n19661), .ZN(
        n19613) );
  AOI22_X1 U22635 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19637), .B1(
        n19662), .B2(n19636), .ZN(n19612) );
  OAI211_X1 U22636 ( .C1(n19614), .C2(n19706), .A(n19613), .B(n19612), .ZN(
        P2_U3161) );
  AOI22_X1 U22637 ( .A1(n19669), .A2(n19629), .B1(n19667), .B2(n19633), .ZN(
        n19616) );
  AOI22_X1 U22638 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19637), .B1(
        n19668), .B2(n19636), .ZN(n19615) );
  OAI211_X1 U22639 ( .C1(n19672), .C2(n19632), .A(n19616), .B(n19615), .ZN(
        P2_U3162) );
  AOI22_X1 U22640 ( .A1(n19617), .A2(n19634), .B1(n19673), .B2(n19633), .ZN(
        n19619) );
  AOI22_X1 U22641 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19637), .B1(
        n19674), .B2(n19636), .ZN(n19618) );
  OAI211_X1 U22642 ( .C1(n19620), .C2(n19706), .A(n19619), .B(n19618), .ZN(
        P2_U3163) );
  AOI22_X1 U22643 ( .A1(n19621), .A2(n19634), .B1(n19679), .B2(n19633), .ZN(
        n19623) );
  AOI22_X1 U22644 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19637), .B1(
        n19680), .B2(n19636), .ZN(n19622) );
  OAI211_X1 U22645 ( .C1(n19624), .C2(n19706), .A(n19623), .B(n19622), .ZN(
        P2_U3164) );
  AOI22_X1 U22646 ( .A1(n19625), .A2(n19634), .B1(n19633), .B2(n19685), .ZN(
        n19627) );
  AOI22_X1 U22647 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19637), .B1(
        n19686), .B2(n19636), .ZN(n19626) );
  OAI211_X1 U22648 ( .C1(n19628), .C2(n19706), .A(n19627), .B(n19626), .ZN(
        P2_U3165) );
  AOI22_X1 U22649 ( .A1(n19693), .A2(n19629), .B1(n19691), .B2(n19633), .ZN(
        n19631) );
  AOI22_X1 U22650 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19637), .B1(
        n19692), .B2(n19636), .ZN(n19630) );
  OAI211_X1 U22651 ( .C1(n19696), .C2(n19632), .A(n19631), .B(n19630), .ZN(
        P2_U3166) );
  AOI22_X1 U22652 ( .A1(n19635), .A2(n19634), .B1(n19633), .B2(n19697), .ZN(
        n19639) );
  AOI22_X1 U22653 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19637), .B1(
        n19699), .B2(n19636), .ZN(n19638) );
  OAI211_X1 U22654 ( .C1(n19640), .C2(n19706), .A(n19639), .B(n19638), .ZN(
        P2_U3167) );
  NOR2_X1 U22655 ( .A1(n19811), .A2(n19641), .ZN(n19656) );
  INV_X1 U22656 ( .A(n19656), .ZN(n19642) );
  OR2_X1 U22657 ( .A1(n19642), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19644) );
  NAND2_X1 U22658 ( .A1(n19648), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19643) );
  NOR2_X1 U22659 ( .A1(n13296), .A2(n19643), .ZN(n19652) );
  AOI21_X1 U22660 ( .B1(n19852), .B2(n19644), .A(n19652), .ZN(n19700) );
  INV_X1 U22661 ( .A(n19648), .ZN(n19698) );
  AOI22_X1 U22662 ( .A1(n19700), .A2(n19646), .B1(n19698), .B2(n19645), .ZN(
        n19659) );
  INV_X1 U22663 ( .A(n19798), .ZN(n19655) );
  INV_X1 U22664 ( .A(n19647), .ZN(n19654) );
  AND2_X1 U22665 ( .A1(n19648), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19649) );
  OR2_X1 U22666 ( .A1(n19650), .A2(n19649), .ZN(n19651) );
  NOR2_X1 U22667 ( .A1(n19652), .A2(n19651), .ZN(n19653) );
  OAI221_X1 U22668 ( .B1(n19656), .B2(n19655), .C1(n19656), .C2(n19654), .A(
        n19653), .ZN(n19703) );
  AOI22_X1 U22669 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19703), .B1(
        n19702), .B2(n19657), .ZN(n19658) );
  OAI211_X1 U22670 ( .C1(n19660), .C2(n19706), .A(n19659), .B(n19658), .ZN(
        P2_U3168) );
  AOI22_X1 U22671 ( .A1(n19700), .A2(n19662), .B1(n19698), .B2(n19661), .ZN(
        n19665) );
  AOI22_X1 U22672 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19703), .B1(
        n19702), .B2(n19663), .ZN(n19664) );
  OAI211_X1 U22673 ( .C1(n19666), .C2(n19706), .A(n19665), .B(n19664), .ZN(
        P2_U3169) );
  AOI22_X1 U22674 ( .A1(n19700), .A2(n19668), .B1(n19698), .B2(n19667), .ZN(
        n19671) );
  AOI22_X1 U22675 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19703), .B1(
        n19702), .B2(n19669), .ZN(n19670) );
  OAI211_X1 U22676 ( .C1(n19672), .C2(n19706), .A(n19671), .B(n19670), .ZN(
        P2_U3170) );
  AOI22_X1 U22677 ( .A1(n19700), .A2(n19674), .B1(n19698), .B2(n19673), .ZN(
        n19677) );
  AOI22_X1 U22678 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19703), .B1(
        n19702), .B2(n19675), .ZN(n19676) );
  OAI211_X1 U22679 ( .C1(n19678), .C2(n19706), .A(n19677), .B(n19676), .ZN(
        P2_U3171) );
  AOI22_X1 U22680 ( .A1(n19700), .A2(n19680), .B1(n19698), .B2(n19679), .ZN(
        n19683) );
  AOI22_X1 U22681 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19703), .B1(
        n19702), .B2(n19681), .ZN(n19682) );
  OAI211_X1 U22682 ( .C1(n19684), .C2(n19706), .A(n19683), .B(n19682), .ZN(
        P2_U3172) );
  AOI22_X1 U22683 ( .A1(n19700), .A2(n19686), .B1(n19698), .B2(n19685), .ZN(
        n19689) );
  AOI22_X1 U22684 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19703), .B1(
        n19702), .B2(n19687), .ZN(n19688) );
  OAI211_X1 U22685 ( .C1(n19690), .C2(n19706), .A(n19689), .B(n19688), .ZN(
        P2_U3173) );
  AOI22_X1 U22686 ( .A1(n19700), .A2(n19692), .B1(n19698), .B2(n19691), .ZN(
        n19695) );
  AOI22_X1 U22687 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19703), .B1(
        n19702), .B2(n19693), .ZN(n19694) );
  OAI211_X1 U22688 ( .C1(n19696), .C2(n19706), .A(n19695), .B(n19694), .ZN(
        P2_U3174) );
  AOI22_X1 U22689 ( .A1(n19700), .A2(n19699), .B1(n19698), .B2(n19697), .ZN(
        n19705) );
  AOI22_X1 U22690 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19703), .B1(
        n19702), .B2(n19701), .ZN(n19704) );
  OAI211_X1 U22691 ( .C1(n19707), .C2(n19706), .A(n19705), .B(n19704), .ZN(
        P2_U3175) );
  AOI21_X1 U22692 ( .B1(n19710), .B2(n19709), .A(n19708), .ZN(n19714) );
  OAI211_X1 U22693 ( .C1(n19715), .C2(n19711), .A(n19717), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19712) );
  OAI211_X1 U22694 ( .C1(n19715), .C2(n19714), .A(n19713), .B(n19712), .ZN(
        P2_U3177) );
  AND2_X1 U22695 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19716), .ZN(
        P2_U3179) );
  AND2_X1 U22696 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19716), .ZN(
        P2_U3180) );
  AND2_X1 U22697 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19716), .ZN(
        P2_U3181) );
  AND2_X1 U22698 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19716), .ZN(
        P2_U3182) );
  AND2_X1 U22699 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19716), .ZN(
        P2_U3183) );
  AND2_X1 U22700 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19716), .ZN(
        P2_U3184) );
  AND2_X1 U22701 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19716), .ZN(
        P2_U3185) );
  AND2_X1 U22702 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19716), .ZN(
        P2_U3186) );
  AND2_X1 U22703 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19716), .ZN(
        P2_U3187) );
  AND2_X1 U22704 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19716), .ZN(
        P2_U3188) );
  AND2_X1 U22705 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19716), .ZN(
        P2_U3189) );
  AND2_X1 U22706 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19716), .ZN(
        P2_U3190) );
  AND2_X1 U22707 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19716), .ZN(
        P2_U3191) );
  AND2_X1 U22708 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19716), .ZN(
        P2_U3192) );
  AND2_X1 U22709 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19716), .ZN(
        P2_U3193) );
  AND2_X1 U22710 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19716), .ZN(
        P2_U3194) );
  AND2_X1 U22711 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19716), .ZN(
        P2_U3195) );
  AND2_X1 U22712 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19716), .ZN(
        P2_U3196) );
  AND2_X1 U22713 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19716), .ZN(
        P2_U3197) );
  AND2_X1 U22714 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19716), .ZN(
        P2_U3198) );
  AND2_X1 U22715 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19716), .ZN(
        P2_U3199) );
  INV_X1 U22716 ( .A(P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20895) );
  NOR2_X1 U22717 ( .A1(n20895), .A2(n19797), .ZN(P2_U3200) );
  AND2_X1 U22718 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19716), .ZN(P2_U3201) );
  AND2_X1 U22719 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19716), .ZN(P2_U3202) );
  AND2_X1 U22720 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19716), .ZN(P2_U3203) );
  AND2_X1 U22721 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19716), .ZN(P2_U3204) );
  AND2_X1 U22722 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19716), .ZN(P2_U3205) );
  AND2_X1 U22723 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19716), .ZN(P2_U3206) );
  AND2_X1 U22724 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19716), .ZN(P2_U3207) );
  AND2_X1 U22725 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19716), .ZN(P2_U3208) );
  INV_X1 U22726 ( .A(NA), .ZN(n20663) );
  OAI21_X1 U22727 ( .B1(n20663), .B2(n19722), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19732) );
  INV_X1 U22728 ( .A(n19732), .ZN(n19720) );
  NAND2_X1 U22729 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19717), .ZN(n19730) );
  INV_X1 U22730 ( .A(n19730), .ZN(n19726) );
  INV_X1 U22731 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19871) );
  NOR3_X1 U22732 ( .A1(n19726), .A2(n19871), .A3(n19721), .ZN(n19719) );
  OAI211_X1 U22733 ( .C1(HOLD), .C2(n19871), .A(n19872), .B(n19727), .ZN(
        n19718) );
  OAI21_X1 U22734 ( .B1(n19720), .B2(n19719), .A(n19718), .ZN(P2_U3209) );
  NOR2_X1 U22735 ( .A1(HOLD), .A2(n19721), .ZN(n19731) );
  AOI21_X1 U22736 ( .B1(n19733), .B2(n19722), .A(n19731), .ZN(n19724) );
  OAI22_X1 U22737 ( .A1(n19724), .A2(n19871), .B1(n20668), .B2(n19723), .ZN(
        n19725) );
  OR3_X1 U22738 ( .A1(n19866), .A2(n19726), .A3(n19725), .ZN(P2_U3210) );
  OAI22_X1 U22739 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19727), .B1(NA), 
        .B2(n19730), .ZN(n19728) );
  OAI211_X1 U22740 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19728), .ZN(n19729) );
  OAI221_X1 U22741 ( .B1(n19732), .B2(n19731), .C1(n19732), .C2(n19730), .A(
        n19729), .ZN(P2_U3211) );
  OAI222_X1 U22742 ( .A1(n19787), .A2(n19736), .B1(n19735), .B2(n19780), .C1(
        n19734), .C2(n19784), .ZN(P2_U3212) );
  OAI222_X1 U22743 ( .A1(n19787), .A2(n13370), .B1(n19737), .B2(n19780), .C1(
        n19736), .C2(n19784), .ZN(P2_U3213) );
  INV_X1 U22744 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n20899) );
  OAI222_X1 U22745 ( .A1(n19787), .A2(n20899), .B1(n19738), .B2(n19780), .C1(
        n13370), .C2(n19784), .ZN(P2_U3214) );
  OAI222_X1 U22746 ( .A1(n19787), .A2(n13582), .B1(n19739), .B2(n19780), .C1(
        n20899), .C2(n19784), .ZN(P2_U3215) );
  OAI222_X1 U22747 ( .A1(n19787), .A2(n19741), .B1(n19740), .B2(n19780), .C1(
        n13582), .C2(n19784), .ZN(P2_U3216) );
  OAI222_X1 U22748 ( .A1(n19787), .A2(n19743), .B1(n19742), .B2(n19780), .C1(
        n19741), .C2(n19784), .ZN(P2_U3217) );
  OAI222_X1 U22749 ( .A1(n19787), .A2(n19745), .B1(n19744), .B2(n19780), .C1(
        n19743), .C2(n19784), .ZN(P2_U3218) );
  OAI222_X1 U22750 ( .A1(n19787), .A2(n19747), .B1(n19746), .B2(n19780), .C1(
        n19745), .C2(n19784), .ZN(P2_U3219) );
  OAI222_X1 U22751 ( .A1(n19787), .A2(n19749), .B1(n19748), .B2(n19780), .C1(
        n19747), .C2(n19784), .ZN(P2_U3220) );
  OAI222_X1 U22752 ( .A1(n19787), .A2(n15520), .B1(n19750), .B2(n19780), .C1(
        n19749), .C2(n19784), .ZN(P2_U3221) );
  OAI222_X1 U22753 ( .A1(n19787), .A2(n19752), .B1(n19751), .B2(n19780), .C1(
        n15520), .C2(n19784), .ZN(P2_U3222) );
  INV_X1 U22754 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n19754) );
  OAI222_X1 U22755 ( .A1(n19787), .A2(n19754), .B1(n19753), .B2(n19780), .C1(
        n19752), .C2(n19784), .ZN(P2_U3223) );
  OAI222_X1 U22756 ( .A1(n19787), .A2(n19756), .B1(n19755), .B2(n19780), .C1(
        n19754), .C2(n19784), .ZN(P2_U3224) );
  OAI222_X1 U22757 ( .A1(n19787), .A2(n15266), .B1(n19757), .B2(n19780), .C1(
        n19756), .C2(n19784), .ZN(P2_U3225) );
  INV_X1 U22758 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20814) );
  OAI222_X1 U22759 ( .A1(n19787), .A2(n20814), .B1(n19758), .B2(n19780), .C1(
        n15266), .C2(n19784), .ZN(P2_U3226) );
  INV_X1 U22760 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19760) );
  OAI222_X1 U22761 ( .A1(n19787), .A2(n19760), .B1(n19759), .B2(n19780), .C1(
        n20814), .C2(n19784), .ZN(P2_U3227) );
  INV_X1 U22762 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19762) );
  OAI222_X1 U22763 ( .A1(n19787), .A2(n19762), .B1(n19761), .B2(n19780), .C1(
        n19760), .C2(n19784), .ZN(P2_U3228) );
  OAI222_X1 U22764 ( .A1(n19787), .A2(n19764), .B1(n19763), .B2(n19780), .C1(
        n19762), .C2(n19784), .ZN(P2_U3229) );
  INV_X1 U22765 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19766) );
  OAI222_X1 U22766 ( .A1(n19787), .A2(n19766), .B1(n19765), .B2(n19780), .C1(
        n19764), .C2(n19784), .ZN(P2_U3230) );
  OAI222_X1 U22767 ( .A1(n19787), .A2(n19767), .B1(n20892), .B2(n19780), .C1(
        n19766), .C2(n19784), .ZN(P2_U3231) );
  INV_X1 U22768 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19769) );
  OAI222_X1 U22769 ( .A1(n19787), .A2(n19769), .B1(n19768), .B2(n19780), .C1(
        n19767), .C2(n19784), .ZN(P2_U3232) );
  OAI222_X1 U22770 ( .A1(n19787), .A2(n20860), .B1(n19770), .B2(n19780), .C1(
        n19769), .C2(n19784), .ZN(P2_U3233) );
  OAI222_X1 U22771 ( .A1(n19787), .A2(n19772), .B1(n19771), .B2(n19780), .C1(
        n20860), .C2(n19784), .ZN(P2_U3234) );
  OAI222_X1 U22772 ( .A1(n19787), .A2(n19774), .B1(n19773), .B2(n19780), .C1(
        n19772), .C2(n19784), .ZN(P2_U3235) );
  OAI222_X1 U22773 ( .A1(n19787), .A2(n15161), .B1(n19775), .B2(n19780), .C1(
        n19774), .C2(n19784), .ZN(P2_U3236) );
  OAI222_X1 U22774 ( .A1(n19787), .A2(n19778), .B1(n19776), .B2(n19780), .C1(
        n15161), .C2(n19784), .ZN(P2_U3237) );
  OAI222_X1 U22775 ( .A1(n19784), .A2(n19778), .B1(n19777), .B2(n19780), .C1(
        n19779), .C2(n19787), .ZN(P2_U3238) );
  OAI222_X1 U22776 ( .A1(n19787), .A2(n19782), .B1(n19781), .B2(n19780), .C1(
        n19779), .C2(n19784), .ZN(P2_U3239) );
  OAI222_X1 U22777 ( .A1(n19787), .A2(n13951), .B1(n19783), .B2(n19780), .C1(
        n19782), .C2(n19784), .ZN(P2_U3240) );
  OAI222_X1 U22778 ( .A1(n19787), .A2(n19786), .B1(n19785), .B2(n19780), .C1(
        n13951), .C2(n19784), .ZN(P2_U3241) );
  INV_X1 U22779 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19788) );
  AOI22_X1 U22780 ( .A1(n19780), .A2(n19789), .B1(n19788), .B2(n19872), .ZN(
        P2_U3585) );
  MUX2_X1 U22781 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n19780), .Z(P2_U3586) );
  INV_X1 U22782 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n19790) );
  AOI22_X1 U22783 ( .A1(n19780), .A2(n19791), .B1(n19790), .B2(n19872), .ZN(
        P2_U3587) );
  INV_X1 U22784 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n19792) );
  AOI22_X1 U22785 ( .A1(n19780), .A2(n19793), .B1(n19792), .B2(n19872), .ZN(
        P2_U3588) );
  OAI21_X1 U22786 ( .B1(n19797), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19795), 
        .ZN(n19794) );
  INV_X1 U22787 ( .A(n19794), .ZN(P2_U3591) );
  OAI21_X1 U22788 ( .B1(n19797), .B2(n19796), .A(n19795), .ZN(P2_U3592) );
  NAND2_X1 U22789 ( .A1(n19798), .A2(n19812), .ZN(n19802) );
  AND2_X1 U22790 ( .A1(n19800), .A2(n19799), .ZN(n19801) );
  NAND2_X1 U22791 ( .A1(n19802), .A2(n19801), .ZN(n19816) );
  NAND2_X1 U22792 ( .A1(n19816), .A2(n19803), .ZN(n19806) );
  NAND2_X1 U22793 ( .A1(n19804), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19805) );
  OAI211_X1 U22794 ( .C1(n19808), .C2(n19807), .A(n19806), .B(n19805), .ZN(
        n19809) );
  INV_X1 U22795 ( .A(n19809), .ZN(n19810) );
  AOI22_X1 U22796 ( .A1(n19837), .A2(n19811), .B1(n19810), .B2(n19838), .ZN(
        P2_U3602) );
  NAND2_X1 U22797 ( .A1(n19812), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19823) );
  OAI21_X1 U22798 ( .B1(n19814), .B2(n19823), .A(n19813), .ZN(n19815) );
  AOI22_X1 U22799 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19817), .B1(n19816), 
        .B2(n19815), .ZN(n19818) );
  AOI22_X1 U22800 ( .A1(n19837), .A2(n19819), .B1(n19818), .B2(n19838), .ZN(
        P2_U3603) );
  INV_X1 U22801 ( .A(n19820), .ZN(n19821) );
  NAND3_X1 U22802 ( .A1(n19824), .A2(n19829), .A3(n19821), .ZN(n19822) );
  OAI21_X1 U22803 ( .B1(n19824), .B2(n19823), .A(n19822), .ZN(n19825) );
  AOI21_X1 U22804 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19826), .A(n19825), 
        .ZN(n19827) );
  AOI22_X1 U22805 ( .A1(n19837), .A2(n19828), .B1(n19827), .B2(n19838), .ZN(
        P2_U3604) );
  INV_X1 U22806 ( .A(n19829), .ZN(n19833) );
  INV_X1 U22807 ( .A(n19830), .ZN(n19832) );
  OAI22_X1 U22808 ( .A1(n19834), .A2(n19833), .B1(n19832), .B2(n19831), .ZN(
        n19835) );
  AOI21_X1 U22809 ( .B1(n19839), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19835), 
        .ZN(n19836) );
  OAI22_X1 U22810 ( .A1(n19839), .A2(n19838), .B1(n19837), .B2(n19836), .ZN(
        P2_U3605) );
  INV_X1 U22811 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19840) );
  AOI22_X1 U22812 ( .A1(n19780), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19840), 
        .B2(n19872), .ZN(P2_U3608) );
  INV_X1 U22813 ( .A(n19841), .ZN(n19845) );
  INV_X1 U22814 ( .A(n19842), .ZN(n19843) );
  OAI21_X1 U22815 ( .B1(n19845), .B2(n19844), .A(n19843), .ZN(n19846) );
  OAI211_X1 U22816 ( .C1(n19849), .C2(n19848), .A(n19847), .B(n19846), .ZN(
        n19851) );
  MUX2_X1 U22817 ( .A(P2_MORE_REG_SCAN_IN), .B(n19851), .S(n19850), .Z(
        P2_U3609) );
  NOR2_X1 U22818 ( .A1(n19853), .A2(n19852), .ZN(n19854) );
  NOR2_X1 U22819 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19854), .ZN(n19857) );
  INV_X1 U22820 ( .A(n19855), .ZN(n19856) );
  AOI211_X1 U22821 ( .C1(n19858), .C2(n19859), .A(n19857), .B(n19856), .ZN(
        n19870) );
  NAND2_X1 U22822 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19859), .ZN(n19862) );
  NOR4_X1 U22823 ( .A1(n19860), .A2(n11798), .A3(n19866), .A4(n11587), .ZN(
        n19861) );
  AOI21_X1 U22824 ( .B1(n19863), .B2(n19862), .A(n19861), .ZN(n19869) );
  AOI211_X1 U22825 ( .C1(P2_STATEBS16_REG_SCAN_IN), .C2(n19866), .A(n19865), 
        .B(n19864), .ZN(n19867) );
  NOR2_X1 U22826 ( .A1(n19870), .A2(n19867), .ZN(n19868) );
  AOI22_X1 U22827 ( .A1(n19871), .A2(n19870), .B1(n19869), .B2(n19868), .ZN(
        P2_U3610) );
  INV_X1 U22828 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n19873) );
  AOI22_X1 U22829 ( .A1(n19780), .A2(n19874), .B1(n19873), .B2(n19872), .ZN(
        P2_U3611) );
  INV_X1 U22830 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n19875) );
  OAI21_X1 U22831 ( .B1(n19875), .B2(P1_STATE_REG_2__SCAN_IN), .A(
        P1_STATE_REG_0__SCAN_IN), .ZN(n19883) );
  OR2_X1 U22832 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n19875), .ZN(n20753) );
  OAI21_X1 U22833 ( .B1(n19883), .B2(P1_ADS_N_REG_SCAN_IN), .A(n20753), .ZN(
        n19876) );
  INV_X1 U22834 ( .A(n19876), .ZN(P1_U2802) );
  NAND2_X1 U22835 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n19877), .ZN(n19881) );
  OAI21_X1 U22836 ( .B1(n19879), .B2(n19878), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19880) );
  OAI21_X1 U22837 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n19881), .A(n19880), 
        .ZN(P1_U2803) );
  NOR2_X1 U22838 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19884) );
  OAI21_X1 U22839 ( .B1(n19884), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20753), .ZN(
        n19882) );
  OAI21_X1 U22840 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20753), .A(n19882), 
        .ZN(P1_U2804) );
  AND2_X1 U22841 ( .A1(n20753), .A2(n19883), .ZN(n20733) );
  OAI21_X1 U22842 ( .B1(BS16), .B2(n19884), .A(n20733), .ZN(n20731) );
  OAI21_X1 U22843 ( .B1(n20733), .B2(n20515), .A(n20731), .ZN(P1_U2805) );
  OAI21_X1 U22844 ( .B1(n19886), .B2(n19885), .A(n20030), .ZN(P1_U2806) );
  NOR4_X1 U22845 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19890) );
  NOR4_X1 U22846 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19889) );
  NOR4_X1 U22847 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19888) );
  NOR4_X1 U22848 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19887) );
  NAND4_X1 U22849 ( .A1(n19890), .A2(n19889), .A3(n19888), .A4(n19887), .ZN(
        n19896) );
  NOR4_X1 U22850 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19894) );
  AOI211_X1 U22851 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_15__SCAN_IN), .B(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19893) );
  NOR4_X1 U22852 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19892) );
  NOR4_X1 U22853 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19891) );
  NAND4_X1 U22854 ( .A1(n19894), .A2(n19893), .A3(n19892), .A4(n19891), .ZN(
        n19895) );
  NOR2_X1 U22855 ( .A1(n19896), .A2(n19895), .ZN(n20748) );
  INV_X1 U22856 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20726) );
  NOR3_X1 U22857 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19898) );
  OAI21_X1 U22858 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19898), .A(n20748), .ZN(
        n19897) );
  OAI21_X1 U22859 ( .B1(n20748), .B2(n20726), .A(n19897), .ZN(P1_U2807) );
  INV_X1 U22860 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20744) );
  INV_X1 U22861 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20732) );
  AOI21_X1 U22862 ( .B1(n20744), .B2(n20732), .A(n19898), .ZN(n19899) );
  INV_X1 U22863 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20723) );
  INV_X1 U22864 ( .A(n20748), .ZN(n20751) );
  AOI22_X1 U22865 ( .A1(n20748), .A2(n19899), .B1(n20723), .B2(n20751), .ZN(
        P1_U2808) );
  AOI21_X1 U22866 ( .B1(n19972), .B2(n19913), .A(n19959), .ZN(n19922) );
  AOI22_X1 U22867 ( .A1(n19967), .A2(P1_EBX_REG_9__SCAN_IN), .B1(n19961), .B2(
        n19900), .ZN(n19910) );
  INV_X1 U22868 ( .A(n19901), .ZN(n19908) );
  AOI22_X1 U22869 ( .A1(n19948), .A2(n19903), .B1(n19902), .B2(n13654), .ZN(
        n19904) );
  OAI211_X1 U22870 ( .C1(n19906), .C2(n19905), .A(n19904), .B(n20036), .ZN(
        n19907) );
  AOI21_X1 U22871 ( .B1(n19908), .B2(n19942), .A(n19907), .ZN(n19909) );
  OAI211_X1 U22872 ( .C1(n19922), .C2(n13654), .A(n19910), .B(n19909), .ZN(
        P1_U2831) );
  INV_X1 U22873 ( .A(n19911), .ZN(n19912) );
  AOI22_X1 U22874 ( .A1(n19967), .A2(P1_EBX_REG_8__SCAN_IN), .B1(n19912), .B2(
        n19961), .ZN(n19921) );
  AND2_X1 U22875 ( .A1(n19913), .A2(n19972), .ZN(n19914) );
  AOI22_X1 U22876 ( .A1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19962), .B1(
        n19915), .B2(n19914), .ZN(n19916) );
  OAI211_X1 U22877 ( .C1(n19917), .C2(n19976), .A(n19916), .B(n20036), .ZN(
        n19918) );
  AOI21_X1 U22878 ( .B1(n19919), .B2(n19942), .A(n19918), .ZN(n19920) );
  OAI211_X1 U22879 ( .C1(n19922), .C2(n20679), .A(n19921), .B(n19920), .ZN(
        P1_U2832) );
  AOI21_X1 U22880 ( .B1(n19972), .B2(n19923), .A(n19959), .ZN(n19945) );
  NOR3_X1 U22881 ( .A1(n19924), .A2(P1_REIP_REG_7__SCAN_IN), .A3(n19923), .ZN(
        n19925) );
  AOI21_X1 U22882 ( .B1(n19967), .B2(P1_EBX_REG_7__SCAN_IN), .A(n19925), .ZN(
        n19934) );
  NAND2_X1 U22883 ( .A1(n19962), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n19926) );
  OAI211_X1 U22884 ( .C1(n19950), .C2(n19927), .A(n20036), .B(n19926), .ZN(
        n19931) );
  NOR2_X1 U22885 ( .A1(n19929), .A2(n19928), .ZN(n19930) );
  AOI211_X1 U22886 ( .C1(n19932), .C2(n19948), .A(n19931), .B(n19930), .ZN(
        n19933) );
  OAI211_X1 U22887 ( .C1(n19945), .C2(n20678), .A(n19934), .B(n19933), .ZN(
        P1_U2833) );
  NAND2_X1 U22888 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n19935), .ZN(n19946) );
  INV_X1 U22889 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20676) );
  AOI21_X1 U22890 ( .B1(n19962), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n10704), .ZN(n19936) );
  OAI21_X1 U22891 ( .B1(n19950), .B2(n19937), .A(n19936), .ZN(n19938) );
  AOI21_X1 U22892 ( .B1(n19967), .B2(P1_EBX_REG_6__SCAN_IN), .A(n19938), .ZN(
        n19939) );
  OAI21_X1 U22893 ( .B1(n19940), .B2(n19976), .A(n19939), .ZN(n19941) );
  AOI21_X1 U22894 ( .B1(n19943), .B2(n19942), .A(n19941), .ZN(n19944) );
  OAI221_X1 U22895 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(n19946), .C1(n20676), 
        .C2(n19945), .A(n19944), .ZN(P1_U2834) );
  INV_X1 U22896 ( .A(n20037), .ZN(n19947) );
  AOI22_X1 U22897 ( .A1(n19967), .A2(P1_EBX_REG_4__SCAN_IN), .B1(n19948), .B2(
        n19947), .ZN(n19958) );
  OAI22_X1 U22898 ( .A1(n20022), .A2(n19950), .B1(n19949), .B2(n19965), .ZN(
        n19951) );
  AOI211_X1 U22899 ( .C1(n19962), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n10704), .B(n19951), .ZN(n19957) );
  NAND2_X1 U22900 ( .A1(n20672), .A2(n19952), .ZN(n19954) );
  AOI22_X1 U22901 ( .A1(n20018), .A2(n19955), .B1(n19954), .B2(n19953), .ZN(
        n19956) );
  NAND3_X1 U22902 ( .A1(n19958), .A2(n19957), .A3(n19956), .ZN(P1_U2836) );
  AOI22_X1 U22903 ( .A1(n19961), .A2(n19960), .B1(n19959), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n19964) );
  NAND2_X1 U22904 ( .A1(n19962), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n19963) );
  OAI211_X1 U22905 ( .C1(n12997), .C2(n19965), .A(n19964), .B(n19963), .ZN(
        n19966) );
  AOI21_X1 U22906 ( .B1(n19967), .B2(P1_EBX_REG_1__SCAN_IN), .A(n19966), .ZN(
        n19968) );
  OAI21_X1 U22907 ( .B1(n19970), .B2(n19969), .A(n19968), .ZN(n19971) );
  INV_X1 U22908 ( .A(n19971), .ZN(n19974) );
  NAND2_X1 U22909 ( .A1(n19972), .A2(n20744), .ZN(n19973) );
  OAI211_X1 U22910 ( .C1(n19976), .C2(n19975), .A(n19974), .B(n19973), .ZN(
        P1_U2839) );
  AOI22_X1 U22911 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n19979), .B1(n20008), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19977) );
  OAI21_X1 U22912 ( .B1(n20758), .B2(n19978), .A(n19977), .ZN(P1_U2921) );
  AOI22_X1 U22913 ( .A1(n20009), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20008), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19980) );
  OAI21_X1 U22914 ( .B1(n19981), .B2(n20011), .A(n19980), .ZN(P1_U2922) );
  AOI22_X1 U22915 ( .A1(n20009), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20008), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19982) );
  OAI21_X1 U22916 ( .B1(n19983), .B2(n20011), .A(n19982), .ZN(P1_U2923) );
  AOI22_X1 U22917 ( .A1(n20009), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20008), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19984) );
  OAI21_X1 U22918 ( .B1(n19985), .B2(n20011), .A(n19984), .ZN(P1_U2924) );
  AOI22_X1 U22919 ( .A1(n20009), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20008), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19986) );
  OAI21_X1 U22920 ( .B1(n19987), .B2(n20011), .A(n19986), .ZN(P1_U2925) );
  AOI22_X1 U22921 ( .A1(n20009), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n19999), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19988) );
  OAI21_X1 U22922 ( .B1(n19989), .B2(n20011), .A(n19988), .ZN(P1_U2926) );
  AOI22_X1 U22923 ( .A1(n20009), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n19999), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19990) );
  OAI21_X1 U22924 ( .B1(n19991), .B2(n20011), .A(n19990), .ZN(P1_U2927) );
  AOI22_X1 U22925 ( .A1(n20009), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n19999), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19992) );
  OAI21_X1 U22926 ( .B1(n19993), .B2(n20011), .A(n19992), .ZN(P1_U2928) );
  AOI22_X1 U22927 ( .A1(n20009), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n19999), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19994) );
  OAI21_X1 U22928 ( .B1(n19995), .B2(n20011), .A(n19994), .ZN(P1_U2929) );
  AOI22_X1 U22929 ( .A1(n20009), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20008), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19996) );
  OAI21_X1 U22930 ( .B1(n19997), .B2(n20011), .A(n19996), .ZN(P1_U2930) );
  AOI22_X1 U22931 ( .A1(n20009), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20008), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19998) );
  OAI21_X1 U22932 ( .B1(n11111), .B2(n20011), .A(n19998), .ZN(P1_U2931) );
  AOI22_X1 U22933 ( .A1(n20009), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n19999), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20000) );
  OAI21_X1 U22934 ( .B1(n20001), .B2(n20011), .A(n20000), .ZN(P1_U2932) );
  AOI22_X1 U22935 ( .A1(n20009), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20008), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20002) );
  OAI21_X1 U22936 ( .B1(n20003), .B2(n20011), .A(n20002), .ZN(P1_U2933) );
  AOI22_X1 U22937 ( .A1(n20009), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20008), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20004) );
  OAI21_X1 U22938 ( .B1(n20005), .B2(n20011), .A(n20004), .ZN(P1_U2934) );
  AOI22_X1 U22939 ( .A1(n20009), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20008), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20006) );
  OAI21_X1 U22940 ( .B1(n20007), .B2(n20011), .A(n20006), .ZN(P1_U2935) );
  AOI22_X1 U22941 ( .A1(n20009), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20008), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20010) );
  OAI21_X1 U22942 ( .B1(n20012), .B2(n20011), .A(n20010), .ZN(P1_U2936) );
  AOI22_X1 U22943 ( .A1(n20013), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n10704), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20021) );
  OAI21_X1 U22944 ( .B1(n20016), .B2(n20015), .A(n20014), .ZN(n20017) );
  INV_X1 U22945 ( .A(n20017), .ZN(n20042) );
  AOI22_X1 U22946 ( .A1(n20042), .A2(n20019), .B1(n14447), .B2(n20018), .ZN(
        n20020) );
  OAI211_X1 U22947 ( .C1(n20023), .C2(n20022), .A(n20021), .B(n20020), .ZN(
        P1_U2995) );
  NAND2_X1 U22948 ( .A1(n20025), .A2(n20024), .ZN(n20026) );
  AOI22_X1 U22949 ( .A1(n14447), .A2(n20027), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20026), .ZN(n20029) );
  NAND2_X1 U22950 ( .A1(n10704), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n20028) );
  OAI211_X1 U22951 ( .C1(n20031), .C2(n20030), .A(n20029), .B(n20028), .ZN(
        P1_U2999) );
  NOR2_X1 U22952 ( .A1(n20056), .A2(n20032), .ZN(n20057) );
  OAI21_X1 U22953 ( .B1(n20034), .B2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n20033), .ZN(n20062) );
  AOI211_X1 U22954 ( .C1(n20067), .C2(n20035), .A(n20057), .B(n20062), .ZN(
        n20053) );
  OAI22_X1 U22955 ( .A1(n20038), .A2(n20037), .B1(n20672), .B2(n20036), .ZN(
        n20041) );
  AOI211_X1 U22956 ( .C1(n20044), .C2(n20052), .A(n20039), .B(n20047), .ZN(
        n20040) );
  AOI211_X1 U22957 ( .C1(n20042), .C2(n20063), .A(n20041), .B(n20040), .ZN(
        n20043) );
  OAI21_X1 U22958 ( .B1(n20053), .B2(n20044), .A(n20043), .ZN(P1_U3027) );
  AOI21_X1 U22959 ( .B1(n20059), .B2(n20046), .A(n20045), .ZN(n20051) );
  INV_X1 U22960 ( .A(n20047), .ZN(n20048) );
  AOI22_X1 U22961 ( .A1(n20049), .A2(n20063), .B1(n20052), .B2(n20048), .ZN(
        n20050) );
  OAI211_X1 U22962 ( .C1(n20053), .C2(n20052), .A(n20051), .B(n20050), .ZN(
        P1_U3028) );
  NOR3_X1 U22963 ( .A1(n20056), .A2(n20055), .A3(n20054), .ZN(n20058) );
  AOI211_X1 U22964 ( .C1(n20060), .C2(n20059), .A(n20058), .B(n20057), .ZN(
        n20071) );
  INV_X1 U22965 ( .A(n20061), .ZN(n20064) );
  AOI22_X1 U22966 ( .A1(n20064), .A2(n20063), .B1(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20062), .ZN(n20070) );
  NAND2_X1 U22967 ( .A1(n10704), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n20069) );
  NAND3_X1 U22968 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20067), .A3(
        n20066), .ZN(n20068) );
  NAND4_X1 U22969 ( .A1(n20071), .A2(n20070), .A3(n20069), .A4(n20068), .ZN(
        P1_U3029) );
  NOR2_X1 U22970 ( .A1(n20072), .A2(n20740), .ZN(P1_U3032) );
  AND2_X1 U22971 ( .A1(n20074), .A2(n20104), .ZN(n20587) );
  OAI22_X1 U22972 ( .A1(n20629), .A2(n20598), .B1(n20106), .B2(n20396), .ZN(
        n20075) );
  INV_X1 U22973 ( .A(n20075), .ZN(n20078) );
  NOR2_X2 U22974 ( .A1(n20076), .A2(n20224), .ZN(n20588) );
  AOI22_X1 U22975 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20109), .B1(DATAI_16_), 
        .B2(n13388), .ZN(n20554) );
  INV_X1 U22976 ( .A(n20554), .ZN(n20595) );
  AOI22_X1 U22977 ( .A1(n20588), .A2(n20110), .B1(n20127), .B2(n20595), .ZN(
        n20077) );
  OAI211_X1 U22978 ( .C1(n20114), .C2(n20079), .A(n20078), .B(n20077), .ZN(
        P1_U3033) );
  AOI22_X1 U22979 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20109), .B1(DATAI_25_), 
        .B2(n13388), .ZN(n20491) );
  INV_X1 U22980 ( .A(n20599), .ZN(n20410) );
  OAI22_X1 U22981 ( .A1(n20629), .A2(n20491), .B1(n20106), .B2(n20410), .ZN(
        n20081) );
  INV_X1 U22982 ( .A(n20081), .ZN(n20084) );
  NOR2_X2 U22983 ( .A1(n20082), .A2(n20224), .ZN(n20600) );
  INV_X1 U22984 ( .A(n20604), .ZN(n20488) );
  AOI22_X1 U22985 ( .A1(n20600), .A2(n20110), .B1(n20127), .B2(n20488), .ZN(
        n20083) );
  OAI211_X1 U22986 ( .C1(n20114), .C2(n20085), .A(n20084), .B(n20083), .ZN(
        P1_U3034) );
  AOI22_X1 U22987 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20109), .B1(DATAI_27_), 
        .B2(n13388), .ZN(n20616) );
  INV_X1 U22988 ( .A(n20611), .ZN(n20418) );
  OAI22_X1 U22989 ( .A1(n20629), .A2(n20616), .B1(n20106), .B2(n20418), .ZN(
        n20087) );
  INV_X1 U22990 ( .A(n20087), .ZN(n20090) );
  NOR2_X2 U22991 ( .A1(n20088), .A2(n20224), .ZN(n20612) );
  AOI22_X1 U22992 ( .A1(DATAI_19_), .A2(n13388), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n20109), .ZN(n20564) );
  INV_X1 U22993 ( .A(n20564), .ZN(n20613) );
  AOI22_X1 U22994 ( .A1(n20612), .A2(n20110), .B1(n20127), .B2(n20613), .ZN(
        n20089) );
  OAI211_X1 U22995 ( .C1(n20114), .C2(n20091), .A(n20090), .B(n20089), .ZN(
        P1_U3036) );
  AOI22_X1 U22996 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20109), .B1(DATAI_29_), 
        .B2(n13388), .ZN(n20501) );
  AND2_X1 U22997 ( .A1(n20092), .A2(n20104), .ZN(n20623) );
  INV_X1 U22998 ( .A(n20623), .ZN(n20426) );
  OAI22_X1 U22999 ( .A1(n20629), .A2(n20501), .B1(n20106), .B2(n20426), .ZN(
        n20093) );
  INV_X1 U23000 ( .A(n20093), .ZN(n20096) );
  NOR2_X2 U23001 ( .A1(n20094), .A2(n20224), .ZN(n20624) );
  AOI22_X1 U23002 ( .A1(DATAI_21_), .A2(n13388), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20109), .ZN(n20630) );
  INV_X1 U23003 ( .A(n20630), .ZN(n20498) );
  AOI22_X1 U23004 ( .A1(n20624), .A2(n20110), .B1(n20127), .B2(n20498), .ZN(
        n20095) );
  OAI211_X1 U23005 ( .C1(n20114), .C2(n20097), .A(n20096), .B(n20095), .ZN(
        P1_U3038) );
  INV_X1 U23006 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n20103) );
  OAI22_X1 U23007 ( .A1(n20629), .A2(n20636), .B1(n20106), .B2(n20430), .ZN(
        n20099) );
  INV_X1 U23008 ( .A(n20099), .ZN(n20102) );
  NOR2_X2 U23009 ( .A1(n20100), .A2(n20224), .ZN(n20632) );
  AOI22_X1 U23010 ( .A1(DATAI_22_), .A2(n13388), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n20109), .ZN(n20533) );
  INV_X1 U23011 ( .A(n20533), .ZN(n20633) );
  AOI22_X1 U23012 ( .A1(n20632), .A2(n20110), .B1(n20127), .B2(n20633), .ZN(
        n20101) );
  OAI211_X1 U23013 ( .C1(n20114), .C2(n20103), .A(n20102), .B(n20101), .ZN(
        P1_U3039) );
  OAI22_X1 U23014 ( .A1(n20629), .A2(n20647), .B1(n20106), .B2(n20435), .ZN(
        n20107) );
  INV_X1 U23015 ( .A(n20107), .ZN(n20112) );
  NOR2_X2 U23016 ( .A1(n20108), .A2(n20224), .ZN(n20640) );
  AOI22_X1 U23017 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20109), .B1(DATAI_23_), 
        .B2(n13388), .ZN(n20581) );
  INV_X1 U23018 ( .A(n20581), .ZN(n20641) );
  AOI22_X1 U23019 ( .A1(n20640), .A2(n20110), .B1(n20127), .B2(n20641), .ZN(
        n20111) );
  OAI211_X1 U23020 ( .C1(n20114), .C2(n20113), .A(n20112), .B(n20111), .ZN(
        P1_U3040) );
  INV_X1 U23021 ( .A(n20739), .ZN(n20510) );
  INV_X1 U23022 ( .A(n20115), .ZN(n20512) );
  NOR2_X1 U23023 ( .A1(n20742), .A2(n20116), .ZN(n20136) );
  AOI21_X1 U23024 ( .B1(n20184), .B2(n20512), .A(n20136), .ZN(n20118) );
  OAI22_X1 U23025 ( .A1(n20118), .A2(n20586), .B1(n20116), .B2(n20652), .ZN(
        n20137) );
  AOI22_X1 U23026 ( .A1(n20588), .A2(n20137), .B1(n20587), .B2(n20136), .ZN(
        n20122) );
  INV_X1 U23027 ( .A(n20116), .ZN(n20120) );
  OAI21_X1 U23028 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n20481), .A(
        n20117), .ZN(n20185) );
  OAI211_X1 U23029 ( .C1(n20180), .C2(n20515), .A(n20369), .B(n20118), .ZN(
        n20119) );
  OAI211_X1 U23030 ( .C1(n20369), .C2(n20120), .A(n20593), .B(n20119), .ZN(
        n20138) );
  INV_X1 U23031 ( .A(n20598), .ZN(n20551) );
  AOI22_X1 U23032 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20138), .B1(
        n20127), .B2(n20551), .ZN(n20121) );
  OAI211_X1 U23033 ( .C1(n20554), .C2(n20177), .A(n20122), .B(n20121), .ZN(
        P1_U3041) );
  AOI22_X1 U23034 ( .A1(n20600), .A2(n20137), .B1(n20599), .B2(n20136), .ZN(
        n20124) );
  INV_X1 U23035 ( .A(n20491), .ZN(n20601) );
  AOI22_X1 U23036 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20138), .B1(
        n20127), .B2(n20601), .ZN(n20123) );
  OAI211_X1 U23037 ( .C1(n20604), .C2(n20177), .A(n20124), .B(n20123), .ZN(
        P1_U3042) );
  AOI22_X1 U23038 ( .A1(n20606), .A2(n20137), .B1(n20605), .B2(n20136), .ZN(
        n20126) );
  INV_X1 U23039 ( .A(n20560), .ZN(n20607) );
  AOI22_X1 U23040 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20138), .B1(
        n20143), .B2(n20607), .ZN(n20125) );
  OAI211_X1 U23041 ( .C1(n20610), .C2(n20141), .A(n20126), .B(n20125), .ZN(
        P1_U3043) );
  AOI22_X1 U23042 ( .A1(n20612), .A2(n20137), .B1(n20611), .B2(n20136), .ZN(
        n20129) );
  INV_X1 U23043 ( .A(n20616), .ZN(n20561) );
  AOI22_X1 U23044 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20138), .B1(
        n20127), .B2(n20561), .ZN(n20128) );
  OAI211_X1 U23045 ( .C1(n20564), .C2(n20177), .A(n20129), .B(n20128), .ZN(
        P1_U3044) );
  AOI22_X1 U23046 ( .A1(n20137), .A2(n20618), .B1(n20617), .B2(n20136), .ZN(
        n20131) );
  INV_X1 U23047 ( .A(n20568), .ZN(n20619) );
  AOI22_X1 U23048 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20138), .B1(
        n20143), .B2(n20619), .ZN(n20130) );
  OAI211_X1 U23049 ( .C1(n20622), .C2(n20141), .A(n20131), .B(n20130), .ZN(
        P1_U3045) );
  AOI22_X1 U23050 ( .A1(n20624), .A2(n20137), .B1(n20623), .B2(n20136), .ZN(
        n20133) );
  AOI22_X1 U23051 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20138), .B1(
        n20143), .B2(n20498), .ZN(n20132) );
  OAI211_X1 U23052 ( .C1(n20501), .C2(n20141), .A(n20133), .B(n20132), .ZN(
        P1_U3046) );
  AOI22_X1 U23053 ( .A1(n20632), .A2(n20137), .B1(n20631), .B2(n20136), .ZN(
        n20135) );
  AOI22_X1 U23054 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20138), .B1(
        n20143), .B2(n20633), .ZN(n20134) );
  OAI211_X1 U23055 ( .C1(n20636), .C2(n20141), .A(n20135), .B(n20134), .ZN(
        P1_U3047) );
  AOI22_X1 U23056 ( .A1(n20640), .A2(n20137), .B1(n20637), .B2(n20136), .ZN(
        n20140) );
  AOI22_X1 U23057 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20138), .B1(
        n20143), .B2(n20641), .ZN(n20139) );
  OAI211_X1 U23058 ( .C1(n20647), .C2(n20141), .A(n20140), .B(n20139), .ZN(
        P1_U3048) );
  NAND3_X1 U23059 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20442), .A3(
        n20395), .ZN(n20188) );
  OR2_X1 U23060 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20188), .ZN(
        n20171) );
  OAI22_X1 U23061 ( .A1(n20212), .A2(n20554), .B1(n20396), .B2(n20171), .ZN(
        n20142) );
  INV_X1 U23062 ( .A(n20142), .ZN(n20152) );
  INV_X1 U23063 ( .A(n20212), .ZN(n20144) );
  OAI21_X1 U23064 ( .B1(n20144), .B2(n20143), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20145) );
  NAND2_X1 U23065 ( .A1(n20145), .A2(n20369), .ZN(n20150) );
  NOR2_X1 U23066 ( .A1(n20146), .A2(n12997), .ZN(n20148) );
  OR2_X1 U23067 ( .A1(n20399), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20280) );
  AND2_X1 U23068 ( .A1(n20280), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20276) );
  AOI211_X1 U23069 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20171), .A(n20276), 
        .B(n20342), .ZN(n20147) );
  INV_X1 U23070 ( .A(n20148), .ZN(n20149) );
  OAI22_X1 U23071 ( .A1(n20150), .A2(n20149), .B1(n20405), .B2(n20280), .ZN(
        n20173) );
  AOI22_X1 U23072 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20174), .B1(
        n20588), .B2(n20173), .ZN(n20151) );
  OAI211_X1 U23073 ( .C1(n20598), .C2(n20177), .A(n20152), .B(n20151), .ZN(
        P1_U3049) );
  OAI22_X1 U23074 ( .A1(n20177), .A2(n20491), .B1(n20410), .B2(n20171), .ZN(
        n20153) );
  INV_X1 U23075 ( .A(n20153), .ZN(n20155) );
  AOI22_X1 U23076 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20174), .B1(
        n20600), .B2(n20173), .ZN(n20154) );
  OAI211_X1 U23077 ( .C1(n20604), .C2(n20212), .A(n20155), .B(n20154), .ZN(
        P1_U3050) );
  INV_X1 U23078 ( .A(n20605), .ZN(n20414) );
  OAI22_X1 U23079 ( .A1(n20212), .A2(n20560), .B1(n20171), .B2(n20414), .ZN(
        n20156) );
  INV_X1 U23080 ( .A(n20156), .ZN(n20158) );
  AOI22_X1 U23081 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20174), .B1(
        n20606), .B2(n20173), .ZN(n20157) );
  OAI211_X1 U23082 ( .C1(n20610), .C2(n20177), .A(n20158), .B(n20157), .ZN(
        P1_U3051) );
  OAI22_X1 U23083 ( .A1(n20177), .A2(n20616), .B1(n20171), .B2(n20418), .ZN(
        n20159) );
  INV_X1 U23084 ( .A(n20159), .ZN(n20161) );
  AOI22_X1 U23085 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20174), .B1(
        n20612), .B2(n20173), .ZN(n20160) );
  OAI211_X1 U23086 ( .C1(n20564), .C2(n20212), .A(n20161), .B(n20160), .ZN(
        P1_U3052) );
  INV_X1 U23087 ( .A(n20617), .ZN(n20422) );
  OAI22_X1 U23088 ( .A1(n20212), .A2(n20568), .B1(n20171), .B2(n20422), .ZN(
        n20162) );
  INV_X1 U23089 ( .A(n20162), .ZN(n20164) );
  AOI22_X1 U23090 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20174), .B1(
        n20618), .B2(n20173), .ZN(n20163) );
  OAI211_X1 U23091 ( .C1(n20622), .C2(n20177), .A(n20164), .B(n20163), .ZN(
        P1_U3053) );
  OAI22_X1 U23092 ( .A1(n20212), .A2(n20630), .B1(n20426), .B2(n20171), .ZN(
        n20165) );
  INV_X1 U23093 ( .A(n20165), .ZN(n20167) );
  AOI22_X1 U23094 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20174), .B1(
        n20624), .B2(n20173), .ZN(n20166) );
  OAI211_X1 U23095 ( .C1(n20501), .C2(n20177), .A(n20167), .B(n20166), .ZN(
        P1_U3054) );
  OAI22_X1 U23096 ( .A1(n20212), .A2(n20533), .B1(n20171), .B2(n20430), .ZN(
        n20168) );
  INV_X1 U23097 ( .A(n20168), .ZN(n20170) );
  AOI22_X1 U23098 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20174), .B1(
        n20632), .B2(n20173), .ZN(n20169) );
  OAI211_X1 U23099 ( .C1(n20636), .C2(n20177), .A(n20170), .B(n20169), .ZN(
        P1_U3055) );
  OAI22_X1 U23100 ( .A1(n20212), .A2(n20581), .B1(n20171), .B2(n20435), .ZN(
        n20172) );
  INV_X1 U23101 ( .A(n20172), .ZN(n20176) );
  AOI22_X1 U23102 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20174), .B1(
        n20640), .B2(n20173), .ZN(n20175) );
  OAI211_X1 U23103 ( .C1(n20647), .C2(n20177), .A(n20176), .B(n20175), .ZN(
        P1_U3056) );
  INV_X1 U23104 ( .A(n20312), .ZN(n20449) );
  INV_X1 U23105 ( .A(n20443), .ZN(n20178) );
  NAND2_X1 U23106 ( .A1(n20178), .A2(n20442), .ZN(n20211) );
  OAI22_X1 U23107 ( .A1(n20246), .A2(n20554), .B1(n20396), .B2(n20211), .ZN(
        n20179) );
  INV_X1 U23108 ( .A(n20179), .ZN(n20192) );
  OAI21_X1 U23109 ( .B1(n20180), .B2(n20590), .A(n20369), .ZN(n20189) );
  AND2_X1 U23110 ( .A1(n20182), .A2(n20181), .ZN(n20583) );
  INV_X1 U23111 ( .A(n20211), .ZN(n20183) );
  AOI21_X1 U23112 ( .B1(n20184), .B2(n20583), .A(n20183), .ZN(n20190) );
  INV_X1 U23113 ( .A(n20190), .ZN(n20187) );
  AOI21_X1 U23114 ( .B1(n20586), .B2(n20188), .A(n20185), .ZN(n20186) );
  OAI21_X1 U23115 ( .B1(n20189), .B2(n20187), .A(n20186), .ZN(n20215) );
  OAI22_X1 U23116 ( .A1(n20190), .A2(n20189), .B1(n20652), .B2(n20188), .ZN(
        n20214) );
  AOI22_X1 U23117 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20215), .B1(
        n20588), .B2(n20214), .ZN(n20191) );
  OAI211_X1 U23118 ( .C1(n20598), .C2(n20212), .A(n20192), .B(n20191), .ZN(
        P1_U3057) );
  OAI22_X1 U23119 ( .A1(n20246), .A2(n20604), .B1(n20211), .B2(n20410), .ZN(
        n20193) );
  INV_X1 U23120 ( .A(n20193), .ZN(n20195) );
  AOI22_X1 U23121 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20215), .B1(
        n20600), .B2(n20214), .ZN(n20194) );
  OAI211_X1 U23122 ( .C1(n20491), .C2(n20212), .A(n20195), .B(n20194), .ZN(
        P1_U3058) );
  OAI22_X1 U23123 ( .A1(n20246), .A2(n20560), .B1(n20211), .B2(n20414), .ZN(
        n20196) );
  INV_X1 U23124 ( .A(n20196), .ZN(n20198) );
  AOI22_X1 U23125 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20215), .B1(
        n20606), .B2(n20214), .ZN(n20197) );
  OAI211_X1 U23126 ( .C1(n20610), .C2(n20212), .A(n20198), .B(n20197), .ZN(
        P1_U3059) );
  OAI22_X1 U23127 ( .A1(n20212), .A2(n20616), .B1(n20211), .B2(n20418), .ZN(
        n20199) );
  INV_X1 U23128 ( .A(n20199), .ZN(n20201) );
  AOI22_X1 U23129 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20215), .B1(
        n20612), .B2(n20214), .ZN(n20200) );
  OAI211_X1 U23130 ( .C1(n20564), .C2(n20246), .A(n20201), .B(n20200), .ZN(
        P1_U3060) );
  OAI22_X1 U23131 ( .A1(n20246), .A2(n20568), .B1(n20211), .B2(n20422), .ZN(
        n20202) );
  INV_X1 U23132 ( .A(n20202), .ZN(n20204) );
  AOI22_X1 U23133 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20215), .B1(
        n20618), .B2(n20214), .ZN(n20203) );
  OAI211_X1 U23134 ( .C1(n20622), .C2(n20212), .A(n20204), .B(n20203), .ZN(
        P1_U3061) );
  OAI22_X1 U23135 ( .A1(n20246), .A2(n20630), .B1(n20211), .B2(n20426), .ZN(
        n20205) );
  INV_X1 U23136 ( .A(n20205), .ZN(n20207) );
  AOI22_X1 U23137 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20215), .B1(
        n20624), .B2(n20214), .ZN(n20206) );
  OAI211_X1 U23138 ( .C1(n20501), .C2(n20212), .A(n20207), .B(n20206), .ZN(
        P1_U3062) );
  OAI22_X1 U23139 ( .A1(n20212), .A2(n20636), .B1(n20211), .B2(n20430), .ZN(
        n20208) );
  INV_X1 U23140 ( .A(n20208), .ZN(n20210) );
  AOI22_X1 U23141 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20215), .B1(
        n20632), .B2(n20214), .ZN(n20209) );
  OAI211_X1 U23142 ( .C1(n20533), .C2(n20246), .A(n20210), .B(n20209), .ZN(
        P1_U3063) );
  OAI22_X1 U23143 ( .A1(n20212), .A2(n20647), .B1(n20211), .B2(n20435), .ZN(
        n20213) );
  INV_X1 U23144 ( .A(n20213), .ZN(n20217) );
  AOI22_X1 U23145 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20215), .B1(
        n20640), .B2(n20214), .ZN(n20216) );
  OAI211_X1 U23146 ( .C1(n20581), .C2(n20246), .A(n20217), .B(n20216), .ZN(
        P1_U3064) );
  NOR2_X1 U23147 ( .A1(n12944), .A2(n20218), .ZN(n20315) );
  NAND3_X1 U23148 ( .A1(n20315), .A2(n20738), .A3(n12997), .ZN(n20219) );
  OAI21_X1 U23149 ( .B1(n20544), .B2(n20220), .A(n20219), .ZN(n20242) );
  NAND3_X1 U23150 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20442), .A3(
        n20475), .ZN(n20247) );
  NOR2_X1 U23151 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20247), .ZN(
        n20241) );
  AOI22_X1 U23152 ( .A1(n20588), .A2(n20242), .B1(n20587), .B2(n20241), .ZN(
        n20227) );
  AOI21_X1 U23153 ( .B1(n20246), .B2(n20271), .A(n20515), .ZN(n20221) );
  AOI21_X1 U23154 ( .B1(n20315), .B2(n12997), .A(n20221), .ZN(n20222) );
  NOR2_X1 U23155 ( .A1(n20222), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20225) );
  AOI22_X1 U23156 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20243), .B1(
        n20261), .B2(n20595), .ZN(n20226) );
  OAI211_X1 U23157 ( .C1(n20598), .C2(n20246), .A(n20227), .B(n20226), .ZN(
        P1_U3065) );
  AOI22_X1 U23158 ( .A1(n20600), .A2(n20242), .B1(n20599), .B2(n20241), .ZN(
        n20229) );
  INV_X1 U23159 ( .A(n20246), .ZN(n20232) );
  AOI22_X1 U23160 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20243), .B1(
        n20232), .B2(n20601), .ZN(n20228) );
  OAI211_X1 U23161 ( .C1(n20604), .C2(n20271), .A(n20229), .B(n20228), .ZN(
        P1_U3066) );
  AOI22_X1 U23162 ( .A1(n20606), .A2(n20242), .B1(n20605), .B2(n20241), .ZN(
        n20231) );
  AOI22_X1 U23163 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20243), .B1(
        n20261), .B2(n20607), .ZN(n20230) );
  OAI211_X1 U23164 ( .C1(n20610), .C2(n20246), .A(n20231), .B(n20230), .ZN(
        P1_U3067) );
  AOI22_X1 U23165 ( .A1(n20612), .A2(n20242), .B1(n20611), .B2(n20241), .ZN(
        n20234) );
  AOI22_X1 U23166 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20243), .B1(
        n20232), .B2(n20561), .ZN(n20233) );
  OAI211_X1 U23167 ( .C1(n20564), .C2(n20271), .A(n20234), .B(n20233), .ZN(
        P1_U3068) );
  AOI22_X1 U23168 ( .A1(n20242), .A2(n20618), .B1(n20617), .B2(n20241), .ZN(
        n20236) );
  AOI22_X1 U23169 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20243), .B1(
        n20261), .B2(n20619), .ZN(n20235) );
  OAI211_X1 U23170 ( .C1(n20622), .C2(n20246), .A(n20236), .B(n20235), .ZN(
        P1_U3069) );
  AOI22_X1 U23171 ( .A1(n20624), .A2(n20242), .B1(n20623), .B2(n20241), .ZN(
        n20238) );
  AOI22_X1 U23172 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20243), .B1(
        n20261), .B2(n20498), .ZN(n20237) );
  OAI211_X1 U23173 ( .C1(n20501), .C2(n20246), .A(n20238), .B(n20237), .ZN(
        P1_U3070) );
  AOI22_X1 U23174 ( .A1(n20632), .A2(n20242), .B1(n20631), .B2(n20241), .ZN(
        n20240) );
  AOI22_X1 U23175 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20243), .B1(
        n20261), .B2(n20633), .ZN(n20239) );
  OAI211_X1 U23176 ( .C1(n20636), .C2(n20246), .A(n20240), .B(n20239), .ZN(
        P1_U3071) );
  AOI22_X1 U23177 ( .A1(n20640), .A2(n20242), .B1(n20637), .B2(n20241), .ZN(
        n20245) );
  AOI22_X1 U23178 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20243), .B1(
        n20261), .B2(n20641), .ZN(n20244) );
  OAI211_X1 U23179 ( .C1(n20647), .C2(n20246), .A(n20245), .B(n20244), .ZN(
        P1_U3072) );
  NOR2_X1 U23180 ( .A1(n20742), .A2(n20247), .ZN(n20266) );
  AOI21_X1 U23181 ( .B1(n20315), .B2(n20512), .A(n20266), .ZN(n20248) );
  OAI22_X1 U23182 ( .A1(n20248), .A2(n20586), .B1(n20247), .B2(n20652), .ZN(
        n20267) );
  AOI22_X1 U23183 ( .A1(n20588), .A2(n20267), .B1(n20587), .B2(n20266), .ZN(
        n20252) );
  INV_X1 U23184 ( .A(n20247), .ZN(n20250) );
  OAI21_X1 U23185 ( .B1(n20311), .B2(n20515), .A(n20248), .ZN(n20249) );
  OAI221_X1 U23186 ( .B1(n20738), .B2(n20250), .C1(n20586), .C2(n20249), .A(
        n20593), .ZN(n20268) );
  AOI22_X1 U23187 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20268), .B1(
        n20261), .B2(n20551), .ZN(n20251) );
  OAI211_X1 U23188 ( .C1(n20554), .C2(n20304), .A(n20252), .B(n20251), .ZN(
        P1_U3073) );
  AOI22_X1 U23189 ( .A1(n20600), .A2(n20267), .B1(n20599), .B2(n20266), .ZN(
        n20254) );
  AOI22_X1 U23190 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20268), .B1(
        n20273), .B2(n20488), .ZN(n20253) );
  OAI211_X1 U23191 ( .C1(n20491), .C2(n20271), .A(n20254), .B(n20253), .ZN(
        P1_U3074) );
  AOI22_X1 U23192 ( .A1(n20606), .A2(n20267), .B1(n20605), .B2(n20266), .ZN(
        n20256) );
  AOI22_X1 U23193 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20268), .B1(
        n20273), .B2(n20607), .ZN(n20255) );
  OAI211_X1 U23194 ( .C1(n20610), .C2(n20271), .A(n20256), .B(n20255), .ZN(
        P1_U3075) );
  AOI22_X1 U23195 ( .A1(n20612), .A2(n20267), .B1(n20611), .B2(n20266), .ZN(
        n20258) );
  AOI22_X1 U23196 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20268), .B1(
        n20273), .B2(n20613), .ZN(n20257) );
  OAI211_X1 U23197 ( .C1(n20616), .C2(n20271), .A(n20258), .B(n20257), .ZN(
        P1_U3076) );
  AOI22_X1 U23198 ( .A1(n20267), .A2(n20618), .B1(n20617), .B2(n20266), .ZN(
        n20260) );
  AOI22_X1 U23199 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20268), .B1(
        n20261), .B2(n20565), .ZN(n20259) );
  OAI211_X1 U23200 ( .C1(n20568), .C2(n20304), .A(n20260), .B(n20259), .ZN(
        P1_U3077) );
  AOI22_X1 U23201 ( .A1(n20624), .A2(n20267), .B1(n20623), .B2(n20266), .ZN(
        n20263) );
  INV_X1 U23202 ( .A(n20501), .ZN(n20625) );
  AOI22_X1 U23203 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20268), .B1(
        n20261), .B2(n20625), .ZN(n20262) );
  OAI211_X1 U23204 ( .C1(n20630), .C2(n20304), .A(n20263), .B(n20262), .ZN(
        P1_U3078) );
  AOI22_X1 U23205 ( .A1(n20632), .A2(n20267), .B1(n20631), .B2(n20266), .ZN(
        n20265) );
  AOI22_X1 U23206 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20268), .B1(
        n20273), .B2(n20633), .ZN(n20264) );
  OAI211_X1 U23207 ( .C1(n20636), .C2(n20271), .A(n20265), .B(n20264), .ZN(
        P1_U3079) );
  AOI22_X1 U23208 ( .A1(n20640), .A2(n20267), .B1(n20637), .B2(n20266), .ZN(
        n20270) );
  AOI22_X1 U23209 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20268), .B1(
        n20273), .B2(n20641), .ZN(n20269) );
  OAI211_X1 U23210 ( .C1(n20647), .C2(n20271), .A(n20270), .B(n20269), .ZN(
        P1_U3080) );
  INV_X1 U23211 ( .A(n20319), .ZN(n20316) );
  NOR2_X1 U23212 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20316), .ZN(
        n20279) );
  INV_X1 U23213 ( .A(n20279), .ZN(n20303) );
  OAI22_X1 U23214 ( .A1(n20304), .A2(n20598), .B1(n20396), .B2(n20303), .ZN(
        n20272) );
  INV_X1 U23215 ( .A(n20272), .ZN(n20284) );
  NOR3_X1 U23216 ( .A1(n20336), .A2(n20273), .A3(n20586), .ZN(n20275) );
  INV_X1 U23217 ( .A(n20477), .ZN(n20274) );
  NOR2_X1 U23218 ( .A1(n20275), .A2(n20274), .ZN(n20282) );
  INV_X1 U23219 ( .A(n20282), .ZN(n20277) );
  NAND2_X1 U23220 ( .A1(n20315), .A2(n20543), .ZN(n20281) );
  AOI21_X1 U23221 ( .B1(n20277), .B2(n20281), .A(n20276), .ZN(n20278) );
  OAI211_X1 U23222 ( .C1(n20279), .C2(n20481), .A(n20549), .B(n20278), .ZN(
        n20307) );
  OAI22_X1 U23223 ( .A1(n20282), .A2(n20281), .B1(n20280), .B2(n20544), .ZN(
        n20306) );
  AOI22_X1 U23224 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20307), .B1(
        n20588), .B2(n20306), .ZN(n20283) );
  OAI211_X1 U23225 ( .C1(n20554), .C2(n20310), .A(n20284), .B(n20283), .ZN(
        P1_U3081) );
  OAI22_X1 U23226 ( .A1(n20304), .A2(n20491), .B1(n20410), .B2(n20303), .ZN(
        n20285) );
  INV_X1 U23227 ( .A(n20285), .ZN(n20287) );
  AOI22_X1 U23228 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20307), .B1(
        n20600), .B2(n20306), .ZN(n20286) );
  OAI211_X1 U23229 ( .C1(n20604), .C2(n20310), .A(n20287), .B(n20286), .ZN(
        P1_U3082) );
  OAI22_X1 U23230 ( .A1(n20310), .A2(n20560), .B1(n20303), .B2(n20414), .ZN(
        n20288) );
  INV_X1 U23231 ( .A(n20288), .ZN(n20290) );
  AOI22_X1 U23232 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20307), .B1(
        n20606), .B2(n20306), .ZN(n20289) );
  OAI211_X1 U23233 ( .C1(n20610), .C2(n20304), .A(n20290), .B(n20289), .ZN(
        P1_U3083) );
  OAI22_X1 U23234 ( .A1(n20304), .A2(n20616), .B1(n20418), .B2(n20303), .ZN(
        n20291) );
  INV_X1 U23235 ( .A(n20291), .ZN(n20293) );
  AOI22_X1 U23236 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20307), .B1(
        n20612), .B2(n20306), .ZN(n20292) );
  OAI211_X1 U23237 ( .C1(n20564), .C2(n20310), .A(n20293), .B(n20292), .ZN(
        P1_U3084) );
  OAI22_X1 U23238 ( .A1(n20304), .A2(n20622), .B1(n20303), .B2(n20422), .ZN(
        n20294) );
  INV_X1 U23239 ( .A(n20294), .ZN(n20296) );
  AOI22_X1 U23240 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20307), .B1(
        n20618), .B2(n20306), .ZN(n20295) );
  OAI211_X1 U23241 ( .C1(n20568), .C2(n20310), .A(n20296), .B(n20295), .ZN(
        P1_U3085) );
  OAI22_X1 U23242 ( .A1(n20304), .A2(n20501), .B1(n20426), .B2(n20303), .ZN(
        n20297) );
  INV_X1 U23243 ( .A(n20297), .ZN(n20299) );
  AOI22_X1 U23244 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20307), .B1(
        n20624), .B2(n20306), .ZN(n20298) );
  OAI211_X1 U23245 ( .C1(n20630), .C2(n20310), .A(n20299), .B(n20298), .ZN(
        P1_U3086) );
  OAI22_X1 U23246 ( .A1(n20310), .A2(n20533), .B1(n20303), .B2(n20430), .ZN(
        n20300) );
  INV_X1 U23247 ( .A(n20300), .ZN(n20302) );
  AOI22_X1 U23248 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20307), .B1(
        n20632), .B2(n20306), .ZN(n20301) );
  OAI211_X1 U23249 ( .C1(n20636), .C2(n20304), .A(n20302), .B(n20301), .ZN(
        P1_U3087) );
  OAI22_X1 U23250 ( .A1(n20304), .A2(n20647), .B1(n20435), .B2(n20303), .ZN(
        n20305) );
  INV_X1 U23251 ( .A(n20305), .ZN(n20309) );
  AOI22_X1 U23252 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20307), .B1(
        n20640), .B2(n20306), .ZN(n20308) );
  OAI211_X1 U23253 ( .C1(n20581), .C2(n20310), .A(n20309), .B(n20308), .ZN(
        P1_U3088) );
  INV_X1 U23254 ( .A(n20311), .ZN(n20313) );
  INV_X1 U23255 ( .A(n20314), .ZN(n20334) );
  AOI21_X1 U23256 ( .B1(n20315), .B2(n20583), .A(n20334), .ZN(n20317) );
  OAI22_X1 U23257 ( .A1(n20317), .A2(n20586), .B1(n20316), .B2(n20652), .ZN(
        n20335) );
  AOI22_X1 U23258 ( .A1(n20588), .A2(n20335), .B1(n20334), .B2(n20587), .ZN(
        n20321) );
  OAI21_X1 U23259 ( .B1(n20319), .B2(n20318), .A(n20593), .ZN(n20337) );
  AOI22_X1 U23260 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20337), .B1(
        n20336), .B2(n20551), .ZN(n20320) );
  OAI211_X1 U23261 ( .C1(n20554), .C2(n20366), .A(n20321), .B(n20320), .ZN(
        P1_U3089) );
  AOI22_X1 U23262 ( .A1(n20600), .A2(n20335), .B1(n20334), .B2(n20599), .ZN(
        n20323) );
  AOI22_X1 U23263 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20337), .B1(
        n20336), .B2(n20601), .ZN(n20322) );
  OAI211_X1 U23264 ( .C1(n20604), .C2(n20366), .A(n20323), .B(n20322), .ZN(
        P1_U3090) );
  AOI22_X1 U23265 ( .A1(n20606), .A2(n20335), .B1(n20334), .B2(n20605), .ZN(
        n20325) );
  AOI22_X1 U23266 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20337), .B1(
        n20336), .B2(n20557), .ZN(n20324) );
  OAI211_X1 U23267 ( .C1(n20560), .C2(n20366), .A(n20325), .B(n20324), .ZN(
        P1_U3091) );
  AOI22_X1 U23268 ( .A1(n20612), .A2(n20335), .B1(n20334), .B2(n20611), .ZN(
        n20327) );
  AOI22_X1 U23269 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20337), .B1(
        n20336), .B2(n20561), .ZN(n20326) );
  OAI211_X1 U23270 ( .C1(n20564), .C2(n20366), .A(n20327), .B(n20326), .ZN(
        P1_U3092) );
  AOI22_X1 U23271 ( .A1(n20335), .A2(n20618), .B1(n20334), .B2(n20617), .ZN(
        n20329) );
  AOI22_X1 U23272 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20337), .B1(
        n20336), .B2(n20565), .ZN(n20328) );
  OAI211_X1 U23273 ( .C1(n20568), .C2(n20366), .A(n20329), .B(n20328), .ZN(
        P1_U3093) );
  AOI22_X1 U23274 ( .A1(n20624), .A2(n20335), .B1(n20334), .B2(n20623), .ZN(
        n20331) );
  AOI22_X1 U23275 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20337), .B1(
        n20336), .B2(n20625), .ZN(n20330) );
  OAI211_X1 U23276 ( .C1(n20630), .C2(n20366), .A(n20331), .B(n20330), .ZN(
        P1_U3094) );
  AOI22_X1 U23277 ( .A1(n20632), .A2(n20335), .B1(n20334), .B2(n20631), .ZN(
        n20333) );
  INV_X1 U23278 ( .A(n20636), .ZN(n20530) );
  AOI22_X1 U23279 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20337), .B1(
        n20336), .B2(n20530), .ZN(n20332) );
  OAI211_X1 U23280 ( .C1(n20533), .C2(n20366), .A(n20333), .B(n20332), .ZN(
        P1_U3095) );
  AOI22_X1 U23281 ( .A1(n20640), .A2(n20335), .B1(n20334), .B2(n20637), .ZN(
        n20339) );
  INV_X1 U23282 ( .A(n20647), .ZN(n20576) );
  AOI22_X1 U23283 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20337), .B1(
        n20336), .B2(n20576), .ZN(n20338) );
  OAI211_X1 U23284 ( .C1(n20581), .C2(n20366), .A(n20339), .B(n20338), .ZN(
        P1_U3096) );
  AND2_X1 U23285 ( .A1(n12956), .A2(n12944), .ZN(n20444) );
  NAND3_X1 U23286 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20395), .A3(
        n20475), .ZN(n20367) );
  NOR2_X1 U23287 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20367), .ZN(
        n20361) );
  AOI21_X1 U23288 ( .B1(n20444), .B2(n12997), .A(n20361), .ZN(n20344) );
  INV_X1 U23289 ( .A(n20340), .ZN(n20341) );
  NAND2_X1 U23290 ( .A1(n20341), .A2(n20399), .ZN(n20483) );
  OAI22_X1 U23291 ( .A1(n20344), .A2(n20586), .B1(n20405), .B2(n20483), .ZN(
        n20362) );
  AOI22_X1 U23292 ( .A1(n20588), .A2(n20362), .B1(n20587), .B2(n20361), .ZN(
        n20348) );
  INV_X1 U23293 ( .A(n20342), .ZN(n20400) );
  INV_X1 U23294 ( .A(n20366), .ZN(n20343) );
  OAI21_X1 U23295 ( .B1(n20381), .B2(n20343), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20345) );
  NAND2_X1 U23296 ( .A1(n20345), .A2(n20344), .ZN(n20346) );
  AOI22_X1 U23297 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20363), .B1(
        n20381), .B2(n20595), .ZN(n20347) );
  OAI211_X1 U23298 ( .C1(n20598), .C2(n20366), .A(n20348), .B(n20347), .ZN(
        P1_U3097) );
  AOI22_X1 U23299 ( .A1(n20600), .A2(n20362), .B1(n20599), .B2(n20361), .ZN(
        n20350) );
  AOI22_X1 U23300 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20363), .B1(
        n20381), .B2(n20488), .ZN(n20349) );
  OAI211_X1 U23301 ( .C1(n20491), .C2(n20366), .A(n20350), .B(n20349), .ZN(
        P1_U3098) );
  AOI22_X1 U23302 ( .A1(n20606), .A2(n20362), .B1(n20605), .B2(n20361), .ZN(
        n20352) );
  AOI22_X1 U23303 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20363), .B1(
        n20381), .B2(n20607), .ZN(n20351) );
  OAI211_X1 U23304 ( .C1(n20610), .C2(n20366), .A(n20352), .B(n20351), .ZN(
        P1_U3099) );
  AOI22_X1 U23305 ( .A1(n20612), .A2(n20362), .B1(n20611), .B2(n20361), .ZN(
        n20354) );
  AOI22_X1 U23306 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20363), .B1(
        n20381), .B2(n20613), .ZN(n20353) );
  OAI211_X1 U23307 ( .C1(n20616), .C2(n20366), .A(n20354), .B(n20353), .ZN(
        P1_U3100) );
  AOI22_X1 U23308 ( .A1(n20362), .A2(n20618), .B1(n20617), .B2(n20361), .ZN(
        n20356) );
  AOI22_X1 U23309 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20363), .B1(
        n20381), .B2(n20619), .ZN(n20355) );
  OAI211_X1 U23310 ( .C1(n20622), .C2(n20366), .A(n20356), .B(n20355), .ZN(
        P1_U3101) );
  AOI22_X1 U23311 ( .A1(n20624), .A2(n20362), .B1(n20623), .B2(n20361), .ZN(
        n20358) );
  AOI22_X1 U23312 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20363), .B1(
        n20381), .B2(n20498), .ZN(n20357) );
  OAI211_X1 U23313 ( .C1(n20501), .C2(n20366), .A(n20358), .B(n20357), .ZN(
        P1_U3102) );
  AOI22_X1 U23314 ( .A1(n20632), .A2(n20362), .B1(n20631), .B2(n20361), .ZN(
        n20360) );
  AOI22_X1 U23315 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20363), .B1(
        n20381), .B2(n20633), .ZN(n20359) );
  OAI211_X1 U23316 ( .C1(n20636), .C2(n20366), .A(n20360), .B(n20359), .ZN(
        P1_U3103) );
  AOI22_X1 U23317 ( .A1(n20640), .A2(n20362), .B1(n20637), .B2(n20361), .ZN(
        n20365) );
  AOI22_X1 U23318 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20363), .B1(
        n20381), .B2(n20641), .ZN(n20364) );
  OAI211_X1 U23319 ( .C1(n20647), .C2(n20366), .A(n20365), .B(n20364), .ZN(
        P1_U3104) );
  NOR2_X1 U23320 ( .A1(n20742), .A2(n20367), .ZN(n20388) );
  AOI21_X1 U23321 ( .B1(n20444), .B2(n20512), .A(n20388), .ZN(n20368) );
  OAI22_X1 U23322 ( .A1(n20368), .A2(n20586), .B1(n20367), .B2(n20652), .ZN(
        n20389) );
  AOI22_X1 U23323 ( .A1(n20588), .A2(n20389), .B1(n20587), .B2(n20388), .ZN(
        n20374) );
  INV_X1 U23324 ( .A(n20367), .ZN(n20371) );
  OAI211_X1 U23325 ( .C1(n20450), .C2(n20515), .A(n20369), .B(n20368), .ZN(
        n20370) );
  OAI211_X1 U23326 ( .C1(n20369), .C2(n20371), .A(n20593), .B(n20370), .ZN(
        n20391) );
  INV_X1 U23327 ( .A(n20441), .ZN(n20390) );
  AOI22_X1 U23328 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20391), .B1(
        n20390), .B2(n20595), .ZN(n20373) );
  OAI211_X1 U23329 ( .C1(n20598), .C2(n20394), .A(n20374), .B(n20373), .ZN(
        P1_U3105) );
  AOI22_X1 U23330 ( .A1(n20600), .A2(n20389), .B1(n20599), .B2(n20388), .ZN(
        n20376) );
  AOI22_X1 U23331 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20391), .B1(
        n20381), .B2(n20601), .ZN(n20375) );
  OAI211_X1 U23332 ( .C1(n20604), .C2(n20441), .A(n20376), .B(n20375), .ZN(
        P1_U3106) );
  AOI22_X1 U23333 ( .A1(n20606), .A2(n20389), .B1(n20605), .B2(n20388), .ZN(
        n20378) );
  AOI22_X1 U23334 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20391), .B1(
        n20390), .B2(n20607), .ZN(n20377) );
  OAI211_X1 U23335 ( .C1(n20610), .C2(n20394), .A(n20378), .B(n20377), .ZN(
        P1_U3107) );
  AOI22_X1 U23336 ( .A1(n20612), .A2(n20389), .B1(n20611), .B2(n20388), .ZN(
        n20380) );
  AOI22_X1 U23337 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20391), .B1(
        n20381), .B2(n20561), .ZN(n20379) );
  OAI211_X1 U23338 ( .C1(n20564), .C2(n20441), .A(n20380), .B(n20379), .ZN(
        P1_U3108) );
  AOI22_X1 U23339 ( .A1(n20389), .A2(n20618), .B1(n20617), .B2(n20388), .ZN(
        n20383) );
  AOI22_X1 U23340 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20391), .B1(
        n20381), .B2(n20565), .ZN(n20382) );
  OAI211_X1 U23341 ( .C1(n20568), .C2(n20441), .A(n20383), .B(n20382), .ZN(
        P1_U3109) );
  AOI22_X1 U23342 ( .A1(n20624), .A2(n20389), .B1(n20623), .B2(n20388), .ZN(
        n20385) );
  AOI22_X1 U23343 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20391), .B1(
        n20390), .B2(n20498), .ZN(n20384) );
  OAI211_X1 U23344 ( .C1(n20501), .C2(n20394), .A(n20385), .B(n20384), .ZN(
        P1_U3110) );
  AOI22_X1 U23345 ( .A1(n20632), .A2(n20389), .B1(n20631), .B2(n20388), .ZN(
        n20387) );
  AOI22_X1 U23346 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20391), .B1(
        n20390), .B2(n20633), .ZN(n20386) );
  OAI211_X1 U23347 ( .C1(n20636), .C2(n20394), .A(n20387), .B(n20386), .ZN(
        P1_U3111) );
  AOI22_X1 U23348 ( .A1(n20640), .A2(n20389), .B1(n20637), .B2(n20388), .ZN(
        n20393) );
  AOI22_X1 U23349 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20391), .B1(
        n20390), .B2(n20641), .ZN(n20392) );
  OAI211_X1 U23350 ( .C1(n20647), .C2(n20394), .A(n20393), .B(n20392), .ZN(
        P1_U3112) );
  NAND3_X1 U23351 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n20395), .ZN(n20445) );
  NOR2_X1 U23352 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20445), .ZN(
        n20401) );
  INV_X1 U23353 ( .A(n20401), .ZN(n20434) );
  OAI22_X1 U23354 ( .A1(n20472), .A2(n20554), .B1(n20396), .B2(n20434), .ZN(
        n20397) );
  INV_X1 U23355 ( .A(n20397), .ZN(n20409) );
  NAND3_X1 U23356 ( .A1(n20472), .A2(n20441), .A3(n20738), .ZN(n20398) );
  NAND2_X1 U23357 ( .A1(n20398), .A2(n20477), .ZN(n20404) );
  NAND2_X1 U23358 ( .A1(n20444), .A2(n20543), .ZN(n20406) );
  OR2_X1 U23359 ( .A1(n20399), .A2(n20442), .ZN(n20545) );
  NAND2_X1 U23360 ( .A1(n20545), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20548) );
  OAI211_X1 U23361 ( .C1(n20481), .C2(n20401), .A(n20548), .B(n20400), .ZN(
        n20402) );
  AOI21_X1 U23362 ( .B1(n20404), .B2(n20406), .A(n20402), .ZN(n20403) );
  INV_X1 U23363 ( .A(n20404), .ZN(n20407) );
  OAI22_X1 U23364 ( .A1(n20407), .A2(n20406), .B1(n20405), .B2(n20545), .ZN(
        n20437) );
  AOI22_X1 U23365 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20438), .B1(
        n20588), .B2(n20437), .ZN(n20408) );
  OAI211_X1 U23366 ( .C1(n20598), .C2(n20441), .A(n20409), .B(n20408), .ZN(
        P1_U3113) );
  OAI22_X1 U23367 ( .A1(n20441), .A2(n20491), .B1(n20410), .B2(n20434), .ZN(
        n20411) );
  INV_X1 U23368 ( .A(n20411), .ZN(n20413) );
  AOI22_X1 U23369 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20438), .B1(
        n20600), .B2(n20437), .ZN(n20412) );
  OAI211_X1 U23370 ( .C1(n20604), .C2(n20472), .A(n20413), .B(n20412), .ZN(
        P1_U3114) );
  OAI22_X1 U23371 ( .A1(n20441), .A2(n20610), .B1(n20434), .B2(n20414), .ZN(
        n20415) );
  INV_X1 U23372 ( .A(n20415), .ZN(n20417) );
  AOI22_X1 U23373 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20438), .B1(
        n20606), .B2(n20437), .ZN(n20416) );
  OAI211_X1 U23374 ( .C1(n20560), .C2(n20472), .A(n20417), .B(n20416), .ZN(
        P1_U3115) );
  OAI22_X1 U23375 ( .A1(n20472), .A2(n20564), .B1(n20418), .B2(n20434), .ZN(
        n20419) );
  INV_X1 U23376 ( .A(n20419), .ZN(n20421) );
  AOI22_X1 U23377 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20438), .B1(
        n20612), .B2(n20437), .ZN(n20420) );
  OAI211_X1 U23378 ( .C1(n20616), .C2(n20441), .A(n20421), .B(n20420), .ZN(
        P1_U3116) );
  OAI22_X1 U23379 ( .A1(n20441), .A2(n20622), .B1(n20434), .B2(n20422), .ZN(
        n20423) );
  INV_X1 U23380 ( .A(n20423), .ZN(n20425) );
  AOI22_X1 U23381 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20438), .B1(
        n20618), .B2(n20437), .ZN(n20424) );
  OAI211_X1 U23382 ( .C1(n20568), .C2(n20472), .A(n20425), .B(n20424), .ZN(
        P1_U3117) );
  OAI22_X1 U23383 ( .A1(n20441), .A2(n20501), .B1(n20426), .B2(n20434), .ZN(
        n20427) );
  INV_X1 U23384 ( .A(n20427), .ZN(n20429) );
  AOI22_X1 U23385 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20438), .B1(
        n20624), .B2(n20437), .ZN(n20428) );
  OAI211_X1 U23386 ( .C1(n20630), .C2(n20472), .A(n20429), .B(n20428), .ZN(
        P1_U3118) );
  OAI22_X1 U23387 ( .A1(n20472), .A2(n20533), .B1(n20430), .B2(n20434), .ZN(
        n20431) );
  INV_X1 U23388 ( .A(n20431), .ZN(n20433) );
  AOI22_X1 U23389 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20438), .B1(
        n20632), .B2(n20437), .ZN(n20432) );
  OAI211_X1 U23390 ( .C1(n20636), .C2(n20441), .A(n20433), .B(n20432), .ZN(
        P1_U3119) );
  OAI22_X1 U23391 ( .A1(n20472), .A2(n20581), .B1(n20435), .B2(n20434), .ZN(
        n20436) );
  INV_X1 U23392 ( .A(n20436), .ZN(n20440) );
  AOI22_X1 U23393 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20438), .B1(
        n20640), .B2(n20437), .ZN(n20439) );
  OAI211_X1 U23394 ( .C1(n20647), .C2(n20441), .A(n20440), .B(n20439), .ZN(
        P1_U3120) );
  NOR2_X1 U23395 ( .A1(n20443), .A2(n20442), .ZN(n20466) );
  AOI21_X1 U23396 ( .B1(n20444), .B2(n20583), .A(n20466), .ZN(n20446) );
  OAI22_X1 U23397 ( .A1(n20446), .A2(n20586), .B1(n20445), .B2(n20652), .ZN(
        n20467) );
  AOI22_X1 U23398 ( .A1(n20588), .A2(n20467), .B1(n20587), .B2(n20466), .ZN(
        n20452) );
  INV_X1 U23399 ( .A(n20445), .ZN(n20448) );
  OAI211_X1 U23400 ( .C1(n20450), .C2(n20590), .A(n20738), .B(n20446), .ZN(
        n20447) );
  OAI211_X1 U23401 ( .C1(n20738), .C2(n20448), .A(n20593), .B(n20447), .ZN(
        n20469) );
  INV_X1 U23402 ( .A(n20509), .ZN(n20468) );
  AOI22_X1 U23403 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20469), .B1(
        n20468), .B2(n20595), .ZN(n20451) );
  OAI211_X1 U23404 ( .C1(n20598), .C2(n20472), .A(n20452), .B(n20451), .ZN(
        P1_U3121) );
  AOI22_X1 U23405 ( .A1(n20600), .A2(n20467), .B1(n20599), .B2(n20466), .ZN(
        n20454) );
  AOI22_X1 U23406 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20469), .B1(
        n20468), .B2(n20488), .ZN(n20453) );
  OAI211_X1 U23407 ( .C1(n20491), .C2(n20472), .A(n20454), .B(n20453), .ZN(
        P1_U3122) );
  AOI22_X1 U23408 ( .A1(n20606), .A2(n20467), .B1(n20605), .B2(n20466), .ZN(
        n20456) );
  INV_X1 U23409 ( .A(n20472), .ZN(n20463) );
  AOI22_X1 U23410 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20469), .B1(
        n20463), .B2(n20557), .ZN(n20455) );
  OAI211_X1 U23411 ( .C1(n20560), .C2(n20509), .A(n20456), .B(n20455), .ZN(
        P1_U3123) );
  AOI22_X1 U23412 ( .A1(n20612), .A2(n20467), .B1(n20611), .B2(n20466), .ZN(
        n20458) );
  AOI22_X1 U23413 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20469), .B1(
        n20468), .B2(n20613), .ZN(n20457) );
  OAI211_X1 U23414 ( .C1(n20616), .C2(n20472), .A(n20458), .B(n20457), .ZN(
        P1_U3124) );
  AOI22_X1 U23415 ( .A1(n20467), .A2(n20618), .B1(n20617), .B2(n20466), .ZN(
        n20460) );
  AOI22_X1 U23416 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20469), .B1(
        n20463), .B2(n20565), .ZN(n20459) );
  OAI211_X1 U23417 ( .C1(n20568), .C2(n20509), .A(n20460), .B(n20459), .ZN(
        P1_U3125) );
  AOI22_X1 U23418 ( .A1(n20624), .A2(n20467), .B1(n20623), .B2(n20466), .ZN(
        n20462) );
  AOI22_X1 U23419 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20469), .B1(
        n20463), .B2(n20625), .ZN(n20461) );
  OAI211_X1 U23420 ( .C1(n20630), .C2(n20509), .A(n20462), .B(n20461), .ZN(
        P1_U3126) );
  AOI22_X1 U23421 ( .A1(n20632), .A2(n20467), .B1(n20631), .B2(n20466), .ZN(
        n20465) );
  AOI22_X1 U23422 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20469), .B1(
        n20463), .B2(n20530), .ZN(n20464) );
  OAI211_X1 U23423 ( .C1(n20533), .C2(n20509), .A(n20465), .B(n20464), .ZN(
        P1_U3127) );
  AOI22_X1 U23424 ( .A1(n20640), .A2(n20467), .B1(n20637), .B2(n20466), .ZN(
        n20471) );
  AOI22_X1 U23425 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20469), .B1(
        n20468), .B2(n20641), .ZN(n20470) );
  OAI211_X1 U23426 ( .C1(n20647), .C2(n20472), .A(n20471), .B(n20470), .ZN(
        P1_U3128) );
  INV_X1 U23427 ( .A(n20473), .ZN(n20474) );
  NAND3_X1 U23428 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20475), .ZN(n20513) );
  NOR2_X1 U23429 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20513), .ZN(
        n20504) );
  AOI22_X1 U23430 ( .A1(n20536), .A2(n20595), .B1(n20587), .B2(n20504), .ZN(
        n20487) );
  INV_X1 U23431 ( .A(n20536), .ZN(n20476) );
  NAND3_X1 U23432 ( .A1(n20476), .A2(n20738), .A3(n20509), .ZN(n20478) );
  NAND2_X1 U23433 ( .A1(n20478), .A2(n20477), .ZN(n20482) );
  NOR2_X1 U23434 ( .A1(n12944), .A2(n20479), .ZN(n20584) );
  NAND2_X1 U23435 ( .A1(n20584), .A2(n12997), .ZN(n20484) );
  AOI22_X1 U23436 ( .A1(n20482), .A2(n20484), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20483), .ZN(n20480) );
  OAI211_X1 U23437 ( .C1(n20504), .C2(n20481), .A(n20549), .B(n20480), .ZN(
        n20506) );
  INV_X1 U23438 ( .A(n20482), .ZN(n20485) );
  OAI22_X1 U23439 ( .A1(n20485), .A2(n20484), .B1(n20544), .B2(n20483), .ZN(
        n20505) );
  AOI22_X1 U23440 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20506), .B1(
        n20588), .B2(n20505), .ZN(n20486) );
  OAI211_X1 U23441 ( .C1(n20598), .C2(n20509), .A(n20487), .B(n20486), .ZN(
        P1_U3129) );
  AOI22_X1 U23442 ( .A1(n20536), .A2(n20488), .B1(n20599), .B2(n20504), .ZN(
        n20490) );
  AOI22_X1 U23443 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20506), .B1(
        n20600), .B2(n20505), .ZN(n20489) );
  OAI211_X1 U23444 ( .C1(n20491), .C2(n20509), .A(n20490), .B(n20489), .ZN(
        P1_U3130) );
  AOI22_X1 U23445 ( .A1(n20536), .A2(n20607), .B1(n20504), .B2(n20605), .ZN(
        n20493) );
  AOI22_X1 U23446 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20506), .B1(
        n20606), .B2(n20505), .ZN(n20492) );
  OAI211_X1 U23447 ( .C1(n20610), .C2(n20509), .A(n20493), .B(n20492), .ZN(
        P1_U3131) );
  AOI22_X1 U23448 ( .A1(n20536), .A2(n20613), .B1(n20611), .B2(n20504), .ZN(
        n20495) );
  AOI22_X1 U23449 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20506), .B1(
        n20612), .B2(n20505), .ZN(n20494) );
  OAI211_X1 U23450 ( .C1(n20616), .C2(n20509), .A(n20495), .B(n20494), .ZN(
        P1_U3132) );
  AOI22_X1 U23451 ( .A1(n20536), .A2(n20619), .B1(n20504), .B2(n20617), .ZN(
        n20497) );
  AOI22_X1 U23452 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20506), .B1(
        n20618), .B2(n20505), .ZN(n20496) );
  OAI211_X1 U23453 ( .C1(n20622), .C2(n20509), .A(n20497), .B(n20496), .ZN(
        P1_U3133) );
  AOI22_X1 U23454 ( .A1(n20536), .A2(n20498), .B1(n20623), .B2(n20504), .ZN(
        n20500) );
  AOI22_X1 U23455 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20506), .B1(
        n20624), .B2(n20505), .ZN(n20499) );
  OAI211_X1 U23456 ( .C1(n20501), .C2(n20509), .A(n20500), .B(n20499), .ZN(
        P1_U3134) );
  AOI22_X1 U23457 ( .A1(n20536), .A2(n20633), .B1(n20631), .B2(n20504), .ZN(
        n20503) );
  AOI22_X1 U23458 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20506), .B1(
        n20632), .B2(n20505), .ZN(n20502) );
  OAI211_X1 U23459 ( .C1(n20636), .C2(n20509), .A(n20503), .B(n20502), .ZN(
        P1_U3135) );
  AOI22_X1 U23460 ( .A1(n20536), .A2(n20641), .B1(n20637), .B2(n20504), .ZN(
        n20508) );
  AOI22_X1 U23461 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20506), .B1(
        n20640), .B2(n20505), .ZN(n20507) );
  OAI211_X1 U23462 ( .C1(n20647), .C2(n20509), .A(n20508), .B(n20507), .ZN(
        P1_U3136) );
  NOR2_X1 U23463 ( .A1(n20742), .A2(n20513), .ZN(n20534) );
  AOI21_X1 U23464 ( .B1(n20584), .B2(n20512), .A(n20534), .ZN(n20514) );
  OAI22_X1 U23465 ( .A1(n20514), .A2(n20586), .B1(n20513), .B2(n20652), .ZN(
        n20535) );
  AOI22_X1 U23466 ( .A1(n20588), .A2(n20535), .B1(n20587), .B2(n20534), .ZN(
        n20519) );
  INV_X1 U23467 ( .A(n20513), .ZN(n20517) );
  INV_X1 U23468 ( .A(n20542), .ZN(n20591) );
  OAI211_X1 U23469 ( .C1(n20591), .C2(n20515), .A(n20369), .B(n20514), .ZN(
        n20516) );
  OAI211_X1 U23470 ( .C1(n20738), .C2(n20517), .A(n20593), .B(n20516), .ZN(
        n20537) );
  AOI22_X1 U23471 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20537), .B1(
        n20536), .B2(n20551), .ZN(n20518) );
  OAI211_X1 U23472 ( .C1(n20554), .C2(n20573), .A(n20519), .B(n20518), .ZN(
        P1_U3137) );
  AOI22_X1 U23473 ( .A1(n20600), .A2(n20535), .B1(n20599), .B2(n20534), .ZN(
        n20521) );
  AOI22_X1 U23474 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20537), .B1(
        n20536), .B2(n20601), .ZN(n20520) );
  OAI211_X1 U23475 ( .C1(n20604), .C2(n20573), .A(n20521), .B(n20520), .ZN(
        P1_U3138) );
  AOI22_X1 U23476 ( .A1(n20606), .A2(n20535), .B1(n20605), .B2(n20534), .ZN(
        n20523) );
  AOI22_X1 U23477 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20537), .B1(
        n20536), .B2(n20557), .ZN(n20522) );
  OAI211_X1 U23478 ( .C1(n20560), .C2(n20573), .A(n20523), .B(n20522), .ZN(
        P1_U3139) );
  AOI22_X1 U23479 ( .A1(n20612), .A2(n20535), .B1(n20611), .B2(n20534), .ZN(
        n20525) );
  AOI22_X1 U23480 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20537), .B1(
        n20536), .B2(n20561), .ZN(n20524) );
  OAI211_X1 U23481 ( .C1(n20564), .C2(n20573), .A(n20525), .B(n20524), .ZN(
        P1_U3140) );
  AOI22_X1 U23482 ( .A1(n20535), .A2(n20618), .B1(n20617), .B2(n20534), .ZN(
        n20527) );
  AOI22_X1 U23483 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20537), .B1(
        n20536), .B2(n20565), .ZN(n20526) );
  OAI211_X1 U23484 ( .C1(n20568), .C2(n20573), .A(n20527), .B(n20526), .ZN(
        P1_U3141) );
  AOI22_X1 U23485 ( .A1(n20624), .A2(n20535), .B1(n20623), .B2(n20534), .ZN(
        n20529) );
  AOI22_X1 U23486 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20537), .B1(
        n20536), .B2(n20625), .ZN(n20528) );
  OAI211_X1 U23487 ( .C1(n20630), .C2(n20573), .A(n20529), .B(n20528), .ZN(
        P1_U3142) );
  AOI22_X1 U23488 ( .A1(n20632), .A2(n20535), .B1(n20631), .B2(n20534), .ZN(
        n20532) );
  AOI22_X1 U23489 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20537), .B1(
        n20536), .B2(n20530), .ZN(n20531) );
  OAI211_X1 U23490 ( .C1(n20533), .C2(n20573), .A(n20532), .B(n20531), .ZN(
        P1_U3143) );
  AOI22_X1 U23491 ( .A1(n20640), .A2(n20535), .B1(n20637), .B2(n20534), .ZN(
        n20539) );
  AOI22_X1 U23492 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20537), .B1(
        n20536), .B2(n20576), .ZN(n20538) );
  OAI211_X1 U23493 ( .C1(n20581), .C2(n20573), .A(n20539), .B(n20538), .ZN(
        P1_U3144) );
  INV_X1 U23494 ( .A(n20540), .ZN(n20541) );
  NAND2_X1 U23495 ( .A1(n20584), .A2(n20543), .ZN(n20546) );
  OAI22_X1 U23496 ( .A1(n20546), .A2(n20586), .B1(n20545), .B2(n20544), .ZN(
        n20575) );
  NOR2_X1 U23497 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20585), .ZN(
        n20574) );
  AOI22_X1 U23498 ( .A1(n20588), .A2(n20575), .B1(n20587), .B2(n20574), .ZN(
        n20553) );
  INV_X1 U23499 ( .A(n20646), .ZN(n20626) );
  OAI21_X1 U23500 ( .B1(n20577), .B2(n20626), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20547) );
  AOI21_X1 U23501 ( .B1(n20547), .B2(n20546), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20550) );
  AOI22_X1 U23502 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20551), .ZN(n20552) );
  OAI211_X1 U23503 ( .C1(n20554), .C2(n20646), .A(n20553), .B(n20552), .ZN(
        P1_U3145) );
  AOI22_X1 U23504 ( .A1(n20600), .A2(n20575), .B1(n20599), .B2(n20574), .ZN(
        n20556) );
  AOI22_X1 U23505 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20601), .ZN(n20555) );
  OAI211_X1 U23506 ( .C1(n20604), .C2(n20646), .A(n20556), .B(n20555), .ZN(
        P1_U3146) );
  AOI22_X1 U23507 ( .A1(n20606), .A2(n20575), .B1(n20605), .B2(n20574), .ZN(
        n20559) );
  AOI22_X1 U23508 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20557), .ZN(n20558) );
  OAI211_X1 U23509 ( .C1(n20560), .C2(n20646), .A(n20559), .B(n20558), .ZN(
        P1_U3147) );
  AOI22_X1 U23510 ( .A1(n20612), .A2(n20575), .B1(n20611), .B2(n20574), .ZN(
        n20563) );
  AOI22_X1 U23511 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20561), .ZN(n20562) );
  OAI211_X1 U23512 ( .C1(n20564), .C2(n20646), .A(n20563), .B(n20562), .ZN(
        P1_U3148) );
  AOI22_X1 U23513 ( .A1(n20575), .A2(n20618), .B1(n20617), .B2(n20574), .ZN(
        n20567) );
  AOI22_X1 U23514 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20565), .ZN(n20566) );
  OAI211_X1 U23515 ( .C1(n20568), .C2(n20646), .A(n20567), .B(n20566), .ZN(
        P1_U3149) );
  AOI22_X1 U23516 ( .A1(n20624), .A2(n20575), .B1(n20623), .B2(n20574), .ZN(
        n20570) );
  AOI22_X1 U23517 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20625), .ZN(n20569) );
  OAI211_X1 U23518 ( .C1(n20630), .C2(n20646), .A(n20570), .B(n20569), .ZN(
        P1_U3150) );
  AOI22_X1 U23519 ( .A1(n20632), .A2(n20575), .B1(n20631), .B2(n20574), .ZN(
        n20572) );
  AOI22_X1 U23520 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20578), .B1(
        n20626), .B2(n20633), .ZN(n20571) );
  OAI211_X1 U23521 ( .C1(n20636), .C2(n20573), .A(n20572), .B(n20571), .ZN(
        P1_U3151) );
  AOI22_X1 U23522 ( .A1(n20640), .A2(n20575), .B1(n20637), .B2(n20574), .ZN(
        n20580) );
  AOI22_X1 U23523 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20576), .ZN(n20579) );
  OAI211_X1 U23524 ( .C1(n20581), .C2(n20646), .A(n20580), .B(n20579), .ZN(
        P1_U3152) );
  INV_X1 U23525 ( .A(n20582), .ZN(n20638) );
  AOI21_X1 U23526 ( .B1(n20584), .B2(n20583), .A(n20638), .ZN(n20589) );
  OAI22_X1 U23527 ( .A1(n20589), .A2(n20586), .B1(n20585), .B2(n20652), .ZN(
        n20639) );
  AOI22_X1 U23528 ( .A1(n20588), .A2(n20639), .B1(n20638), .B2(n20587), .ZN(
        n20597) );
  OAI211_X1 U23529 ( .C1(n20591), .C2(n20590), .A(n20369), .B(n20589), .ZN(
        n20592) );
  OAI211_X1 U23530 ( .C1(n20594), .C2(n20369), .A(n20593), .B(n20592), .ZN(
        n20643) );
  AOI22_X1 U23531 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20643), .B1(
        n20642), .B2(n20595), .ZN(n20596) );
  OAI211_X1 U23532 ( .C1(n20598), .C2(n20646), .A(n20597), .B(n20596), .ZN(
        P1_U3153) );
  AOI22_X1 U23533 ( .A1(n20600), .A2(n20639), .B1(n20638), .B2(n20599), .ZN(
        n20603) );
  AOI22_X1 U23534 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20643), .B1(
        n20626), .B2(n20601), .ZN(n20602) );
  OAI211_X1 U23535 ( .C1(n20604), .C2(n20629), .A(n20603), .B(n20602), .ZN(
        P1_U3154) );
  AOI22_X1 U23536 ( .A1(n20606), .A2(n20639), .B1(n20638), .B2(n20605), .ZN(
        n20609) );
  AOI22_X1 U23537 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20643), .B1(
        n20642), .B2(n20607), .ZN(n20608) );
  OAI211_X1 U23538 ( .C1(n20610), .C2(n20646), .A(n20609), .B(n20608), .ZN(
        P1_U3155) );
  AOI22_X1 U23539 ( .A1(n20612), .A2(n20639), .B1(n20638), .B2(n20611), .ZN(
        n20615) );
  AOI22_X1 U23540 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20643), .B1(
        n20642), .B2(n20613), .ZN(n20614) );
  OAI211_X1 U23541 ( .C1(n20616), .C2(n20646), .A(n20615), .B(n20614), .ZN(
        P1_U3156) );
  AOI22_X1 U23542 ( .A1(n20639), .A2(n20618), .B1(n20638), .B2(n20617), .ZN(
        n20621) );
  AOI22_X1 U23543 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20643), .B1(
        n20642), .B2(n20619), .ZN(n20620) );
  OAI211_X1 U23544 ( .C1(n20622), .C2(n20646), .A(n20621), .B(n20620), .ZN(
        P1_U3157) );
  AOI22_X1 U23545 ( .A1(n20624), .A2(n20639), .B1(n20638), .B2(n20623), .ZN(
        n20628) );
  AOI22_X1 U23546 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20643), .B1(
        n20626), .B2(n20625), .ZN(n20627) );
  OAI211_X1 U23547 ( .C1(n20630), .C2(n20629), .A(n20628), .B(n20627), .ZN(
        P1_U3158) );
  AOI22_X1 U23548 ( .A1(n20632), .A2(n20639), .B1(n20638), .B2(n20631), .ZN(
        n20635) );
  AOI22_X1 U23549 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20643), .B1(
        n20642), .B2(n20633), .ZN(n20634) );
  OAI211_X1 U23550 ( .C1(n20636), .C2(n20646), .A(n20635), .B(n20634), .ZN(
        P1_U3159) );
  AOI22_X1 U23551 ( .A1(n20640), .A2(n20639), .B1(n20638), .B2(n20637), .ZN(
        n20645) );
  AOI22_X1 U23552 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20643), .B1(
        n20642), .B2(n20641), .ZN(n20644) );
  OAI211_X1 U23553 ( .C1(n20647), .C2(n20646), .A(n20645), .B(n20644), .ZN(
        P1_U3160) );
  NOR2_X1 U23554 ( .A1(n20649), .A2(n20648), .ZN(n20653) );
  INV_X1 U23555 ( .A(n20650), .ZN(n20651) );
  OAI21_X1 U23556 ( .B1(n20653), .B2(n20652), .A(n20651), .ZN(P1_U3163) );
  INV_X1 U23557 ( .A(n20733), .ZN(n20729) );
  AND2_X1 U23558 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20729), .ZN(
        P1_U3164) );
  AND2_X1 U23559 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20729), .ZN(
        P1_U3165) );
  AND2_X1 U23560 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20729), .ZN(
        P1_U3166) );
  AND2_X1 U23561 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20729), .ZN(
        P1_U3167) );
  AND2_X1 U23562 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20729), .ZN(
        P1_U3168) );
  AND2_X1 U23563 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20729), .ZN(
        P1_U3169) );
  AND2_X1 U23564 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20729), .ZN(
        P1_U3170) );
  AND2_X1 U23565 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20729), .ZN(
        P1_U3171) );
  AND2_X1 U23566 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20729), .ZN(
        P1_U3172) );
  AND2_X1 U23567 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20729), .ZN(
        P1_U3173) );
  AND2_X1 U23568 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20729), .ZN(
        P1_U3174) );
  AND2_X1 U23569 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20729), .ZN(
        P1_U3175) );
  AND2_X1 U23570 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20729), .ZN(
        P1_U3176) );
  AND2_X1 U23571 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20729), .ZN(
        P1_U3177) );
  AND2_X1 U23572 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20729), .ZN(
        P1_U3178) );
  AND2_X1 U23573 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20729), .ZN(
        P1_U3179) );
  AND2_X1 U23574 ( .A1(n20729), .A2(P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(
        P1_U3180) );
  AND2_X1 U23575 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20729), .ZN(
        P1_U3181) );
  AND2_X1 U23576 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20729), .ZN(
        P1_U3182) );
  AND2_X1 U23577 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20729), .ZN(
        P1_U3183) );
  AND2_X1 U23578 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20729), .ZN(
        P1_U3184) );
  AND2_X1 U23579 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20729), .ZN(
        P1_U3185) );
  AND2_X1 U23580 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20729), .ZN(P1_U3186) );
  AND2_X1 U23581 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20729), .ZN(P1_U3187) );
  AND2_X1 U23582 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20729), .ZN(P1_U3188) );
  AND2_X1 U23583 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20729), .ZN(P1_U3189) );
  AND2_X1 U23584 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20729), .ZN(P1_U3190) );
  AND2_X1 U23585 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20729), .ZN(P1_U3191) );
  AND2_X1 U23586 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20729), .ZN(P1_U3192) );
  AND2_X1 U23587 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20729), .ZN(P1_U3193) );
  NAND2_X1 U23588 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20662), .ZN(n20661) );
  INV_X1 U23589 ( .A(n20661), .ZN(n20657) );
  INV_X2 U23590 ( .A(n20753), .ZN(n20768) );
  OAI21_X1 U23591 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20663), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20654) );
  AOI211_X1 U23592 ( .C1(HOLD), .C2(P1_STATE_REG_1__SCAN_IN), .A(n20655), .B(
        n20654), .ZN(n20656) );
  OAI22_X1 U23593 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20657), .B1(n20768), 
        .B2(n20656), .ZN(P1_U3194) );
  INV_X1 U23594 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20766) );
  OAI211_X1 U23595 ( .C1(NA), .C2(n20659), .A(P1_STATE_REG_1__SCAN_IN), .B(
        n20658), .ZN(n20660) );
  OAI211_X1 U23596 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20766), .A(
        P1_STATE_REG_0__SCAN_IN), .B(n20660), .ZN(n20667) );
  OAI211_X1 U23597 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n20663), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20661), .ZN(n20666) );
  INV_X1 U23598 ( .A(n20662), .ZN(n20664) );
  NAND4_X1 U23599 ( .A1(P1_REQUESTPENDING_REG_SCAN_IN), .A2(
        P1_STATE_REG_0__SCAN_IN), .A3(n20664), .A4(n20663), .ZN(n20665) );
  OAI211_X1 U23600 ( .C1(n20668), .C2(n20667), .A(n20666), .B(n20665), .ZN(
        P1_U3196) );
  NAND2_X1 U23601 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20768), .ZN(n20721) );
  NOR2_X1 U23602 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20753), .ZN(n20714) );
  AOI22_X1 U23603 ( .A1(P1_ADDRESS_REG_0__SCAN_IN), .A2(n20753), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n20714), .ZN(n20669) );
  OAI21_X1 U23604 ( .B1(n20744), .B2(n20721), .A(n20669), .ZN(P1_U3197) );
  INV_X1 U23605 ( .A(n20714), .ZN(n20717) );
  INV_X1 U23606 ( .A(n20721), .ZN(n20715) );
  AOI22_X1 U23607 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n20753), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n20715), .ZN(n20670) );
  OAI21_X1 U23608 ( .B1(n13162), .B2(n20717), .A(n20670), .ZN(P1_U3198) );
  INV_X1 U23609 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20846) );
  OAI222_X1 U23610 ( .A1(n20721), .A2(n13162), .B1(n20846), .B2(n20768), .C1(
        n20672), .C2(n20717), .ZN(P1_U3199) );
  OAI222_X1 U23611 ( .A1(n20721), .A2(n20672), .B1(n20671), .B2(n20768), .C1(
        n20674), .C2(n20717), .ZN(P1_U3200) );
  INV_X1 U23612 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20673) );
  OAI222_X1 U23613 ( .A1(n20721), .A2(n20674), .B1(n20673), .B2(n20768), .C1(
        n20676), .C2(n20717), .ZN(P1_U3201) );
  INV_X1 U23614 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n20675) );
  OAI222_X1 U23615 ( .A1(n20721), .A2(n20676), .B1(n20675), .B2(n20768), .C1(
        n20678), .C2(n20717), .ZN(P1_U3202) );
  INV_X1 U23616 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20677) );
  OAI222_X1 U23617 ( .A1(n20721), .A2(n20678), .B1(n20677), .B2(n20768), .C1(
        n20679), .C2(n20717), .ZN(P1_U3203) );
  INV_X1 U23618 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20680) );
  OAI222_X1 U23619 ( .A1(n20717), .A2(n13654), .B1(n20680), .B2(n20768), .C1(
        n20679), .C2(n20721), .ZN(P1_U3204) );
  INV_X1 U23620 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20681) );
  OAI222_X1 U23621 ( .A1(n20721), .A2(n13654), .B1(n20681), .B2(n20768), .C1(
        n20683), .C2(n20717), .ZN(P1_U3205) );
  AOI22_X1 U23622 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(n20753), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n20714), .ZN(n20682) );
  OAI21_X1 U23623 ( .B1(n20683), .B2(n20721), .A(n20682), .ZN(P1_U3206) );
  AOI22_X1 U23624 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n20753), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n20715), .ZN(n20684) );
  OAI21_X1 U23625 ( .B1(n20686), .B2(n20717), .A(n20684), .ZN(P1_U3207) );
  INV_X1 U23626 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n20685) );
  OAI222_X1 U23627 ( .A1(n20721), .A2(n20686), .B1(n20685), .B2(n20768), .C1(
        n20688), .C2(n20717), .ZN(P1_U3208) );
  AOI22_X1 U23628 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20753), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20714), .ZN(n20687) );
  OAI21_X1 U23629 ( .B1(n20688), .B2(n20721), .A(n20687), .ZN(P1_U3209) );
  AOI22_X1 U23630 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n20753), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20715), .ZN(n20689) );
  OAI21_X1 U23631 ( .B1(n20691), .B2(n20717), .A(n20689), .ZN(P1_U3210) );
  INV_X1 U23632 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n20690) );
  OAI222_X1 U23633 ( .A1(n20721), .A2(n20691), .B1(n20690), .B2(n20768), .C1(
        n20693), .C2(n20717), .ZN(P1_U3211) );
  AOI22_X1 U23634 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20753), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20714), .ZN(n20692) );
  OAI21_X1 U23635 ( .B1(n20693), .B2(n20721), .A(n20692), .ZN(P1_U3212) );
  AOI22_X1 U23636 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20753), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20715), .ZN(n20694) );
  OAI21_X1 U23637 ( .B1(n20696), .B2(n20717), .A(n20694), .ZN(P1_U3213) );
  INV_X1 U23638 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20695) );
  OAI222_X1 U23639 ( .A1(n20721), .A2(n20696), .B1(n20695), .B2(n20768), .C1(
        n20698), .C2(n20717), .ZN(P1_U3214) );
  AOI22_X1 U23640 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20753), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20714), .ZN(n20697) );
  OAI21_X1 U23641 ( .B1(n20698), .B2(n20721), .A(n20697), .ZN(P1_U3215) );
  AOI22_X1 U23642 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n20753), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20715), .ZN(n20699) );
  OAI21_X1 U23643 ( .B1(n20701), .B2(n20717), .A(n20699), .ZN(P1_U3216) );
  INV_X1 U23644 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20700) );
  OAI222_X1 U23645 ( .A1(n20721), .A2(n20701), .B1(n20700), .B2(n20768), .C1(
        n20703), .C2(n20717), .ZN(P1_U3217) );
  INV_X1 U23646 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20702) );
  OAI222_X1 U23647 ( .A1(n20721), .A2(n20703), .B1(n20702), .B2(n20768), .C1(
        n20908), .C2(n20717), .ZN(P1_U3218) );
  INV_X1 U23648 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n20704) );
  OAI222_X1 U23649 ( .A1(n20721), .A2(n20908), .B1(n20704), .B2(n20768), .C1(
        n14143), .C2(n20717), .ZN(P1_U3219) );
  INV_X1 U23650 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20705) );
  OAI222_X1 U23651 ( .A1(n20721), .A2(n14143), .B1(n20705), .B2(n20768), .C1(
        n20707), .C2(n20717), .ZN(P1_U3220) );
  INV_X1 U23652 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20706) );
  INV_X1 U23653 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20709) );
  OAI222_X1 U23654 ( .A1(n20721), .A2(n20707), .B1(n20706), .B2(n20768), .C1(
        n20709), .C2(n20717), .ZN(P1_U3221) );
  INV_X1 U23655 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20708) );
  OAI222_X1 U23656 ( .A1(n20721), .A2(n20709), .B1(n20708), .B2(n20768), .C1(
        n20712), .C2(n20717), .ZN(P1_U3222) );
  INV_X1 U23657 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n20711) );
  OAI222_X1 U23658 ( .A1(n20721), .A2(n20712), .B1(n20711), .B2(n20768), .C1(
        n20710), .C2(n20717), .ZN(P1_U3223) );
  AOI222_X1 U23659 ( .A1(n20715), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20753), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20714), .ZN(n20713) );
  INV_X1 U23660 ( .A(n20713), .ZN(P1_U3224) );
  AOI222_X1 U23661 ( .A1(n20715), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20753), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(n20714), .ZN(n20716) );
  INV_X1 U23662 ( .A(n20716), .ZN(P1_U3225) );
  INV_X1 U23663 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20719) );
  OAI222_X1 U23664 ( .A1(n20721), .A2(n20720), .B1(n20719), .B2(n20768), .C1(
        n20718), .C2(n20717), .ZN(P1_U3226) );
  INV_X1 U23665 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20722) );
  AOI22_X1 U23666 ( .A1(n20768), .A2(n20723), .B1(n20722), .B2(n20753), .ZN(
        P1_U3458) );
  INV_X1 U23667 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20746) );
  INV_X1 U23668 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20724) );
  AOI22_X1 U23669 ( .A1(n20768), .A2(n20746), .B1(n20724), .B2(n20753), .ZN(
        P1_U3459) );
  INV_X1 U23670 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20725) );
  AOI22_X1 U23671 ( .A1(n20768), .A2(n20726), .B1(n20725), .B2(n20753), .ZN(
        P1_U3460) );
  INV_X1 U23672 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20752) );
  INV_X1 U23673 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20727) );
  AOI22_X1 U23674 ( .A1(n20768), .A2(n20752), .B1(n20727), .B2(n20753), .ZN(
        P1_U3461) );
  INV_X1 U23675 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20730) );
  INV_X1 U23676 ( .A(n20731), .ZN(n20728) );
  AOI21_X1 U23677 ( .B1(n20730), .B2(n20729), .A(n20728), .ZN(P1_U3464) );
  OAI21_X1 U23678 ( .B1(n20733), .B2(n20732), .A(n20731), .ZN(P1_U3465) );
  OAI21_X1 U23679 ( .B1(n20736), .B2(n20735), .A(n20734), .ZN(n20737) );
  AOI21_X1 U23680 ( .B1(n20739), .B2(n20738), .A(n20737), .ZN(n20741) );
  AOI22_X1 U23681 ( .A1(n20743), .A2(n20742), .B1(n20741), .B2(n20740), .ZN(
        P1_U3478) );
  AOI21_X1 U23682 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20745) );
  AOI22_X1 U23683 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20745), .B2(n20744), .ZN(n20747) );
  AOI22_X1 U23684 ( .A1(n20748), .A2(n20747), .B1(n20746), .B2(n20751), .ZN(
        P1_U3481) );
  NOR2_X1 U23685 ( .A1(n20751), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20749) );
  AOI22_X1 U23686 ( .A1(n20752), .A2(n20751), .B1(n20750), .B2(n20749), .ZN(
        P1_U3482) );
  AOI22_X1 U23687 ( .A1(n20768), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20754), 
        .B2(n20753), .ZN(P1_U3483) );
  INV_X1 U23688 ( .A(n20755), .ZN(n20756) );
  OAI211_X1 U23689 ( .C1(n20759), .C2(n20758), .A(n20757), .B(n20756), .ZN(
        n20767) );
  NOR2_X1 U23690 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20760), .ZN(n20765) );
  OAI211_X1 U23691 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20762), .A(n20761), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20763) );
  NAND2_X1 U23692 ( .A1(n20767), .A2(n20763), .ZN(n20764) );
  OAI22_X1 U23693 ( .A1(n20767), .A2(n20766), .B1(n20765), .B2(n20764), .ZN(
        P1_U3485) );
  MUX2_X1 U23694 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n20768), .Z(P1_U3486) );
  NAND4_X1 U23695 ( .A1(keyinput29), .A2(keyinput19), .A3(keyinput47), .A4(
        keyinput56), .ZN(n20791) );
  NOR3_X1 U23696 ( .A1(keyinput52), .A2(keyinput7), .A3(keyinput54), .ZN(
        n20772) );
  NOR4_X1 U23697 ( .A1(keyinput9), .A2(keyinput49), .A3(keyinput36), .A4(
        keyinput18), .ZN(n20771) );
  INV_X1 U23698 ( .A(keyinput1), .ZN(n20769) );
  NOR4_X1 U23699 ( .A1(keyinput60), .A2(keyinput50), .A3(keyinput22), .A4(
        n20769), .ZN(n20770) );
  NAND4_X1 U23700 ( .A1(keyinput58), .A2(n20772), .A3(n20771), .A4(n20770), 
        .ZN(n20790) );
  NOR4_X1 U23701 ( .A1(keyinput63), .A2(keyinput62), .A3(keyinput38), .A4(
        keyinput34), .ZN(n20776) );
  NOR4_X1 U23702 ( .A1(keyinput30), .A2(keyinput27), .A3(keyinput23), .A4(
        keyinput14), .ZN(n20775) );
  NOR4_X1 U23703 ( .A1(keyinput10), .A2(keyinput5), .A3(keyinput13), .A4(
        keyinput32), .ZN(n20774) );
  NOR4_X1 U23704 ( .A1(keyinput8), .A2(keyinput20), .A3(keyinput12), .A4(
        keyinput24), .ZN(n20773) );
  NAND4_X1 U23705 ( .A1(n20776), .A2(n20775), .A3(n20774), .A4(n20773), .ZN(
        n20789) );
  NOR3_X1 U23706 ( .A1(keyinput28), .A2(keyinput0), .A3(keyinput31), .ZN(
        n20787) );
  NAND3_X1 U23707 ( .A1(keyinput40), .A2(keyinput43), .A3(keyinput6), .ZN(
        n20780) );
  NOR3_X1 U23708 ( .A1(keyinput2), .A2(keyinput42), .A3(keyinput17), .ZN(
        n20778) );
  NOR3_X1 U23709 ( .A1(keyinput15), .A2(keyinput48), .A3(keyinput21), .ZN(
        n20777) );
  NAND4_X1 U23710 ( .A1(keyinput61), .A2(n20778), .A3(keyinput55), .A4(n20777), 
        .ZN(n20779) );
  NOR3_X1 U23711 ( .A1(keyinput45), .A2(n20780), .A3(n20779), .ZN(n20786) );
  NAND4_X1 U23712 ( .A1(keyinput44), .A2(keyinput59), .A3(keyinput51), .A4(
        keyinput39), .ZN(n20784) );
  NAND4_X1 U23713 ( .A1(keyinput26), .A2(keyinput35), .A3(keyinput11), .A4(
        keyinput3), .ZN(n20783) );
  NAND4_X1 U23714 ( .A1(keyinput33), .A2(keyinput41), .A3(keyinput37), .A4(
        keyinput53), .ZN(n20782) );
  NAND4_X1 U23715 ( .A1(keyinput57), .A2(keyinput25), .A3(keyinput16), .A4(
        keyinput4), .ZN(n20781) );
  NOR4_X1 U23716 ( .A1(n20784), .A2(n20783), .A3(n20782), .A4(n20781), .ZN(
        n20785) );
  NAND4_X1 U23717 ( .A1(keyinput46), .A2(n20787), .A3(n20786), .A4(n20785), 
        .ZN(n20788) );
  NOR4_X1 U23718 ( .A1(n20791), .A2(n20790), .A3(n20789), .A4(n20788), .ZN(
        n20924) );
  OAI22_X1 U23719 ( .A1(n20794), .A2(keyinput29), .B1(n20793), .B2(keyinput19), 
        .ZN(n20792) );
  AOI221_X1 U23720 ( .B1(n20794), .B2(keyinput29), .C1(keyinput19), .C2(n20793), .A(n20792), .ZN(n20807) );
  OAI22_X1 U23721 ( .A1(n20797), .A2(keyinput52), .B1(n20796), .B2(keyinput58), 
        .ZN(n20795) );
  AOI221_X1 U23722 ( .B1(n20797), .B2(keyinput52), .C1(keyinput58), .C2(n20796), .A(n20795), .ZN(n20806) );
  INV_X1 U23723 ( .A(keyinput56), .ZN(n20799) );
  OAI22_X1 U23724 ( .A1(keyinput47), .A2(n20800), .B1(n20799), .B2(
        P3_LWORD_REG_1__SCAN_IN), .ZN(n20798) );
  AOI221_X1 U23725 ( .B1(n20800), .B2(keyinput47), .C1(n20799), .C2(
        P3_LWORD_REG_1__SCAN_IN), .A(n20798), .ZN(n20805) );
  XOR2_X1 U23726 ( .A(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B(keyinput54), .Z(
        n20803) );
  INV_X1 U23727 ( .A(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n20801) );
  XNOR2_X1 U23728 ( .A(keyinput7), .B(n20801), .ZN(n20802) );
  NOR2_X1 U23729 ( .A1(n20803), .A2(n20802), .ZN(n20804) );
  NAND4_X1 U23730 ( .A1(n20807), .A2(n20806), .A3(n20805), .A4(n20804), .ZN(
        n20923) );
  INV_X1 U23731 ( .A(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n20809) );
  AOI22_X1 U23732 ( .A1(n20810), .A2(keyinput40), .B1(n20809), .B2(keyinput43), 
        .ZN(n20808) );
  OAI221_X1 U23733 ( .B1(n20810), .B2(keyinput40), .C1(n20809), .C2(keyinput43), .A(n20808), .ZN(n20822) );
  INV_X1 U23734 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n20812) );
  AOI22_X1 U23735 ( .A1(n20812), .A2(keyinput6), .B1(keyinput45), .B2(n11940), 
        .ZN(n20811) );
  OAI221_X1 U23736 ( .B1(n20812), .B2(keyinput6), .C1(n11940), .C2(keyinput45), 
        .A(n20811), .ZN(n20821) );
  AOI22_X1 U23737 ( .A1(n20815), .A2(keyinput28), .B1(n20814), .B2(keyinput0), 
        .ZN(n20813) );
  OAI221_X1 U23738 ( .B1(n20815), .B2(keyinput28), .C1(n20814), .C2(keyinput0), 
        .A(n20813), .ZN(n20820) );
  INV_X1 U23739 ( .A(READY1), .ZN(n20817) );
  AOI22_X1 U23740 ( .A1(n20818), .A2(keyinput46), .B1(n20817), .B2(keyinput31), 
        .ZN(n20816) );
  OAI221_X1 U23741 ( .B1(n20818), .B2(keyinput46), .C1(n20817), .C2(keyinput31), .A(n20816), .ZN(n20819) );
  NOR4_X1 U23742 ( .A1(n20822), .A2(n20821), .A3(n20820), .A4(n20819), .ZN(
        n20857) );
  INV_X1 U23743 ( .A(keyinput61), .ZN(n20824) );
  AOI22_X1 U23744 ( .A1(n20825), .A2(keyinput17), .B1(P1_UWORD_REG_0__SCAN_IN), 
        .B2(n20824), .ZN(n20823) );
  OAI221_X1 U23745 ( .B1(n20825), .B2(keyinput17), .C1(n20824), .C2(
        P1_UWORD_REG_0__SCAN_IN), .A(n20823), .ZN(n20838) );
  INV_X1 U23746 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n20827) );
  AOI22_X1 U23747 ( .A1(n20828), .A2(keyinput48), .B1(n20827), .B2(keyinput21), 
        .ZN(n20826) );
  OAI221_X1 U23748 ( .B1(n20828), .B2(keyinput48), .C1(n20827), .C2(keyinput21), .A(n20826), .ZN(n20837) );
  INV_X1 U23749 ( .A(keyinput55), .ZN(n20830) );
  AOI22_X1 U23750 ( .A1(n20831), .A2(keyinput15), .B1(P3_LWORD_REG_11__SCAN_IN), .B2(n20830), .ZN(n20829) );
  OAI221_X1 U23751 ( .B1(n20831), .B2(keyinput15), .C1(n20830), .C2(
        P3_LWORD_REG_11__SCAN_IN), .A(n20829), .ZN(n20836) );
  INV_X1 U23752 ( .A(keyinput42), .ZN(n20832) );
  XOR2_X1 U23753 ( .A(P1_UWORD_REG_12__SCAN_IN), .B(n20832), .Z(n20834) );
  XNOR2_X1 U23754 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B(keyinput2), .ZN(
        n20833) );
  NAND2_X1 U23755 ( .A1(n20834), .A2(n20833), .ZN(n20835) );
  NOR4_X1 U23756 ( .A1(n20838), .A2(n20837), .A3(n20836), .A4(n20835), .ZN(
        n20856) );
  INV_X1 U23757 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n20841) );
  INV_X1 U23758 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n20840) );
  AOI22_X1 U23759 ( .A1(n20841), .A2(keyinput9), .B1(keyinput49), .B2(n20840), 
        .ZN(n20839) );
  OAI221_X1 U23760 ( .B1(n20841), .B2(keyinput9), .C1(n20840), .C2(keyinput49), 
        .A(n20839), .ZN(n20854) );
  AOI22_X1 U23761 ( .A1(n20844), .A2(keyinput36), .B1(keyinput18), .B2(n20843), 
        .ZN(n20842) );
  OAI221_X1 U23762 ( .B1(n20844), .B2(keyinput36), .C1(n20843), .C2(keyinput18), .A(n20842), .ZN(n20853) );
  AOI22_X1 U23763 ( .A1(n20847), .A2(keyinput1), .B1(n20846), .B2(keyinput50), 
        .ZN(n20845) );
  OAI221_X1 U23764 ( .B1(n20847), .B2(keyinput1), .C1(n20846), .C2(keyinput50), 
        .A(n20845), .ZN(n20852) );
  INV_X1 U23765 ( .A(keyinput22), .ZN(n20849) );
  AOI22_X1 U23766 ( .A1(n20850), .A2(keyinput60), .B1(P2_LWORD_REG_0__SCAN_IN), 
        .B2(n20849), .ZN(n20848) );
  OAI221_X1 U23767 ( .B1(n20850), .B2(keyinput60), .C1(n20849), .C2(
        P2_LWORD_REG_0__SCAN_IN), .A(n20848), .ZN(n20851) );
  NOR4_X1 U23768 ( .A1(n20854), .A2(n20853), .A3(n20852), .A4(n20851), .ZN(
        n20855) );
  NAND3_X1 U23769 ( .A1(n20857), .A2(n20856), .A3(n20855), .ZN(n20922) );
  AOI22_X1 U23770 ( .A1(n20860), .A2(keyinput38), .B1(keyinput16), .B2(n20859), 
        .ZN(n20858) );
  OAI221_X1 U23771 ( .B1(n20860), .B2(keyinput38), .C1(n20859), .C2(keyinput16), .A(n20858), .ZN(n20871) );
  AOI22_X1 U23772 ( .A1(n20862), .A2(keyinput34), .B1(n14143), .B2(keyinput51), 
        .ZN(n20861) );
  OAI221_X1 U23773 ( .B1(n20862), .B2(keyinput34), .C1(n14143), .C2(keyinput51), .A(n20861), .ZN(n20870) );
  AOI22_X1 U23774 ( .A1(n20864), .A2(keyinput8), .B1(n11898), .B2(keyinput24), 
        .ZN(n20863) );
  OAI221_X1 U23775 ( .B1(n20864), .B2(keyinput8), .C1(n11898), .C2(keyinput24), 
        .A(n20863), .ZN(n20869) );
  INV_X1 U23776 ( .A(DATAI_6_), .ZN(n20866) );
  AOI22_X1 U23777 ( .A1(n20867), .A2(keyinput20), .B1(keyinput57), .B2(n20866), 
        .ZN(n20865) );
  OAI221_X1 U23778 ( .B1(n20867), .B2(keyinput20), .C1(n20866), .C2(keyinput57), .A(n20865), .ZN(n20868) );
  NOR4_X1 U23779 ( .A1(n20871), .A2(n20870), .A3(n20869), .A4(n20868), .ZN(
        n20920) );
  INV_X1 U23780 ( .A(keyinput14), .ZN(n20874) );
  INV_X1 U23781 ( .A(keyinput37), .ZN(n20873) );
  AOI22_X1 U23782 ( .A1(n20874), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n20873), .ZN(n20872) );
  OAI221_X1 U23783 ( .B1(n20874), .B2(P1_DATAO_REG_17__SCAN_IN), .C1(n20873), 
        .C2(P1_DATAO_REG_22__SCAN_IN), .A(n20872), .ZN(n20887) );
  AOI22_X1 U23784 ( .A1(n20877), .A2(keyinput23), .B1(n20876), .B2(keyinput44), 
        .ZN(n20875) );
  OAI221_X1 U23785 ( .B1(n20877), .B2(keyinput23), .C1(n20876), .C2(keyinput44), .A(n20875), .ZN(n20886) );
  INV_X1 U23786 ( .A(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n20879) );
  AOI22_X1 U23787 ( .A1(n20880), .A2(keyinput12), .B1(n20879), .B2(keyinput25), 
        .ZN(n20878) );
  OAI221_X1 U23788 ( .B1(n20880), .B2(keyinput12), .C1(n20879), .C2(keyinput25), .A(n20878), .ZN(n20885) );
  INV_X1 U23789 ( .A(keyinput10), .ZN(n20881) );
  XOR2_X1 U23790 ( .A(P1_DATAWIDTH_REG_15__SCAN_IN), .B(n20881), .Z(n20883) );
  XNOR2_X1 U23791 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B(keyinput32), .ZN(
        n20882) );
  NAND2_X1 U23792 ( .A1(n20883), .A2(n20882), .ZN(n20884) );
  NOR4_X1 U23793 ( .A1(n20887), .A2(n20886), .A3(n20885), .A4(n20884), .ZN(
        n20919) );
  INV_X1 U23794 ( .A(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n20889) );
  AOI22_X1 U23795 ( .A1(n20890), .A2(keyinput62), .B1(n20889), .B2(keyinput59), 
        .ZN(n20888) );
  OAI221_X1 U23796 ( .B1(n20890), .B2(keyinput62), .C1(n20889), .C2(keyinput59), .A(n20888), .ZN(n20903) );
  INV_X1 U23797 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n20893) );
  AOI22_X1 U23798 ( .A1(n20893), .A2(keyinput26), .B1(n20892), .B2(keyinput53), 
        .ZN(n20891) );
  OAI221_X1 U23799 ( .B1(n20893), .B2(keyinput26), .C1(n20892), .C2(keyinput53), .A(n20891), .ZN(n20902) );
  INV_X1 U23800 ( .A(keyinput63), .ZN(n20896) );
  AOI22_X1 U23801 ( .A1(n20896), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(keyinput27), 
        .B2(n20895), .ZN(n20894) );
  OAI221_X1 U23802 ( .B1(n20896), .B2(P3_UWORD_REG_8__SCAN_IN), .C1(n20895), 
        .C2(keyinput27), .A(n20894), .ZN(n20901) );
  AOI22_X1 U23803 ( .A1(n20899), .A2(keyinput30), .B1(keyinput5), .B2(n9743), 
        .ZN(n20897) );
  OAI221_X1 U23804 ( .B1(n20899), .B2(keyinput30), .C1(n20898), .C2(keyinput5), 
        .A(n20897), .ZN(n20900) );
  NOR4_X1 U23805 ( .A1(n20903), .A2(n20902), .A3(n20901), .A4(n20900), .ZN(
        n20918) );
  INV_X1 U23806 ( .A(keyinput39), .ZN(n20905) );
  AOI22_X1 U23807 ( .A1(n15128), .A2(keyinput13), .B1(P3_DATAO_REG_9__SCAN_IN), 
        .B2(n20905), .ZN(n20904) );
  OAI221_X1 U23808 ( .B1(n15128), .B2(keyinput13), .C1(n20905), .C2(
        P3_DATAO_REG_9__SCAN_IN), .A(n20904), .ZN(n20916) );
  INV_X1 U23809 ( .A(keyinput33), .ZN(n20907) );
  AOI22_X1 U23810 ( .A1(n20908), .A2(keyinput3), .B1(P3_DATAO_REG_19__SCAN_IN), 
        .B2(n20907), .ZN(n20906) );
  OAI221_X1 U23811 ( .B1(n20908), .B2(keyinput3), .C1(n20907), .C2(
        P3_DATAO_REG_19__SCAN_IN), .A(n20906), .ZN(n20915) );
  AOI22_X1 U23812 ( .A1(n15130), .A2(keyinput11), .B1(n11967), .B2(keyinput4), 
        .ZN(n20909) );
  OAI221_X1 U23813 ( .B1(n15130), .B2(keyinput11), .C1(n11967), .C2(keyinput4), 
        .A(n20909), .ZN(n20914) );
  AOI22_X1 U23814 ( .A1(n20912), .A2(keyinput35), .B1(n20911), .B2(keyinput41), 
        .ZN(n20910) );
  OAI221_X1 U23815 ( .B1(n20912), .B2(keyinput35), .C1(n20911), .C2(keyinput41), .A(n20910), .ZN(n20913) );
  NOR4_X1 U23816 ( .A1(n20916), .A2(n20915), .A3(n20914), .A4(n20913), .ZN(
        n20917) );
  NAND4_X1 U23817 ( .A1(n20920), .A2(n20919), .A3(n20918), .A4(n20917), .ZN(
        n20921) );
  NOR4_X1 U23818 ( .A1(n20924), .A2(n20923), .A3(n20922), .A4(n20921), .ZN(
        n20934) );
  AOI21_X1 U23819 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n20926), .A(n20925), .ZN(
        n20929) );
  OAI222_X1 U23820 ( .A1(n20932), .A2(n20931), .B1(n20930), .B2(n20929), .C1(
        n20928), .C2(n20927), .ZN(n20933) );
  XOR2_X1 U23821 ( .A(n20934), .B(n20933), .Z(P3_U2729) );
  AND4_X1 U12969 ( .A1(n10140), .A2(n10139), .A3(n10138), .A4(n10137), .ZN(
        n10171) );
  BUF_X2 U12404 ( .A(n11756), .Z(n14787) );
  AND4_X2 U11089 ( .A1(n10174), .A2(n10173), .A3(n10172), .A4(n10171), .ZN(
        n12635) );
  CLKBUF_X1 U11095 ( .A(n10761), .Z(n17050) );
  CLKBUF_X1 U11130 ( .A(n14072), .Z(n14073) );
  INV_X2 U11131 ( .A(n10510), .ZN(n15980) );
  CLKBUF_X1 U11132 ( .A(n11851), .Z(n14020) );
  CLKBUF_X1 U11865 ( .A(n13215), .Z(n13188) );
  CLKBUF_X1 U11883 ( .A(n11766), .Z(n13344) );
  CLKBUF_X1 U12107 ( .A(n14095), .Z(n14109) );
  CLKBUF_X1 U12171 ( .A(n19114), .Z(n19111) );
  CLKBUF_X1 U12194 ( .A(n10815), .Z(n17300) );
  CLKBUF_X1 U12198 ( .A(n16447), .Z(n16445) );
  CLKBUF_X1 U12226 ( .A(n18747), .Z(n17340) );
endmodule

