

module b20_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852;

  INV_X4 U5014 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NAND2_X1 U5015 ( .A1(n9321), .A2(n9305), .ZN(n9357) );
  AND2_X1 U5016 ( .A1(n6777), .A2(n6776), .ZN(n10439) );
  OAI21_X1 U5017 ( .B1(n6780), .B2(n6779), .A(n6778), .ZN(n6784) );
  NAND2_X1 U5018 ( .A1(n6771), .A2(n6770), .ZN(n6780) );
  OAI21_X1 U5019 ( .B1(n9562), .B2(n9141), .A(n9259), .ZN(n9552) );
  OR2_X1 U5020 ( .A1(n8515), .A2(n8516), .ZN(n8635) );
  CLKBUF_X2 U5021 ( .A(n10211), .Z(n4961) );
  XNOR2_X1 U5022 ( .A(n6009), .B(n6008), .ZN(n6007) );
  INV_X1 U5023 ( .A(n7150), .ZN(n7179) );
  INV_X2 U5024 ( .A(n7028), .ZN(n7150) );
  INV_X1 U5025 ( .A(n7625), .ZN(n9393) );
  AND4_X1 U5026 ( .A1(n6235), .A2(n6234), .A3(n6233), .A4(n6232), .ZN(n7625)
         );
  NAND2_X1 U5027 ( .A1(n7316), .A2(n4965), .ZN(n5659) );
  BUF_X2 U5028 ( .A(n5617), .Z(n4965) );
  CLKBUF_X2 U5029 ( .A(n5617), .Z(n4964) );
  NOR2_X1 U5030 ( .A1(n6214), .A2(n6197), .ZN(n5221) );
  NOR2_X1 U5031 ( .A1(n6260), .A2(n6213), .ZN(n5220) );
  NAND2_X2 U5032 ( .A1(n5071), .A2(n5460), .ZN(n5617) );
  CLKBUF_X1 U5033 ( .A(n10852), .Z(P1_U3973) );
  AND2_X1 U5034 ( .A1(n7255), .A2(n7319), .ZN(n10852) );
  NAND2_X1 U5035 ( .A1(n9588), .A2(n4955), .ZN(n4952) );
  AND2_X2 U5036 ( .A1(n4952), .A2(n4953), .ZN(n9562) );
  OR2_X1 U5037 ( .A1(n4954), .A2(n5360), .ZN(n4953) );
  INV_X1 U5038 ( .A(n9247), .ZN(n4954) );
  AND2_X1 U5039 ( .A1(n9572), .A2(n9247), .ZN(n4955) );
  AND3_X2 U5041 ( .A1(n5107), .A2(n5028), .A3(n5106), .ZN(n4957) );
  INV_X4 U5042 ( .A(n10328), .ZN(n10335) );
  BUF_X1 U5043 ( .A(n6970), .Z(n7176) );
  OR2_X1 U5044 ( .A1(n10211), .A2(n10360), .ZN(n10185) );
  CLKBUF_X2 U5045 ( .A(n7269), .Z(n7270) );
  INV_X1 U5047 ( .A(n6599), .ZN(n6457) );
  NAND2_X1 U5048 ( .A1(n10185), .A2(n6745), .ZN(n10201) );
  INV_X2 U5049 ( .A(n5659), .ZN(n6785) );
  XNOR2_X1 U5050 ( .A(n6219), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9464) );
  NAND2_X1 U5051 ( .A1(n5652), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5598) );
  XNOR2_X1 U5052 ( .A(n5591), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5597) );
  XNOR2_X1 U5053 ( .A(n6218), .B(n6217), .ZN(n6221) );
  OAI21_X2 U5054 ( .B1(n5847), .B2(n5480), .A(n5477), .ZN(n5903) );
  NAND2_X2 U5055 ( .A1(n5845), .A2(n5844), .ZN(n5847) );
  XNOR2_X2 U5056 ( .A(n8076), .B(n10044), .ZN(n6119) );
  AOI211_X2 U5057 ( .C1(n9257), .C2(n9565), .A(n9264), .B(n9555), .ZN(n5298)
         );
  BUF_X4 U5058 ( .A(n5631), .Z(n4958) );
  AND2_X1 U5059 ( .A1(n5597), .A2(n10481), .ZN(n5631) );
  NAND2_X2 U5060 ( .A1(n6117), .A2(n8218), .ZN(n6950) );
  NAND2_X1 U5061 ( .A1(n7264), .A2(n7263), .ZN(n4959) );
  NAND2_X1 U5062 ( .A1(n7264), .A2(n7263), .ZN(n4960) );
  NAND2_X1 U5063 ( .A1(n7264), .A2(n7263), .ZN(n7269) );
  INV_X2 U5064 ( .A(n7269), .ZN(n8966) );
  NAND2_X2 U5065 ( .A1(n6012), .A2(n6011), .ZN(n10234) );
  NAND2_X1 U5066 ( .A1(n7709), .A2(n5540), .ZN(n7795) );
  OAI21_X1 U5067 ( .B1(n6512), .B2(n5659), .A(n6050), .ZN(n10211) );
  OAI21_X2 U5068 ( .B1(n6007), .B2(SI_22_), .A(n6010), .ZN(n6022) );
  NOR4_X2 U5069 ( .A1(n9355), .A2(n9354), .A3(n9353), .A4(n9352), .ZN(n9361)
         );
  OAI21_X1 U5070 ( .B1(n6766), .B2(n10143), .A(n6765), .ZN(n6794) );
  OAI21_X1 U5071 ( .B1(n5078), .B2(n5076), .A(n5073), .ZN(n10202) );
  OR3_X1 U5072 ( .A1(n10201), .A2(n6843), .A3(n6802), .ZN(n6659) );
  AOI21_X1 U5073 ( .B1(n6736), .B2(n6802), .A(n10256), .ZN(n5274) );
  AND2_X1 U5074 ( .A1(n8634), .A2(n4983), .ZN(n10322) );
  AND2_X1 U5075 ( .A1(n8398), .A2(n8437), .ZN(n8474) );
  OR2_X1 U5076 ( .A1(n7855), .A2(n7856), .ZN(n7857) );
  OR2_X1 U5077 ( .A1(n8289), .A2(n8288), .ZN(n8270) );
  OAI21_X1 U5078 ( .B1(n7397), .B2(n5659), .A(n5776), .ZN(n8269) );
  INV_X1 U5079 ( .A(n8347), .ZN(n7848) );
  NAND2_X2 U5080 ( .A1(n6674), .A2(n6876), .ZN(n8128) );
  INV_X4 U5082 ( .A(n9269), .ZN(n9284) );
  NAND2_X1 U5083 ( .A1(n6945), .A2(n8088), .ZN(n6876) );
  NAND2_X1 U5084 ( .A1(n8078), .A2(n6813), .ZN(n6121) );
  INV_X1 U5085 ( .A(n9392), .ZN(n6284) );
  INV_X1 U5086 ( .A(n6802), .ZN(n4963) );
  INV_X1 U5087 ( .A(n8088), .ZN(n10043) );
  INV_X2 U5088 ( .A(n6145), .ZN(n5609) );
  XNOR2_X1 U5090 ( .A(n5534), .B(P2_IR_REG_30__SCAN_IN), .ZN(n9838) );
  NAND2_X1 U5091 ( .A1(n6113), .A2(n6112), .ZN(n6114) );
  NOR2_X1 U5092 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n6208) );
  AOI21_X1 U5093 ( .B1(n8916), .B2(n10842), .A(n5247), .ZN(n8918) );
  OAI21_X1 U5094 ( .B1(n8916), .B2(n10843), .A(n5185), .ZN(n6194) );
  INV_X1 U5095 ( .A(n7186), .ZN(n7213) );
  AOI21_X1 U5096 ( .B1(n5188), .B2(n10838), .A(n6153), .ZN(n5187) );
  NAND2_X1 U5097 ( .A1(n5105), .A2(n5005), .ZN(n7186) );
  OR3_X1 U5098 ( .A1(n9715), .A2(n9714), .A3(n9713), .ZN(n9797) );
  OAI21_X1 U5099 ( .B1(n10353), .B2(n10425), .A(n5085), .ZN(n5084) );
  AND2_X1 U5100 ( .A1(n10350), .A2(n10349), .ZN(n10351) );
  XNOR2_X1 U5101 ( .A(n5087), .B(n10168), .ZN(n10353) );
  OAI21_X1 U5102 ( .B1(n5183), .B2(n8902), .A(n5181), .ZN(n10165) );
  AOI22_X1 U5103 ( .A1(n10140), .A2(n10312), .B1(n10139), .B2(n10138), .ZN(
        n10350) );
  OR2_X1 U5104 ( .A1(n6852), .A2(n10127), .ZN(n6930) );
  NAND2_X1 U5105 ( .A1(n9552), .A2(n6587), .ZN(n5309) );
  OR2_X1 U5106 ( .A1(n10439), .A2(n10138), .ZN(n6808) );
  NAND2_X1 U5107 ( .A1(n10186), .A2(n5378), .ZN(n10169) );
  OR2_X1 U5108 ( .A1(n6152), .A2(n10147), .ZN(n10156) );
  NAND2_X1 U5109 ( .A1(n6789), .A2(n6788), .ZN(n6852) );
  AND2_X1 U5110 ( .A1(n8980), .A2(n8977), .ZN(n5542) );
  OAI21_X1 U5111 ( .B1(n6524), .B2(n5385), .A(n5383), .ZN(n7221) );
  NAND2_X1 U5112 ( .A1(n10184), .A2(n5168), .ZN(n10186) );
  NAND2_X1 U5113 ( .A1(n5158), .A2(n5524), .ZN(n8967) );
  NAND2_X1 U5114 ( .A1(n10203), .A2(n10204), .ZN(n10184) );
  NAND2_X1 U5115 ( .A1(n10269), .A2(n5967), .ZN(n10257) );
  NAND2_X1 U5116 ( .A1(n8921), .A2(n6135), .ZN(n10203) );
  OAI21_X1 U5117 ( .B1(n5335), .B2(n5334), .A(n7231), .ZN(n5333) );
  NAND2_X1 U5118 ( .A1(n7224), .A2(n7223), .ZN(n7243) );
  OAI21_X1 U5119 ( .B1(n5272), .B2(n6828), .A(n5271), .ZN(n6742) );
  XNOR2_X1 U5120 ( .A(n6780), .B(n6779), .ZN(n9289) );
  AOI21_X1 U5121 ( .B1(n5275), .B2(n5274), .A(n5273), .ZN(n5272) );
  AND2_X1 U5122 ( .A1(n6590), .A2(n8978), .ZN(n5335) );
  AND2_X1 U5123 ( .A1(n9312), .A2(n9314), .ZN(n9351) );
  NAND2_X1 U5124 ( .A1(n10220), .A2(n10221), .ZN(n10219) );
  NAND2_X1 U5125 ( .A1(n10289), .A2(n5952), .ZN(n10288) );
  AND2_X1 U5126 ( .A1(n6834), .A2(n6746), .ZN(n10190) );
  NAND2_X1 U5127 ( .A1(n5242), .A2(n6149), .ZN(n5241) );
  AND2_X1 U5128 ( .A1(n10171), .A2(n6746), .ZN(n5378) );
  OR2_X1 U5129 ( .A1(n9282), .A2(n9499), .ZN(n9312) );
  OR2_X1 U5130 ( .A1(n6767), .A2(n8763), .ZN(n6771) );
  AND2_X1 U5131 ( .A1(n6835), .A2(n6833), .ZN(n10171) );
  AOI21_X1 U5132 ( .B1(n5079), .B2(n5075), .A(n5074), .ZN(n5073) );
  INV_X1 U5133 ( .A(n9515), .ZN(n9703) );
  NAND2_X1 U5134 ( .A1(n6544), .A2(n6543), .ZN(n9282) );
  AND2_X1 U5135 ( .A1(n9308), .A2(n5003), .ZN(n9494) );
  OR2_X1 U5136 ( .A1(n10177), .A2(n7203), .ZN(n6835) );
  INV_X1 U5137 ( .A(n10177), .ZN(n6149) );
  AND2_X1 U5138 ( .A1(n6526), .A2(n6525), .ZN(n9515) );
  OR2_X1 U5139 ( .A1(n8992), .A2(n9122), .ZN(n9308) );
  AND2_X1 U5140 ( .A1(n6135), .A2(n6841), .ZN(n8922) );
  NAND2_X1 U5141 ( .A1(n6515), .A2(n6514), .ZN(n9518) );
  NOR2_X1 U5142 ( .A1(n9547), .A2(n9262), .ZN(n5197) );
  NAND2_X1 U5143 ( .A1(n6536), .A2(n6535), .ZN(n8992) );
  OR2_X1 U5144 ( .A1(n6512), .A2(n6513), .ZN(n6515) );
  OR2_X2 U5145 ( .A1(n9263), .A2(n9262), .ZN(n9555) );
  NAND2_X1 U5146 ( .A1(n6082), .A2(n6081), .ZN(n10177) );
  NAND2_X1 U5147 ( .A1(n5083), .A2(n5082), .ZN(n8643) );
  NAND2_X1 U5148 ( .A1(n5530), .A2(n5006), .ZN(n9048) );
  AND2_X1 U5149 ( .A1(n5204), .A2(n5359), .ZN(n5203) );
  NAND2_X1 U5150 ( .A1(n6028), .A2(n6027), .ZN(n10372) );
  NOR2_X1 U5151 ( .A1(n9084), .A2(n5528), .ZN(n5527) );
  AOI21_X1 U5152 ( .B1(n5362), .B2(n5365), .A(n5360), .ZN(n5359) );
  OR2_X1 U5153 ( .A1(n9142), .A2(n9141), .ZN(n9565) );
  NAND2_X1 U5154 ( .A1(n6504), .A2(n6503), .ZN(n9531) );
  NAND2_X1 U5155 ( .A1(n5362), .A2(n5205), .ZN(n5204) );
  NAND2_X1 U5156 ( .A1(n8592), .A2(n8591), .ZN(n8938) );
  AND2_X1 U5157 ( .A1(n6915), .A2(n6737), .ZN(n10252) );
  NAND2_X1 U5158 ( .A1(n9639), .A2(n9638), .ZN(n9637) );
  AND2_X2 U5159 ( .A1(n6496), .A2(n6495), .ZN(n9801) );
  NAND2_X1 U5160 ( .A1(n5995), .A2(n5994), .ZN(n10383) );
  NAND2_X1 U5161 ( .A1(n6484), .A2(n6483), .ZN(n9258) );
  OR2_X1 U5162 ( .A1(n10390), .A2(n7120), .ZN(n6915) );
  INV_X1 U5163 ( .A(n5151), .ZN(n8592) );
  OR2_X1 U5164 ( .A1(n9577), .A2(n9376), .ZN(n9247) );
  AND2_X1 U5165 ( .A1(n5162), .A2(n5389), .ZN(n5161) );
  OAI21_X1 U5166 ( .B1(n8629), .B2(n8628), .A(n6898), .ZN(n8614) );
  NAND2_X1 U5167 ( .A1(n5981), .A2(n5980), .ZN(n10390) );
  INV_X1 U5168 ( .A(n9328), .ZN(n5366) );
  AOI21_X1 U5169 ( .B1(n5122), .B2(n5120), .A(n5119), .ZN(n5118) );
  NAND2_X1 U5170 ( .A1(n6476), .A2(n6475), .ZN(n9577) );
  NAND2_X1 U5171 ( .A1(n8575), .A2(n5154), .ZN(n9091) );
  NAND2_X1 U5172 ( .A1(n8285), .A2(n5761), .ZN(n8268) );
  OR2_X1 U5173 ( .A1(n9594), .A2(n9603), .ZN(n9248) );
  NOR2_X1 U5174 ( .A1(n8908), .A2(n5237), .ZN(n5236) );
  AND2_X1 U5175 ( .A1(n6728), .A2(n6910), .ZN(n10300) );
  OR2_X1 U5176 ( .A1(n9014), .A2(n9378), .ZN(n8956) );
  AND2_X1 U5177 ( .A1(n6902), .A2(n6709), .ZN(n8617) );
  AND2_X1 U5178 ( .A1(n9237), .A2(n9232), .ZN(n9615) );
  NAND2_X1 U5179 ( .A1(n5959), .A2(n5958), .ZN(n10273) );
  NAND2_X1 U5180 ( .A1(n6467), .A2(n6466), .ZN(n9594) );
  NAND2_X1 U5181 ( .A1(n5944), .A2(n5943), .ZN(n10296) );
  NOR2_X1 U5182 ( .A1(n10024), .A2(n10422), .ZN(n5238) );
  INV_X1 U5183 ( .A(n6902), .ZN(n5167) );
  OAI21_X1 U5184 ( .B1(n4990), .B2(n5141), .A(n9000), .ZN(n5140) );
  OR2_X1 U5185 ( .A1(n9106), .A2(n9623), .ZN(n9237) );
  AOI22_X1 U5186 ( .A1(n5404), .A2(n5401), .B1(n5408), .B2(n5400), .ZN(n5399)
         );
  NAND2_X1 U5187 ( .A1(n6459), .A2(n6458), .ZN(n9014) );
  NAND2_X1 U5188 ( .A1(n6448), .A2(n6447), .ZN(n9106) );
  AND2_X1 U5189 ( .A1(n9226), .A2(n9225), .ZN(n9638) );
  AND2_X1 U5190 ( .A1(n6408), .A2(n6407), .ZN(n9834) );
  AND2_X1 U5191 ( .A1(n9206), .A2(n9207), .ZN(n9344) );
  AND2_X1 U5192 ( .A1(n9216), .A2(n6402), .ZN(n9664) );
  OAI21_X1 U5193 ( .B1(n8309), .B2(n5452), .A(n5451), .ZN(n10634) );
  AND2_X1 U5194 ( .A1(n5407), .A2(n8378), .ZN(n5406) );
  NAND2_X1 U5195 ( .A1(n6435), .A2(n6434), .ZN(n9234) );
  OAI21_X1 U5196 ( .B1(n5935), .B2(n5476), .A(n5937), .ZN(n5957) );
  OR2_X1 U5197 ( .A1(n10427), .A2(n10021), .ZN(n6898) );
  OR2_X1 U5198 ( .A1(n8941), .A2(n9383), .ZN(n5552) );
  AND2_X1 U5199 ( .A1(n5818), .A2(n5817), .ZN(n10836) );
  NAND2_X1 U5200 ( .A1(n6396), .A2(n6395), .ZN(n9757) );
  NAND2_X1 U5201 ( .A1(n5891), .A2(n5890), .ZN(n10422) );
  NAND2_X1 U5202 ( .A1(n5852), .A2(n5851), .ZN(n10427) );
  NOR2_X2 U5203 ( .A1(n8270), .A2(n8269), .ZN(n8398) );
  NOR2_X1 U5204 ( .A1(n4989), .A2(n5327), .ZN(n5326) );
  NAND2_X1 U5205 ( .A1(n6384), .A2(n6383), .ZN(n9677) );
  NAND2_X1 U5206 ( .A1(n5791), .A2(n5790), .ZN(n8572) );
  NAND2_X1 U5207 ( .A1(n5833), .A2(n5832), .ZN(n8516) );
  AND2_X1 U5208 ( .A1(n8111), .A2(n8370), .ZN(n8251) );
  AND2_X1 U5209 ( .A1(n6884), .A2(n8224), .ZN(n8102) );
  NOR2_X1 U5210 ( .A1(n8125), .A2(n5243), .ZN(n8111) );
  AND2_X1 U5211 ( .A1(n6691), .A2(n8226), .ZN(n8225) );
  OR2_X1 U5212 ( .A1(n8426), .A2(n8577), .ZN(n9194) );
  NAND2_X1 U5213 ( .A1(n5175), .A2(n5753), .ZN(n8288) );
  AND2_X1 U5214 ( .A1(n6334), .A2(n6333), .ZN(n8193) );
  INV_X2 U5215 ( .A(n9672), .ZN(n9694) );
  NAND2_X1 U5216 ( .A1(n5770), .A2(n5769), .ZN(n5786) );
  AND2_X1 U5217 ( .A1(n5722), .A2(n5721), .ZN(n8370) );
  XNOR2_X1 U5218 ( .A(n5765), .B(n5764), .ZN(n7398) );
  NAND2_X2 U5219 ( .A1(n7647), .A2(n9669), .ZN(n9672) );
  OAI21_X1 U5220 ( .B1(n7375), .B2(n6513), .A(n6327), .ZN(n8180) );
  NAND2_X1 U5221 ( .A1(n7301), .A2(n9284), .ZN(n9685) );
  OAI211_X1 U5222 ( .C1(n6513), .C2(n7371), .A(n6306), .B(n6305), .ZN(n7915)
         );
  NAND2_X1 U5223 ( .A1(n5717), .A2(n5716), .ZN(n5733) );
  AND2_X1 U5224 ( .A1(n6956), .A2(n6955), .ZN(n6964) );
  NAND2_X1 U5225 ( .A1(n6121), .A2(n6120), .ZN(n8127) );
  AND3_X1 U5226 ( .A1(n5669), .A2(n5668), .A3(n5667), .ZN(n10784) );
  NAND3_X1 U5227 ( .A1(n5112), .A2(n5711), .A3(n5111), .ZN(n5717) );
  INV_X1 U5228 ( .A(n7895), .ZN(n6283) );
  NAND2_X1 U5229 ( .A1(n5700), .A2(n5089), .ZN(n7371) );
  AND3_X1 U5230 ( .A1(n6282), .A2(n6281), .A3(n6280), .ZN(n7895) );
  INV_X2 U5231 ( .A(n7380), .ZN(n7400) );
  INV_X2 U5233 ( .A(n6970), .ZN(n7163) );
  AND4_X1 U5234 ( .A1(n6291), .A2(n6290), .A3(n6289), .A4(n6288), .ZN(n7908)
         );
  AND2_X1 U5235 ( .A1(n6246), .A2(n5192), .ZN(n7265) );
  AND4_X1 U5236 ( .A1(n5613), .A2(n5612), .A3(n5611), .A4(n5610), .ZN(n8088)
         );
  AND2_X1 U5237 ( .A1(n8019), .A2(n6949), .ZN(n7001) );
  NAND2_X1 U5238 ( .A1(n6947), .A2(n10116), .ZN(n8014) );
  XNOR2_X1 U5239 ( .A(n6172), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6947) );
  INV_X1 U5240 ( .A(n6115), .ZN(n10116) );
  OAI21_X1 U5241 ( .B1(n6204), .B2(P2_IR_REG_19__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6218) );
  AND2_X2 U5242 ( .A1(n6252), .A2(n7346), .ZN(n6275) );
  NAND2_X1 U5243 ( .A1(n5395), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6172) );
  AOI21_X1 U5244 ( .B1(n5559), .B2(n5456), .A(n5455), .ZN(n5454) );
  NAND2_X1 U5246 ( .A1(n5597), .A2(n5596), .ZN(n6145) );
  OAI21_X1 U5247 ( .B1(n5684), .B2(n5115), .A(n5704), .ZN(n5114) );
  INV_X1 U5248 ( .A(n5596), .ZN(n10481) );
  AND2_X1 U5249 ( .A1(n5595), .A2(n10475), .ZN(n5596) );
  XNOR2_X1 U5250 ( .A(n6166), .B(n5388), .ZN(n10490) );
  AND2_X1 U5251 ( .A1(n5660), .A2(n5645), .ZN(n5646) );
  NAND2_X2 U5252 ( .A1(n5354), .A2(n5351), .ZN(n6601) );
  NAND2_X1 U5253 ( .A1(n7316), .A2(n7346), .ZN(n6787) );
  NAND2_X1 U5254 ( .A1(n6614), .A2(n4969), .ZN(n8610) );
  OAI21_X2 U5255 ( .B1(n6114), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6162) );
  XNOR2_X1 U5256 ( .A(n6114), .B(P1_IR_REG_20__SCAN_IN), .ZN(n8218) );
  OR2_X1 U5257 ( .A1(n5594), .A2(n10474), .ZN(n5591) );
  NAND2_X1 U5258 ( .A1(n5576), .A2(n5575), .ZN(n7316) );
  MUX2_X1 U5259 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6613), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n6614) );
  NAND2_X1 U5260 ( .A1(n6229), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5534) );
  AND2_X1 U5261 ( .A1(n5070), .A2(SI_0_), .ZN(n5585) );
  NOR2_X1 U5262 ( .A1(n5353), .A2(n5352), .ZN(n5351) );
  AND2_X1 U5263 ( .A1(n5522), .A2(n5719), .ZN(n6154) );
  NAND2_X1 U5264 ( .A1(n5428), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6113) );
  NAND2_X1 U5265 ( .A1(n5155), .A2(n6612), .ZN(n6639) );
  AND2_X1 U5266 ( .A1(n5523), .A2(n4972), .ZN(n5522) );
  OR2_X1 U5267 ( .A1(n6197), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5544) );
  AND3_X1 U5268 ( .A1(n6116), .A2(n6171), .A3(n6174), .ZN(n6159) );
  AND2_X1 U5269 ( .A1(n5323), .A2(n6222), .ZN(n5318) );
  NAND2_X1 U5270 ( .A1(n6198), .A2(n5292), .ZN(n5291) );
  NAND3_X1 U5271 ( .A1(n10776), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5460) );
  NOR2_X1 U5272 ( .A1(P1_RD_REG_SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n5579) );
  INV_X1 U5273 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6324) );
  NOR2_X1 U5274 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5339) );
  INV_X1 U5275 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6404) );
  NOR2_X1 U5276 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n6196) );
  INV_X1 U5277 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6313) );
  INV_X1 U5278 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6302) );
  NOR2_X1 U5279 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n6110) );
  XNOR2_X1 U5280 ( .A(n6784), .B(n6783), .ZN(n9835) );
  XNOR2_X1 U5281 ( .A(n6090), .B(n6089), .ZN(n10486) );
  AND2_X4 U5282 ( .A1(n9842), .A2(n6230), .ZN(n6267) );
  NAND2_X4 U5283 ( .A1(n6959), .A2(n6970), .ZN(n6966) );
  AOI21_X1 U5284 ( .B1(n9841), .B2(n6785), .A(n6763), .ZN(n10152) );
  NAND2_X1 U5285 ( .A1(n5354), .A2(n5351), .ZN(n4967) );
  NAND2_X2 U5286 ( .A1(n6600), .A2(n4967), .ZN(n6252) );
  NAND2_X1 U5287 ( .A1(n5266), .A2(n5265), .ZN(n6706) );
  NAND2_X1 U5288 ( .A1(n10634), .A2(n5058), .ZN(n5056) );
  OR2_X1 U5289 ( .A1(n10634), .A2(n5041), .ZN(n5053) );
  NAND2_X1 U5290 ( .A1(n8188), .A2(n8189), .ZN(n6567) );
  NOR2_X1 U5291 ( .A1(n5382), .A2(n9624), .ZN(n5381) );
  INV_X1 U5292 ( .A(n9225), .ZN(n5382) );
  AND2_X1 U5293 ( .A1(n6231), .A2(n9838), .ZN(n6269) );
  NAND2_X1 U5294 ( .A1(n6236), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6238) );
  NAND2_X1 U5295 ( .A1(n5262), .A2(n4992), .ZN(n5261) );
  NAND2_X1 U5296 ( .A1(n5264), .A2(n5263), .ZN(n5262) );
  NAND2_X1 U5297 ( .A1(n6721), .A2(n6897), .ZN(n5264) );
  AOI21_X1 U5298 ( .B1(n6584), .B2(n6585), .A(n5123), .ZN(n5122) );
  INV_X1 U5299 ( .A(n8955), .ZN(n5123) );
  NAND2_X1 U5300 ( .A1(n7630), .A2(n9393), .ZN(n9150) );
  NOR2_X1 U5301 ( .A1(n5526), .A2(n5160), .ZN(n5159) );
  INV_X1 U5302 ( .A(n8961), .ZN(n5160) );
  INV_X1 U5303 ( .A(n5527), .ZN(n5526) );
  INV_X1 U5304 ( .A(n5140), .ZN(n5139) );
  INV_X1 U5305 ( .A(n9838), .ZN(n6230) );
  NAND2_X1 U5306 ( .A1(n7584), .A2(n7583), .ZN(n7679) );
  NAND2_X1 U5307 ( .A1(n7569), .A2(n5439), .ZN(n7574) );
  NAND2_X1 U5308 ( .A1(n5441), .A2(n5440), .ZN(n5439) );
  NAND2_X1 U5309 ( .A1(n10572), .A2(n7573), .ZN(n7575) );
  AND2_X1 U5310 ( .A1(n5441), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5438) );
  NAND2_X1 U5311 ( .A1(n5065), .A2(n7652), .ZN(n5064) );
  NOR2_X1 U5312 ( .A1(n5289), .A2(n6260), .ZN(n5287) );
  NAND2_X1 U5313 ( .A1(n5290), .A2(n6207), .ZN(n5289) );
  NAND2_X1 U5314 ( .A1(n5052), .A2(n5040), .ZN(n5051) );
  INV_X1 U5315 ( .A(n5448), .ZN(n5050) );
  INV_X1 U5316 ( .A(n6574), .ZN(n5307) );
  AOI21_X1 U5317 ( .B1(n5212), .B2(n5216), .A(n5210), .ZN(n5209) );
  INV_X1 U5318 ( .A(n9194), .ZN(n5210) );
  XNOR2_X1 U5319 ( .A(n8610), .B(P2_B_REG_SCAN_IN), .ZN(n5157) );
  NOR2_X1 U5320 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n5549) );
  INV_X1 U5321 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6222) );
  NAND2_X1 U5322 ( .A1(n5325), .A2(n5324), .ZN(n6611) );
  INV_X1 U5323 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5325) );
  INV_X1 U5324 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5324) );
  AND2_X1 U5325 ( .A1(n5405), .A2(n8488), .ZN(n5404) );
  NAND2_X1 U5326 ( .A1(n5406), .A2(n8377), .ZN(n5405) );
  AND2_X1 U5327 ( .A1(n5409), .A2(n8489), .ZN(n5408) );
  NAND2_X1 U5328 ( .A1(n8377), .A2(n8378), .ZN(n5409) );
  NOR2_X1 U5329 ( .A1(n6128), .A2(n5174), .ZN(n5173) );
  INV_X1 U5330 ( .A(n6729), .ZN(n5174) );
  AND2_X1 U5331 ( .A1(n10273), .A2(n10302), .ZN(n6129) );
  INV_X1 U5332 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5429) );
  XNOR2_X1 U5333 ( .A(n8966), .B(n7880), .ZN(n7273) );
  AOI21_X1 U5334 ( .B1(n4987), .B2(n8051), .A(n4979), .ZN(n5546) );
  OR2_X1 U5335 ( .A1(n8576), .A2(n8577), .ZN(n5154) );
  INV_X1 U5336 ( .A(n7620), .ZN(n5537) );
  INV_X1 U5337 ( .A(n5384), .ZN(n5383) );
  OAI21_X1 U5338 ( .B1(n4970), .B2(n5385), .A(n9308), .ZN(n5384) );
  NAND2_X1 U5339 ( .A1(n9508), .A2(n5003), .ZN(n5385) );
  INV_X1 U5340 ( .A(n5367), .ZN(n5364) );
  NAND2_X1 U5341 ( .A1(n5366), .A2(n9241), .ZN(n5365) );
  NOR2_X1 U5342 ( .A1(n5368), .A2(n9243), .ZN(n5367) );
  INV_X1 U5343 ( .A(n9237), .ZN(n5368) );
  NAND2_X1 U5344 ( .A1(n5227), .A2(n5225), .ZN(n9639) );
  AOI21_X1 U5345 ( .B1(n5228), .B2(n9664), .A(n5226), .ZN(n5225) );
  INV_X1 U5346 ( .A(n6416), .ZN(n5226) );
  NAND2_X1 U5347 ( .A1(n8481), .A2(n9200), .ZN(n8528) );
  NAND2_X1 U5348 ( .A1(n6563), .A2(n6562), .ZN(n8068) );
  NOR2_X1 U5349 ( .A1(n4980), .A2(n5315), .ZN(n5310) );
  NAND2_X1 U5350 ( .A1(n6275), .A2(n5357), .ZN(n5356) );
  INV_X1 U5351 ( .A(n7373), .ZN(n5357) );
  INV_X1 U5352 ( .A(n6275), .ZN(n6513) );
  MUX2_X1 U5353 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6225), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n6228) );
  INV_X1 U5354 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6174) );
  INV_X1 U5355 ( .A(n7212), .ZN(n5413) );
  AND2_X1 U5356 ( .A1(n5399), .A2(n7030), .ZN(n5103) );
  OR2_X1 U5357 ( .A1(n6099), .A2(n6098), .ZN(n10149) );
  INV_X1 U5358 ( .A(n10135), .ZN(n5375) );
  NOR3_X2 U5359 ( .A1(n10195), .A2(n5241), .A3(n10157), .ZN(n10147) );
  AND2_X1 U5360 ( .A1(n10190), .A2(n10185), .ZN(n5168) );
  OAI21_X1 U5361 ( .B1(n10202), .B2(n6059), .A(n6058), .ZN(n10191) );
  NAND2_X1 U5362 ( .A1(n10219), .A2(n6134), .ZN(n8921) );
  INV_X1 U5363 ( .A(n8922), .ZN(n6133) );
  INV_X1 U5364 ( .A(n5080), .ZN(n5079) );
  OAI21_X1 U5365 ( .B1(n6828), .B2(n5081), .A(n6020), .ZN(n5080) );
  OR2_X1 U5366 ( .A1(n10273), .A2(n10302), .ZN(n6729) );
  NAND2_X1 U5367 ( .A1(n5501), .A2(n5502), .ZN(n10289) );
  NAND2_X1 U5368 ( .A1(n5018), .A2(n4973), .ZN(n5502) );
  NAND2_X1 U5369 ( .A1(n5493), .A2(n4996), .ZN(n5083) );
  NAND2_X1 U5370 ( .A1(n8507), .A2(n6719), .ZN(n8629) );
  AOI21_X1 U5371 ( .B1(n5507), .B2(n5509), .A(n5010), .ZN(n5506) );
  NAND2_X1 U5372 ( .A1(n8268), .A2(n5507), .ZN(n5072) );
  AND2_X1 U5373 ( .A1(n6087), .A2(n6086), .ZN(n7203) );
  NAND2_X1 U5374 ( .A1(n5454), .A2(n5045), .ZN(n5685) );
  INV_X1 U5375 ( .A(n5680), .ZN(n5455) );
  OR2_X1 U5376 ( .A1(n7663), .A2(n7662), .ZN(n5062) );
  MUX2_X1 U5377 ( .A(P2_U3893), .B(n7593), .S(n6600), .Z(n10737) );
  NAND2_X1 U5378 ( .A1(n8127), .A2(n6814), .ZN(n6672) );
  NAND2_X1 U5379 ( .A1(n6669), .A2(n4963), .ZN(n5269) );
  NAND2_X1 U5380 ( .A1(n6735), .A2(n4963), .ZN(n5275) );
  INV_X1 U5381 ( .A(n6591), .ZN(n5334) );
  NOR2_X1 U5382 ( .A1(n5331), .A2(n5334), .ZN(n5330) );
  INV_X1 U5383 ( .A(n8981), .ZN(n5331) );
  NAND2_X1 U5384 ( .A1(n6748), .A2(n6802), .ZN(n5254) );
  INV_X1 U5385 ( .A(n5291), .ZN(n5290) );
  INV_X1 U5386 ( .A(n9184), .ZN(n5213) );
  NOR2_X1 U5387 ( .A1(n5956), .A2(n5475), .ZN(n5474) );
  INV_X1 U5388 ( .A(n5937), .ZN(n5475) );
  INV_X1 U5389 ( .A(n5484), .ZN(n5479) );
  INV_X1 U5390 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8857) );
  NAND2_X1 U5391 ( .A1(n10577), .A2(n7582), .ZN(n7583) );
  NAND2_X1 U5392 ( .A1(n5436), .A2(n5435), .ZN(n7657) );
  NAND2_X1 U5393 ( .A1(n5438), .A2(n5437), .ZN(n5435) );
  NAND2_X1 U5394 ( .A1(n7733), .A2(n7682), .ZN(n10593) );
  OR2_X1 U5395 ( .A1(n7735), .A2(n7657), .ZN(n5065) );
  NAND2_X1 U5396 ( .A1(n5279), .A2(n5278), .ZN(n7685) );
  NAND2_X1 U5397 ( .A1(n7658), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U5398 ( .A1(n10593), .A2(n5280), .ZN(n5279) );
  INV_X1 U5399 ( .A(n10592), .ZN(n5280) );
  AND2_X1 U5400 ( .A1(n5049), .A2(n5048), .ZN(n9412) );
  NAND2_X1 U5401 ( .A1(n8308), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5048) );
  XNOR2_X1 U5402 ( .A(n9412), .B(n9413), .ZN(n8309) );
  INV_X1 U5403 ( .A(n5197), .ZN(n5196) );
  INV_X1 U5404 ( .A(n6585), .ZN(n5120) );
  INV_X1 U5405 ( .A(n8956), .ZN(n5119) );
  INV_X1 U5406 ( .A(n5122), .ZN(n5121) );
  OAI21_X1 U5407 ( .B1(n9209), .B2(n5307), .A(n6575), .ZN(n5306) );
  NAND2_X1 U5408 ( .A1(n7908), .A2(n7966), .ZN(n9160) );
  NAND2_X1 U5409 ( .A1(n6284), .A2(n6283), .ZN(n7783) );
  NAND2_X1 U5410 ( .A1(n6273), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6234) );
  INV_X1 U5411 ( .A(n5212), .ZN(n5211) );
  AND4_X1 U5412 ( .A1(n6208), .A2(n6199), .A3(n6404), .A4(n6392), .ZN(n6200)
         );
  INV_X1 U5413 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6199) );
  NOR2_X1 U5414 ( .A1(n6260), .A2(n6197), .ZN(n6341) );
  INV_X1 U5415 ( .A(n5099), .ZN(n5098) );
  AOI21_X1 U5416 ( .B1(n5419), .B2(n9899), .A(n5009), .ZN(n5099) );
  OAI22_X1 U5417 ( .A1(n8129), .A2(n7028), .B1(n7848), .B2(n6983), .ZN(n6984)
         );
  NAND2_X1 U5418 ( .A1(n7310), .A2(n6965), .ZN(n6973) );
  XNOR2_X1 U5419 ( .A(n6971), .B(n7176), .ZN(n6974) );
  INV_X1 U5420 ( .A(n9920), .ZN(n5426) );
  NOR2_X1 U5421 ( .A1(n5512), .A2(n6038), .ZN(n5075) );
  NOR2_X1 U5422 ( .A1(n10372), .A2(n10205), .ZN(n5074) );
  INV_X1 U5423 ( .A(n6038), .ZN(n5077) );
  INV_X1 U5424 ( .A(n6845), .ZN(n6841) );
  NAND2_X1 U5425 ( .A1(n6839), .A2(n5172), .ZN(n5171) );
  INV_X1 U5426 ( .A(n5173), .ZN(n5172) );
  NAND2_X1 U5427 ( .A1(n10238), .A2(n10243), .ZN(n10230) );
  NOR2_X1 U5428 ( .A1(n6126), .A2(n5392), .ZN(n5391) );
  INV_X1 U5429 ( .A(n6905), .ZN(n5392) );
  NOR2_X1 U5430 ( .A1(n5842), .A2(n5500), .ZN(n5499) );
  INV_X1 U5431 ( .A(n5826), .ZN(n5500) );
  INV_X1 U5432 ( .A(n6810), .ZN(n5177) );
  OR2_X1 U5433 ( .A1(n6888), .A2(n5341), .ZN(n5340) );
  OR2_X1 U5434 ( .A1(n8288), .A2(n8494), .ZN(n6663) );
  INV_X1 U5435 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5574) );
  INV_X1 U5436 ( .A(n6060), .ZN(n5488) );
  INV_X1 U5437 ( .A(n5573), .ZN(n5510) );
  AND2_X1 U5438 ( .A1(n5490), .A2(n6044), .ZN(n5489) );
  INV_X1 U5439 ( .A(n6047), .ZN(n5490) );
  NAND2_X1 U5440 ( .A1(n5562), .A2(n5234), .ZN(n5233) );
  INV_X1 U5441 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5234) );
  NOR2_X1 U5442 ( .A1(n5863), .A2(n5485), .ZN(n5484) );
  INV_X1 U5443 ( .A(n5846), .ZN(n5485) );
  INV_X1 U5444 ( .A(n5465), .ZN(n5464) );
  AOI21_X1 U5445 ( .B1(n5463), .B2(n5465), .A(n5462), .ZN(n5461) );
  INV_X1 U5446 ( .A(n5828), .ZN(n5462) );
  NOR2_X1 U5447 ( .A1(n5802), .A2(n5471), .ZN(n5470) );
  INV_X1 U5448 ( .A(n5785), .ZN(n5471) );
  OR2_X1 U5449 ( .A1(n6460), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6469) );
  AOI21_X1 U5450 ( .B1(n5150), .B2(n8994), .A(n8984), .ZN(n5149) );
  INV_X1 U5451 ( .A(n8982), .ZN(n5150) );
  INV_X1 U5452 ( .A(n5149), .ZN(n5147) );
  XNOR2_X1 U5453 ( .A(n9351), .B(n7270), .ZN(n8985) );
  XNOR2_X1 U5454 ( .A(n9518), .B(n7270), .ZN(n8976) );
  INV_X1 U5455 ( .A(n8947), .ZN(n5533) );
  NOR2_X1 U5456 ( .A1(n4975), .A2(n9128), .ZN(n5531) );
  AOI21_X1 U5457 ( .B1(n5527), .B2(n5525), .A(n5014), .ZN(n5524) );
  INV_X1 U5458 ( .A(n9024), .ZN(n5525) );
  NAND2_X1 U5459 ( .A1(n9030), .A2(n9031), .ZN(n5543) );
  NAND2_X1 U5460 ( .A1(n5138), .A2(n8944), .ZN(n5137) );
  NAND2_X1 U5461 ( .A1(n5139), .A2(n5141), .ZN(n5138) );
  OR2_X1 U5462 ( .A1(n7260), .A2(n6648), .ZN(n7299) );
  NAND2_X1 U5463 ( .A1(n5043), .A2(n9356), .ZN(n9306) );
  OAI21_X1 U5464 ( .B1(n9296), .B2(n5044), .A(n9322), .ZN(n5043) );
  OR2_X1 U5465 ( .A1(n9295), .A2(n9355), .ZN(n5044) );
  NAND2_X1 U5466 ( .A1(n9325), .A2(n9324), .ZN(n5224) );
  INV_X1 U5467 ( .A(n9323), .ZN(n9324) );
  AND4_X1 U5468 ( .A1(n6521), .A2(n6520), .A3(n6519), .A4(n6518), .ZN(n8975)
         );
  AND4_X1 U5469 ( .A1(n6301), .A2(n6300), .A3(n6299), .A4(n6298), .ZN(n8070)
         );
  OAI21_X1 U5470 ( .B1(n10571), .B2(n7571), .A(n7573), .ZN(n10574) );
  AND2_X1 U5471 ( .A1(n7575), .A2(n7574), .ZN(n7653) );
  NAND2_X1 U5472 ( .A1(n5062), .A2(n5061), .ZN(n5060) );
  NAND2_X1 U5473 ( .A1(n7978), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5061) );
  OR2_X1 U5474 ( .A1(n7984), .A2(n7983), .ZN(n5049) );
  NAND2_X1 U5475 ( .A1(n8037), .A2(n8003), .ZN(n8004) );
  NAND2_X1 U5476 ( .A1(n8004), .A2(n8005), .ZN(n8296) );
  NAND2_X1 U5477 ( .A1(n5035), .A2(n5056), .ZN(n10651) );
  NAND2_X1 U5478 ( .A1(n9419), .A2(n5450), .ZN(n5448) );
  NOR2_X1 U5479 ( .A1(n5449), .A2(n5055), .ZN(n5054) );
  INV_X1 U5480 ( .A(n5057), .ZN(n5055) );
  NAND2_X1 U5481 ( .A1(n5450), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5449) );
  NOR2_X1 U5482 ( .A1(n10651), .A2(n10650), .ZN(n10649) );
  XNOR2_X1 U5483 ( .A(n9420), .B(n10673), .ZN(n10683) );
  OR2_X1 U5484 ( .A1(n10683), .A2(n10682), .ZN(n5445) );
  INV_X1 U5485 ( .A(n9421), .ZN(n5444) );
  OR2_X1 U5486 ( .A1(n10683), .A2(n5443), .ZN(n5069) );
  NAND2_X1 U5487 ( .A1(n5446), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5443) );
  NAND2_X1 U5488 ( .A1(n9421), .A2(n5446), .ZN(n5442) );
  OAI21_X1 U5489 ( .B1(n10715), .B2(n5447), .A(n5066), .ZN(n10730) );
  NAND2_X1 U5490 ( .A1(n9425), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U5491 ( .A1(n9423), .A2(n9425), .ZN(n5066) );
  NAND2_X1 U5492 ( .A1(n6524), .A2(n4970), .ZN(n9511) );
  NAND2_X1 U5493 ( .A1(n6494), .A2(n5199), .ZN(n5198) );
  AOI21_X1 U5494 ( .B1(n5204), .B2(n4978), .A(n5011), .ZN(n5201) );
  NAND2_X1 U5495 ( .A1(n9614), .A2(n9615), .ZN(n6456) );
  NOR2_X1 U5496 ( .A1(n9649), .A2(n5229), .ZN(n5228) );
  INV_X1 U5497 ( .A(n6403), .ZN(n5229) );
  AOI21_X1 U5498 ( .B1(n9690), .B2(n5371), .A(n5008), .ZN(n5370) );
  OR2_X1 U5499 ( .A1(n9659), .A2(n9664), .ZN(n9660) );
  NAND2_X1 U5500 ( .A1(n8529), .A2(n9209), .ZN(n8530) );
  INV_X1 U5501 ( .A(n9387), .ZN(n8415) );
  NAND2_X1 U5502 ( .A1(n5302), .A2(n9336), .ZN(n5135) );
  AND4_X1 U5503 ( .A1(n6312), .A2(n6311), .A3(n6310), .A4(n6309), .ZN(n7907)
         );
  NAND2_X1 U5504 ( .A1(n6560), .A2(n5312), .ZN(n5311) );
  INV_X1 U5505 ( .A(n6559), .ZN(n5313) );
  NAND2_X1 U5506 ( .A1(n6252), .A2(n5191), .ZN(n5192) );
  NAND2_X1 U5507 ( .A1(n5019), .A2(n4982), .ZN(n5191) );
  INV_X1 U5508 ( .A(n9540), .ZN(n9684) );
  AND2_X1 U5509 ( .A1(n6221), .A2(n9464), .ZN(n7259) );
  NOR2_X1 U5510 ( .A1(n9773), .A2(n7361), .ZN(n7642) );
  NAND2_X1 U5511 ( .A1(n7240), .A2(n8545), .ZN(n5393) );
  NOR2_X1 U5512 ( .A1(n5133), .A2(n5129), .ZN(n5128) );
  INV_X1 U5513 ( .A(n6605), .ZN(n5129) );
  AND2_X1 U5514 ( .A1(n9491), .A2(n9778), .ZN(n5133) );
  NAND2_X1 U5515 ( .A1(n9143), .A2(n8505), .ZN(n9773) );
  OR2_X1 U5516 ( .A1(n9269), .A2(n6607), .ZN(n7295) );
  AND2_X1 U5517 ( .A1(n7291), .A2(n7357), .ZN(n7354) );
  NAND2_X1 U5518 ( .A1(n5219), .A2(n5318), .ZN(n5317) );
  AND2_X1 U5519 ( .A1(n5549), .A2(n6237), .ZN(n5548) );
  NOR2_X1 U5520 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5352) );
  NAND2_X1 U5521 ( .A1(n6205), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6206) );
  AOI21_X1 U5522 ( .B1(n6204), .B2(P2_IR_REG_31__SCAN_IN), .A(n5285), .ZN(
        n5284) );
  NAND2_X1 U5523 ( .A1(n5093), .A2(n5092), .ZN(n5424) );
  AOI21_X1 U5524 ( .B1(n5094), .B2(n4968), .A(n5017), .ZN(n5092) );
  NOR2_X1 U5525 ( .A1(n7030), .A2(n5422), .ZN(n5421) );
  INV_X1 U5526 ( .A(n7024), .ZN(n5422) );
  INV_X1 U5527 ( .A(n8562), .ZN(n5398) );
  NOR2_X1 U5528 ( .A1(n7136), .A2(n7135), .ZN(n7137) );
  NOR2_X1 U5529 ( .A1(n9869), .A2(n9977), .ZN(n7135) );
  NAND2_X1 U5530 ( .A1(n7031), .A2(n7030), .ZN(n8359) );
  NAND2_X1 U5531 ( .A1(n8360), .A2(n8358), .ZN(n8357) );
  NAND2_X1 U5532 ( .A1(n5100), .A2(n7055), .ZN(n9896) );
  INV_X1 U5533 ( .A(n9898), .ZN(n5100) );
  INV_X1 U5534 ( .A(n8378), .ZN(n5400) );
  INV_X1 U5535 ( .A(n5406), .ZN(n5401) );
  NOR2_X1 U5536 ( .A1(n5404), .A2(n5408), .ZN(n5402) );
  NAND2_X1 U5537 ( .A1(n6945), .A2(n7001), .ZN(n6953) );
  OAI22_X1 U5538 ( .A1(n8088), .A2(n7028), .B1(n5629), .B2(n6983), .ZN(n6952)
         );
  OR2_X1 U5539 ( .A1(n9945), .A2(n5415), .ZN(n5105) );
  NAND2_X1 U5540 ( .A1(n6799), .A2(n6798), .ZN(n6801) );
  AND2_X1 U5541 ( .A1(n5989), .A2(n5988), .ZN(n7120) );
  NOR2_X1 U5542 ( .A1(n10171), .A2(n5519), .ZN(n5518) );
  AND2_X1 U5543 ( .A1(n6100), .A2(n10149), .ZN(n10158) );
  NAND2_X1 U5544 ( .A1(n10169), .A2(n5556), .ZN(n10136) );
  NAND2_X1 U5545 ( .A1(n10280), .A2(n5173), .ZN(n5380) );
  INV_X1 U5546 ( .A(n6129), .ZN(n10250) );
  AND2_X1 U5547 ( .A1(n6729), .A2(n10250), .ZN(n10279) );
  NAND2_X1 U5548 ( .A1(n10288), .A2(n5520), .ZN(n10269) );
  AND2_X1 U5549 ( .A1(n5966), .A2(n5953), .ZN(n5520) );
  INV_X1 U5550 ( .A(n10279), .ZN(n5966) );
  INV_X1 U5551 ( .A(n5164), .ZN(n8647) );
  AOI21_X1 U5552 ( .B1(n8614), .B2(n8617), .A(n5167), .ZN(n5164) );
  OR2_X1 U5553 ( .A1(n8647), .A2(n8648), .ZN(n8645) );
  AND2_X1 U5554 ( .A1(n8648), .A2(n4977), .ZN(n5082) );
  AOI21_X1 U5555 ( .B1(n4974), .B2(n5498), .A(n4998), .ZN(n5494) );
  INV_X1 U5556 ( .A(n5841), .ZN(n5498) );
  NAND2_X1 U5557 ( .A1(n8472), .A2(n5825), .ZN(n5827) );
  AND2_X1 U5558 ( .A1(n6897), .A2(n6719), .ZN(n8509) );
  NAND2_X1 U5559 ( .A1(n8260), .A2(n6666), .ZN(n5180) );
  AND4_X1 U5560 ( .A1(n5799), .A2(n5798), .A3(n5797), .A4(n5796), .ZN(n8469)
         );
  NAND2_X1 U5561 ( .A1(n5342), .A2(n5343), .ZN(n8260) );
  NAND2_X1 U5562 ( .A1(n8268), .A2(n8267), .ZN(n8266) );
  OR2_X1 U5563 ( .A1(n6950), .A2(n10116), .ZN(n7934) );
  NAND2_X1 U5564 ( .A1(n8133), .A2(n5692), .ZN(n8106) );
  NAND2_X1 U5565 ( .A1(n6882), .A2(n6683), .ZN(n8134) );
  NAND2_X1 U5566 ( .A1(n8128), .A2(n6876), .ZN(n5348) );
  NOR2_X1 U5567 ( .A1(n8125), .A2(n8347), .ZN(n8085) );
  INV_X1 U5568 ( .A(n6120), .ZN(n5350) );
  INV_X1 U5569 ( .A(n6967), .ZN(n8076) );
  NAND2_X1 U5570 ( .A1(n7315), .A2(n10485), .ZN(n10315) );
  AND2_X1 U5571 ( .A1(n7315), .A2(n7321), .ZN(n10389) );
  NOR2_X2 U5572 ( .A1(n8011), .A2(n6150), .ZN(n10292) );
  INV_X1 U5573 ( .A(n7316), .ZN(n5941) );
  AND2_X1 U5574 ( .A1(n6167), .A2(n6191), .ZN(n7417) );
  NOR2_X1 U5575 ( .A1(n5569), .A2(n5568), .ZN(n5570) );
  NOR2_X1 U5576 ( .A1(n5866), .A2(n5482), .ZN(n5481) );
  INV_X1 U5577 ( .A(n5862), .ZN(n5482) );
  NOR2_X1 U5578 ( .A1(n5466), .A2(n5805), .ZN(n5465) );
  INV_X1 U5579 ( .A(n5468), .ZN(n5466) );
  NAND2_X1 U5580 ( .A1(n5786), .A2(n5470), .ZN(n5467) );
  NAND2_X1 U5581 ( .A1(n5469), .A2(n8755), .ZN(n5468) );
  INV_X1 U5582 ( .A(n5801), .ZN(n5469) );
  NAND2_X1 U5583 ( .A1(n5733), .A2(n5732), .ZN(n5745) );
  INV_X1 U5584 ( .A(n5114), .ZN(n5113) );
  INV_X1 U5585 ( .A(n5699), .ZN(n5115) );
  INV_X1 U5586 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U5587 ( .A1(n5184), .A2(n8805), .ZN(n5663) );
  INV_X1 U5588 ( .A(n5662), .ZN(n5184) );
  NAND2_X1 U5589 ( .A1(n5646), .A2(n5647), .ZN(n5661) );
  INV_X1 U5590 ( .A(n9801), .ZN(n9011) );
  AND4_X1 U5591 ( .A1(n6372), .A2(n6371), .A3(n6370), .A4(n6369), .ZN(n9094)
         );
  INV_X1 U5592 ( .A(n7272), .ZN(n5538) );
  AND4_X1 U5593 ( .A1(n6351), .A2(n6350), .A3(n6349), .A4(n6348), .ZN(n8577)
         );
  AND4_X1 U5594 ( .A1(n6511), .A2(n6510), .A3(n6509), .A4(n6508), .ZN(n9554)
         );
  AND4_X1 U5595 ( .A1(n6362), .A2(n6361), .A3(n6360), .A4(n6359), .ZN(n9100)
         );
  AND4_X1 U5596 ( .A1(n6465), .A2(n6464), .A3(n6463), .A4(n6462), .ZN(n9613)
         );
  INV_X1 U5597 ( .A(n9539), .ZN(n9564) );
  AND4_X1 U5598 ( .A1(n6542), .A2(n6541), .A3(n6540), .A4(n6539), .ZN(n9122)
         );
  INV_X1 U5599 ( .A(n7907), .ZN(n9389) );
  NAND2_X1 U5600 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n6277) );
  NOR2_X1 U5601 ( .A1(n10611), .A2(n7660), .ZN(n7663) );
  XNOR2_X1 U5602 ( .A(n5060), .B(n5059), .ZN(n8036) );
  XNOR2_X1 U5603 ( .A(n10761), .B(n10760), .ZN(n10770) );
  AND2_X1 U5604 ( .A1(n10759), .A2(n10758), .ZN(n10761) );
  AND2_X1 U5605 ( .A1(n10768), .A2(n10767), .ZN(n10769) );
  XNOR2_X1 U5606 ( .A(n10754), .B(n10753), .ZN(n5282) );
  AOI21_X1 U5607 ( .B1(n10757), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n10756), .ZN(
        n5283) );
  XNOR2_X1 U5608 ( .A(n5431), .B(n5430), .ZN(n5558) );
  INV_X1 U5609 ( .A(n9432), .ZN(n5430) );
  OAI21_X1 U5610 ( .B1(n10759), .B2(n10760), .A(n5432), .ZN(n5431) );
  AOI21_X1 U5611 ( .B1(n9428), .B2(n10771), .A(n5433), .ZN(n5432) );
  NAND2_X1 U5612 ( .A1(n9466), .A2(n9465), .ZN(n9467) );
  NAND2_X1 U5613 ( .A1(n9460), .A2(n10772), .ZN(n9466) );
  OR2_X1 U5614 ( .A1(n7609), .A2(n6513), .ZN(n6408) );
  NAND2_X1 U5615 ( .A1(n10851), .A2(n9771), .ZN(n9833) );
  XNOR2_X1 U5616 ( .A(n6175), .B(n6174), .ZN(n7319) );
  AOI21_X1 U5617 ( .B1(n4994), .B2(n5415), .A(n5412), .ZN(n5411) );
  INV_X1 U5618 ( .A(n7211), .ZN(n5412) );
  AND4_X1 U5619 ( .A1(n5840), .A2(n5839), .A3(n5838), .A4(n5837), .ZN(n9904)
         );
  INV_X1 U5620 ( .A(n10033), .ZN(n9925) );
  AND2_X1 U5621 ( .A1(n6019), .A2(n6018), .ZN(n9948) );
  NOR2_X1 U5622 ( .A1(n7191), .A2(n7185), .ZN(n10002) );
  INV_X1 U5623 ( .A(n10360), .ZN(n10030) );
  INV_X1 U5624 ( .A(n9948), .ZN(n10245) );
  OR2_X1 U5625 ( .A1(n5934), .A2(n5933), .ZN(n10031) );
  AOI21_X1 U5626 ( .B1(n5556), .B2(n5376), .A(n5375), .ZN(n5374) );
  NAND2_X1 U5627 ( .A1(n6075), .A2(n6074), .ZN(n5087) );
  AND2_X1 U5628 ( .A1(n6005), .A2(n6004), .ZN(n10377) );
  AND3_X1 U5629 ( .A1(n5965), .A2(n5964), .A3(n5963), .ZN(n10302) );
  NAND2_X1 U5630 ( .A1(n10157), .A2(n8917), .ZN(n5249) );
  NAND2_X1 U5631 ( .A1(n5250), .A2(n5187), .ZN(n8916) );
  INV_X1 U5632 ( .A(n10165), .ZN(n5250) );
  AND2_X1 U5633 ( .A1(n10846), .A2(n10428), .ZN(n8435) );
  NAND2_X1 U5634 ( .A1(n9189), .A2(n9188), .ZN(n9199) );
  NAND2_X1 U5635 ( .A1(n5268), .A2(n5267), .ZN(n5266) );
  NOR2_X1 U5636 ( .A1(n6896), .A2(n4963), .ZN(n5267) );
  NAND2_X1 U5637 ( .A1(n6703), .A2(n8278), .ZN(n5268) );
  NAND2_X1 U5638 ( .A1(n5296), .A2(n9227), .ZN(n9235) );
  NAND2_X1 U5639 ( .A1(n5296), .A2(n5294), .ZN(n9233) );
  INV_X1 U5640 ( .A(n9227), .ZN(n5295) );
  OAI211_X1 U5641 ( .C1(n6724), .C2(n6723), .A(n5261), .B(n6722), .ZN(n5260)
         );
  NAND2_X1 U5642 ( .A1(n9265), .A2(n9535), .ZN(n5297) );
  OAI21_X1 U5643 ( .B1(n6747), .B2(n6847), .A(n6834), .ZN(n5252) );
  NOR2_X1 U5644 ( .A1(n9285), .A2(n9284), .ZN(n9286) );
  OR2_X1 U5645 ( .A1(n9293), .A2(n9499), .ZN(n5047) );
  AND2_X1 U5646 ( .A1(n9319), .A2(n9284), .ZN(n9292) );
  NAND2_X1 U5647 ( .A1(n8321), .A2(n5109), .ZN(n5108) );
  INV_X1 U5648 ( .A(n6566), .ZN(n5109) );
  INV_X1 U5649 ( .A(n6568), .ZN(n5327) );
  INV_X1 U5650 ( .A(n5333), .ZN(n5332) );
  NAND2_X1 U5651 ( .A1(n6951), .A2(n8014), .ZN(n6970) );
  NOR2_X1 U5652 ( .A1(n6818), .A2(n5337), .ZN(n6820) );
  OR2_X1 U5653 ( .A1(n7945), .A2(n5338), .ZN(n5337) );
  INV_X1 U5654 ( .A(n6891), .ZN(n5341) );
  NOR2_X1 U5655 ( .A1(n10234), .A2(n10230), .ZN(n8926) );
  NAND2_X1 U5656 ( .A1(n6761), .A2(n6760), .ZN(n6769) );
  INV_X1 U5657 ( .A(SI_20_), .ZN(n8778) );
  INV_X1 U5658 ( .A(SI_18_), .ZN(n8777) );
  INV_X1 U5659 ( .A(SI_16_), .ZN(n8788) );
  INV_X1 U5660 ( .A(SI_17_), .ZN(n8784) );
  INV_X1 U5661 ( .A(n5470), .ZN(n5463) );
  INV_X1 U5662 ( .A(n5552), .ZN(n5141) );
  NAND2_X1 U5663 ( .A1(n5276), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10577) );
  NAND2_X1 U5664 ( .A1(n7679), .A2(n5001), .ZN(n7681) );
  NAND2_X1 U5665 ( .A1(n10607), .A2(n7686), .ZN(n7688) );
  NAND2_X1 U5666 ( .A1(n7688), .A2(n7687), .ZN(n7999) );
  INV_X1 U5667 ( .A(n10667), .ZN(n5450) );
  NAND2_X1 U5668 ( .A1(n5036), .A2(n5058), .ZN(n5057) );
  INV_X1 U5669 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5292) );
  NAND2_X1 U5670 ( .A1(n10658), .A2(n5038), .ZN(n9404) );
  INV_X1 U5671 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6392) );
  INV_X1 U5672 ( .A(n10699), .ZN(n5446) );
  NAND3_X1 U5673 ( .A1(n5069), .A2(n5068), .A3(n5442), .ZN(n5067) );
  NAND2_X1 U5674 ( .A1(n9437), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5068) );
  OR2_X1 U5675 ( .A1(n6497), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6506) );
  INV_X1 U5676 ( .A(n9615), .ZN(n5205) );
  INV_X1 U5677 ( .A(n6469), .ZN(n6468) );
  INV_X1 U5678 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8851) );
  NOR2_X1 U5679 ( .A1(n6409), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6426) );
  INV_X1 U5680 ( .A(n9834), .ZN(n9220) );
  INV_X1 U5681 ( .A(n9207), .ZN(n5371) );
  INV_X1 U5682 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8823) );
  NOR2_X1 U5683 ( .A1(n5303), .A2(n6564), .ZN(n5302) );
  INV_X1 U5684 ( .A(n5305), .ZN(n5303) );
  NAND2_X1 U5685 ( .A1(n6564), .A2(n6565), .ZN(n5305) );
  AND3_X1 U5686 ( .A1(n4988), .A2(n5318), .A3(n5549), .ZN(n5217) );
  NAND2_X1 U5687 ( .A1(n6616), .A2(n6223), .ZN(n6239) );
  INV_X1 U5688 ( .A(n6236), .ZN(n5353) );
  NAND2_X1 U5689 ( .A1(n5286), .A2(n6217), .ZN(n5285) );
  NAND2_X1 U5690 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), 
        .ZN(n5286) );
  INV_X1 U5691 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6116) );
  NOR2_X1 U5692 ( .A1(n5755), .A2(n5754), .ZN(n5777) );
  INV_X1 U5693 ( .A(n8489), .ZN(n5407) );
  NAND2_X1 U5694 ( .A1(n7857), .A2(n7000), .ZN(n7005) );
  NAND3_X1 U5695 ( .A1(n6948), .A2(n7934), .A3(n6949), .ZN(n6959) );
  OR2_X1 U5696 ( .A1(n6947), .A2(n6946), .ZN(n6948) );
  INV_X1 U5697 ( .A(n5380), .ZN(n6842) );
  INV_X1 U5698 ( .A(n6809), .ZN(n6838) );
  INV_X1 U5699 ( .A(n5914), .ZN(n5504) );
  AND2_X1 U5700 ( .A1(n8900), .A2(n4973), .ZN(n5503) );
  NAND2_X1 U5701 ( .A1(n5165), .A2(n5167), .ZN(n5162) );
  NAND2_X1 U5702 ( .A1(n5391), .A2(n8648), .ZN(n5390) );
  AND2_X1 U5703 ( .A1(n5927), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5945) );
  NOR2_X1 U5704 ( .A1(n5908), .A2(n5907), .ZN(n5927) );
  INV_X1 U5705 ( .A(n5238), .ZN(n5237) );
  NAND2_X1 U5706 ( .A1(n5497), .A2(n5841), .ZN(n5496) );
  INV_X1 U5707 ( .A(n5499), .ZN(n5497) );
  INV_X1 U5708 ( .A(n5508), .ZN(n5507) );
  OAI21_X1 U5709 ( .B1(n8267), .B2(n5509), .A(n5800), .ZN(n5508) );
  INV_X1 U5710 ( .A(n5784), .ZN(n5509) );
  NOR2_X1 U5711 ( .A1(n5350), .A2(n5349), .ZN(n5347) );
  NAND2_X1 U5712 ( .A1(n8634), .A2(n8899), .ZN(n8650) );
  NAND4_X1 U5713 ( .A1(n5523), .A2(n4972), .A3(n5231), .A4(n5230), .ZN(n5573)
         );
  AND2_X1 U5714 ( .A1(n5232), .A2(n4993), .ZN(n5231) );
  INV_X1 U5715 ( .A(n5686), .ZN(n5230) );
  INV_X1 U5716 ( .A(n5233), .ZN(n5232) );
  NOR2_X1 U5717 ( .A1(n5387), .A2(n5590), .ZN(n5386) );
  INV_X1 U5718 ( .A(n4993), .ZN(n5387) );
  XNOR2_X1 U5719 ( .A(n6769), .B(n6768), .ZN(n6767) );
  INV_X1 U5720 ( .A(SI_27_), .ZN(n8761) );
  NAND2_X1 U5721 ( .A1(n5573), .A2(n5511), .ZN(n6861) );
  NOR2_X1 U5722 ( .A1(n10474), .A2(n6146), .ZN(n5511) );
  INV_X1 U5723 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5572) );
  INV_X1 U5724 ( .A(SI_23_), .ZN(n8771) );
  AOI21_X1 U5725 ( .B1(n5476), .B2(n5474), .A(n5034), .ZN(n5473) );
  XNOR2_X1 U5726 ( .A(n5968), .B(n8778), .ZN(n5970) );
  NAND2_X1 U5727 ( .A1(n5921), .A2(SI_18_), .ZN(n5937) );
  INV_X1 U5728 ( .A(n5936), .ZN(n5476) );
  INV_X1 U5729 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5564) );
  NOR2_X1 U5730 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5565) );
  INV_X1 U5731 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5567) );
  INV_X1 U5732 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5872) );
  INV_X1 U5733 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5848) );
  INV_X1 U5734 ( .A(n5481), .ZN(n5480) );
  AOI21_X1 U5735 ( .B1(n5479), .B2(n5481), .A(n5478), .ZN(n5477) );
  INV_X1 U5736 ( .A(n5886), .ZN(n5478) );
  NOR2_X1 U5737 ( .A1(n5815), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5849) );
  INV_X1 U5738 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5809) );
  INV_X1 U5739 ( .A(n5660), .ZN(n5456) );
  AOI21_X1 U5740 ( .B1(n5460), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n5458), .ZN(
        n5457) );
  XNOR2_X1 U5741 ( .A(n8992), .B(n7270), .ZN(n8983) );
  AND2_X1 U5742 ( .A1(n6335), .A2(n8750), .ZN(n6346) );
  INV_X1 U5743 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8750) );
  XNOR2_X1 U5744 ( .A(n7265), .B(n4959), .ZN(n7266) );
  INV_X1 U5745 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8846) );
  XNOR2_X1 U5746 ( .A(n9531), .B(n7270), .ZN(n8972) );
  XNOR2_X1 U5747 ( .A(n8966), .B(n7821), .ZN(n7274) );
  NAND2_X1 U5748 ( .A1(n8938), .A2(n4990), .ZN(n9072) );
  INV_X1 U5749 ( .A(n8963), .ZN(n5528) );
  NAND2_X1 U5750 ( .A1(n9023), .A2(n9024), .ZN(n5529) );
  OR2_X1 U5751 ( .A1(n6477), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6486) );
  NAND2_X1 U5752 ( .A1(n6485), .A2(n8866), .ZN(n6497) );
  INV_X1 U5753 ( .A(n6486), .ZN(n6485) );
  OR2_X1 U5754 ( .A1(n6357), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6367) );
  NOR2_X1 U5755 ( .A1(n6367), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6376) );
  NAND2_X1 U5756 ( .A1(n6449), .A2(n8745), .ZN(n6460) );
  OR2_X1 U5757 ( .A1(n8050), .A2(n8051), .ZN(n5547) );
  NAND2_X1 U5758 ( .A1(n8823), .A2(n6397), .ZN(n6409) );
  NAND2_X1 U5759 ( .A1(n7572), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10572) );
  NOR2_X1 U5760 ( .A1(n7653), .A2(n5438), .ZN(n7654) );
  INV_X1 U5761 ( .A(n5064), .ZN(n10589) );
  INV_X1 U5762 ( .A(n5065), .ZN(n10591) );
  XNOR2_X1 U5763 ( .A(n7659), .B(n10610), .ZN(n10613) );
  XNOR2_X1 U5764 ( .A(n7685), .B(n10610), .ZN(n10608) );
  AND2_X1 U5765 ( .A1(n5064), .A2(n5063), .ZN(n7659) );
  NAND2_X1 U5766 ( .A1(n7658), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5063) );
  NAND2_X1 U5767 ( .A1(n7999), .A2(n5277), .ZN(n8002) );
  NAND2_X1 U5768 ( .A1(n7978), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5277) );
  NAND2_X1 U5769 ( .A1(n8296), .A2(n8297), .ZN(n9396) );
  NAND2_X1 U5770 ( .A1(n5453), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U5771 ( .A1(n9415), .A2(n5453), .ZN(n5451) );
  INV_X1 U5772 ( .A(n10635), .ZN(n5453) );
  NOR2_X1 U5773 ( .A1(n8309), .A2(n8324), .ZN(n9414) );
  NAND2_X1 U5774 ( .A1(n10645), .A2(n9402), .ZN(n10659) );
  NAND2_X1 U5775 ( .A1(n10659), .A2(n10660), .ZN(n10658) );
  XNOR2_X1 U5776 ( .A(n9404), .B(n10673), .ZN(n10675) );
  XNOR2_X1 U5777 ( .A(n5067), .B(n9435), .ZN(n10715) );
  NOR2_X1 U5778 ( .A1(n10715), .A2(n10714), .ZN(n10713) );
  NAND2_X1 U5779 ( .A1(n9426), .A2(n10738), .ZN(n5434) );
  INV_X1 U5780 ( .A(n6601), .ZN(n7577) );
  NOR2_X1 U5781 ( .A1(n10758), .A2(n9427), .ZN(n5433) );
  NAND2_X1 U5782 ( .A1(n10758), .A2(n9427), .ZN(n9428) );
  NAND2_X1 U5783 ( .A1(n4981), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n10759) );
  INV_X1 U5784 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n9461) );
  OR2_X1 U5785 ( .A1(n6545), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n9473) );
  AOI21_X1 U5786 ( .B1(n5200), .B2(n5197), .A(n5195), .ZN(n5194) );
  INV_X1 U5787 ( .A(n9266), .ZN(n5195) );
  NAND2_X1 U5788 ( .A1(n6505), .A2(n8732), .ZN(n6516) );
  INV_X1 U5789 ( .A(n6506), .ZN(n6505) );
  OR2_X1 U5790 ( .A1(n6516), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6528) );
  NAND2_X1 U5791 ( .A1(n5309), .A2(n5308), .ZN(n9537) );
  AND2_X1 U5792 ( .A1(n9547), .A2(n6588), .ZN(n5308) );
  NAND2_X1 U5793 ( .A1(n5117), .A2(n5116), .ZN(n9588) );
  AOI21_X1 U5794 ( .B1(n5118), .B2(n5121), .A(n5366), .ZN(n5116) );
  INV_X1 U5795 ( .A(n5306), .ZN(n5125) );
  NOR2_X1 U5796 ( .A1(n6385), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6397) );
  NAND2_X1 U5797 ( .A1(n8846), .A2(n6376), .ZN(n6385) );
  NAND2_X1 U5798 ( .A1(n7819), .A2(n9160), .ZN(n7865) );
  NAND2_X1 U5799 ( .A1(n7629), .A2(n9148), .ZN(n7717) );
  NAND2_X1 U5800 ( .A1(n5190), .A2(n5189), .ZN(n7629) );
  OR3_X1 U5801 ( .A1(n7643), .A2(n9464), .A3(n6220), .ZN(n7878) );
  NAND2_X1 U5802 ( .A1(n7641), .A2(n7640), .ZN(n7647) );
  NAND2_X1 U5803 ( .A1(n6267), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6233) );
  XNOR2_X1 U5804 ( .A(n7232), .B(n6592), .ZN(n6606) );
  INV_X1 U5805 ( .A(n9351), .ZN(n6592) );
  NAND2_X1 U5806 ( .A1(n9495), .A2(n6591), .ZN(n7232) );
  NAND2_X1 U5807 ( .A1(n9291), .A2(n9290), .ZN(n9298) );
  AND2_X1 U5808 ( .A1(n7259), .A2(n8505), .ZN(n7241) );
  NAND2_X1 U5809 ( .A1(n9637), .A2(n9225), .ZN(n9625) );
  OAI21_X1 U5810 ( .B1(n8029), .B2(n5211), .A(n5209), .ZN(n8462) );
  NAND2_X1 U5811 ( .A1(n6560), .A2(n6559), .ZN(n7822) );
  INV_X1 U5812 ( .A(n6635), .ZN(n5155) );
  AND2_X1 U5813 ( .A1(n6215), .A2(n5320), .ZN(n5319) );
  NOR2_X1 U5814 ( .A1(n5321), .A2(n6260), .ZN(n5320) );
  NAND2_X1 U5815 ( .A1(n5322), .A2(n5323), .ZN(n5321) );
  INV_X1 U5816 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6202) );
  NAND2_X1 U5817 ( .A1(n6260), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6303) );
  NAND2_X1 U5818 ( .A1(n4971), .A2(n5416), .ZN(n5415) );
  INV_X1 U5819 ( .A(n7149), .ZN(n5416) );
  AND2_X1 U5820 ( .A1(n7172), .A2(n7171), .ZN(n7212) );
  INV_X1 U5821 ( .A(n6959), .ZN(n7173) );
  AND2_X1 U5822 ( .A1(n10011), .A2(n5426), .ZN(n5097) );
  INV_X1 U5823 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5754) );
  OR2_X1 U5824 ( .A1(n6949), .A2(n6957), .ZN(n6958) );
  NAND2_X1 U5825 ( .A1(n7115), .A2(n9955), .ZN(n9958) );
  INV_X1 U5826 ( .A(n7060), .ZN(n5420) );
  OR2_X1 U5827 ( .A1(n5819), .A2(n7545), .ZN(n5835) );
  OR2_X1 U5828 ( .A1(n5835), .A2(n5834), .ZN(n5853) );
  NAND2_X1 U5829 ( .A1(n6976), .A2(n6975), .ZN(n5394) );
  INV_X1 U5830 ( .A(n7088), .ZN(n5096) );
  INV_X1 U5831 ( .A(n5095), .ZN(n5094) );
  OAI21_X1 U5832 ( .B1(n4968), .B2(n5426), .A(n7093), .ZN(n5095) );
  OR2_X1 U5833 ( .A1(n9930), .A2(n9929), .ZN(n7093) );
  NAND2_X1 U5834 ( .A1(n4971), .A2(n9909), .ZN(n5414) );
  AND2_X1 U5835 ( .A1(n6947), .A2(n6117), .ZN(n7315) );
  OAI21_X1 U5836 ( .B1(n6794), .B2(n10439), .A(n5258), .ZN(n5257) );
  AND2_X1 U5837 ( .A1(n6793), .A2(n5259), .ZN(n5258) );
  NAND2_X1 U5838 ( .A1(n10439), .A2(n4963), .ZN(n5259) );
  AND2_X1 U5839 ( .A1(n6852), .A2(n10138), .ZN(n6793) );
  INV_X1 U5840 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7449) );
  INV_X1 U5841 ( .A(n5378), .ZN(n5376) );
  INV_X1 U5842 ( .A(n5556), .ZN(n5377) );
  NOR2_X1 U5843 ( .A1(n6750), .A2(n5516), .ZN(n5515) );
  INV_X1 U5844 ( .A(n6088), .ZN(n5516) );
  AND2_X1 U5845 ( .A1(n6106), .A2(n6105), .ZN(n10172) );
  AND2_X1 U5846 ( .A1(n10186), .A2(n6746), .ZN(n10170) );
  NAND2_X1 U5847 ( .A1(n5079), .A2(n5077), .ZN(n5076) );
  INV_X1 U5848 ( .A(n10237), .ZN(n5078) );
  AND2_X1 U5849 ( .A1(n6037), .A2(n6036), .ZN(n10222) );
  INV_X1 U5850 ( .A(n5379), .ZN(n10220) );
  OR2_X1 U5851 ( .A1(n6828), .A2(n5171), .ZN(n5169) );
  INV_X1 U5852 ( .A(n10252), .ZN(n10256) );
  NAND2_X1 U5853 ( .A1(n8645), .A2(n5391), .ZN(n10309) );
  NAND2_X1 U5854 ( .A1(n8634), .A2(n5236), .ZN(n10323) );
  OR2_X1 U5855 ( .A1(n5892), .A2(n8455), .ZN(n5908) );
  NAND2_X1 U5856 ( .A1(n5495), .A2(n5841), .ZN(n8627) );
  NAND2_X1 U5857 ( .A1(n5827), .A2(n5499), .ZN(n5495) );
  AND2_X1 U5858 ( .A1(n5021), .A2(n6812), .ZN(n5179) );
  AND2_X1 U5859 ( .A1(n6889), .A2(n8391), .ZN(n8261) );
  NAND2_X1 U5860 ( .A1(n7398), .A2(n6785), .ZN(n5175) );
  AND2_X1 U5861 ( .A1(n6663), .A2(n6819), .ZN(n8281) );
  INV_X1 U5862 ( .A(n6694), .ZN(n8231) );
  INV_X1 U5863 ( .A(n8225), .ZN(n8244) );
  INV_X1 U5864 ( .A(n10038), .ZN(n8229) );
  OR2_X1 U5865 ( .A1(n8125), .A2(n5246), .ZN(n8136) );
  INV_X1 U5866 ( .A(n5245), .ZN(n5246) );
  OR2_X1 U5867 ( .A1(n8125), .A2(n5244), .ZN(n8137) );
  NAND2_X1 U5868 ( .A1(n5245), .A2(n7890), .ZN(n5244) );
  AND4_X1 U5869 ( .A1(n5698), .A2(n5697), .A3(n5696), .A4(n5695), .ZN(n8243)
         );
  INV_X1 U5870 ( .A(n8134), .ZN(n8140) );
  NAND2_X1 U5871 ( .A1(n7938), .A2(n5670), .ZN(n8135) );
  NAND2_X1 U5872 ( .A1(n8135), .A2(n8134), .ZN(n8133) );
  AND4_X1 U5873 ( .A1(n5678), .A2(n5677), .A3(n5676), .A4(n5675), .ZN(n8107)
         );
  NAND2_X1 U5874 ( .A1(n7939), .A2(n7945), .ZN(n7938) );
  OR2_X1 U5875 ( .A1(n8123), .A2(n6945), .ZN(n8125) );
  AND4_X1 U5876 ( .A1(n5635), .A2(n5634), .A3(n5633), .A4(n5632), .ZN(n8129)
         );
  NAND2_X1 U5877 ( .A1(n6192), .A2(n10473), .ZN(n7970) );
  INV_X1 U5878 ( .A(n10167), .ZN(n5188) );
  INV_X1 U5879 ( .A(n6787), .ZN(n5942) );
  INV_X1 U5880 ( .A(n10292), .ZN(n10803) );
  OR2_X1 U5881 ( .A1(n6189), .A2(n7931), .ZN(n7971) );
  NOR2_X1 U5882 ( .A1(n8011), .A2(n6934), .ZN(n10428) );
  OR2_X1 U5883 ( .A1(n6947), .A2(n6117), .ZN(n8011) );
  XNOR2_X1 U5884 ( .A(n6147), .B(P1_IR_REG_28__SCAN_IN), .ZN(n7321) );
  INV_X1 U5885 ( .A(n5487), .ZN(n5486) );
  OAI21_X1 U5886 ( .B1(n5489), .B2(n5037), .A(n6078), .ZN(n5487) );
  NAND2_X1 U5887 ( .A1(n6061), .A2(n6060), .ZN(n6080) );
  NAND2_X1 U5888 ( .A1(n5939), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U5889 ( .A1(n5847), .A2(n5846), .ZN(n5864) );
  INV_X1 U5890 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5810) );
  INV_X1 U5891 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8745) );
  NAND2_X1 U5892 ( .A1(n5113), .A2(n5115), .ZN(n5111) );
  NAND2_X1 U5893 ( .A1(n5579), .A2(n7845), .ZN(n5071) );
  AND2_X1 U5894 ( .A1(n5547), .A2(n4986), .ZN(n8177) );
  NAND2_X1 U5895 ( .A1(n5547), .A2(n4987), .ZN(n8175) );
  NAND2_X1 U5896 ( .A1(n8995), .A2(n8994), .ZN(n8993) );
  INV_X1 U5897 ( .A(n9381), .ZN(n9667) );
  NAND2_X1 U5898 ( .A1(n9072), .A2(n5552), .ZN(n9001) );
  NAND2_X1 U5899 ( .A1(n9017), .A2(n9016), .ZN(n9015) );
  OR2_X1 U5900 ( .A1(n9119), .A2(n5148), .ZN(n5143) );
  NAND2_X1 U5901 ( .A1(n8994), .A2(n8985), .ZN(n5148) );
  NOR2_X1 U5902 ( .A1(n8985), .A2(n5147), .ZN(n5146) );
  OAI22_X1 U5903 ( .A1(n5147), .A2(n5145), .B1(n8985), .B2(n5149), .ZN(n5144)
         );
  NOR2_X1 U5904 ( .A1(n8985), .A2(n8994), .ZN(n5145) );
  NOR2_X1 U5905 ( .A1(n7612), .A2(n7613), .ZN(n7611) );
  AND4_X1 U5906 ( .A1(n6474), .A2(n6473), .A3(n6472), .A4(n6471), .ZN(n9603)
         );
  NAND2_X1 U5907 ( .A1(n9063), .A2(n8961), .ZN(n9023) );
  OAI21_X1 U5908 ( .B1(n9091), .B2(n5153), .A(n5152), .ZN(n5151) );
  INV_X1 U5909 ( .A(n8590), .ZN(n5153) );
  INV_X1 U5910 ( .A(n8589), .ZN(n5152) );
  AND4_X1 U5911 ( .A1(n6455), .A2(n6454), .A3(n6453), .A4(n6452), .ZN(n9623)
         );
  AOI21_X1 U5912 ( .B1(n9038), .B2(n9380), .A(n5533), .ZN(n5532) );
  NAND2_X1 U5913 ( .A1(n5541), .A2(n9391), .ZN(n5540) );
  AOI21_X1 U5914 ( .B1(n8418), .B2(n8417), .A(n5554), .ZN(n8420) );
  NAND2_X1 U5915 ( .A1(n8420), .A2(n8419), .ZN(n8575) );
  INV_X1 U5916 ( .A(n9134), .ZN(n9111) );
  NAND2_X1 U5917 ( .A1(n9015), .A2(n8958), .ZN(n9065) );
  NAND2_X1 U5918 ( .A1(n8938), .A2(n8937), .ZN(n9074) );
  AND2_X1 U5919 ( .A1(n7290), .A2(n7642), .ZN(n9079) );
  NAND2_X1 U5920 ( .A1(n5529), .A2(n5527), .ZN(n9085) );
  INV_X1 U5921 ( .A(n5539), .ZN(n7618) );
  AND4_X1 U5922 ( .A1(n6443), .A2(n6442), .A3(n6441), .A4(n6440), .ZN(n9636)
         );
  INV_X1 U5923 ( .A(n9132), .ZN(n9113) );
  AND2_X1 U5924 ( .A1(n7303), .A2(n7302), .ZN(n9132) );
  NAND2_X1 U5925 ( .A1(n5543), .A2(n8977), .ZN(n9117) );
  NAND2_X1 U5926 ( .A1(n7303), .A2(n7301), .ZN(n9134) );
  NAND2_X1 U5927 ( .A1(n7298), .A2(n7297), .ZN(n9136) );
  NAND2_X1 U5928 ( .A1(n5224), .A2(n9327), .ZN(n5223) );
  XNOR2_X1 U5929 ( .A(n6216), .B(P2_IR_REG_22__SCAN_IN), .ZN(n9369) );
  INV_X1 U5930 ( .A(n8975), .ZN(n9542) );
  INV_X1 U5931 ( .A(n9576), .ZN(n9375) );
  INV_X1 U5932 ( .A(n9613), .ZN(n9378) );
  INV_X1 U5933 ( .A(n9623), .ZN(n8952) );
  INV_X1 U5934 ( .A(n8070), .ZN(n9390) );
  INV_X1 U5935 ( .A(P2_U3893), .ZN(n10766) );
  NAND4_X1 U5936 ( .A1(n6250), .A2(n6249), .A3(n6248), .A4(n6247), .ZN(n6552)
         );
  INV_X1 U5937 ( .A(n7652), .ZN(n10590) );
  XNOR2_X1 U5938 ( .A(n8002), .B(n7979), .ZN(n8038) );
  NOR2_X1 U5939 ( .A1(n8034), .A2(n7981), .ZN(n7984) );
  INV_X1 U5940 ( .A(n5060), .ZN(n7980) );
  INV_X1 U5941 ( .A(n5049), .ZN(n8307) );
  XNOR2_X1 U5942 ( .A(n9396), .B(n9413), .ZN(n8298) );
  NOR2_X1 U5943 ( .A1(n5544), .A2(n6260), .ZN(n6353) );
  NAND2_X1 U5944 ( .A1(n5448), .A2(n5052), .ZN(n10666) );
  INV_X1 U5945 ( .A(n5445), .ZN(n10681) );
  NAND2_X1 U5946 ( .A1(n5069), .A2(n5442), .ZN(n10698) );
  AND2_X1 U5947 ( .A1(n6432), .A2(n6422), .ZN(n10721) );
  XNOR2_X1 U5948 ( .A(n7225), .B(n9353), .ZN(n7240) );
  NOR2_X1 U5949 ( .A1(n6604), .A2(n6603), .ZN(n6605) );
  NAND2_X1 U5950 ( .A1(n9511), .A2(n9508), .ZN(n9493) );
  NAND2_X1 U5951 ( .A1(n9261), .A2(n5198), .ZN(n9548) );
  NAND2_X1 U5952 ( .A1(n5198), .A2(n5197), .ZN(n9712) );
  NAND2_X1 U5953 ( .A1(n6494), .A2(n6493), .ZN(n9556) );
  NAND2_X1 U5954 ( .A1(n5358), .A2(n5362), .ZN(n9581) );
  OR2_X1 U5955 ( .A1(n6456), .A2(n5365), .ZN(n5358) );
  NAND2_X1 U5956 ( .A1(n6456), .A2(n5367), .ZN(n5361) );
  NAND2_X1 U5957 ( .A1(n9660), .A2(n5228), .ZN(n9650) );
  NAND2_X1 U5958 ( .A1(n9691), .A2(n9690), .ZN(n9689) );
  NAND2_X1 U5959 ( .A1(n5372), .A2(n9207), .ZN(n9691) );
  NAND2_X1 U5960 ( .A1(n8528), .A2(n9344), .ZN(n5372) );
  NAND2_X1 U5961 ( .A1(n8530), .A2(n6574), .ZN(n9680) );
  NAND2_X1 U5962 ( .A1(n5328), .A2(n6568), .ZN(n8460) );
  NAND2_X1 U5963 ( .A1(n8320), .A2(n8321), .ZN(n5328) );
  NAND2_X1 U5964 ( .A1(n5214), .A2(n9184), .ZN(n8326) );
  NAND2_X1 U5965 ( .A1(n8029), .A2(n5215), .ZN(n5214) );
  NAND2_X1 U5966 ( .A1(n8029), .A2(n9191), .ZN(n8192) );
  OAI21_X1 U5967 ( .B1(n8068), .B2(n6565), .A(n6564), .ZN(n8023) );
  NAND2_X1 U5968 ( .A1(n5311), .A2(n5314), .ZN(n7866) );
  OR2_X1 U5969 ( .A1(n7647), .A2(n9678), .ZN(n9652) );
  INV_X1 U5970 ( .A(n9669), .ZN(n9688) );
  NAND2_X1 U5971 ( .A1(n7642), .A2(n7259), .ZN(n9669) );
  NAND2_X1 U5972 ( .A1(n6606), .A2(n5128), .ZN(n5127) );
  INV_X1 U5973 ( .A(n9298), .ZN(n9787) );
  INV_X1 U5974 ( .A(n8992), .ZN(n9791) );
  INV_X1 U5975 ( .A(n9258), .ZN(n9805) );
  INV_X1 U5976 ( .A(n9106), .ZN(n9821) );
  OAI21_X1 U5977 ( .B1(n7289), .B2(n6652), .A(n6651), .ZN(n6653) );
  INV_X1 U5978 ( .A(n7354), .ZN(n7361) );
  INV_X1 U5979 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6226) );
  INV_X1 U5980 ( .A(n9369), .ZN(n8505) );
  INV_X1 U5981 ( .A(n7262), .ZN(n9143) );
  INV_X1 U5982 ( .A(n10689), .ZN(n9437) );
  INV_X1 U5983 ( .A(n10623), .ZN(n9417) );
  INV_X1 U5984 ( .A(n7998), .ZN(n8308) );
  AND2_X1 U5985 ( .A1(n4965), .A2(P2_U3151), .ZN(n9846) );
  INV_X1 U5986 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5581) );
  NAND2_X1 U5987 ( .A1(n6244), .A2(n6243), .ZN(n10571) );
  MUX2_X1 U5988 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6241), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n6244) );
  NAND2_X1 U5989 ( .A1(n5403), .A2(n8378), .ZN(n8491) );
  OR2_X1 U5990 ( .A1(n8381), .A2(n8377), .ZN(n5403) );
  NAND2_X1 U5991 ( .A1(n5424), .A2(n5425), .ZN(n9880) );
  AND4_X1 U5992 ( .A1(n5760), .A2(n5759), .A3(n5758), .A4(n5757), .ZN(n8494)
         );
  AOI21_X1 U5993 ( .B1(n5402), .B2(n5399), .A(n5398), .ZN(n5397) );
  NAND2_X1 U5994 ( .A1(n7031), .A2(n5103), .ZN(n5102) );
  NAND2_X1 U5995 ( .A1(n5427), .A2(n10011), .ZN(n9919) );
  NAND2_X1 U5996 ( .A1(n9917), .A2(n7088), .ZN(n9932) );
  AND2_X1 U5997 ( .A1(n7142), .A2(n9941), .ZN(n7147) );
  AND4_X1 U5998 ( .A1(n5743), .A2(n5742), .A3(n5741), .A4(n5740), .ZN(n8385)
         );
  NAND2_X1 U5999 ( .A1(n9896), .A2(n7060), .ZN(n9966) );
  INV_X1 U6000 ( .A(n10017), .ZN(n9991) );
  OR2_X1 U6001 ( .A1(n8381), .A2(n5402), .ZN(n5396) );
  OAI211_X1 U6002 ( .C1(n10011), .C2(n4968), .A(n5091), .B(n5094), .ZN(n9990)
         );
  OR2_X1 U6003 ( .A1(n5427), .A2(n4968), .ZN(n5091) );
  INV_X1 U6004 ( .A(n10020), .ZN(n10003) );
  NAND2_X1 U6005 ( .A1(n7200), .A2(n7749), .ZN(n10015) );
  INV_X1 U6006 ( .A(n10002), .ZN(n10026) );
  AOI21_X1 U6007 ( .B1(n5256), .B2(n5255), .A(n6803), .ZN(n6870) );
  NOR2_X1 U6008 ( .A1(n6800), .A2(n6805), .ZN(n5255) );
  OAI21_X1 U6009 ( .B1(n6854), .B2(n4963), .A(n6117), .ZN(n6803) );
  NAND2_X1 U6010 ( .A1(n6801), .A2(n5257), .ZN(n5256) );
  INV_X1 U6011 ( .A(n7203), .ZN(n10188) );
  INV_X1 U6012 ( .A(n10208), .ZN(n7768) );
  INV_X1 U6013 ( .A(n10222), .ZN(n10205) );
  INV_X1 U6014 ( .A(n8469), .ZN(n10036) );
  AND2_X1 U6015 ( .A1(n7343), .A2(n7342), .ZN(n10560) );
  OR2_X1 U6016 ( .A1(n10563), .A2(n10554), .ZN(n10122) );
  INV_X1 U6017 ( .A(n5182), .ZN(n5181) );
  AND2_X1 U6018 ( .A1(n6057), .A2(n6056), .ZN(n10360) );
  OAI21_X1 U6019 ( .B1(n10237), .B2(n5081), .A(n5079), .ZN(n8919) );
  NAND2_X1 U6020 ( .A1(n5513), .A2(n6006), .ZN(n10226) );
  NAND2_X1 U6021 ( .A1(n10237), .A2(n6828), .ZN(n5513) );
  NAND2_X1 U6022 ( .A1(n5380), .A2(n6839), .ZN(n10244) );
  OR2_X1 U6023 ( .A1(n8220), .A2(n5659), .ZN(n5981) );
  NAND2_X1 U6024 ( .A1(n10280), .A2(n6729), .ZN(n10251) );
  AND3_X1 U6025 ( .A1(n5951), .A2(n5950), .A3(n5949), .ZN(n10396) );
  NAND2_X1 U6026 ( .A1(n10288), .A2(n5953), .ZN(n10271) );
  NAND2_X1 U6027 ( .A1(n8905), .A2(n8900), .ZN(n5505) );
  NAND2_X1 U6028 ( .A1(n8645), .A2(n6905), .ZN(n8901) );
  AND2_X1 U6029 ( .A1(n5083), .A2(n4977), .ZN(n8644) );
  AND4_X1 U6030 ( .A1(n5858), .A2(n5857), .A3(n5856), .A4(n5855), .ZN(n10021)
         );
  NAND2_X1 U6031 ( .A1(n5827), .A2(n5826), .ZN(n8506) );
  NAND2_X1 U6032 ( .A1(n5180), .A2(n6812), .ZN(n8468) );
  AND4_X1 U6033 ( .A1(n5783), .A2(n5782), .A3(n5781), .A4(n5780), .ZN(n8431)
         );
  NAND2_X1 U6034 ( .A1(n8266), .A2(n5784), .ZN(n8395) );
  NAND2_X1 U6035 ( .A1(n10328), .A2(n7940), .ZN(n10325) );
  OAI21_X1 U6036 ( .B1(n6121), .B2(n8128), .A(n5345), .ZN(n8090) );
  AOI21_X1 U6037 ( .B1(n6814), .B2(n5350), .A(n5349), .ZN(n5345) );
  OR2_X1 U6038 ( .A1(n7941), .A2(n4966), .ZN(n10264) );
  INV_X1 U6039 ( .A(n10325), .ZN(n10297) );
  NAND2_X1 U6040 ( .A1(n7941), .A2(n10326), .ZN(n10328) );
  AND2_X1 U6041 ( .A1(n10842), .A2(n10428), .ZN(n8917) );
  INV_X1 U6042 ( .A(n6852), .ZN(n10435) );
  AND2_X1 U6043 ( .A1(n10348), .A2(n10347), .ZN(n10349) );
  INV_X1 U6044 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n5186) );
  INV_X1 U6045 ( .A(n5084), .ZN(n10441) );
  NOR2_X1 U6046 ( .A1(n10354), .A2(n5086), .ZN(n5085) );
  AND2_X1 U6047 ( .A1(n10355), .A2(n10292), .ZN(n5086) );
  INV_X1 U6048 ( .A(n10234), .ZN(n10455) );
  INV_X1 U6049 ( .A(n8516), .ZN(n9975) );
  INV_X1 U6050 ( .A(n8435), .ZN(n10469) );
  AND2_X1 U6051 ( .A1(n5691), .A2(n5022), .ZN(n5088) );
  OR2_X1 U6052 ( .A1(n6787), .A2(n7366), .ZN(n5649) );
  INV_X1 U6053 ( .A(n5492), .ZN(n5491) );
  OR2_X1 U6054 ( .A1(n5659), .A2(n7352), .ZN(n5589) );
  OAI22_X1 U6055 ( .A1(n6787), .A2(n5458), .B1(n7316), .B2(n7349), .ZN(n5492)
         );
  INV_X2 U6056 ( .A(n10843), .ZN(n10846) );
  NAND2_X1 U6057 ( .A1(n7418), .A2(n7750), .ZN(n10497) );
  NAND2_X1 U6058 ( .A1(n5719), .A2(n5523), .ZN(n5924) );
  NAND2_X1 U6059 ( .A1(n5483), .A2(n5481), .ZN(n5887) );
  NAND2_X1 U6060 ( .A1(n5467), .A2(n5465), .ZN(n5829) );
  NAND2_X1 U6061 ( .A1(n5467), .A2(n5468), .ZN(n5806) );
  NAND2_X1 U6062 ( .A1(n5786), .A2(n5785), .ZN(n5803) );
  NAND2_X1 U6063 ( .A1(n5773), .A2(n5786), .ZN(n7397) );
  NAND2_X1 U6064 ( .A1(n5700), .A2(n5699), .ZN(n5705) );
  NAND2_X1 U6065 ( .A1(n5660), .A2(n5661), .ZN(n5679) );
  INV_X1 U6066 ( .A(n5062), .ZN(n7977) );
  NAND2_X1 U6067 ( .A1(n5282), .A2(n10745), .ZN(n5281) );
  AOI21_X1 U6068 ( .B1(n5558), .B2(n9468), .A(n9467), .ZN(n9469) );
  NAND2_X1 U6069 ( .A1(n5132), .A2(n5130), .ZN(P2_U3487) );
  NOR2_X1 U6070 ( .A1(n5030), .A2(n5131), .ZN(n5130) );
  NAND2_X1 U6071 ( .A1(n5127), .A2(n5126), .ZN(n5132) );
  NOR2_X1 U6072 ( .A1(n9781), .A2(n6643), .ZN(n5131) );
  OAI21_X1 U6073 ( .B1(n9480), .B2(n9833), .A(n7245), .ZN(n7246) );
  OAI21_X1 U6074 ( .B1(n6149), .B2(n10009), .A(n7217), .ZN(n7218) );
  NAND2_X1 U6075 ( .A1(n5249), .A2(n5248), .ZN(n5247) );
  NAND2_X1 U6076 ( .A1(n10840), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5248) );
  NAND2_X1 U6077 ( .A1(n10843), .A2(n5186), .ZN(n5185) );
  XNOR2_X1 U6078 ( .A(n6206), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7262) );
  OR2_X1 U6079 ( .A1(n7094), .A2(n5096), .ZN(n4968) );
  NAND2_X1 U6080 ( .A1(n5319), .A2(n4988), .ZN(n4969) );
  INV_X1 U6081 ( .A(n7001), .ZN(n7028) );
  OAI21_X1 U6082 ( .B1(n7371), .B2(n5659), .A(n5088), .ZN(n8172) );
  NAND2_X1 U6083 ( .A1(n5589), .A2(n5491), .ZN(n6967) );
  INV_X1 U6084 ( .A(n6828), .ZN(n5514) );
  AND2_X1 U6085 ( .A1(n6523), .A2(n9277), .ZN(n4970) );
  INV_X1 U6086 ( .A(n8128), .ZN(n6814) );
  NOR2_X1 U6087 ( .A1(n6279), .A2(n6278), .ZN(n7680) );
  NOR2_X1 U6088 ( .A1(n9998), .A2(n9999), .ZN(n4971) );
  AND3_X1 U6089 ( .A1(n6159), .A2(n5571), .A3(n6110), .ZN(n4972) );
  OR2_X1 U6090 ( .A1(n10324), .A2(n10031), .ZN(n4973) );
  AND2_X1 U6091 ( .A1(n8628), .A2(n5496), .ZN(n4974) );
  NOR2_X1 U6092 ( .A1(n9038), .A2(n9380), .ZN(n4975) );
  OR2_X1 U6093 ( .A1(n10195), .A2(n10198), .ZN(n4976) );
  NAND2_X1 U6094 ( .A1(n8899), .A2(n9925), .ZN(n4977) );
  AND2_X1 U6095 ( .A1(n5359), .A2(n5206), .ZN(n4978) );
  NOR2_X1 U6096 ( .A1(n9965), .A2(n5420), .ZN(n5419) );
  AND2_X1 U6097 ( .A1(n7279), .A2(n8191), .ZN(n4979) );
  NOR2_X1 U6098 ( .A1(n9390), .A2(n7915), .ZN(n4980) );
  AND2_X1 U6099 ( .A1(n10758), .A2(n5434), .ZN(n4981) );
  NAND2_X1 U6100 ( .A1(n4964), .A2(n5581), .ZN(n4982) );
  INV_X1 U6101 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6223) );
  INV_X1 U6102 ( .A(n7628), .ZN(n5190) );
  AND2_X1 U6103 ( .A1(n5236), .A2(n5235), .ZN(n4983) );
  AND2_X1 U6104 ( .A1(n8959), .A2(n8958), .ZN(n4984) );
  INV_X1 U6105 ( .A(n8001), .ZN(n7978) );
  INV_X1 U6106 ( .A(n7979), .ZN(n5059) );
  NAND2_X1 U6107 ( .A1(n5136), .A2(n8945), .ZN(n9129) );
  OR3_X1 U6108 ( .A1(n5544), .A2(n6260), .A3(P2_IR_REG_10__SCAN_IN), .ZN(n4985) );
  INV_X2 U6109 ( .A(n10840), .ZN(n10842) );
  INV_X1 U6110 ( .A(n10641), .ZN(n5058) );
  AND2_X1 U6111 ( .A1(n9167), .A2(n9160), .ZN(n7816) );
  NAND2_X1 U6112 ( .A1(n7278), .A2(n9389), .ZN(n4986) );
  AND2_X1 U6113 ( .A1(n4986), .A2(n8176), .ZN(n4987) );
  INV_X1 U6114 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5323) );
  OAI211_X1 U6115 ( .C1(n7316), .C2(n10061), .A(n5650), .B(n5649), .ZN(n8347)
         );
  NAND2_X1 U6116 ( .A1(n6170), .A2(n6169), .ZN(n6949) );
  NAND2_X1 U6117 ( .A1(n6242), .A2(n6195), .ZN(n6261) );
  NAND2_X1 U6118 ( .A1(n6154), .A2(n5572), .ZN(n6157) );
  INV_X1 U6119 ( .A(n5617), .ZN(n7346) );
  NOR2_X1 U6120 ( .A1(n6611), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n4988) );
  NOR2_X1 U6121 ( .A1(n8583), .A2(n9386), .ZN(n4989) );
  AND2_X1 U6122 ( .A1(n8939), .A2(n8937), .ZN(n4990) );
  NOR2_X1 U6123 ( .A1(n5686), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5688) );
  NAND2_X1 U6124 ( .A1(n5719), .A2(n5563), .ZN(n5734) );
  AND3_X1 U6125 ( .A1(n6272), .A2(n6271), .A3(n6270), .ZN(n4991) );
  INV_X1 U6126 ( .A(n8628), .ZN(n5263) );
  AND4_X1 U6127 ( .A1(n6907), .A2(n6802), .A3(n6898), .A4(n6902), .ZN(n4992)
         );
  XNOR2_X1 U6128 ( .A(n6767), .B(SI_29_), .ZN(n9841) );
  AND2_X1 U6129 ( .A1(n5572), .A2(n5388), .ZN(n4993) );
  XNOR2_X1 U6130 ( .A(n8967), .B(n8968), .ZN(n9007) );
  AND2_X1 U6131 ( .A1(n5414), .A2(n5413), .ZN(n4994) );
  NAND2_X1 U6132 ( .A1(n5355), .A2(n6292), .ZN(n7966) );
  OR2_X1 U6133 ( .A1(n8583), .A2(n9100), .ZN(n4995) );
  INV_X1 U6134 ( .A(n7880), .ZN(n7713) );
  AND3_X1 U6135 ( .A1(n6266), .A2(n6265), .A3(n6264), .ZN(n7880) );
  XNOR2_X1 U6136 ( .A(n6618), .B(P2_IR_REG_26__SCAN_IN), .ZN(n6633) );
  INV_X1 U6137 ( .A(n6633), .ZN(n5156) );
  INV_X1 U6138 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6352) );
  NAND2_X1 U6139 ( .A1(n6061), .A2(n6049), .ZN(n6512) );
  NAND2_X1 U6140 ( .A1(n6063), .A2(n6062), .ZN(n10198) );
  INV_X1 U6141 ( .A(n10198), .ZN(n5242) );
  INV_X1 U6142 ( .A(n9580), .ZN(n5360) );
  AND2_X1 U6143 ( .A1(n5876), .A2(n5875), .ZN(n8899) );
  NAND2_X1 U6144 ( .A1(n5529), .A2(n8963), .ZN(n9083) );
  INV_X1 U6145 ( .A(n9909), .ZN(n5417) );
  NAND3_X1 U6146 ( .A1(n5614), .A2(n5521), .A3(n5561), .ZN(n5686) );
  AND2_X1 U6147 ( .A1(n6263), .A2(n6260), .ZN(n7745) );
  INV_X1 U6148 ( .A(n7745), .ZN(n5437) );
  AND2_X1 U6149 ( .A1(n5494), .A2(n5885), .ZN(n4996) );
  AND2_X1 U6150 ( .A1(n7187), .A2(n10002), .ZN(n4997) );
  AND2_X1 U6151 ( .A1(n10427), .A2(n8511), .ZN(n4998) );
  NAND2_X1 U6152 ( .A1(n5309), .A2(n6588), .ZN(n9534) );
  NAND2_X1 U6153 ( .A1(n5614), .A2(n5521), .ZN(n5665) );
  NAND4_X1 U6154 ( .A1(n6257), .A2(n6256), .A3(n6255), .A4(n6254), .ZN(n9391)
         );
  NOR2_X1 U6155 ( .A1(n10713), .A2(n9423), .ZN(n4999) );
  INV_X1 U6156 ( .A(n8191), .ZN(n9388) );
  AND4_X1 U6157 ( .A1(n6323), .A2(n6322), .A3(n6321), .A4(n6320), .ZN(n8191)
         );
  AND2_X1 U6158 ( .A1(n5134), .A2(n6605), .ZN(n5000) );
  OR2_X1 U6159 ( .A1(n7680), .A2(n7578), .ZN(n5001) );
  NOR2_X1 U6160 ( .A1(n7211), .A2(n7212), .ZN(n5002) );
  NAND2_X1 U6161 ( .A1(n8992), .A2(n9122), .ZN(n5003) );
  NAND2_X1 U6162 ( .A1(n6107), .A2(n10135), .ZN(n6831) );
  INV_X1 U6163 ( .A(n6831), .ZN(n6750) );
  AND2_X1 U6164 ( .A1(n9362), .A2(n6609), .ZN(n5004) );
  INV_X1 U6165 ( .A(n8908), .ZN(n10470) );
  NAND2_X1 U6166 ( .A1(n5906), .A2(n5905), .ZN(n8908) );
  NAND2_X1 U6167 ( .A1(n9011), .A2(n9564), .ZN(n9261) );
  INV_X1 U6168 ( .A(n6876), .ZN(n5349) );
  AND2_X1 U6169 ( .A1(n5414), .A2(n5002), .ZN(n5005) );
  OR2_X1 U6170 ( .A1(n4975), .A2(n5532), .ZN(n5006) );
  INV_X1 U6171 ( .A(n5216), .ZN(n5215) );
  NAND2_X1 U6172 ( .A1(n9174), .A2(n9191), .ZN(n5216) );
  AND2_X1 U6173 ( .A1(n7107), .A2(n5425), .ZN(n5007) );
  INV_X1 U6174 ( .A(n5315), .ZN(n5314) );
  AND2_X1 U6175 ( .A1(n9677), .A2(n9666), .ZN(n5008) );
  INV_X1 U6176 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10474) );
  NOR2_X1 U6177 ( .A1(n7066), .A2(n7065), .ZN(n5009) );
  NOR2_X1 U6178 ( .A1(n8572), .A2(n10036), .ZN(n5010) );
  INV_X1 U6179 ( .A(n5240), .ZN(n10176) );
  NOR2_X1 U6180 ( .A1(n10195), .A2(n5241), .ZN(n5240) );
  NOR2_X1 U6181 ( .A1(n9577), .A2(n9592), .ZN(n5011) );
  INV_X1 U6182 ( .A(n5512), .ZN(n5081) );
  AND2_X1 U6183 ( .A1(n5550), .A2(n6006), .ZN(n5512) );
  AND2_X1 U6184 ( .A1(n10324), .A2(n10031), .ZN(n5012) );
  AND2_X1 U6185 ( .A1(n5363), .A2(n9248), .ZN(n5362) );
  INV_X1 U6186 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6146) );
  AND3_X1 U6187 ( .A1(n5221), .A2(n5220), .A3(n5218), .ZN(n6616) );
  AND2_X1 U6188 ( .A1(n5410), .A2(n5411), .ZN(n5013) );
  AND2_X1 U6189 ( .A1(n8965), .A2(n9375), .ZN(n5014) );
  NAND2_X1 U6190 ( .A1(n8191), .A2(n8212), .ZN(n5015) );
  AND2_X1 U6191 ( .A1(n5105), .A2(n5414), .ZN(n5016) );
  INV_X1 U6192 ( .A(n5200), .ZN(n5199) );
  NAND2_X1 U6193 ( .A1(n9140), .A2(n6493), .ZN(n5200) );
  NOR2_X1 U6194 ( .A1(n9987), .A2(n9988), .ZN(n5017) );
  OR2_X1 U6195 ( .A1(n5012), .A2(n5504), .ZN(n5018) );
  NAND2_X1 U6196 ( .A1(n7352), .A2(n7346), .ZN(n5019) );
  AND2_X1 U6197 ( .A1(n5134), .A2(n5128), .ZN(n5020) );
  NAND2_X1 U6198 ( .A1(n10836), .A2(n10035), .ZN(n5021) );
  OR2_X1 U6199 ( .A1(n6787), .A2(n7372), .ZN(n5022) );
  OR2_X1 U6200 ( .A1(n10738), .A2(n9426), .ZN(n10758) );
  AND2_X1 U6201 ( .A1(n5747), .A2(n5732), .ZN(n5023) );
  AND2_X1 U6202 ( .A1(n9287), .A2(n9316), .ZN(n5024) );
  AND2_X1 U6203 ( .A1(n10774), .A2(n5283), .ZN(n5025) );
  INV_X1 U6204 ( .A(n5166), .ZN(n5165) );
  OAI21_X1 U6205 ( .B1(n8617), .B2(n5167), .A(n5391), .ZN(n5166) );
  AND2_X1 U6206 ( .A1(n9690), .A2(n9344), .ZN(n5026) );
  AND2_X1 U6207 ( .A1(n5108), .A2(n5110), .ZN(n5027) );
  NAND2_X1 U6208 ( .A1(n8583), .A2(n9386), .ZN(n5028) );
  INV_X1 U6209 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6195) );
  AND2_X1 U6210 ( .A1(n6619), .A2(n7355), .ZN(n7260) );
  INV_X1 U6211 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5458) );
  OAI21_X1 U6212 ( .B1(n9614), .B2(n5206), .A(n5203), .ZN(n9582) );
  AOI21_X1 U6213 ( .B1(n5157), .B2(n8624), .A(n5156), .ZN(n6621) );
  OR3_X1 U6214 ( .A1(n5544), .A2(n6260), .A3(n5291), .ZN(n5029) );
  NAND2_X1 U6215 ( .A1(n5396), .A2(n5399), .ZN(n8564) );
  NAND2_X1 U6216 ( .A1(n5072), .A2(n5506), .ZN(n8472) );
  NAND2_X1 U6217 ( .A1(n5361), .A2(n9241), .ZN(n9593) );
  NAND2_X1 U6218 ( .A1(n5505), .A2(n5914), .ZN(n10319) );
  NAND2_X1 U6219 ( .A1(n5124), .A2(n6576), .ZN(n9663) );
  NAND2_X1 U6220 ( .A1(n9129), .A2(n8947), .ZN(n9037) );
  NAND2_X1 U6221 ( .A1(n6456), .A2(n9237), .ZN(n9604) );
  NAND2_X1 U6222 ( .A1(n5493), .A2(n5494), .ZN(n8616) );
  INV_X1 U6223 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5388) );
  NAND2_X1 U6224 ( .A1(n5424), .A2(n5007), .ZN(n9879) );
  AOI21_X1 U6225 ( .B1(n8938), .B2(n5139), .A(n5137), .ZN(n5136) );
  NAND2_X1 U6226 ( .A1(n9896), .A2(n5419), .ZN(n9967) );
  NOR2_X1 U6227 ( .A1(n9489), .A2(n9753), .ZN(n5030) );
  NOR2_X1 U6228 ( .A1(n10649), .A2(n9419), .ZN(n5031) );
  NAND2_X1 U6229 ( .A1(n8634), .A2(n5238), .ZN(n5239) );
  AND2_X1 U6230 ( .A1(n9660), .A2(n6403), .ZN(n5032) );
  AND2_X1 U6231 ( .A1(n5445), .A2(n5444), .ZN(n5033) );
  NAND2_X1 U6232 ( .A1(n5097), .A2(n5427), .ZN(n9917) );
  INV_X1 U6233 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6198) );
  AND2_X1 U6234 ( .A1(n5955), .A2(n8775), .ZN(n5034) );
  AND2_X1 U6235 ( .A1(n5053), .A2(n5057), .ZN(n5035) );
  OR2_X1 U6236 ( .A1(n7971), .A2(n7184), .ZN(n10843) );
  AND2_X1 U6237 ( .A1(n10784), .A2(n7848), .ZN(n5245) );
  NAND2_X1 U6238 ( .A1(n5926), .A2(n5925), .ZN(n10324) );
  INV_X1 U6239 ( .A(n10324), .ZN(n5235) );
  AND2_X1 U6240 ( .A1(n9417), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5036) );
  NAND2_X1 U6241 ( .A1(n8103), .A2(n6884), .ZN(n8223) );
  OR2_X1 U6242 ( .A1(n6079), .A2(n5488), .ZN(n5037) );
  OAI211_X1 U6243 ( .C1(n5304), .C2(n8068), .A(n5015), .B(n5135), .ZN(n8188)
         );
  OR2_X1 U6244 ( .A1(n10657), .A2(n9403), .ZN(n5038) );
  NAND2_X1 U6245 ( .A1(n6567), .A2(n6566), .ZN(n8320) );
  NAND2_X1 U6246 ( .A1(n5090), .A2(n7017), .ZN(n8059) );
  NAND2_X1 U6247 ( .A1(n7009), .A2(n7887), .ZN(n7951) );
  AND2_X1 U6248 ( .A1(n6572), .A2(n6573), .ZN(n8529) );
  NOR2_X1 U6249 ( .A1(n9414), .A2(n9415), .ZN(n5039) );
  OR2_X1 U6250 ( .A1(n10657), .A2(n8534), .ZN(n5040) );
  INV_X1 U6251 ( .A(n6823), .ZN(n6888) );
  OR2_X1 U6252 ( .A1(n5036), .A2(n5058), .ZN(n5041) );
  XNOR2_X1 U6253 ( .A(n6238), .B(n6237), .ZN(n6600) );
  BUF_X1 U6254 ( .A(n6252), .Z(n6599) );
  NAND2_X1 U6255 ( .A1(n6138), .A2(n6137), .ZN(n10312) );
  NAND2_X1 U6256 ( .A1(n8501), .A2(n4966), .ZN(n6802) );
  NAND2_X1 U6258 ( .A1(n6554), .A2(n6553), .ZN(n7720) );
  INV_X1 U6259 ( .A(n10838), .ZN(n10425) );
  NAND2_X1 U6260 ( .A1(n7936), .A2(n10793), .ZN(n10838) );
  INV_X1 U6261 ( .A(n9144), .ZN(n5189) );
  OR2_X1 U6262 ( .A1(n5510), .A2(n10474), .ZN(n5042) );
  INV_X1 U6263 ( .A(n10576), .ZN(n5276) );
  INV_X1 U6264 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7845) );
  INV_X1 U6265 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5440) );
  AOI21_X1 U6266 ( .B1(n5128), .B2(n9682), .A(n7250), .ZN(n5126) );
  OR2_X1 U6267 ( .A1(n6606), .A2(n9682), .ZN(n5134) );
  OAI21_X1 U6268 ( .B1(n9272), .B2(n9271), .A(n9270), .ZN(n9273) );
  AND2_X1 U6269 ( .A1(n5222), .A2(n5223), .ZN(n9364) );
  OR2_X1 U6270 ( .A1(n9649), .A2(n9215), .ZN(n9219) );
  AOI21_X2 U6271 ( .B1(n5765), .B2(n5764), .A(n5763), .ZN(n5770) );
  NAND2_X1 U6272 ( .A1(n5483), .A2(n5862), .ZN(n5867) );
  NAND3_X1 U6273 ( .A1(n5293), .A2(n9638), .A3(n9224), .ZN(n5296) );
  NAND3_X1 U6274 ( .A1(n5647), .A2(n5646), .A3(n5559), .ZN(n5045) );
  INV_X1 U6275 ( .A(n5460), .ZN(n5459) );
  OAI21_X1 U6276 ( .B1(n5617), .B2(n5581), .A(n5580), .ZN(n5582) );
  NAND2_X1 U6277 ( .A1(n5751), .A2(n5750), .ZN(n5765) );
  OR2_X1 U6278 ( .A1(n5582), .A2(SI_1_), .ZN(n5583) );
  NAND3_X1 U6279 ( .A1(n5046), .A2(n9288), .A3(n5024), .ZN(n9296) );
  NAND3_X1 U6280 ( .A1(n9286), .A2(n9319), .A3(n5047), .ZN(n5046) );
  OAI21_X1 U6281 ( .B1(n5298), .B2(n5297), .A(n9268), .ZN(n9272) );
  AOI21_X1 U6282 ( .B1(n9363), .B2(n6221), .A(n5004), .ZN(n5222) );
  NOR2_X1 U6283 ( .A1(n5051), .A2(n5050), .ZN(n9420) );
  NOR2_X1 U6284 ( .A1(n10634), .A2(n5036), .ZN(n9418) );
  NAND3_X1 U6285 ( .A1(n5056), .A2(n5054), .A3(n5053), .ZN(n5052) );
  AND2_X1 U6286 ( .A1(n5067), .A2(n9435), .ZN(n9423) );
  MUX2_X1 U6287 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(P2_DATAO_REG_0__SCAN_IN), 
        .S(n5617), .Z(n5070) );
  OR2_X1 U6288 ( .A1(n5685), .A2(n5684), .ZN(n5089) );
  NAND2_X1 U6289 ( .A1(n8059), .A2(n8060), .ZN(n5423) );
  NAND2_X1 U6290 ( .A1(n7951), .A2(n7952), .ZN(n5090) );
  NAND2_X1 U6291 ( .A1(n7005), .A2(n7006), .ZN(n7886) );
  NAND3_X1 U6292 ( .A1(n5427), .A2(n10011), .A3(n5094), .ZN(n5093) );
  AOI21_X2 U6293 ( .B1(n9898), .B2(n5419), .A(n5098), .ZN(n7072) );
  NOR2_X2 U6294 ( .A1(n5686), .A2(n5233), .ZN(n5719) );
  AND2_X2 U6295 ( .A1(n5570), .A2(n5563), .ZN(n5523) );
  NAND2_X1 U6296 ( .A1(n8360), .A2(n5101), .ZN(n5104) );
  AND2_X1 U6297 ( .A1(n5399), .A2(n8358), .ZN(n5101) );
  NAND3_X1 U6298 ( .A1(n5104), .A2(n5102), .A3(n5397), .ZN(n7051) );
  NAND2_X1 U6299 ( .A1(n8357), .A2(n8359), .ZN(n8381) );
  NAND3_X1 U6300 ( .A1(n6567), .A2(n5108), .A3(n5326), .ZN(n5107) );
  NAND3_X1 U6301 ( .A1(n5107), .A2(n5028), .A3(n5106), .ZN(n6571) );
  NAND2_X1 U6302 ( .A1(n5027), .A2(n5326), .ZN(n5106) );
  INV_X1 U6303 ( .A(n8321), .ZN(n5110) );
  NAND2_X1 U6304 ( .A1(n5685), .A2(n5684), .ZN(n5700) );
  OAI21_X1 U6305 ( .B1(n5685), .B2(n5115), .A(n5113), .ZN(n5712) );
  NAND2_X1 U6306 ( .A1(n5685), .A2(n5113), .ZN(n5112) );
  OAI21_X1 U6307 ( .B1(n9611), .B2(n5121), .A(n5118), .ZN(n9587) );
  NAND2_X1 U6308 ( .A1(n9611), .A2(n5118), .ZN(n5117) );
  OAI21_X1 U6309 ( .B1(n9611), .B2(n6584), .A(n6585), .ZN(n9601) );
  NAND2_X1 U6310 ( .A1(n9663), .A2(n9664), .ZN(n6577) );
  OAI21_X1 U6311 ( .B1(n8529), .B2(n5307), .A(n5125), .ZN(n5124) );
  INV_X1 U6312 ( .A(n8180), .ZN(n8212) );
  NAND2_X1 U6313 ( .A1(n5718), .A2(n5733), .ZN(n7375) );
  INV_X1 U6314 ( .A(n5136), .ZN(n9126) );
  NAND3_X1 U6315 ( .A1(n5143), .A2(n5142), .A3(n5144), .ZN(n8991) );
  NAND2_X1 U6316 ( .A1(n9119), .A2(n5146), .ZN(n5142) );
  NAND2_X1 U6317 ( .A1(n9119), .A2(n8982), .ZN(n8995) );
  MUX2_X1 U6318 ( .A(n8979), .B(n9509), .S(n8966), .Z(n9118) );
  NAND3_X1 U6319 ( .A1(n6341), .A2(n5323), .A3(n6215), .ZN(n6635) );
  NAND2_X1 U6320 ( .A1(n9063), .A2(n5159), .ZN(n5158) );
  INV_X1 U6321 ( .A(n8614), .ZN(n5163) );
  OAI21_X1 U6322 ( .B1(n5163), .B2(n5166), .A(n5161), .ZN(n6127) );
  OAI211_X1 U6323 ( .C1(n10280), .C2(n5170), .A(n6661), .B(n5169), .ZN(n5379)
         );
  OR2_X1 U6324 ( .A1(n6828), .A2(n6131), .ZN(n5170) );
  NAND2_X1 U6325 ( .A1(n5178), .A2(n5176), .ZN(n8508) );
  AOI21_X1 U6326 ( .B1(n6893), .B2(n5179), .A(n5177), .ZN(n5176) );
  NAND3_X1 U6327 ( .A1(n5342), .A2(n5179), .A3(n5343), .ZN(n5178) );
  OAI21_X1 U6328 ( .B1(n10136), .B2(n8902), .A(n6148), .ZN(n5182) );
  NAND2_X1 U6329 ( .A1(n6136), .A2(n6831), .ZN(n5183) );
  MUX2_X1 U6330 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n4964), .Z(n5662) );
  NOR2_X4 U6331 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6242) );
  NAND2_X1 U6332 ( .A1(n9150), .A2(n9148), .ZN(n7628) );
  AND2_X2 U6333 ( .A1(n6252), .A2(n4964), .ZN(n6258) );
  OR2_X1 U6334 ( .A1(n6494), .A2(n5196), .ZN(n5193) );
  NAND2_X1 U6335 ( .A1(n5193), .A2(n5194), .ZN(n9527) );
  NAND2_X1 U6336 ( .A1(n9614), .A2(n5203), .ZN(n5202) );
  NAND2_X1 U6337 ( .A1(n5202), .A2(n5201), .ZN(n9566) );
  INV_X1 U6338 ( .A(n5362), .ZN(n5206) );
  NAND3_X1 U6339 ( .A1(n5209), .A2(n4995), .A3(n8029), .ZN(n5208) );
  NAND3_X1 U6340 ( .A1(n5208), .A2(n5207), .A3(n9197), .ZN(n8482) );
  NAND3_X1 U6341 ( .A1(n5209), .A2(n5211), .A3(n4995), .ZN(n5207) );
  NOR2_X1 U6342 ( .A1(n8321), .A2(n5213), .ZN(n5212) );
  AND2_X1 U6343 ( .A1(n4988), .A2(n5318), .ZN(n5218) );
  NOR2_X1 U6344 ( .A1(n6260), .A2(n6197), .ZN(n5219) );
  INV_X1 U6345 ( .A(n6197), .ZN(n5322) );
  NAND3_X1 U6346 ( .A1(n5221), .A2(n5220), .A3(n5217), .ZN(n6236) );
  NOR2_X2 U6347 ( .A1(n6213), .A2(n6214), .ZN(n6215) );
  NAND2_X1 U6348 ( .A1(n9659), .A2(n5228), .ZN(n5227) );
  INV_X1 U6349 ( .A(n5239), .ZN(n8906) );
  NAND3_X1 U6350 ( .A1(n10795), .A2(n5245), .A3(n7890), .ZN(n5243) );
  NAND2_X1 U6351 ( .A1(n5254), .A2(n5251), .ZN(n6751) );
  NAND2_X1 U6352 ( .A1(n5252), .A2(n4963), .ZN(n5251) );
  NAND2_X1 U6353 ( .A1(n5253), .A2(n6834), .ZN(n6747) );
  NAND2_X1 U6354 ( .A1(n6743), .A2(n6744), .ZN(n5253) );
  AND2_X2 U6355 ( .A1(n5260), .A2(n8904), .ZN(n6732) );
  NAND2_X1 U6356 ( .A1(n6671), .A2(n4963), .ZN(n5265) );
  NAND2_X1 U6357 ( .A1(n5270), .A2(n5269), .ZN(n6703) );
  OR3_X1 U6358 ( .A1(n6893), .A2(n6668), .A3(n4963), .ZN(n5270) );
  INV_X1 U6359 ( .A(n6739), .ZN(n5271) );
  INV_X1 U6360 ( .A(n6738), .ZN(n5273) );
  MUX2_X1 U6361 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n7346), .Z(n5643) );
  MUX2_X1 U6362 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n7346), .Z(n5681) );
  MUX2_X1 U6363 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n7346), .Z(n5701) );
  NAND3_X1 U6364 ( .A1(n10775), .A2(n5025), .A3(n5281), .ZN(P2_U3200) );
  INV_X1 U6365 ( .A(n5284), .ZN(n6205) );
  NAND2_X1 U6366 ( .A1(n6204), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6219) );
  INV_X1 U6367 ( .A(n5544), .ZN(n5288) );
  NAND2_X1 U6368 ( .A1(n5288), .A2(n5287), .ZN(n6382) );
  NAND2_X1 U6369 ( .A1(n9218), .A2(n9217), .ZN(n5293) );
  NOR2_X1 U6370 ( .A1(n9229), .A2(n5295), .ZN(n5294) );
  AND2_X1 U6371 ( .A1(n5300), .A2(n5299), .ZN(n5301) );
  NAND3_X1 U6372 ( .A1(n9284), .A2(n9333), .A3(n9152), .ZN(n5299) );
  NAND3_X1 U6373 ( .A1(n9153), .A2(n9333), .A3(n9269), .ZN(n5300) );
  NAND2_X1 U6374 ( .A1(n9158), .A2(n5301), .ZN(n9166) );
  NAND2_X1 U6375 ( .A1(n10299), .A2(n10300), .ZN(n10298) );
  NAND2_X1 U6376 ( .A1(n8508), .A2(n8509), .ZN(n8507) );
  NAND4_X2 U6377 ( .A1(n6196), .A2(n6324), .A3(n6313), .A4(n6302), .ZN(n6197)
         );
  OR2_X2 U6378 ( .A1(n10291), .A2(n10273), .ZN(n10261) );
  NAND2_X1 U6379 ( .A1(n9336), .A2(n5305), .ZN(n5304) );
  NAND2_X1 U6380 ( .A1(n5311), .A2(n5310), .ZN(n6563) );
  NOR2_X1 U6381 ( .A1(n6561), .A2(n5313), .ZN(n5312) );
  NOR2_X1 U6382 ( .A1(n7428), .A2(n7966), .ZN(n5315) );
  NOR2_X2 U6383 ( .A1(n5316), .A2(n5317), .ZN(n6227) );
  NAND3_X1 U6384 ( .A1(n4988), .A2(n6215), .A3(n5548), .ZN(n5316) );
  NAND2_X1 U6385 ( .A1(n9505), .A2(n8981), .ZN(n5336) );
  NAND2_X1 U6386 ( .A1(n5329), .A2(n5332), .ZN(n7234) );
  NAND2_X1 U6387 ( .A1(n9505), .A2(n5330), .ZN(n5329) );
  NAND2_X1 U6388 ( .A1(n5336), .A2(n5335), .ZN(n9495) );
  AND2_X1 U6389 ( .A1(n5336), .A2(n8978), .ZN(n9496) );
  OAI21_X1 U6390 ( .B1(n6119), .B2(n8074), .A(n8073), .ZN(n8343) );
  NAND2_X1 U6391 ( .A1(n6884), .A2(n8078), .ZN(n5338) );
  INV_X1 U6392 ( .A(n6119), .ZN(n8078) );
  NAND2_X2 U6393 ( .A1(n6242), .A2(n5339), .ZN(n6260) );
  AOI21_X1 U6394 ( .B1(n6888), .B2(n6817), .A(n5341), .ZN(n5344) );
  AND2_X1 U6395 ( .A1(n5340), .A2(n8261), .ZN(n5342) );
  OAI21_X1 U6396 ( .B1(n8103), .B2(n6823), .A(n5344), .ZN(n8262) );
  NAND2_X1 U6397 ( .A1(n8103), .A2(n5344), .ZN(n5343) );
  NAND2_X1 U6398 ( .A1(n6121), .A2(n5347), .ZN(n5346) );
  NAND3_X1 U6399 ( .A1(n6815), .A2(n5348), .A3(n5346), .ZN(n6122) );
  AND2_X1 U6401 ( .A1(n5356), .A2(n6293), .ZN(n5355) );
  NAND3_X1 U6402 ( .A1(n5364), .A2(n5366), .A3(n9241), .ZN(n5363) );
  NAND2_X1 U6403 ( .A1(n8528), .A2(n5026), .ZN(n5369) );
  NAND2_X1 U6404 ( .A1(n5369), .A2(n5370), .ZN(n9659) );
  OR2_X1 U6405 ( .A1(n10186), .A2(n5377), .ZN(n5373) );
  NAND2_X1 U6406 ( .A1(n5373), .A2(n5374), .ZN(n10137) );
  NAND2_X1 U6407 ( .A1(n9637), .A2(n5381), .ZN(n9627) );
  NAND2_X1 U6408 ( .A1(n6524), .A2(n6523), .ZN(n9307) );
  NAND3_X1 U6409 ( .A1(n5522), .A2(n5386), .A3(n5719), .ZN(n5592) );
  AND2_X1 U6410 ( .A1(n6730), .A2(n5390), .ZN(n5389) );
  NAND3_X1 U6411 ( .A1(n7239), .A2(n7230), .A3(n5393), .ZN(n9479) );
  NAND2_X1 U6412 ( .A1(n6977), .A2(n5394), .ZN(n7755) );
  NAND2_X1 U6413 ( .A1(n7760), .A2(n5394), .ZN(n7762) );
  NAND2_X1 U6414 ( .A1(n6162), .A2(n6116), .ZN(n5395) );
  NAND2_X1 U6415 ( .A1(n9945), .A2(n4994), .ZN(n5410) );
  OR2_X1 U6416 ( .A1(n9945), .A2(n7149), .ZN(n5418) );
  AND2_X2 U6417 ( .A1(n5418), .A2(n5417), .ZN(n10000) );
  INV_X1 U6418 ( .A(n5418), .ZN(n9910) );
  NAND2_X1 U6419 ( .A1(n5423), .A2(n7024), .ZN(n7031) );
  NAND2_X1 U6420 ( .A1(n5423), .A2(n5421), .ZN(n8360) );
  NAND2_X1 U6421 ( .A1(n9987), .A2(n9988), .ZN(n5425) );
  NAND2_X1 U6422 ( .A1(n10010), .A2(n10013), .ZN(n5427) );
  NAND2_X1 U6423 ( .A1(n7081), .A2(n7080), .ZN(n10011) );
  NAND4_X1 U6424 ( .A1(n5523), .A2(n5688), .A3(n5429), .A4(n5562), .ZN(n5428)
         );
  NAND3_X1 U6425 ( .A1(n7575), .A2(n7574), .A3(n5437), .ZN(n5436) );
  INV_X1 U6426 ( .A(n7680), .ZN(n5441) );
  OAI21_X1 U6427 ( .B1(n5579), .B2(n5459), .A(n5457), .ZN(n5580) );
  OAI21_X2 U6428 ( .B1(n5786), .B2(n5464), .A(n5461), .ZN(n5845) );
  NAND2_X1 U6429 ( .A1(n5935), .A2(n5474), .ZN(n5472) );
  NAND2_X1 U6430 ( .A1(n5472), .A2(n5473), .ZN(n5971) );
  NAND2_X1 U6431 ( .A1(n5847), .A2(n5484), .ZN(n5483) );
  NAND2_X1 U6432 ( .A1(n6022), .A2(n6021), .ZN(n6026) );
  NAND2_X1 U6433 ( .A1(n5733), .A2(n5023), .ZN(n5751) );
  NAND2_X1 U6434 ( .A1(n6045), .A2(n5489), .ZN(n6061) );
  NAND2_X1 U6435 ( .A1(n6045), .A2(n6044), .ZN(n6048) );
  OAI21_X2 U6436 ( .B1(n6045), .B2(n5037), .A(n5486), .ZN(n6090) );
  NAND2_X1 U6437 ( .A1(n5827), .A2(n4974), .ZN(n5493) );
  NAND2_X1 U6438 ( .A1(n8905), .A2(n5503), .ZN(n5501) );
  NAND2_X1 U6439 ( .A1(n6861), .A2(n5590), .ZN(n5576) );
  NAND2_X1 U6440 ( .A1(n6075), .A2(n5518), .ZN(n5517) );
  NAND2_X1 U6441 ( .A1(n5517), .A2(n5515), .ZN(n10142) );
  NAND2_X1 U6442 ( .A1(n5517), .A2(n6088), .ZN(n6108) );
  INV_X1 U6443 ( .A(n6074), .ZN(n5519) );
  NOR2_X2 U6444 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5521) );
  NOR2_X2 U6445 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5614) );
  NAND2_X1 U6446 ( .A1(n5136), .A2(n5531), .ZN(n5530) );
  NAND2_X1 U6447 ( .A1(n5536), .A2(n5539), .ZN(n7709) );
  NAND2_X1 U6448 ( .A1(n5535), .A2(n5537), .ZN(n5539) );
  INV_X1 U6449 ( .A(n7619), .ZN(n5535) );
  AND2_X1 U6450 ( .A1(n7710), .A2(n5538), .ZN(n5536) );
  NOR2_X1 U6451 ( .A1(n7618), .A2(n7272), .ZN(n7711) );
  INV_X1 U6452 ( .A(n7273), .ZN(n5541) );
  NAND2_X1 U6453 ( .A1(n9015), .A2(n4984), .ZN(n9063) );
  NAND2_X1 U6455 ( .A1(n8050), .A2(n4987), .ZN(n5545) );
  NAND2_X1 U6456 ( .A1(n5545), .A2(n5546), .ZN(n8418) );
  INV_X1 U6457 ( .A(n5547), .ZN(n8049) );
  INV_X1 U6458 ( .A(n9353), .ZN(n7235) );
  MUX2_X2 U6459 ( .A(n6654), .B(n5020), .S(n10851), .Z(n6655) );
  NAND2_X1 U6460 ( .A1(n5654), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5601) );
  AND2_X1 U6461 ( .A1(n6949), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6176) );
  INV_X1 U6462 ( .A(n6973), .ZN(n6976) );
  XNOR2_X1 U6463 ( .A(n6164), .B(n6163), .ZN(n6170) );
  AND2_X2 U6464 ( .A1(n8932), .A2(n5596), .ZN(n5654) );
  OR2_X1 U6465 ( .A1(n6009), .A2(n6008), .ZN(n6010) );
  NAND2_X1 U6466 ( .A1(n5654), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5602) );
  OAI21_X1 U6467 ( .B1(n9322), .B2(n9784), .A(n9357), .ZN(n9323) );
  INV_X1 U6468 ( .A(n8218), .ZN(n6150) );
  NAND2_X1 U6469 ( .A1(n10116), .A2(n8218), .ZN(n6946) );
  XNOR2_X1 U6470 ( .A(n6756), .B(n6755), .ZN(n9844) );
  NAND2_X1 U6471 ( .A1(n10142), .A2(n6109), .ZN(n10167) );
  INV_X1 U6472 ( .A(n5597), .ZN(n8932) );
  AOI21_X2 U6473 ( .B1(n5971), .B2(n5970), .A(n5969), .ZN(n5976) );
  INV_X1 U6474 ( .A(n6552), .ZN(n7633) );
  OR2_X1 U6475 ( .A1(n6252), .A2(n6245), .ZN(n6246) );
  OAI21_X1 U6476 ( .B1(n7625), .B2(n7266), .A(n7267), .ZN(n7612) );
  NAND2_X1 U6477 ( .A1(n7266), .A2(n7625), .ZN(n7267) );
  AND4_X1 U6478 ( .A1(n6431), .A2(n6430), .A3(n6429), .A4(n6428), .ZN(n9648)
         );
  OR2_X1 U6479 ( .A1(n10234), .A2(n10245), .ZN(n5550) );
  AND2_X1 U6480 ( .A1(n10028), .A2(n10138), .ZN(n5551) );
  AND3_X1 U6481 ( .A1(n6792), .A2(n6791), .A3(n6790), .ZN(n6806) );
  INV_X1 U6482 ( .A(n6806), .ZN(n10138) );
  INV_X1 U6483 ( .A(n6221), .ZN(n6609) );
  OR2_X1 U6484 ( .A1(n9391), .A2(n7713), .ZN(n5553) );
  AND2_X1 U6485 ( .A1(n8416), .A2(n8415), .ZN(n5554) );
  AND3_X1 U6486 ( .A1(n7205), .A2(n10002), .A3(n7204), .ZN(n5555) );
  AND2_X1 U6487 ( .A1(n6750), .A2(n6835), .ZN(n5556) );
  OR2_X1 U6488 ( .A1(n10564), .A2(n6601), .ZN(n10747) );
  INV_X1 U6489 ( .A(n10747), .ZN(n9468) );
  XNOR2_X1 U6490 ( .A(n6615), .B(P2_IR_REG_25__SCAN_IN), .ZN(n6632) );
  AND2_X1 U6491 ( .A1(n9433), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5557) );
  AND2_X1 U6492 ( .A1(n5680), .A2(n5663), .ZN(n5559) );
  INV_X1 U6493 ( .A(n9282), .ZN(n9489) );
  INV_X1 U6494 ( .A(n9494), .ZN(n6590) );
  AND2_X1 U6495 ( .A1(n9672), .A2(n7879), .ZN(n9692) );
  NAND2_X1 U6496 ( .A1(n7078), .A2(n7079), .ZN(n10010) );
  OR2_X1 U6497 ( .A1(n9489), .A2(n9833), .ZN(n5560) );
  INV_X1 U6498 ( .A(n9781), .ZN(n7250) );
  INV_X1 U6499 ( .A(n10851), .ZN(n7244) );
  AND2_X1 U6500 ( .A1(n9326), .A2(n6646), .ZN(n9682) );
  NAND2_X1 U6501 ( .A1(n7072), .A2(n7073), .ZN(n9858) );
  INV_X1 U6502 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6207) );
  INV_X1 U6503 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5566) );
  INV_X1 U6504 ( .A(n9382), .ZN(n8943) );
  INV_X1 U6505 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5563) );
  NOR3_X1 U6506 ( .A1(n9294), .A2(n9489), .A3(n9293), .ZN(n9295) );
  INV_X1 U6507 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6224) );
  INV_X1 U6508 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6345) );
  INV_X1 U6509 ( .A(n7783), .ZN(n9154) );
  INV_X1 U6510 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6237) );
  INV_X1 U6511 ( .A(n8920), .ZN(n6132) );
  INV_X1 U6512 ( .A(n8089), .ZN(n6815) );
  INV_X1 U6513 ( .A(n9118), .ZN(n8980) );
  NAND2_X1 U6514 ( .A1(n6468), .A2(n8857), .ZN(n6477) );
  NAND2_X1 U6515 ( .A1(n6346), .A2(n6345), .ZN(n6357) );
  NAND2_X1 U6516 ( .A1(n6558), .A2(n5553), .ZN(n6560) );
  NOR2_X1 U6517 ( .A1(n5982), .A2(n9891), .ZN(n5996) );
  AOI21_X1 U6518 ( .B1(n6804), .B2(n6802), .A(n5551), .ZN(n6798) );
  NOR2_X1 U6519 ( .A1(n5853), .A2(n7809), .ZN(n5877) );
  NOR2_X1 U6520 ( .A1(n6133), .A2(n6132), .ZN(n6134) );
  OR2_X1 U6521 ( .A1(n6769), .A2(n6768), .ZN(n6770) );
  INV_X1 U6522 ( .A(SI_19_), .ZN(n8775) );
  OR2_X1 U6523 ( .A1(n5869), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5870) );
  INV_X1 U6524 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5562) );
  NOR2_X1 U6525 ( .A1(n6318), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6335) );
  INV_X1 U6526 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6296) );
  NOR2_X1 U6527 ( .A1(n9122), .A2(n9684), .ZN(n6603) );
  NAND2_X1 U6528 ( .A1(n9703), .A2(n9521), .ZN(n8981) );
  INV_X1 U6529 ( .A(n6611), .ZN(n6612) );
  INV_X1 U6530 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6171) );
  AND2_X1 U6531 ( .A1(n5777), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5792) );
  INV_X1 U6532 ( .A(n9899), .ZN(n7055) );
  AND2_X1 U6533 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5671) );
  OR2_X1 U6534 ( .A1(n6013), .A2(n9874), .ZN(n6030) );
  INV_X1 U6535 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5834) );
  NOR2_X1 U6536 ( .A1(n6051), .A2(n9911), .ZN(n6064) );
  INV_X1 U6537 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7467) );
  INV_X1 U6538 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7809) );
  NAND2_X1 U6539 ( .A1(n10152), .A2(n10029), .ZN(n6809) );
  NAND2_X1 U6540 ( .A1(n5945), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5961) );
  INV_X1 U6541 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5907) );
  AND2_X1 U6542 ( .A1(n6670), .A2(n6695), .ZN(n6694) );
  OAI21_X1 U6543 ( .B1(n7946), .B2(n6682), .A(n6881), .ZN(n8141) );
  INV_X1 U6544 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6163) );
  OR2_X1 U6545 ( .A1(n5812), .A2(n5811), .ZN(n5815) );
  OR2_X1 U6546 ( .A1(n6537), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6545) );
  OR2_X1 U6547 ( .A1(n6307), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6318) );
  NAND2_X1 U6548 ( .A1(n7783), .A2(n6555), .ZN(n7716) );
  OR2_X1 U6549 ( .A1(n7636), .A2(n7638), .ZN(n6644) );
  AND2_X1 U6550 ( .A1(n9202), .A2(n9200), .ZN(n9343) );
  AND2_X1 U6551 ( .A1(n9162), .A2(n9173), .ZN(n9332) );
  INV_X1 U6552 ( .A(n7241), .ZN(n8540) );
  INV_X1 U6553 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6217) );
  OR2_X1 U6554 ( .A1(n5738), .A2(n7467), .ZN(n5755) );
  OR2_X1 U6555 ( .A1(n6030), .A2(n6029), .ZN(n6051) );
  OR2_X1 U6556 ( .A1(n5961), .A2(n5960), .ZN(n5982) );
  INV_X1 U6557 ( .A(n10035), .ZN(n8570) );
  INV_X1 U6558 ( .A(n5654), .ZN(n6142) );
  INV_X1 U6559 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7545) );
  INV_X1 U6560 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8455) );
  INV_X1 U6561 ( .A(n10143), .ZN(n10144) );
  AND2_X1 U6562 ( .A1(n6072), .A2(n6071), .ZN(n10208) );
  INV_X1 U6563 ( .A(n10300), .ZN(n5952) );
  AND4_X1 U6564 ( .A1(n5913), .A2(n5912), .A3(n5911), .A4(n5910), .ZN(n10314)
         );
  OR2_X1 U6565 ( .A1(n10127), .A2(n10126), .ZN(n10340) );
  INV_X1 U6566 ( .A(n10238), .ZN(n10262) );
  NAND2_X1 U6567 ( .A1(n6675), .A2(n6879), .ZN(n8089) );
  INV_X1 U6568 ( .A(n10389), .ZN(n10395) );
  AND2_X1 U6569 ( .A1(n5937), .A2(n5923), .ZN(n5936) );
  INV_X1 U6570 ( .A(n7294), .ZN(n7287) );
  INV_X1 U6571 ( .A(n9127), .ZN(n9109) );
  AND4_X1 U6572 ( .A1(n6551), .A2(n6550), .A3(n6549), .A4(n6548), .ZN(n9499)
         );
  AND4_X1 U6573 ( .A1(n6491), .A2(n6490), .A3(n6489), .A4(n6488), .ZN(n9576)
         );
  AND4_X1 U6574 ( .A1(n6381), .A2(n6380), .A3(n6379), .A4(n6378), .ZN(n9683)
         );
  INV_X1 U6575 ( .A(n10755), .ZN(n10745) );
  AND2_X1 U6576 ( .A1(P2_U3893), .A2(n6600), .ZN(n10772) );
  OR2_X1 U6577 ( .A1(n9773), .A2(n7259), .ZN(n9678) );
  INV_X1 U6578 ( .A(n9344), .ZN(n9209) );
  AND2_X1 U6579 ( .A1(n7302), .A2(n9284), .ZN(n9540) );
  AND2_X1 U6580 ( .A1(n6644), .A2(n6640), .ZN(n7640) );
  INV_X1 U6581 ( .A(n9773), .ZN(n9771) );
  NAND2_X1 U6582 ( .A1(n7878), .A2(n8540), .ZN(n9778) );
  NAND2_X1 U6583 ( .A1(n6639), .A2(n6638), .ZN(n7296) );
  NAND2_X1 U6584 ( .A1(n7051), .A2(n8563), .ZN(n9898) );
  NAND2_X1 U6585 ( .A1(n6964), .A2(n6958), .ZN(n7312) );
  AND4_X1 U6586 ( .A1(n5897), .A2(n5896), .A3(n5895), .A4(n5894), .ZN(n9935)
         );
  INV_X1 U6587 ( .A(n10122), .ZN(n10072) );
  INV_X1 U6588 ( .A(n10117), .ZN(n10076) );
  INV_X1 U6589 ( .A(n10171), .ZN(n10168) );
  INV_X1 U6590 ( .A(n10315), .ZN(n10282) );
  INV_X1 U6591 ( .A(n10264), .ZN(n10286) );
  NAND2_X1 U6592 ( .A1(n8639), .A2(n7937), .ZN(n10321) );
  OR2_X1 U6593 ( .A1(n7189), .A2(n7188), .ZN(n10326) );
  OR2_X1 U6594 ( .A1(n6802), .A2(n6150), .ZN(n10793) );
  AND2_X1 U6595 ( .A1(n6176), .A2(n7319), .ZN(n7750) );
  AND2_X1 U6596 ( .A1(n5690), .A2(n5689), .ZN(n10078) );
  AND2_X1 U6597 ( .A1(n4965), .A2(P1_U3086), .ZN(n8886) );
  OR2_X1 U6598 ( .A1(n7291), .A2(n7256), .ZN(n7566) );
  INV_X1 U6599 ( .A(n6569), .ZN(n9774) );
  NAND2_X1 U6600 ( .A1(n7287), .A2(n7286), .ZN(n9127) );
  AND4_X1 U6601 ( .A1(n9304), .A2(n6598), .A3(n6597), .A4(n6596), .ZN(n8988)
         );
  INV_X1 U6602 ( .A(n9554), .ZN(n9522) );
  OR2_X1 U6603 ( .A1(P2_U3150), .A2(n7567), .ZN(n10605) );
  AOI21_X1 U6604 ( .B1(n10770), .B2(n9468), .A(n10769), .ZN(n10775) );
  INV_X1 U6605 ( .A(n9692), .ZN(n9676) );
  NAND2_X1 U6606 ( .A1(n9781), .A2(n9771), .ZN(n9753) );
  AND3_X2 U6607 ( .A1(n6642), .A2(n7640), .A3(n6641), .ZN(n9781) );
  INV_X1 U6608 ( .A(n9014), .ZN(n9817) );
  AND2_X2 U6609 ( .A1(n6653), .A2(n7354), .ZN(n10851) );
  INV_X1 U6610 ( .A(n10721), .ZN(n9433) );
  INV_X1 U6611 ( .A(n9846), .ZN(n9855) );
  NAND2_X1 U6612 ( .A1(n7213), .A2(n4997), .ZN(n7209) );
  INV_X1 U6613 ( .A(n10372), .ZN(n9953) );
  INV_X1 U6614 ( .A(n10023), .ZN(n10009) );
  INV_X1 U6615 ( .A(n10172), .ZN(n10345) );
  INV_X1 U6616 ( .A(n7120), .ZN(n10281) );
  INV_X1 U6617 ( .A(n9904), .ZN(n10034) );
  OR2_X1 U6618 ( .A1(n7342), .A2(n7341), .ZN(n10563) );
  OR2_X1 U6619 ( .A1(n10563), .A2(n10124), .ZN(n10090) );
  OR2_X1 U6620 ( .A1(n10563), .A2(n7321), .ZN(n10117) );
  INV_X1 U6621 ( .A(n10321), .ZN(n10307) );
  INV_X1 U6622 ( .A(n8917), .ZN(n10419) );
  OR2_X1 U6623 ( .A1(n7971), .A2(n7970), .ZN(n10840) );
  INV_X1 U6624 ( .A(n10296), .ZN(n10462) );
  INV_X1 U6625 ( .A(n8442), .ZN(n8447) );
  NOR2_X2 U6626 ( .A1(n7566), .A2(P2_U3151), .ZN(P2_U3893) );
  NAND2_X1 U6627 ( .A1(n6194), .A2(n6193), .ZN(P1_U3518) );
  NAND4_X1 U6628 ( .A1(n5565), .A2(n5564), .A3(n5810), .A4(n5809), .ZN(n5569)
         );
  NAND4_X1 U6629 ( .A1(n5848), .A2(n5872), .A3(n5567), .A4(n5566), .ZN(n5568)
         );
  NOR3_X1 U6630 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .A3(
        P1_IR_REG_24__SCAN_IN), .ZN(n5571) );
  NAND2_X1 U6631 ( .A1(n5574), .A2(n6146), .ZN(n5590) );
  NAND3_X1 U6632 ( .A1(n5573), .A2(P1_IR_REG_31__SCAN_IN), .A3(n5574), .ZN(
        n5575) );
  INV_X1 U6633 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U6634 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5577) );
  XNOR2_X1 U6635 ( .A(n5578), .B(n5577), .ZN(n7349) );
  NAND2_X1 U6636 ( .A1(n5582), .A2(SI_1_), .ZN(n5615) );
  NAND2_X1 U6637 ( .A1(n5583), .A2(n5615), .ZN(n5587) );
  INV_X1 U6638 ( .A(n5587), .ZN(n5584) );
  INV_X1 U6639 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U6640 ( .A1(n5584), .A2(n5585), .ZN(n5616) );
  INV_X1 U6641 ( .A(n5585), .ZN(n5586) );
  NAND2_X1 U6642 ( .A1(n5587), .A2(n5586), .ZN(n5588) );
  NAND2_X1 U6643 ( .A1(n5616), .A2(n5588), .ZN(n7352) );
  NOR2_X2 U6644 ( .A1(n5592), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U6645 ( .A1(n5592), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5593) );
  MUX2_X1 U6646 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5593), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5595) );
  INV_X1 U6647 ( .A(n5594), .ZN(n10475) );
  NAND2_X1 U6648 ( .A1(n5631), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U6649 ( .A1(n5609), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5599) );
  AND2_X2 U6650 ( .A1(n8932), .A2(n10481), .ZN(n5652) );
  NAND4_X4 U6651 ( .A1(n5601), .A2(n5600), .A3(n5599), .A4(n5598), .ZN(n10044)
         );
  NAND2_X1 U6652 ( .A1(n5609), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5605) );
  NAND2_X1 U6653 ( .A1(n4958), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5604) );
  NAND2_X1 U6654 ( .A1(n5652), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5603) );
  NAND4_X1 U6655 ( .A1(n5605), .A2(n5604), .A3(n5603), .A4(n5602), .ZN(n6960)
         );
  INV_X1 U6656 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10557) );
  NAND2_X1 U6657 ( .A1(n4965), .A2(SI_0_), .ZN(n5607) );
  XNOR2_X1 U6658 ( .A(n5607), .B(n5606), .ZN(n10495) );
  MUX2_X1 U6659 ( .A(n10557), .B(n10495), .S(n7316), .Z(n8075) );
  INV_X1 U6660 ( .A(n8075), .ZN(n8010) );
  NAND2_X1 U6661 ( .A1(n6960), .A2(n8010), .ZN(n8074) );
  NAND2_X1 U6662 ( .A1(n6119), .A2(n8074), .ZN(n8073) );
  INV_X1 U6663 ( .A(n10044), .ZN(n8126) );
  NAND2_X1 U6664 ( .A1(n8126), .A2(n8076), .ZN(n5608) );
  NAND2_X1 U6665 ( .A1(n8073), .A2(n5608), .ZN(n8122) );
  NAND2_X1 U6666 ( .A1(n4958), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U6667 ( .A1(n5654), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5612) );
  NAND2_X1 U6668 ( .A1(n5609), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U6669 ( .A1(n5652), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5610) );
  OR2_X1 U6670 ( .A1(n5614), .A2(n10474), .ZN(n5637) );
  INV_X1 U6671 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5636) );
  XNOR2_X1 U6672 ( .A(n5637), .B(n5636), .ZN(n7367) );
  NAND2_X1 U6673 ( .A1(n5616), .A2(n5615), .ZN(n5623) );
  MUX2_X1 U6674 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5617), .Z(n5618) );
  NAND2_X1 U6675 ( .A1(n5618), .A2(SI_2_), .ZN(n5641) );
  INV_X1 U6676 ( .A(n5618), .ZN(n5620) );
  INV_X1 U6677 ( .A(SI_2_), .ZN(n5619) );
  NAND2_X1 U6678 ( .A1(n5620), .A2(n5619), .ZN(n5621) );
  NAND2_X1 U6679 ( .A1(n5641), .A2(n5621), .ZN(n5624) );
  INV_X1 U6680 ( .A(n5624), .ZN(n5622) );
  NAND2_X1 U6681 ( .A1(n5623), .A2(n5622), .ZN(n5642) );
  INV_X1 U6682 ( .A(n5623), .ZN(n5625) );
  NAND2_X1 U6683 ( .A1(n5625), .A2(n5624), .ZN(n5626) );
  AND2_X1 U6684 ( .A1(n5642), .A2(n5626), .ZN(n7350) );
  NAND2_X1 U6685 ( .A1(n6785), .A2(n7350), .ZN(n5628) );
  INV_X1 U6686 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7369) );
  OR2_X1 U6687 ( .A1(n6787), .A2(n7369), .ZN(n5627) );
  OAI211_X1 U6688 ( .C1(n7316), .C2(n7367), .A(n5628), .B(n5627), .ZN(n6945)
         );
  INV_X1 U6689 ( .A(n6945), .ZN(n5629) );
  NAND2_X1 U6690 ( .A1(n10043), .A2(n5629), .ZN(n6674) );
  NAND2_X1 U6691 ( .A1(n8122), .A2(n8128), .ZN(n8121) );
  NAND2_X1 U6692 ( .A1(n8088), .A2(n5629), .ZN(n5630) );
  NAND2_X1 U6693 ( .A1(n8121), .A2(n5630), .ZN(n8084) );
  INV_X1 U6694 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n8348) );
  NAND2_X1 U6695 ( .A1(n5609), .A2(n8348), .ZN(n5635) );
  NAND2_X1 U6696 ( .A1(n4958), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5634) );
  NAND2_X1 U6697 ( .A1(n5654), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5633) );
  NAND2_X1 U6698 ( .A1(n5652), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5632) );
  INV_X1 U6699 ( .A(n8129), .ZN(n10042) );
  NAND2_X1 U6700 ( .A1(n5637), .A2(n5636), .ZN(n5638) );
  NAND2_X1 U6701 ( .A1(n5638), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5640) );
  INV_X1 U6702 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5639) );
  XNOR2_X1 U6703 ( .A(n5640), .B(n5639), .ZN(n10061) );
  NAND2_X1 U6704 ( .A1(n5642), .A2(n5641), .ZN(n5647) );
  NAND2_X1 U6705 ( .A1(n5643), .A2(SI_3_), .ZN(n5660) );
  INV_X1 U6706 ( .A(n5643), .ZN(n5644) );
  INV_X1 U6707 ( .A(SI_3_), .ZN(n8810) );
  NAND2_X1 U6708 ( .A1(n5644), .A2(n8810), .ZN(n5645) );
  OR2_X1 U6709 ( .A1(n5647), .A2(n5646), .ZN(n5648) );
  AND2_X1 U6710 ( .A1(n5661), .A2(n5648), .ZN(n6259) );
  INV_X1 U6711 ( .A(n6259), .ZN(n7365) );
  OR2_X1 U6712 ( .A1(n5659), .A2(n7365), .ZN(n5650) );
  INV_X1 U6713 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7366) );
  NAND2_X1 U6714 ( .A1(n10042), .A2(n7848), .ZN(n6675) );
  NAND2_X1 U6715 ( .A1(n8129), .A2(n8347), .ZN(n6879) );
  NAND2_X1 U6716 ( .A1(n8084), .A2(n8089), .ZN(n8083) );
  NAND2_X1 U6717 ( .A1(n8129), .A2(n7848), .ZN(n5651) );
  NAND2_X1 U6718 ( .A1(n8083), .A2(n5651), .ZN(n7939) );
  NAND2_X1 U6719 ( .A1(n5652), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5658) );
  NAND2_X1 U6720 ( .A1(n4958), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5657) );
  INV_X1 U6721 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5653) );
  XNOR2_X1 U6722 ( .A(n5653), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n7942) );
  NAND2_X1 U6723 ( .A1(n5609), .A2(n7942), .ZN(n5656) );
  NAND2_X1 U6724 ( .A1(n5654), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5655) );
  NAND4_X1 U6725 ( .A1(n5658), .A2(n5657), .A3(n5656), .A4(n5655), .ZN(n10041)
         );
  NAND2_X1 U6726 ( .A1(n5662), .A2(SI_4_), .ZN(n5680) );
  INV_X1 U6727 ( .A(SI_4_), .ZN(n8805) );
  XNOR2_X1 U6728 ( .A(n5679), .B(n5559), .ZN(n7373) );
  OR2_X1 U6729 ( .A1(n5659), .A2(n7373), .ZN(n5669) );
  INV_X1 U6730 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n5664) );
  OR2_X1 U6731 ( .A1(n6787), .A2(n5664), .ZN(n5668) );
  NAND2_X1 U6732 ( .A1(n5665), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5666) );
  XNOR2_X1 U6733 ( .A(n5666), .B(P1_IR_REG_4__SCAN_IN), .ZN(n7433) );
  NAND2_X1 U6734 ( .A1(n5941), .A2(n7433), .ZN(n5667) );
  NOR2_X1 U6735 ( .A1(n10041), .A2(n10784), .ZN(n6682) );
  INV_X1 U6736 ( .A(n6682), .ZN(n6676) );
  NAND2_X1 U6737 ( .A1(n10041), .A2(n10784), .ZN(n6881) );
  NAND2_X1 U6738 ( .A1(n6676), .A2(n6881), .ZN(n7945) );
  INV_X1 U6739 ( .A(n10041), .ZN(n8139) );
  NAND2_X1 U6740 ( .A1(n8139), .A2(n10784), .ZN(n5670) );
  NAND2_X1 U6741 ( .A1(n4958), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U6742 ( .A1(n5654), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5677) );
  NAND2_X1 U6743 ( .A1(n5671), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5693) );
  INV_X1 U6744 ( .A(n5671), .ZN(n5673) );
  INV_X1 U6745 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5672) );
  NAND2_X1 U6746 ( .A1(n5673), .A2(n5672), .ZN(n5674) );
  AND2_X1 U6747 ( .A1(n5693), .A2(n5674), .ZN(n8162) );
  NAND2_X1 U6748 ( .A1(n5609), .A2(n8162), .ZN(n5676) );
  NAND2_X1 U6749 ( .A1(n5652), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5675) );
  INV_X1 U6750 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7372) );
  NAND2_X1 U6751 ( .A1(n5681), .A2(SI_5_), .ZN(n5699) );
  INV_X1 U6752 ( .A(n5681), .ZN(n5682) );
  INV_X1 U6753 ( .A(SI_5_), .ZN(n8802) );
  NAND2_X1 U6754 ( .A1(n5682), .A2(n8802), .ZN(n5683) );
  AND2_X1 U6755 ( .A1(n5699), .A2(n5683), .ZN(n5684) );
  NAND2_X1 U6756 ( .A1(n5686), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5687) );
  MUX2_X1 U6757 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5687), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5690) );
  INV_X1 U6758 ( .A(n5688), .ZN(n5689) );
  NAND2_X1 U6759 ( .A1(n5941), .A2(n10078), .ZN(n5691) );
  NAND2_X1 U6760 ( .A1(n8107), .A2(n8172), .ZN(n6683) );
  INV_X1 U6761 ( .A(n8107), .ZN(n10040) );
  INV_X1 U6762 ( .A(n8172), .ZN(n7890) );
  NAND2_X1 U6763 ( .A1(n10040), .A2(n7890), .ZN(n6882) );
  NAND2_X1 U6764 ( .A1(n8107), .A2(n7890), .ZN(n5692) );
  NAND2_X1 U6765 ( .A1(n4958), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5698) );
  NAND2_X1 U6766 ( .A1(n5652), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5697) );
  NOR2_X1 U6767 ( .A1(n5693), .A2(n7449), .ZN(n5723) );
  INV_X1 U6768 ( .A(n5723), .ZN(n5725) );
  NAND2_X1 U6769 ( .A1(n5693), .A2(n7449), .ZN(n5694) );
  AND2_X1 U6770 ( .A1(n5725), .A2(n5694), .ZN(n8113) );
  NAND2_X1 U6771 ( .A1(n5609), .A2(n8113), .ZN(n5696) );
  NAND2_X1 U6772 ( .A1(n5654), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5695) );
  NAND2_X1 U6773 ( .A1(n5701), .A2(SI_6_), .ZN(n5711) );
  INV_X1 U6774 ( .A(n5701), .ZN(n5702) );
  INV_X1 U6775 ( .A(SI_6_), .ZN(n8806) );
  NAND2_X1 U6776 ( .A1(n5702), .A2(n8806), .ZN(n5703) );
  AND2_X1 U6777 ( .A1(n5711), .A2(n5703), .ZN(n5704) );
  OR2_X1 U6778 ( .A1(n5705), .A2(n5704), .ZN(n5706) );
  NAND2_X1 U6779 ( .A1(n5712), .A2(n5706), .ZN(n7363) );
  OR2_X1 U6780 ( .A1(n7363), .A2(n5659), .ZN(n5709) );
  OR2_X1 U6781 ( .A1(n5688), .A2(n10474), .ZN(n5707) );
  XNOR2_X1 U6782 ( .A(n5707), .B(P1_IR_REG_6__SCAN_IN), .ZN(n7461) );
  AOI22_X1 U6783 ( .A1(n5942), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5941), .B2(
        n7461), .ZN(n5708) );
  NAND2_X1 U6784 ( .A1(n5709), .A2(n5708), .ZN(n8114) );
  NAND2_X1 U6785 ( .A1(n8243), .A2(n8114), .ZN(n6884) );
  INV_X1 U6786 ( .A(n8114), .ZN(n10795) );
  INV_X1 U6787 ( .A(n8243), .ZN(n10039) );
  AND2_X1 U6788 ( .A1(n10795), .A2(n10039), .ZN(n8245) );
  INV_X1 U6789 ( .A(n8245), .ZN(n8224) );
  INV_X1 U6790 ( .A(n8102), .ZN(n8105) );
  NAND2_X1 U6791 ( .A1(n8106), .A2(n8105), .ZN(n8104) );
  NAND2_X1 U6792 ( .A1(n8243), .A2(n10795), .ZN(n5710) );
  NAND2_X1 U6793 ( .A1(n8104), .A2(n5710), .ZN(n8242) );
  MUX2_X1 U6794 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4965), .Z(n5713) );
  NAND2_X1 U6795 ( .A1(n5713), .A2(SI_7_), .ZN(n5732) );
  INV_X1 U6796 ( .A(n5713), .ZN(n5714) );
  INV_X1 U6797 ( .A(SI_7_), .ZN(n8803) );
  NAND2_X1 U6798 ( .A1(n5714), .A2(n8803), .ZN(n5715) );
  AND2_X1 U6799 ( .A1(n5732), .A2(n5715), .ZN(n5716) );
  OR2_X1 U6800 ( .A1(n5717), .A2(n5716), .ZN(n5718) );
  OR2_X1 U6801 ( .A1(n7375), .A2(n5659), .ZN(n5722) );
  OR2_X1 U6802 ( .A1(n5719), .A2(n10474), .ZN(n5720) );
  XNOR2_X1 U6803 ( .A(n5720), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7460) );
  AOI22_X1 U6804 ( .A1(n5942), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5941), .B2(
        n7460), .ZN(n5721) );
  NAND2_X1 U6805 ( .A1(n5652), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5730) );
  NAND2_X1 U6806 ( .A1(n4958), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5729) );
  NAND2_X1 U6807 ( .A1(n5723), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5738) );
  INV_X1 U6808 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5724) );
  NAND2_X1 U6809 ( .A1(n5725), .A2(n5724), .ZN(n5726) );
  AND2_X1 U6810 ( .A1(n5738), .A2(n5726), .ZN(n8368) );
  NAND2_X1 U6811 ( .A1(n5609), .A2(n8368), .ZN(n5728) );
  NAND2_X1 U6812 ( .A1(n5654), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5727) );
  NAND4_X1 U6813 ( .A1(n5730), .A2(n5729), .A3(n5728), .A4(n5727), .ZN(n10038)
         );
  AND2_X1 U6814 ( .A1(n8370), .A2(n10038), .ZN(n6688) );
  INV_X1 U6815 ( .A(n6688), .ZN(n6691) );
  INV_X1 U6816 ( .A(n8370), .ZN(n8253) );
  NAND2_X1 U6817 ( .A1(n8253), .A2(n8229), .ZN(n8226) );
  NAND2_X1 U6818 ( .A1(n8242), .A2(n8244), .ZN(n8241) );
  NAND2_X1 U6819 ( .A1(n8370), .A2(n8229), .ZN(n5731) );
  NAND2_X1 U6820 ( .A1(n8241), .A2(n5731), .ZN(n8232) );
  MUX2_X1 U6821 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n4965), .Z(n5748) );
  XNOR2_X1 U6822 ( .A(n5748), .B(SI_8_), .ZN(n5746) );
  XNOR2_X1 U6823 ( .A(n5745), .B(n5746), .ZN(n7377) );
  NAND2_X1 U6824 ( .A1(n7377), .A2(n6785), .ZN(n5737) );
  NAND2_X1 U6825 ( .A1(n5734), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5735) );
  XNOR2_X1 U6826 ( .A(n5735), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7492) );
  AOI22_X1 U6827 ( .A1(n5942), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5941), .B2(
        n7492), .ZN(n5736) );
  NAND2_X1 U6828 ( .A1(n5737), .A2(n5736), .ZN(n8234) );
  NAND2_X1 U6829 ( .A1(n4958), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5743) );
  NAND2_X1 U6830 ( .A1(n5652), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5742) );
  NAND2_X1 U6831 ( .A1(n5738), .A2(n7467), .ZN(n5739) );
  AND2_X1 U6832 ( .A1(n5755), .A2(n5739), .ZN(n8365) );
  NAND2_X1 U6833 ( .A1(n5609), .A2(n8365), .ZN(n5741) );
  NAND2_X1 U6834 ( .A1(n5654), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5740) );
  OR2_X1 U6835 ( .A1(n8234), .A2(n8385), .ZN(n6670) );
  NAND2_X1 U6836 ( .A1(n8234), .A2(n8385), .ZN(n6695) );
  NAND2_X1 U6837 ( .A1(n8232), .A2(n8231), .ZN(n8230) );
  INV_X1 U6838 ( .A(n8385), .ZN(n8283) );
  OR2_X1 U6839 ( .A1(n8234), .A2(n8283), .ZN(n5744) );
  NAND2_X1 U6840 ( .A1(n8230), .A2(n5744), .ZN(n8287) );
  INV_X1 U6841 ( .A(n5746), .ZN(n5747) );
  INV_X1 U6842 ( .A(n5748), .ZN(n5749) );
  INV_X1 U6843 ( .A(SI_8_), .ZN(n8689) );
  NAND2_X1 U6844 ( .A1(n5749), .A2(n8689), .ZN(n5750) );
  MUX2_X1 U6845 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n4964), .Z(n5762) );
  INV_X1 U6846 ( .A(SI_9_), .ZN(n5752) );
  XNOR2_X1 U6847 ( .A(n5762), .B(n5752), .ZN(n5764) );
  OR2_X1 U6848 ( .A1(n5734), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5812) );
  NAND2_X1 U6849 ( .A1(n5812), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5774) );
  XNOR2_X1 U6850 ( .A(n5774), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7500) );
  AOI22_X1 U6851 ( .A1(n5942), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5941), .B2(
        n7500), .ZN(n5753) );
  NAND2_X1 U6852 ( .A1(n4958), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5760) );
  NAND2_X1 U6853 ( .A1(n5652), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5759) );
  INV_X1 U6854 ( .A(n5777), .ZN(n5778) );
  NAND2_X1 U6855 ( .A1(n5755), .A2(n5754), .ZN(n5756) );
  AND2_X1 U6856 ( .A1(n5778), .A2(n5756), .ZN(n8388) );
  NAND2_X1 U6857 ( .A1(n5609), .A2(n8388), .ZN(n5758) );
  NAND2_X1 U6858 ( .A1(n5654), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5757) );
  NAND2_X1 U6859 ( .A1(n8288), .A2(n8494), .ZN(n6819) );
  INV_X1 U6860 ( .A(n8281), .ZN(n8286) );
  NAND2_X1 U6861 ( .A1(n8287), .A2(n8286), .ZN(n8285) );
  INV_X1 U6862 ( .A(n8494), .ZN(n7600) );
  OR2_X1 U6863 ( .A1(n8288), .A2(n7600), .ZN(n5761) );
  NOR2_X1 U6864 ( .A1(n5762), .A2(SI_9_), .ZN(n5763) );
  MUX2_X1 U6865 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n4965), .Z(n5766) );
  NAND2_X1 U6866 ( .A1(n5766), .A2(SI_10_), .ZN(n5785) );
  INV_X1 U6867 ( .A(n5766), .ZN(n5767) );
  INV_X1 U6868 ( .A(SI_10_), .ZN(n8754) );
  NAND2_X1 U6869 ( .A1(n5767), .A2(n8754), .ZN(n5768) );
  NAND2_X1 U6870 ( .A1(n5785), .A2(n5768), .ZN(n5771) );
  INV_X1 U6871 ( .A(n5771), .ZN(n5769) );
  INV_X1 U6872 ( .A(n5770), .ZN(n5772) );
  NAND2_X1 U6873 ( .A1(n5772), .A2(n5771), .ZN(n5773) );
  NAND2_X1 U6874 ( .A1(n5774), .A2(n5809), .ZN(n5775) );
  NAND2_X1 U6875 ( .A1(n5775), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5787) );
  XNOR2_X1 U6876 ( .A(n5787), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7531) );
  AOI22_X1 U6877 ( .A1(n5942), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5941), .B2(
        n7531), .ZN(n5776) );
  NAND2_X1 U6878 ( .A1(n5652), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5783) );
  NAND2_X1 U6879 ( .A1(n4958), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5782) );
  INV_X1 U6880 ( .A(n5792), .ZN(n5794) );
  INV_X1 U6881 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7522) );
  NAND2_X1 U6882 ( .A1(n5778), .A2(n7522), .ZN(n5779) );
  AND2_X1 U6883 ( .A1(n5794), .A2(n5779), .ZN(n8497) );
  NAND2_X1 U6884 ( .A1(n5609), .A2(n8497), .ZN(n5781) );
  NAND2_X1 U6885 ( .A1(n5654), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5780) );
  OR2_X1 U6886 ( .A1(n8269), .A2(n8431), .ZN(n6889) );
  NAND2_X1 U6887 ( .A1(n8269), .A2(n8431), .ZN(n8391) );
  INV_X1 U6888 ( .A(n8261), .ZN(n8267) );
  INV_X1 U6889 ( .A(n8431), .ZN(n10037) );
  OR2_X1 U6890 ( .A1(n8269), .A2(n10037), .ZN(n5784) );
  MUX2_X1 U6891 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n4965), .Z(n5801) );
  XNOR2_X1 U6892 ( .A(n5801), .B(SI_11_), .ZN(n5802) );
  XNOR2_X1 U6893 ( .A(n5803), .B(n5802), .ZN(n8887) );
  NAND2_X1 U6894 ( .A1(n8887), .A2(n6785), .ZN(n5791) );
  NAND2_X1 U6895 ( .A1(n5787), .A2(n5810), .ZN(n5788) );
  NAND2_X1 U6896 ( .A1(n5788), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5789) );
  XNOR2_X1 U6897 ( .A(n5789), .B(P1_IR_REG_11__SCAN_IN), .ZN(n8885) );
  AOI22_X1 U6898 ( .A1(n5942), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5941), .B2(
        n8885), .ZN(n5790) );
  NAND2_X1 U6899 ( .A1(n5652), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5799) );
  NAND2_X1 U6900 ( .A1(n4958), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5798) );
  NAND2_X1 U6901 ( .A1(n5792), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5819) );
  INV_X1 U6902 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5793) );
  NAND2_X1 U6903 ( .A1(n5794), .A2(n5793), .ZN(n5795) );
  AND2_X1 U6904 ( .A1(n5819), .A2(n5795), .ZN(n8567) );
  NAND2_X1 U6905 ( .A1(n5609), .A2(n8567), .ZN(n5797) );
  NAND2_X1 U6906 ( .A1(n5654), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5796) );
  NAND2_X1 U6907 ( .A1(n8572), .A2(n10036), .ZN(n5800) );
  MUX2_X1 U6908 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n4965), .Z(n5804) );
  NAND2_X1 U6909 ( .A1(n5804), .A2(SI_12_), .ZN(n5828) );
  OAI21_X1 U6910 ( .B1(n5804), .B2(SI_12_), .A(n5828), .ZN(n5805) );
  NAND2_X1 U6911 ( .A1(n5806), .A2(n5805), .ZN(n5807) );
  NAND2_X1 U6912 ( .A1(n5807), .A2(n5829), .ZN(n7432) );
  OR2_X1 U6913 ( .A1(n7432), .A2(n5659), .ZN(n5818) );
  INV_X1 U6914 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5808) );
  NAND3_X1 U6915 ( .A1(n5810), .A2(n5809), .A3(n5808), .ZN(n5811) );
  NAND2_X1 U6916 ( .A1(n5815), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5813) );
  MUX2_X1 U6917 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5813), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n5814) );
  INV_X1 U6918 ( .A(n5814), .ZN(n5816) );
  NOR2_X1 U6919 ( .A1(n5816), .A2(n5849), .ZN(n7700) );
  AOI22_X1 U6920 ( .A1(n5942), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5941), .B2(
        n7700), .ZN(n5817) );
  NAND2_X1 U6921 ( .A1(n4958), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5824) );
  NAND2_X1 U6922 ( .A1(n5652), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5823) );
  NAND2_X1 U6923 ( .A1(n5819), .A2(n7545), .ZN(n5820) );
  AND2_X1 U6924 ( .A1(n5835), .A2(n5820), .ZN(n9901) );
  NAND2_X1 U6925 ( .A1(n5609), .A2(n9901), .ZN(n5822) );
  NAND2_X1 U6926 ( .A1(n5654), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5821) );
  NAND4_X1 U6927 ( .A1(n5824), .A2(n5823), .A3(n5822), .A4(n5821), .ZN(n10035)
         );
  OR2_X1 U6928 ( .A1(n10836), .A2(n8570), .ZN(n5825) );
  NAND2_X1 U6929 ( .A1(n10836), .A2(n8570), .ZN(n5826) );
  MUX2_X1 U6930 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n4965), .Z(n5830) );
  NAND2_X1 U6931 ( .A1(n5830), .A2(SI_13_), .ZN(n5846) );
  OAI21_X1 U6932 ( .B1(n5830), .B2(SI_13_), .A(n5846), .ZN(n5843) );
  XNOR2_X1 U6933 ( .A(n5845), .B(n5843), .ZN(n7515) );
  NAND2_X1 U6934 ( .A1(n7515), .A2(n6785), .ZN(n5833) );
  OR2_X1 U6935 ( .A1(n5849), .A2(n10474), .ZN(n5831) );
  XNOR2_X1 U6936 ( .A(n5831), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7801) );
  AOI22_X1 U6937 ( .A1(n5942), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5941), .B2(
        n7801), .ZN(n5832) );
  NAND2_X1 U6938 ( .A1(n5652), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5840) );
  NAND2_X1 U6939 ( .A1(n5631), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U6940 ( .A1(n5835), .A2(n5834), .ZN(n5836) );
  AND2_X1 U6941 ( .A1(n5853), .A2(n5836), .ZN(n9972) );
  NAND2_X1 U6942 ( .A1(n5609), .A2(n9972), .ZN(n5838) );
  NAND2_X1 U6943 ( .A1(n5654), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5837) );
  NOR2_X1 U6944 ( .A1(n8516), .A2(n10034), .ZN(n5842) );
  NAND2_X1 U6945 ( .A1(n8516), .A2(n10034), .ZN(n5841) );
  INV_X1 U6946 ( .A(n5843), .ZN(n5844) );
  MUX2_X1 U6947 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4965), .Z(n5859) );
  XNOR2_X1 U6948 ( .A(n5859), .B(SI_14_), .ZN(n5863) );
  XNOR2_X1 U6949 ( .A(n5864), .B(n5863), .ZN(n7533) );
  NAND2_X1 U6950 ( .A1(n7533), .A2(n6785), .ZN(n5852) );
  NAND2_X1 U6951 ( .A1(n5849), .A2(n5848), .ZN(n5869) );
  NAND2_X1 U6952 ( .A1(n5869), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5850) );
  XNOR2_X1 U6953 ( .A(n5850), .B(P1_IR_REG_14__SCAN_IN), .ZN(n8146) );
  AOI22_X1 U6954 ( .A1(n5942), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5941), .B2(
        n8146), .ZN(n5851) );
  NAND2_X1 U6955 ( .A1(n5652), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5858) );
  NAND2_X1 U6956 ( .A1(n4958), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5857) );
  INV_X1 U6957 ( .A(n5877), .ZN(n5879) );
  NAND2_X1 U6958 ( .A1(n5853), .A2(n7809), .ZN(n5854) );
  AND2_X1 U6959 ( .A1(n5879), .A2(n5854), .ZN(n9863) );
  NAND2_X1 U6960 ( .A1(n5609), .A2(n9863), .ZN(n5856) );
  NAND2_X1 U6961 ( .A1(n5654), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5855) );
  NAND2_X1 U6962 ( .A1(n10427), .A2(n10021), .ZN(n6708) );
  NAND2_X1 U6963 ( .A1(n6898), .A2(n6708), .ZN(n8628) );
  INV_X1 U6964 ( .A(n10021), .ZN(n8511) );
  INV_X1 U6965 ( .A(n5859), .ZN(n5861) );
  INV_X1 U6966 ( .A(SI_14_), .ZN(n5860) );
  NAND2_X1 U6967 ( .A1(n5861), .A2(n5860), .ZN(n5862) );
  MUX2_X1 U6968 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n4964), .Z(n5865) );
  NAND2_X1 U6969 ( .A1(n5865), .A2(SI_15_), .ZN(n5886) );
  OAI21_X1 U6970 ( .B1(n5865), .B2(SI_15_), .A(n5886), .ZN(n5866) );
  NAND2_X1 U6971 ( .A1(n5867), .A2(n5866), .ZN(n5868) );
  NAND2_X1 U6972 ( .A1(n5887), .A2(n5868), .ZN(n7609) );
  OR2_X1 U6973 ( .A1(n7609), .A2(n5659), .ZN(n5876) );
  NAND2_X1 U6974 ( .A1(n5870), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5873) );
  INV_X1 U6975 ( .A(n5873), .ZN(n5871) );
  NAND2_X1 U6976 ( .A1(n5871), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U6977 ( .A1(n5873), .A2(n5872), .ZN(n5888) );
  AND2_X1 U6978 ( .A1(n5874), .A2(n5888), .ZN(n8442) );
  AOI22_X1 U6979 ( .A1(n5942), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8442), .B2(
        n5941), .ZN(n5875) );
  NAND2_X1 U6980 ( .A1(n5631), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5884) );
  NAND2_X1 U6981 ( .A1(n5652), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5883) );
  NAND2_X1 U6982 ( .A1(n5877), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5892) );
  INV_X1 U6983 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U6984 ( .A1(n5879), .A2(n5878), .ZN(n5880) );
  AND2_X1 U6985 ( .A1(n5892), .A2(n5880), .ZN(n10014) );
  NAND2_X1 U6986 ( .A1(n5609), .A2(n10014), .ZN(n5882) );
  NAND2_X1 U6987 ( .A1(n5654), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5881) );
  NAND4_X1 U6988 ( .A1(n5884), .A2(n5883), .A3(n5882), .A4(n5881), .ZN(n10033)
         );
  NAND2_X1 U6989 ( .A1(n8899), .A2(n10033), .ZN(n6902) );
  INV_X1 U6990 ( .A(n8899), .ZN(n10024) );
  NAND2_X1 U6991 ( .A1(n10024), .A2(n9925), .ZN(n6709) );
  INV_X1 U6992 ( .A(n8617), .ZN(n5885) );
  MUX2_X1 U6993 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n4965), .Z(n5899) );
  XNOR2_X1 U6994 ( .A(n5899), .B(SI_16_), .ZN(n5902) );
  XNOR2_X1 U6995 ( .A(n5903), .B(n5902), .ZN(n7726) );
  NAND2_X1 U6996 ( .A1(n7726), .A2(n6785), .ZN(n5891) );
  NAND2_X1 U6997 ( .A1(n5888), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5889) );
  XNOR2_X1 U6998 ( .A(n5889), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8555) );
  AOI22_X1 U6999 ( .A1(n8555), .A2(n5941), .B1(n5942), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U7000 ( .A1(n4958), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5897) );
  NAND2_X1 U7001 ( .A1(n5654), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U7002 ( .A1(n5892), .A2(n8455), .ZN(n5893) );
  AND2_X1 U7003 ( .A1(n5908), .A2(n5893), .ZN(n9921) );
  NAND2_X1 U7004 ( .A1(n5609), .A2(n9921), .ZN(n5895) );
  NAND2_X1 U7005 ( .A1(n5652), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5894) );
  OR2_X1 U7006 ( .A1(n10422), .A2(n9935), .ZN(n6907) );
  NAND2_X1 U7007 ( .A1(n10422), .A2(n9935), .ZN(n6905) );
  NAND2_X1 U7008 ( .A1(n6907), .A2(n6905), .ZN(n8648) );
  INV_X1 U7009 ( .A(n9935), .ZN(n10032) );
  NAND2_X1 U7010 ( .A1(n10422), .A2(n10032), .ZN(n5898) );
  NAND2_X1 U7011 ( .A1(n8643), .A2(n5898), .ZN(n8905) );
  INV_X1 U7012 ( .A(n5899), .ZN(n5900) );
  NAND2_X1 U7013 ( .A1(n5900), .A2(n8788), .ZN(n5901) );
  OAI21_X1 U7014 ( .B1(n5903), .B2(n5902), .A(n5901), .ZN(n5916) );
  MUX2_X1 U7015 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n4965), .Z(n5917) );
  XNOR2_X1 U7016 ( .A(n5917), .B(n8784), .ZN(n5915) );
  XNOR2_X1 U7017 ( .A(n5916), .B(n5915), .ZN(n7792) );
  NAND2_X1 U7018 ( .A1(n7792), .A2(n6785), .ZN(n5906) );
  NAND2_X1 U7019 ( .A1(n5924), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5904) );
  XNOR2_X1 U7020 ( .A(n5904), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10096) );
  AOI22_X1 U7021 ( .A1(n5942), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5941), .B2(
        n10096), .ZN(n5905) );
  NAND2_X1 U7022 ( .A1(n4958), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U7023 ( .A1(n5652), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5912) );
  INV_X1 U7024 ( .A(n5927), .ZN(n5929) );
  NAND2_X1 U7025 ( .A1(n5908), .A2(n5907), .ZN(n5909) );
  AND2_X1 U7026 ( .A1(n5929), .A2(n5909), .ZN(n9938) );
  NAND2_X1 U7027 ( .A1(n5609), .A2(n9938), .ZN(n5911) );
  NAND2_X1 U7028 ( .A1(n5654), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5910) );
  OR2_X1 U7029 ( .A1(n8908), .A2(n10314), .ZN(n10308) );
  AND2_X1 U7030 ( .A1(n8908), .A2(n10314), .ZN(n6126) );
  INV_X1 U7031 ( .A(n6126), .ZN(n6725) );
  NAND2_X1 U7032 ( .A1(n10308), .A2(n6725), .ZN(n8900) );
  INV_X1 U7033 ( .A(n10314), .ZN(n9993) );
  NAND2_X1 U7034 ( .A1(n8908), .A2(n9993), .ZN(n5914) );
  NAND2_X1 U7035 ( .A1(n5916), .A2(n5915), .ZN(n5920) );
  INV_X1 U7036 ( .A(n5917), .ZN(n5918) );
  NAND2_X1 U7037 ( .A1(n5918), .A2(n8784), .ZN(n5919) );
  NAND2_X1 U7038 ( .A1(n5920), .A2(n5919), .ZN(n5935) );
  MUX2_X1 U7039 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4965), .Z(n5921) );
  INV_X1 U7040 ( .A(n5921), .ZN(n5922) );
  NAND2_X1 U7041 ( .A1(n5922), .A2(n8777), .ZN(n5923) );
  XNOR2_X1 U7042 ( .A(n5935), .B(n5936), .ZN(n7927) );
  NAND2_X1 U7043 ( .A1(n7927), .A2(n6785), .ZN(n5926) );
  XNOR2_X1 U7044 ( .A(n6113), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10111) );
  AOI22_X1 U7045 ( .A1(n5942), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5941), .B2(
        n10111), .ZN(n5925) );
  INV_X1 U7046 ( .A(n5945), .ZN(n5947) );
  INV_X1 U7047 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U7048 ( .A1(n5929), .A2(n5928), .ZN(n5930) );
  NAND2_X1 U7049 ( .A1(n5947), .A2(n5930), .ZN(n10327) );
  INV_X1 U7050 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10412) );
  OAI22_X1 U7051 ( .A1(n10327), .A2(n6145), .B1(n6142), .B2(n10412), .ZN(n5934) );
  NAND2_X1 U7052 ( .A1(n5652), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5932) );
  NAND2_X1 U7053 ( .A1(n4958), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U7054 ( .A1(n5932), .A2(n5931), .ZN(n5933) );
  MUX2_X1 U7055 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n4965), .Z(n5954) );
  XNOR2_X1 U7056 ( .A(n5954), .B(SI_19_), .ZN(n5956) );
  XNOR2_X1 U7057 ( .A(n5957), .B(n5956), .ZN(n7974) );
  NAND2_X1 U7058 ( .A1(n7974), .A2(n6785), .ZN(n5944) );
  INV_X1 U7059 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5938) );
  NAND2_X1 U7060 ( .A1(n6113), .A2(n5938), .ZN(n5939) );
  XNOR2_X1 U7061 ( .A(n5940), .B(P1_IR_REG_19__SCAN_IN), .ZN(n6115) );
  AOI22_X1 U7062 ( .A1(n5942), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5941), .B2(
        n4966), .ZN(n5943) );
  INV_X1 U7063 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U7064 ( .A1(n5947), .A2(n5946), .ZN(n5948) );
  NAND2_X1 U7065 ( .A1(n5961), .A2(n5948), .ZN(n10290) );
  OR2_X1 U7066 ( .A1(n10290), .A2(n6145), .ZN(n5951) );
  AOI22_X1 U7067 ( .A1(n5631), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n5652), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n5950) );
  NAND2_X1 U7068 ( .A1(n5654), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5949) );
  OR2_X1 U7069 ( .A1(n10296), .A2(n10396), .ZN(n6728) );
  NAND2_X1 U7070 ( .A1(n10296), .A2(n10396), .ZN(n6910) );
  INV_X1 U7071 ( .A(n10396), .ZN(n7604) );
  NAND2_X1 U7072 ( .A1(n10296), .A2(n7604), .ZN(n5953) );
  INV_X1 U7073 ( .A(n5954), .ZN(n5955) );
  MUX2_X1 U7074 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n4965), .Z(n5968) );
  XNOR2_X1 U7075 ( .A(n5971), .B(n5970), .ZN(n8217) );
  NAND2_X1 U7076 ( .A1(n8217), .A2(n6785), .ZN(n5959) );
  INV_X1 U7077 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8219) );
  OR2_X1 U7078 ( .A1(n6787), .A2(n8219), .ZN(n5958) );
  INV_X1 U7079 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5960) );
  NAND2_X1 U7080 ( .A1(n5961), .A2(n5960), .ZN(n5962) );
  AND2_X1 U7081 ( .A1(n5982), .A2(n5962), .ZN(n10275) );
  NAND2_X1 U7082 ( .A1(n10275), .A2(n5609), .ZN(n5965) );
  AOI22_X1 U7083 ( .A1(n5654), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n4958), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U7084 ( .A1(n5652), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5963) );
  INV_X1 U7085 ( .A(n10302), .ZN(n10388) );
  OR2_X1 U7086 ( .A1(n10273), .A2(n10388), .ZN(n5967) );
  NOR2_X1 U7087 ( .A1(n5968), .A2(SI_20_), .ZN(n5969) );
  MUX2_X1 U7088 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n4964), .Z(n5972) );
  NAND2_X1 U7089 ( .A1(n5972), .A2(SI_21_), .ZN(n5992) );
  INV_X1 U7090 ( .A(n5972), .ZN(n5973) );
  INV_X1 U7091 ( .A(SI_21_), .ZN(n8774) );
  NAND2_X1 U7092 ( .A1(n5973), .A2(n8774), .ZN(n5974) );
  NAND2_X1 U7093 ( .A1(n5992), .A2(n5974), .ZN(n5977) );
  INV_X1 U7094 ( .A(n5977), .ZN(n5975) );
  NAND2_X1 U7095 ( .A1(n5976), .A2(n5975), .ZN(n5993) );
  INV_X1 U7096 ( .A(n5976), .ZN(n5978) );
  NAND2_X1 U7097 ( .A1(n5978), .A2(n5977), .ZN(n5979) );
  NAND2_X1 U7098 ( .A1(n5993), .A2(n5979), .ZN(n8220) );
  INV_X1 U7099 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8222) );
  OR2_X1 U7100 ( .A1(n6787), .A2(n8222), .ZN(n5980) );
  INV_X1 U7101 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9891) );
  INV_X1 U7102 ( .A(n5996), .ZN(n5998) );
  NAND2_X1 U7103 ( .A1(n5982), .A2(n9891), .ZN(n5983) );
  NAND2_X1 U7104 ( .A1(n5998), .A2(n5983), .ZN(n10258) );
  OR2_X1 U7105 ( .A1(n10258), .A2(n6145), .ZN(n5989) );
  INV_X1 U7106 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7107 ( .A1(n5652), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5985) );
  NAND2_X1 U7108 ( .A1(n4958), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5984) );
  OAI211_X1 U7109 ( .C1(n5986), .C2(n6142), .A(n5985), .B(n5984), .ZN(n5987)
         );
  INV_X1 U7110 ( .A(n5987), .ZN(n5988) );
  NAND2_X1 U7111 ( .A1(n10390), .A2(n7120), .ZN(n6737) );
  NAND2_X1 U7112 ( .A1(n10257), .A2(n10256), .ZN(n5991) );
  OR2_X1 U7113 ( .A1(n10390), .A2(n10281), .ZN(n5990) );
  NAND2_X1 U7114 ( .A1(n5991), .A2(n5990), .ZN(n10237) );
  NAND2_X1 U7115 ( .A1(n5993), .A2(n5992), .ZN(n6009) );
  MUX2_X1 U7116 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n4965), .Z(n6008) );
  XNOR2_X1 U7117 ( .A(n6007), .B(SI_22_), .ZN(n8500) );
  NAND2_X1 U7118 ( .A1(n8500), .A2(n6785), .ZN(n5995) );
  INV_X1 U7119 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8502) );
  OR2_X1 U7120 ( .A1(n6787), .A2(n8502), .ZN(n5994) );
  NAND2_X1 U7121 ( .A1(n5996), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6013) );
  INV_X1 U7122 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5997) );
  NAND2_X1 U7123 ( .A1(n5998), .A2(n5997), .ZN(n5999) );
  NAND2_X1 U7124 ( .A1(n6013), .A2(n5999), .ZN(n10240) );
  OR2_X1 U7125 ( .A1(n10240), .A2(n6145), .ZN(n6005) );
  INV_X1 U7126 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U7127 ( .A1(n5652), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U7128 ( .A1(n5631), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6000) );
  OAI211_X1 U7129 ( .C1(n6002), .C2(n6142), .A(n6001), .B(n6000), .ZN(n6003)
         );
  INV_X1 U7130 ( .A(n6003), .ZN(n6004) );
  XNOR2_X1 U7131 ( .A(n10383), .B(n10377), .ZN(n6828) );
  INV_X1 U7132 ( .A(n10377), .ZN(n10254) );
  OR2_X1 U7133 ( .A1(n10383), .A2(n10254), .ZN(n6006) );
  MUX2_X1 U7134 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n4964), .Z(n6023) );
  XNOR2_X1 U7135 ( .A(n6023), .B(n8771), .ZN(n6021) );
  XNOR2_X1 U7136 ( .A(n6022), .B(n6021), .ZN(n8524) );
  NAND2_X1 U7137 ( .A1(n8524), .A2(n6785), .ZN(n6012) );
  INV_X1 U7138 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8527) );
  OR2_X1 U7139 ( .A1(n6787), .A2(n8527), .ZN(n6011) );
  INV_X1 U7140 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9874) );
  NAND2_X1 U7141 ( .A1(n6013), .A2(n9874), .ZN(n6014) );
  NAND2_X1 U7142 ( .A1(n6030), .A2(n6014), .ZN(n10227) );
  OR2_X1 U7143 ( .A1(n10227), .A2(n6145), .ZN(n6019) );
  INV_X1 U7144 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10380) );
  NAND2_X1 U7145 ( .A1(n5652), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U7146 ( .A1(n4958), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6015) );
  OAI211_X1 U7147 ( .C1(n10380), .C2(n6142), .A(n6016), .B(n6015), .ZN(n6017)
         );
  INV_X1 U7148 ( .A(n6017), .ZN(n6018) );
  NAND2_X1 U7149 ( .A1(n10234), .A2(n10245), .ZN(n6020) );
  INV_X1 U7150 ( .A(n6023), .ZN(n6024) );
  NAND2_X1 U7151 ( .A1(n6024), .A2(n8771), .ZN(n6025) );
  NAND2_X1 U7152 ( .A1(n6026), .A2(n6025), .ZN(n6040) );
  MUX2_X1 U7153 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n4965), .Z(n6041) );
  INV_X1 U7154 ( .A(SI_24_), .ZN(n6042) );
  XNOR2_X1 U7155 ( .A(n6041), .B(n6042), .ZN(n6039) );
  XNOR2_X1 U7156 ( .A(n6040), .B(n6039), .ZN(n8608) );
  NAND2_X1 U7157 ( .A1(n8608), .A2(n6785), .ZN(n6028) );
  INV_X1 U7158 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8613) );
  OR2_X1 U7159 ( .A1(n6787), .A2(n8613), .ZN(n6027) );
  INV_X1 U7160 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6029) );
  NAND2_X1 U7161 ( .A1(n6030), .A2(n6029), .ZN(n6031) );
  AND2_X1 U7162 ( .A1(n6051), .A2(n6031), .ZN(n9950) );
  NAND2_X1 U7163 ( .A1(n9950), .A2(n5609), .ZN(n6037) );
  INV_X1 U7164 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7165 ( .A1(n4958), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6033) );
  NAND2_X1 U7166 ( .A1(n5652), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6032) );
  OAI211_X1 U7167 ( .C1(n6034), .C2(n6142), .A(n6033), .B(n6032), .ZN(n6035)
         );
  INV_X1 U7168 ( .A(n6035), .ZN(n6036) );
  AND2_X1 U7169 ( .A1(n10372), .A2(n10205), .ZN(n6038) );
  NAND2_X1 U7170 ( .A1(n6040), .A2(n6039), .ZN(n6045) );
  INV_X1 U7171 ( .A(n6041), .ZN(n6043) );
  NAND2_X1 U7172 ( .A1(n6043), .A2(n6042), .ZN(n6044) );
  MUX2_X1 U7173 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(P2_DATAO_REG_25__SCAN_IN), 
        .S(n4965), .Z(n6046) );
  NAND2_X1 U7174 ( .A1(n6046), .A2(SI_25_), .ZN(n6060) );
  OAI21_X1 U7175 ( .B1(n6046), .B2(SI_25_), .A(n6060), .ZN(n6047) );
  NAND2_X1 U7176 ( .A1(n6048), .A2(n6047), .ZN(n6049) );
  INV_X1 U7177 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8625) );
  OR2_X1 U7178 ( .A1(n6787), .A2(n8625), .ZN(n6050) );
  INV_X1 U7179 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9911) );
  INV_X1 U7180 ( .A(n6064), .ZN(n6066) );
  NAND2_X1 U7181 ( .A1(n6051), .A2(n9911), .ZN(n6052) );
  NAND2_X1 U7182 ( .A1(n6066), .A2(n6052), .ZN(n10212) );
  OR2_X1 U7183 ( .A1(n10212), .A2(n6145), .ZN(n6057) );
  INV_X1 U7184 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n10368) );
  NAND2_X1 U7185 ( .A1(n5631), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6054) );
  NAND2_X1 U7186 ( .A1(n5652), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6053) );
  OAI211_X1 U7187 ( .C1(n6142), .C2(n10368), .A(n6054), .B(n6053), .ZN(n6055)
         );
  INV_X1 U7188 ( .A(n6055), .ZN(n6056) );
  NOR2_X1 U7189 ( .A1(n4961), .A2(n10030), .ZN(n6059) );
  NAND2_X1 U7190 ( .A1(n4961), .A2(n10030), .ZN(n6058) );
  MUX2_X1 U7191 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .S(n4965), .Z(n6076) );
  XNOR2_X1 U7192 ( .A(n6076), .B(SI_26_), .ZN(n6079) );
  XNOR2_X1 U7193 ( .A(n6080), .B(n6079), .ZN(n9853) );
  NAND2_X1 U7194 ( .A1(n9853), .A2(n6785), .ZN(n6063) );
  INV_X1 U7195 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10493) );
  OR2_X1 U7196 ( .A1(n6787), .A2(n10493), .ZN(n6062) );
  NAND2_X1 U7197 ( .A1(n6064), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6099) );
  INV_X1 U7198 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7199 ( .A1(n6066), .A2(n6065), .ZN(n6067) );
  NAND2_X1 U7200 ( .A1(n6099), .A2(n6067), .ZN(n10192) );
  OR2_X1 U7201 ( .A1(n10192), .A2(n6145), .ZN(n6072) );
  INV_X1 U7202 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10363) );
  NAND2_X1 U7203 ( .A1(n5631), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7204 ( .A1(n5652), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6068) );
  OAI211_X1 U7205 ( .C1(n6142), .C2(n10363), .A(n6069), .B(n6068), .ZN(n6070)
         );
  INV_X1 U7206 ( .A(n6070), .ZN(n6071) );
  OR2_X1 U7207 ( .A1(n10198), .A2(n10208), .ZN(n6834) );
  NAND2_X1 U7208 ( .A1(n10198), .A2(n10208), .ZN(n6746) );
  INV_X1 U7209 ( .A(n10190), .ZN(n6073) );
  NAND2_X1 U7210 ( .A1(n10191), .A2(n6073), .ZN(n6075) );
  NAND2_X1 U7211 ( .A1(n10198), .A2(n7768), .ZN(n6074) );
  INV_X1 U7212 ( .A(n6076), .ZN(n6077) );
  INV_X1 U7213 ( .A(SI_26_), .ZN(n8757) );
  NAND2_X1 U7214 ( .A1(n6077), .A2(n8757), .ZN(n6078) );
  MUX2_X1 U7215 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n4965), .Z(n6091) );
  XNOR2_X1 U7216 ( .A(n6091), .B(n8761), .ZN(n6089) );
  NAND2_X1 U7217 ( .A1(n10486), .A2(n6785), .ZN(n6082) );
  INV_X1 U7218 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10487) );
  OR2_X1 U7219 ( .A1(n6787), .A2(n10487), .ZN(n6081) );
  XNOR2_X1 U7220 ( .A(n6099), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n10179) );
  NAND2_X1 U7221 ( .A1(n10179), .A2(n5609), .ZN(n6087) );
  INV_X1 U7222 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10356) );
  NAND2_X1 U7223 ( .A1(n4958), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6084) );
  NAND2_X1 U7224 ( .A1(n5652), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6083) );
  OAI211_X1 U7225 ( .C1(n6142), .C2(n10356), .A(n6084), .B(n6083), .ZN(n6085)
         );
  INV_X1 U7226 ( .A(n6085), .ZN(n6086) );
  NAND2_X1 U7227 ( .A1(n10177), .A2(n7203), .ZN(n6833) );
  OR2_X1 U7228 ( .A1(n10177), .A2(n10188), .ZN(n6088) );
  NAND2_X1 U7229 ( .A1(n6090), .A2(n6089), .ZN(n6094) );
  INV_X1 U7230 ( .A(n6091), .ZN(n6092) );
  NAND2_X1 U7231 ( .A1(n6092), .A2(n8761), .ZN(n6093) );
  NAND2_X1 U7232 ( .A1(n6094), .A2(n6093), .ZN(n6756) );
  MUX2_X1 U7233 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n4965), .Z(n6757) );
  INV_X1 U7234 ( .A(SI_28_), .ZN(n6758) );
  XNOR2_X1 U7235 ( .A(n6757), .B(n6758), .ZN(n6755) );
  NAND2_X1 U7236 ( .A1(n9844), .A2(n6785), .ZN(n6096) );
  INV_X1 U7237 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10483) );
  OR2_X1 U7238 ( .A1(n6787), .A2(n10483), .ZN(n6095) );
  NAND2_X2 U7239 ( .A1(n6096), .A2(n6095), .ZN(n10157) );
  INV_X1 U7240 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n7214) );
  INV_X1 U7241 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6097) );
  OAI21_X1 U7242 ( .B1(n6099), .B2(n7214), .A(n6097), .ZN(n6100) );
  NAND2_X1 U7243 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6098) );
  NAND2_X1 U7244 ( .A1(n10158), .A2(n5609), .ZN(n6106) );
  INV_X1 U7245 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7246 ( .A1(n5631), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6102) );
  NAND2_X1 U7247 ( .A1(n5652), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6101) );
  OAI211_X1 U7248 ( .C1(n6103), .C2(n6142), .A(n6102), .B(n6101), .ZN(n6104)
         );
  INV_X1 U7249 ( .A(n6104), .ZN(n6105) );
  NOR2_X1 U7250 ( .A1(n10157), .A2(n10172), .ZN(n6837) );
  INV_X1 U7251 ( .A(n6837), .ZN(n6107) );
  NAND2_X1 U7252 ( .A1(n10157), .A2(n10172), .ZN(n10135) );
  NAND2_X1 U7253 ( .A1(n6108), .A2(n6750), .ZN(n6109) );
  INV_X1 U7254 ( .A(n6110), .ZN(n6111) );
  NAND2_X1 U7255 ( .A1(n6111), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6112) );
  XNOR2_X1 U7256 ( .A(n6162), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6117) );
  INV_X1 U7257 ( .A(n6946), .ZN(n6934) );
  MUX2_X1 U7258 ( .A(n6950), .B(n6934), .S(n8014), .Z(n6118) );
  NAND2_X1 U7259 ( .A1(n6118), .A2(n8011), .ZN(n7936) );
  INV_X1 U7260 ( .A(n6947), .ZN(n8501) );
  NOR2_X1 U7261 ( .A1(n6960), .A2(n8075), .ZN(n6813) );
  NAND2_X1 U7262 ( .A1(n8126), .A2(n6967), .ZN(n6120) );
  NAND2_X1 U7263 ( .A1(n6122), .A2(n6879), .ZN(n7946) );
  NAND2_X1 U7264 ( .A1(n8141), .A2(n8140), .ZN(n6123) );
  NAND2_X1 U7265 ( .A1(n6123), .A2(n6882), .ZN(n8103) );
  NAND2_X1 U7266 ( .A1(n6663), .A2(n6670), .ZN(n6124) );
  OR3_X1 U7267 ( .A1(n6124), .A2(n6688), .A3(n8245), .ZN(n6823) );
  AND2_X1 U7268 ( .A1(n6695), .A2(n8226), .ZN(n6821) );
  OR2_X1 U7269 ( .A1(n6124), .A2(n6821), .ZN(n6125) );
  AND2_X1 U7270 ( .A1(n6125), .A2(n6819), .ZN(n6891) );
  NAND2_X1 U7271 ( .A1(n8572), .A2(n8469), .ZN(n6811) );
  AND2_X1 U7272 ( .A1(n6811), .A2(n8391), .ZN(n6666) );
  OR2_X1 U7273 ( .A1(n8572), .A2(n8469), .ZN(n6812) );
  INV_X1 U7274 ( .A(n10836), .ZN(n9906) );
  NAND2_X1 U7275 ( .A1(n9906), .A2(n8570), .ZN(n6810) );
  OR2_X1 U7276 ( .A1(n8516), .A2(n9904), .ZN(n6897) );
  NAND2_X1 U7277 ( .A1(n8516), .A2(n9904), .ZN(n6719) );
  INV_X1 U7278 ( .A(n10031), .ZN(n10301) );
  OR2_X1 U7279 ( .A1(n10324), .A2(n10301), .ZN(n6916) );
  AND2_X1 U7280 ( .A1(n6916), .A2(n10308), .ZN(n6730) );
  NAND2_X1 U7281 ( .A1(n10324), .A2(n10301), .ZN(n6731) );
  NAND2_X1 U7282 ( .A1(n6127), .A2(n6731), .ZN(n10299) );
  NAND2_X1 U7283 ( .A1(n10298), .A2(n6910), .ZN(n10280) );
  INV_X1 U7284 ( .A(n6915), .ZN(n6128) );
  NAND2_X1 U7285 ( .A1(n6915), .A2(n6129), .ZN(n6130) );
  AND2_X1 U7286 ( .A1(n6130), .A2(n6737), .ZN(n6839) );
  INV_X1 U7287 ( .A(n6839), .ZN(n6131) );
  OR2_X1 U7288 ( .A1(n10383), .A2(n10377), .ZN(n6661) );
  OR2_X1 U7289 ( .A1(n10234), .A2(n9948), .ZN(n6740) );
  NAND2_X1 U7290 ( .A1(n10234), .A2(n9948), .ZN(n8920) );
  NAND2_X1 U7291 ( .A1(n6740), .A2(n8920), .ZN(n10225) );
  INV_X1 U7292 ( .A(n10225), .ZN(n10221) );
  NOR2_X1 U7293 ( .A1(n10372), .A2(n10222), .ZN(n6843) );
  INV_X1 U7294 ( .A(n6843), .ZN(n6135) );
  AND2_X1 U7295 ( .A1(n10372), .A2(n10222), .ZN(n6845) );
  NAND2_X1 U7296 ( .A1(n4961), .A2(n10360), .ZN(n6745) );
  INV_X1 U7297 ( .A(n10201), .ZN(n10204) );
  NAND2_X1 U7298 ( .A1(n10169), .A2(n6835), .ZN(n6136) );
  NAND2_X1 U7299 ( .A1(n6947), .A2(n4966), .ZN(n6138) );
  NAND2_X1 U7300 ( .A1(n6117), .A2(n6150), .ZN(n6137) );
  INV_X1 U7301 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U7302 ( .A1(n4958), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7303 ( .A1(n5652), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6139) );
  OAI211_X1 U7304 ( .C1(n6142), .C2(n6141), .A(n6140), .B(n6139), .ZN(n6143)
         );
  INV_X1 U7305 ( .A(n6143), .ZN(n6144) );
  OAI21_X1 U7306 ( .B1(n10149), .B2(n6145), .A(n6144), .ZN(n10029) );
  NAND2_X1 U7307 ( .A1(n5042), .A2(n6146), .ZN(n6860) );
  NAND2_X1 U7308 ( .A1(n6860), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6147) );
  INV_X1 U7309 ( .A(n7321), .ZN(n10485) );
  NAND2_X1 U7310 ( .A1(n10029), .A2(n10282), .ZN(n6148) );
  NAND2_X1 U7311 ( .A1(n8076), .A2(n8075), .ZN(n8123) );
  INV_X1 U7312 ( .A(n8234), .ZN(n10802) );
  NAND2_X1 U7313 ( .A1(n8251), .A2(n10802), .ZN(n8289) );
  INV_X1 U7314 ( .A(n8572), .ZN(n8437) );
  NAND2_X1 U7315 ( .A1(n8474), .A2(n10836), .ZN(n8515) );
  NOR2_X4 U7316 ( .A1(n8635), .A2(n10427), .ZN(n8634) );
  NAND2_X1 U7317 ( .A1(n10462), .A2(n10322), .ZN(n10291) );
  NOR2_X2 U7318 ( .A1(n10261), .A2(n10390), .ZN(n10238) );
  NAND2_X1 U7319 ( .A1(n9953), .A2(n8926), .ZN(n10210) );
  OR2_X2 U7320 ( .A1(n4961), .A2(n10210), .ZN(n10195) );
  NAND2_X1 U7321 ( .A1(n10157), .A2(n10176), .ZN(n6151) );
  NAND2_X1 U7322 ( .A1(n6151), .A2(n10292), .ZN(n6152) );
  OAI21_X1 U7323 ( .B1(n7203), .B2(n10395), .A(n10156), .ZN(n6153) );
  INV_X1 U7324 ( .A(n6154), .ZN(n6155) );
  NAND2_X1 U7325 ( .A1(n6155), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6156) );
  MUX2_X1 U7326 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6156), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n6158) );
  NAND2_X1 U7327 ( .A1(n6158), .A2(n6157), .ZN(n8626) );
  NAND2_X1 U7328 ( .A1(n8626), .A2(P1_B_REG_SCAN_IN), .ZN(n6165) );
  INV_X1 U7329 ( .A(n6159), .ZN(n6160) );
  NAND2_X1 U7330 ( .A1(n6160), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U7331 ( .A1(n6162), .A2(n6161), .ZN(n6164) );
  MUX2_X1 U7332 ( .A(n6165), .B(P1_B_REG_SCAN_IN), .S(n6170), .Z(n6167) );
  NAND2_X1 U7333 ( .A1(n6157), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6166) );
  INV_X1 U7334 ( .A(n10490), .ZN(n6191) );
  INV_X1 U7335 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n7421) );
  NAND2_X1 U7336 ( .A1(n7417), .A2(n7421), .ZN(n6168) );
  NAND2_X1 U7337 ( .A1(n10490), .A2(n8626), .ZN(n7419) );
  NAND2_X1 U7338 ( .A1(n6168), .A2(n7419), .ZN(n7182) );
  NAND2_X1 U7339 ( .A1(n10292), .A2(n4966), .ZN(n7189) );
  NAND2_X1 U7340 ( .A1(n7182), .A2(n7189), .ZN(n6189) );
  NOR2_X1 U7341 ( .A1(n10490), .A2(n8626), .ZN(n6169) );
  NAND2_X1 U7342 ( .A1(n6172), .A2(n6171), .ZN(n6173) );
  NAND2_X1 U7343 ( .A1(n6173), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U7344 ( .A1(n7315), .A2(n6946), .ZN(n7195) );
  AND2_X1 U7345 ( .A1(n7750), .A2(n7195), .ZN(n6188) );
  NOR4_X1 U7346 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6180) );
  NOR4_X1 U7347 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6179) );
  NOR4_X1 U7348 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6178) );
  NOR4_X1 U7349 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6177) );
  AND4_X1 U7350 ( .A1(n6180), .A2(n6179), .A3(n6178), .A4(n6177), .ZN(n6186)
         );
  NOR2_X1 U7351 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n6184) );
  NOR4_X1 U7352 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6183) );
  NOR4_X1 U7353 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6182) );
  NOR4_X1 U7354 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6181) );
  AND4_X1 U7355 ( .A1(n6184), .A2(n6183), .A3(n6182), .A4(n6181), .ZN(n6185)
         );
  NAND2_X1 U7356 ( .A1(n6186), .A2(n6185), .ZN(n6187) );
  NAND2_X1 U7357 ( .A1(n7417), .A2(n6187), .ZN(n7183) );
  NAND2_X1 U7358 ( .A1(n6188), .A2(n7183), .ZN(n7931) );
  INV_X1 U7359 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U7360 ( .A1(n7417), .A2(n6190), .ZN(n6192) );
  OR2_X1 U7361 ( .A1(n6170), .A2(n6191), .ZN(n10473) );
  INV_X1 U7362 ( .A(n7970), .ZN(n7184) );
  NAND2_X1 U7363 ( .A1(n10157), .A2(n8435), .ZN(n6193) );
  INV_X1 U7364 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6643) );
  INV_X1 U7365 ( .A(n6382), .ZN(n6201) );
  NAND2_X1 U7366 ( .A1(n6201), .A2(n6200), .ZN(n6445) );
  INV_X1 U7367 ( .A(n6445), .ZN(n6203) );
  NAND2_X1 U7368 ( .A1(n6203), .A2(n6202), .ZN(n6204) );
  NAND3_X1 U7369 ( .A1(n6208), .A2(n6404), .A3(n6207), .ZN(n6214) );
  NOR2_X1 U7370 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n6212) );
  NOR2_X1 U7371 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n6211) );
  NOR2_X1 U7372 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n6210) );
  NOR2_X1 U7373 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n6209) );
  NAND4_X1 U7374 ( .A1(n6212), .A2(n6211), .A3(n6210), .A4(n6209), .ZN(n6213)
         );
  NAND2_X1 U7375 ( .A1(n6635), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6216) );
  INV_X1 U7376 ( .A(n9464), .ZN(n7976) );
  NAND2_X1 U7377 ( .A1(n6221), .A2(n7976), .ZN(n6607) );
  NAND2_X1 U7378 ( .A1(n7295), .A2(n9773), .ZN(n7643) );
  AND2_X1 U7379 ( .A1(n6609), .A2(n8505), .ZN(n6220) );
  OR2_X1 U7380 ( .A1(n6227), .A2(n6352), .ZN(n6225) );
  NAND2_X1 U7381 ( .A1(n6227), .A2(n6226), .ZN(n6229) );
  NAND2_X1 U7382 ( .A1(n6228), .A2(n6229), .ZN(n6231) );
  NAND2_X1 U7383 ( .A1(n6269), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6235) );
  INV_X1 U7384 ( .A(n6231), .ZN(n9842) );
  AND2_X2 U7385 ( .A1(n9842), .A2(n9838), .ZN(n6273) );
  AND2_X2 U7386 ( .A1(n6231), .A2(n6230), .ZN(n6253) );
  NAND2_X1 U7387 ( .A1(n6253), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U7388 ( .A1(n6239), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6240) );
  NAND2_X1 U7389 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6241) );
  INV_X1 U7390 ( .A(n6242), .ZN(n6243) );
  INV_X1 U7391 ( .A(n10571), .ZN(n6245) );
  INV_X1 U7392 ( .A(n7265), .ZN(n7630) );
  NAND2_X1 U7393 ( .A1(n7625), .A2(n7265), .ZN(n9148) );
  NAND2_X1 U7394 ( .A1(n6253), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6250) );
  NAND2_X1 U7395 ( .A1(n6273), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6249) );
  NAND2_X1 U7396 ( .A1(n6269), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6248) );
  NAND2_X1 U7397 ( .A1(n6267), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U7398 ( .A1(n7346), .A2(SI_0_), .ZN(n6251) );
  XNOR2_X1 U7399 ( .A(n6251), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9857) );
  MUX2_X1 U7400 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9857), .S(n6599), .Z(n7648) );
  NAND2_X1 U7401 ( .A1(n7633), .A2(n7648), .ZN(n9144) );
  NAND2_X1 U7402 ( .A1(n6267), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6257) );
  INV_X1 U7403 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8833) );
  NAND2_X1 U7404 ( .A1(n6273), .A2(n8833), .ZN(n6256) );
  NAND2_X1 U7405 ( .A1(n6269), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6255) );
  INV_X1 U7406 ( .A(n6253), .ZN(n6268) );
  NAND2_X1 U7407 ( .A1(n6547), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6254) );
  NAND2_X1 U7408 ( .A1(n6258), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6266) );
  NAND2_X1 U7409 ( .A1(n6275), .A2(n6259), .ZN(n6265) );
  NAND2_X1 U7410 ( .A1(n6261), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6262) );
  MUX2_X1 U7411 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6262), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n6263) );
  NAND2_X1 U7412 ( .A1(n6457), .A2(n7745), .ZN(n6264) );
  NAND2_X1 U7413 ( .A1(n9391), .A2(n7880), .ZN(n9159) );
  NAND2_X1 U7414 ( .A1(n6267), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6272) );
  NAND2_X1 U7415 ( .A1(n6253), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6271) );
  NAND2_X1 U7416 ( .A1(n6269), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U7417 ( .A1(n6273), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6274) );
  NAND2_X1 U7418 ( .A1(n4991), .A2(n6274), .ZN(n9392) );
  NAND2_X1 U7419 ( .A1(n6258), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6282) );
  NAND2_X1 U7420 ( .A1(n6275), .A2(n7350), .ZN(n6281) );
  NAND2_X1 U7421 ( .A1(n6352), .A2(n6195), .ZN(n6276) );
  OAI21_X1 U7422 ( .B1(n6242), .B2(n6277), .A(n6276), .ZN(n6279) );
  INV_X1 U7423 ( .A(n6261), .ZN(n6278) );
  OR2_X1 U7424 ( .A1(n6599), .A2(n5441), .ZN(n6280) );
  NAND2_X1 U7425 ( .A1(n9392), .A2(n7895), .ZN(n6555) );
  AND2_X1 U7426 ( .A1(n9159), .A2(n6555), .ZN(n9157) );
  NAND2_X1 U7427 ( .A1(n7717), .A2(n9157), .ZN(n6286) );
  NOR2_X1 U7428 ( .A1(n9391), .A2(n7880), .ZN(n9155) );
  AOI21_X1 U7429 ( .B1(n9154), .B2(n9159), .A(n9155), .ZN(n6285) );
  NAND2_X1 U7430 ( .A1(n6286), .A2(n6285), .ZN(n6294) );
  NAND2_X1 U7431 ( .A1(n6269), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6291) );
  NAND2_X1 U7432 ( .A1(n6267), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6290) );
  AND2_X1 U7433 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6287) );
  NOR2_X1 U7434 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6295) );
  OR2_X1 U7435 ( .A1(n6287), .A2(n6295), .ZN(n7965) );
  NAND2_X1 U7436 ( .A1(n6273), .A2(n7965), .ZN(n6289) );
  NAND2_X1 U7437 ( .A1(n6547), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U7438 ( .A1(n6258), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6293) );
  XNOR2_X1 U7439 ( .A(n6303), .B(P2_IR_REG_4__SCAN_IN), .ZN(n10599) );
  NAND2_X1 U7440 ( .A1(n6457), .A2(n10599), .ZN(n6292) );
  INV_X1 U7441 ( .A(n7908), .ZN(n7428) );
  INV_X1 U7442 ( .A(n7966), .ZN(n7821) );
  NAND2_X1 U7443 ( .A1(n7428), .A2(n7821), .ZN(n9167) );
  NAND2_X1 U7444 ( .A1(n6294), .A2(n7816), .ZN(n7819) );
  NAND2_X1 U7445 ( .A1(n6269), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U7446 ( .A1(n6267), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6300) );
  NAND2_X1 U7447 ( .A1(n6295), .A2(n6296), .ZN(n6307) );
  OR2_X1 U7448 ( .A1(n6296), .A2(n6295), .ZN(n6297) );
  NAND2_X1 U7449 ( .A1(n6307), .A2(n6297), .ZN(n7914) );
  NAND2_X1 U7450 ( .A1(n6273), .A2(n7914), .ZN(n6299) );
  NAND2_X1 U7451 ( .A1(n6547), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6298) );
  NAND2_X1 U7452 ( .A1(n6258), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n6306) );
  NAND2_X1 U7453 ( .A1(n6303), .A2(n6302), .ZN(n6304) );
  NAND2_X1 U7454 ( .A1(n6304), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6314) );
  XNOR2_X1 U7455 ( .A(n6314), .B(P2_IR_REG_5__SCAN_IN), .ZN(n10610) );
  NAND2_X1 U7456 ( .A1(n6457), .A2(n10610), .ZN(n6305) );
  NAND2_X1 U7457 ( .A1(n8070), .A2(n7915), .ZN(n9162) );
  INV_X1 U7458 ( .A(n7915), .ZN(n7872) );
  NAND2_X1 U7459 ( .A1(n9390), .A2(n7872), .ZN(n9173) );
  NAND2_X1 U7460 ( .A1(n7865), .A2(n9332), .ZN(n7864) );
  NAND2_X1 U7461 ( .A1(n7864), .A2(n9162), .ZN(n8066) );
  NAND2_X1 U7462 ( .A1(n6595), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6312) );
  NAND2_X1 U7463 ( .A1(n6267), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6311) );
  NAND2_X1 U7464 ( .A1(n6307), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6308) );
  NAND2_X1 U7465 ( .A1(n6318), .A2(n6308), .ZN(n8097) );
  NAND2_X1 U7466 ( .A1(n6273), .A2(n8097), .ZN(n6310) );
  NAND2_X1 U7467 ( .A1(n6253), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6309) );
  NAND2_X1 U7468 ( .A1(n6258), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6317) );
  NAND2_X1 U7469 ( .A1(n6314), .A2(n6313), .ZN(n6315) );
  NAND2_X1 U7470 ( .A1(n6315), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6325) );
  XNOR2_X1 U7471 ( .A(n6325), .B(P2_IR_REG_6__SCAN_IN), .ZN(n8001) );
  NAND2_X1 U7472 ( .A1(n6457), .A2(n8001), .ZN(n6316) );
  OAI211_X1 U7473 ( .C1(n6513), .C2(n7363), .A(n6317), .B(n6316), .ZN(n8098)
         );
  NAND2_X1 U7474 ( .A1(n7907), .A2(n8098), .ZN(n9177) );
  INV_X1 U7475 ( .A(n8098), .ZN(n8067) );
  NAND2_X1 U7476 ( .A1(n9389), .A2(n8067), .ZN(n9172) );
  AND2_X1 U7477 ( .A1(n9177), .A2(n9172), .ZN(n9329) );
  NAND2_X1 U7478 ( .A1(n8066), .A2(n9329), .ZN(n8026) );
  NAND2_X1 U7479 ( .A1(n6267), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6323) );
  NAND2_X1 U7480 ( .A1(n6595), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6322) );
  AND2_X1 U7481 ( .A1(n6318), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6319) );
  OR2_X1 U7482 ( .A1(n6319), .A2(n6335), .ZN(n8179) );
  NAND2_X1 U7483 ( .A1(n6594), .A2(n8179), .ZN(n6321) );
  NAND2_X1 U7484 ( .A1(n6253), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6320) );
  NAND2_X1 U7485 ( .A1(n6325), .A2(n6324), .ZN(n6326) );
  NAND2_X1 U7486 ( .A1(n6326), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6330) );
  XNOR2_X1 U7487 ( .A(n6330), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7979) );
  AOI22_X1 U7488 ( .A1(n6258), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6457), .B2(
        n7979), .ZN(n6327) );
  NAND2_X1 U7489 ( .A1(n8191), .A2(n8180), .ZN(n9183) );
  NAND2_X1 U7490 ( .A1(n9388), .A2(n8212), .ZN(n9191) );
  NAND2_X1 U7491 ( .A1(n9183), .A2(n9191), .ZN(n9336) );
  INV_X1 U7492 ( .A(n9177), .ZN(n8027) );
  NOR2_X1 U7493 ( .A1(n9336), .A2(n8027), .ZN(n6328) );
  NAND2_X1 U7494 ( .A1(n8026), .A2(n6328), .ZN(n8029) );
  NAND2_X1 U7495 ( .A1(n7377), .A2(n6275), .ZN(n6334) );
  INV_X1 U7496 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6329) );
  NAND2_X1 U7497 ( .A1(n6330), .A2(n6329), .ZN(n6331) );
  NAND2_X1 U7498 ( .A1(n6331), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6332) );
  XNOR2_X1 U7499 ( .A(n6332), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7998) );
  AOI22_X1 U7500 ( .A1(n6258), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6457), .B2(
        n7998), .ZN(n6333) );
  NAND2_X1 U7501 ( .A1(n6267), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6340) );
  NOR2_X1 U7502 ( .A1(n6335), .A2(n8750), .ZN(n6336) );
  OR2_X1 U7503 ( .A1(n6346), .A2(n6336), .ZN(n8198) );
  NAND2_X1 U7504 ( .A1(n6273), .A2(n8198), .ZN(n6339) );
  INV_X2 U7505 ( .A(n6268), .ZN(n6547) );
  NAND2_X1 U7506 ( .A1(n6547), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6338) );
  NAND2_X1 U7507 ( .A1(n6595), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6337) );
  NAND4_X1 U7508 ( .A1(n6340), .A2(n6339), .A3(n6338), .A4(n6337), .ZN(n9387)
         );
  AND2_X1 U7509 ( .A1(n8193), .A2(n9387), .ZN(n9193) );
  INV_X1 U7510 ( .A(n8193), .ZN(n8202) );
  NAND2_X1 U7511 ( .A1(n8415), .A2(n8202), .ZN(n9184) );
  NAND2_X1 U7512 ( .A1(n7398), .A2(n6275), .ZN(n6344) );
  OR2_X1 U7513 ( .A1(n6341), .A2(n6352), .ZN(n6342) );
  XNOR2_X1 U7514 ( .A(n6342), .B(P2_IR_REG_9__SCAN_IN), .ZN(n9413) );
  AOI22_X1 U7515 ( .A1(n6258), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6457), .B2(
        n9413), .ZN(n6343) );
  NAND2_X1 U7516 ( .A1(n6344), .A2(n6343), .ZN(n8426) );
  NAND2_X1 U7517 ( .A1(n6595), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6351) );
  NAND2_X1 U7518 ( .A1(n6267), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6350) );
  OR2_X1 U7519 ( .A1(n6346), .A2(n6345), .ZN(n6347) );
  NAND2_X1 U7520 ( .A1(n6357), .A2(n6347), .ZN(n8421) );
  NAND2_X1 U7521 ( .A1(n6273), .A2(n8421), .ZN(n6349) );
  NAND2_X1 U7522 ( .A1(n6253), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6348) );
  NAND2_X1 U7523 ( .A1(n8426), .A2(n8577), .ZN(n9185) );
  NAND2_X1 U7524 ( .A1(n9194), .A2(n9185), .ZN(n8321) );
  OR2_X1 U7525 ( .A1(n7397), .A2(n6513), .ZN(n6356) );
  OR2_X1 U7526 ( .A1(n6353), .A2(n6352), .ZN(n6354) );
  XNOR2_X1 U7527 ( .A(n6354), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10623) );
  AOI22_X1 U7528 ( .A1(n6258), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6457), .B2(
        n10623), .ZN(n6355) );
  NAND2_X1 U7529 ( .A1(n6356), .A2(n6355), .ZN(n8583) );
  NAND2_X1 U7530 ( .A1(n6267), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6362) );
  NAND2_X1 U7531 ( .A1(n6253), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6361) );
  NAND2_X1 U7532 ( .A1(n6357), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6358) );
  NAND2_X1 U7533 ( .A1(n6367), .A2(n6358), .ZN(n8579) );
  NAND2_X1 U7534 ( .A1(n6273), .A2(n8579), .ZN(n6360) );
  NAND2_X1 U7535 ( .A1(n6595), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6359) );
  NAND2_X1 U7536 ( .A1(n8583), .A2(n9100), .ZN(n9197) );
  NAND2_X1 U7537 ( .A1(n8887), .A2(n6275), .ZN(n6366) );
  NAND2_X1 U7538 ( .A1(n4985), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6363) );
  MUX2_X1 U7539 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6363), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n6364) );
  AND2_X1 U7540 ( .A1(n6364), .A2(n5029), .ZN(n10641) );
  AOI22_X1 U7541 ( .A1(n6258), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6457), .B2(
        n10641), .ZN(n6365) );
  NAND2_X1 U7542 ( .A1(n6366), .A2(n6365), .ZN(n6569) );
  NAND2_X1 U7543 ( .A1(n6595), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6372) );
  NAND2_X1 U7544 ( .A1(n6267), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6371) );
  AND2_X1 U7545 ( .A1(n6367), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6368) );
  OR2_X1 U7546 ( .A1(n6376), .A2(n6368), .ZN(n9103) );
  NAND2_X1 U7547 ( .A1(n6273), .A2(n9103), .ZN(n6370) );
  NAND2_X1 U7548 ( .A1(n6253), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6369) );
  OR2_X1 U7549 ( .A1(n6569), .A2(n9094), .ZN(n9202) );
  NAND2_X1 U7550 ( .A1(n6569), .A2(n9094), .ZN(n9200) );
  NAND2_X1 U7551 ( .A1(n8482), .A2(n9343), .ZN(n8481) );
  OR2_X1 U7552 ( .A1(n7432), .A2(n6513), .ZN(n6375) );
  NAND2_X1 U7553 ( .A1(n5029), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6373) );
  XNOR2_X1 U7554 ( .A(n6373), .B(P2_IR_REG_12__SCAN_IN), .ZN(n10657) );
  AOI22_X1 U7555 ( .A1(n6258), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6457), .B2(
        n10657), .ZN(n6374) );
  NAND2_X1 U7556 ( .A1(n6375), .A2(n6374), .ZN(n9770) );
  NAND2_X1 U7557 ( .A1(n6595), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6381) );
  NAND2_X1 U7558 ( .A1(n6267), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6380) );
  OR2_X1 U7559 ( .A1(n6376), .A2(n8846), .ZN(n6377) );
  NAND2_X1 U7560 ( .A1(n6377), .A2(n6385), .ZN(n8596) );
  NAND2_X1 U7561 ( .A1(n6273), .A2(n8596), .ZN(n6379) );
  NAND2_X1 U7562 ( .A1(n6253), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6378) );
  OR2_X1 U7563 ( .A1(n9770), .A2(n9683), .ZN(n9206) );
  NAND2_X1 U7564 ( .A1(n9770), .A2(n9683), .ZN(n9207) );
  NAND2_X1 U7565 ( .A1(n7515), .A2(n6275), .ZN(n6384) );
  NAND2_X1 U7566 ( .A1(n6382), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6393) );
  XNOR2_X1 U7567 ( .A(n6393), .B(P2_IR_REG_13__SCAN_IN), .ZN(n10673) );
  AOI22_X1 U7568 ( .A1(n6258), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6457), .B2(
        n10673), .ZN(n6383) );
  NAND2_X1 U7569 ( .A1(n6267), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6391) );
  NAND2_X1 U7570 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(n6385), .ZN(n6387) );
  INV_X1 U7571 ( .A(n6397), .ZN(n6386) );
  NAND2_X1 U7572 ( .A1(n6387), .A2(n6386), .ZN(n9687) );
  NAND2_X1 U7573 ( .A1(n6273), .A2(n9687), .ZN(n6390) );
  NAND2_X1 U7574 ( .A1(n6595), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6389) );
  NAND2_X1 U7575 ( .A1(n6253), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6388) );
  NAND4_X1 U7576 ( .A1(n6391), .A2(n6390), .A3(n6389), .A4(n6388), .ZN(n9383)
         );
  XNOR2_X1 U7577 ( .A(n9677), .B(n9383), .ZN(n9690) );
  INV_X1 U7578 ( .A(n9383), .ZN(n9666) );
  NAND2_X1 U7579 ( .A1(n7533), .A2(n6275), .ZN(n6396) );
  NAND2_X1 U7580 ( .A1(n6393), .A2(n6392), .ZN(n6394) );
  NAND2_X1 U7581 ( .A1(n6394), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6405) );
  XNOR2_X1 U7582 ( .A(n6405), .B(P2_IR_REG_14__SCAN_IN), .ZN(n10689) );
  AOI22_X1 U7583 ( .A1(n6258), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6457), .B2(
        n10689), .ZN(n6395) );
  NAND2_X1 U7584 ( .A1(n6267), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6401) );
  OAI21_X1 U7585 ( .B1(n8823), .B2(n6397), .A(n6409), .ZN(n9668) );
  NAND2_X1 U7586 ( .A1(n6273), .A2(n9668), .ZN(n6400) );
  NAND2_X1 U7587 ( .A1(n6595), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6399) );
  NAND2_X1 U7588 ( .A1(n6253), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6398) );
  NAND4_X1 U7589 ( .A1(n6401), .A2(n6400), .A3(n6399), .A4(n6398), .ZN(n9382)
         );
  NAND2_X1 U7590 ( .A1(n9757), .A2(n9382), .ZN(n9216) );
  OR2_X1 U7591 ( .A1(n9757), .A2(n9382), .ZN(n6402) );
  OR2_X1 U7592 ( .A1(n9757), .A2(n8943), .ZN(n6403) );
  NAND2_X1 U7593 ( .A1(n6405), .A2(n6404), .ZN(n6406) );
  NAND2_X1 U7594 ( .A1(n6406), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6418) );
  XNOR2_X1 U7595 ( .A(n6418), .B(P2_IR_REG_15__SCAN_IN), .ZN(n10705) );
  AOI22_X1 U7596 ( .A1(n6258), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6457), .B2(
        n10705), .ZN(n6407) );
  NAND2_X1 U7597 ( .A1(n6267), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6414) );
  NAND2_X1 U7598 ( .A1(n6409), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6410) );
  INV_X1 U7599 ( .A(n6426), .ZN(n6425) );
  NAND2_X1 U7600 ( .A1(n6410), .A2(n6425), .ZN(n9653) );
  NAND2_X1 U7601 ( .A1(n6594), .A2(n9653), .ZN(n6413) );
  NAND2_X1 U7602 ( .A1(n6595), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6412) );
  NAND2_X1 U7603 ( .A1(n6253), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6411) );
  NAND4_X1 U7604 ( .A1(n6414), .A2(n6413), .A3(n6412), .A4(n6411), .ZN(n9381)
         );
  NAND2_X1 U7605 ( .A1(n9834), .A2(n9381), .ZN(n6415) );
  NAND2_X1 U7606 ( .A1(n9220), .A2(n9667), .ZN(n6416) );
  NAND2_X1 U7607 ( .A1(n6415), .A2(n6416), .ZN(n9649) );
  NAND2_X1 U7608 ( .A1(n7726), .A2(n6275), .ZN(n6424) );
  INV_X1 U7609 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6417) );
  NAND2_X1 U7610 ( .A1(n6418), .A2(n6417), .ZN(n6419) );
  NAND2_X1 U7611 ( .A1(n6419), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6421) );
  INV_X1 U7612 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6420) );
  NAND2_X1 U7613 ( .A1(n6421), .A2(n6420), .ZN(n6432) );
  OR2_X1 U7614 ( .A1(n6421), .A2(n6420), .ZN(n6422) );
  AOI22_X1 U7615 ( .A1(n6258), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6457), .B2(
        n10721), .ZN(n6423) );
  NAND2_X1 U7616 ( .A1(n6424), .A2(n6423), .ZN(n9640) );
  NAND2_X1 U7617 ( .A1(n6595), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6431) );
  NAND2_X1 U7618 ( .A1(n6267), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6430) );
  NAND2_X1 U7619 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(n6425), .ZN(n6427) );
  NAND2_X1 U7620 ( .A1(n8851), .A2(n6426), .ZN(n6438) );
  NAND2_X1 U7621 ( .A1(n6427), .A2(n6438), .ZN(n9641) );
  NAND2_X1 U7622 ( .A1(n6594), .A2(n9641), .ZN(n6429) );
  NAND2_X1 U7623 ( .A1(n6547), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6428) );
  OR2_X1 U7624 ( .A1(n9640), .A2(n9648), .ZN(n9226) );
  NAND2_X1 U7625 ( .A1(n9640), .A2(n9648), .ZN(n9225) );
  NAND2_X1 U7626 ( .A1(n7792), .A2(n6275), .ZN(n6435) );
  NAND2_X1 U7627 ( .A1(n6432), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6433) );
  XNOR2_X1 U7628 ( .A(n6433), .B(P2_IR_REG_17__SCAN_IN), .ZN(n10738) );
  AOI22_X1 U7629 ( .A1(n6258), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6457), .B2(
        n10738), .ZN(n6434) );
  NAND2_X1 U7630 ( .A1(n6595), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6443) );
  NAND2_X1 U7631 ( .A1(n6267), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6442) );
  INV_X1 U7632 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6437) );
  INV_X1 U7633 ( .A(n6438), .ZN(n6436) );
  NAND2_X1 U7634 ( .A1(n6437), .A2(n6436), .ZN(n6450) );
  NAND2_X1 U7635 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(n6438), .ZN(n6439) );
  NAND2_X1 U7636 ( .A1(n6450), .A2(n6439), .ZN(n9628) );
  NAND2_X1 U7637 ( .A1(n6273), .A2(n9628), .ZN(n6441) );
  NAND2_X1 U7638 ( .A1(n6547), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6440) );
  XNOR2_X1 U7639 ( .A(n9234), .B(n9636), .ZN(n9624) );
  OR2_X1 U7640 ( .A1(n9234), .A2(n9636), .ZN(n6444) );
  NAND2_X1 U7641 ( .A1(n9627), .A2(n6444), .ZN(n9614) );
  NAND2_X1 U7642 ( .A1(n7927), .A2(n6275), .ZN(n6448) );
  NAND2_X1 U7643 ( .A1(n6445), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6446) );
  XNOR2_X1 U7644 ( .A(n6446), .B(P2_IR_REG_18__SCAN_IN), .ZN(n10767) );
  AOI22_X1 U7645 ( .A1(n6258), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6457), .B2(
        n10767), .ZN(n6447) );
  NAND2_X1 U7646 ( .A1(n6595), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6455) );
  NAND2_X1 U7647 ( .A1(n6267), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6454) );
  INV_X1 U7648 ( .A(n6450), .ZN(n6449) );
  NAND2_X1 U7649 ( .A1(n6450), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6451) );
  NAND2_X1 U7650 ( .A1(n6460), .A2(n6451), .ZN(n9616) );
  NAND2_X1 U7651 ( .A1(n6594), .A2(n9616), .ZN(n6453) );
  NAND2_X1 U7652 ( .A1(n6547), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6452) );
  NAND2_X1 U7653 ( .A1(n9106), .A2(n9623), .ZN(n9232) );
  NAND2_X1 U7654 ( .A1(n7974), .A2(n6275), .ZN(n6459) );
  AOI22_X1 U7655 ( .A1(n6258), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9464), .B2(
        n6457), .ZN(n6458) );
  NAND2_X1 U7656 ( .A1(n6267), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6465) );
  NAND2_X1 U7657 ( .A1(n6595), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6464) );
  NAND2_X1 U7658 ( .A1(n6460), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6461) );
  NAND2_X1 U7659 ( .A1(n6469), .A2(n6461), .ZN(n9606) );
  NAND2_X1 U7660 ( .A1(n6273), .A2(n9606), .ZN(n6463) );
  NAND2_X1 U7661 ( .A1(n6547), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6462) );
  NOR2_X1 U7662 ( .A1(n9014), .A2(n9613), .ZN(n9243) );
  NAND2_X1 U7663 ( .A1(n9014), .A2(n9613), .ZN(n9241) );
  NAND2_X1 U7664 ( .A1(n8217), .A2(n6275), .ZN(n6467) );
  NAND2_X1 U7665 ( .A1(n6258), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6466) );
  NAND2_X1 U7666 ( .A1(n6267), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6474) );
  NAND2_X1 U7667 ( .A1(n6595), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6473) );
  NAND2_X1 U7668 ( .A1(n6469), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6470) );
  NAND2_X1 U7669 ( .A1(n6477), .A2(n6470), .ZN(n9595) );
  NAND2_X1 U7670 ( .A1(n6273), .A2(n9595), .ZN(n6472) );
  NAND2_X1 U7671 ( .A1(n6253), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6471) );
  NAND2_X1 U7672 ( .A1(n9594), .A2(n9603), .ZN(n9249) );
  NAND2_X1 U7673 ( .A1(n9248), .A2(n9249), .ZN(n9328) );
  OR2_X1 U7674 ( .A1(n8220), .A2(n6513), .ZN(n6476) );
  NAND2_X1 U7675 ( .A1(n6258), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6475) );
  NAND2_X1 U7676 ( .A1(n6267), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6482) );
  NAND2_X1 U7677 ( .A1(n6477), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6478) );
  NAND2_X1 U7678 ( .A1(n6486), .A2(n6478), .ZN(n9578) );
  NAND2_X1 U7679 ( .A1(n6594), .A2(n9578), .ZN(n6481) );
  NAND2_X1 U7680 ( .A1(n6595), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6480) );
  NAND2_X1 U7681 ( .A1(n6547), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6479) );
  NAND4_X1 U7682 ( .A1(n6482), .A2(n6481), .A3(n6480), .A4(n6479), .ZN(n9376)
         );
  NAND2_X1 U7683 ( .A1(n9577), .A2(n9376), .ZN(n9254) );
  NAND2_X1 U7684 ( .A1(n9247), .A2(n9254), .ZN(n9580) );
  INV_X1 U7685 ( .A(n9376), .ZN(n9592) );
  NAND2_X1 U7686 ( .A1(n8500), .A2(n6275), .ZN(n6484) );
  NAND2_X1 U7687 ( .A1(n6258), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6483) );
  NAND2_X1 U7688 ( .A1(n6595), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6491) );
  NAND2_X1 U7689 ( .A1(n6267), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6490) );
  INV_X1 U7690 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8866) );
  NAND2_X1 U7691 ( .A1(n6486), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6487) );
  NAND2_X1 U7692 ( .A1(n6497), .A2(n6487), .ZN(n9567) );
  NAND2_X1 U7693 ( .A1(n6594), .A2(n9567), .ZN(n6489) );
  NAND2_X1 U7694 ( .A1(n6547), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6488) );
  NAND2_X1 U7695 ( .A1(n9258), .A2(n9576), .ZN(n6492) );
  NAND2_X1 U7696 ( .A1(n9566), .A2(n6492), .ZN(n6494) );
  OR2_X1 U7697 ( .A1(n9258), .A2(n9576), .ZN(n6493) );
  NAND2_X1 U7698 ( .A1(n8524), .A2(n6275), .ZN(n6496) );
  NAND2_X1 U7699 ( .A1(n6258), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6495) );
  NAND2_X1 U7700 ( .A1(n6267), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6502) );
  NAND2_X1 U7701 ( .A1(n6497), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6498) );
  NAND2_X1 U7702 ( .A1(n6506), .A2(n6498), .ZN(n9557) );
  NAND2_X1 U7703 ( .A1(n6594), .A2(n9557), .ZN(n6501) );
  NAND2_X1 U7704 ( .A1(n6253), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6500) );
  NAND2_X1 U7705 ( .A1(n6595), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6499) );
  NAND4_X1 U7706 ( .A1(n6502), .A2(n6501), .A3(n6500), .A4(n6499), .ZN(n9539)
         );
  AND2_X1 U7707 ( .A1(n9801), .A2(n9539), .ZN(n9263) );
  NAND2_X1 U7708 ( .A1(n8608), .A2(n6275), .ZN(n6504) );
  NAND2_X1 U7709 ( .A1(n6258), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6503) );
  NAND2_X1 U7710 ( .A1(n6595), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6511) );
  NAND2_X1 U7711 ( .A1(n6267), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6510) );
  INV_X1 U7712 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8732) );
  NAND2_X1 U7713 ( .A1(n6506), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6507) );
  NAND2_X1 U7714 ( .A1(n6516), .A2(n6507), .ZN(n9532) );
  NAND2_X1 U7715 ( .A1(n6273), .A2(n9532), .ZN(n6509) );
  NAND2_X1 U7716 ( .A1(n6547), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6508) );
  XNOR2_X1 U7717 ( .A(n9531), .B(n9554), .ZN(n9547) );
  OR2_X1 U7718 ( .A1(n9531), .A2(n9554), .ZN(n9266) );
  NAND2_X1 U7719 ( .A1(n6258), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6514) );
  NAND2_X1 U7720 ( .A1(n6595), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6521) );
  NAND2_X1 U7721 ( .A1(n6267), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6520) );
  NAND2_X1 U7722 ( .A1(n6516), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6517) );
  NAND2_X1 U7723 ( .A1(n6528), .A2(n6517), .ZN(n9526) );
  NAND2_X1 U7724 ( .A1(n6594), .A2(n9526), .ZN(n6519) );
  NAND2_X1 U7725 ( .A1(n6253), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6518) );
  NAND2_X1 U7726 ( .A1(n9518), .A2(n8975), .ZN(n6522) );
  NAND2_X1 U7727 ( .A1(n9527), .A2(n6522), .ZN(n6524) );
  OR2_X1 U7728 ( .A1(n9518), .A2(n8975), .ZN(n6523) );
  NAND2_X1 U7729 ( .A1(n9853), .A2(n6275), .ZN(n6526) );
  NAND2_X1 U7730 ( .A1(n6258), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6525) );
  NAND2_X1 U7731 ( .A1(n6267), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6533) );
  INV_X1 U7732 ( .A(n6528), .ZN(n6527) );
  INV_X1 U7733 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8876) );
  NAND2_X1 U7734 ( .A1(n6527), .A2(n8876), .ZN(n6537) );
  NAND2_X1 U7735 ( .A1(n6528), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6529) );
  NAND2_X1 U7736 ( .A1(n6537), .A2(n6529), .ZN(n9513) );
  NAND2_X1 U7737 ( .A1(n6594), .A2(n9513), .ZN(n6532) );
  NAND2_X1 U7738 ( .A1(n6547), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6531) );
  NAND2_X1 U7739 ( .A1(n6595), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6530) );
  NAND4_X1 U7740 ( .A1(n6533), .A2(n6532), .A3(n6531), .A4(n6530), .ZN(n9521)
         );
  AND2_X1 U7741 ( .A1(n9515), .A2(n9521), .ZN(n9309) );
  INV_X1 U7742 ( .A(n9521), .ZN(n6534) );
  NAND2_X1 U7743 ( .A1(n9703), .A2(n6534), .ZN(n9508) );
  NAND2_X1 U7744 ( .A1(n10486), .A2(n6275), .ZN(n6536) );
  NAND2_X1 U7745 ( .A1(n6258), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6535) );
  NAND2_X1 U7746 ( .A1(n6595), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6542) );
  NAND2_X1 U7747 ( .A1(n6267), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6541) );
  NAND2_X1 U7748 ( .A1(n6537), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6538) );
  NAND2_X1 U7749 ( .A1(n6545), .A2(n6538), .ZN(n9500) );
  NAND2_X1 U7750 ( .A1(n6594), .A2(n9500), .ZN(n6540) );
  NAND2_X1 U7751 ( .A1(n6547), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6539) );
  NAND2_X1 U7752 ( .A1(n9844), .A2(n6275), .ZN(n6544) );
  NAND2_X1 U7753 ( .A1(n6258), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6543) );
  NAND2_X1 U7754 ( .A1(n6595), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6551) );
  NAND2_X1 U7755 ( .A1(n6267), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6550) );
  NAND2_X1 U7756 ( .A1(n6545), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U7757 ( .A1(n9473), .A2(n6546), .ZN(n9487) );
  NAND2_X1 U7758 ( .A1(n6594), .A2(n9487), .ZN(n6549) );
  NAND2_X1 U7759 ( .A1(n6547), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6548) );
  NAND2_X1 U7760 ( .A1(n9282), .A2(n9499), .ZN(n9314) );
  XOR2_X1 U7761 ( .A(n7221), .B(n9351), .Z(n9491) );
  NAND2_X1 U7762 ( .A1(n6552), .A2(n7648), .ZN(n7631) );
  NAND2_X1 U7763 ( .A1(n7628), .A2(n7631), .ZN(n6554) );
  NAND2_X1 U7764 ( .A1(n7625), .A2(n7630), .ZN(n6553) );
  NAND2_X1 U7765 ( .A1(n7720), .A2(n7716), .ZN(n6557) );
  NAND2_X1 U7766 ( .A1(n6284), .A2(n7895), .ZN(n6556) );
  NAND2_X1 U7767 ( .A1(n6557), .A2(n6556), .ZN(n7787) );
  INV_X1 U7768 ( .A(n7787), .ZN(n6558) );
  NAND2_X1 U7769 ( .A1(n9391), .A2(n7713), .ZN(n6559) );
  AND2_X1 U7770 ( .A1(n7428), .A2(n7966), .ZN(n6561) );
  NAND2_X1 U7771 ( .A1(n9390), .A2(n7915), .ZN(n6562) );
  AND2_X1 U7772 ( .A1(n9389), .A2(n8098), .ZN(n6565) );
  NAND2_X1 U7773 ( .A1(n7907), .A2(n8067), .ZN(n6564) );
  INV_X1 U7774 ( .A(n9193), .ZN(n9174) );
  NAND2_X1 U7775 ( .A1(n9174), .A2(n9184), .ZN(n8189) );
  NAND2_X1 U7776 ( .A1(n8193), .A2(n8415), .ZN(n6566) );
  INV_X1 U7777 ( .A(n8577), .ZN(n8578) );
  OR2_X1 U7778 ( .A1(n8426), .A2(n8578), .ZN(n6568) );
  INV_X1 U7779 ( .A(n9100), .ZN(n9386) );
  INV_X1 U7780 ( .A(n9094), .ZN(n9385) );
  NAND2_X1 U7781 ( .A1(n6571), .A2(n9385), .ZN(n6570) );
  NAND2_X1 U7782 ( .A1(n6570), .A2(n9774), .ZN(n6573) );
  NAND2_X1 U7783 ( .A1(n4957), .A2(n9094), .ZN(n6572) );
  INV_X1 U7784 ( .A(n9683), .ZN(n9384) );
  NAND2_X1 U7785 ( .A1(n9770), .A2(n9384), .ZN(n6574) );
  OR2_X1 U7786 ( .A1(n9677), .A2(n9383), .ZN(n6575) );
  NAND2_X1 U7787 ( .A1(n9677), .A2(n9383), .ZN(n6576) );
  NAND2_X1 U7788 ( .A1(n6577), .A2(n9216), .ZN(n9646) );
  NAND2_X1 U7789 ( .A1(n9646), .A2(n9649), .ZN(n6579) );
  NAND2_X1 U7790 ( .A1(n9220), .A2(n9381), .ZN(n6578) );
  NAND2_X1 U7791 ( .A1(n6579), .A2(n6578), .ZN(n9633) );
  INV_X1 U7792 ( .A(n9638), .ZN(n9634) );
  NAND2_X1 U7793 ( .A1(n9633), .A2(n9634), .ZN(n6581) );
  INV_X1 U7794 ( .A(n9648), .ZN(n9380) );
  NAND2_X1 U7795 ( .A1(n9640), .A2(n9380), .ZN(n6580) );
  NAND2_X1 U7796 ( .A1(n6581), .A2(n6580), .ZN(n9621) );
  NAND2_X1 U7797 ( .A1(n9621), .A2(n9624), .ZN(n6583) );
  INV_X1 U7798 ( .A(n9636), .ZN(n9379) );
  NAND2_X1 U7799 ( .A1(n9234), .A2(n9379), .ZN(n6582) );
  NAND2_X1 U7800 ( .A1(n6583), .A2(n6582), .ZN(n9611) );
  AND2_X1 U7801 ( .A1(n9106), .A2(n8952), .ZN(n6584) );
  OR2_X1 U7802 ( .A1(n9106), .A2(n8952), .ZN(n6585) );
  NAND2_X1 U7803 ( .A1(n9014), .A2(n9378), .ZN(n8955) );
  INV_X1 U7804 ( .A(n9603), .ZN(n9377) );
  OR2_X1 U7805 ( .A1(n9594), .A2(n9377), .ZN(n9572) );
  NAND2_X1 U7806 ( .A1(n9588), .A2(n9572), .ZN(n6586) );
  NAND2_X1 U7807 ( .A1(n6586), .A2(n5360), .ZN(n9574) );
  NOR2_X1 U7808 ( .A1(n9258), .A2(n9375), .ZN(n9141) );
  NAND2_X1 U7809 ( .A1(n9258), .A2(n9375), .ZN(n9259) );
  OR2_X1 U7810 ( .A1(n9539), .A2(n9011), .ZN(n6587) );
  NAND2_X1 U7811 ( .A1(n9011), .A2(n9539), .ZN(n6588) );
  INV_X1 U7812 ( .A(n9547), .ZN(n9535) );
  OR2_X1 U7813 ( .A1(n9531), .A2(n9522), .ZN(n6589) );
  NAND2_X1 U7814 ( .A1(n9537), .A2(n6589), .ZN(n9520) );
  XNOR2_X1 U7815 ( .A(n9518), .B(n8975), .ZN(n9528) );
  NAND2_X1 U7816 ( .A1(n9520), .A2(n9528), .ZN(n9519) );
  OR2_X1 U7817 ( .A1(n9518), .A2(n9542), .ZN(n9274) );
  NAND2_X1 U7818 ( .A1(n9519), .A2(n9274), .ZN(n9505) );
  OR2_X1 U7819 ( .A1(n9703), .A2(n9521), .ZN(n8978) );
  INV_X1 U7820 ( .A(n9122), .ZN(n9506) );
  NAND2_X1 U7821 ( .A1(n8992), .A2(n9506), .ZN(n6591) );
  NAND2_X1 U7822 ( .A1(n7262), .A2(n6609), .ZN(n9326) );
  NAND2_X1 U7823 ( .A1(n9464), .A2(n9369), .ZN(n6646) );
  INV_X1 U7824 ( .A(n9473), .ZN(n6593) );
  NAND2_X1 U7825 ( .A1(n6594), .A2(n6593), .ZN(n9304) );
  NAND2_X1 U7826 ( .A1(n6267), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6598) );
  NAND2_X1 U7827 ( .A1(n6253), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6597) );
  NAND2_X1 U7828 ( .A1(n6595), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6596) );
  INV_X1 U7829 ( .A(n6600), .ZN(n9366) );
  NAND2_X1 U7830 ( .A1(n9366), .A2(n7577), .ZN(n6602) );
  NAND2_X1 U7831 ( .A1(n6599), .A2(n6602), .ZN(n7301) );
  NOR2_X1 U7832 ( .A1(n8988), .A2(n9685), .ZN(n6604) );
  INV_X1 U7833 ( .A(n7301), .ZN(n7302) );
  INV_X1 U7834 ( .A(n6607), .ZN(n6608) );
  OR2_X1 U7835 ( .A1(n9269), .A2(n6608), .ZN(n7292) );
  NAND3_X1 U7836 ( .A1(n6609), .A2(n9369), .A3(n7976), .ZN(n6610) );
  NAND2_X1 U7837 ( .A1(n9269), .A2(n6610), .ZN(n7637) );
  NAND2_X1 U7838 ( .A1(n7292), .A2(n7637), .ZN(n7639) );
  NAND2_X1 U7839 ( .A1(n6639), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6613) );
  NAND2_X1 U7840 ( .A1(n4969), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6615) );
  INV_X1 U7841 ( .A(n6616), .ZN(n6617) );
  NAND2_X1 U7842 ( .A1(n6617), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6618) );
  INV_X1 U7843 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n7358) );
  NAND2_X1 U7844 ( .A1(n6621), .A2(n7358), .ZN(n6619) );
  NAND2_X1 U7845 ( .A1(n5156), .A2(n8610), .ZN(n7355) );
  OAI21_X1 U7846 ( .B1(n7262), .B2(n8540), .A(n7260), .ZN(n6620) );
  NAND2_X1 U7847 ( .A1(n7639), .A2(n6620), .ZN(n6642) );
  INV_X1 U7848 ( .A(n6621), .ZN(n7353) );
  OAI22_X1 U7849 ( .A1(n7353), .A2(P2_D_REG_1__SCAN_IN), .B1(n6633), .B2(n6632), .ZN(n7636) );
  INV_X1 U7850 ( .A(n7260), .ZN(n7638) );
  NOR2_X1 U7851 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6625) );
  NOR4_X1 U7852 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6624) );
  NOR4_X1 U7853 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6623) );
  NOR4_X1 U7854 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6622) );
  NAND4_X1 U7855 ( .A1(n6625), .A2(n6624), .A3(n6623), .A4(n6622), .ZN(n6631)
         );
  NOR4_X1 U7856 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6629) );
  NOR4_X1 U7857 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6628) );
  NOR4_X1 U7858 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6627) );
  NOR4_X1 U7859 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6626) );
  NAND4_X1 U7860 ( .A1(n6629), .A2(n6628), .A3(n6627), .A4(n6626), .ZN(n6630)
         );
  OAI21_X1 U7861 ( .B1(n6631), .B2(n6630), .A(n6621), .ZN(n6647) );
  INV_X1 U7862 ( .A(n6632), .ZN(n8624) );
  NOR2_X1 U7863 ( .A1(n8624), .A2(n8610), .ZN(n6634) );
  NAND2_X1 U7864 ( .A1(n6634), .A2(n6633), .ZN(n7291) );
  OR2_X1 U7865 ( .A1(n6635), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n6636) );
  NAND2_X1 U7866 ( .A1(n6636), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6637) );
  MUX2_X1 U7867 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6637), .S(
        P2_IR_REG_23__SCAN_IN), .Z(n6638) );
  AND2_X1 U7868 ( .A1(n7296), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7357) );
  AND2_X1 U7869 ( .A1(n6647), .A2(n7354), .ZN(n6640) );
  NAND2_X1 U7870 ( .A1(n7637), .A2(n7636), .ZN(n6641) );
  INV_X1 U7871 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6654) );
  INV_X1 U7872 ( .A(n6644), .ZN(n6645) );
  NAND2_X1 U7873 ( .A1(n6645), .A2(n6647), .ZN(n7289) );
  OR3_X1 U7874 ( .A1(n7262), .A2(n6221), .A3(n6646), .ZN(n7282) );
  AND2_X1 U7875 ( .A1(n7295), .A2(n7282), .ZN(n6652) );
  NAND2_X1 U7876 ( .A1(n7636), .A2(n6647), .ZN(n6648) );
  INV_X1 U7877 ( .A(n7299), .ZN(n6650) );
  NAND3_X1 U7878 ( .A1(n9269), .A2(n7282), .A3(n9773), .ZN(n6649) );
  NAND2_X1 U7879 ( .A1(n9678), .A2(n6649), .ZN(n7281) );
  NAND2_X1 U7880 ( .A1(n6650), .A2(n7281), .ZN(n6651) );
  NAND2_X1 U7881 ( .A1(n6655), .A2(n5560), .ZN(P2_U3455) );
  NAND2_X1 U7882 ( .A1(n6841), .A2(n10030), .ZN(n6656) );
  NAND2_X1 U7883 ( .A1(n6656), .A2(n4961), .ZN(n6657) );
  OAI211_X1 U7884 ( .C1(n10030), .C2(n6841), .A(n6657), .B(n6802), .ZN(n6658)
         );
  NAND2_X1 U7885 ( .A1(n6659), .A2(n6658), .ZN(n6744) );
  NAND2_X1 U7886 ( .A1(n10383), .A2(n10377), .ZN(n6660) );
  AND2_X1 U7887 ( .A1(n8920), .A2(n6660), .ZN(n6840) );
  INV_X1 U7888 ( .A(n6840), .ZN(n6662) );
  NAND2_X1 U7889 ( .A1(n6740), .A2(n6661), .ZN(n6844) );
  MUX2_X1 U7890 ( .A(n6662), .B(n6844), .S(n4963), .Z(n6739) );
  INV_X1 U7891 ( .A(n8900), .ZN(n8904) );
  AND2_X1 U7892 ( .A1(n6810), .A2(n6811), .ZN(n6671) );
  INV_X1 U7893 ( .A(n6663), .ZN(n6664) );
  NAND2_X1 U7894 ( .A1(n8391), .A2(n6664), .ZN(n6665) );
  AND2_X1 U7895 ( .A1(n6665), .A2(n6889), .ZN(n6669) );
  INV_X1 U7896 ( .A(n6666), .ZN(n6893) );
  INV_X1 U7897 ( .A(n6819), .ZN(n6667) );
  AND2_X1 U7898 ( .A1(n6889), .A2(n6667), .ZN(n6668) );
  INV_X1 U7899 ( .A(n6670), .ZN(n8278) );
  NAND2_X1 U7900 ( .A1(n5021), .A2(n6812), .ZN(n6896) );
  NAND3_X1 U7901 ( .A1(n6672), .A2(n6876), .A3(n6879), .ZN(n6673) );
  NAND3_X1 U7902 ( .A1(n6673), .A2(n6881), .A3(n6675), .ZN(n6681) );
  AND2_X1 U7903 ( .A1(n6675), .A2(n6674), .ZN(n6877) );
  OAI21_X1 U7904 ( .B1(n8127), .B2(n8128), .A(n6877), .ZN(n6679) );
  AND2_X1 U7905 ( .A1(n6879), .A2(n6676), .ZN(n6678) );
  INV_X1 U7906 ( .A(n6881), .ZN(n6677) );
  AOI21_X1 U7907 ( .B1(n6679), .B2(n6678), .A(n6677), .ZN(n6680) );
  MUX2_X1 U7908 ( .A(n6681), .B(n6680), .S(n4963), .Z(n6686) );
  NAND2_X1 U7909 ( .A1(n6682), .A2(n6882), .ZN(n6684) );
  AND2_X1 U7910 ( .A1(n6684), .A2(n6683), .ZN(n6885) );
  MUX2_X1 U7911 ( .A(n6882), .B(n6885), .S(n6802), .Z(n6685) );
  OAI211_X1 U7912 ( .C1(n6686), .C2(n8134), .A(n8102), .B(n6685), .ZN(n6687)
         );
  NAND2_X1 U7913 ( .A1(n6687), .A2(n8225), .ZN(n6690) );
  NAND2_X1 U7914 ( .A1(n6688), .A2(n4963), .ZN(n6689) );
  NAND2_X1 U7915 ( .A1(n6690), .A2(n6689), .ZN(n6693) );
  INV_X1 U7916 ( .A(n6884), .ZN(n6817) );
  NAND3_X1 U7917 ( .A1(n6691), .A2(n4963), .A3(n6817), .ZN(n6692) );
  NAND2_X1 U7918 ( .A1(n6693), .A2(n6692), .ZN(n6700) );
  NAND2_X1 U7919 ( .A1(n6700), .A2(n6694), .ZN(n6696) );
  NAND3_X1 U7920 ( .A1(n6696), .A2(n8391), .A3(n6695), .ZN(n6697) );
  NAND2_X1 U7921 ( .A1(n6697), .A2(n4963), .ZN(n6702) );
  NOR2_X1 U7922 ( .A1(n8224), .A2(n4963), .ZN(n6699) );
  INV_X1 U7923 ( .A(n8226), .ZN(n6698) );
  NOR2_X1 U7924 ( .A1(n8231), .A2(n6698), .ZN(n8279) );
  OAI21_X1 U7925 ( .B1(n6700), .B2(n6699), .A(n8279), .ZN(n6701) );
  NAND4_X1 U7926 ( .A1(n6702), .A2(n8281), .A3(n6889), .A4(n6701), .ZN(n6704)
         );
  NAND3_X1 U7927 ( .A1(n6704), .A2(n6703), .A3(n6812), .ZN(n6705) );
  NAND2_X1 U7928 ( .A1(n6706), .A2(n6705), .ZN(n6720) );
  NAND3_X1 U7929 ( .A1(n6720), .A2(n6897), .A3(n5021), .ZN(n6707) );
  AOI21_X1 U7930 ( .B1(n6707), .B2(n6719), .A(n8628), .ZN(n6724) );
  AND2_X1 U7931 ( .A1(n6709), .A2(n6708), .ZN(n6871) );
  NAND3_X1 U7932 ( .A1(n6905), .A2(n4963), .A3(n6871), .ZN(n6723) );
  NAND3_X1 U7933 ( .A1(n10024), .A2(n9925), .A3(n6802), .ZN(n6710) );
  NAND2_X1 U7934 ( .A1(n9935), .A2(n6802), .ZN(n6711) );
  NAND2_X1 U7935 ( .A1(n6710), .A2(n6711), .ZN(n6714) );
  NAND2_X1 U7936 ( .A1(n10032), .A2(n4963), .ZN(n6715) );
  OAI21_X1 U7937 ( .B1(n9925), .B2(n6715), .A(n8899), .ZN(n6713) );
  OAI21_X1 U7938 ( .B1(n10033), .B2(n6711), .A(n10024), .ZN(n6712) );
  AOI22_X1 U7939 ( .A1(n10422), .A2(n6714), .B1(n6713), .B2(n6712), .ZN(n6718)
         );
  OAI21_X1 U7940 ( .B1(n6902), .B2(n6802), .A(n6715), .ZN(n6716) );
  INV_X1 U7941 ( .A(n10422), .ZN(n8653) );
  NAND2_X1 U7942 ( .A1(n6716), .A2(n8653), .ZN(n6717) );
  AND2_X1 U7943 ( .A1(n6718), .A2(n6717), .ZN(n6722) );
  AND2_X1 U7944 ( .A1(n6719), .A2(n6810), .ZN(n6872) );
  NAND2_X1 U7945 ( .A1(n6720), .A2(n6872), .ZN(n6721) );
  NAND2_X1 U7946 ( .A1(n6731), .A2(n6725), .ZN(n6909) );
  OAI211_X1 U7947 ( .C1(n6732), .C2(n6909), .A(n10300), .B(n6916), .ZN(n6726)
         );
  NAND3_X1 U7948 ( .A1(n6726), .A2(n6910), .A3(n10250), .ZN(n6727) );
  NAND2_X1 U7949 ( .A1(n6727), .A2(n6729), .ZN(n6736) );
  NAND2_X1 U7950 ( .A1(n6729), .A2(n6728), .ZN(n6921) );
  INV_X1 U7951 ( .A(n6730), .ZN(n6913) );
  OAI211_X1 U7952 ( .C1(n6913), .C2(n6732), .A(n6731), .B(n6910), .ZN(n6733)
         );
  INV_X1 U7953 ( .A(n6733), .ZN(n6734) );
  OAI21_X1 U7954 ( .B1(n6921), .B2(n6734), .A(n10250), .ZN(n6735) );
  MUX2_X1 U7955 ( .A(n6915), .B(n6737), .S(n6802), .Z(n6738) );
  MUX2_X1 U7956 ( .A(n8920), .B(n6740), .S(n6802), .Z(n6741) );
  NAND4_X1 U7957 ( .A1(n6742), .A2(n8922), .A3(n10185), .A4(n6741), .ZN(n6743)
         );
  NAND2_X1 U7958 ( .A1(n6746), .A2(n6745), .ZN(n6847) );
  NAND2_X1 U7959 ( .A1(n6747), .A2(n6746), .ZN(n6748) );
  MUX2_X1 U7960 ( .A(n6833), .B(n6835), .S(n6802), .Z(n6749) );
  OAI211_X1 U7961 ( .C1(n6751), .C2(n10168), .A(n6750), .B(n6749), .ZN(n6754)
         );
  MUX2_X1 U7962 ( .A(n10345), .B(n10157), .S(n6802), .Z(n6752) );
  NAND2_X1 U7963 ( .A1(n10157), .A2(n10345), .ZN(n10141) );
  NAND2_X1 U7964 ( .A1(n6752), .A2(n10141), .ZN(n6753) );
  NAND2_X1 U7965 ( .A1(n6754), .A2(n6753), .ZN(n6766) );
  NAND2_X1 U7966 ( .A1(n6756), .A2(n6755), .ZN(n6761) );
  INV_X1 U7967 ( .A(n6757), .ZN(n6759) );
  NAND2_X1 U7968 ( .A1(n6759), .A2(n6758), .ZN(n6760) );
  INV_X1 U7969 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n6762) );
  INV_X1 U7970 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10482) );
  MUX2_X1 U7971 ( .A(n6762), .B(n10482), .S(n4964), .Z(n6768) );
  NOR2_X1 U7972 ( .A1(n6787), .A2(n10482), .ZN(n6763) );
  INV_X1 U7973 ( .A(n10152), .ZN(n10346) );
  INV_X1 U7974 ( .A(n10029), .ZN(n6764) );
  NAND2_X1 U7975 ( .A1(n10346), .A2(n6764), .ZN(n6807) );
  NAND2_X1 U7976 ( .A1(n6809), .A2(n6807), .ZN(n10143) );
  MUX2_X1 U7977 ( .A(n6807), .B(n6809), .S(n6802), .Z(n6765) );
  INV_X1 U7978 ( .A(SI_29_), .ZN(n8763) );
  INV_X1 U7979 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n6772) );
  INV_X1 U7980 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8933) );
  MUX2_X1 U7981 ( .A(n6772), .B(n8933), .S(n4965), .Z(n6773) );
  INV_X1 U7982 ( .A(SI_30_), .ZN(n8764) );
  NAND2_X1 U7983 ( .A1(n6773), .A2(n8764), .ZN(n6778) );
  INV_X1 U7984 ( .A(n6773), .ZN(n6774) );
  NAND2_X1 U7985 ( .A1(n6774), .A2(SI_30_), .ZN(n6775) );
  NAND2_X1 U7986 ( .A1(n6778), .A2(n6775), .ZN(n6779) );
  NAND2_X1 U7987 ( .A1(n9289), .A2(n6785), .ZN(n6777) );
  OR2_X1 U7988 ( .A1(n6787), .A2(n8933), .ZN(n6776) );
  INV_X1 U7989 ( .A(n10439), .ZN(n6804) );
  MUX2_X1 U7990 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n4965), .Z(n6782) );
  INV_X1 U7991 ( .A(SI_31_), .ZN(n6781) );
  XNOR2_X1 U7992 ( .A(n6782), .B(n6781), .ZN(n6783) );
  NAND2_X1 U7993 ( .A1(n9835), .A2(n6785), .ZN(n6789) );
  INV_X1 U7994 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6786) );
  OR2_X1 U7995 ( .A1(n6787), .A2(n6786), .ZN(n6788) );
  NAND2_X1 U7996 ( .A1(n5654), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6792) );
  NAND2_X1 U7997 ( .A1(n4958), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6791) );
  NAND2_X1 U7998 ( .A1(n5652), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6790) );
  OR2_X2 U7999 ( .A1(n6794), .A2(n6804), .ZN(n6799) );
  NAND2_X1 U8000 ( .A1(n5654), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6797) );
  NAND2_X1 U8001 ( .A1(n5631), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6796) );
  NAND2_X1 U8002 ( .A1(n5652), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6795) );
  AND3_X1 U8003 ( .A1(n6797), .A2(n6796), .A3(n6795), .ZN(n10127) );
  INV_X1 U8004 ( .A(n10127), .ZN(n10028) );
  INV_X1 U8005 ( .A(n6930), .ZN(n6800) );
  AND2_X1 U8006 ( .A1(n6852), .A2(n10127), .ZN(n6805) );
  INV_X1 U8007 ( .A(n6805), .ZN(n6854) );
  INV_X1 U8008 ( .A(n6117), .ZN(n8221) );
  NOR2_X1 U8009 ( .A1(n6804), .A2(n6806), .ZN(n6853) );
  NOR2_X1 U8010 ( .A1(n6805), .A2(n6853), .ZN(n6929) );
  NAND2_X1 U8011 ( .A1(n6808), .A2(n6807), .ZN(n6926) );
  NAND2_X1 U8012 ( .A1(n5021), .A2(n6810), .ZN(n8473) );
  NAND2_X1 U8013 ( .A1(n6812), .A2(n6811), .ZN(n8394) );
  INV_X1 U8014 ( .A(n6813), .ZN(n8079) );
  NAND2_X1 U8015 ( .A1(n6960), .A2(n8075), .ZN(n6874) );
  NAND2_X1 U8016 ( .A1(n8079), .A2(n6874), .ZN(n8012) );
  NOR2_X1 U8017 ( .A1(n8012), .A2(n6117), .ZN(n6816) );
  NAND4_X1 U8018 ( .A1(n6816), .A2(n8140), .A3(n6815), .A4(n6814), .ZN(n6818)
         );
  NAND4_X1 U8019 ( .A1(n8261), .A2(n6821), .A3(n6820), .A4(n6819), .ZN(n6822)
         );
  NOR4_X1 U8020 ( .A1(n8473), .A2(n8394), .A3(n6823), .A4(n6822), .ZN(n6824)
         );
  NAND4_X1 U8021 ( .A1(n8617), .A2(n5263), .A3(n8509), .A4(n6824), .ZN(n6825)
         );
  NOR4_X1 U8022 ( .A1(n5952), .A2(n8900), .A3(n8648), .A4(n6825), .ZN(n6826)
         );
  XNOR2_X1 U8023 ( .A(n10324), .B(n10031), .ZN(n10320) );
  NAND4_X1 U8024 ( .A1(n10252), .A2(n10279), .A3(n6826), .A4(n10320), .ZN(
        n6827) );
  NOR4_X1 U8025 ( .A1(n10201), .A2(n6828), .A3(n10225), .A4(n6827), .ZN(n6829)
         );
  NAND4_X1 U8026 ( .A1(n10171), .A2(n8922), .A3(n10190), .A4(n6829), .ZN(n6830) );
  NOR4_X1 U8027 ( .A1(n6926), .A2(n6838), .A3(n6831), .A4(n6830), .ZN(n6832)
         );
  NAND3_X1 U8028 ( .A1(n6929), .A2(n6832), .A3(n6930), .ZN(n6856) );
  OAI211_X1 U8029 ( .C1(n6947), .C2(n8221), .A(n6856), .B(n4966), .ZN(n6868)
         );
  NAND2_X1 U8030 ( .A1(n10135), .A2(n6833), .ZN(n6848) );
  AOI21_X1 U8031 ( .B1(n6835), .B2(n6834), .A(n6848), .ZN(n6836) );
  NOR3_X1 U8032 ( .A1(n6838), .A2(n6837), .A3(n6836), .ZN(n6928) );
  NAND3_X1 U8033 ( .A1(n6841), .A2(n6840), .A3(n6839), .ZN(n6918) );
  NOR2_X1 U8034 ( .A1(n6918), .A2(n6842), .ZN(n6849) );
  AOI21_X1 U8035 ( .B1(n8920), .B2(n6844), .A(n6843), .ZN(n6846) );
  OAI21_X1 U8036 ( .B1(n6846), .B2(n6845), .A(n10185), .ZN(n6924) );
  NOR2_X1 U8037 ( .A1(n6848), .A2(n6847), .ZN(n6923) );
  OAI21_X1 U8038 ( .B1(n6849), .B2(n6924), .A(n6923), .ZN(n6851) );
  AOI21_X1 U8039 ( .B1(n10127), .B2(n10439), .A(n6852), .ZN(n6850) );
  AOI211_X1 U8040 ( .C1(n6928), .C2(n6851), .A(n6926), .B(n6850), .ZN(n6858)
         );
  INV_X1 U8041 ( .A(n6853), .ZN(n6855) );
  OAI211_X1 U8042 ( .C1(n10435), .C2(n6855), .A(n7315), .B(n6854), .ZN(n6857)
         );
  OAI21_X1 U8043 ( .B1(n6858), .B2(n6857), .A(n6856), .ZN(n6866) );
  NOR2_X1 U8044 ( .A1(n8014), .A2(n6950), .ZN(n6859) );
  NAND2_X1 U8045 ( .A1(n7750), .A2(n6859), .ZN(n7192) );
  AND2_X1 U8046 ( .A1(n6861), .A2(n6860), .ZN(n10124) );
  NAND2_X1 U8047 ( .A1(n7321), .A2(n10124), .ZN(n10554) );
  OR2_X1 U8048 ( .A1(n7192), .A2(n10554), .ZN(n6865) );
  INV_X1 U8049 ( .A(n7319), .ZN(n6862) );
  AND2_X1 U8050 ( .A1(n6862), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6937) );
  INV_X1 U8051 ( .A(P1_B_REG_SCAN_IN), .ZN(n6863) );
  AOI21_X1 U8052 ( .B1(n6937), .B2(n8501), .A(n6863), .ZN(n6864) );
  AND2_X1 U8053 ( .A1(n6865), .A2(n6864), .ZN(n6933) );
  AOI211_X1 U8054 ( .C1(n6866), .C2(n10116), .A(n6933), .B(n8218), .ZN(n6867)
         );
  OAI21_X1 U8055 ( .B1(n6870), .B2(n6868), .A(n6867), .ZN(n6869) );
  INV_X1 U8056 ( .A(n6869), .ZN(n6944) );
  OAI211_X1 U8057 ( .C1(n10116), .C2(n6930), .A(n6870), .B(n8501), .ZN(n6943)
         );
  INV_X1 U8058 ( .A(n6910), .ZN(n6917) );
  INV_X1 U8059 ( .A(n6871), .ZN(n6904) );
  INV_X1 U8060 ( .A(n6872), .ZN(n6900) );
  NAND2_X1 U8061 ( .A1(n10044), .A2(n8076), .ZN(n6873) );
  NAND3_X1 U8062 ( .A1(n6874), .A2(n6117), .A3(n6873), .ZN(n6875) );
  NAND2_X1 U8063 ( .A1(n6876), .A2(n6875), .ZN(n6878) );
  OAI21_X1 U8064 ( .B1(n8127), .B2(n6878), .A(n6877), .ZN(n6880) );
  NAND2_X1 U8065 ( .A1(n6880), .A2(n6879), .ZN(n6883) );
  NAND3_X1 U8066 ( .A1(n6883), .A2(n6882), .A3(n6881), .ZN(n6886) );
  NAND3_X1 U8067 ( .A1(n6886), .A2(n6885), .A3(n6884), .ZN(n6887) );
  NAND2_X1 U8068 ( .A1(n6888), .A2(n6887), .ZN(n6892) );
  INV_X1 U8069 ( .A(n6889), .ZN(n6890) );
  AOI21_X1 U8070 ( .B1(n6892), .B2(n6891), .A(n6890), .ZN(n6894) );
  NOR2_X1 U8071 ( .A1(n6894), .A2(n6893), .ZN(n6895) );
  NOR2_X1 U8072 ( .A1(n6896), .A2(n6895), .ZN(n6899) );
  OAI211_X1 U8073 ( .C1(n6900), .C2(n6899), .A(n6898), .B(n6897), .ZN(n6901)
         );
  INV_X1 U8074 ( .A(n6901), .ZN(n6903) );
  OAI21_X1 U8075 ( .B1(n6904), .B2(n6903), .A(n6902), .ZN(n6906) );
  NAND2_X1 U8076 ( .A1(n6906), .A2(n6905), .ZN(n6908) );
  NAND2_X1 U8077 ( .A1(n6908), .A2(n6907), .ZN(n6912) );
  INV_X1 U8078 ( .A(n6909), .ZN(n6911) );
  OAI211_X1 U8079 ( .C1(n6913), .C2(n6912), .A(n6911), .B(n6910), .ZN(n6914)
         );
  OAI211_X1 U8080 ( .C1(n6917), .C2(n6916), .A(n6915), .B(n6914), .ZN(n6920)
         );
  INV_X1 U8081 ( .A(n6918), .ZN(n6919) );
  OAI21_X1 U8082 ( .B1(n6921), .B2(n6920), .A(n6919), .ZN(n6922) );
  INV_X1 U8083 ( .A(n6922), .ZN(n6925) );
  OAI21_X1 U8084 ( .B1(n6925), .B2(n6924), .A(n6923), .ZN(n6927) );
  AOI21_X1 U8085 ( .B1(n6928), .B2(n6927), .A(n6926), .ZN(n6932) );
  INV_X1 U8086 ( .A(n6929), .ZN(n6931) );
  OAI21_X1 U8087 ( .B1(n6932), .B2(n6931), .A(n6930), .ZN(n6936) );
  INV_X1 U8088 ( .A(n6936), .ZN(n6935) );
  INV_X1 U8089 ( .A(n6933), .ZN(n6938) );
  NAND3_X1 U8090 ( .A1(n6935), .A2(n6934), .A3(n6938), .ZN(n6941) );
  NAND4_X1 U8091 ( .A1(n6936), .A2(n8218), .A3(n4966), .A4(n6938), .ZN(n6940)
         );
  INV_X1 U8092 ( .A(n6937), .ZN(n8525) );
  NAND2_X1 U8093 ( .A1(n6938), .A2(n8525), .ZN(n6939) );
  NAND3_X1 U8094 ( .A1(n6941), .A2(n6940), .A3(n6939), .ZN(n6942) );
  AOI21_X1 U8095 ( .B1(n6944), .B2(n6943), .A(n6942), .ZN(P1_U3242) );
  INV_X1 U8096 ( .A(n6950), .ZN(n8019) );
  AND2_X1 U8097 ( .A1(n6950), .A2(n6949), .ZN(n6951) );
  XNOR2_X1 U8098 ( .A(n6952), .B(n7163), .ZN(n6980) );
  OR2_X1 U8099 ( .A1(n8088), .A2(n7165), .ZN(n6954) );
  NAND2_X1 U8100 ( .A1(n6954), .A2(n6953), .ZN(n6978) );
  XNOR2_X1 U8101 ( .A(n6980), .B(n6978), .ZN(n7756) );
  NAND2_X1 U8102 ( .A1(n6960), .A2(n7001), .ZN(n6956) );
  NAND2_X1 U8103 ( .A1(n6966), .A2(n8010), .ZN(n6955) );
  INV_X1 U8104 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6957) );
  NAND2_X1 U8105 ( .A1(n6960), .A2(n7173), .ZN(n6963) );
  OAI22_X1 U8106 ( .A1(n8075), .A2(n7028), .B1(n10557), .B2(n6949), .ZN(n6961)
         );
  INV_X1 U8107 ( .A(n6961), .ZN(n6962) );
  NAND2_X1 U8108 ( .A1(n6963), .A2(n6962), .ZN(n7311) );
  NAND2_X1 U8109 ( .A1(n7312), .A2(n7311), .ZN(n7310) );
  NAND2_X1 U8110 ( .A1(n6964), .A2(n7163), .ZN(n6965) );
  NAND2_X1 U8111 ( .A1(n10044), .A2(n7001), .ZN(n6969) );
  NAND2_X1 U8112 ( .A1(n6966), .A2(n6967), .ZN(n6968) );
  NAND2_X1 U8113 ( .A1(n6969), .A2(n6968), .ZN(n6971) );
  NAND2_X1 U8114 ( .A1(n6973), .A2(n6974), .ZN(n7760) );
  AND2_X1 U8115 ( .A1(n6967), .A2(n7001), .ZN(n6972) );
  AOI21_X1 U8116 ( .B1(n10044), .B2(n7173), .A(n6972), .ZN(n7761) );
  NAND2_X1 U8117 ( .A1(n7760), .A2(n7761), .ZN(n6977) );
  INV_X1 U8118 ( .A(n6974), .ZN(n6975) );
  NAND2_X1 U8119 ( .A1(n7756), .A2(n7755), .ZN(n6982) );
  INV_X1 U8120 ( .A(n6978), .ZN(n6979) );
  NAND2_X1 U8121 ( .A1(n6980), .A2(n6979), .ZN(n6981) );
  NAND2_X1 U8122 ( .A1(n6982), .A2(n6981), .ZN(n7850) );
  XNOR2_X1 U8123 ( .A(n6984), .B(n7163), .ZN(n6989) );
  OR2_X1 U8124 ( .A1(n8129), .A2(n7165), .ZN(n6986) );
  NAND2_X1 U8125 ( .A1(n8347), .A2(n7150), .ZN(n6985) );
  NAND2_X1 U8126 ( .A1(n6986), .A2(n6985), .ZN(n6987) );
  XNOR2_X1 U8127 ( .A(n6989), .B(n6987), .ZN(n7851) );
  NAND2_X1 U8128 ( .A1(n7850), .A2(n7851), .ZN(n6991) );
  INV_X1 U8129 ( .A(n6987), .ZN(n6988) );
  NAND2_X1 U8130 ( .A1(n6989), .A2(n6988), .ZN(n6990) );
  NAND2_X1 U8131 ( .A1(n6991), .A2(n6990), .ZN(n7855) );
  NAND2_X1 U8132 ( .A1(n10041), .A2(n7150), .ZN(n6993) );
  INV_X1 U8133 ( .A(n10784), .ZN(n6995) );
  NAND2_X1 U8134 ( .A1(n6995), .A2(n6966), .ZN(n6992) );
  NAND2_X1 U8135 ( .A1(n6993), .A2(n6992), .ZN(n6994) );
  XNOR2_X1 U8136 ( .A(n6994), .B(n7163), .ZN(n6996) );
  AOI22_X1 U8137 ( .A1(n10041), .A2(n7173), .B1(n7150), .B2(n6995), .ZN(n6997)
         );
  XNOR2_X1 U8138 ( .A(n6996), .B(n6997), .ZN(n7856) );
  INV_X1 U8139 ( .A(n6996), .ZN(n6999) );
  INV_X1 U8140 ( .A(n6997), .ZN(n6998) );
  NAND2_X1 U8141 ( .A1(n6999), .A2(n6998), .ZN(n7000) );
  OAI22_X1 U8142 ( .A1(n8107), .A2(n7179), .B1(n7890), .B2(n6983), .ZN(n7002)
         );
  XNOR2_X1 U8143 ( .A(n7002), .B(n7176), .ZN(n7006) );
  OR2_X1 U8144 ( .A1(n8107), .A2(n7165), .ZN(n7004) );
  NAND2_X1 U8145 ( .A1(n8172), .A2(n7150), .ZN(n7003) );
  AND2_X1 U8146 ( .A1(n7004), .A2(n7003), .ZN(n7888) );
  NAND2_X1 U8147 ( .A1(n7886), .A2(n7888), .ZN(n7009) );
  INV_X1 U8148 ( .A(n7005), .ZN(n7008) );
  INV_X1 U8149 ( .A(n7006), .ZN(n7007) );
  NAND2_X1 U8150 ( .A1(n7008), .A2(n7007), .ZN(n7887) );
  NAND2_X1 U8151 ( .A1(n8114), .A2(n6966), .ZN(n7010) );
  OAI21_X1 U8152 ( .B1(n8243), .B2(n7179), .A(n7010), .ZN(n7011) );
  XNOR2_X1 U8153 ( .A(n7011), .B(n7163), .ZN(n7016) );
  OR2_X1 U8154 ( .A1(n8243), .A2(n7165), .ZN(n7013) );
  NAND2_X1 U8155 ( .A1(n8114), .A2(n7150), .ZN(n7012) );
  NAND2_X1 U8156 ( .A1(n7013), .A2(n7012), .ZN(n7014) );
  XNOR2_X1 U8157 ( .A(n7016), .B(n7014), .ZN(n7952) );
  INV_X1 U8158 ( .A(n7014), .ZN(n7015) );
  NAND2_X1 U8159 ( .A1(n7016), .A2(n7015), .ZN(n7017) );
  OAI22_X1 U8160 ( .A1(n8370), .A2(n6983), .B1(n8229), .B2(n7179), .ZN(n7018)
         );
  XNOR2_X1 U8161 ( .A(n7018), .B(n7163), .ZN(n7023) );
  OR2_X1 U8162 ( .A1(n8370), .A2(n7179), .ZN(n7020) );
  NAND2_X1 U8163 ( .A1(n10038), .A2(n7173), .ZN(n7019) );
  NAND2_X1 U8164 ( .A1(n7020), .A2(n7019), .ZN(n7021) );
  XNOR2_X1 U8165 ( .A(n7023), .B(n7021), .ZN(n8060) );
  INV_X1 U8166 ( .A(n7021), .ZN(n7022) );
  NAND2_X1 U8167 ( .A1(n7023), .A2(n7022), .ZN(n7024) );
  NAND2_X1 U8168 ( .A1(n8234), .A2(n6966), .ZN(n7026) );
  OR2_X1 U8169 ( .A1(n8385), .A2(n7179), .ZN(n7025) );
  NAND2_X1 U8170 ( .A1(n7026), .A2(n7025), .ZN(n7027) );
  XNOR2_X1 U8171 ( .A(n7027), .B(n7163), .ZN(n7030) );
  NOR2_X1 U8172 ( .A1(n8385), .A2(n7165), .ZN(n7029) );
  AOI21_X1 U8173 ( .B1(n8234), .B2(n7150), .A(n7029), .ZN(n8358) );
  NAND2_X1 U8174 ( .A1(n8288), .A2(n6966), .ZN(n7033) );
  OR2_X1 U8175 ( .A1(n8494), .A2(n7028), .ZN(n7032) );
  NAND2_X1 U8176 ( .A1(n7033), .A2(n7032), .ZN(n7034) );
  XNOR2_X1 U8177 ( .A(n7034), .B(n7163), .ZN(n7036) );
  NOR2_X1 U8178 ( .A1(n8494), .A2(n7165), .ZN(n7035) );
  AOI21_X1 U8179 ( .B1(n8288), .B2(n7150), .A(n7035), .ZN(n7037) );
  AND2_X1 U8180 ( .A1(n7036), .A2(n7037), .ZN(n8377) );
  INV_X1 U8181 ( .A(n7036), .ZN(n7039) );
  INV_X1 U8182 ( .A(n7037), .ZN(n7038) );
  NAND2_X1 U8183 ( .A1(n7039), .A2(n7038), .ZN(n8378) );
  NAND2_X1 U8184 ( .A1(n8269), .A2(n7150), .ZN(n7041) );
  OR2_X1 U8185 ( .A1(n8431), .A2(n7165), .ZN(n7040) );
  NAND2_X1 U8186 ( .A1(n7041), .A2(n7040), .ZN(n8489) );
  NAND2_X1 U8187 ( .A1(n8269), .A2(n6966), .ZN(n7043) );
  OR2_X1 U8188 ( .A1(n8431), .A2(n7179), .ZN(n7042) );
  NAND2_X1 U8189 ( .A1(n7043), .A2(n7042), .ZN(n7044) );
  XNOR2_X1 U8190 ( .A(n7044), .B(n7176), .ZN(n8488) );
  NAND2_X1 U8191 ( .A1(n8572), .A2(n6966), .ZN(n7046) );
  OR2_X1 U8192 ( .A1(n8469), .A2(n7179), .ZN(n7045) );
  NAND2_X1 U8193 ( .A1(n7046), .A2(n7045), .ZN(n7047) );
  XNOR2_X1 U8194 ( .A(n7047), .B(n7163), .ZN(n7050) );
  NOR2_X1 U8195 ( .A1(n8469), .A2(n7165), .ZN(n7048) );
  AOI21_X1 U8196 ( .B1(n8572), .B2(n7150), .A(n7048), .ZN(n7049) );
  NAND2_X1 U8197 ( .A1(n7050), .A2(n7049), .ZN(n8562) );
  OR2_X1 U8198 ( .A1(n7050), .A2(n7049), .ZN(n8563) );
  OAI22_X1 U8199 ( .A1(n10836), .A2(n6983), .B1(n8570), .B2(n7179), .ZN(n7052)
         );
  XNOR2_X1 U8200 ( .A(n7052), .B(n7176), .ZN(n7056) );
  OR2_X1 U8201 ( .A1(n10836), .A2(n7179), .ZN(n7054) );
  NAND2_X1 U8202 ( .A1(n10035), .A2(n7173), .ZN(n7053) );
  NAND2_X1 U8203 ( .A1(n7054), .A2(n7053), .ZN(n7057) );
  XNOR2_X1 U8204 ( .A(n7056), .B(n7057), .ZN(n9899) );
  INV_X1 U8205 ( .A(n7056), .ZN(n7059) );
  INV_X1 U8206 ( .A(n7057), .ZN(n7058) );
  NAND2_X1 U8207 ( .A1(n7059), .A2(n7058), .ZN(n7060) );
  NAND2_X1 U8208 ( .A1(n8516), .A2(n6966), .ZN(n7062) );
  OR2_X1 U8209 ( .A1(n9904), .A2(n7179), .ZN(n7061) );
  NAND2_X1 U8210 ( .A1(n7062), .A2(n7061), .ZN(n7063) );
  XNOR2_X1 U8211 ( .A(n7063), .B(n7163), .ZN(n7066) );
  NOR2_X1 U8212 ( .A1(n9904), .A2(n7165), .ZN(n7064) );
  AOI21_X1 U8213 ( .B1(n8516), .B2(n7150), .A(n7064), .ZN(n7065) );
  XNOR2_X1 U8214 ( .A(n7066), .B(n7065), .ZN(n9965) );
  NAND2_X1 U8215 ( .A1(n10427), .A2(n6966), .ZN(n7068) );
  OR2_X1 U8216 ( .A1(n10021), .A2(n7179), .ZN(n7067) );
  NAND2_X1 U8217 ( .A1(n7068), .A2(n7067), .ZN(n7069) );
  XNOR2_X1 U8218 ( .A(n7069), .B(n7163), .ZN(n7073) );
  NAND2_X1 U8219 ( .A1(n10427), .A2(n7150), .ZN(n7071) );
  OR2_X1 U8220 ( .A1(n10021), .A2(n7165), .ZN(n7070) );
  NAND2_X1 U8221 ( .A1(n7071), .A2(n7070), .ZN(n9861) );
  NAND2_X1 U8222 ( .A1(n9858), .A2(n9861), .ZN(n7076) );
  INV_X1 U8223 ( .A(n7072), .ZN(n7075) );
  INV_X1 U8224 ( .A(n7073), .ZN(n7074) );
  NAND2_X1 U8225 ( .A1(n7075), .A2(n7074), .ZN(n9859) );
  AND2_X2 U8226 ( .A1(n7076), .A2(n9859), .ZN(n7078) );
  OAI22_X1 U8227 ( .A1(n8899), .A2(n6983), .B1(n9925), .B2(n7179), .ZN(n7077)
         );
  XNOR2_X1 U8228 ( .A(n7077), .B(n7163), .ZN(n7079) );
  OAI22_X1 U8229 ( .A1(n8899), .A2(n7179), .B1(n9925), .B2(n7165), .ZN(n10013)
         );
  INV_X1 U8230 ( .A(n7078), .ZN(n7081) );
  INV_X1 U8231 ( .A(n7079), .ZN(n7080) );
  NAND2_X1 U8232 ( .A1(n10422), .A2(n6966), .ZN(n7083) );
  OR2_X1 U8233 ( .A1(n9935), .A2(n7179), .ZN(n7082) );
  NAND2_X1 U8234 ( .A1(n7083), .A2(n7082), .ZN(n7084) );
  XNOR2_X1 U8235 ( .A(n7084), .B(n7163), .ZN(n7087) );
  NOR2_X1 U8236 ( .A1(n9935), .A2(n7165), .ZN(n7085) );
  AOI21_X1 U8237 ( .B1(n10422), .B2(n7150), .A(n7085), .ZN(n7086) );
  XNOR2_X1 U8238 ( .A(n7087), .B(n7086), .ZN(n9920) );
  NAND2_X1 U8239 ( .A1(n7087), .A2(n7086), .ZN(n7088) );
  NAND2_X1 U8240 ( .A1(n8908), .A2(n6966), .ZN(n7090) );
  OR2_X1 U8241 ( .A1(n10314), .A2(n7179), .ZN(n7089) );
  NAND2_X1 U8242 ( .A1(n7090), .A2(n7089), .ZN(n7091) );
  XNOR2_X1 U8243 ( .A(n7091), .B(n7163), .ZN(n9930) );
  NOR2_X1 U8244 ( .A1(n10314), .A2(n7165), .ZN(n7092) );
  AOI21_X1 U8245 ( .B1(n8908), .B2(n7150), .A(n7092), .ZN(n9929) );
  AND2_X1 U8246 ( .A1(n9930), .A2(n9929), .ZN(n7094) );
  NAND2_X1 U8247 ( .A1(n10324), .A2(n7150), .ZN(n7096) );
  NAND2_X1 U8248 ( .A1(n10031), .A2(n7173), .ZN(n7095) );
  NAND2_X1 U8249 ( .A1(n7096), .A2(n7095), .ZN(n9988) );
  NAND2_X1 U8250 ( .A1(n10324), .A2(n6966), .ZN(n7098) );
  NAND2_X1 U8251 ( .A1(n10031), .A2(n7150), .ZN(n7097) );
  NAND2_X1 U8252 ( .A1(n7098), .A2(n7097), .ZN(n7099) );
  XNOR2_X1 U8253 ( .A(n7099), .B(n7176), .ZN(n9987) );
  NAND2_X1 U8254 ( .A1(n10296), .A2(n6966), .ZN(n7101) );
  NAND2_X1 U8255 ( .A1(n7604), .A2(n7150), .ZN(n7100) );
  NAND2_X1 U8256 ( .A1(n7101), .A2(n7100), .ZN(n7102) );
  XNOR2_X1 U8257 ( .A(n7102), .B(n7163), .ZN(n7105) );
  NOR2_X1 U8258 ( .A1(n10396), .A2(n7165), .ZN(n7103) );
  AOI21_X1 U8259 ( .B1(n10296), .B2(n7150), .A(n7103), .ZN(n7104) );
  NAND2_X1 U8260 ( .A1(n7105), .A2(n7104), .ZN(n9954) );
  OR2_X1 U8261 ( .A1(n7105), .A2(n7104), .ZN(n7106) );
  NAND2_X1 U8262 ( .A1(n9954), .A2(n7106), .ZN(n9881) );
  INV_X1 U8263 ( .A(n9881), .ZN(n7107) );
  NAND2_X1 U8264 ( .A1(n9879), .A2(n9954), .ZN(n7115) );
  NAND2_X1 U8265 ( .A1(n10273), .A2(n6966), .ZN(n7109) );
  OR2_X1 U8266 ( .A1(n10302), .A2(n7179), .ZN(n7108) );
  NAND2_X1 U8267 ( .A1(n7109), .A2(n7108), .ZN(n7110) );
  XNOR2_X1 U8268 ( .A(n7110), .B(n7163), .ZN(n7113) );
  NOR2_X1 U8269 ( .A1(n10302), .A2(n7165), .ZN(n7111) );
  AOI21_X1 U8270 ( .B1(n10273), .B2(n7150), .A(n7111), .ZN(n7112) );
  NAND2_X1 U8271 ( .A1(n7113), .A2(n7112), .ZN(n7116) );
  OR2_X1 U8272 ( .A1(n7113), .A2(n7112), .ZN(n7114) );
  AND2_X1 U8273 ( .A1(n7116), .A2(n7114), .ZN(n9955) );
  NAND2_X1 U8274 ( .A1(n9958), .A2(n7116), .ZN(n9888) );
  NAND2_X1 U8275 ( .A1(n10390), .A2(n6966), .ZN(n7118) );
  NAND2_X1 U8276 ( .A1(n10281), .A2(n7150), .ZN(n7117) );
  NAND2_X1 U8277 ( .A1(n7118), .A2(n7117), .ZN(n7119) );
  XNOR2_X1 U8278 ( .A(n7119), .B(n7176), .ZN(n7122) );
  NOR2_X1 U8279 ( .A1(n7120), .A2(n7165), .ZN(n7121) );
  AOI21_X1 U8280 ( .B1(n10390), .B2(n7150), .A(n7121), .ZN(n7123) );
  XNOR2_X1 U8281 ( .A(n7122), .B(n7123), .ZN(n9889) );
  NAND2_X1 U8282 ( .A1(n9888), .A2(n9889), .ZN(n9887) );
  INV_X1 U8283 ( .A(n7122), .ZN(n7124) );
  NAND2_X1 U8284 ( .A1(n7124), .A2(n7123), .ZN(n7125) );
  NAND2_X1 U8285 ( .A1(n9887), .A2(n7125), .ZN(n9870) );
  NAND2_X1 U8286 ( .A1(n10234), .A2(n6966), .ZN(n7127) );
  NAND2_X1 U8287 ( .A1(n10245), .A2(n7150), .ZN(n7126) );
  NAND2_X1 U8288 ( .A1(n7127), .A2(n7126), .ZN(n7128) );
  XNOR2_X1 U8289 ( .A(n7128), .B(n7176), .ZN(n7138) );
  NAND2_X1 U8290 ( .A1(n10234), .A2(n7150), .ZN(n7130) );
  NAND2_X1 U8291 ( .A1(n10245), .A2(n7173), .ZN(n7129) );
  NAND2_X1 U8292 ( .A1(n7130), .A2(n7129), .ZN(n7139) );
  NAND2_X1 U8293 ( .A1(n7138), .A2(n7139), .ZN(n9871) );
  INV_X1 U8294 ( .A(n9871), .ZN(n7136) );
  NAND2_X1 U8295 ( .A1(n10383), .A2(n6966), .ZN(n7132) );
  OR2_X1 U8296 ( .A1(n10377), .A2(n7179), .ZN(n7131) );
  NAND2_X1 U8297 ( .A1(n7132), .A2(n7131), .ZN(n7133) );
  XNOR2_X1 U8298 ( .A(n7133), .B(n7163), .ZN(n9869) );
  NOR2_X1 U8299 ( .A1(n10377), .A2(n7165), .ZN(n7134) );
  AOI21_X1 U8300 ( .B1(n10383), .B2(n7150), .A(n7134), .ZN(n9977) );
  NAND2_X1 U8301 ( .A1(n9870), .A2(n7137), .ZN(n7148) );
  NAND3_X1 U8302 ( .A1(n9871), .A2(n9977), .A3(n9869), .ZN(n7142) );
  INV_X1 U8303 ( .A(n7138), .ZN(n7141) );
  INV_X1 U8304 ( .A(n7139), .ZN(n7140) );
  NAND2_X1 U8305 ( .A1(n7141), .A2(n7140), .ZN(n9941) );
  AOI22_X1 U8306 ( .A1(n10372), .A2(n6966), .B1(n7150), .B2(n10205), .ZN(n7143) );
  XOR2_X1 U8307 ( .A(n7176), .B(n7143), .Z(n7145) );
  OAI22_X1 U8308 ( .A1(n9953), .A2(n7179), .B1(n10222), .B2(n7165), .ZN(n7144)
         );
  NOR2_X1 U8309 ( .A1(n7145), .A2(n7144), .ZN(n7149) );
  AOI21_X1 U8310 ( .B1(n7145), .B2(n7144), .A(n7149), .ZN(n9942) );
  INV_X1 U8311 ( .A(n9942), .ZN(n7146) );
  AOI21_X2 U8312 ( .B1(n7148), .B2(n7147), .A(n7146), .ZN(n9945) );
  AOI22_X1 U8313 ( .A1(n4961), .A2(n7150), .B1(n7173), .B2(n10030), .ZN(n7158)
         );
  NAND2_X1 U8314 ( .A1(n4961), .A2(n6966), .ZN(n7152) );
  NAND2_X1 U8315 ( .A1(n10030), .A2(n7150), .ZN(n7151) );
  NAND2_X1 U8316 ( .A1(n7152), .A2(n7151), .ZN(n7153) );
  XNOR2_X1 U8317 ( .A(n7153), .B(n7176), .ZN(n7160) );
  XOR2_X1 U8318 ( .A(n7158), .B(n7160), .Z(n9909) );
  NAND2_X1 U8319 ( .A1(n10198), .A2(n6966), .ZN(n7155) );
  NAND2_X1 U8320 ( .A1(n7768), .A2(n7150), .ZN(n7154) );
  NAND2_X1 U8321 ( .A1(n7155), .A2(n7154), .ZN(n7156) );
  XNOR2_X1 U8322 ( .A(n7156), .B(n7163), .ZN(n7169) );
  NOR2_X1 U8323 ( .A1(n10208), .A2(n7165), .ZN(n7157) );
  AOI21_X1 U8324 ( .B1(n10198), .B2(n7150), .A(n7157), .ZN(n7170) );
  XNOR2_X1 U8325 ( .A(n7169), .B(n7170), .ZN(n9998) );
  INV_X1 U8326 ( .A(n7158), .ZN(n7159) );
  NOR2_X1 U8327 ( .A1(n7160), .A2(n7159), .ZN(n9999) );
  NAND2_X1 U8328 ( .A1(n10177), .A2(n6966), .ZN(n7162) );
  OR2_X1 U8329 ( .A1(n7203), .A2(n7179), .ZN(n7161) );
  NAND2_X1 U8330 ( .A1(n7162), .A2(n7161), .ZN(n7164) );
  XNOR2_X1 U8331 ( .A(n7164), .B(n7163), .ZN(n7168) );
  NOR2_X1 U8332 ( .A1(n7203), .A2(n7165), .ZN(n7166) );
  AOI21_X1 U8333 ( .B1(n10177), .B2(n7150), .A(n7166), .ZN(n7167) );
  NAND2_X1 U8334 ( .A1(n7168), .A2(n7167), .ZN(n7204) );
  OAI21_X1 U8335 ( .B1(n7168), .B2(n7167), .A(n7204), .ZN(n7211) );
  INV_X1 U8336 ( .A(n7169), .ZN(n7172) );
  INV_X1 U8337 ( .A(n7170), .ZN(n7171) );
  NAND2_X1 U8338 ( .A1(n10157), .A2(n7150), .ZN(n7175) );
  NAND2_X1 U8339 ( .A1(n10345), .A2(n7173), .ZN(n7174) );
  NAND2_X1 U8340 ( .A1(n7175), .A2(n7174), .ZN(n7177) );
  XNOR2_X1 U8341 ( .A(n7177), .B(n7176), .ZN(n7181) );
  NAND2_X1 U8342 ( .A1(n10157), .A2(n6966), .ZN(n7178) );
  OAI21_X1 U8343 ( .B1(n10172), .B2(n7179), .A(n7178), .ZN(n7180) );
  XNOR2_X1 U8344 ( .A(n7181), .B(n7180), .ZN(n7205) );
  INV_X1 U8345 ( .A(n7182), .ZN(n7932) );
  NAND3_X1 U8346 ( .A1(n7184), .A2(n7932), .A3(n7183), .ZN(n7199) );
  INV_X1 U8347 ( .A(n7750), .ZN(n7188) );
  OR2_X1 U8348 ( .A1(n7199), .A2(n7188), .ZN(n7191) );
  OR2_X1 U8349 ( .A1(n10428), .A2(n7315), .ZN(n7185) );
  NAND2_X1 U8350 ( .A1(n7186), .A2(n5555), .ZN(n7210) );
  INV_X1 U8351 ( .A(n7205), .ZN(n7187) );
  NOR2_X1 U8352 ( .A1(n8011), .A2(n8218), .ZN(n7940) );
  INV_X1 U8353 ( .A(n7940), .ZN(n7190) );
  OAI21_X2 U8354 ( .B1(n7191), .B2(n7190), .A(n10326), .ZN(n10023) );
  OR2_X1 U8355 ( .A1(n7199), .A2(n7192), .ZN(n7194) );
  INV_X1 U8356 ( .A(n7194), .ZN(n7193) );
  NAND2_X1 U8357 ( .A1(n7193), .A2(n7321), .ZN(n10020) );
  NOR2_X2 U8358 ( .A1(n7194), .A2(n7321), .ZN(n10017) );
  AOI22_X1 U8359 ( .A1(n10029), .A2(n10017), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n7202) );
  INV_X1 U8360 ( .A(n10428), .ZN(n10835) );
  NAND2_X1 U8361 ( .A1(n7199), .A2(n10835), .ZN(n7196) );
  NAND2_X1 U8362 ( .A1(n7196), .A2(n7195), .ZN(n7748) );
  NAND2_X1 U8363 ( .A1(n7319), .A2(n6949), .ZN(n7197) );
  OAI21_X1 U8364 ( .B1(n7748), .B2(n7197), .A(P1_STATE_REG_SCAN_IN), .ZN(n7200) );
  AND2_X1 U8365 ( .A1(n7940), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7198) );
  NAND2_X1 U8366 ( .A1(n7199), .A2(n7198), .ZN(n7749) );
  NAND2_X1 U8367 ( .A1(n10158), .A2(n10015), .ZN(n7201) );
  OAI211_X1 U8368 ( .C1(n7203), .C2(n10020), .A(n7202), .B(n7201), .ZN(n7207)
         );
  NOR3_X1 U8369 ( .A1(n7205), .A2(n10026), .A3(n7204), .ZN(n7206) );
  AOI211_X1 U8370 ( .C1(n10157), .C2(n10023), .A(n7207), .B(n7206), .ZN(n7208)
         );
  NAND3_X1 U8371 ( .A1(n7210), .A2(n7209), .A3(n7208), .ZN(P1_U3220) );
  OAI21_X1 U8372 ( .B1(n7213), .B2(n5013), .A(n10002), .ZN(n7220) );
  OAI22_X1 U8373 ( .A1(n10208), .A2(n10020), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7214), .ZN(n7216) );
  NOR2_X1 U8374 ( .A1(n10172), .A2(n9991), .ZN(n7215) );
  AOI211_X1 U8375 ( .C1(n10179), .C2(n10015), .A(n7216), .B(n7215), .ZN(n7217)
         );
  INV_X1 U8376 ( .A(n7218), .ZN(n7219) );
  NAND2_X1 U8377 ( .A1(n7220), .A2(n7219), .ZN(P1_U3214) );
  NAND2_X1 U8378 ( .A1(n7221), .A2(n9351), .ZN(n7222) );
  NAND2_X1 U8379 ( .A1(n7222), .A2(n9312), .ZN(n7225) );
  NAND2_X1 U8380 ( .A1(n9841), .A2(n6275), .ZN(n7224) );
  NAND2_X1 U8381 ( .A1(n6258), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7223) );
  OR2_X2 U8382 ( .A1(n7243), .A2(n8988), .ZN(n9319) );
  NAND2_X1 U8383 ( .A1(n7243), .A2(n8988), .ZN(n9316) );
  NAND2_X1 U8384 ( .A1(n9319), .A2(n9316), .ZN(n9353) );
  INV_X1 U8385 ( .A(n7878), .ZN(n8545) );
  INV_X1 U8386 ( .A(n9499), .ZN(n9374) );
  NAND2_X1 U8387 ( .A1(n6267), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n7228) );
  NAND2_X1 U8388 ( .A1(n6595), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7227) );
  NAND2_X1 U8389 ( .A1(n6547), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n7226) );
  NAND4_X1 U8390 ( .A1(n9304), .A2(n7228), .A3(n7227), .A4(n7226), .ZN(n9373)
         );
  AND2_X1 U8391 ( .A1(n6252), .A2(P2_B_REG_SCAN_IN), .ZN(n7229) );
  NOR2_X1 U8392 ( .A1(n9685), .A2(n7229), .ZN(n9471) );
  AOI22_X1 U8393 ( .A1(n9540), .A2(n9374), .B1(n9373), .B2(n9471), .ZN(n7230)
         );
  NAND2_X1 U8394 ( .A1(n9489), .A2(n9499), .ZN(n7231) );
  NAND2_X1 U8395 ( .A1(n9282), .A2(n9374), .ZN(n7233) );
  NAND2_X1 U8396 ( .A1(n7234), .A2(n7233), .ZN(n7236) );
  XNOR2_X1 U8397 ( .A(n7236), .B(n7235), .ZN(n7238) );
  INV_X1 U8398 ( .A(n9682), .ZN(n7237) );
  NAND2_X1 U8399 ( .A1(n7238), .A2(n7237), .ZN(n7239) );
  AND2_X1 U8400 ( .A1(n7240), .A2(n7241), .ZN(n7242) );
  NOR2_X1 U8401 ( .A1(n9479), .A2(n7242), .ZN(n7249) );
  OR2_X1 U8402 ( .A1(n7249), .A2(n7244), .ZN(n7248) );
  INV_X1 U8403 ( .A(n7243), .ZN(n9480) );
  NAND2_X1 U8404 ( .A1(n7244), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7245) );
  INV_X1 U8405 ( .A(n7246), .ZN(n7247) );
  NAND2_X1 U8406 ( .A1(n7248), .A2(n7247), .ZN(P2_U3456) );
  OR2_X1 U8407 ( .A1(n7249), .A2(n7250), .ZN(n7254) );
  NAND2_X1 U8408 ( .A1(n7250), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n7251) );
  OAI21_X1 U8409 ( .B1(n9480), .B2(n9753), .A(n7251), .ZN(n7252) );
  INV_X1 U8410 ( .A(n7252), .ZN(n7253) );
  NAND2_X1 U8411 ( .A1(n7254), .A2(n7253), .ZN(P2_U3488) );
  NOR2_X1 U8412 ( .A1(n6949), .A2(P1_U3086), .ZN(n7255) );
  INV_X4 U8413 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U8414 ( .A(n7296), .ZN(n7256) );
  NAND2_X1 U8415 ( .A1(n9269), .A2(n7291), .ZN(n7257) );
  NAND2_X1 U8416 ( .A1(n7257), .A2(n7296), .ZN(n7592) );
  NAND2_X1 U8417 ( .A1(n7592), .A2(n6599), .ZN(n7258) );
  NAND2_X1 U8418 ( .A1(n7258), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NOR2_X1 U8419 ( .A1(n7259), .A2(n7262), .ZN(n7261) );
  NAND2_X1 U8420 ( .A1(n7261), .A2(n7260), .ZN(n7264) );
  NAND2_X1 U8421 ( .A1(n7262), .A2(n6221), .ZN(n7263) );
  XNOR2_X1 U8422 ( .A(n7915), .B(n8966), .ZN(n7276) );
  INV_X1 U8423 ( .A(n9391), .ZN(n7824) );
  OAI21_X1 U8424 ( .B1(n7648), .B2(n8966), .A(n7631), .ZN(n7613) );
  INV_X1 U8425 ( .A(n7267), .ZN(n7268) );
  NOR2_X1 U8426 ( .A1(n7611), .A2(n7268), .ZN(n7619) );
  XNOR2_X1 U8427 ( .A(n4960), .B(n7895), .ZN(n7271) );
  XNOR2_X1 U8428 ( .A(n7271), .B(n9392), .ZN(n7620) );
  NOR2_X1 U8429 ( .A1(n9392), .A2(n7271), .ZN(n7272) );
  XNOR2_X1 U8430 ( .A(n7273), .B(n9391), .ZN(n7710) );
  NAND2_X1 U8431 ( .A1(n7908), .A2(n7274), .ZN(n7275) );
  OAI21_X1 U8432 ( .B1(n7908), .B2(n7274), .A(n7275), .ZN(n7794) );
  NOR2_X1 U8433 ( .A1(n7795), .A2(n7794), .ZN(n7904) );
  INV_X1 U8434 ( .A(n7275), .ZN(n7903) );
  XNOR2_X1 U8435 ( .A(n8070), .B(n7276), .ZN(n7902) );
  OAI21_X2 U8436 ( .B1(n7904), .B2(n7903), .A(n7902), .ZN(n7901) );
  OAI21_X1 U8437 ( .B1(n7276), .B2(n9390), .A(n7901), .ZN(n8050) );
  XNOR2_X1 U8438 ( .A(n8098), .B(n7269), .ZN(n7277) );
  XNOR2_X1 U8439 ( .A(n7907), .B(n7277), .ZN(n8051) );
  INV_X1 U8440 ( .A(n7277), .ZN(n7278) );
  XNOR2_X1 U8441 ( .A(n8180), .B(n7269), .ZN(n7279) );
  XNOR2_X1 U8442 ( .A(n9388), .B(n7279), .ZN(n8176) );
  XNOR2_X1 U8443 ( .A(n8193), .B(n7270), .ZN(n8414) );
  XNOR2_X1 U8444 ( .A(n8414), .B(n9387), .ZN(n7280) );
  XNOR2_X1 U8445 ( .A(n8418), .B(n7280), .ZN(n7288) );
  NAND2_X1 U8446 ( .A1(n7289), .A2(n7281), .ZN(n7285) );
  INV_X1 U8447 ( .A(n7282), .ZN(n7283) );
  NAND2_X1 U8448 ( .A1(n7299), .A2(n7283), .ZN(n7284) );
  NAND2_X1 U8449 ( .A1(n7285), .A2(n7284), .ZN(n7294) );
  AND3_X1 U8450 ( .A1(n9269), .A2(n9773), .A3(n7354), .ZN(n7286) );
  NOR2_X1 U8451 ( .A1(n7288), .A2(n9127), .ZN(n7308) );
  INV_X1 U8452 ( .A(n7259), .ZN(n9546) );
  NAND2_X1 U8453 ( .A1(n7289), .A2(n9546), .ZN(n7290) );
  INV_X1 U8454 ( .A(n9079), .ZN(n9139) );
  NOR2_X1 U8455 ( .A1(n8193), .A2(n9139), .ZN(n7307) );
  NAND2_X1 U8456 ( .A1(n7292), .A2(n7291), .ZN(n7293) );
  OAI21_X1 U8457 ( .B1(n7294), .B2(n7293), .A(P2_STATE_REG_SCAN_IN), .ZN(n7298) );
  OR2_X1 U8458 ( .A1(n7295), .A2(n7361), .ZN(n7300) );
  INV_X1 U8459 ( .A(n7300), .ZN(n9367) );
  NOR2_X1 U8460 ( .A1(n7296), .A2(P2_U3151), .ZN(n9365) );
  AOI21_X1 U8461 ( .B1(n9367), .B2(n7299), .A(n9365), .ZN(n7297) );
  AND2_X1 U8462 ( .A1(n9136), .A2(n8198), .ZN(n7306) );
  NOR2_X1 U8463 ( .A1(n7300), .A2(n7299), .ZN(n7303) );
  NAND2_X1 U8464 ( .A1(n9388), .A2(n9132), .ZN(n7304) );
  OR2_X1 U8465 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8750), .ZN(n7994) );
  OAI211_X1 U8466 ( .C1(n8577), .C2(n9134), .A(n7304), .B(n7994), .ZN(n7305)
         );
  OR4_X1 U8467 ( .A1(n7308), .A2(n7307), .A3(n7306), .A4(n7305), .ZN(P2_U3161)
         );
  INV_X1 U8468 ( .A(n10124), .ZN(n10489) );
  AND2_X1 U8469 ( .A1(n7321), .A2(n10489), .ZN(n10553) );
  INV_X1 U8470 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10555) );
  NOR2_X1 U8471 ( .A1(n10485), .A2(n10555), .ZN(n7309) );
  XNOR2_X1 U8472 ( .A(n7309), .B(n10557), .ZN(n7314) );
  OAI21_X1 U8473 ( .B1(n7312), .B2(n7311), .A(n7310), .ZN(n7754) );
  NAND2_X1 U8474 ( .A1(n7754), .A2(n10553), .ZN(n7313) );
  OAI211_X1 U8475 ( .C1(n10553), .C2(n7314), .A(n7313), .B(n10852), .ZN(n7551)
         );
  NAND2_X1 U8476 ( .A1(n7315), .A2(n7319), .ZN(n7317) );
  NAND2_X1 U8477 ( .A1(n7317), .A2(n7316), .ZN(n7342) );
  INV_X1 U8478 ( .A(n6949), .ZN(n7318) );
  NAND2_X1 U8479 ( .A1(n7319), .A2(n7318), .ZN(n7320) );
  NAND2_X1 U8480 ( .A1(n7320), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7341) );
  AND2_X1 U8481 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7860) );
  AOI21_X1 U8482 ( .B1(n10076), .B2(n7433), .A(n7860), .ZN(n7340) );
  INV_X1 U8483 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7322) );
  MUX2_X1 U8484 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7322), .S(n7433), .Z(n7327)
         );
  XNOR2_X1 U8485 ( .A(n7367), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n7556) );
  XNOR2_X1 U8486 ( .A(n7349), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n10047) );
  AND2_X1 U8487 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n10046) );
  NAND2_X1 U8488 ( .A1(n10047), .A2(n10046), .ZN(n10045) );
  INV_X1 U8489 ( .A(n7349), .ZN(n10051) );
  NAND2_X1 U8490 ( .A1(n10051), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7323) );
  NAND2_X1 U8491 ( .A1(n10045), .A2(n7323), .ZN(n7555) );
  NAND2_X1 U8492 ( .A1(n7556), .A2(n7555), .ZN(n7554) );
  INV_X1 U8493 ( .A(n7367), .ZN(n7557) );
  NAND2_X1 U8494 ( .A1(n7557), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7324) );
  NAND2_X1 U8495 ( .A1(n7554), .A2(n7324), .ZN(n10059) );
  XNOR2_X1 U8496 ( .A(n10061), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n10060) );
  NAND2_X1 U8497 ( .A1(n10059), .A2(n10060), .ZN(n10058) );
  INV_X1 U8498 ( .A(n10061), .ZN(n7334) );
  NAND2_X1 U8499 ( .A1(n7334), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7325) );
  NAND2_X1 U8500 ( .A1(n10058), .A2(n7325), .ZN(n7326) );
  NAND2_X1 U8501 ( .A1(n7326), .A2(n7327), .ZN(n7435) );
  OAI211_X1 U8502 ( .C1(n7327), .C2(n7326), .A(n10072), .B(n7435), .ZN(n7339)
         );
  INV_X1 U8503 ( .A(n10090), .ZN(n10120) );
  INV_X1 U8504 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n7328) );
  MUX2_X1 U8505 ( .A(n7328), .B(P1_REG1_REG_2__SCAN_IN), .S(n7367), .Z(n7553)
         );
  INV_X1 U8506 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7329) );
  MUX2_X1 U8507 ( .A(n7329), .B(P1_REG1_REG_1__SCAN_IN), .S(n7349), .Z(n10049)
         );
  AND2_X1 U8508 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n10050) );
  NAND2_X1 U8509 ( .A1(n10049), .A2(n10050), .ZN(n10048) );
  NAND2_X1 U8510 ( .A1(n10051), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7330) );
  NAND2_X1 U8511 ( .A1(n10048), .A2(n7330), .ZN(n7552) );
  NAND2_X1 U8512 ( .A1(n7553), .A2(n7552), .ZN(n10063) );
  NAND2_X1 U8513 ( .A1(n7557), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n10062) );
  NAND2_X1 U8514 ( .A1(n10063), .A2(n10062), .ZN(n7333) );
  INV_X1 U8515 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7331) );
  MUX2_X1 U8516 ( .A(n7331), .B(P1_REG1_REG_3__SCAN_IN), .S(n10061), .Z(n7332)
         );
  NAND2_X1 U8517 ( .A1(n7333), .A2(n7332), .ZN(n10066) );
  NAND2_X1 U8518 ( .A1(n7334), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7336) );
  INV_X1 U8519 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10788) );
  MUX2_X1 U8520 ( .A(n10788), .B(P1_REG1_REG_4__SCAN_IN), .S(n7433), .Z(n7335)
         );
  AOI21_X1 U8521 ( .B1(n10066), .B2(n7336), .A(n7335), .ZN(n7445) );
  INV_X1 U8522 ( .A(n7445), .ZN(n10081) );
  NAND3_X1 U8523 ( .A1(n10066), .A2(n7336), .A3(n7335), .ZN(n7337) );
  NAND3_X1 U8524 ( .A1(n10120), .A2(n10081), .A3(n7337), .ZN(n7338) );
  NAND4_X1 U8525 ( .A1(n7551), .A2(n7340), .A3(n7339), .A4(n7338), .ZN(n7345)
         );
  INV_X1 U8526 ( .A(n7341), .ZN(n7343) );
  AND2_X1 U8527 ( .A1(n10560), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n7344) );
  OR2_X1 U8528 ( .A1(n7345), .A2(n7344), .ZN(P1_U3247) );
  AND2_X1 U8529 ( .A1(n7346), .A2(P2_U3151), .ZN(n9848) );
  INV_X2 U8530 ( .A(n9848), .ZN(n9856) );
  AOI22_X1 U8531 ( .A1(n7745), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n9846), .ZN(n7347) );
  OAI21_X1 U8532 ( .B1(n7365), .B2(n9856), .A(n7347), .ZN(P2_U3292) );
  AOI22_X1 U8533 ( .A1(n10599), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n9846), .ZN(n7348) );
  OAI21_X1 U8534 ( .B1(n7373), .B2(n9856), .A(n7348), .ZN(P2_U3291) );
  NOR2_X1 U8535 ( .A1(n4964), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10477) );
  INV_X2 U8536 ( .A(n10477), .ZN(n10494) );
  INV_X2 U8537 ( .A(n8886), .ZN(n10492) );
  OAI222_X1 U8538 ( .A1(n10494), .A2(n5458), .B1(n10492), .B2(n7352), .C1(
        n7349), .C2(P1_U3086), .ZN(P1_U3354) );
  INV_X1 U8539 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n7351) );
  INV_X1 U8540 ( .A(n7350), .ZN(n7368) );
  OAI222_X1 U8541 ( .A1(n9855), .A2(n7351), .B1(n9856), .B2(n7368), .C1(
        P2_U3151), .C2(n5441), .ZN(P2_U3293) );
  OAI222_X1 U8542 ( .A1(n10571), .A2(P2_U3151), .B1(n9855), .B2(n5581), .C1(
        n9856), .C2(n7352), .ZN(P2_U3294) );
  NAND2_X1 U8543 ( .A1(n7354), .A2(n7353), .ZN(n7380) );
  INV_X1 U8544 ( .A(n7355), .ZN(n7356) );
  AOI22_X1 U8545 ( .A1(n7380), .A2(n7358), .B1(n7357), .B2(n7356), .ZN(
        P2_U3376) );
  INV_X1 U8546 ( .A(n10610), .ZN(n7684) );
  INV_X1 U8547 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7359) );
  OAI222_X1 U8548 ( .A1(P2_U3151), .A2(n7684), .B1(n9856), .B2(n7371), .C1(
        n7359), .C2(n9855), .ZN(P2_U3290) );
  NAND2_X1 U8549 ( .A1(n7361), .A2(P2_D_REG_1__SCAN_IN), .ZN(n7360) );
  OAI21_X1 U8550 ( .B1(n7636), .B2(n7361), .A(n7360), .ZN(P2_U3377) );
  INV_X1 U8551 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7362) );
  OAI222_X1 U8552 ( .A1(P2_U3151), .A2(n7978), .B1(n9856), .B2(n7363), .C1(
        n7362), .C2(n9855), .ZN(P2_U3289) );
  INV_X1 U8553 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7364) );
  INV_X1 U8554 ( .A(n7461), .ZN(n7452) );
  OAI222_X1 U8555 ( .A1(n10494), .A2(n7364), .B1(n10492), .B2(n7363), .C1(
        n7452), .C2(P1_U3086), .ZN(P1_U3349) );
  OAI222_X1 U8556 ( .A1(n10494), .A2(n7366), .B1(n10492), .B2(n7365), .C1(
        n10061), .C2(P1_U3086), .ZN(P1_U3352) );
  OAI222_X1 U8557 ( .A1(n10494), .A2(n7369), .B1(n10492), .B2(n7368), .C1(
        n7367), .C2(P1_U3086), .ZN(P1_U3353) );
  INV_X1 U8558 ( .A(n10078), .ZN(n7370) );
  OAI222_X1 U8559 ( .A1(n10494), .A2(n7372), .B1(n10492), .B2(n7371), .C1(
        n7370), .C2(P1_U3086), .ZN(P1_U3350) );
  INV_X1 U8560 ( .A(n7433), .ZN(n7442) );
  OAI222_X1 U8561 ( .A1(P1_U3086), .A2(n7442), .B1(n10492), .B2(n7373), .C1(
        n10494), .C2(n5664), .ZN(P1_U3351) );
  INV_X1 U8562 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7374) );
  OAI222_X1 U8563 ( .A1(P2_U3151), .A2(n5059), .B1(n9856), .B2(n7375), .C1(
        n7374), .C2(n9855), .ZN(P2_U3288) );
  INV_X1 U8564 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7376) );
  INV_X1 U8565 ( .A(n7460), .ZN(n7481) );
  OAI222_X1 U8566 ( .A1(n10494), .A2(n7376), .B1(n10492), .B2(n7375), .C1(
        n7481), .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U8567 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7378) );
  INV_X1 U8568 ( .A(n7377), .ZN(n7379) );
  INV_X1 U8569 ( .A(n7492), .ZN(n7486) );
  OAI222_X1 U8570 ( .A1(n10494), .A2(n7378), .B1(n10492), .B2(n7379), .C1(
        P1_U3086), .C2(n7486), .ZN(P1_U3347) );
  INV_X1 U8571 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7599) );
  OAI222_X1 U8572 ( .A1(n8308), .A2(P2_U3151), .B1(n9856), .B2(n7379), .C1(
        n9855), .C2(n7599), .ZN(P2_U3287) );
  INV_X1 U8573 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n7381) );
  NOR2_X1 U8574 ( .A1(n7400), .A2(n7381), .ZN(P2_U3252) );
  INV_X1 U8575 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n7382) );
  NOR2_X1 U8576 ( .A1(n7400), .A2(n7382), .ZN(P2_U3244) );
  INV_X1 U8577 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n7383) );
  NOR2_X1 U8578 ( .A1(n7400), .A2(n7383), .ZN(P2_U3246) );
  INV_X1 U8579 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n7384) );
  NOR2_X1 U8580 ( .A1(n7400), .A2(n7384), .ZN(P2_U3247) );
  INV_X1 U8581 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n7385) );
  NOR2_X1 U8582 ( .A1(n7400), .A2(n7385), .ZN(P2_U3248) );
  INV_X1 U8583 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n7386) );
  NOR2_X1 U8584 ( .A1(n7400), .A2(n7386), .ZN(P2_U3249) );
  INV_X1 U8585 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n7387) );
  NOR2_X1 U8586 ( .A1(n7400), .A2(n7387), .ZN(P2_U3250) );
  INV_X1 U8587 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n7388) );
  NOR2_X1 U8588 ( .A1(n7400), .A2(n7388), .ZN(P2_U3251) );
  INV_X1 U8589 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n7389) );
  NOR2_X1 U8590 ( .A1(n7400), .A2(n7389), .ZN(P2_U3239) );
  INV_X1 U8591 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n7390) );
  NOR2_X1 U8592 ( .A1(n7400), .A2(n7390), .ZN(P2_U3254) );
  INV_X1 U8593 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n7391) );
  NOR2_X1 U8594 ( .A1(n7400), .A2(n7391), .ZN(P2_U3240) );
  INV_X1 U8595 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n7392) );
  NOR2_X1 U8596 ( .A1(n7400), .A2(n7392), .ZN(P2_U3241) );
  INV_X1 U8597 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n7393) );
  NOR2_X1 U8598 ( .A1(n7400), .A2(n7393), .ZN(P2_U3242) );
  INV_X1 U8599 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n7394) );
  NOR2_X1 U8600 ( .A1(n7400), .A2(n7394), .ZN(P2_U3253) );
  INV_X1 U8601 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7395) );
  INV_X1 U8602 ( .A(n7531), .ZN(n7508) );
  OAI222_X1 U8603 ( .A1(n10494), .A2(n7395), .B1(n10492), .B2(n7397), .C1(
        n7508), .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U8604 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7396) );
  OAI222_X1 U8605 ( .A1(P2_U3151), .A2(n9417), .B1(n9856), .B2(n7397), .C1(
        n7396), .C2(n9855), .ZN(P2_U3285) );
  INV_X1 U8606 ( .A(n7500), .ZN(n7507) );
  INV_X1 U8607 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7427) );
  INV_X1 U8608 ( .A(n7398), .ZN(n7399) );
  OAI222_X1 U8609 ( .A1(P1_U3086), .A2(n7507), .B1(n10494), .B2(n7427), .C1(
        n7399), .C2(n10492), .ZN(P1_U3346) );
  INV_X1 U8610 ( .A(n9413), .ZN(n9397) );
  INV_X1 U8611 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7602) );
  OAI222_X1 U8612 ( .A1(n9397), .A2(P2_U3151), .B1(n9855), .B2(n7602), .C1(
        n7399), .C2(n9856), .ZN(P2_U3286) );
  INV_X1 U8613 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n7401) );
  NOR2_X1 U8614 ( .A1(n7400), .A2(n7401), .ZN(P2_U3243) );
  INV_X1 U8615 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n7402) );
  NOR2_X1 U8616 ( .A1(n7400), .A2(n7402), .ZN(P2_U3257) );
  INV_X1 U8617 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n7403) );
  NOR2_X1 U8618 ( .A1(n7400), .A2(n7403), .ZN(P2_U3245) );
  INV_X1 U8619 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n7404) );
  NOR2_X1 U8620 ( .A1(n7400), .A2(n7404), .ZN(P2_U3259) );
  INV_X1 U8621 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n7405) );
  NOR2_X1 U8622 ( .A1(n7400), .A2(n7405), .ZN(P2_U3260) );
  INV_X1 U8623 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n7406) );
  NOR2_X1 U8624 ( .A1(n7400), .A2(n7406), .ZN(P2_U3256) );
  INV_X1 U8625 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n7407) );
  NOR2_X1 U8626 ( .A1(n7400), .A2(n7407), .ZN(P2_U3235) );
  INV_X1 U8627 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n7408) );
  NOR2_X1 U8628 ( .A1(n7400), .A2(n7408), .ZN(P2_U3236) );
  INV_X1 U8629 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n7409) );
  NOR2_X1 U8630 ( .A1(n7400), .A2(n7409), .ZN(P2_U3258) );
  INV_X1 U8631 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n7410) );
  NOR2_X1 U8632 ( .A1(n7400), .A2(n7410), .ZN(P2_U3238) );
  INV_X1 U8633 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n7411) );
  NOR2_X1 U8634 ( .A1(n7400), .A2(n7411), .ZN(P2_U3255) );
  INV_X1 U8635 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n7412) );
  NOR2_X1 U8636 ( .A1(n7400), .A2(n7412), .ZN(P2_U3261) );
  INV_X1 U8637 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n7413) );
  NOR2_X1 U8638 ( .A1(n7400), .A2(n7413), .ZN(P2_U3262) );
  INV_X1 U8639 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n7414) );
  NOR2_X1 U8640 ( .A1(n7400), .A2(n7414), .ZN(P2_U3263) );
  INV_X1 U8641 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n7415) );
  NOR2_X1 U8642 ( .A1(n7400), .A2(n7415), .ZN(P2_U3234) );
  INV_X1 U8643 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n7416) );
  NOR2_X1 U8644 ( .A1(n7400), .A2(n7416), .ZN(P2_U3237) );
  INV_X1 U8645 ( .A(n7417), .ZN(n7418) );
  INV_X1 U8646 ( .A(n10497), .ZN(n7422) );
  NAND2_X1 U8647 ( .A1(n7422), .A2(n7419), .ZN(n7420) );
  OAI21_X1 U8648 ( .B1(n7422), .B2(n7421), .A(n7420), .ZN(P1_U3440) );
  INV_X1 U8649 ( .A(n8887), .ZN(n7424) );
  INV_X1 U8650 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7423) );
  OAI222_X1 U8651 ( .A1(n5058), .A2(P2_U3151), .B1(n9856), .B2(n7424), .C1(
        n7423), .C2(n9855), .ZN(P2_U3284) );
  INV_X1 U8652 ( .A(n10766), .ZN(n9394) );
  INV_X1 U8653 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7930) );
  NAND2_X1 U8654 ( .A1(n8952), .A2(n9394), .ZN(n7425) );
  OAI21_X1 U8655 ( .B1(n9394), .B2(n7930), .A(n7425), .ZN(P2_U3509) );
  NAND2_X1 U8656 ( .A1(n8578), .A2(n9394), .ZN(n7426) );
  OAI21_X1 U8657 ( .B1(n9394), .B2(n7427), .A(n7426), .ZN(P2_U3500) );
  NAND2_X1 U8658 ( .A1(n7428), .A2(n9394), .ZN(n7429) );
  OAI21_X1 U8659 ( .B1(n9394), .B2(n5664), .A(n7429), .ZN(P2_U3495) );
  INV_X1 U8660 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7430) );
  INV_X1 U8661 ( .A(n7700), .ZN(n7546) );
  OAI222_X1 U8662 ( .A1(n10494), .A2(n7430), .B1(n10492), .B2(n7432), .C1(
        n7546), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U8663 ( .A(n10657), .ZN(n9441) );
  INV_X1 U8664 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7431) );
  OAI222_X1 U8665 ( .A1(P2_U3151), .A2(n9441), .B1(n9856), .B2(n7432), .C1(
        n7431), .C2(n9855), .ZN(P2_U3283) );
  NAND2_X1 U8666 ( .A1(n7433), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7434) );
  NAND2_X1 U8667 ( .A1(n7435), .A2(n7434), .ZN(n10073) );
  NAND2_X1 U8668 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n10078), .ZN(n7436) );
  OAI21_X1 U8669 ( .B1(n10078), .B2(P1_REG2_REG_5__SCAN_IN), .A(n7436), .ZN(
        n7437) );
  INV_X1 U8670 ( .A(n7437), .ZN(n10074) );
  AND2_X1 U8671 ( .A1(n10073), .A2(n10074), .ZN(n10070) );
  AOI21_X1 U8672 ( .B1(n10078), .B2(P1_REG2_REG_5__SCAN_IN), .A(n10070), .ZN(
        n7440) );
  NAND2_X1 U8673 ( .A1(n7461), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7438) );
  OAI21_X1 U8674 ( .B1(n7461), .B2(P1_REG2_REG_6__SCAN_IN), .A(n7438), .ZN(
        n7439) );
  NOR2_X1 U8675 ( .A1(n7440), .A2(n7439), .ZN(n7455) );
  AOI211_X1 U8676 ( .C1(n7440), .C2(n7439), .A(n7455), .B(n10122), .ZN(n7454)
         );
  INV_X1 U8677 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7441) );
  MUX2_X1 U8678 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n7441), .S(n7461), .Z(n7448)
         );
  NOR2_X1 U8679 ( .A1(n7442), .A2(n10788), .ZN(n10077) );
  INV_X1 U8680 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7443) );
  MUX2_X1 U8681 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n7443), .S(n10078), .Z(n7444)
         );
  OAI21_X1 U8682 ( .B1(n7445), .B2(n10077), .A(n7444), .ZN(n10083) );
  NAND2_X1 U8683 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n10078), .ZN(n7446) );
  NAND2_X1 U8684 ( .A1(n10083), .A2(n7446), .ZN(n7447) );
  NAND2_X1 U8685 ( .A1(n7448), .A2(n7447), .ZN(n7462) );
  OAI211_X1 U8686 ( .C1(n7448), .C2(n7447), .A(n10120), .B(n7462), .ZN(n7451)
         );
  NOR2_X1 U8687 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7449), .ZN(n7954) );
  AOI21_X1 U8688 ( .B1(n10560), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n7954), .ZN(
        n7450) );
  OAI211_X1 U8689 ( .C1(n10117), .C2(n7452), .A(n7451), .B(n7450), .ZN(n7453)
         );
  OR2_X1 U8690 ( .A1(n7454), .A2(n7453), .ZN(P1_U3249) );
  AOI21_X1 U8691 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n7461), .A(n7455), .ZN(
        n7475) );
  NAND2_X1 U8692 ( .A1(n7460), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7456) );
  OAI21_X1 U8693 ( .B1(n7460), .B2(P1_REG2_REG_7__SCAN_IN), .A(n7456), .ZN(
        n7474) );
  NOR2_X1 U8694 ( .A1(n7475), .A2(n7474), .ZN(n7473) );
  AOI21_X1 U8695 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n7460), .A(n7473), .ZN(
        n7459) );
  NAND2_X1 U8696 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n7492), .ZN(n7457) );
  OAI21_X1 U8697 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n7492), .A(n7457), .ZN(
        n7458) );
  NOR2_X1 U8698 ( .A1(n7459), .A2(n7458), .ZN(n7491) );
  AOI211_X1 U8699 ( .C1(n7459), .C2(n7458), .A(n7491), .B(n10122), .ZN(n7472)
         );
  INV_X1 U8700 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n8256) );
  MUX2_X1 U8701 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n8256), .S(n7460), .Z(n7477)
         );
  NAND2_X1 U8702 ( .A1(n7461), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7463) );
  NAND2_X1 U8703 ( .A1(n7463), .A2(n7462), .ZN(n7478) );
  NAND2_X1 U8704 ( .A1(n7477), .A2(n7478), .ZN(n7476) );
  OAI21_X1 U8705 ( .B1(n7481), .B2(n8256), .A(n7476), .ZN(n7466) );
  INV_X1 U8706 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7464) );
  MUX2_X1 U8707 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n7464), .S(n7492), .Z(n7465)
         );
  NAND2_X1 U8708 ( .A1(n7465), .A2(n7466), .ZN(n7485) );
  OAI211_X1 U8709 ( .C1(n7466), .C2(n7465), .A(n10120), .B(n7485), .ZN(n7470)
         );
  NOR2_X1 U8710 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7467), .ZN(n7468) );
  AOI21_X1 U8711 ( .B1(n10560), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n7468), .ZN(
        n7469) );
  OAI211_X1 U8712 ( .C1(n10117), .C2(n7486), .A(n7470), .B(n7469), .ZN(n7471)
         );
  OR2_X1 U8713 ( .A1(n7472), .A2(n7471), .ZN(P1_U3251) );
  AOI211_X1 U8714 ( .C1(n7475), .C2(n7474), .A(n7473), .B(n10122), .ZN(n7483)
         );
  OAI211_X1 U8715 ( .C1(n7478), .C2(n7477), .A(n10120), .B(n7476), .ZN(n7480)
         );
  AND2_X1 U8716 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8062) );
  AOI21_X1 U8717 ( .B1(n10560), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n8062), .ZN(
        n7479) );
  OAI211_X1 U8718 ( .C1(n10117), .C2(n7481), .A(n7480), .B(n7479), .ZN(n7482)
         );
  OR2_X1 U8719 ( .A1(n7483), .A2(n7482), .ZN(P1_U3250) );
  INV_X1 U8720 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7484) );
  MUX2_X1 U8721 ( .A(n7484), .B(P1_REG1_REG_9__SCAN_IN), .S(n7500), .Z(n7488)
         );
  OAI21_X1 U8722 ( .B1(n7486), .B2(n7464), .A(n7485), .ZN(n7487) );
  NOR2_X1 U8723 ( .A1(n7488), .A2(n7487), .ZN(n7506) );
  AOI21_X1 U8724 ( .B1(n7488), .B2(n7487), .A(n7506), .ZN(n7490) );
  AND2_X1 U8725 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n8382) );
  AOI21_X1 U8726 ( .B1(n10560), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n8382), .ZN(
        n7489) );
  OAI21_X1 U8727 ( .B1(n7490), .B2(n10090), .A(n7489), .ZN(n7497) );
  AOI21_X1 U8728 ( .B1(n7492), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7491), .ZN(
        n7495) );
  NOR2_X1 U8729 ( .A1(n7500), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7493) );
  AOI21_X1 U8730 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n7500), .A(n7493), .ZN(
        n7494) );
  NAND2_X1 U8731 ( .A1(n7494), .A2(n7495), .ZN(n7499) );
  AOI221_X1 U8732 ( .B1(n7495), .B2(n7499), .C1(n7494), .C2(n7499), .A(n10122), 
        .ZN(n7496) );
  AOI211_X1 U8733 ( .C1(n10076), .C2(n7500), .A(n7497), .B(n7496), .ZN(n7498)
         );
  INV_X1 U8734 ( .A(n7498), .ZN(P1_U3252) );
  OAI21_X1 U8735 ( .B1(n7500), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7499), .ZN(
        n7528) );
  INV_X1 U8736 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7501) );
  AOI22_X1 U8737 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n7508), .B1(n7531), .B2(
        n7501), .ZN(n7527) );
  NOR2_X1 U8738 ( .A1(n7528), .A2(n7527), .ZN(n7526) );
  AOI21_X1 U8739 ( .B1(n7531), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7526), .ZN(
        n7504) );
  INV_X1 U8740 ( .A(n8885), .ZN(n7537) );
  INV_X1 U8741 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7502) );
  AOI22_X1 U8742 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n7537), .B1(n8885), .B2(
        n7502), .ZN(n7503) );
  NOR2_X1 U8743 ( .A1(n7504), .A2(n7503), .ZN(n7541) );
  AOI211_X1 U8744 ( .C1(n7504), .C2(n7503), .A(n7541), .B(n10122), .ZN(n7514)
         );
  INV_X1 U8745 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7505) );
  MUX2_X1 U8746 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n7505), .S(n8885), .Z(n7510)
         );
  INV_X1 U8747 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10824) );
  MUX2_X1 U8748 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n10824), .S(n7531), .Z(n7520) );
  AOI21_X1 U8749 ( .B1(n7507), .B2(n7484), .A(n7506), .ZN(n7521) );
  NAND2_X1 U8750 ( .A1(n7520), .A2(n7521), .ZN(n7519) );
  OAI21_X1 U8751 ( .B1(n7508), .B2(n10824), .A(n7519), .ZN(n7509) );
  NAND2_X1 U8752 ( .A1(n7510), .A2(n7509), .ZN(n7536) );
  OAI211_X1 U8753 ( .C1(n7510), .C2(n7509), .A(n10120), .B(n7536), .ZN(n7512)
         );
  AND2_X1 U8754 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8566) );
  AOI21_X1 U8755 ( .B1(n10560), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n8566), .ZN(
        n7511) );
  OAI211_X1 U8756 ( .C1(n10117), .C2(n7537), .A(n7512), .B(n7511), .ZN(n7513)
         );
  OR2_X1 U8757 ( .A1(n7514), .A2(n7513), .ZN(P1_U3254) );
  INV_X1 U8758 ( .A(n10673), .ZN(n9439) );
  INV_X1 U8759 ( .A(n7515), .ZN(n7518) );
  INV_X1 U8760 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7516) );
  OAI222_X1 U8761 ( .A1(n9439), .A2(P2_U3151), .B1(n9856), .B2(n7518), .C1(
        n7516), .C2(n9855), .ZN(P2_U3282) );
  INV_X1 U8762 ( .A(n7801), .ZN(n7806) );
  INV_X1 U8763 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7517) );
  OAI222_X1 U8764 ( .A1(P1_U3086), .A2(n7806), .B1(n10492), .B2(n7518), .C1(
        n10494), .C2(n7517), .ZN(P1_U3342) );
  INV_X1 U8765 ( .A(n10560), .ZN(n7525) );
  INV_X1 U8766 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7524) );
  OAI211_X1 U8767 ( .C1(n7521), .C2(n7520), .A(n10120), .B(n7519), .ZN(n7523)
         );
  OR2_X1 U8768 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7522), .ZN(n8492) );
  OAI211_X1 U8769 ( .C1(n7525), .C2(n7524), .A(n7523), .B(n8492), .ZN(n7530)
         );
  AOI211_X1 U8770 ( .C1(n7528), .C2(n7527), .A(n7526), .B(n10122), .ZN(n7529)
         );
  AOI211_X1 U8771 ( .C1(n10076), .C2(n7531), .A(n7530), .B(n7529), .ZN(n7532)
         );
  INV_X1 U8772 ( .A(n7532), .ZN(P1_U3253) );
  INV_X1 U8773 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7534) );
  INV_X1 U8774 ( .A(n7533), .ZN(n7535) );
  INV_X1 U8775 ( .A(n8146), .ZN(n8151) );
  OAI222_X1 U8776 ( .A1(n10494), .A2(n7534), .B1(n10492), .B2(n7535), .C1(
        P1_U3086), .C2(n8151), .ZN(P1_U3341) );
  INV_X1 U8777 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7607) );
  OAI222_X1 U8778 ( .A1(n9437), .A2(P2_U3151), .B1(n9856), .B2(n7535), .C1(
        n9855), .C2(n7607), .ZN(P2_U3281) );
  NOR2_X1 U8779 ( .A1(n10560), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8780 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10841) );
  AOI22_X1 U8781 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n7546), .B1(n7700), .B2(
        n10841), .ZN(n7539) );
  OAI21_X1 U8782 ( .B1(n7537), .B2(n7505), .A(n7536), .ZN(n7538) );
  NOR2_X1 U8783 ( .A1(n7539), .A2(n7538), .ZN(n7702) );
  AOI21_X1 U8784 ( .B1(n7539), .B2(n7538), .A(n7702), .ZN(n7550) );
  NOR2_X1 U8785 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7700), .ZN(n7540) );
  AOI21_X1 U8786 ( .B1(n7700), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7540), .ZN(
        n7543) );
  AOI21_X1 U8787 ( .B1(n8885), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7541), .ZN(
        n7542) );
  NAND2_X1 U8788 ( .A1(n7543), .A2(n7542), .ZN(n7697) );
  OAI21_X1 U8789 ( .B1(n7543), .B2(n7542), .A(n7697), .ZN(n7544) );
  NAND2_X1 U8790 ( .A1(n7544), .A2(n10072), .ZN(n7549) );
  NOR2_X1 U8791 ( .A1(n7545), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9900) );
  NOR2_X1 U8792 ( .A1(n10117), .A2(n7546), .ZN(n7547) );
  AOI211_X1 U8793 ( .C1(n10560), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n9900), .B(
        n7547), .ZN(n7548) );
  OAI211_X1 U8794 ( .C1(n7550), .C2(n10090), .A(n7549), .B(n7548), .ZN(
        P1_U3255) );
  INV_X1 U8795 ( .A(n7551), .ZN(n7563) );
  OAI211_X1 U8796 ( .C1(n7553), .C2(n7552), .A(n10120), .B(n10063), .ZN(n7561)
         );
  OAI211_X1 U8797 ( .C1(n7556), .C2(n7555), .A(n10072), .B(n7554), .ZN(n7560)
         );
  AOI22_X1 U8798 ( .A1(n10560), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n7559) );
  NAND2_X1 U8799 ( .A1(n10076), .A2(n7557), .ZN(n7558) );
  NAND4_X1 U8800 ( .A1(n7561), .A2(n7560), .A3(n7559), .A4(n7558), .ZN(n7562)
         );
  OR2_X1 U8801 ( .A1(n7563), .A2(n7562), .ZN(P1_U3245) );
  MUX2_X1 U8802 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n6601), .Z(n7565) );
  XOR2_X1 U8803 ( .A(n10571), .B(n7565), .Z(n10584) );
  INV_X1 U8804 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7570) );
  INV_X1 U8805 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7564) );
  MUX2_X1 U8806 ( .A(n7570), .B(n7564), .S(n6601), .Z(n10565) );
  NAND2_X1 U8807 ( .A1(n10565), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n10583) );
  AOI22_X1 U8808 ( .A1(n10584), .A2(n10583), .B1(n7565), .B2(n10571), .ZN(
        n7671) );
  MUX2_X1 U8809 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n6601), .Z(n7668) );
  XOR2_X1 U8810 ( .A(n7680), .B(n7668), .Z(n7670) );
  XNOR2_X1 U8811 ( .A(n7671), .B(n7670), .ZN(n7596) );
  INV_X1 U8812 ( .A(n10772), .ZN(n8314) );
  INV_X1 U8813 ( .A(n7566), .ZN(n7567) );
  INV_X1 U8814 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7568) );
  NOR2_X1 U8815 ( .A1(n10605), .A2(n7568), .ZN(n7591) );
  NOR2_X1 U8816 ( .A1(n6600), .A2(P2_U3151), .ZN(n9845) );
  NAND2_X1 U8817 ( .A1(n7592), .A2(n9845), .ZN(n10564) );
  NAND2_X1 U8818 ( .A1(n7680), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7569) );
  NOR2_X1 U8819 ( .A1(n7570), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7571) );
  NAND2_X1 U8820 ( .A1(n6242), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7573) );
  INV_X1 U8821 ( .A(n10574), .ZN(n7572) );
  INV_X1 U8822 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10575) );
  NOR2_X1 U8823 ( .A1(n7574), .A2(n7575), .ZN(n7576) );
  NOR2_X1 U8824 ( .A1(n7576), .A2(n7653), .ZN(n7589) );
  OR2_X1 U8825 ( .A1(n10564), .A2(n7577), .ZN(n10755) );
  INV_X1 U8826 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7578) );
  MUX2_X1 U8827 ( .A(n7578), .B(P2_REG1_REG_2__SCAN_IN), .S(n7680), .Z(n7584)
         );
  INV_X1 U8828 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7579) );
  AND2_X1 U8829 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n7579), .ZN(n7580) );
  NAND2_X1 U8830 ( .A1(n6242), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7582) );
  OAI21_X1 U8831 ( .B1(n10571), .B2(n7580), .A(n7582), .ZN(n10576) );
  INV_X1 U8832 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7581) );
  OAI21_X1 U8833 ( .B1(n7584), .B2(n7583), .A(n7679), .ZN(n7585) );
  INV_X1 U8834 ( .A(n7585), .ZN(n7586) );
  OR2_X1 U8835 ( .A1(n10755), .A2(n7586), .ZN(n7588) );
  NAND2_X1 U8836 ( .A1(P2_U3151), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7587) );
  OAI211_X1 U8837 ( .C1(n10747), .C2(n7589), .A(n7588), .B(n7587), .ZN(n7590)
         );
  NOR2_X1 U8838 ( .A1(n7591), .A2(n7590), .ZN(n7595) );
  NOR2_X1 U8839 ( .A1(n6601), .A2(P2_U3151), .ZN(n9849) );
  AND2_X1 U8840 ( .A1(n7592), .A2(n9849), .ZN(n7593) );
  NAND2_X1 U8841 ( .A1(n10737), .A2(n7680), .ZN(n7594) );
  OAI211_X1 U8842 ( .C1(n7596), .C2(n8314), .A(n7595), .B(n7594), .ZN(P2_U3184) );
  INV_X1 U8843 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8915) );
  NAND2_X1 U8844 ( .A1(n10388), .A2(P1_U3973), .ZN(n7597) );
  OAI21_X1 U8845 ( .B1(n8915), .B2(P1_U3973), .A(n7597), .ZN(P1_U3574) );
  NAND2_X1 U8846 ( .A1(n8283), .A2(P1_U3973), .ZN(n7598) );
  OAI21_X1 U8847 ( .B1(P1_U3973), .B2(n7599), .A(n7598), .ZN(P1_U3562) );
  NAND2_X1 U8848 ( .A1(n7600), .A2(P1_U3973), .ZN(n7601) );
  OAI21_X1 U8849 ( .B1(n7602), .B2(P1_U3973), .A(n7601), .ZN(P1_U3563) );
  INV_X1 U8850 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7815) );
  NAND2_X1 U8851 ( .A1(n9993), .A2(P1_U3973), .ZN(n7603) );
  OAI21_X1 U8852 ( .B1(n7815), .B2(P1_U3973), .A(n7603), .ZN(P1_U3571) );
  INV_X1 U8853 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7975) );
  NAND2_X1 U8854 ( .A1(n7604), .A2(P1_U3973), .ZN(n7605) );
  OAI21_X1 U8855 ( .B1(n7975), .B2(P1_U3973), .A(n7605), .ZN(P1_U3573) );
  NAND2_X1 U8856 ( .A1(n8511), .A2(P1_U3973), .ZN(n7606) );
  OAI21_X1 U8857 ( .B1(n7607), .B2(P1_U3973), .A(n7606), .ZN(P1_U3568) );
  INV_X1 U8858 ( .A(n10705), .ZN(n9435) );
  INV_X1 U8859 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7608) );
  OAI222_X1 U8860 ( .A1(P2_U3151), .A2(n9435), .B1(n9856), .B2(n7609), .C1(
        n7608), .C2(n9855), .ZN(P2_U3280) );
  INV_X1 U8861 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7610) );
  OAI222_X1 U8862 ( .A1(n10494), .A2(n7610), .B1(n10492), .B2(n7609), .C1(
        n8447), .C2(P1_U3086), .ZN(P1_U3340) );
  AOI21_X1 U8863 ( .B1(n7613), .B2(n7612), .A(n7611), .ZN(n7617) );
  INV_X1 U8864 ( .A(n9136), .ZN(n8057) );
  NAND2_X1 U8865 ( .A1(n8057), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7770) );
  AOI22_X1 U8866 ( .A1(n6552), .A2(n9132), .B1(n7265), .B2(n9079), .ZN(n7614)
         );
  OAI21_X1 U8867 ( .B1(n6284), .B2(n9134), .A(n7614), .ZN(n7615) );
  AOI21_X1 U8868 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7770), .A(n7615), .ZN(
        n7616) );
  OAI21_X1 U8869 ( .B1(n7617), .B2(n9127), .A(n7616), .ZN(P2_U3162) );
  AOI21_X1 U8870 ( .B1(n7620), .B2(n7619), .A(n7618), .ZN(n7624) );
  AOI22_X1 U8871 ( .A1(n9393), .A2(n9132), .B1(n9079), .B2(n6283), .ZN(n7621)
         );
  OAI21_X1 U8872 ( .B1(n7824), .B2(n9134), .A(n7621), .ZN(n7622) );
  AOI21_X1 U8873 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n7770), .A(n7622), .ZN(
        n7623) );
  OAI21_X1 U8874 ( .B1(n7624), .B2(n9127), .A(n7623), .ZN(P2_U3177) );
  INV_X1 U8875 ( .A(n9778), .ZN(n9766) );
  INV_X1 U8876 ( .A(n7648), .ZN(n7775) );
  NAND2_X1 U8877 ( .A1(n6552), .A2(n7775), .ZN(n9147) );
  AND2_X1 U8878 ( .A1(n9147), .A2(n9144), .ZN(n9331) );
  AOI21_X1 U8879 ( .B1(n9682), .B2(n9766), .A(n9331), .ZN(n7626) );
  NOR2_X1 U8880 ( .A1(n7625), .A2(n9685), .ZN(n7646) );
  NOR2_X1 U8881 ( .A1(n7626), .A2(n7646), .ZN(n7778) );
  INV_X1 U8882 ( .A(n9753), .ZN(n8407) );
  AOI22_X1 U8883 ( .A1(n8407), .A2(n7648), .B1(n7250), .B2(
        P2_REG1_REG_0__SCAN_IN), .ZN(n7627) );
  OAI21_X1 U8884 ( .B1(n7778), .B2(n7250), .A(n7627), .ZN(P2_U3459) );
  OAI21_X1 U8885 ( .B1(n5190), .B2(n5189), .A(n7629), .ZN(n7924) );
  NOR2_X1 U8886 ( .A1(n7630), .A2(n9773), .ZN(n7634) );
  XNOR2_X1 U8887 ( .A(n7631), .B(n5190), .ZN(n7632) );
  OAI222_X1 U8888 ( .A1(n9684), .A2(n7633), .B1(n9685), .B2(n6284), .C1(n9682), 
        .C2(n7632), .ZN(n7921) );
  AOI211_X1 U8889 ( .C1(n9778), .C2(n7924), .A(n7634), .B(n7921), .ZN(n10778)
         );
  OR2_X1 U8890 ( .A1(n10778), .A2(n7250), .ZN(n7635) );
  OAI21_X1 U8891 ( .B1(n9781), .B2(n7581), .A(n7635), .ZN(P2_U3460) );
  OAI22_X1 U8892 ( .A1(n7639), .A2(n7638), .B1(n7637), .B2(n7636), .ZN(n7641)
         );
  INV_X1 U8893 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10570) );
  NOR2_X1 U8894 ( .A1(n9669), .A2(n10570), .ZN(n7645) );
  NOR3_X1 U8895 ( .A1(n9331), .A2(n7643), .A3(n7647), .ZN(n7644) );
  AOI211_X1 U8896 ( .C1(n7646), .C2(n9672), .A(n7645), .B(n7644), .ZN(n7650)
         );
  INV_X1 U8897 ( .A(n9652), .ZN(n8536) );
  NAND2_X1 U8898 ( .A1(n8536), .A2(n7648), .ZN(n7649) );
  OAI211_X1 U8899 ( .C1(n7570), .C2(n9672), .A(n7650), .B(n7649), .ZN(P2_U3233) );
  INV_X1 U8900 ( .A(n10599), .ZN(n7658) );
  INV_X1 U8901 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7651) );
  MUX2_X1 U8902 ( .A(n7651), .B(P2_REG2_REG_4__SCAN_IN), .S(n10599), .Z(n7652)
         );
  INV_X1 U8903 ( .A(n7657), .ZN(n7656) );
  NAND2_X1 U8904 ( .A1(n7654), .A2(n7745), .ZN(n7655) );
  NAND2_X1 U8905 ( .A1(n7656), .A2(n7655), .ZN(n7737) );
  INV_X1 U8906 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7736) );
  NOR2_X1 U8907 ( .A1(n7737), .A2(n7736), .ZN(n7735) );
  NOR2_X1 U8908 ( .A1(n10610), .A2(n7659), .ZN(n7660) );
  INV_X1 U8909 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10612) );
  NOR2_X1 U8910 ( .A1(n10613), .A2(n10612), .ZN(n10611) );
  INV_X1 U8911 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7661) );
  AOI22_X1 U8912 ( .A1(n8001), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n7661), .B2(
        n7978), .ZN(n7662) );
  AOI21_X1 U8913 ( .B1(n7663), .B2(n7662), .A(n7977), .ZN(n7695) );
  MUX2_X1 U8914 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n6601), .Z(n7664) );
  INV_X1 U8915 ( .A(n7664), .ZN(n7666) );
  NOR2_X1 U8916 ( .A1(n7664), .A2(n7978), .ZN(n7988) );
  INV_X1 U8917 ( .A(n7988), .ZN(n7665) );
  OAI21_X1 U8918 ( .B1(n8001), .B2(n7666), .A(n7665), .ZN(n7678) );
  MUX2_X1 U8919 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n6601), .Z(n7675) );
  NAND2_X1 U8920 ( .A1(n7675), .A2(n7684), .ZN(n7676) );
  MUX2_X1 U8921 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n6601), .Z(n7673) );
  INV_X1 U8922 ( .A(n7673), .ZN(n7674) );
  MUX2_X1 U8923 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n6601), .Z(n7667) );
  INV_X1 U8924 ( .A(n7667), .ZN(n7672) );
  XOR2_X1 U8925 ( .A(n7745), .B(n7667), .Z(n7731) );
  INV_X1 U8926 ( .A(n7668), .ZN(n7669) );
  OAI22_X1 U8927 ( .A1(n7671), .A2(n7670), .B1(n7680), .B2(n7669), .ZN(n7732)
         );
  NOR2_X1 U8928 ( .A1(n7731), .A2(n7732), .ZN(n7730) );
  AOI21_X1 U8929 ( .B1(n7672), .B2(n7745), .A(n7730), .ZN(n10602) );
  XNOR2_X1 U8930 ( .A(n7673), .B(n10599), .ZN(n10601) );
  NAND2_X1 U8931 ( .A1(n10602), .A2(n10601), .ZN(n10600) );
  OAI21_X1 U8932 ( .B1(n10599), .B2(n7674), .A(n10600), .ZN(n10619) );
  XNOR2_X1 U8933 ( .A(n7675), .B(n10610), .ZN(n10618) );
  NAND2_X1 U8934 ( .A1(n10619), .A2(n10618), .ZN(n10617) );
  NAND2_X1 U8935 ( .A1(n7676), .A2(n10617), .ZN(n7677) );
  NOR2_X1 U8936 ( .A1(n7678), .A2(n7677), .ZN(n7987) );
  AOI21_X1 U8937 ( .B1(n7678), .B2(n7677), .A(n7987), .ZN(n7692) );
  INV_X1 U8938 ( .A(n10605), .ZN(n10757) );
  INV_X1 U8939 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7683) );
  MUX2_X1 U8940 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n7683), .S(n10599), .Z(n10592) );
  NAND2_X1 U8941 ( .A1(n5437), .A2(n7681), .ZN(n7682) );
  XNOR2_X1 U8942 ( .A(n7681), .B(n7745), .ZN(n7734) );
  NAND2_X1 U8943 ( .A1(P2_REG1_REG_3__SCAN_IN), .A2(n7734), .ZN(n7733) );
  NAND2_X1 U8944 ( .A1(n7684), .A2(n7685), .ZN(n7686) );
  NAND2_X1 U8945 ( .A1(P2_REG1_REG_5__SCAN_IN), .A2(n10608), .ZN(n10607) );
  INV_X1 U8946 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n8000) );
  AOI22_X1 U8947 ( .A1(n8001), .A2(n8000), .B1(P2_REG1_REG_6__SCAN_IN), .B2(
        n7978), .ZN(n7687) );
  OAI21_X1 U8948 ( .B1(n7688), .B2(n7687), .A(n7999), .ZN(n7689) );
  AOI22_X1 U8949 ( .A1(n10757), .A2(P2_ADDR_REG_6__SCAN_IN), .B1(n7689), .B2(
        n10745), .ZN(n7691) );
  INV_X1 U8950 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8871) );
  NOR2_X1 U8951 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8871), .ZN(n8054) );
  INV_X1 U8952 ( .A(n8054), .ZN(n7690) );
  OAI211_X1 U8953 ( .C1(n7692), .C2(n8314), .A(n7691), .B(n7690), .ZN(n7693)
         );
  AOI21_X1 U8954 ( .B1(n8001), .B2(n10737), .A(n7693), .ZN(n7694) );
  OAI21_X1 U8955 ( .B1(n7695), .B2(n10747), .A(n7694), .ZN(P2_U3188) );
  INV_X1 U8956 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7696) );
  AOI22_X1 U8957 ( .A1(n7801), .A2(n7696), .B1(P1_REG2_REG_13__SCAN_IN), .B2(
        n7806), .ZN(n7699) );
  OAI21_X1 U8958 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7700), .A(n7697), .ZN(
        n7698) );
  NOR2_X1 U8959 ( .A1(n7699), .A2(n7698), .ZN(n7800) );
  AOI211_X1 U8960 ( .C1(n7699), .C2(n7698), .A(n7800), .B(n10122), .ZN(n7708)
         );
  NOR2_X1 U8961 ( .A1(n7700), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7701) );
  NOR2_X1 U8962 ( .A1(n7702), .A2(n7701), .ZN(n7704) );
  INV_X1 U8963 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n8606) );
  XNOR2_X1 U8964 ( .A(n7801), .B(n8606), .ZN(n7703) );
  NAND2_X1 U8965 ( .A1(n7704), .A2(n7703), .ZN(n7805) );
  OAI211_X1 U8966 ( .C1(n7704), .C2(n7703), .A(n7805), .B(n10120), .ZN(n7706)
         );
  AND2_X1 U8967 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9969) );
  AOI21_X1 U8968 ( .B1(n10560), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n9969), .ZN(
        n7705) );
  OAI211_X1 U8969 ( .C1(n10117), .C2(n7806), .A(n7706), .B(n7705), .ZN(n7707)
         );
  OR2_X1 U8970 ( .A1(n7708), .A2(n7707), .ZN(P1_U3256) );
  OAI211_X1 U8971 ( .C1(n7711), .C2(n7710), .A(n7709), .B(n9109), .ZN(n7715)
         );
  NOR2_X1 U8972 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8833), .ZN(n7740) );
  OAI22_X1 U8973 ( .A1(n6284), .A2(n9113), .B1(n7908), .B2(n9134), .ZN(n7712)
         );
  AOI211_X1 U8974 ( .C1(n9079), .C2(n7713), .A(n7740), .B(n7712), .ZN(n7714)
         );
  OAI211_X1 U8975 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8057), .A(n7715), .B(
        n7714), .ZN(P2_U3158) );
  INV_X1 U8976 ( .A(n7717), .ZN(n7719) );
  INV_X1 U8977 ( .A(n7716), .ZN(n9333) );
  NAND2_X1 U8978 ( .A1(n7717), .A2(n9333), .ZN(n7784) );
  INV_X1 U8979 ( .A(n7784), .ZN(n7718) );
  AOI21_X1 U8980 ( .B1(n7719), .B2(n7716), .A(n7718), .ZN(n7900) );
  INV_X1 U8981 ( .A(n7900), .ZN(n7724) );
  XNOR2_X1 U8982 ( .A(n7716), .B(n7720), .ZN(n7721) );
  NAND2_X1 U8983 ( .A1(n7721), .A2(n7237), .ZN(n7723) );
  INV_X1 U8984 ( .A(n9685), .ZN(n9541) );
  AOI22_X1 U8985 ( .A1(n9393), .A2(n9540), .B1(n9541), .B2(n9391), .ZN(n7722)
         );
  NAND2_X1 U8986 ( .A1(n7723), .A2(n7722), .ZN(n7896) );
  AOI21_X1 U8987 ( .B1(n7724), .B2(n9778), .A(n7896), .ZN(n7782) );
  AOI22_X1 U8988 ( .A1(n8407), .A2(n6283), .B1(n7250), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n7725) );
  OAI21_X1 U8989 ( .B1(n7782), .B2(n7250), .A(n7725), .ZN(P2_U3461) );
  INV_X1 U8990 ( .A(n7726), .ZN(n7728) );
  INV_X1 U8991 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7727) );
  OAI222_X1 U8992 ( .A1(n9433), .A2(P2_U3151), .B1(n9856), .B2(n7728), .C1(
        n7727), .C2(n9855), .ZN(P2_U3279) );
  INV_X1 U8993 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7729) );
  INV_X1 U8994 ( .A(n8555), .ZN(n8549) );
  OAI222_X1 U8995 ( .A1(n10494), .A2(n7729), .B1(n10492), .B2(n7728), .C1(
        P1_U3086), .C2(n8549), .ZN(P1_U3339) );
  AOI21_X1 U8996 ( .B1(n7732), .B2(n7731), .A(n7730), .ZN(n7747) );
  INV_X1 U8997 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n7743) );
  OAI21_X1 U8998 ( .B1(n7734), .B2(P2_REG1_REG_3__SCAN_IN), .A(n7733), .ZN(
        n7741) );
  AOI21_X1 U8999 ( .B1(n7737), .B2(n7736), .A(n7735), .ZN(n7738) );
  NOR2_X1 U9000 ( .A1(n10747), .A2(n7738), .ZN(n7739) );
  AOI211_X1 U9001 ( .C1(n10745), .C2(n7741), .A(n7740), .B(n7739), .ZN(n7742)
         );
  OAI21_X1 U9002 ( .B1(n10605), .B2(n7743), .A(n7742), .ZN(n7744) );
  AOI21_X1 U9003 ( .B1(n7745), .B2(n10737), .A(n7744), .ZN(n7746) );
  OAI21_X1 U9004 ( .B1(n7747), .B2(n8314), .A(n7746), .ZN(P2_U3185) );
  INV_X1 U9005 ( .A(n7748), .ZN(n7751) );
  NAND3_X1 U9006 ( .A1(n7751), .A2(n7750), .A3(n7749), .ZN(n7763) );
  AOI22_X1 U9007 ( .A1(n7763), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n10023), .B2(
        n8010), .ZN(n7753) );
  NAND2_X1 U9008 ( .A1(n10017), .A2(n10044), .ZN(n7752) );
  OAI211_X1 U9009 ( .C1(n10026), .C2(n7754), .A(n7753), .B(n7752), .ZN(
        P1_U3232) );
  XOR2_X1 U9010 ( .A(n7756), .B(n7755), .Z(n7759) );
  AOI22_X1 U9011 ( .A1(n10003), .A2(n10044), .B1(n10017), .B2(n10042), .ZN(
        n7758) );
  AOI22_X1 U9012 ( .A1(n7763), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n10023), .B2(
        n6945), .ZN(n7757) );
  OAI211_X1 U9013 ( .C1(n7759), .C2(n10026), .A(n7758), .B(n7757), .ZN(
        P1_U3237) );
  XNOR2_X1 U9014 ( .A(n7762), .B(n7761), .ZN(n7766) );
  AOI22_X1 U9015 ( .A1(n10003), .A2(n6960), .B1(n10017), .B2(n10043), .ZN(
        n7765) );
  AOI22_X1 U9016 ( .A1(n7763), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n10023), .B2(
        n6967), .ZN(n7764) );
  OAI211_X1 U9017 ( .C1(n7766), .C2(n10026), .A(n7765), .B(n7764), .ZN(
        P1_U3222) );
  INV_X1 U9018 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9852) );
  NAND2_X1 U9019 ( .A1(n10188), .A2(P1_U3973), .ZN(n7767) );
  OAI21_X1 U9020 ( .B1(n9852), .B2(P1_U3973), .A(n7767), .ZN(P1_U3581) );
  INV_X1 U9021 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9854) );
  NAND2_X1 U9022 ( .A1(n7768), .A2(P1_U3973), .ZN(n7769) );
  OAI21_X1 U9023 ( .B1(n9854), .B2(P1_U3973), .A(n7769), .ZN(P1_U3580) );
  NAND2_X1 U9024 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(n7770), .ZN(n7771) );
  OAI21_X1 U9025 ( .B1(n9139), .B2(n7775), .A(n7771), .ZN(n7772) );
  AOI21_X1 U9026 ( .B1(n9111), .B2(n9393), .A(n7772), .ZN(n7773) );
  OAI21_X1 U9027 ( .B1(n9331), .B2(n9127), .A(n7773), .ZN(P2_U3172) );
  INV_X1 U9028 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7774) );
  OAI22_X1 U9029 ( .A1(n9833), .A2(n7775), .B1(n10851), .B2(n7774), .ZN(n7776)
         );
  INV_X1 U9030 ( .A(n7776), .ZN(n7777) );
  OAI21_X1 U9031 ( .B1(n7778), .B2(n7244), .A(n7777), .ZN(P2_U3390) );
  INV_X1 U9032 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n7779) );
  OAI22_X1 U9033 ( .A1(n9833), .A2(n7895), .B1(n10851), .B2(n7779), .ZN(n7780)
         );
  INV_X1 U9034 ( .A(n7780), .ZN(n7781) );
  OAI21_X1 U9035 ( .B1(n7782), .B2(n7244), .A(n7781), .ZN(P2_U3396) );
  INV_X1 U9036 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7791) );
  NAND2_X1 U9037 ( .A1(n7784), .A2(n7783), .ZN(n7786) );
  INV_X1 U9038 ( .A(n9159), .ZN(n7785) );
  NOR2_X1 U9039 ( .A1(n9155), .A2(n7785), .ZN(n9330) );
  NAND2_X1 U9040 ( .A1(n7786), .A2(n9330), .ZN(n7818) );
  OAI21_X1 U9041 ( .B1(n7786), .B2(n9330), .A(n7818), .ZN(n7884) );
  NOR2_X1 U9042 ( .A1(n7880), .A2(n9773), .ZN(n7789) );
  XNOR2_X1 U9043 ( .A(n7787), .B(n9330), .ZN(n7788) );
  OAI222_X1 U9044 ( .A1(n9685), .A2(n7908), .B1(n9684), .B2(n6284), .C1(n9682), 
        .C2(n7788), .ZN(n7881) );
  AOI211_X1 U9045 ( .C1(n9778), .C2(n7884), .A(n7789), .B(n7881), .ZN(n10780)
         );
  OR2_X1 U9046 ( .A1(n10780), .A2(n7250), .ZN(n7790) );
  OAI21_X1 U9047 ( .B1(n9781), .B2(n7791), .A(n7790), .ZN(P2_U3462) );
  INV_X1 U9048 ( .A(n7792), .ZN(n7814) );
  AOI22_X1 U9049 ( .A1(n10096), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10477), .ZN(n7793) );
  OAI21_X1 U9050 ( .B1(n7814), .B2(n10492), .A(n7793), .ZN(P1_U3338) );
  AOI21_X1 U9051 ( .B1(n7795), .B2(n7794), .A(n7904), .ZN(n7799) );
  INV_X1 U9052 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n8861) );
  NOR2_X1 U9053 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8861), .ZN(n10594) );
  OAI22_X1 U9054 ( .A1(n7824), .A2(n9113), .B1(n8070), .B2(n9134), .ZN(n7796)
         );
  AOI211_X1 U9055 ( .C1(n9079), .C2(n7966), .A(n10594), .B(n7796), .ZN(n7798)
         );
  NAND2_X1 U9056 ( .A1(n9136), .A2(n7965), .ZN(n7797) );
  OAI211_X1 U9057 ( .C1(n7799), .C2(n9127), .A(n7798), .B(n7797), .ZN(P2_U3170) );
  AOI21_X1 U9058 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n7801), .A(n7800), .ZN(
        n7804) );
  NAND2_X1 U9059 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n8146), .ZN(n7802) );
  OAI21_X1 U9060 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n8146), .A(n7802), .ZN(
        n7803) );
  NOR2_X1 U9061 ( .A1(n7804), .A2(n7803), .ZN(n8145) );
  AOI211_X1 U9062 ( .C1(n7804), .C2(n7803), .A(n8145), .B(n10122), .ZN(n7813)
         );
  XNOR2_X1 U9063 ( .A(n8151), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n7808) );
  OAI21_X1 U9064 ( .B1(n7806), .B2(n8606), .A(n7805), .ZN(n7807) );
  NAND2_X1 U9065 ( .A1(n7808), .A2(n7807), .ZN(n8149) );
  OAI211_X1 U9066 ( .C1(n7808), .C2(n7807), .A(n10120), .B(n8149), .ZN(n7811)
         );
  NOR2_X1 U9067 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7809), .ZN(n9862) );
  AOI21_X1 U9068 ( .B1(n10560), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n9862), .ZN(
        n7810) );
  OAI211_X1 U9069 ( .C1(n10117), .C2(n8151), .A(n7811), .B(n7810), .ZN(n7812)
         );
  OR2_X1 U9070 ( .A1(n7813), .A2(n7812), .ZN(P1_U3257) );
  INV_X1 U9071 ( .A(n10738), .ZN(n9455) );
  OAI222_X1 U9072 ( .A1(n9455), .A2(P2_U3151), .B1(n9855), .B2(n7815), .C1(
        n7814), .C2(n9856), .ZN(P2_U3278) );
  INV_X1 U9073 ( .A(n9155), .ZN(n9165) );
  INV_X1 U9074 ( .A(n7816), .ZN(n7817) );
  NAND3_X1 U9075 ( .A1(n7818), .A2(n9165), .A3(n7817), .ZN(n7820) );
  NAND2_X1 U9076 ( .A1(n7820), .A2(n7819), .ZN(n7962) );
  NOR2_X1 U9077 ( .A1(n7821), .A2(n9773), .ZN(n7825) );
  XOR2_X1 U9078 ( .A(n7816), .B(n7822), .Z(n7823) );
  OAI222_X1 U9079 ( .A1(n9685), .A2(n8070), .B1(n9684), .B2(n7824), .C1(n7823), 
        .C2(n9682), .ZN(n7963) );
  AOI211_X1 U9080 ( .C1(n9778), .C2(n7962), .A(n7825), .B(n7963), .ZN(n10782)
         );
  NAND2_X1 U9081 ( .A1(n7250), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7826) );
  OAI21_X1 U9082 ( .B1(n10782), .B2(n7250), .A(n7826), .ZN(P2_U3463) );
  NOR2_X1 U9083 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n7827) );
  AOI21_X1 U9084 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(P2_ADDR_REG_18__SCAN_IN), 
        .A(n7827), .ZN(n10552) );
  NOR2_X1 U9085 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7828) );
  AOI21_X1 U9086 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7828), .ZN(n10549) );
  NOR2_X1 U9087 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7829) );
  AOI21_X1 U9088 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7829), .ZN(n10546) );
  NOR2_X1 U9089 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7830) );
  AOI21_X1 U9090 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7830), .ZN(n10543) );
  NOR2_X1 U9091 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7831) );
  AOI21_X1 U9092 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7831), .ZN(n10540) );
  NOR2_X1 U9093 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7832) );
  AOI21_X1 U9094 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7832), .ZN(n10537) );
  NOR2_X1 U9095 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7833) );
  AOI21_X1 U9096 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7833), .ZN(n10534) );
  NOR2_X1 U9097 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7834) );
  AOI21_X1 U9098 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7834), .ZN(n10531) );
  NOR2_X1 U9099 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7835) );
  AOI21_X1 U9100 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7835), .ZN(n10528) );
  NOR2_X1 U9101 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7836) );
  AOI21_X1 U9102 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7836), .ZN(n10525) );
  NOR2_X1 U9103 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7837) );
  AOI21_X1 U9104 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7837), .ZN(n10522) );
  NOR2_X1 U9105 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7838) );
  AOI21_X1 U9106 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7838), .ZN(n10519) );
  NOR2_X1 U9107 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7839) );
  AOI21_X1 U9108 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7839), .ZN(n10516) );
  NOR2_X1 U9109 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7840) );
  AOI21_X1 U9110 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7840), .ZN(n10513) );
  AND2_X1 U9111 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .ZN(n7841) );
  NOR2_X1 U9112 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7841), .ZN(n10499) );
  INV_X1 U9113 ( .A(n10499), .ZN(n10500) );
  INV_X1 U9114 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10588) );
  NAND3_X1 U9115 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10501) );
  NAND2_X1 U9116 ( .A1(n10588), .A2(n10501), .ZN(n10498) );
  NAND2_X1 U9117 ( .A1(n10500), .A2(n10498), .ZN(n10504) );
  NAND2_X1 U9118 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7842) );
  OAI21_X1 U9119 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7842), .ZN(n10503) );
  NOR2_X1 U9120 ( .A1(n10504), .A2(n10503), .ZN(n10502) );
  AOI21_X1 U9121 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10502), .ZN(n10507) );
  NAND2_X1 U9122 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7843) );
  OAI21_X1 U9123 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n7843), .ZN(n10506) );
  NOR2_X1 U9124 ( .A1(n10507), .A2(n10506), .ZN(n10505) );
  AOI21_X1 U9125 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10505), .ZN(n10510) );
  NOR2_X1 U9126 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7844) );
  AOI21_X1 U9127 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7844), .ZN(n10509) );
  NAND2_X1 U9128 ( .A1(n10510), .A2(n10509), .ZN(n10508) );
  OAI21_X1 U9129 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10508), .ZN(n10512) );
  NAND2_X1 U9130 ( .A1(n10513), .A2(n10512), .ZN(n10511) );
  OAI21_X1 U9131 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10511), .ZN(n10515) );
  NAND2_X1 U9132 ( .A1(n10516), .A2(n10515), .ZN(n10514) );
  OAI21_X1 U9133 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10514), .ZN(n10518) );
  NAND2_X1 U9134 ( .A1(n10519), .A2(n10518), .ZN(n10517) );
  OAI21_X1 U9135 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10517), .ZN(n10521) );
  NAND2_X1 U9136 ( .A1(n10522), .A2(n10521), .ZN(n10520) );
  OAI21_X1 U9137 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10520), .ZN(n10524) );
  NAND2_X1 U9138 ( .A1(n10525), .A2(n10524), .ZN(n10523) );
  OAI21_X1 U9139 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10523), .ZN(n10527) );
  NAND2_X1 U9140 ( .A1(n10528), .A2(n10527), .ZN(n10526) );
  OAI21_X1 U9141 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10526), .ZN(n10530) );
  NAND2_X1 U9142 ( .A1(n10531), .A2(n10530), .ZN(n10529) );
  OAI21_X1 U9143 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10529), .ZN(n10533) );
  NAND2_X1 U9144 ( .A1(n10534), .A2(n10533), .ZN(n10532) );
  OAI21_X1 U9145 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10532), .ZN(n10536) );
  NAND2_X1 U9146 ( .A1(n10537), .A2(n10536), .ZN(n10535) );
  OAI21_X1 U9147 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10535), .ZN(n10539) );
  NAND2_X1 U9148 ( .A1(n10540), .A2(n10539), .ZN(n10538) );
  OAI21_X1 U9149 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10538), .ZN(n10542) );
  NAND2_X1 U9150 ( .A1(n10543), .A2(n10542), .ZN(n10541) );
  OAI21_X1 U9151 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10541), .ZN(n10545) );
  NAND2_X1 U9152 ( .A1(n10546), .A2(n10545), .ZN(n10544) );
  OAI21_X1 U9153 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10544), .ZN(n10548) );
  NAND2_X1 U9154 ( .A1(n10549), .A2(n10548), .ZN(n10547) );
  OAI21_X1 U9155 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10547), .ZN(n10551) );
  NAND2_X1 U9156 ( .A1(n10552), .A2(n10551), .ZN(n10550) );
  OAI21_X1 U9157 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(P1_ADDR_REG_18__SCAN_IN), 
        .A(n10550), .ZN(n7847) );
  XNOR2_X1 U9158 ( .A(n7845), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7846) );
  XNOR2_X1 U9159 ( .A(n7847), .B(n7846), .ZN(ADD_1068_U4) );
  INV_X1 U9160 ( .A(n10015), .ZN(n10005) );
  AND2_X1 U9161 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10057) );
  OAI22_X1 U9162 ( .A1(n7848), .A2(n10009), .B1(n9991), .B2(n8139), .ZN(n7849)
         );
  AOI211_X1 U9163 ( .C1(n10003), .C2(n10043), .A(n10057), .B(n7849), .ZN(n7854) );
  XNOR2_X1 U9164 ( .A(n7851), .B(n7850), .ZN(n7852) );
  NAND2_X1 U9165 ( .A1(n7852), .A2(n10002), .ZN(n7853) );
  OAI211_X1 U9166 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n10005), .A(n7854), .B(
        n7853), .ZN(P1_U3218) );
  INV_X1 U9167 ( .A(n7942), .ZN(n7863) );
  AOI21_X1 U9168 ( .B1(n7855), .B2(n7856), .A(n10026), .ZN(n7858) );
  NAND2_X1 U9169 ( .A1(n7858), .A2(n7857), .ZN(n7862) );
  OAI22_X1 U9170 ( .A1(n10784), .A2(n10009), .B1(n9991), .B2(n8107), .ZN(n7859) );
  AOI211_X1 U9171 ( .C1(n10003), .C2(n10042), .A(n7860), .B(n7859), .ZN(n7861)
         );
  OAI211_X1 U9172 ( .C1(n10005), .C2(n7863), .A(n7862), .B(n7861), .ZN(
        P1_U3230) );
  OAI21_X1 U9173 ( .B1(n7865), .B2(n9332), .A(n7864), .ZN(n7918) );
  XNOR2_X1 U9174 ( .A(n7866), .B(n9332), .ZN(n7867) );
  OAI222_X1 U9175 ( .A1(n9684), .A2(n7908), .B1(n9685), .B2(n7907), .C1(n9682), 
        .C2(n7867), .ZN(n7913) );
  AOI21_X1 U9176 ( .B1(n9778), .B2(n7918), .A(n7913), .ZN(n7875) );
  INV_X1 U9177 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7868) );
  OAI22_X1 U9178 ( .A1(n9833), .A2(n7872), .B1(n10851), .B2(n7868), .ZN(n7869)
         );
  INV_X1 U9179 ( .A(n7869), .ZN(n7870) );
  OAI21_X1 U9180 ( .B1(n7875), .B2(n7244), .A(n7870), .ZN(P2_U3405) );
  INV_X1 U9181 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7871) );
  OAI22_X1 U9182 ( .A1(n9753), .A2(n7872), .B1(n9781), .B2(n7871), .ZN(n7873)
         );
  INV_X1 U9183 ( .A(n7873), .ZN(n7874) );
  OAI21_X1 U9184 ( .B1(n7875), .B2(n7250), .A(n7874), .ZN(P2_U3464) );
  NAND2_X1 U9185 ( .A1(n10766), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7876) );
  OAI21_X1 U9186 ( .B1(n8988), .B2(n10766), .A(n7876), .ZN(P2_U3520) );
  AND2_X1 U9187 ( .A1(n7259), .A2(n7262), .ZN(n9478) );
  INV_X1 U9188 ( .A(n9478), .ZN(n7877) );
  NAND2_X1 U9189 ( .A1(n7878), .A2(n7877), .ZN(n7879) );
  OAI22_X1 U9190 ( .A1(n9652), .A2(n7880), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9669), .ZN(n7883) );
  MUX2_X1 U9191 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n7881), .S(n9672), .Z(n7882)
         );
  AOI211_X1 U9192 ( .C1(n9692), .C2(n7884), .A(n7883), .B(n7882), .ZN(n7885)
         );
  INV_X1 U9193 ( .A(n7885), .ZN(P2_U3230) );
  NAND2_X1 U9194 ( .A1(n7887), .A2(n7886), .ZN(n7889) );
  XNOR2_X1 U9195 ( .A(n7889), .B(n7888), .ZN(n7894) );
  AND2_X1 U9196 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10075) );
  OAI22_X1 U9197 ( .A1(n7890), .A2(n10009), .B1(n9991), .B2(n8243), .ZN(n7891)
         );
  AOI211_X1 U9198 ( .C1(n10003), .C2(n10041), .A(n10075), .B(n7891), .ZN(n7893) );
  NAND2_X1 U9199 ( .A1(n10015), .A2(n8162), .ZN(n7892) );
  OAI211_X1 U9200 ( .C1(n7894), .C2(n10026), .A(n7893), .B(n7892), .ZN(
        P1_U3227) );
  NOR2_X1 U9201 ( .A1(n7895), .A2(n9678), .ZN(n7897) );
  AOI211_X1 U9202 ( .C1(n9688), .C2(P2_REG3_REG_2__SCAN_IN), .A(n7897), .B(
        n7896), .ZN(n7898) );
  MUX2_X1 U9203 ( .A(n5440), .B(n7898), .S(n9672), .Z(n7899) );
  OAI21_X1 U9204 ( .B1(n9676), .B2(n7900), .A(n7899), .ZN(P2_U3231) );
  INV_X1 U9205 ( .A(n7914), .ZN(n7912) );
  INV_X1 U9206 ( .A(n7901), .ZN(n7906) );
  NOR3_X1 U9207 ( .A1(n7904), .A2(n7903), .A3(n7902), .ZN(n7905) );
  OAI21_X1 U9208 ( .B1(n7906), .B2(n7905), .A(n9109), .ZN(n7911) );
  AND2_X1 U9209 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10616) );
  OAI22_X1 U9210 ( .A1(n7908), .A2(n9113), .B1(n7907), .B2(n9134), .ZN(n7909)
         );
  AOI211_X1 U9211 ( .C1(n9079), .C2(n7915), .A(n10616), .B(n7909), .ZN(n7910)
         );
  OAI211_X1 U9212 ( .C1(n7912), .C2(n8057), .A(n7911), .B(n7910), .ZN(P2_U3167) );
  INV_X1 U9213 ( .A(n7913), .ZN(n7920) );
  AOI22_X1 U9214 ( .A1(n8536), .A2(n7915), .B1(n9688), .B2(n7914), .ZN(n7916)
         );
  OAI21_X1 U9215 ( .B1(n10612), .B2(n9672), .A(n7916), .ZN(n7917) );
  AOI21_X1 U9216 ( .B1(n7918), .B2(n9692), .A(n7917), .ZN(n7919) );
  OAI21_X1 U9217 ( .B1(n7920), .B2(n9694), .A(n7919), .ZN(P2_U3228) );
  INV_X1 U9218 ( .A(n7921), .ZN(n7926) );
  AOI22_X1 U9219 ( .A1(n8536), .A2(n7265), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9688), .ZN(n7922) );
  OAI21_X1 U9220 ( .B1(n10575), .B2(n9672), .A(n7922), .ZN(n7923) );
  AOI21_X1 U9221 ( .B1(n7924), .B2(n9692), .A(n7923), .ZN(n7925) );
  OAI21_X1 U9222 ( .B1(n7926), .B2(n9694), .A(n7925), .ZN(P2_U3232) );
  INV_X1 U9223 ( .A(n10767), .ZN(n10771) );
  INV_X1 U9224 ( .A(n7927), .ZN(n7929) );
  INV_X1 U9225 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7928) );
  OAI222_X1 U9226 ( .A1(P2_U3151), .A2(n10771), .B1(n9856), .B2(n7929), .C1(
        n7928), .C2(n9855), .ZN(P2_U3277) );
  INV_X1 U9227 ( .A(n10111), .ZN(n10105) );
  OAI222_X1 U9228 ( .A1(P1_U3086), .A2(n10105), .B1(n10494), .B2(n7930), .C1(
        n7929), .C2(n10492), .ZN(P1_U3337) );
  INV_X1 U9229 ( .A(n7931), .ZN(n7933) );
  NAND3_X1 U9230 ( .A1(n7933), .A2(n7932), .A3(n7970), .ZN(n7941) );
  INV_X1 U9231 ( .A(n7934), .ZN(n7935) );
  NAND2_X1 U9232 ( .A1(n10328), .A2(n7935), .ZN(n8639) );
  INV_X1 U9233 ( .A(n7936), .ZN(n8633) );
  NAND2_X1 U9234 ( .A1(n10328), .A2(n8633), .ZN(n7937) );
  OAI21_X1 U9235 ( .B1(n7939), .B2(n7945), .A(n7938), .ZN(n10787) );
  OAI211_X1 U9236 ( .C1(n8085), .C2(n10784), .A(n8136), .B(n10292), .ZN(n10783) );
  INV_X1 U9237 ( .A(n10783), .ZN(n7943) );
  INV_X2 U9238 ( .A(n10326), .ZN(n10274) );
  AOI22_X1 U9239 ( .A1(n7943), .A2(n10286), .B1(n7942), .B2(n10274), .ZN(n7944) );
  OAI21_X1 U9240 ( .B1(n10784), .B2(n10325), .A(n7944), .ZN(n7949) );
  XNOR2_X1 U9241 ( .A(n7946), .B(n7945), .ZN(n7947) );
  INV_X1 U9242 ( .A(n10312), .ZN(n8902) );
  OAI222_X1 U9243 ( .A1(n10315), .A2(n8107), .B1(n10395), .B2(n8129), .C1(
        n7947), .C2(n8902), .ZN(n10785) );
  MUX2_X1 U9244 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10785), .S(n10328), .Z(n7948) );
  AOI211_X1 U9245 ( .C1(n10321), .C2(n10787), .A(n7949), .B(n7948), .ZN(n7950)
         );
  INV_X1 U9246 ( .A(n7950), .ZN(P1_U3289) );
  XOR2_X1 U9247 ( .A(n7951), .B(n7952), .Z(n7957) );
  OAI22_X1 U9248 ( .A1(n10795), .A2(n10009), .B1(n9991), .B2(n8229), .ZN(n7953) );
  AOI211_X1 U9249 ( .C1(n10003), .C2(n10040), .A(n7954), .B(n7953), .ZN(n7956)
         );
  NAND2_X1 U9250 ( .A1(n10015), .A2(n8113), .ZN(n7955) );
  OAI211_X1 U9251 ( .C1(n7957), .C2(n10026), .A(n7956), .B(n7955), .ZN(
        P1_U3239) );
  INV_X1 U9252 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7961) );
  OAI21_X1 U9253 ( .B1(n10312), .B2(n10838), .A(n8012), .ZN(n7959) );
  NOR2_X1 U9254 ( .A1(n8126), .A2(n10315), .ZN(n8013) );
  INV_X1 U9255 ( .A(n8013), .ZN(n7958) );
  OAI211_X1 U9256 ( .C1(n8011), .C2(n8075), .A(n7959), .B(n7958), .ZN(n7972)
         );
  NAND2_X1 U9257 ( .A1(n7972), .A2(n10846), .ZN(n7960) );
  OAI21_X1 U9258 ( .B1(n10846), .B2(n7961), .A(n7960), .ZN(P1_U3453) );
  INV_X1 U9259 ( .A(n7962), .ZN(n7969) );
  INV_X1 U9260 ( .A(n7963), .ZN(n7964) );
  MUX2_X1 U9261 ( .A(n7651), .B(n7964), .S(n9672), .Z(n7968) );
  AOI22_X1 U9262 ( .A1(n8536), .A2(n7966), .B1(n9688), .B2(n7965), .ZN(n7967)
         );
  OAI211_X1 U9263 ( .C1(n7969), .C2(n9676), .A(n7968), .B(n7967), .ZN(P2_U3229) );
  NAND2_X1 U9264 ( .A1(n7972), .A2(n10842), .ZN(n7973) );
  OAI21_X1 U9265 ( .B1(n10842), .B2(n6957), .A(n7973), .ZN(P1_U3522) );
  INV_X1 U9266 ( .A(n7974), .ZN(n8934) );
  OAI222_X1 U9267 ( .A1(n7976), .A2(P2_U3151), .B1(n9856), .B2(n8934), .C1(
        n9855), .C2(n7975), .ZN(P2_U3276) );
  NOR2_X1 U9268 ( .A1(n7979), .A2(n7980), .ZN(n7981) );
  INV_X1 U9269 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n8035) );
  NOR2_X1 U9270 ( .A1(n8035), .A2(n8036), .ZN(n8034) );
  NAND2_X1 U9271 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n8308), .ZN(n7982) );
  OAI21_X1 U9272 ( .B1(n8308), .B2(P2_REG2_REG_8__SCAN_IN), .A(n7982), .ZN(
        n7983) );
  AOI21_X1 U9273 ( .B1(n7984), .B2(n7983), .A(n8307), .ZN(n8009) );
  MUX2_X1 U9274 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n6601), .Z(n7985) );
  NOR2_X1 U9275 ( .A1(n7985), .A2(n8308), .ZN(n8304) );
  AOI21_X1 U9276 ( .B1(n7985), .B2(n8308), .A(n8304), .ZN(n7986) );
  INV_X1 U9277 ( .A(n7986), .ZN(n7993) );
  MUX2_X1 U9278 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n6601), .Z(n7989) );
  NOR2_X1 U9279 ( .A1(n7989), .A2(n5059), .ZN(n7991) );
  NOR2_X1 U9280 ( .A1(n7988), .A2(n7987), .ZN(n8040) );
  AOI21_X1 U9281 ( .B1(n7989), .B2(n5059), .A(n7991), .ZN(n7990) );
  INV_X1 U9282 ( .A(n7990), .ZN(n8041) );
  NOR2_X1 U9283 ( .A1(n8040), .A2(n8041), .ZN(n8039) );
  NOR2_X1 U9284 ( .A1(n7991), .A2(n8039), .ZN(n7992) );
  NOR2_X1 U9285 ( .A1(n7992), .A2(n7993), .ZN(n8303) );
  AOI21_X1 U9286 ( .B1(n7993), .B2(n7992), .A(n8303), .ZN(n7996) );
  NAND2_X1 U9287 ( .A1(n10757), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7995) );
  OAI211_X1 U9288 ( .C1(n7996), .C2(n8314), .A(n7995), .B(n7994), .ZN(n7997)
         );
  AOI21_X1 U9289 ( .B1(n7998), .B2(n10737), .A(n7997), .ZN(n8008) );
  INV_X1 U9290 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n8195) );
  AOI22_X1 U9291 ( .A1(n7998), .A2(n8195), .B1(P2_REG1_REG_8__SCAN_IN), .B2(
        n8308), .ZN(n8005) );
  NAND2_X1 U9292 ( .A1(n5059), .A2(n8002), .ZN(n8003) );
  NAND2_X1 U9293 ( .A1(P2_REG1_REG_7__SCAN_IN), .A2(n8038), .ZN(n8037) );
  OAI21_X1 U9294 ( .B1(n8005), .B2(n8004), .A(n8296), .ZN(n8006) );
  NAND2_X1 U9295 ( .A1(n8006), .A2(n10745), .ZN(n8007) );
  OAI211_X1 U9296 ( .C1(n8009), .C2(n10747), .A(n8008), .B(n8007), .ZN(
        P2_U3190) );
  NOR2_X1 U9297 ( .A1(n10264), .A2(n10803), .ZN(n10178) );
  OAI21_X1 U9298 ( .B1(n10178), .B2(n10297), .A(n8010), .ZN(n8022) );
  AND2_X1 U9299 ( .A1(n8012), .A2(n8011), .ZN(n8015) );
  INV_X1 U9300 ( .A(n8015), .ZN(n8018) );
  AOI21_X1 U9301 ( .B1(n10274), .B2(P1_REG3_REG_0__SCAN_IN), .A(n8013), .ZN(
        n8017) );
  NAND2_X1 U9302 ( .A1(n8015), .A2(n8014), .ZN(n8016) );
  OAI211_X1 U9303 ( .C1(n8019), .C2(n8018), .A(n8017), .B(n8016), .ZN(n8020)
         );
  NAND2_X1 U9304 ( .A1(n8020), .A2(n10328), .ZN(n8021) );
  OAI211_X1 U9305 ( .C1(n10555), .C2(n10328), .A(n8022), .B(n8021), .ZN(
        P1_U3293) );
  XNOR2_X1 U9306 ( .A(n8023), .B(n9336), .ZN(n8024) );
  AOI222_X1 U9307 ( .A1(n7237), .A2(n8024), .B1(n9387), .B2(n9541), .C1(n9389), 
        .C2(n9540), .ZN(n8206) );
  INV_X1 U9308 ( .A(n8179), .ZN(n8025) );
  OAI22_X1 U9309 ( .A1(n9672), .A2(n8035), .B1(n8025), .B2(n9669), .ZN(n8032)
         );
  INV_X1 U9310 ( .A(n8026), .ZN(n8028) );
  OAI21_X1 U9311 ( .B1(n8028), .B2(n8027), .A(n9336), .ZN(n8030) );
  NAND2_X1 U9312 ( .A1(n8030), .A2(n8029), .ZN(n8207) );
  NOR2_X1 U9313 ( .A1(n8207), .A2(n9676), .ZN(n8031) );
  AOI211_X1 U9314 ( .C1(n8536), .C2(n8180), .A(n8032), .B(n8031), .ZN(n8033)
         );
  OAI21_X1 U9315 ( .B1(n8206), .B2(n9694), .A(n8033), .ZN(P2_U3226) );
  AOI21_X1 U9316 ( .B1(n8036), .B2(n8035), .A(n8034), .ZN(n8048) );
  OAI21_X1 U9317 ( .B1(P2_REG1_REG_7__SCAN_IN), .B2(n8038), .A(n8037), .ZN(
        n8046) );
  INV_X1 U9318 ( .A(n10737), .ZN(n10765) );
  INV_X1 U9319 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8752) );
  NOR2_X1 U9320 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8752), .ZN(n8178) );
  AOI21_X1 U9321 ( .B1(n8041), .B2(n8040), .A(n8039), .ZN(n8042) );
  NOR2_X1 U9322 ( .A1(n8042), .A2(n8314), .ZN(n8043) );
  AOI211_X1 U9323 ( .C1(n10757), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n8178), .B(
        n8043), .ZN(n8044) );
  OAI21_X1 U9324 ( .B1(n5059), .B2(n10765), .A(n8044), .ZN(n8045) );
  AOI21_X1 U9325 ( .B1(n10745), .B2(n8046), .A(n8045), .ZN(n8047) );
  OAI21_X1 U9326 ( .B1(n8048), .B2(n10747), .A(n8047), .ZN(P2_U3189) );
  INV_X1 U9327 ( .A(n8097), .ZN(n8058) );
  AOI211_X1 U9328 ( .C1(n8051), .C2(n8050), .A(n9127), .B(n8049), .ZN(n8052)
         );
  INV_X1 U9329 ( .A(n8052), .ZN(n8056) );
  OAI22_X1 U9330 ( .A1(n8191), .A2(n9134), .B1(n9139), .B2(n8067), .ZN(n8053)
         );
  AOI211_X1 U9331 ( .C1(n9132), .C2(n9390), .A(n8054), .B(n8053), .ZN(n8055)
         );
  OAI211_X1 U9332 ( .C1(n8058), .C2(n8057), .A(n8056), .B(n8055), .ZN(P2_U3179) );
  XOR2_X1 U9333 ( .A(n8059), .B(n8060), .Z(n8065) );
  OAI22_X1 U9334 ( .A1(n8370), .A2(n10009), .B1(n9991), .B2(n8385), .ZN(n8061)
         );
  AOI211_X1 U9335 ( .C1(n10003), .C2(n10039), .A(n8062), .B(n8061), .ZN(n8064)
         );
  NAND2_X1 U9336 ( .A1(n10015), .A2(n8368), .ZN(n8063) );
  OAI211_X1 U9337 ( .C1(n8065), .C2(n10026), .A(n8064), .B(n8063), .ZN(
        P1_U3213) );
  OAI21_X1 U9338 ( .B1(n8066), .B2(n9329), .A(n8026), .ZN(n8094) );
  NOR2_X1 U9339 ( .A1(n8067), .A2(n9773), .ZN(n8071) );
  XOR2_X1 U9340 ( .A(n9329), .B(n8068), .Z(n8069) );
  OAI222_X1 U9341 ( .A1(n9685), .A2(n8191), .B1(n9684), .B2(n8070), .C1(n8069), 
        .C2(n9682), .ZN(n8095) );
  AOI211_X1 U9342 ( .C1(n9778), .C2(n8094), .A(n8071), .B(n8095), .ZN(n10792)
         );
  NAND2_X1 U9343 ( .A1(n7250), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8072) );
  OAI21_X1 U9344 ( .B1(n10792), .B2(n7250), .A(n8072), .ZN(P2_U3465) );
  INV_X1 U9345 ( .A(n6960), .ZN(n8077) );
  OAI211_X1 U9346 ( .C1(n8076), .C2(n8075), .A(n10292), .B(n8123), .ZN(n8341)
         );
  OAI21_X1 U9347 ( .B1(n8077), .B2(n10395), .A(n8341), .ZN(n8081) );
  XNOR2_X1 U9348 ( .A(n8079), .B(n8078), .ZN(n8080) );
  OAI22_X1 U9349 ( .A1(n8080), .A2(n8902), .B1(n8088), .B2(n10315), .ZN(n8338)
         );
  AOI211_X1 U9350 ( .C1(n10838), .C2(n8343), .A(n8081), .B(n8338), .ZN(n8158)
         );
  AOI22_X1 U9351 ( .A1(n8435), .A2(n6967), .B1(n10843), .B2(
        P1_REG0_REG_1__SCAN_IN), .ZN(n8082) );
  OAI21_X1 U9352 ( .B1(n8158), .B2(n10843), .A(n8082), .ZN(P1_U3456) );
  OAI21_X1 U9353 ( .B1(n8084), .B2(n8089), .A(n8083), .ZN(n8353) );
  INV_X1 U9354 ( .A(n8085), .ZN(n8087) );
  AOI21_X1 U9355 ( .B1(n8125), .B2(n8347), .A(n10803), .ZN(n8086) );
  NAND2_X1 U9356 ( .A1(n8087), .A2(n8086), .ZN(n8351) );
  OAI21_X1 U9357 ( .B1(n8088), .B2(n10395), .A(n8351), .ZN(n8092) );
  XNOR2_X1 U9358 ( .A(n8090), .B(n8089), .ZN(n8091) );
  OAI22_X1 U9359 ( .A1(n8091), .A2(n8902), .B1(n8139), .B2(n10315), .ZN(n8346)
         );
  AOI211_X1 U9360 ( .C1(n10838), .C2(n8353), .A(n8092), .B(n8346), .ZN(n8160)
         );
  AOI22_X1 U9361 ( .A1(n8435), .A2(n8347), .B1(n10843), .B2(
        P1_REG0_REG_3__SCAN_IN), .ZN(n8093) );
  OAI21_X1 U9362 ( .B1(n8160), .B2(n10843), .A(n8093), .ZN(P1_U3462) );
  INV_X1 U9363 ( .A(n8094), .ZN(n8101) );
  INV_X1 U9364 ( .A(n8095), .ZN(n8096) );
  MUX2_X1 U9365 ( .A(n7661), .B(n8096), .S(n9672), .Z(n8100) );
  AOI22_X1 U9366 ( .A1(n8536), .A2(n8098), .B1(n9688), .B2(n8097), .ZN(n8099)
         );
  OAI211_X1 U9367 ( .C1(n8101), .C2(n9676), .A(n8100), .B(n8099), .ZN(P2_U3227) );
  XNOR2_X1 U9368 ( .A(n8103), .B(n8102), .ZN(n8110) );
  OAI21_X1 U9369 ( .B1(n8106), .B2(n8105), .A(n8104), .ZN(n10798) );
  OAI22_X1 U9370 ( .A1(n8229), .A2(n10315), .B1(n8107), .B2(n10395), .ZN(n8108) );
  AOI21_X1 U9371 ( .B1(n10798), .B2(n8633), .A(n8108), .ZN(n8109) );
  OAI21_X1 U9372 ( .B1(n8902), .B2(n8110), .A(n8109), .ZN(n10796) );
  INV_X1 U9373 ( .A(n10796), .ZN(n8120) );
  INV_X1 U9374 ( .A(n8639), .ZN(n8118) );
  INV_X1 U9375 ( .A(n8137), .ZN(n8112) );
  INV_X1 U9376 ( .A(n8111), .ZN(n8252) );
  OAI211_X1 U9377 ( .C1(n10795), .C2(n8112), .A(n8252), .B(n10292), .ZN(n10794) );
  AOI22_X1 U9378 ( .A1(n10335), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n8113), .B2(
        n10274), .ZN(n8116) );
  NAND2_X1 U9379 ( .A1(n10297), .A2(n8114), .ZN(n8115) );
  OAI211_X1 U9380 ( .C1(n10794), .C2(n10264), .A(n8116), .B(n8115), .ZN(n8117)
         );
  AOI21_X1 U9381 ( .B1(n10798), .B2(n8118), .A(n8117), .ZN(n8119) );
  OAI21_X1 U9382 ( .B1(n8120), .B2(n10335), .A(n8119), .ZN(P1_U3287) );
  OAI21_X1 U9383 ( .B1(n8122), .B2(n8128), .A(n8121), .ZN(n8335) );
  NAND2_X1 U9384 ( .A1(n8123), .A2(n6945), .ZN(n8124) );
  NAND3_X1 U9385 ( .A1(n8125), .A2(n10292), .A3(n8124), .ZN(n8333) );
  OAI21_X1 U9386 ( .B1(n8126), .B2(n10395), .A(n8333), .ZN(n8131) );
  XNOR2_X1 U9387 ( .A(n8128), .B(n8127), .ZN(n8130) );
  OAI22_X1 U9388 ( .A1(n8130), .A2(n8902), .B1(n8129), .B2(n10315), .ZN(n8330)
         );
  AOI211_X1 U9389 ( .C1(n10838), .C2(n8335), .A(n8131), .B(n8330), .ZN(n8171)
         );
  AOI22_X1 U9390 ( .A1(n8435), .A2(n6945), .B1(n10843), .B2(
        P1_REG0_REG_2__SCAN_IN), .ZN(n8132) );
  OAI21_X1 U9391 ( .B1(n8171), .B2(n10843), .A(n8132), .ZN(P1_U3459) );
  OAI21_X1 U9392 ( .B1(n8135), .B2(n8134), .A(n8133), .ZN(n8167) );
  AOI21_X1 U9393 ( .B1(n8136), .B2(n8172), .A(n10803), .ZN(n8138) );
  NAND2_X1 U9394 ( .A1(n8138), .A2(n8137), .ZN(n8165) );
  OAI21_X1 U9395 ( .B1(n8139), .B2(n10395), .A(n8165), .ZN(n8143) );
  XNOR2_X1 U9396 ( .A(n8141), .B(n8140), .ZN(n8142) );
  OAI22_X1 U9397 ( .A1(n8142), .A2(n8902), .B1(n8243), .B2(n10315), .ZN(n8161)
         );
  AOI211_X1 U9398 ( .C1(n10838), .C2(n8167), .A(n8143), .B(n8161), .ZN(n8174)
         );
  AOI22_X1 U9399 ( .A1(n8435), .A2(n8172), .B1(n10843), .B2(
        P1_REG0_REG_5__SCAN_IN), .ZN(n8144) );
  OAI21_X1 U9400 ( .B1(n8174), .B2(n10843), .A(n8144), .ZN(P1_U3468) );
  INV_X1 U9401 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8148) );
  AOI21_X1 U9402 ( .B1(n8146), .B2(P1_REG2_REG_14__SCAN_IN), .A(n8145), .ZN(
        n8448) );
  XNOR2_X1 U9403 ( .A(n8447), .B(n8448), .ZN(n8147) );
  NOR2_X1 U9404 ( .A1(n8148), .A2(n8147), .ZN(n8449) );
  AOI211_X1 U9405 ( .C1(n8148), .C2(n8147), .A(n8449), .B(n10122), .ZN(n8156)
         );
  INV_X1 U9406 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8150) );
  OAI21_X1 U9407 ( .B1(n8151), .B2(n8150), .A(n8149), .ZN(n8441) );
  XNOR2_X1 U9408 ( .A(n8447), .B(n8441), .ZN(n8152) );
  NAND2_X1 U9409 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n8152), .ZN(n8443) );
  OAI211_X1 U9410 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n8152), .A(n10120), .B(
        n8443), .ZN(n8154) );
  AND2_X1 U9411 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10016) );
  AOI21_X1 U9412 ( .B1(n10560), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n10016), .ZN(
        n8153) );
  OAI211_X1 U9413 ( .C1(n10117), .C2(n8447), .A(n8154), .B(n8153), .ZN(n8155)
         );
  OR2_X1 U9414 ( .A1(n8156), .A2(n8155), .ZN(P1_U3258) );
  AOI22_X1 U9415 ( .A1(n8917), .A2(n6967), .B1(n10840), .B2(
        P1_REG1_REG_1__SCAN_IN), .ZN(n8157) );
  OAI21_X1 U9416 ( .B1(n8158), .B2(n10840), .A(n8157), .ZN(P1_U3523) );
  AOI22_X1 U9417 ( .A1(n8917), .A2(n8347), .B1(n10840), .B2(
        P1_REG1_REG_3__SCAN_IN), .ZN(n8159) );
  OAI21_X1 U9418 ( .B1(n8160), .B2(n10840), .A(n8159), .ZN(P1_U3525) );
  INV_X1 U9419 ( .A(n8161), .ZN(n8169) );
  AND2_X1 U9420 ( .A1(n10328), .A2(n10389), .ZN(n10159) );
  AOI22_X1 U9421 ( .A1(n10297), .A2(n8172), .B1(n10159), .B2(n10041), .ZN(
        n8164) );
  AOI22_X1 U9422 ( .A1(n10335), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n8162), .B2(
        n10274), .ZN(n8163) );
  OAI211_X1 U9423 ( .C1(n10264), .C2(n8165), .A(n8164), .B(n8163), .ZN(n8166)
         );
  AOI21_X1 U9424 ( .B1(n8167), .B2(n10321), .A(n8166), .ZN(n8168) );
  OAI21_X1 U9425 ( .B1(n8169), .B2(n10335), .A(n8168), .ZN(P1_U3288) );
  AOI22_X1 U9426 ( .A1(n8917), .A2(n6945), .B1(n10840), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n8170) );
  OAI21_X1 U9427 ( .B1(n8171), .B2(n10840), .A(n8170), .ZN(P1_U3524) );
  AOI22_X1 U9428 ( .A1(n8917), .A2(n8172), .B1(n10840), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n8173) );
  OAI21_X1 U9429 ( .B1(n8174), .B2(n10840), .A(n8173), .ZN(P1_U3527) );
  OAI21_X1 U9430 ( .B1(n8177), .B2(n8176), .A(n8175), .ZN(n8186) );
  AOI21_X1 U9431 ( .B1(n9389), .B2(n9132), .A(n8178), .ZN(n8184) );
  NAND2_X1 U9432 ( .A1(n9136), .A2(n8179), .ZN(n8183) );
  NAND2_X1 U9433 ( .A1(n9079), .A2(n8180), .ZN(n8182) );
  NAND2_X1 U9434 ( .A1(n9111), .A2(n9387), .ZN(n8181) );
  NAND4_X1 U9435 ( .A1(n8184), .A2(n8183), .A3(n8182), .A4(n8181), .ZN(n8185)
         );
  AOI21_X1 U9436 ( .B1(n8186), .B2(n9109), .A(n8185), .ZN(n8187) );
  INV_X1 U9437 ( .A(n8187), .ZN(P2_U3153) );
  INV_X1 U9438 ( .A(n8189), .ZN(n9337) );
  XNOR2_X1 U9439 ( .A(n8188), .B(n9337), .ZN(n8190) );
  OAI222_X1 U9440 ( .A1(n9685), .A2(n8577), .B1(n9684), .B2(n8191), .C1(n9682), 
        .C2(n8190), .ZN(n8197) );
  XNOR2_X1 U9441 ( .A(n8192), .B(n9337), .ZN(n8205) );
  OAI22_X1 U9442 ( .A1(n8205), .A2(n9766), .B1(n8193), .B2(n9773), .ZN(n8194)
         );
  NOR2_X1 U9443 ( .A1(n8197), .A2(n8194), .ZN(n10811) );
  OR2_X1 U9444 ( .A1(n9781), .A2(n8195), .ZN(n8196) );
  OAI21_X1 U9445 ( .B1(n10811), .B2(n7250), .A(n8196), .ZN(P2_U3467) );
  NAND2_X1 U9446 ( .A1(n8197), .A2(n9672), .ZN(n8204) );
  INV_X1 U9447 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n8200) );
  INV_X1 U9448 ( .A(n8198), .ZN(n8199) );
  OAI22_X1 U9449 ( .A1(n9672), .A2(n8200), .B1(n8199), .B2(n9669), .ZN(n8201)
         );
  AOI21_X1 U9450 ( .B1(n8536), .B2(n8202), .A(n8201), .ZN(n8203) );
  OAI211_X1 U9451 ( .C1(n8205), .C2(n9676), .A(n8204), .B(n8203), .ZN(P2_U3225) );
  OAI21_X1 U9452 ( .B1(n9766), .B2(n8207), .A(n8206), .ZN(n8214) );
  INV_X1 U9453 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n8208) );
  OAI22_X1 U9454 ( .A1(n9753), .A2(n8212), .B1(n9781), .B2(n8208), .ZN(n8209)
         );
  AOI21_X1 U9455 ( .B1(n8214), .B2(n9781), .A(n8209), .ZN(n8210) );
  INV_X1 U9456 ( .A(n8210), .ZN(P2_U3466) );
  INV_X1 U9457 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n8211) );
  OAI22_X1 U9458 ( .A1(n9833), .A2(n8212), .B1(n10851), .B2(n8211), .ZN(n8213)
         );
  AOI21_X1 U9459 ( .B1(n8214), .B2(n10851), .A(n8213), .ZN(n8215) );
  INV_X1 U9460 ( .A(n8215), .ZN(P2_U3411) );
  INV_X1 U9461 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8216) );
  OAI222_X1 U9462 ( .A1(P2_U3151), .A2(n9143), .B1(n9856), .B2(n8220), .C1(
        n8216), .C2(n9855), .ZN(P2_U3274) );
  INV_X1 U9463 ( .A(n8217), .ZN(n8914) );
  OAI222_X1 U9464 ( .A1(n10494), .A2(n8219), .B1(P1_U3086), .B2(n8218), .C1(
        n8914), .C2(n10492), .ZN(P1_U3335) );
  OAI222_X1 U9465 ( .A1(n10494), .A2(n8222), .B1(P1_U3086), .B2(n8221), .C1(
        n10492), .C2(n8220), .ZN(P1_U3334) );
  NAND3_X1 U9466 ( .A1(n8223), .A2(n8225), .A3(n8224), .ZN(n8280) );
  NAND2_X1 U9467 ( .A1(n8280), .A2(n8226), .ZN(n8227) );
  XNOR2_X1 U9468 ( .A(n8227), .B(n8231), .ZN(n8228) );
  OAI222_X1 U9469 ( .A1(n10315), .A2(n8494), .B1(n10395), .B2(n8229), .C1(
        n8228), .C2(n8902), .ZN(n10805) );
  INV_X1 U9470 ( .A(n10805), .ZN(n8240) );
  OAI21_X1 U9471 ( .B1(n8232), .B2(n8231), .A(n8230), .ZN(n10807) );
  OR2_X1 U9472 ( .A1(n8251), .A2(n10802), .ZN(n8233) );
  NAND2_X1 U9473 ( .A1(n8289), .A2(n8233), .ZN(n10804) );
  INV_X1 U9474 ( .A(n10178), .ZN(n8237) );
  AOI22_X1 U9475 ( .A1(n10335), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n8365), .B2(
        n10274), .ZN(n8236) );
  NAND2_X1 U9476 ( .A1(n10297), .A2(n8234), .ZN(n8235) );
  OAI211_X1 U9477 ( .C1(n10804), .C2(n8237), .A(n8236), .B(n8235), .ZN(n8238)
         );
  AOI21_X1 U9478 ( .B1(n10807), .B2(n10321), .A(n8238), .ZN(n8239) );
  OAI21_X1 U9479 ( .B1(n8240), .B2(n10335), .A(n8239), .ZN(P1_U3285) );
  OAI21_X1 U9480 ( .B1(n8242), .B2(n8244), .A(n8241), .ZN(n8250) );
  INV_X1 U9481 ( .A(n8250), .ZN(n8371) );
  OAI22_X1 U9482 ( .A1(n8243), .A2(n10395), .B1(n8385), .B2(n10315), .ZN(n8249) );
  INV_X1 U9483 ( .A(n8223), .ZN(n8246) );
  OAI21_X1 U9484 ( .B1(n8246), .B2(n8245), .A(n8244), .ZN(n8247) );
  AOI21_X1 U9485 ( .B1(n8247), .B2(n8280), .A(n8902), .ZN(n8248) );
  AOI211_X1 U9486 ( .C1(n8633), .C2(n8250), .A(n8249), .B(n8248), .ZN(n8376)
         );
  AOI21_X1 U9487 ( .B1(n8253), .B2(n8252), .A(n8251), .ZN(n8374) );
  AOI22_X1 U9488 ( .A1(n8374), .A2(n10292), .B1(n10428), .B2(n8253), .ZN(n8254) );
  OAI211_X1 U9489 ( .C1(n8371), .C2(n10793), .A(n8376), .B(n8254), .ZN(n8257)
         );
  NAND2_X1 U9490 ( .A1(n8257), .A2(n10842), .ZN(n8255) );
  OAI21_X1 U9491 ( .B1(n10842), .B2(n8256), .A(n8255), .ZN(P1_U3529) );
  INV_X1 U9492 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n8259) );
  NAND2_X1 U9493 ( .A1(n8257), .A2(n10846), .ZN(n8258) );
  OAI21_X1 U9494 ( .B1(n10846), .B2(n8259), .A(n8258), .ZN(P1_U3474) );
  OR2_X1 U9495 ( .A1(n8262), .A2(n8261), .ZN(n8263) );
  NAND2_X1 U9496 ( .A1(n8260), .A2(n8263), .ZN(n8265) );
  OAI22_X1 U9497 ( .A1(n8494), .A2(n10395), .B1(n8469), .B2(n10315), .ZN(n8264) );
  AOI21_X1 U9498 ( .B1(n8265), .B2(n10312), .A(n8264), .ZN(n10820) );
  OAI21_X1 U9499 ( .B1(n8268), .B2(n8267), .A(n8266), .ZN(n10823) );
  NAND2_X1 U9500 ( .A1(n10823), .A2(n10321), .ZN(n8277) );
  INV_X1 U9501 ( .A(n8269), .ZN(n10821) );
  INV_X1 U9502 ( .A(n8270), .ZN(n8272) );
  INV_X1 U9503 ( .A(n8398), .ZN(n8271) );
  OAI211_X1 U9504 ( .C1(n10821), .C2(n8272), .A(n8271), .B(n10292), .ZN(n10819) );
  INV_X1 U9505 ( .A(n10819), .ZN(n8275) );
  AOI22_X1 U9506 ( .A1(n10335), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n8497), .B2(
        n10274), .ZN(n8273) );
  OAI21_X1 U9507 ( .B1(n10821), .B2(n10325), .A(n8273), .ZN(n8274) );
  AOI21_X1 U9508 ( .B1(n8275), .B2(n10286), .A(n8274), .ZN(n8276) );
  OAI211_X1 U9509 ( .C1(n10335), .C2(n10820), .A(n8277), .B(n8276), .ZN(
        P1_U3283) );
  AOI21_X1 U9510 ( .B1(n8280), .B2(n8279), .A(n8278), .ZN(n8282) );
  XNOR2_X1 U9511 ( .A(n8282), .B(n8281), .ZN(n8284) );
  AOI22_X1 U9512 ( .A1(n8284), .A2(n10312), .B1(n10389), .B2(n8283), .ZN(
        n10813) );
  OAI21_X1 U9513 ( .B1(n8287), .B2(n8286), .A(n8285), .ZN(n10816) );
  NAND2_X1 U9514 ( .A1(n10816), .A2(n10321), .ZN(n8295) );
  INV_X1 U9515 ( .A(n8288), .ZN(n10814) );
  XNOR2_X1 U9516 ( .A(n8289), .B(n10814), .ZN(n8290) );
  AOI22_X1 U9517 ( .A1(n8290), .A2(n10292), .B1(n10282), .B2(n10037), .ZN(
        n10812) );
  INV_X1 U9518 ( .A(n10812), .ZN(n8293) );
  AOI22_X1 U9519 ( .A1(n10335), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n8388), .B2(
        n10274), .ZN(n8291) );
  OAI21_X1 U9520 ( .B1(n10814), .B2(n10325), .A(n8291), .ZN(n8292) );
  AOI21_X1 U9521 ( .B1(n8293), .B2(n10286), .A(n8292), .ZN(n8294) );
  OAI211_X1 U9522 ( .C1(n10335), .C2(n10813), .A(n8295), .B(n8294), .ZN(
        P1_U3284) );
  NAND2_X1 U9523 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n8308), .ZN(n8297) );
  NAND2_X1 U9524 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(n8298), .ZN(n9398) );
  OAI21_X1 U9525 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n8298), .A(n9398), .ZN(
        n8299) );
  NAND2_X1 U9526 ( .A1(n8299), .A2(n10745), .ZN(n8319) );
  NOR2_X1 U9527 ( .A1(n10765), .A2(n9397), .ZN(n8317) );
  MUX2_X1 U9528 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n6601), .Z(n8300) );
  INV_X1 U9529 ( .A(n8300), .ZN(n8302) );
  NOR2_X1 U9530 ( .A1(n8300), .A2(n9397), .ZN(n9444) );
  INV_X1 U9531 ( .A(n9444), .ZN(n8301) );
  OAI21_X1 U9532 ( .B1(n9413), .B2(n8302), .A(n8301), .ZN(n8306) );
  NOR2_X1 U9533 ( .A1(n8304), .A2(n8303), .ZN(n8305) );
  NOR2_X1 U9534 ( .A1(n8305), .A2(n8306), .ZN(n9443) );
  AOI21_X1 U9535 ( .B1(n8306), .B2(n8305), .A(n9443), .ZN(n8315) );
  INV_X1 U9536 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n8324) );
  AOI21_X1 U9537 ( .B1(n8309), .B2(n8324), .A(n9414), .ZN(n8311) );
  NOR2_X1 U9538 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6345), .ZN(n8422) );
  INV_X1 U9539 ( .A(n8422), .ZN(n8310) );
  OAI21_X1 U9540 ( .B1(n10747), .B2(n8311), .A(n8310), .ZN(n8312) );
  INV_X1 U9541 ( .A(n8312), .ZN(n8313) );
  OAI21_X1 U9542 ( .B1(n8315), .B2(n8314), .A(n8313), .ZN(n8316) );
  AOI211_X1 U9543 ( .C1(n10757), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n8317), .B(
        n8316), .ZN(n8318) );
  NAND2_X1 U9544 ( .A1(n8319), .A2(n8318), .ZN(P2_U3191) );
  XNOR2_X1 U9545 ( .A(n8320), .B(n5110), .ZN(n8322) );
  OAI222_X1 U9546 ( .A1(n9685), .A2(n9100), .B1(n9684), .B2(n8415), .C1(n9682), 
        .C2(n8322), .ZN(n8403) );
  INV_X1 U9547 ( .A(n8403), .ZN(n8329) );
  INV_X1 U9548 ( .A(n8421), .ZN(n8323) );
  OAI22_X1 U9549 ( .A1(n9672), .A2(n8324), .B1(n8323), .B2(n9669), .ZN(n8325)
         );
  AOI21_X1 U9550 ( .B1(n8426), .B2(n8536), .A(n8325), .ZN(n8328) );
  XNOR2_X1 U9551 ( .A(n8326), .B(n5110), .ZN(n8404) );
  NAND2_X1 U9552 ( .A1(n8404), .A2(n9692), .ZN(n8327) );
  OAI211_X1 U9553 ( .C1(n8329), .C2(n9694), .A(n8328), .B(n8327), .ZN(P2_U3224) );
  INV_X1 U9554 ( .A(n8330), .ZN(n8337) );
  AOI22_X1 U9555 ( .A1(n10297), .A2(n6945), .B1(n10159), .B2(n10044), .ZN(
        n8332) );
  AOI22_X1 U9556 ( .A1(n10335), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10274), .ZN(n8331) );
  OAI211_X1 U9557 ( .C1(n10264), .C2(n8333), .A(n8332), .B(n8331), .ZN(n8334)
         );
  AOI21_X1 U9558 ( .B1(n10321), .B2(n8335), .A(n8334), .ZN(n8336) );
  OAI21_X1 U9559 ( .B1(n10335), .B2(n8337), .A(n8336), .ZN(P1_U3291) );
  INV_X1 U9560 ( .A(n8338), .ZN(n8345) );
  AOI22_X1 U9561 ( .A1(n10297), .A2(n6967), .B1(n10159), .B2(n6960), .ZN(n8340) );
  AOI22_X1 U9562 ( .A1(n10335), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n10274), .ZN(n8339) );
  OAI211_X1 U9563 ( .C1(n10264), .C2(n8341), .A(n8340), .B(n8339), .ZN(n8342)
         );
  AOI21_X1 U9564 ( .B1(n10321), .B2(n8343), .A(n8342), .ZN(n8344) );
  OAI21_X1 U9565 ( .B1(n10335), .B2(n8345), .A(n8344), .ZN(P1_U3292) );
  INV_X1 U9566 ( .A(n8346), .ZN(n8355) );
  AOI22_X1 U9567 ( .A1(n10297), .A2(n8347), .B1(n10159), .B2(n10043), .ZN(
        n8350) );
  AOI22_X1 U9568 ( .A1(n10335), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10274), .B2(
        n8348), .ZN(n8349) );
  OAI211_X1 U9569 ( .C1(n10264), .C2(n8351), .A(n8350), .B(n8349), .ZN(n8352)
         );
  AOI21_X1 U9570 ( .B1(n8353), .B2(n10321), .A(n8352), .ZN(n8354) );
  OAI21_X1 U9571 ( .B1(n8355), .B2(n10335), .A(n8354), .ZN(P1_U3290) );
  INV_X1 U9572 ( .A(n8359), .ZN(n8356) );
  NOR2_X1 U9573 ( .A1(n8357), .A2(n8356), .ZN(n8362) );
  AOI21_X1 U9574 ( .B1(n8360), .B2(n8359), .A(n8358), .ZN(n8361) );
  OAI21_X1 U9575 ( .B1(n8362), .B2(n8361), .A(n10002), .ZN(n8367) );
  AOI22_X1 U9576 ( .A1(n10003), .A2(n10038), .B1(P1_REG3_REG_8__SCAN_IN), .B2(
        P1_U3086), .ZN(n8363) );
  OAI21_X1 U9577 ( .B1(n8494), .B2(n9991), .A(n8363), .ZN(n8364) );
  AOI21_X1 U9578 ( .B1(n8365), .B2(n10015), .A(n8364), .ZN(n8366) );
  OAI211_X1 U9579 ( .C1(n10802), .C2(n10009), .A(n8367), .B(n8366), .ZN(
        P1_U3221) );
  AOI22_X1 U9580 ( .A1(n10335), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n8368), .B2(
        n10274), .ZN(n8369) );
  OAI21_X1 U9581 ( .B1(n8370), .B2(n10325), .A(n8369), .ZN(n8373) );
  NOR2_X1 U9582 ( .A1(n8371), .A2(n8639), .ZN(n8372) );
  AOI211_X1 U9583 ( .C1(n8374), .C2(n10178), .A(n8373), .B(n8372), .ZN(n8375)
         );
  OAI21_X1 U9584 ( .B1(n10335), .B2(n8376), .A(n8375), .ZN(P1_U3286) );
  INV_X1 U9585 ( .A(n8377), .ZN(n8379) );
  NAND2_X1 U9586 ( .A1(n8379), .A2(n8378), .ZN(n8380) );
  XNOR2_X1 U9587 ( .A(n8381), .B(n8380), .ZN(n8390) );
  NAND2_X1 U9588 ( .A1(n10017), .A2(n10037), .ZN(n8384) );
  INV_X1 U9589 ( .A(n8382), .ZN(n8383) );
  OAI211_X1 U9590 ( .C1(n10020), .C2(n8385), .A(n8384), .B(n8383), .ZN(n8387)
         );
  NOR2_X1 U9591 ( .A1(n10009), .A2(n10814), .ZN(n8386) );
  AOI211_X1 U9592 ( .C1(n8388), .C2(n10015), .A(n8387), .B(n8386), .ZN(n8389)
         );
  OAI21_X1 U9593 ( .B1(n8390), .B2(n10026), .A(n8389), .ZN(P1_U3231) );
  NAND2_X1 U9594 ( .A1(n8260), .A2(n8391), .ZN(n8392) );
  XOR2_X1 U9595 ( .A(n8394), .B(n8392), .Z(n8393) );
  AOI22_X1 U9596 ( .A1(n8393), .A2(n10312), .B1(n10282), .B2(n10035), .ZN(
        n8430) );
  XNOR2_X1 U9597 ( .A(n8395), .B(n8394), .ZN(n8433) );
  NAND2_X1 U9598 ( .A1(n8433), .A2(n10321), .ZN(n8402) );
  INV_X1 U9599 ( .A(n10159), .ZN(n10278) );
  AOI22_X1 U9600 ( .A1(n10335), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n8567), .B2(
        n10274), .ZN(n8396) );
  OAI21_X1 U9601 ( .B1(n10278), .B2(n8431), .A(n8396), .ZN(n8400) );
  INV_X1 U9602 ( .A(n8474), .ZN(n8397) );
  OAI211_X1 U9603 ( .C1(n8437), .C2(n8398), .A(n8397), .B(n10292), .ZN(n8429)
         );
  NOR2_X1 U9604 ( .A1(n8429), .A2(n10264), .ZN(n8399) );
  AOI211_X1 U9605 ( .C1(n10297), .C2(n8572), .A(n8400), .B(n8399), .ZN(n8401)
         );
  OAI211_X1 U9606 ( .C1(n10335), .C2(n8430), .A(n8402), .B(n8401), .ZN(
        P1_U3282) );
  AOI21_X1 U9607 ( .B1(n8404), .B2(n9778), .A(n8403), .ZN(n8413) );
  INV_X1 U9608 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n8405) );
  NOR2_X1 U9609 ( .A1(n9781), .A2(n8405), .ZN(n8406) );
  AOI21_X1 U9610 ( .B1(n8426), .B2(n8407), .A(n8406), .ZN(n8408) );
  OAI21_X1 U9611 ( .B1(n8413), .B2(n7250), .A(n8408), .ZN(P2_U3468) );
  INV_X1 U9612 ( .A(n9833), .ZN(n8411) );
  INV_X1 U9613 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n8409) );
  NOR2_X1 U9614 ( .A1(n10851), .A2(n8409), .ZN(n8410) );
  AOI21_X1 U9615 ( .B1(n8426), .B2(n8411), .A(n8410), .ZN(n8412) );
  OAI21_X1 U9616 ( .B1(n8413), .B2(n7244), .A(n8412), .ZN(P2_U3417) );
  NAND2_X1 U9617 ( .A1(n8414), .A2(n9387), .ZN(n8417) );
  INV_X1 U9618 ( .A(n8414), .ZN(n8416) );
  XNOR2_X1 U9619 ( .A(n8426), .B(n7270), .ZN(n8576) );
  XNOR2_X1 U9620 ( .A(n8576), .B(n8578), .ZN(n8419) );
  OAI211_X1 U9621 ( .C1(n8420), .C2(n8419), .A(n8575), .B(n9109), .ZN(n8428)
         );
  NAND2_X1 U9622 ( .A1(n9136), .A2(n8421), .ZN(n8424) );
  AOI21_X1 U9623 ( .B1(n9387), .B2(n9132), .A(n8422), .ZN(n8423) );
  OAI211_X1 U9624 ( .C1(n9100), .C2(n9134), .A(n8424), .B(n8423), .ZN(n8425)
         );
  AOI21_X1 U9625 ( .B1(n9079), .B2(n8426), .A(n8425), .ZN(n8427) );
  NAND2_X1 U9626 ( .A1(n8428), .A2(n8427), .ZN(P2_U3171) );
  OAI211_X1 U9627 ( .C1(n8431), .C2(n10395), .A(n8430), .B(n8429), .ZN(n8432)
         );
  AOI21_X1 U9628 ( .B1(n8433), .B2(n10838), .A(n8432), .ZN(n8440) );
  AOI22_X1 U9629 ( .A1(n8572), .A2(n8917), .B1(n10840), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n8434) );
  OAI21_X1 U9630 ( .B1(n8440), .B2(n10840), .A(n8434), .ZN(P1_U3533) );
  INV_X1 U9631 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n8436) );
  OAI22_X1 U9632 ( .A1(n8437), .A2(n10469), .B1(n10846), .B2(n8436), .ZN(n8438) );
  INV_X1 U9633 ( .A(n8438), .ZN(n8439) );
  OAI21_X1 U9634 ( .B1(n8440), .B2(n10843), .A(n8439), .ZN(P1_U3486) );
  NAND2_X1 U9635 ( .A1(n8442), .A2(n8441), .ZN(n8444) );
  NAND2_X1 U9636 ( .A1(n8444), .A2(n8443), .ZN(n8446) );
  XNOR2_X1 U9637 ( .A(n8555), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n8445) );
  NOR2_X1 U9638 ( .A1(n8445), .A2(n8446), .ZN(n8547) );
  AOI21_X1 U9639 ( .B1(n8446), .B2(n8445), .A(n8547), .ZN(n8459) );
  NOR2_X1 U9640 ( .A1(n8448), .A2(n8447), .ZN(n8450) );
  NOR2_X1 U9641 ( .A1(n8450), .A2(n8449), .ZN(n8453) );
  NAND2_X1 U9642 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n8555), .ZN(n8451) );
  OAI21_X1 U9643 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n8555), .A(n8451), .ZN(
        n8452) );
  NOR2_X1 U9644 ( .A1(n8453), .A2(n8452), .ZN(n8554) );
  AOI211_X1 U9645 ( .C1(n8453), .C2(n8452), .A(n8554), .B(n10122), .ZN(n8454)
         );
  INV_X1 U9646 ( .A(n8454), .ZN(n8458) );
  NOR2_X1 U9647 ( .A1(n8455), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9922) );
  NOR2_X1 U9648 ( .A1(n10117), .A2(n8549), .ZN(n8456) );
  AOI211_X1 U9649 ( .C1(n10560), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9922), .B(
        n8456), .ZN(n8457) );
  OAI211_X1 U9650 ( .C1(n8459), .C2(n10090), .A(n8458), .B(n8457), .ZN(
        P1_U3259) );
  XNOR2_X1 U9651 ( .A(n8583), .B(n9100), .ZN(n9340) );
  XOR2_X1 U9652 ( .A(n8460), .B(n9340), .Z(n8461) );
  OAI222_X1 U9653 ( .A1(n9685), .A2(n9094), .B1(n9684), .B2(n8577), .C1(n8461), 
        .C2(n9682), .ZN(n8542) );
  INV_X1 U9654 ( .A(n8542), .ZN(n8467) );
  INV_X1 U9655 ( .A(n9340), .ZN(n8463) );
  XNOR2_X1 U9656 ( .A(n8462), .B(n8463), .ZN(n8541) );
  INV_X1 U9657 ( .A(n8541), .ZN(n8544) );
  INV_X1 U9658 ( .A(n8583), .ZN(n8539) );
  AOI22_X1 U9659 ( .A1(n9694), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n9688), .B2(
        n8579), .ZN(n8464) );
  OAI21_X1 U9660 ( .B1(n8539), .B2(n9652), .A(n8464), .ZN(n8465) );
  AOI21_X1 U9661 ( .B1(n8544), .B2(n9692), .A(n8465), .ZN(n8466) );
  OAI21_X1 U9662 ( .B1(n8467), .B2(n9694), .A(n8466), .ZN(P2_U3223) );
  XNOR2_X1 U9663 ( .A(n8468), .B(n8473), .ZN(n8471) );
  OAI22_X1 U9664 ( .A1(n8469), .A2(n10395), .B1(n9904), .B2(n10315), .ZN(n8470) );
  AOI21_X1 U9665 ( .B1(n8471), .B2(n10312), .A(n8470), .ZN(n10834) );
  XNOR2_X1 U9666 ( .A(n8472), .B(n8473), .ZN(n10839) );
  NAND2_X1 U9667 ( .A1(n10839), .A2(n10321), .ZN(n8479) );
  OAI211_X1 U9668 ( .C1(n8474), .C2(n10836), .A(n10292), .B(n8515), .ZN(n10833) );
  INV_X1 U9669 ( .A(n10833), .ZN(n8477) );
  NAND2_X1 U9670 ( .A1(n10328), .A2(n10116), .ZN(n10293) );
  INV_X1 U9671 ( .A(n10293), .ZN(n10331) );
  AOI22_X1 U9672 ( .A1(n10335), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n9901), .B2(
        n10274), .ZN(n8475) );
  OAI21_X1 U9673 ( .B1(n10836), .B2(n10325), .A(n8475), .ZN(n8476) );
  AOI21_X1 U9674 ( .B1(n8477), .B2(n10331), .A(n8476), .ZN(n8478) );
  OAI211_X1 U9675 ( .C1(n10335), .C2(n10834), .A(n8479), .B(n8478), .ZN(
        P1_U3281) );
  XNOR2_X1 U9676 ( .A(n4957), .B(n9343), .ZN(n8480) );
  OAI222_X1 U9677 ( .A1(n9685), .A2(n9683), .B1(n9684), .B2(n9100), .C1(n8480), 
        .C2(n9682), .ZN(n9775) );
  INV_X1 U9678 ( .A(n9775), .ZN(n8487) );
  OAI21_X1 U9679 ( .B1(n8482), .B2(n9343), .A(n8481), .ZN(n9777) );
  NOR2_X1 U9680 ( .A1(n9774), .A2(n9652), .ZN(n8485) );
  INV_X1 U9681 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10650) );
  INV_X1 U9682 ( .A(n9103), .ZN(n8483) );
  OAI22_X1 U9683 ( .A1(n9672), .A2(n10650), .B1(n8483), .B2(n9669), .ZN(n8484)
         );
  AOI211_X1 U9684 ( .C1(n9777), .C2(n9692), .A(n8485), .B(n8484), .ZN(n8486)
         );
  OAI21_X1 U9685 ( .B1(n8487), .B2(n9694), .A(n8486), .ZN(P2_U3222) );
  XOR2_X1 U9686 ( .A(n8489), .B(n8488), .Z(n8490) );
  XNOR2_X1 U9687 ( .A(n8491), .B(n8490), .ZN(n8499) );
  NAND2_X1 U9688 ( .A1(n10017), .A2(n10036), .ZN(n8493) );
  OAI211_X1 U9689 ( .C1(n10020), .C2(n8494), .A(n8493), .B(n8492), .ZN(n8496)
         );
  NOR2_X1 U9690 ( .A1(n10821), .A2(n10009), .ZN(n8495) );
  AOI211_X1 U9691 ( .C1(n8497), .C2(n10015), .A(n8496), .B(n8495), .ZN(n8498)
         );
  OAI21_X1 U9692 ( .B1(n8499), .B2(n10026), .A(n8498), .ZN(P1_U3217) );
  INV_X1 U9693 ( .A(n8500), .ZN(n8504) );
  OAI222_X1 U9694 ( .A1(n10494), .A2(n8502), .B1(n10492), .B2(n8504), .C1(
        n8501), .C2(P1_U3086), .ZN(P1_U3333) );
  INV_X1 U9695 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8503) );
  OAI222_X1 U9696 ( .A1(n8505), .A2(P2_U3151), .B1(n9856), .B2(n8504), .C1(
        n8503), .C2(n9855), .ZN(P2_U3273) );
  XOR2_X1 U9697 ( .A(n8509), .B(n8506), .Z(n8602) );
  INV_X1 U9698 ( .A(n8602), .ZN(n8521) );
  OAI21_X1 U9699 ( .B1(n8509), .B2(n8508), .A(n8507), .ZN(n8510) );
  NAND2_X1 U9700 ( .A1(n8510), .A2(n10312), .ZN(n8513) );
  AOI22_X1 U9701 ( .A1(n8511), .A2(n10282), .B1(n10389), .B2(n10035), .ZN(
        n8512) );
  NAND2_X1 U9702 ( .A1(n8513), .A2(n8512), .ZN(n8600) );
  INV_X1 U9703 ( .A(n8635), .ZN(n8514) );
  AOI211_X1 U9704 ( .C1(n8516), .C2(n8515), .A(n10803), .B(n8514), .ZN(n8601)
         );
  NAND2_X1 U9705 ( .A1(n8601), .A2(n10286), .ZN(n8518) );
  AOI22_X1 U9706 ( .A1(n10335), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9972), .B2(
        n10274), .ZN(n8517) );
  OAI211_X1 U9707 ( .C1(n9975), .C2(n10325), .A(n8518), .B(n8517), .ZN(n8519)
         );
  AOI21_X1 U9708 ( .B1(n10328), .B2(n8600), .A(n8519), .ZN(n8520) );
  OAI21_X1 U9709 ( .B1(n8521), .B2(n10307), .A(n8520), .ZN(P1_U3280) );
  INV_X1 U9710 ( .A(n8524), .ZN(n8523) );
  AOI21_X1 U9711 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n9846), .A(n9365), .ZN(
        n8522) );
  OAI21_X1 U9712 ( .B1(n8523), .B2(n9856), .A(n8522), .ZN(P2_U3272) );
  NAND2_X1 U9713 ( .A1(n8524), .A2(n8886), .ZN(n8526) );
  OAI211_X1 U9714 ( .C1(n8527), .C2(n10494), .A(n8526), .B(n8525), .ZN(
        P1_U3332) );
  XNOR2_X1 U9715 ( .A(n8528), .B(n9209), .ZN(n9767) );
  OAI211_X1 U9716 ( .C1(n8529), .C2(n9209), .A(n8530), .B(n7237), .ZN(n8532)
         );
  AOI22_X1 U9717 ( .A1(n9385), .A2(n9540), .B1(n9541), .B2(n9383), .ZN(n8531)
         );
  NAND2_X1 U9718 ( .A1(n8532), .A2(n8531), .ZN(n9768) );
  NAND2_X1 U9719 ( .A1(n9768), .A2(n9672), .ZN(n8538) );
  INV_X1 U9720 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8534) );
  INV_X1 U9721 ( .A(n8596), .ZN(n8533) );
  OAI22_X1 U9722 ( .A1(n9672), .A2(n8534), .B1(n8533), .B2(n9669), .ZN(n8535)
         );
  AOI21_X1 U9723 ( .B1(n9770), .B2(n8536), .A(n8535), .ZN(n8537) );
  OAI211_X1 U9724 ( .C1(n9767), .C2(n9676), .A(n8538), .B(n8537), .ZN(P2_U3221) );
  INV_X1 U9725 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9395) );
  OAI22_X1 U9726 ( .A1(n8541), .A2(n8540), .B1(n8539), .B2(n9773), .ZN(n8543)
         );
  AOI211_X1 U9727 ( .C1(n8545), .C2(n8544), .A(n8543), .B(n8542), .ZN(n10828)
         );
  OR2_X1 U9728 ( .A1(n10828), .A2(n7250), .ZN(n8546) );
  OAI21_X1 U9729 ( .B1(n9781), .B2(n9395), .A(n8546), .ZN(P2_U3469) );
  INV_X1 U9730 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n8548) );
  AOI21_X1 U9731 ( .B1(n8549), .B2(n8548), .A(n8547), .ZN(n8551) );
  XNOR2_X1 U9732 ( .A(n10096), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n8550) );
  NOR2_X1 U9733 ( .A1(n8551), .A2(n8550), .ZN(n10088) );
  AOI21_X1 U9734 ( .B1(n8551), .B2(n8550), .A(n10088), .ZN(n8553) );
  NAND2_X1 U9735 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9933) );
  NAND2_X1 U9736 ( .A1(n10560), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n8552) );
  OAI211_X1 U9737 ( .C1(n8553), .C2(n10090), .A(n9933), .B(n8552), .ZN(n8560)
         );
  AOI21_X1 U9738 ( .B1(n8555), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8554), .ZN(
        n8558) );
  NOR2_X1 U9739 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n10096), .ZN(n8556) );
  AOI21_X1 U9740 ( .B1(n10096), .B2(P1_REG2_REG_17__SCAN_IN), .A(n8556), .ZN(
        n8557) );
  NAND2_X1 U9741 ( .A1(n8557), .A2(n8558), .ZN(n10095) );
  AOI221_X1 U9742 ( .B1(n8558), .B2(n10095), .C1(n8557), .C2(n10095), .A(
        n10122), .ZN(n8559) );
  AOI211_X1 U9743 ( .C1(n10076), .C2(n10096), .A(n8560), .B(n8559), .ZN(n8561)
         );
  INV_X1 U9744 ( .A(n8561), .ZN(P1_U3260) );
  NAND2_X1 U9745 ( .A1(n8563), .A2(n8562), .ZN(n8565) );
  XOR2_X1 U9746 ( .A(n8565), .B(n8564), .Z(n8574) );
  AOI21_X1 U9747 ( .B1(n10003), .B2(n10037), .A(n8566), .ZN(n8569) );
  NAND2_X1 U9748 ( .A1(n10015), .A2(n8567), .ZN(n8568) );
  OAI211_X1 U9749 ( .C1(n8570), .C2(n9991), .A(n8569), .B(n8568), .ZN(n8571)
         );
  AOI21_X1 U9750 ( .B1(n8572), .B2(n10023), .A(n8571), .ZN(n8573) );
  OAI21_X1 U9751 ( .B1(n8574), .B2(n10026), .A(n8573), .ZN(P1_U3236) );
  XNOR2_X1 U9752 ( .A(n8583), .B(n8966), .ZN(n9092) );
  XNOR2_X1 U9753 ( .A(n9091), .B(n9092), .ZN(n9093) );
  XNOR2_X1 U9754 ( .A(n9093), .B(n9100), .ZN(n8585) );
  AOI22_X1 U9755 ( .A1(n8578), .A2(n9132), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3151), .ZN(n8581) );
  NAND2_X1 U9756 ( .A1(n9136), .A2(n8579), .ZN(n8580) );
  OAI211_X1 U9757 ( .C1(n9094), .C2(n9134), .A(n8581), .B(n8580), .ZN(n8582)
         );
  AOI21_X1 U9758 ( .B1(n9079), .B2(n8583), .A(n8582), .ZN(n8584) );
  OAI21_X1 U9759 ( .B1(n8585), .B2(n9127), .A(n8584), .ZN(P2_U3157) );
  INV_X1 U9760 ( .A(n9770), .ZN(n8599) );
  XNOR2_X1 U9761 ( .A(n9774), .B(n7270), .ZN(n9095) );
  AOI22_X1 U9762 ( .A1(n9095), .A2(n9385), .B1(n9092), .B2(n9386), .ZN(n8590)
         );
  INV_X1 U9763 ( .A(n9092), .ZN(n8586) );
  AOI21_X1 U9764 ( .B1(n8586), .B2(n9100), .A(n9094), .ZN(n8588) );
  NAND3_X1 U9765 ( .A1(n8586), .A2(n9100), .A3(n9094), .ZN(n8587) );
  OAI21_X1 U9766 ( .B1(n9095), .B2(n8588), .A(n8587), .ZN(n8589) );
  XNOR2_X1 U9767 ( .A(n9770), .B(n7270), .ZN(n8936) );
  XNOR2_X1 U9768 ( .A(n8936), .B(n9384), .ZN(n8591) );
  OAI211_X1 U9769 ( .C1(n8592), .C2(n8591), .A(n8938), .B(n9109), .ZN(n8598)
         );
  NAND2_X1 U9770 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n10670) );
  INV_X1 U9771 ( .A(n10670), .ZN(n8593) );
  AOI21_X1 U9772 ( .B1(n9385), .B2(n9132), .A(n8593), .ZN(n8594) );
  OAI21_X1 U9773 ( .B1(n9666), .B2(n9134), .A(n8594), .ZN(n8595) );
  AOI21_X1 U9774 ( .B1(n8596), .B2(n9136), .A(n8595), .ZN(n8597) );
  OAI211_X1 U9775 ( .C1(n8599), .C2(n9139), .A(n8598), .B(n8597), .ZN(P2_U3164) );
  INV_X1 U9776 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n8603) );
  AOI211_X1 U9777 ( .C1(n8602), .C2(n10838), .A(n8601), .B(n8600), .ZN(n8605)
         );
  MUX2_X1 U9778 ( .A(n8603), .B(n8605), .S(n10846), .Z(n8604) );
  OAI21_X1 U9779 ( .B1(n9975), .B2(n10469), .A(n8604), .ZN(P1_U3492) );
  MUX2_X1 U9780 ( .A(n8606), .B(n8605), .S(n10842), .Z(n8607) );
  OAI21_X1 U9781 ( .B1(n9975), .B2(n10419), .A(n8607), .ZN(P1_U3535) );
  INV_X1 U9782 ( .A(n8608), .ZN(n8611) );
  INV_X1 U9783 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8609) );
  OAI222_X1 U9784 ( .A1(n8610), .A2(P2_U3151), .B1(n9856), .B2(n8611), .C1(
        n8609), .C2(n9855), .ZN(P2_U3271) );
  INV_X1 U9785 ( .A(n6170), .ZN(n8612) );
  OAI222_X1 U9786 ( .A1(n10494), .A2(n8613), .B1(P1_U3086), .B2(n8612), .C1(
        n8611), .C2(n10492), .ZN(P1_U3331) );
  XOR2_X1 U9787 ( .A(n8617), .B(n8614), .Z(n8615) );
  AOI22_X1 U9788 ( .A1(n8615), .A2(n10312), .B1(n10282), .B2(n10032), .ZN(
        n8891) );
  XNOR2_X1 U9789 ( .A(n8616), .B(n8617), .ZN(n8893) );
  NAND2_X1 U9790 ( .A1(n8893), .A2(n10321), .ZN(n8622) );
  AOI22_X1 U9791 ( .A1(n10335), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n10014), 
        .B2(n10274), .ZN(n8618) );
  OAI21_X1 U9792 ( .B1(n10278), .B2(n10021), .A(n8618), .ZN(n8620) );
  OAI211_X1 U9793 ( .C1(n8634), .C2(n8899), .A(n8650), .B(n10292), .ZN(n8890)
         );
  NOR2_X1 U9794 ( .A1(n8890), .A2(n10264), .ZN(n8619) );
  AOI211_X1 U9795 ( .C1(n10297), .C2(n10024), .A(n8620), .B(n8619), .ZN(n8621)
         );
  OAI211_X1 U9796 ( .C1(n10335), .C2(n8891), .A(n8622), .B(n8621), .ZN(
        P1_U3278) );
  INV_X1 U9797 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8623) );
  OAI222_X1 U9798 ( .A1(n8624), .A2(P2_U3151), .B1(n9856), .B2(n6512), .C1(
        n8623), .C2(n9855), .ZN(P2_U3270) );
  OAI222_X1 U9799 ( .A1(n8626), .A2(P1_U3086), .B1(n10492), .B2(n6512), .C1(
        n8625), .C2(n10494), .ZN(P1_U3330) );
  XNOR2_X1 U9800 ( .A(n8627), .B(n5263), .ZN(n8638) );
  XNOR2_X1 U9801 ( .A(n8629), .B(n8628), .ZN(n8631) );
  AOI22_X1 U9802 ( .A1(n10034), .A2(n10389), .B1(n10282), .B2(n10033), .ZN(
        n8630) );
  OAI21_X1 U9803 ( .B1(n8631), .B2(n8902), .A(n8630), .ZN(n8632) );
  AOI21_X1 U9804 ( .B1(n8638), .B2(n8633), .A(n8632), .ZN(n10430) );
  AOI211_X1 U9805 ( .C1(n10427), .C2(n8635), .A(n10803), .B(n8634), .ZN(n10426) );
  INV_X1 U9806 ( .A(n10427), .ZN(n8637) );
  AOI22_X1 U9807 ( .A1(n10335), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9863), .B2(
        n10274), .ZN(n8636) );
  OAI21_X1 U9808 ( .B1(n8637), .B2(n10325), .A(n8636), .ZN(n8641) );
  INV_X1 U9809 ( .A(n8638), .ZN(n10431) );
  NOR2_X1 U9810 ( .A1(n10431), .A2(n8639), .ZN(n8640) );
  AOI211_X1 U9811 ( .C1(n10426), .C2(n10286), .A(n8641), .B(n8640), .ZN(n8642)
         );
  OAI21_X1 U9812 ( .B1(n10335), .B2(n10430), .A(n8642), .ZN(P1_U3279) );
  OAI21_X1 U9813 ( .B1(n8644), .B2(n8648), .A(n8643), .ZN(n10424) );
  INV_X1 U9814 ( .A(n8645), .ZN(n8646) );
  AOI21_X1 U9815 ( .B1(n8648), .B2(n8647), .A(n8646), .ZN(n8649) );
  OAI222_X1 U9816 ( .A1(n10315), .A2(n10314), .B1(n10395), .B2(n9925), .C1(
        n8902), .C2(n8649), .ZN(n10420) );
  AOI211_X1 U9817 ( .C1(n10422), .C2(n8650), .A(n10803), .B(n8906), .ZN(n10421) );
  NAND2_X1 U9818 ( .A1(n10421), .A2(n10286), .ZN(n8652) );
  AOI22_X1 U9819 ( .A1(n10335), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9921), .B2(
        n10274), .ZN(n8651) );
  OAI211_X1 U9820 ( .C1(n8653), .C2(n10325), .A(n8652), .B(n8651), .ZN(n8654)
         );
  AOI21_X1 U9821 ( .B1(n10420), .B2(n10328), .A(n8654), .ZN(n8655) );
  OAI21_X1 U9822 ( .B1(n10424), .B2(n10307), .A(n8655), .ZN(P1_U3277) );
  XOR2_X1 U9823 ( .A(n8876), .B(keyinput_62), .Z(n8884) );
  INV_X1 U9824 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9099) );
  INV_X1 U9825 ( .A(keyinput_58), .ZN(n8743) );
  INV_X1 U9826 ( .A(keyinput_57), .ZN(n8741) );
  INV_X1 U9827 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9076) );
  INV_X1 U9828 ( .A(keyinput_56), .ZN(n8739) );
  AOI22_X1 U9829 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_49), .B1(n6437), 
        .B2(keyinput_50), .ZN(n8656) );
  OAI221_X1 U9830 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_49), .C1(n6437), 
        .C2(keyinput_50), .A(n8656), .ZN(n8730) );
  INV_X1 U9831 ( .A(keyinput_48), .ZN(n8728) );
  INV_X1 U9832 ( .A(keyinput_47), .ZN(n8726) );
  INV_X1 U9833 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8848) );
  INV_X1 U9834 ( .A(keyinput_46), .ZN(n8724) );
  INV_X1 U9835 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8842) );
  INV_X1 U9836 ( .A(keyinput_45), .ZN(n8722) );
  INV_X1 U9837 ( .A(keyinput_44), .ZN(n8720) );
  INV_X1 U9838 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n8839) );
  INV_X1 U9839 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8837) );
  OAI22_X1 U9840 ( .A1(n8837), .A2(keyinput_42), .B1(keyinput_41), .B2(
        P2_REG3_REG_19__SCAN_IN), .ZN(n8657) );
  AOI221_X1 U9841 ( .B1(n8837), .B2(keyinput_42), .C1(P2_REG3_REG_19__SCAN_IN), 
        .C2(keyinput_41), .A(n8657), .ZN(n8717) );
  INV_X1 U9842 ( .A(keyinput_40), .ZN(n8715) );
  INV_X1 U9843 ( .A(keyinput_39), .ZN(n8713) );
  INV_X1 U9844 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8830) );
  INV_X1 U9845 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8826) );
  INV_X1 U9846 ( .A(keyinput_38), .ZN(n8711) );
  INV_X1 U9847 ( .A(keyinput_37), .ZN(n8709) );
  OAI22_X1 U9848 ( .A1(P2_U3151), .A2(keyinput_34), .B1(keyinput_35), .B2(
        P2_REG3_REG_7__SCAN_IN), .ZN(n8658) );
  AOI221_X1 U9849 ( .B1(P2_U3151), .B2(keyinput_34), .C1(
        P2_REG3_REG_7__SCAN_IN), .C2(keyinput_35), .A(n8658), .ZN(n8706) );
  INV_X1 U9850 ( .A(SI_11_), .ZN(n8755) );
  OAI22_X1 U9851 ( .A1(n8755), .A2(keyinput_21), .B1(SI_10_), .B2(keyinput_22), 
        .ZN(n8659) );
  AOI221_X1 U9852 ( .B1(n8755), .B2(keyinput_21), .C1(keyinput_22), .C2(SI_10_), .A(n8659), .ZN(n8692) );
  INV_X1 U9853 ( .A(SI_15_), .ZN(n8791) );
  INV_X1 U9854 ( .A(keyinput_17), .ZN(n8682) );
  INV_X1 U9855 ( .A(keyinput_16), .ZN(n8680) );
  INV_X1 U9856 ( .A(keyinput_15), .ZN(n8678) );
  AOI22_X1 U9857 ( .A1(SI_25_), .A2(keyinput_7), .B1(SI_26_), .B2(keyinput_6), 
        .ZN(n8660) );
  OAI221_X1 U9858 ( .B1(SI_25_), .B2(keyinput_7), .C1(SI_26_), .C2(keyinput_6), 
        .A(n8660), .ZN(n8668) );
  AOI22_X1 U9859 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_0), .B1(SI_30_), .B2(
        keyinput_2), .ZN(n8661) );
  OAI221_X1 U9860 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_0), .C1(SI_30_), .C2(
        keyinput_2), .A(n8661), .ZN(n8666) );
  AOI22_X1 U9861 ( .A1(SI_28_), .A2(keyinput_4), .B1(SI_27_), .B2(keyinput_5), 
        .ZN(n8662) );
  OAI221_X1 U9862 ( .B1(SI_28_), .B2(keyinput_4), .C1(SI_27_), .C2(keyinput_5), 
        .A(n8662), .ZN(n8665) );
  AOI22_X1 U9863 ( .A1(SI_31_), .A2(keyinput_1), .B1(SI_29_), .B2(keyinput_3), 
        .ZN(n8663) );
  OAI221_X1 U9864 ( .B1(SI_31_), .B2(keyinput_1), .C1(SI_29_), .C2(keyinput_3), 
        .A(n8663), .ZN(n8664) );
  NOR3_X1 U9865 ( .A1(n8666), .A2(n8665), .A3(n8664), .ZN(n8667) );
  OAI22_X1 U9866 ( .A1(n8668), .A2(n8667), .B1(SI_22_), .B2(keyinput_10), .ZN(
        n8669) );
  AOI21_X1 U9867 ( .B1(SI_22_), .B2(keyinput_10), .A(n8669), .ZN(n8676) );
  OAI22_X1 U9868 ( .A1(SI_24_), .A2(keyinput_8), .B1(keyinput_9), .B2(SI_23_), 
        .ZN(n8670) );
  AOI221_X1 U9869 ( .B1(SI_24_), .B2(keyinput_8), .C1(SI_23_), .C2(keyinput_9), 
        .A(n8670), .ZN(n8675) );
  AOI22_X1 U9870 ( .A1(n8775), .A2(keyinput_13), .B1(n8778), .B2(keyinput_12), 
        .ZN(n8671) );
  OAI221_X1 U9871 ( .B1(n8775), .B2(keyinput_13), .C1(n8778), .C2(keyinput_12), 
        .A(n8671), .ZN(n8674) );
  AOI22_X1 U9872 ( .A1(SI_18_), .A2(keyinput_14), .B1(SI_21_), .B2(keyinput_11), .ZN(n8672) );
  OAI221_X1 U9873 ( .B1(SI_18_), .B2(keyinput_14), .C1(SI_21_), .C2(
        keyinput_11), .A(n8672), .ZN(n8673) );
  AOI211_X1 U9874 ( .C1(n8676), .C2(n8675), .A(n8674), .B(n8673), .ZN(n8677)
         );
  AOI221_X1 U9875 ( .B1(SI_17_), .B2(keyinput_15), .C1(n8784), .C2(n8678), .A(
        n8677), .ZN(n8679) );
  AOI221_X1 U9876 ( .B1(SI_16_), .B2(keyinput_16), .C1(n8788), .C2(n8680), .A(
        n8679), .ZN(n8681) );
  AOI221_X1 U9877 ( .B1(SI_15_), .B2(keyinput_17), .C1(n8791), .C2(n8682), .A(
        n8681), .ZN(n8686) );
  INV_X1 U9878 ( .A(SI_13_), .ZN(n8793) );
  INV_X1 U9879 ( .A(SI_12_), .ZN(n8684) );
  AOI22_X1 U9880 ( .A1(n8793), .A2(keyinput_19), .B1(keyinput_20), .B2(n8684), 
        .ZN(n8683) );
  OAI221_X1 U9881 ( .B1(n8793), .B2(keyinput_19), .C1(n8684), .C2(keyinput_20), 
        .A(n8683), .ZN(n8685) );
  AOI211_X1 U9882 ( .C1(SI_14_), .C2(keyinput_18), .A(n8686), .B(n8685), .ZN(
        n8687) );
  OAI21_X1 U9883 ( .B1(SI_14_), .B2(keyinput_18), .A(n8687), .ZN(n8691) );
  AOI22_X1 U9884 ( .A1(SI_9_), .A2(keyinput_23), .B1(n8689), .B2(keyinput_24), 
        .ZN(n8688) );
  OAI221_X1 U9885 ( .B1(SI_9_), .B2(keyinput_23), .C1(n8689), .C2(keyinput_24), 
        .A(n8688), .ZN(n8690) );
  AOI21_X1 U9886 ( .B1(n8692), .B2(n8691), .A(n8690), .ZN(n8699) );
  AOI22_X1 U9887 ( .A1(n8810), .A2(keyinput_29), .B1(n8805), .B2(keyinput_28), 
        .ZN(n8693) );
  OAI221_X1 U9888 ( .B1(n8810), .B2(keyinput_29), .C1(n8805), .C2(keyinput_28), 
        .A(n8693), .ZN(n8696) );
  AOI22_X1 U9889 ( .A1(n8803), .A2(keyinput_25), .B1(keyinput_27), .B2(n8802), 
        .ZN(n8694) );
  OAI221_X1 U9890 ( .B1(n8803), .B2(keyinput_25), .C1(n8802), .C2(keyinput_27), 
        .A(n8694), .ZN(n8695) );
  AOI211_X1 U9891 ( .C1(keyinput_26), .C2(SI_6_), .A(n8696), .B(n8695), .ZN(
        n8697) );
  OAI21_X1 U9892 ( .B1(keyinput_26), .B2(SI_6_), .A(n8697), .ZN(n8698) );
  OR2_X1 U9893 ( .A1(n8699), .A2(n8698), .ZN(n8704) );
  OAI22_X1 U9894 ( .A1(SI_1_), .A2(keyinput_31), .B1(SI_0_), .B2(keyinput_32), 
        .ZN(n8700) );
  AOI221_X1 U9895 ( .B1(SI_1_), .B2(keyinput_31), .C1(keyinput_32), .C2(SI_0_), 
        .A(n8700), .ZN(n8703) );
  INV_X1 U9896 ( .A(P2_RD_REG_SCAN_IN), .ZN(n10776) );
  XNOR2_X1 U9897 ( .A(keyinput_33), .B(P2_RD_REG_SCAN_IN), .ZN(n8702) );
  XNOR2_X1 U9898 ( .A(SI_2_), .B(keyinput_30), .ZN(n8701) );
  NAND4_X1 U9899 ( .A1(n8704), .A2(n8703), .A3(n8702), .A4(n8701), .ZN(n8705)
         );
  AOI22_X1 U9900 ( .A1(n8706), .A2(n8705), .B1(keyinput_36), .B2(
        P2_REG3_REG_27__SCAN_IN), .ZN(n8707) );
  OAI21_X1 U9901 ( .B1(keyinput_36), .B2(P2_REG3_REG_27__SCAN_IN), .A(n8707), 
        .ZN(n8708) );
  OAI221_X1 U9902 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(n8709), .C1(n8823), .C2(
        keyinput_37), .A(n8708), .ZN(n8710) );
  OAI221_X1 U9903 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_38), .C1(n8826), 
        .C2(n8711), .A(n8710), .ZN(n8712) );
  OAI221_X1 U9904 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(n8713), .C1(n8830), .C2(
        keyinput_39), .A(n8712), .ZN(n8714) );
  OAI221_X1 U9905 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n8715), .C1(n8833), .C2(
        keyinput_40), .A(n8714), .ZN(n8716) );
  OAI211_X1 U9906 ( .C1(n8750), .C2(keyinput_43), .A(n8717), .B(n8716), .ZN(
        n8718) );
  AOI21_X1 U9907 ( .B1(n8750), .B2(keyinput_43), .A(n8718), .ZN(n8719) );
  AOI221_X1 U9908 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n8720), .C1(n8839), .C2(
        keyinput_44), .A(n8719), .ZN(n8721) );
  AOI221_X1 U9909 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_45), .C1(n8842), 
        .C2(n8722), .A(n8721), .ZN(n8723) );
  AOI221_X1 U9910 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(n8724), .C1(n8846), .C2(
        keyinput_46), .A(n8723), .ZN(n8725) );
  AOI221_X1 U9911 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(n8726), .C1(n8848), .C2(
        keyinput_47), .A(n8725), .ZN(n8727) );
  AOI221_X1 U9912 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_48), .C1(n8851), 
        .C2(n8728), .A(n8727), .ZN(n8729) );
  OAI22_X1 U9913 ( .A1(keyinput_51), .A2(n8732), .B1(n8730), .B2(n8729), .ZN(
        n8731) );
  AOI21_X1 U9914 ( .B1(keyinput_51), .B2(n8732), .A(n8731), .ZN(n8737) );
  AOI22_X1 U9915 ( .A1(n6345), .A2(keyinput_53), .B1(n8857), .B2(keyinput_55), 
        .ZN(n8733) );
  OAI221_X1 U9916 ( .B1(n6345), .B2(keyinput_53), .C1(n8857), .C2(keyinput_55), 
        .A(n8733), .ZN(n8736) );
  AOI22_X1 U9917 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_54), .B1(
        P2_REG3_REG_4__SCAN_IN), .B2(keyinput_52), .ZN(n8734) );
  OAI221_X1 U9918 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_54), .C1(
        P2_REG3_REG_4__SCAN_IN), .C2(keyinput_52), .A(n8734), .ZN(n8735) );
  NOR3_X1 U9919 ( .A1(n8737), .A2(n8736), .A3(n8735), .ZN(n8738) );
  AOI221_X1 U9920 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_56), .C1(n9076), 
        .C2(n8739), .A(n8738), .ZN(n8740) );
  AOI221_X1 U9921 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_57), .C1(n8866), 
        .C2(n8741), .A(n8740), .ZN(n8742) );
  AOI221_X1 U9922 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_58), .C1(n9099), 
        .C2(n8743), .A(n8742), .ZN(n8747) );
  AOI22_X1 U9923 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_59), .B1(n8745), 
        .B2(keyinput_60), .ZN(n8744) );
  OAI221_X1 U9924 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_59), .C1(n8745), 
        .C2(keyinput_60), .A(n8744), .ZN(n8746) );
  AOI211_X1 U9925 ( .C1(P2_REG3_REG_6__SCAN_IN), .C2(keyinput_61), .A(n8747), 
        .B(n8746), .ZN(n8748) );
  OAI21_X1 U9926 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_61), .A(n8748), 
        .ZN(n8883) );
  INV_X1 U9927 ( .A(keyinput_126), .ZN(n8877) );
  INV_X1 U9928 ( .A(keyinput_122), .ZN(n8869) );
  INV_X1 U9929 ( .A(keyinput_121), .ZN(n8867) );
  INV_X1 U9930 ( .A(keyinput_112), .ZN(n8852) );
  INV_X1 U9931 ( .A(keyinput_111), .ZN(n8849) );
  INV_X1 U9932 ( .A(keyinput_110), .ZN(n8845) );
  INV_X1 U9933 ( .A(keyinput_109), .ZN(n8843) );
  INV_X1 U9934 ( .A(keyinput_108), .ZN(n8840) );
  INV_X1 U9935 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9018) );
  OAI22_X1 U9936 ( .A1(n9018), .A2(keyinput_105), .B1(n8750), .B2(keyinput_107), .ZN(n8749) );
  AOI221_X1 U9937 ( .B1(n9018), .B2(keyinput_105), .C1(keyinput_107), .C2(
        n8750), .A(n8749), .ZN(n8835) );
  INV_X1 U9938 ( .A(keyinput_104), .ZN(n8832) );
  INV_X1 U9939 ( .A(keyinput_103), .ZN(n8829) );
  INV_X1 U9940 ( .A(keyinput_102), .ZN(n8827) );
  INV_X1 U9941 ( .A(keyinput_101), .ZN(n8824) );
  INV_X1 U9942 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8821) );
  OAI22_X1 U9943 ( .A1(n8752), .A2(keyinput_99), .B1(keyinput_98), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n8751) );
  AOI221_X1 U9944 ( .B1(n8752), .B2(keyinput_99), .C1(P2_STATE_REG_SCAN_IN), 
        .C2(keyinput_98), .A(n8751), .ZN(n8819) );
  OAI22_X1 U9945 ( .A1(n8755), .A2(keyinput_85), .B1(n8754), .B2(keyinput_86), 
        .ZN(n8753) );
  AOI221_X1 U9946 ( .B1(n8755), .B2(keyinput_85), .C1(keyinput_86), .C2(n8754), 
        .A(n8753), .ZN(n8800) );
  INV_X1 U9947 ( .A(keyinput_81), .ZN(n8790) );
  INV_X1 U9948 ( .A(keyinput_80), .ZN(n8787) );
  INV_X1 U9949 ( .A(keyinput_79), .ZN(n8785) );
  INV_X1 U9950 ( .A(SI_25_), .ZN(n8758) );
  AOI22_X1 U9951 ( .A1(n8758), .A2(keyinput_71), .B1(n8757), .B2(keyinput_70), 
        .ZN(n8756) );
  OAI221_X1 U9952 ( .B1(n8758), .B2(keyinput_71), .C1(n8757), .C2(keyinput_70), 
        .A(n8756), .ZN(n8769) );
  AOI22_X1 U9953 ( .A1(SI_31_), .A2(keyinput_65), .B1(SI_28_), .B2(keyinput_68), .ZN(n8759) );
  OAI221_X1 U9954 ( .B1(SI_31_), .B2(keyinput_65), .C1(SI_28_), .C2(
        keyinput_68), .A(n8759), .ZN(n8767) );
  AOI22_X1 U9955 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_64), .B1(n8761), .B2(
        keyinput_69), .ZN(n8760) );
  OAI221_X1 U9956 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_64), .C1(n8761), .C2(
        keyinput_69), .A(n8760), .ZN(n8766) );
  AOI22_X1 U9957 ( .A1(n8764), .A2(keyinput_66), .B1(n8763), .B2(keyinput_67), 
        .ZN(n8762) );
  OAI221_X1 U9958 ( .B1(n8764), .B2(keyinput_66), .C1(n8763), .C2(keyinput_67), 
        .A(n8762), .ZN(n8765) );
  NOR3_X1 U9959 ( .A1(n8767), .A2(n8766), .A3(n8765), .ZN(n8768) );
  OAI22_X1 U9960 ( .A1(n8769), .A2(n8768), .B1(n8771), .B2(keyinput_73), .ZN(
        n8770) );
  AOI21_X1 U9961 ( .B1(n8771), .B2(keyinput_73), .A(n8770), .ZN(n8782) );
  OAI22_X1 U9962 ( .A1(SI_24_), .A2(keyinput_72), .B1(keyinput_74), .B2(SI_22_), .ZN(n8772) );
  AOI221_X1 U9963 ( .B1(SI_24_), .B2(keyinput_72), .C1(SI_22_), .C2(
        keyinput_74), .A(n8772), .ZN(n8781) );
  AOI22_X1 U9964 ( .A1(n8775), .A2(keyinput_77), .B1(n8774), .B2(keyinput_75), 
        .ZN(n8773) );
  OAI221_X1 U9965 ( .B1(n8775), .B2(keyinput_77), .C1(n8774), .C2(keyinput_75), 
        .A(n8773), .ZN(n8780) );
  AOI22_X1 U9966 ( .A1(n8778), .A2(keyinput_76), .B1(keyinput_78), .B2(n8777), 
        .ZN(n8776) );
  OAI221_X1 U9967 ( .B1(n8778), .B2(keyinput_76), .C1(n8777), .C2(keyinput_78), 
        .A(n8776), .ZN(n8779) );
  AOI211_X1 U9968 ( .C1(n8782), .C2(n8781), .A(n8780), .B(n8779), .ZN(n8783)
         );
  AOI221_X1 U9969 ( .B1(SI_17_), .B2(n8785), .C1(n8784), .C2(keyinput_79), .A(
        n8783), .ZN(n8786) );
  AOI221_X1 U9970 ( .B1(SI_16_), .B2(keyinput_80), .C1(n8788), .C2(n8787), .A(
        n8786), .ZN(n8789) );
  AOI221_X1 U9971 ( .B1(SI_15_), .B2(keyinput_81), .C1(n8791), .C2(n8790), .A(
        n8789), .ZN(n8795) );
  AOI22_X1 U9972 ( .A1(SI_12_), .A2(keyinput_84), .B1(n8793), .B2(keyinput_83), 
        .ZN(n8792) );
  OAI221_X1 U9973 ( .B1(SI_12_), .B2(keyinput_84), .C1(n8793), .C2(keyinput_83), .A(n8792), .ZN(n8794) );
  AOI211_X1 U9974 ( .C1(SI_14_), .C2(keyinput_82), .A(n8795), .B(n8794), .ZN(
        n8796) );
  OAI21_X1 U9975 ( .B1(SI_14_), .B2(keyinput_82), .A(n8796), .ZN(n8799) );
  AOI22_X1 U9976 ( .A1(SI_8_), .A2(keyinput_88), .B1(SI_9_), .B2(keyinput_87), 
        .ZN(n8797) );
  OAI221_X1 U9977 ( .B1(SI_8_), .B2(keyinput_88), .C1(SI_9_), .C2(keyinput_87), 
        .A(n8797), .ZN(n8798) );
  AOI21_X1 U9978 ( .B1(n8800), .B2(n8799), .A(n8798), .ZN(n8812) );
  OAI22_X1 U9979 ( .A1(n8803), .A2(keyinput_89), .B1(n8802), .B2(keyinput_91), 
        .ZN(n8801) );
  AOI221_X1 U9980 ( .B1(n8803), .B2(keyinput_89), .C1(keyinput_91), .C2(n8802), 
        .A(n8801), .ZN(n8809) );
  AOI22_X1 U9981 ( .A1(n8806), .A2(keyinput_90), .B1(keyinput_92), .B2(n8805), 
        .ZN(n8804) );
  OAI221_X1 U9982 ( .B1(n8806), .B2(keyinput_90), .C1(n8805), .C2(keyinput_92), 
        .A(n8804), .ZN(n8807) );
  AOI21_X1 U9983 ( .B1(keyinput_93), .B2(n8810), .A(n8807), .ZN(n8808) );
  OAI211_X1 U9984 ( .C1(keyinput_93), .C2(n8810), .A(n8809), .B(n8808), .ZN(
        n8811) );
  OR2_X1 U9985 ( .A1(n8812), .A2(n8811), .ZN(n8817) );
  OAI22_X1 U9986 ( .A1(n10776), .A2(keyinput_97), .B1(SI_1_), .B2(keyinput_95), 
        .ZN(n8813) );
  AOI221_X1 U9987 ( .B1(n10776), .B2(keyinput_97), .C1(keyinput_95), .C2(SI_1_), .A(n8813), .ZN(n8816) );
  XNOR2_X1 U9988 ( .A(keyinput_96), .B(SI_0_), .ZN(n8815) );
  XNOR2_X1 U9989 ( .A(SI_2_), .B(keyinput_94), .ZN(n8814) );
  NAND4_X1 U9990 ( .A1(n8817), .A2(n8816), .A3(n8815), .A4(n8814), .ZN(n8818)
         );
  AOI22_X1 U9991 ( .A1(keyinput_100), .A2(n8821), .B1(n8819), .B2(n8818), .ZN(
        n8820) );
  OAI21_X1 U9992 ( .B1(n8821), .B2(keyinput_100), .A(n8820), .ZN(n8822) );
  OAI221_X1 U9993 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(n8824), .C1(n8823), .C2(
        keyinput_101), .A(n8822), .ZN(n8825) );
  OAI221_X1 U9994 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(n8827), .C1(n8826), .C2(
        keyinput_102), .A(n8825), .ZN(n8828) );
  OAI221_X1 U9995 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_103), .C1(n8830), .C2(n8829), .A(n8828), .ZN(n8831) );
  OAI221_X1 U9996 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_104), .C1(n8833), 
        .C2(n8832), .A(n8831), .ZN(n8834) );
  OAI211_X1 U9997 ( .C1(n8837), .C2(keyinput_106), .A(n8835), .B(n8834), .ZN(
        n8836) );
  AOI21_X1 U9998 ( .B1(n8837), .B2(keyinput_106), .A(n8836), .ZN(n8838) );
  AOI221_X1 U9999 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n8840), .C1(n8839), .C2(
        keyinput_108), .A(n8838), .ZN(n8841) );
  AOI221_X1 U10000 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(n8843), .C1(n8842), 
        .C2(keyinput_109), .A(n8841), .ZN(n8844) );
  AOI221_X1 U10001 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_110), .C1(
        n8846), .C2(n8845), .A(n8844), .ZN(n8847) );
  AOI221_X1 U10002 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(n8849), .C1(n8848), 
        .C2(keyinput_111), .A(n8847), .ZN(n8850) );
  AOI221_X1 U10003 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(n8852), .C1(n8851), 
        .C2(keyinput_112), .A(n8850), .ZN(n8855) );
  AOI22_X1 U10004 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_113), .B1(n6437), 
        .B2(keyinput_114), .ZN(n8853) );
  OAI221_X1 U10005 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_113), .C1(n6437), .C2(keyinput_114), .A(n8853), .ZN(n8854) );
  OAI22_X1 U10006 ( .A1(n8855), .A2(n8854), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        keyinput_115), .ZN(n8859) );
  OAI22_X1 U10007 ( .A1(n8857), .A2(keyinput_119), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(keyinput_118), .ZN(n8856) );
  AOI221_X1 U10008 ( .B1(n8857), .B2(keyinput_119), .C1(keyinput_118), .C2(
        P2_REG3_REG_0__SCAN_IN), .A(n8856), .ZN(n8858) );
  OAI221_X1 U10009 ( .B1(n8859), .B2(keyinput_115), .C1(n8859), .C2(
        P2_REG3_REG_24__SCAN_IN), .A(n8858), .ZN(n8863) );
  AOI22_X1 U10010 ( .A1(n6345), .A2(keyinput_117), .B1(keyinput_116), .B2(
        n8861), .ZN(n8860) );
  OAI221_X1 U10011 ( .B1(n6345), .B2(keyinput_117), .C1(n8861), .C2(
        keyinput_116), .A(n8860), .ZN(n8862) );
  OAI22_X1 U10012 ( .A1(keyinput_120), .A2(n9076), .B1(n8863), .B2(n8862), 
        .ZN(n8864) );
  AOI21_X1 U10013 ( .B1(keyinput_120), .B2(n9076), .A(n8864), .ZN(n8865) );
  AOI221_X1 U10014 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(n8867), .C1(n8866), 
        .C2(keyinput_121), .A(n8865), .ZN(n8868) );
  AOI221_X1 U10015 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_122), .C1(
        n9099), .C2(n8869), .A(n8868), .ZN(n8873) );
  AOI22_X1 U10016 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_123), .B1(n8871), 
        .B2(keyinput_125), .ZN(n8870) );
  OAI221_X1 U10017 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_123), .C1(n8871), .C2(keyinput_125), .A(n8870), .ZN(n8872) );
  AOI211_X1 U10018 ( .C1(P2_REG3_REG_18__SCAN_IN), .C2(keyinput_124), .A(n8873), .B(n8872), .ZN(n8874) );
  OAI21_X1 U10019 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_124), .A(n8874), 
        .ZN(n8875) );
  OAI221_X1 U10020 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(n8877), .C1(n8876), 
        .C2(keyinput_126), .A(n8875), .ZN(n8879) );
  AOI21_X1 U10021 ( .B1(keyinput_127), .B2(n8879), .A(P2_REG3_REG_15__SCAN_IN), 
        .ZN(n8881) );
  INV_X1 U10022 ( .A(keyinput_127), .ZN(n8878) );
  AOI21_X1 U10023 ( .B1(n8879), .B2(n8878), .A(keyinput_63), .ZN(n8880) );
  AOI22_X1 U10024 ( .A1(keyinput_63), .A2(n8881), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(n8880), .ZN(n8882) );
  AOI21_X1 U10025 ( .B1(n8884), .B2(n8883), .A(n8882), .ZN(n8889) );
  AOI222_X1 U10026 ( .A1(n8887), .A2(n8886), .B1(P2_DATAO_REG_11__SCAN_IN), 
        .B2(n10477), .C1(P1_STATE_REG_SCAN_IN), .C2(n8885), .ZN(n8888) );
  XNOR2_X1 U10027 ( .A(n8889), .B(n8888), .ZN(P1_U3344) );
  INV_X1 U10028 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n8894) );
  OAI211_X1 U10029 ( .C1(n10021), .C2(n10395), .A(n8891), .B(n8890), .ZN(n8892) );
  AOI21_X1 U10030 ( .B1(n8893), .B2(n10838), .A(n8892), .ZN(n8896) );
  MUX2_X1 U10031 ( .A(n8894), .B(n8896), .S(n10846), .Z(n8895) );
  OAI21_X1 U10032 ( .B1(n8899), .B2(n10469), .A(n8895), .ZN(P1_U3498) );
  INV_X1 U10033 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n8897) );
  MUX2_X1 U10034 ( .A(n8897), .B(n8896), .S(n10842), .Z(n8898) );
  OAI21_X1 U10035 ( .B1(n8899), .B2(n10419), .A(n8898), .ZN(P1_U3537) );
  XNOR2_X1 U10036 ( .A(n8901), .B(n8900), .ZN(n8903) );
  OAI222_X1 U10037 ( .A1(n10315), .A2(n10301), .B1(n10395), .B2(n9935), .C1(
        n8903), .C2(n8902), .ZN(n10414) );
  AOI21_X1 U10038 ( .B1(n9938), .B2(n10274), .A(n10414), .ZN(n8913) );
  XNOR2_X1 U10039 ( .A(n8905), .B(n8904), .ZN(n10416) );
  NAND2_X1 U10040 ( .A1(n10416), .A2(n10321), .ZN(n8912) );
  INV_X1 U10041 ( .A(n10323), .ZN(n8907) );
  AOI211_X1 U10042 ( .C1(n8908), .C2(n5239), .A(n10803), .B(n8907), .ZN(n10415) );
  INV_X1 U10043 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8909) );
  OAI22_X1 U10044 ( .A1(n10470), .A2(n10325), .B1(n8909), .B2(n10328), .ZN(
        n8910) );
  AOI21_X1 U10045 ( .B1(n10415), .B2(n10286), .A(n8910), .ZN(n8911) );
  OAI211_X1 U10046 ( .C1(n10335), .C2(n8913), .A(n8912), .B(n8911), .ZN(
        P1_U3276) );
  OAI222_X1 U10047 ( .A1(n6221), .A2(P2_U3151), .B1(n9855), .B2(n8915), .C1(
        n8914), .C2(n9856), .ZN(P2_U3275) );
  INV_X1 U10048 ( .A(n8918), .ZN(P1_U3550) );
  XOR2_X1 U10049 ( .A(n8922), .B(n8919), .Z(n10374) );
  AND2_X1 U10050 ( .A1(n10219), .A2(n8920), .ZN(n8923) );
  OAI211_X1 U10051 ( .C1(n8923), .C2(n8922), .A(n8921), .B(n10312), .ZN(n8925)
         );
  NAND2_X1 U10052 ( .A1(n10245), .A2(n10389), .ZN(n8924) );
  OAI211_X1 U10053 ( .C1(n10360), .C2(n10315), .A(n8925), .B(n8924), .ZN(
        n10371) );
  INV_X1 U10054 ( .A(n8926), .ZN(n10231) );
  INV_X1 U10055 ( .A(n10210), .ZN(n8927) );
  AOI211_X1 U10056 ( .C1(n10372), .C2(n10231), .A(n10803), .B(n8927), .ZN(
        n10370) );
  NAND2_X1 U10057 ( .A1(n10370), .A2(n10286), .ZN(n8929) );
  AOI22_X1 U10058 ( .A1(n9950), .A2(n10274), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10335), .ZN(n8928) );
  OAI211_X1 U10059 ( .C1(n9953), .C2(n10325), .A(n8929), .B(n8928), .ZN(n8930)
         );
  AOI21_X1 U10060 ( .B1(n10328), .B2(n10371), .A(n8930), .ZN(n8931) );
  OAI21_X1 U10061 ( .B1(n10374), .B2(n10307), .A(n8931), .ZN(P1_U3269) );
  INV_X1 U10062 ( .A(n9289), .ZN(n9840) );
  OAI222_X1 U10063 ( .A1(n10494), .A2(n8933), .B1(n10492), .B2(n9840), .C1(
        n8932), .C2(P1_U3086), .ZN(P1_U3325) );
  INV_X1 U10064 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8935) );
  OAI222_X1 U10065 ( .A1(n10494), .A2(n8935), .B1(n10492), .B2(n8934), .C1(
        n10116), .C2(P1_U3086), .ZN(P1_U3336) );
  OR2_X1 U10066 ( .A1(n8936), .A2(n9683), .ZN(n8937) );
  XNOR2_X1 U10067 ( .A(n9677), .B(n7270), .ZN(n8940) );
  XNOR2_X1 U10068 ( .A(n8940), .B(n9666), .ZN(n9075) );
  INV_X1 U10069 ( .A(n9075), .ZN(n8939) );
  INV_X1 U10070 ( .A(n8940), .ZN(n8941) );
  XNOR2_X1 U10071 ( .A(n9757), .B(n7270), .ZN(n8942) );
  XNOR2_X1 U10072 ( .A(n8942), .B(n9382), .ZN(n9000) );
  NAND2_X1 U10073 ( .A1(n8942), .A2(n8943), .ZN(n8944) );
  XNOR2_X1 U10074 ( .A(n9834), .B(n7270), .ZN(n8946) );
  XNOR2_X1 U10075 ( .A(n8946), .B(n9381), .ZN(n9128) );
  INV_X1 U10076 ( .A(n9128), .ZN(n8945) );
  NAND2_X1 U10077 ( .A1(n8946), .A2(n9381), .ZN(n8947) );
  XOR2_X1 U10078 ( .A(n7270), .B(n9640), .Z(n9038) );
  XNOR2_X1 U10079 ( .A(n9234), .B(n7270), .ZN(n8948) );
  NAND2_X1 U10080 ( .A1(n8948), .A2(n9636), .ZN(n9046) );
  NAND2_X1 U10081 ( .A1(n9048), .A2(n9046), .ZN(n8950) );
  INV_X1 U10082 ( .A(n8948), .ZN(n8949) );
  NAND2_X1 U10083 ( .A1(n8949), .A2(n9379), .ZN(n9047) );
  NAND2_X1 U10084 ( .A1(n8950), .A2(n9047), .ZN(n9107) );
  XNOR2_X1 U10085 ( .A(n9106), .B(n7270), .ZN(n8951) );
  XNOR2_X1 U10086 ( .A(n8951), .B(n8952), .ZN(n9110) );
  NAND2_X1 U10087 ( .A1(n9107), .A2(n9110), .ZN(n9108) );
  INV_X1 U10088 ( .A(n8951), .ZN(n8953) );
  NAND2_X1 U10089 ( .A1(n8953), .A2(n8952), .ZN(n8954) );
  NAND2_X1 U10090 ( .A1(n9108), .A2(n8954), .ZN(n9017) );
  NAND2_X1 U10091 ( .A1(n8956), .A2(n8955), .ZN(n9600) );
  XNOR2_X1 U10092 ( .A(n9600), .B(n7270), .ZN(n9016) );
  INV_X1 U10093 ( .A(n9016), .ZN(n8957) );
  NAND2_X1 U10094 ( .A1(n8957), .A2(n9378), .ZN(n8958) );
  XNOR2_X1 U10095 ( .A(n9594), .B(n7270), .ZN(n8960) );
  XNOR2_X1 U10096 ( .A(n8960), .B(n9603), .ZN(n9066) );
  INV_X1 U10097 ( .A(n9066), .ZN(n8959) );
  NAND2_X1 U10098 ( .A1(n8960), .A2(n9603), .ZN(n8961) );
  XNOR2_X1 U10099 ( .A(n9577), .B(n7270), .ZN(n8962) );
  XNOR2_X1 U10100 ( .A(n8962), .B(n9376), .ZN(n9024) );
  NAND2_X1 U10101 ( .A1(n8962), .A2(n9592), .ZN(n8963) );
  XNOR2_X1 U10102 ( .A(n9258), .B(n7270), .ZN(n8964) );
  XNOR2_X1 U10103 ( .A(n8964), .B(n9576), .ZN(n9084) );
  INV_X1 U10104 ( .A(n8964), .ZN(n8965) );
  XNOR2_X1 U10105 ( .A(n9801), .B(n8966), .ZN(n8968) );
  NAND2_X1 U10106 ( .A1(n9007), .A2(n9564), .ZN(n8971) );
  INV_X1 U10107 ( .A(n8967), .ZN(n8969) );
  NAND2_X1 U10108 ( .A1(n8969), .A2(n8968), .ZN(n8970) );
  NAND2_X1 U10109 ( .A1(n8971), .A2(n8970), .ZN(n9056) );
  XNOR2_X1 U10110 ( .A(n8972), .B(n9522), .ZN(n9057) );
  NAND2_X1 U10111 ( .A1(n9056), .A2(n9057), .ZN(n8974) );
  NAND2_X1 U10112 ( .A1(n8972), .A2(n9554), .ZN(n8973) );
  NAND2_X1 U10113 ( .A1(n8974), .A2(n8973), .ZN(n9030) );
  XNOR2_X1 U10114 ( .A(n8976), .B(n9542), .ZN(n9031) );
  NAND2_X1 U10115 ( .A1(n8976), .A2(n8975), .ZN(n8977) );
  NAND2_X1 U10116 ( .A1(n8978), .A2(n8981), .ZN(n9509) );
  INV_X1 U10117 ( .A(n9309), .ZN(n9277) );
  NAND2_X1 U10118 ( .A1(n9277), .A2(n9508), .ZN(n8979) );
  MUX2_X1 U10119 ( .A(n8981), .B(n9277), .S(n7270), .Z(n8982) );
  NOR2_X1 U10120 ( .A1(n8983), .A2(n9122), .ZN(n8984) );
  AOI21_X1 U10121 ( .B1(n9122), .B2(n8983), .A(n8984), .ZN(n8994) );
  AOI22_X1 U10122 ( .A1(n9506), .A2(n9132), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8987) );
  NAND2_X1 U10123 ( .A1(n9136), .A2(n9487), .ZN(n8986) );
  OAI211_X1 U10124 ( .C1(n8988), .C2(n9134), .A(n8987), .B(n8986), .ZN(n8989)
         );
  AOI21_X1 U10125 ( .B1(n9282), .B2(n9079), .A(n8989), .ZN(n8990) );
  OAI21_X1 U10126 ( .B1(n8991), .B2(n9127), .A(n8990), .ZN(P2_U3160) );
  OAI211_X1 U10127 ( .C1(n8995), .C2(n8994), .A(n8993), .B(n9109), .ZN(n8999)
         );
  AOI22_X1 U10128 ( .A1(n9521), .A2(n9132), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8996) );
  OAI21_X1 U10129 ( .B1(n9499), .B2(n9134), .A(n8996), .ZN(n8997) );
  AOI21_X1 U10130 ( .B1(n9500), .B2(n9136), .A(n8997), .ZN(n8998) );
  OAI211_X1 U10131 ( .C1(n9791), .C2(n9139), .A(n8999), .B(n8998), .ZN(
        P2_U3154) );
  XOR2_X1 U10132 ( .A(n9001), .B(n9000), .Z(n9006) );
  AOI22_X1 U10133 ( .A1(n9383), .A2(n9132), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n9003) );
  NAND2_X1 U10134 ( .A1(n9136), .A2(n9668), .ZN(n9002) );
  OAI211_X1 U10135 ( .C1(n9667), .C2(n9134), .A(n9003), .B(n9002), .ZN(n9004)
         );
  AOI21_X1 U10136 ( .B1(n9757), .B2(n9079), .A(n9004), .ZN(n9005) );
  OAI21_X1 U10137 ( .B1(n9006), .B2(n9127), .A(n9005), .ZN(P2_U3155) );
  XNOR2_X1 U10138 ( .A(n9007), .B(n9539), .ZN(n9013) );
  AOI22_X1 U10139 ( .A1(n9522), .A2(n9111), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n9009) );
  NAND2_X1 U10140 ( .A1(n9136), .A2(n9557), .ZN(n9008) );
  OAI211_X1 U10141 ( .C1(n9576), .C2(n9113), .A(n9009), .B(n9008), .ZN(n9010)
         );
  AOI21_X1 U10142 ( .B1(n9011), .B2(n9079), .A(n9010), .ZN(n9012) );
  OAI21_X1 U10143 ( .B1(n9013), .B2(n9127), .A(n9012), .ZN(P2_U3156) );
  OAI211_X1 U10144 ( .C1(n9017), .C2(n9016), .A(n9015), .B(n9109), .ZN(n9022)
         );
  NOR2_X1 U10145 ( .A1(n9018), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9463) );
  AOI21_X1 U10146 ( .B1(n9377), .B2(n9111), .A(n9463), .ZN(n9019) );
  OAI21_X1 U10147 ( .B1(n9623), .B2(n9113), .A(n9019), .ZN(n9020) );
  AOI21_X1 U10148 ( .B1(n9606), .B2(n9136), .A(n9020), .ZN(n9021) );
  OAI211_X1 U10149 ( .C1(n9817), .C2(n9139), .A(n9022), .B(n9021), .ZN(
        P2_U3159) );
  XOR2_X1 U10150 ( .A(n9023), .B(n9024), .Z(n9029) );
  AOI22_X1 U10151 ( .A1(n9375), .A2(n9111), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n9026) );
  NAND2_X1 U10152 ( .A1(n9136), .A2(n9578), .ZN(n9025) );
  OAI211_X1 U10153 ( .C1(n9603), .C2(n9113), .A(n9026), .B(n9025), .ZN(n9027)
         );
  AOI21_X1 U10154 ( .B1(n9577), .B2(n9079), .A(n9027), .ZN(n9028) );
  OAI21_X1 U10155 ( .B1(n9029), .B2(n9127), .A(n9028), .ZN(P2_U3163) );
  XOR2_X1 U10156 ( .A(n9031), .B(n9030), .Z(n9036) );
  AOI22_X1 U10157 ( .A1(n9111), .A2(n9521), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n9033) );
  NAND2_X1 U10158 ( .A1(n9136), .A2(n9526), .ZN(n9032) );
  OAI211_X1 U10159 ( .C1(n9554), .C2(n9113), .A(n9033), .B(n9032), .ZN(n9034)
         );
  AOI21_X1 U10160 ( .B1(n9518), .B2(n9079), .A(n9034), .ZN(n9035) );
  OAI21_X1 U10161 ( .B1(n9036), .B2(n9127), .A(n9035), .ZN(P2_U3165) );
  XNOR2_X1 U10162 ( .A(n9038), .B(n9648), .ZN(n9039) );
  XNOR2_X1 U10163 ( .A(n9037), .B(n9039), .ZN(n9045) );
  NAND2_X1 U10164 ( .A1(n9136), .A2(n9641), .ZN(n9042) );
  NAND2_X1 U10165 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n10734)
         );
  INV_X1 U10166 ( .A(n10734), .ZN(n9040) );
  AOI21_X1 U10167 ( .B1(n9381), .B2(n9132), .A(n9040), .ZN(n9041) );
  OAI211_X1 U10168 ( .C1(n9636), .C2(n9134), .A(n9042), .B(n9041), .ZN(n9043)
         );
  AOI21_X1 U10169 ( .B1(n9640), .B2(n9079), .A(n9043), .ZN(n9044) );
  OAI21_X1 U10170 ( .B1(n9045), .B2(n9127), .A(n9044), .ZN(P2_U3166) );
  NAND2_X1 U10171 ( .A1(n9047), .A2(n9046), .ZN(n9049) );
  XOR2_X1 U10172 ( .A(n9049), .B(n9048), .Z(n9055) );
  NAND2_X1 U10173 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n10750)
         );
  INV_X1 U10174 ( .A(n10750), .ZN(n9050) );
  AOI21_X1 U10175 ( .B1(n9380), .B2(n9132), .A(n9050), .ZN(n9052) );
  NAND2_X1 U10176 ( .A1(n9136), .A2(n9628), .ZN(n9051) );
  OAI211_X1 U10177 ( .C1(n9623), .C2(n9134), .A(n9052), .B(n9051), .ZN(n9053)
         );
  AOI21_X1 U10178 ( .B1(n9234), .B2(n9079), .A(n9053), .ZN(n9054) );
  OAI21_X1 U10179 ( .B1(n9055), .B2(n9127), .A(n9054), .ZN(P2_U3168) );
  XOR2_X1 U10180 ( .A(n9057), .B(n9056), .Z(n9062) );
  AOI22_X1 U10181 ( .A1(n9542), .A2(n9111), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n9059) );
  NAND2_X1 U10182 ( .A1(n9136), .A2(n9532), .ZN(n9058) );
  OAI211_X1 U10183 ( .C1(n9564), .C2(n9113), .A(n9059), .B(n9058), .ZN(n9060)
         );
  AOI21_X1 U10184 ( .B1(n9531), .B2(n9079), .A(n9060), .ZN(n9061) );
  OAI21_X1 U10185 ( .B1(n9062), .B2(n9127), .A(n9061), .ZN(P2_U3169) );
  INV_X1 U10186 ( .A(n9063), .ZN(n9064) );
  AOI21_X1 U10187 ( .B1(n9066), .B2(n9065), .A(n9064), .ZN(n9071) );
  AOI22_X1 U10188 ( .A1(n9111), .A2(n9376), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n9068) );
  NAND2_X1 U10189 ( .A1(n9136), .A2(n9595), .ZN(n9067) );
  OAI211_X1 U10190 ( .C1(n9613), .C2(n9113), .A(n9068), .B(n9067), .ZN(n9069)
         );
  AOI21_X1 U10191 ( .B1(n9594), .B2(n9079), .A(n9069), .ZN(n9070) );
  OAI21_X1 U10192 ( .B1(n9071), .B2(n9127), .A(n9070), .ZN(P2_U3173) );
  INV_X1 U10193 ( .A(n9072), .ZN(n9073) );
  AOI21_X1 U10194 ( .B1(n9075), .B2(n9074), .A(n9073), .ZN(n9082) );
  NOR2_X1 U10195 ( .A1(n8943), .A2(n9134), .ZN(n9078) );
  OAI22_X1 U10196 ( .A1(n9113), .A2(n9683), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9076), .ZN(n9077) );
  AOI211_X1 U10197 ( .C1(n9687), .C2(n9136), .A(n9078), .B(n9077), .ZN(n9081)
         );
  NAND2_X1 U10198 ( .A1(n9677), .A2(n9079), .ZN(n9080) );
  OAI211_X1 U10199 ( .C1(n9082), .C2(n9127), .A(n9081), .B(n9080), .ZN(
        P2_U3174) );
  AOI21_X1 U10200 ( .B1(n9083), .B2(n9084), .A(n9127), .ZN(n9086) );
  NAND2_X1 U10201 ( .A1(n9086), .A2(n9085), .ZN(n9090) );
  AOI22_X1 U10202 ( .A1(n9376), .A2(n9132), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n9087) );
  OAI21_X1 U10203 ( .B1(n9564), .B2(n9134), .A(n9087), .ZN(n9088) );
  AOI21_X1 U10204 ( .B1(n9567), .B2(n9136), .A(n9088), .ZN(n9089) );
  OAI211_X1 U10205 ( .C1(n9805), .C2(n9139), .A(n9090), .B(n9089), .ZN(
        P2_U3175) );
  OAI22_X1 U10206 ( .A1(n9093), .A2(n9386), .B1(n9092), .B2(n9091), .ZN(n9097)
         );
  XNOR2_X1 U10207 ( .A(n9095), .B(n9094), .ZN(n9096) );
  XNOR2_X1 U10208 ( .A(n9097), .B(n9096), .ZN(n9098) );
  NAND2_X1 U10209 ( .A1(n9098), .A2(n9109), .ZN(n9105) );
  NOR2_X1 U10210 ( .A1(n9683), .A2(n9134), .ZN(n9102) );
  OAI22_X1 U10211 ( .A1(n9113), .A2(n9100), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9099), .ZN(n9101) );
  AOI211_X1 U10212 ( .C1(n9103), .C2(n9136), .A(n9102), .B(n9101), .ZN(n9104)
         );
  OAI211_X1 U10213 ( .C1(n9774), .C2(n9139), .A(n9105), .B(n9104), .ZN(
        P2_U3176) );
  OAI211_X1 U10214 ( .C1(n9107), .C2(n9110), .A(n9108), .B(n9109), .ZN(n9116)
         );
  AND2_X1 U10215 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n10756) );
  AOI21_X1 U10216 ( .B1(n9378), .B2(n9111), .A(n10756), .ZN(n9112) );
  OAI21_X1 U10217 ( .B1(n9636), .B2(n9113), .A(n9112), .ZN(n9114) );
  AOI21_X1 U10218 ( .B1(n9616), .B2(n9136), .A(n9114), .ZN(n9115) );
  OAI211_X1 U10219 ( .C1(n9821), .C2(n9139), .A(n9116), .B(n9115), .ZN(
        P2_U3178) );
  AOI21_X1 U10220 ( .B1(n9117), .B2(n9118), .A(n9127), .ZN(n9120) );
  NAND2_X1 U10221 ( .A1(n9120), .A2(n9119), .ZN(n9125) );
  AOI22_X1 U10222 ( .A1(n9542), .A2(n9132), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n9121) );
  OAI21_X1 U10223 ( .B1(n9122), .B2(n9134), .A(n9121), .ZN(n9123) );
  AOI21_X1 U10224 ( .B1(n9513), .B2(n9136), .A(n9123), .ZN(n9124) );
  OAI211_X1 U10225 ( .C1(n9515), .C2(n9139), .A(n9125), .B(n9124), .ZN(
        P2_U3180) );
  AOI21_X1 U10226 ( .B1(n9126), .B2(n9128), .A(n9127), .ZN(n9130) );
  NAND2_X1 U10227 ( .A1(n9130), .A2(n9129), .ZN(n9138) );
  NAND2_X1 U10228 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n10718)
         );
  INV_X1 U10229 ( .A(n10718), .ZN(n9131) );
  AOI21_X1 U10230 ( .B1(n9382), .B2(n9132), .A(n9131), .ZN(n9133) );
  OAI21_X1 U10231 ( .B1(n9648), .B2(n9134), .A(n9133), .ZN(n9135) );
  AOI21_X1 U10232 ( .B1(n9653), .B2(n9136), .A(n9135), .ZN(n9137) );
  OAI211_X1 U10233 ( .C1(n9834), .C2(n9139), .A(n9138), .B(n9137), .ZN(
        P2_U3181) );
  MUX2_X1 U10234 ( .A(n9499), .B(n9489), .S(n9269), .Z(n9283) );
  MUX2_X1 U10235 ( .A(n9308), .B(n5003), .S(n9284), .Z(n9281) );
  INV_X1 U10236 ( .A(n9263), .ZN(n9140) );
  MUX2_X1 U10237 ( .A(n9261), .B(n9140), .S(n9269), .Z(n9265) );
  INV_X1 U10238 ( .A(n9259), .ZN(n9142) );
  NAND2_X1 U10239 ( .A1(n9144), .A2(n9143), .ZN(n9145) );
  NAND3_X1 U10240 ( .A1(n9147), .A2(n9145), .A3(n9150), .ZN(n9146) );
  NAND2_X1 U10241 ( .A1(n9146), .A2(n9148), .ZN(n9153) );
  INV_X1 U10242 ( .A(n9147), .ZN(n9149) );
  NAND2_X1 U10243 ( .A1(n9149), .A2(n9148), .ZN(n9151) );
  NAND2_X1 U10244 ( .A1(n9151), .A2(n9150), .ZN(n9152) );
  NOR2_X1 U10245 ( .A1(n9155), .A2(n9154), .ZN(n9156) );
  MUX2_X1 U10246 ( .A(n9157), .B(n9156), .S(n9269), .Z(n9158) );
  NAND3_X1 U10247 ( .A1(n9166), .A2(n7816), .A3(n9159), .ZN(n9161) );
  NAND3_X1 U10248 ( .A1(n9161), .A2(n9162), .A3(n9160), .ZN(n9164) );
  AND2_X1 U10249 ( .A1(n9162), .A2(n9177), .ZN(n9163) );
  MUX2_X1 U10250 ( .A(n9164), .B(n9163), .S(n9284), .Z(n9171) );
  NAND3_X1 U10251 ( .A1(n9166), .A2(n7816), .A3(n9165), .ZN(n9168) );
  NAND4_X1 U10252 ( .A1(n9168), .A2(n9284), .A3(n9173), .A4(n9167), .ZN(n9170)
         );
  INV_X1 U10253 ( .A(n9172), .ZN(n9169) );
  AOI21_X1 U10254 ( .B1(n9171), .B2(n9170), .A(n9169), .ZN(n9182) );
  AOI21_X1 U10255 ( .B1(n9173), .B2(n9172), .A(n9284), .ZN(n9181) );
  NAND2_X1 U10256 ( .A1(n9174), .A2(n9194), .ZN(n9176) );
  NAND2_X1 U10257 ( .A1(n9185), .A2(n9184), .ZN(n9175) );
  MUX2_X1 U10258 ( .A(n9176), .B(n9175), .S(n9269), .Z(n9196) );
  NOR2_X1 U10259 ( .A1(n9177), .A2(n9284), .ZN(n9178) );
  OR2_X1 U10260 ( .A1(n9336), .A2(n9178), .ZN(n9179) );
  NOR2_X1 U10261 ( .A1(n9196), .A2(n9179), .ZN(n9180) );
  OAI21_X1 U10262 ( .B1(n9182), .B2(n9181), .A(n9180), .ZN(n9189) );
  AND2_X1 U10263 ( .A1(n9184), .A2(n9183), .ZN(n9186) );
  OAI211_X1 U10264 ( .C1(n9196), .C2(n9186), .A(n9197), .B(n9185), .ZN(n9187)
         );
  NAND2_X1 U10265 ( .A1(n9187), .A2(n9284), .ZN(n9188) );
  NAND3_X1 U10266 ( .A1(n9199), .A2(n4995), .A3(n9202), .ZN(n9190) );
  NAND2_X1 U10267 ( .A1(n9190), .A2(n9200), .ZN(n9205) );
  INV_X1 U10268 ( .A(n9191), .ZN(n9192) );
  NOR2_X1 U10269 ( .A1(n9193), .A2(n9192), .ZN(n9195) );
  OAI211_X1 U10270 ( .C1(n9196), .C2(n9195), .A(n4995), .B(n9194), .ZN(n9198)
         );
  OAI21_X1 U10271 ( .B1(n9199), .B2(n9198), .A(n9197), .ZN(n9203) );
  INV_X1 U10272 ( .A(n9200), .ZN(n9201) );
  AOI21_X1 U10273 ( .B1(n9203), .B2(n9202), .A(n9201), .ZN(n9204) );
  MUX2_X1 U10274 ( .A(n9205), .B(n9204), .S(n9269), .Z(n9210) );
  MUX2_X1 U10275 ( .A(n9207), .B(n9206), .S(n9284), .Z(n9208) );
  OAI211_X1 U10276 ( .C1(n9210), .C2(n9209), .A(n9690), .B(n9208), .ZN(n9213)
         );
  MUX2_X1 U10277 ( .A(n9269), .B(n9666), .S(n9677), .Z(n9211) );
  OAI21_X1 U10278 ( .B1(n9284), .B2(n9383), .A(n9211), .ZN(n9212) );
  NAND2_X1 U10279 ( .A1(n9213), .A2(n9212), .ZN(n9218) );
  NAND2_X1 U10280 ( .A1(n9757), .A2(n9269), .ZN(n9214) );
  OAI21_X1 U10281 ( .B1(n8943), .B2(n9269), .A(n9214), .ZN(n9215) );
  OAI21_X1 U10282 ( .B1(n9649), .B2(n9216), .A(n9219), .ZN(n9217) );
  INV_X1 U10283 ( .A(n9219), .ZN(n9223) );
  OAI21_X1 U10284 ( .B1(n9381), .B2(n9269), .A(n9220), .ZN(n9222) );
  OAI21_X1 U10285 ( .B1(n9284), .B2(n9667), .A(n9834), .ZN(n9221) );
  AOI22_X1 U10286 ( .A1(n9223), .A2(n9664), .B1(n9222), .B2(n9221), .ZN(n9224)
         );
  MUX2_X1 U10287 ( .A(n9226), .B(n9225), .S(n9269), .Z(n9227) );
  MUX2_X1 U10288 ( .A(n9379), .B(n9234), .S(n9284), .Z(n9228) );
  INV_X1 U10289 ( .A(n9228), .ZN(n9229) );
  NAND3_X1 U10290 ( .A1(n9233), .A2(n9237), .A3(n9234), .ZN(n9231) );
  NAND3_X1 U10291 ( .A1(n9235), .A2(n9615), .A3(n9636), .ZN(n9230) );
  NAND3_X1 U10292 ( .A1(n9231), .A2(n9232), .A3(n9230), .ZN(n9240) );
  NAND3_X1 U10293 ( .A1(n9233), .A2(n9379), .A3(n9232), .ZN(n9238) );
  INV_X1 U10294 ( .A(n9234), .ZN(n9825) );
  NAND3_X1 U10295 ( .A1(n9235), .A2(n9615), .A3(n9825), .ZN(n9236) );
  NAND3_X1 U10296 ( .A1(n9238), .A2(n9237), .A3(n9236), .ZN(n9239) );
  MUX2_X1 U10297 ( .A(n9240), .B(n9239), .S(n9284), .Z(n9246) );
  INV_X1 U10298 ( .A(n9600), .ZN(n9605) );
  INV_X1 U10299 ( .A(n9241), .ZN(n9242) );
  MUX2_X1 U10300 ( .A(n9243), .B(n9242), .S(n9284), .Z(n9244) );
  NOR2_X1 U10301 ( .A1(n9328), .A2(n9244), .ZN(n9245) );
  OAI21_X1 U10302 ( .B1(n9246), .B2(n9605), .A(n9245), .ZN(n9256) );
  MUX2_X1 U10303 ( .A(n9376), .B(n9577), .S(n9284), .Z(n9253) );
  MUX2_X1 U10305 ( .A(n9249), .B(n9248), .S(n9284), .Z(n9250) );
  OAI21_X1 U10306 ( .B1(n9253), .B2(n4954), .A(n9250), .ZN(n9252) );
  INV_X1 U10307 ( .A(n9252), .ZN(n9255) );
  AOI22_X1 U10308 ( .A1(n9256), .A2(n9255), .B1(n9254), .B2(n9253), .ZN(n9257)
         );
  MUX2_X1 U10309 ( .A(n9375), .B(n9258), .S(n9269), .Z(n9260) );
  AND2_X1 U10310 ( .A1(n9260), .A2(n9259), .ZN(n9264) );
  INV_X1 U10311 ( .A(n9261), .ZN(n9262) );
  NAND2_X1 U10312 ( .A1(n9531), .A2(n9554), .ZN(n9267) );
  MUX2_X1 U10313 ( .A(n9267), .B(n9266), .S(n9284), .Z(n9268) );
  INV_X1 U10314 ( .A(n9272), .ZN(n9275) );
  NAND2_X1 U10315 ( .A1(n9518), .A2(n9542), .ZN(n9271) );
  MUX2_X1 U10316 ( .A(n9542), .B(n9518), .S(n9269), .Z(n9270) );
  OAI21_X1 U10317 ( .B1(n9275), .B2(n9274), .A(n9273), .ZN(n9276) );
  NAND2_X1 U10318 ( .A1(n9276), .A2(n9509), .ZN(n9279) );
  MUX2_X1 U10319 ( .A(n9508), .B(n9277), .S(n9284), .Z(n9278) );
  NAND3_X1 U10320 ( .A1(n9279), .A2(n9494), .A3(n9278), .ZN(n9280) );
  NAND2_X1 U10321 ( .A1(n9281), .A2(n9280), .ZN(n9285) );
  OAI211_X1 U10322 ( .C1(n9283), .C2(n9282), .A(n9292), .B(n9285), .ZN(n9288)
         );
  INV_X1 U10323 ( .A(n9283), .ZN(n9293) );
  NAND3_X1 U10324 ( .A1(n9319), .A2(n9499), .A3(n9293), .ZN(n9287) );
  NAND2_X1 U10325 ( .A1(n9289), .A2(n6275), .ZN(n9291) );
  NAND2_X1 U10326 ( .A1(n6258), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n9290) );
  NOR2_X1 U10327 ( .A1(n9787), .A2(n9373), .ZN(n9355) );
  INV_X1 U10328 ( .A(n9292), .ZN(n9294) );
  INV_X1 U10329 ( .A(n9373), .ZN(n9297) );
  NOR2_X1 U10330 ( .A1(n9298), .A2(n9297), .ZN(n9354) );
  NAND2_X1 U10331 ( .A1(n9835), .A2(n6275), .ZN(n9300) );
  NAND2_X1 U10332 ( .A1(n6258), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n9299) );
  AND2_X2 U10333 ( .A1(n9300), .A2(n9299), .ZN(n9784) );
  NAND2_X1 U10334 ( .A1(n6267), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9303) );
  NAND2_X1 U10335 ( .A1(n6595), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9302) );
  NAND2_X1 U10336 ( .A1(n6547), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9301) );
  NAND4_X1 U10337 ( .A1(n9304), .A2(n9303), .A3(n9302), .A4(n9301), .ZN(n9472)
         );
  NAND2_X1 U10338 ( .A1(n9784), .A2(n9472), .ZN(n9356) );
  INV_X1 U10339 ( .A(n9784), .ZN(n9321) );
  INV_X1 U10340 ( .A(n9472), .ZN(n9305) );
  NAND2_X1 U10341 ( .A1(n9306), .A2(n9357), .ZN(n9363) );
  NAND3_X1 U10342 ( .A1(n9307), .A2(n9508), .A3(n5003), .ZN(n9313) );
  INV_X1 U10343 ( .A(n9308), .ZN(n9310) );
  OAI21_X1 U10344 ( .B1(n9310), .B2(n9309), .A(n5003), .ZN(n9311) );
  NAND3_X1 U10345 ( .A1(n9313), .A2(n9312), .A3(n9311), .ZN(n9315) );
  NAND2_X1 U10346 ( .A1(n9315), .A2(n9314), .ZN(n9318) );
  INV_X1 U10347 ( .A(n9316), .ZN(n9317) );
  AOI211_X1 U10348 ( .C1(n9319), .C2(n9318), .A(n9317), .B(n9355), .ZN(n9320)
         );
  OAI211_X1 U10349 ( .C1(n9787), .C2(n9321), .A(n9320), .B(n9356), .ZN(n9325)
         );
  INV_X1 U10350 ( .A(n9354), .ZN(n9322) );
  INV_X1 U10351 ( .A(n9326), .ZN(n9327) );
  INV_X1 U10352 ( .A(n9690), .ZN(n9679) );
  NAND3_X1 U10353 ( .A1(n9331), .A2(n9330), .A3(n9329), .ZN(n9335) );
  NAND4_X1 U10354 ( .A1(n5190), .A2(n9333), .A3(n7816), .A4(n9332), .ZN(n9334)
         );
  NOR2_X1 U10355 ( .A1(n9335), .A2(n9334), .ZN(n9339) );
  INV_X1 U10356 ( .A(n9336), .ZN(n9338) );
  NAND4_X1 U10357 ( .A1(n9339), .A2(n9338), .A3(n5110), .A4(n9337), .ZN(n9341)
         );
  NOR2_X1 U10358 ( .A1(n9341), .A2(n9340), .ZN(n9342) );
  NAND3_X1 U10359 ( .A1(n9344), .A2(n9343), .A3(n9342), .ZN(n9345) );
  NOR4_X1 U10360 ( .A1(n9649), .A2(n9664), .A3(n9679), .A4(n9345), .ZN(n9346)
         );
  NAND3_X1 U10361 ( .A1(n9615), .A2(n9638), .A3(n9346), .ZN(n9347) );
  NOR4_X1 U10362 ( .A1(n5360), .A2(n9624), .A3(n9605), .A4(n9347), .ZN(n9348)
         );
  NAND3_X1 U10363 ( .A1(n9565), .A2(n5366), .A3(n9348), .ZN(n9349) );
  NOR4_X1 U10364 ( .A1(n9528), .A2(n9547), .A3(n9555), .A4(n9349), .ZN(n9350)
         );
  NAND4_X1 U10365 ( .A1(n9351), .A2(n9494), .A3(n9350), .A4(n9509), .ZN(n9352)
         );
  INV_X1 U10366 ( .A(n9356), .ZN(n9359) );
  INV_X1 U10367 ( .A(n9357), .ZN(n9358) );
  NOR2_X1 U10368 ( .A1(n9359), .A2(n9358), .ZN(n9360) );
  AOI21_X1 U10369 ( .B1(n9361), .B2(n9360), .A(n7262), .ZN(n9362) );
  XNOR2_X1 U10370 ( .A(n9364), .B(n9464), .ZN(n9372) );
  INV_X1 U10371 ( .A(n9365), .ZN(n9371) );
  NAND3_X1 U10372 ( .A1(n9367), .A2(n9366), .A3(n6601), .ZN(n9368) );
  OAI211_X1 U10373 ( .C1(n9369), .C2(n9371), .A(n9368), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9370) );
  OAI21_X1 U10374 ( .B1(n9372), .B2(n9371), .A(n9370), .ZN(P2_U3296) );
  MUX2_X1 U10375 ( .A(n9472), .B(P2_DATAO_REG_31__SCAN_IN), .S(n10766), .Z(
        P2_U3522) );
  MUX2_X1 U10376 ( .A(n9373), .B(P2_DATAO_REG_30__SCAN_IN), .S(n10766), .Z(
        P2_U3521) );
  MUX2_X1 U10377 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n9374), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10378 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n9506), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10379 ( .A(n9521), .B(P2_DATAO_REG_26__SCAN_IN), .S(n10766), .Z(
        P2_U3517) );
  MUX2_X1 U10380 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n9542), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10381 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n9522), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10382 ( .A(n9539), .B(P2_DATAO_REG_23__SCAN_IN), .S(n10766), .Z(
        P2_U3514) );
  MUX2_X1 U10383 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9375), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10384 ( .A(n9376), .B(P2_DATAO_REG_21__SCAN_IN), .S(n10766), .Z(
        P2_U3512) );
  MUX2_X1 U10385 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9377), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10386 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n9378), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10387 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9379), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10388 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9380), .S(n9394), .Z(
        P2_U3507) );
  MUX2_X1 U10389 ( .A(n9381), .B(P2_DATAO_REG_15__SCAN_IN), .S(n10766), .Z(
        P2_U3506) );
  MUX2_X1 U10390 ( .A(n9382), .B(P2_DATAO_REG_14__SCAN_IN), .S(n10766), .Z(
        P2_U3505) );
  MUX2_X1 U10391 ( .A(n9383), .B(P2_DATAO_REG_13__SCAN_IN), .S(n10766), .Z(
        P2_U3504) );
  MUX2_X1 U10392 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n9384), .S(n9394), .Z(
        P2_U3503) );
  MUX2_X1 U10393 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n9385), .S(n9394), .Z(
        P2_U3502) );
  MUX2_X1 U10394 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n9386), .S(n9394), .Z(
        P2_U3501) );
  MUX2_X1 U10395 ( .A(n9387), .B(P2_DATAO_REG_8__SCAN_IN), .S(n10766), .Z(
        P2_U3499) );
  MUX2_X1 U10396 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n9388), .S(n9394), .Z(
        P2_U3498) );
  MUX2_X1 U10397 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n9389), .S(n9394), .Z(
        P2_U3497) );
  MUX2_X1 U10398 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n9390), .S(n9394), .Z(
        P2_U3496) );
  MUX2_X1 U10399 ( .A(n9391), .B(P2_DATAO_REG_3__SCAN_IN), .S(n10766), .Z(
        P2_U3494) );
  MUX2_X1 U10400 ( .A(n9392), .B(P2_DATAO_REG_2__SCAN_IN), .S(n10766), .Z(
        P2_U3493) );
  MUX2_X1 U10401 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n9393), .S(n9394), .Z(
        P2_U3492) );
  MUX2_X1 U10402 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n6552), .S(n9394), .Z(
        P2_U3491) );
  INV_X1 U10403 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9747) );
  AOI22_X1 U10404 ( .A1(n10721), .A2(n9747), .B1(P2_REG1_REG_16__SCAN_IN), 
        .B2(n9433), .ZN(n10724) );
  NAND2_X1 U10405 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n9437), .ZN(n9406) );
  INV_X1 U10406 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9759) );
  AOI22_X1 U10407 ( .A1(n10689), .A2(n9759), .B1(P2_REG1_REG_14__SCAN_IN), 
        .B2(n9437), .ZN(n10692) );
  INV_X1 U10408 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9403) );
  AOI22_X1 U10409 ( .A1(n10657), .A2(n9403), .B1(P2_REG1_REG_12__SCAN_IN), 
        .B2(n9441), .ZN(n10660) );
  NAND2_X1 U10410 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n9417), .ZN(n9400) );
  AOI22_X1 U10411 ( .A1(n10623), .A2(n9395), .B1(P2_REG1_REG_10__SCAN_IN), 
        .B2(n9417), .ZN(n10631) );
  NAND2_X1 U10412 ( .A1(n9397), .A2(n9396), .ZN(n9399) );
  NAND2_X1 U10413 ( .A1(n9399), .A2(n9398), .ZN(n10630) );
  NAND2_X1 U10414 ( .A1(n10631), .A2(n10630), .ZN(n10629) );
  NAND2_X1 U10415 ( .A1(n9400), .A2(n10629), .ZN(n9401) );
  NAND2_X1 U10416 ( .A1(n5058), .A2(n9401), .ZN(n9402) );
  XNOR2_X1 U10417 ( .A(n10641), .B(n9401), .ZN(n10646) );
  NAND2_X1 U10418 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n10646), .ZN(n10645) );
  NAND2_X1 U10419 ( .A1(n9439), .A2(n9404), .ZN(n9405) );
  NAND2_X1 U10420 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n10675), .ZN(n10674) );
  NAND2_X1 U10421 ( .A1(n9405), .A2(n10674), .ZN(n10691) );
  NAND2_X1 U10422 ( .A1(n10692), .A2(n10691), .ZN(n10690) );
  NAND2_X1 U10423 ( .A1(n9406), .A2(n10690), .ZN(n9407) );
  NAND2_X1 U10424 ( .A1(n9435), .A2(n9407), .ZN(n9408) );
  XNOR2_X1 U10425 ( .A(n10705), .B(n9407), .ZN(n10707) );
  NAND2_X1 U10426 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n10707), .ZN(n10706) );
  NAND2_X1 U10427 ( .A1(n9408), .A2(n10706), .ZN(n10723) );
  NAND2_X1 U10428 ( .A1(n10724), .A2(n10723), .ZN(n10722) );
  OAI21_X1 U10429 ( .B1(n10721), .B2(n9747), .A(n10722), .ZN(n9409) );
  NAND2_X1 U10430 ( .A1(n9455), .A2(n9409), .ZN(n9410) );
  XNOR2_X1 U10431 ( .A(n10738), .B(n9409), .ZN(n10740) );
  NAND2_X1 U10432 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n10740), .ZN(n10739) );
  NAND2_X1 U10433 ( .A1(n9410), .A2(n10739), .ZN(n10754) );
  XNOR2_X1 U10434 ( .A(n10767), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n10753) );
  AOI22_X1 U10435 ( .A1(n10754), .A2(n10753), .B1(P2_REG1_REG_18__SCAN_IN), 
        .B2(n10771), .ZN(n9411) );
  XNOR2_X1 U10436 ( .A(n9464), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n9430) );
  XNOR2_X1 U10437 ( .A(n9411), .B(n9430), .ZN(n9470) );
  INV_X1 U10438 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n10714) );
  NOR2_X1 U10439 ( .A1(n9413), .A2(n9412), .ZN(n9415) );
  NAND2_X1 U10440 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n9417), .ZN(n9416) );
  OAI21_X1 U10441 ( .B1(n9417), .B2(P2_REG2_REG_10__SCAN_IN), .A(n9416), .ZN(
        n10635) );
  NOR2_X1 U10442 ( .A1(n10641), .A2(n9418), .ZN(n9419) );
  MUX2_X1 U10443 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n8534), .S(n10657), .Z(
        n10667) );
  NOR2_X1 U10444 ( .A1(n10673), .A2(n9420), .ZN(n9421) );
  INV_X1 U10445 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10682) );
  NAND2_X1 U10446 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n9437), .ZN(n9422) );
  OAI21_X1 U10447 ( .B1(n9437), .B2(P2_REG2_REG_14__SCAN_IN), .A(n9422), .ZN(
        n10699) );
  INV_X1 U10448 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9424) );
  MUX2_X1 U10449 ( .A(n9424), .B(P2_REG2_REG_16__SCAN_IN), .S(n10721), .Z(
        n9425) );
  INV_X1 U10450 ( .A(n9425), .ZN(n10731) );
  NOR2_X1 U10451 ( .A1(n10730), .A2(n5557), .ZN(n9426) );
  MUX2_X1 U10452 ( .A(P2_REG2_REG_18__SCAN_IN), .B(n9427), .S(n10767), .Z(
        n10760) );
  INV_X1 U10453 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9427) );
  INV_X1 U10454 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9429) );
  MUX2_X1 U10455 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n9429), .S(n9464), .Z(n9432) );
  INV_X1 U10456 ( .A(n9430), .ZN(n9431) );
  MUX2_X1 U10457 ( .A(n9432), .B(n9431), .S(n6601), .Z(n9459) );
  MUX2_X1 U10458 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n6601), .Z(n9454) );
  XNOR2_X1 U10459 ( .A(n9454), .B(n10738), .ZN(n10743) );
  MUX2_X1 U10460 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n6601), .Z(n9434) );
  OR2_X1 U10461 ( .A1(n9434), .A2(n9433), .ZN(n9453) );
  XNOR2_X1 U10462 ( .A(n9434), .B(n10721), .ZN(n10727) );
  MUX2_X1 U10463 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n6601), .Z(n9436) );
  OR2_X1 U10464 ( .A1(n9436), .A2(n9435), .ZN(n9452) );
  XNOR2_X1 U10465 ( .A(n9436), .B(n10705), .ZN(n10710) );
  MUX2_X1 U10466 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n6601), .Z(n9438) );
  OR2_X1 U10467 ( .A1(n9438), .A2(n9437), .ZN(n9451) );
  XNOR2_X1 U10468 ( .A(n9438), .B(n10689), .ZN(n10695) );
  MUX2_X1 U10469 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n6601), .Z(n9440) );
  OR2_X1 U10470 ( .A1(n9440), .A2(n9439), .ZN(n9450) );
  XNOR2_X1 U10471 ( .A(n9440), .B(n10673), .ZN(n10678) );
  MUX2_X1 U10472 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n6601), .Z(n9442) );
  OR2_X1 U10473 ( .A1(n9442), .A2(n9441), .ZN(n9449) );
  XNOR2_X1 U10474 ( .A(n9442), .B(n10657), .ZN(n10663) );
  MUX2_X1 U10475 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n6601), .Z(n9447) );
  OR2_X1 U10476 ( .A1(n9447), .A2(n5058), .ZN(n9448) );
  NOR2_X1 U10477 ( .A1(n9444), .A2(n9443), .ZN(n10628) );
  INV_X1 U10478 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9445) );
  MUX2_X1 U10479 ( .A(n9445), .B(n9395), .S(n6601), .Z(n9446) );
  NAND2_X1 U10480 ( .A1(n9446), .A2(n10623), .ZN(n10625) );
  NOR2_X1 U10481 ( .A1(n9446), .A2(n10623), .ZN(n10624) );
  AOI21_X1 U10482 ( .B1(n10628), .B2(n10625), .A(n10624), .ZN(n10644) );
  XNOR2_X1 U10483 ( .A(n9447), .B(n10641), .ZN(n10643) );
  NAND2_X1 U10484 ( .A1(n10644), .A2(n10643), .ZN(n10642) );
  NAND2_X1 U10485 ( .A1(n9448), .A2(n10642), .ZN(n10662) );
  NAND2_X1 U10486 ( .A1(n10663), .A2(n10662), .ZN(n10661) );
  NAND2_X1 U10487 ( .A1(n9449), .A2(n10661), .ZN(n10677) );
  NAND2_X1 U10488 ( .A1(n10678), .A2(n10677), .ZN(n10676) );
  NAND2_X1 U10489 ( .A1(n9450), .A2(n10676), .ZN(n10694) );
  NAND2_X1 U10490 ( .A1(n10695), .A2(n10694), .ZN(n10693) );
  NAND2_X1 U10491 ( .A1(n9451), .A2(n10693), .ZN(n10709) );
  NAND2_X1 U10492 ( .A1(n10710), .A2(n10709), .ZN(n10708) );
  NAND2_X1 U10493 ( .A1(n9452), .A2(n10708), .ZN(n10726) );
  NAND2_X1 U10494 ( .A1(n10727), .A2(n10726), .ZN(n10725) );
  NAND2_X1 U10495 ( .A1(n9453), .A2(n10725), .ZN(n10742) );
  NAND2_X1 U10496 ( .A1(n10743), .A2(n10742), .ZN(n10741) );
  OAI21_X1 U10497 ( .B1(n9455), .B2(n9454), .A(n10741), .ZN(n9457) );
  INV_X1 U10498 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9739) );
  MUX2_X1 U10499 ( .A(n9427), .B(n9739), .S(n6601), .Z(n9456) );
  NOR2_X1 U10500 ( .A1(n9457), .A2(n9456), .ZN(n10762) );
  NAND2_X1 U10501 ( .A1(n9457), .A2(n9456), .ZN(n10763) );
  OAI21_X1 U10502 ( .B1(n10762), .B2(n10771), .A(n10763), .ZN(n9458) );
  XOR2_X1 U10503 ( .A(n9459), .B(n9458), .Z(n9460) );
  NOR2_X1 U10504 ( .A1(n10605), .A2(n9461), .ZN(n9462) );
  AOI211_X1 U10505 ( .C1(n9464), .C2(n10737), .A(n9463), .B(n9462), .ZN(n9465)
         );
  OAI21_X1 U10506 ( .B1(n9470), .B2(n10755), .A(n9469), .ZN(P2_U3201) );
  NAND2_X1 U10507 ( .A1(n9472), .A2(n9471), .ZN(n9782) );
  INV_X1 U10508 ( .A(n9782), .ZN(n9474) );
  NOR2_X1 U10509 ( .A1(n9669), .A2(n9473), .ZN(n9482) );
  NOR3_X1 U10510 ( .A1(n9474), .A2(n9694), .A3(n9482), .ZN(n9477) );
  NOR2_X1 U10511 ( .A1(n9672), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9475) );
  OAI22_X1 U10512 ( .A1(n9784), .A2(n9652), .B1(n9477), .B2(n9475), .ZN(
        P2_U3202) );
  NOR2_X1 U10513 ( .A1(n9672), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9476) );
  OAI22_X1 U10514 ( .A1(n9787), .A2(n9652), .B1(n9477), .B2(n9476), .ZN(
        P2_U3203) );
  INV_X1 U10515 ( .A(n7240), .ZN(n9486) );
  NAND2_X1 U10516 ( .A1(n9672), .A2(n9478), .ZN(n9485) );
  NAND2_X1 U10517 ( .A1(n9479), .A2(n9672), .ZN(n9484) );
  NOR2_X1 U10518 ( .A1(n9480), .A2(n9652), .ZN(n9481) );
  AOI211_X1 U10519 ( .C1(n9694), .C2(P2_REG2_REG_29__SCAN_IN), .A(n9482), .B(
        n9481), .ZN(n9483) );
  OAI211_X1 U10520 ( .C1(n9486), .C2(n9485), .A(n9484), .B(n9483), .ZN(
        P2_U3204) );
  AOI22_X1 U10521 ( .A1(n9694), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n9688), .B2(
        n9487), .ZN(n9488) );
  OAI21_X1 U10522 ( .B1(n9489), .B2(n9652), .A(n9488), .ZN(n9490) );
  AOI21_X1 U10523 ( .B1(n9491), .B2(n9692), .A(n9490), .ZN(n9492) );
  OAI21_X1 U10524 ( .B1(n5000), .B2(n9694), .A(n9492), .ZN(P2_U3205) );
  XNOR2_X1 U10525 ( .A(n9493), .B(n9494), .ZN(n9700) );
  INV_X1 U10526 ( .A(n9700), .ZN(n9504) );
  OAI211_X1 U10527 ( .C1(n9496), .C2(n6590), .A(n7237), .B(n9495), .ZN(n9498)
         );
  NAND2_X1 U10528 ( .A1(n9521), .A2(n9540), .ZN(n9497) );
  OAI211_X1 U10529 ( .C1(n9499), .C2(n9685), .A(n9498), .B(n9497), .ZN(n9699)
         );
  AOI22_X1 U10530 ( .A1(n9694), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n9688), .B2(
        n9500), .ZN(n9501) );
  OAI21_X1 U10531 ( .B1(n9791), .B2(n9652), .A(n9501), .ZN(n9502) );
  AOI21_X1 U10532 ( .B1(n9699), .B2(n9672), .A(n9502), .ZN(n9503) );
  OAI21_X1 U10533 ( .B1(n9504), .B2(n9676), .A(n9503), .ZN(P2_U3206) );
  XOR2_X1 U10534 ( .A(n9505), .B(n9509), .Z(n9507) );
  AOI222_X1 U10535 ( .A1(n7237), .A2(n9507), .B1(n9542), .B2(n9540), .C1(n9506), .C2(n9541), .ZN(n9706) );
  INV_X1 U10536 ( .A(n9508), .ZN(n9512) );
  INV_X1 U10537 ( .A(n9307), .ZN(n9510) );
  OAI22_X1 U10538 ( .A1(n9512), .A2(n9511), .B1(n9510), .B2(n9509), .ZN(n9704)
         );
  AOI22_X1 U10539 ( .A1(n9694), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n9688), .B2(
        n9513), .ZN(n9514) );
  OAI21_X1 U10540 ( .B1(n9515), .B2(n9652), .A(n9514), .ZN(n9516) );
  AOI21_X1 U10541 ( .B1(n9704), .B2(n9692), .A(n9516), .ZN(n9517) );
  OAI21_X1 U10542 ( .B1(n9706), .B2(n9694), .A(n9517), .ZN(P2_U3207) );
  INV_X1 U10543 ( .A(n9518), .ZN(n9796) );
  NOR2_X1 U10544 ( .A1(n9796), .A2(n9678), .ZN(n9525) );
  OAI21_X1 U10545 ( .B1(n9528), .B2(n9520), .A(n9519), .ZN(n9523) );
  AOI222_X1 U10546 ( .A1(n7237), .A2(n9523), .B1(n9522), .B2(n9540), .C1(n9521), .C2(n9541), .ZN(n9524) );
  INV_X1 U10547 ( .A(n9524), .ZN(n9707) );
  AOI211_X1 U10548 ( .C1(n9688), .C2(n9526), .A(n9525), .B(n9707), .ZN(n9530)
         );
  XNOR2_X1 U10549 ( .A(n9527), .B(n9528), .ZN(n9708) );
  AOI22_X1 U10550 ( .A1(n9708), .A2(n9692), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n9694), .ZN(n9529) );
  OAI21_X1 U10551 ( .B1(n9530), .B2(n9694), .A(n9529), .ZN(P2_U3208) );
  AND2_X1 U10552 ( .A1(n9531), .A2(n9771), .ZN(n9713) );
  INV_X1 U10553 ( .A(n9532), .ZN(n9533) );
  NOR2_X1 U10554 ( .A1(n9669), .A2(n9533), .ZN(n9545) );
  NAND2_X1 U10555 ( .A1(n9534), .A2(n9535), .ZN(n9536) );
  NAND2_X1 U10556 ( .A1(n9537), .A2(n9536), .ZN(n9538) );
  NAND2_X1 U10557 ( .A1(n9538), .A2(n7237), .ZN(n9544) );
  AOI22_X1 U10558 ( .A1(n9542), .A2(n9541), .B1(n9540), .B2(n9539), .ZN(n9543)
         );
  NAND2_X1 U10559 ( .A1(n9544), .A2(n9543), .ZN(n9714) );
  AOI211_X1 U10560 ( .C1(n9713), .C2(n9546), .A(n9545), .B(n9714), .ZN(n9551)
         );
  NAND2_X1 U10561 ( .A1(n9548), .A2(n9547), .ZN(n9711) );
  NAND3_X1 U10562 ( .A1(n9712), .A2(n9692), .A3(n9711), .ZN(n9550) );
  NAND2_X1 U10563 ( .A1(n9694), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9549) );
  OAI211_X1 U10564 ( .C1(n9551), .C2(n9694), .A(n9550), .B(n9549), .ZN(
        P2_U3209) );
  XNOR2_X1 U10565 ( .A(n9552), .B(n9555), .ZN(n9553) );
  OAI222_X1 U10566 ( .A1(n9685), .A2(n9554), .B1(n9684), .B2(n9576), .C1(n9553), .C2(n9682), .ZN(n9716) );
  INV_X1 U10567 ( .A(n9716), .ZN(n9561) );
  XNOR2_X1 U10568 ( .A(n9556), .B(n9555), .ZN(n9717) );
  AOI22_X1 U10569 ( .A1(n9694), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n9688), .B2(
        n9557), .ZN(n9558) );
  OAI21_X1 U10570 ( .B1(n9801), .B2(n9652), .A(n9558), .ZN(n9559) );
  AOI21_X1 U10571 ( .B1(n9717), .B2(n9692), .A(n9559), .ZN(n9560) );
  OAI21_X1 U10572 ( .B1(n9561), .B2(n9694), .A(n9560), .ZN(P2_U3210) );
  XNOR2_X1 U10573 ( .A(n9562), .B(n9565), .ZN(n9563) );
  OAI222_X1 U10574 ( .A1(n9685), .A2(n9564), .B1(n9684), .B2(n9592), .C1(n9563), .C2(n9682), .ZN(n9720) );
  INV_X1 U10575 ( .A(n9720), .ZN(n9571) );
  XOR2_X1 U10576 ( .A(n9566), .B(n9565), .Z(n9721) );
  AOI22_X1 U10577 ( .A1(n9694), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9688), .B2(
        n9567), .ZN(n9568) );
  OAI21_X1 U10578 ( .B1(n9805), .B2(n9652), .A(n9568), .ZN(n9569) );
  AOI21_X1 U10579 ( .B1(n9721), .B2(n9692), .A(n9569), .ZN(n9570) );
  OAI21_X1 U10580 ( .B1(n9571), .B2(n9694), .A(n9570), .ZN(P2_U3211) );
  NAND3_X1 U10581 ( .A1(n9588), .A2(n9580), .A3(n9572), .ZN(n9573) );
  AND2_X1 U10582 ( .A1(n9574), .A2(n9573), .ZN(n9575) );
  OAI222_X1 U10583 ( .A1(n9684), .A2(n9603), .B1(n9685), .B2(n9576), .C1(n9682), .C2(n9575), .ZN(n9725) );
  INV_X1 U10584 ( .A(n9577), .ZN(n9809) );
  AOI22_X1 U10585 ( .A1(n9694), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9688), .B2(
        n9578), .ZN(n9579) );
  OAI21_X1 U10586 ( .B1(n9809), .B2(n9652), .A(n9579), .ZN(n9585) );
  NOR2_X1 U10587 ( .A1(n9581), .A2(n9580), .ZN(n9724) );
  INV_X1 U10588 ( .A(n9582), .ZN(n9583) );
  NOR3_X1 U10589 ( .A1(n9724), .A2(n9583), .A3(n9676), .ZN(n9584) );
  AOI211_X1 U10590 ( .C1(n9725), .C2(n9672), .A(n9585), .B(n9584), .ZN(n9586)
         );
  INV_X1 U10591 ( .A(n9586), .ZN(P2_U3212) );
  INV_X1 U10592 ( .A(n9587), .ZN(n9590) );
  INV_X1 U10593 ( .A(n9588), .ZN(n9589) );
  AOI21_X1 U10594 ( .B1(n9590), .B2(n5366), .A(n9589), .ZN(n9591) );
  OAI222_X1 U10595 ( .A1(n9685), .A2(n9592), .B1(n9684), .B2(n9613), .C1(n9682), .C2(n9591), .ZN(n9729) );
  INV_X1 U10596 ( .A(n9729), .ZN(n9599) );
  XNOR2_X1 U10597 ( .A(n9593), .B(n5366), .ZN(n9730) );
  INV_X1 U10598 ( .A(n9594), .ZN(n9813) );
  AOI22_X1 U10599 ( .A1(n9694), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9688), .B2(
        n9595), .ZN(n9596) );
  OAI21_X1 U10600 ( .B1(n9813), .B2(n9652), .A(n9596), .ZN(n9597) );
  AOI21_X1 U10601 ( .B1(n9730), .B2(n9692), .A(n9597), .ZN(n9598) );
  OAI21_X1 U10602 ( .B1(n9599), .B2(n9694), .A(n9598), .ZN(P2_U3213) );
  XNOR2_X1 U10603 ( .A(n9601), .B(n9600), .ZN(n9602) );
  OAI222_X1 U10604 ( .A1(n9685), .A2(n9603), .B1(n9684), .B2(n9623), .C1(n9602), .C2(n9682), .ZN(n9733) );
  INV_X1 U10605 ( .A(n9733), .ZN(n9610) );
  XNOR2_X1 U10606 ( .A(n9604), .B(n9605), .ZN(n9734) );
  AOI22_X1 U10607 ( .A1(n9694), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n9688), .B2(
        n9606), .ZN(n9607) );
  OAI21_X1 U10608 ( .B1(n9817), .B2(n9652), .A(n9607), .ZN(n9608) );
  AOI21_X1 U10609 ( .B1(n9734), .B2(n9692), .A(n9608), .ZN(n9609) );
  OAI21_X1 U10610 ( .B1(n9610), .B2(n9694), .A(n9609), .ZN(P2_U3214) );
  XOR2_X1 U10611 ( .A(n9611), .B(n9615), .Z(n9612) );
  OAI222_X1 U10612 ( .A1(n9685), .A2(n9613), .B1(n9684), .B2(n9636), .C1(n9612), .C2(n9682), .ZN(n9737) );
  INV_X1 U10613 ( .A(n9737), .ZN(n9620) );
  XOR2_X1 U10614 ( .A(n9614), .B(n9615), .Z(n9738) );
  AOI22_X1 U10615 ( .A1(n9694), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9688), .B2(
        n9616), .ZN(n9617) );
  OAI21_X1 U10616 ( .B1(n9821), .B2(n9652), .A(n9617), .ZN(n9618) );
  AOI21_X1 U10617 ( .B1(n9738), .B2(n9692), .A(n9618), .ZN(n9619) );
  OAI21_X1 U10618 ( .B1(n9620), .B2(n9694), .A(n9619), .ZN(P2_U3215) );
  XNOR2_X1 U10619 ( .A(n9621), .B(n9624), .ZN(n9622) );
  OAI222_X1 U10620 ( .A1(n9685), .A2(n9623), .B1(n9684), .B2(n9648), .C1(n9682), .C2(n9622), .ZN(n9741) );
  NAND2_X1 U10621 ( .A1(n9625), .A2(n9624), .ZN(n9626) );
  AND2_X1 U10622 ( .A1(n9627), .A2(n9626), .ZN(n9742) );
  NAND2_X1 U10623 ( .A1(n9742), .A2(n9692), .ZN(n9630) );
  AOI22_X1 U10624 ( .A1(n9694), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n9688), .B2(
        n9628), .ZN(n9629) );
  OAI211_X1 U10625 ( .C1(n9825), .C2(n9652), .A(n9630), .B(n9629), .ZN(n9631)
         );
  AOI21_X1 U10626 ( .B1(n9741), .B2(n9672), .A(n9631), .ZN(n9632) );
  INV_X1 U10627 ( .A(n9632), .ZN(P2_U3216) );
  XNOR2_X1 U10628 ( .A(n9633), .B(n9634), .ZN(n9635) );
  OAI222_X1 U10629 ( .A1(n9685), .A2(n9636), .B1(n9684), .B2(n9667), .C1(n9635), .C2(n9682), .ZN(n9745) );
  INV_X1 U10630 ( .A(n9745), .ZN(n9645) );
  OAI21_X1 U10631 ( .B1(n9639), .B2(n9638), .A(n9637), .ZN(n9746) );
  INV_X1 U10632 ( .A(n9640), .ZN(n9829) );
  AOI22_X1 U10633 ( .A1(n9694), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n9688), .B2(
        n9641), .ZN(n9642) );
  OAI21_X1 U10634 ( .B1(n9829), .B2(n9652), .A(n9642), .ZN(n9643) );
  AOI21_X1 U10635 ( .B1(n9746), .B2(n9692), .A(n9643), .ZN(n9644) );
  OAI21_X1 U10636 ( .B1(n9645), .B2(n9694), .A(n9644), .ZN(P2_U3217) );
  XNOR2_X1 U10637 ( .A(n4956), .B(n9649), .ZN(n9647) );
  OAI222_X1 U10638 ( .A1(n9685), .A2(n9648), .B1(n9684), .B2(n8943), .C1(n9647), .C2(n9682), .ZN(n9749) );
  INV_X1 U10639 ( .A(n9749), .ZN(n9658) );
  INV_X1 U10640 ( .A(n9649), .ZN(n9651) );
  OAI21_X1 U10641 ( .B1(n5032), .B2(n9651), .A(n9650), .ZN(n9750) );
  NOR2_X1 U10642 ( .A1(n9834), .A2(n9652), .ZN(n9656) );
  INV_X1 U10643 ( .A(n9653), .ZN(n9654) );
  OAI22_X1 U10644 ( .A1(n9672), .A2(n10714), .B1(n9654), .B2(n9669), .ZN(n9655) );
  AOI211_X1 U10645 ( .C1(n9750), .C2(n9692), .A(n9656), .B(n9655), .ZN(n9657)
         );
  OAI21_X1 U10646 ( .B1(n9658), .B2(n9694), .A(n9657), .ZN(P2_U3218) );
  INV_X1 U10647 ( .A(n9659), .ZN(n9662) );
  INV_X1 U10648 ( .A(n9664), .ZN(n9661) );
  OAI21_X1 U10649 ( .B1(n9662), .B2(n9661), .A(n9660), .ZN(n9754) );
  XNOR2_X1 U10650 ( .A(n9663), .B(n9664), .ZN(n9665) );
  OAI222_X1 U10651 ( .A1(n9685), .A2(n9667), .B1(n9684), .B2(n9666), .C1(n9682), .C2(n9665), .ZN(n9755) );
  INV_X1 U10652 ( .A(n9757), .ZN(n9671) );
  INV_X1 U10653 ( .A(n9668), .ZN(n9670) );
  OAI22_X1 U10654 ( .A1(n9671), .A2(n9678), .B1(n9670), .B2(n9669), .ZN(n9673)
         );
  OAI21_X1 U10655 ( .B1(n9755), .B2(n9673), .A(n9672), .ZN(n9675) );
  NAND2_X1 U10656 ( .A1(n9694), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n9674) );
  OAI211_X1 U10657 ( .C1(n9754), .C2(n9676), .A(n9675), .B(n9674), .ZN(
        P2_U3219) );
  INV_X1 U10658 ( .A(n9677), .ZN(n9760) );
  NOR2_X1 U10659 ( .A1(n9760), .A2(n9678), .ZN(n9686) );
  XNOR2_X1 U10660 ( .A(n9680), .B(n9679), .ZN(n9681) );
  OAI222_X1 U10661 ( .A1(n9685), .A2(n8943), .B1(n9684), .B2(n9683), .C1(n9682), .C2(n9681), .ZN(n9761) );
  AOI211_X1 U10662 ( .C1(n9688), .C2(n9687), .A(n9686), .B(n9761), .ZN(n9695)
         );
  OAI21_X1 U10663 ( .B1(n9691), .B2(n9690), .A(n9689), .ZN(n9763) );
  AOI22_X1 U10664 ( .A1(n9763), .A2(n9692), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n9694), .ZN(n9693) );
  OAI21_X1 U10665 ( .B1(n9695), .B2(n9694), .A(n9693), .ZN(P2_U3220) );
  NOR2_X1 U10666 ( .A1(n9782), .A2(n7250), .ZN(n9697) );
  AOI21_X1 U10667 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n7250), .A(n9697), .ZN(
        n9696) );
  OAI21_X1 U10668 ( .B1(n9784), .B2(n9753), .A(n9696), .ZN(P2_U3490) );
  AOI21_X1 U10669 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n7250), .A(n9697), .ZN(
        n9698) );
  OAI21_X1 U10670 ( .B1(n9787), .B2(n9753), .A(n9698), .ZN(P2_U3489) );
  INV_X1 U10671 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9701) );
  AOI21_X1 U10672 ( .B1(n9700), .B2(n9778), .A(n9699), .ZN(n9788) );
  MUX2_X1 U10673 ( .A(n9701), .B(n9788), .S(n9781), .Z(n9702) );
  OAI21_X1 U10674 ( .B1(n9791), .B2(n9753), .A(n9702), .ZN(P2_U3486) );
  AOI22_X1 U10675 ( .A1(n9704), .A2(n9778), .B1(n9771), .B2(n9703), .ZN(n9705)
         );
  NAND2_X1 U10676 ( .A1(n9706), .A2(n9705), .ZN(n9792) );
  MUX2_X1 U10677 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9792), .S(n9781), .Z(
        P2_U3485) );
  INV_X1 U10678 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9709) );
  AOI21_X1 U10679 ( .B1(n9708), .B2(n9778), .A(n9707), .ZN(n9793) );
  MUX2_X1 U10680 ( .A(n9709), .B(n9793), .S(n9781), .Z(n9710) );
  OAI21_X1 U10681 ( .B1(n9796), .B2(n9753), .A(n9710), .ZN(P2_U3484) );
  AND3_X1 U10682 ( .A1(n9712), .A2(n9711), .A3(n9778), .ZN(n9715) );
  MUX2_X1 U10683 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9797), .S(n9781), .Z(
        P2_U3483) );
  INV_X1 U10684 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9718) );
  AOI21_X1 U10685 ( .B1(n9778), .B2(n9717), .A(n9716), .ZN(n9798) );
  MUX2_X1 U10686 ( .A(n9718), .B(n9798), .S(n9781), .Z(n9719) );
  OAI21_X1 U10687 ( .B1(n9801), .B2(n9753), .A(n9719), .ZN(P2_U3482) );
  INV_X1 U10688 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9722) );
  AOI21_X1 U10689 ( .B1(n9721), .B2(n9778), .A(n9720), .ZN(n9802) );
  MUX2_X1 U10690 ( .A(n9722), .B(n9802), .S(n9781), .Z(n9723) );
  OAI21_X1 U10691 ( .B1(n9805), .B2(n9753), .A(n9723), .ZN(P2_U3481) );
  INV_X1 U10692 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9727) );
  NOR2_X1 U10693 ( .A1(n9724), .A2(n9766), .ZN(n9726) );
  AOI21_X1 U10694 ( .B1(n9726), .B2(n9582), .A(n9725), .ZN(n9806) );
  MUX2_X1 U10695 ( .A(n9727), .B(n9806), .S(n9781), .Z(n9728) );
  OAI21_X1 U10696 ( .B1(n9809), .B2(n9753), .A(n9728), .ZN(P2_U3480) );
  INV_X1 U10697 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9731) );
  AOI21_X1 U10698 ( .B1(n9730), .B2(n9778), .A(n9729), .ZN(n9810) );
  MUX2_X1 U10699 ( .A(n9731), .B(n9810), .S(n9781), .Z(n9732) );
  OAI21_X1 U10700 ( .B1(n9813), .B2(n9753), .A(n9732), .ZN(P2_U3479) );
  INV_X1 U10701 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9735) );
  AOI21_X1 U10702 ( .B1(n9734), .B2(n9778), .A(n9733), .ZN(n9814) );
  MUX2_X1 U10703 ( .A(n9735), .B(n9814), .S(n9781), .Z(n9736) );
  OAI21_X1 U10704 ( .B1(n9817), .B2(n9753), .A(n9736), .ZN(P2_U3478) );
  AOI21_X1 U10705 ( .B1(n9778), .B2(n9738), .A(n9737), .ZN(n9818) );
  MUX2_X1 U10706 ( .A(n9739), .B(n9818), .S(n9781), .Z(n9740) );
  OAI21_X1 U10707 ( .B1(n9821), .B2(n9753), .A(n9740), .ZN(P2_U3477) );
  INV_X1 U10708 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9743) );
  AOI21_X1 U10709 ( .B1(n9742), .B2(n9778), .A(n9741), .ZN(n9822) );
  MUX2_X1 U10710 ( .A(n9743), .B(n9822), .S(n9781), .Z(n9744) );
  OAI21_X1 U10711 ( .B1(n9825), .B2(n9753), .A(n9744), .ZN(P2_U3476) );
  AOI21_X1 U10712 ( .B1(n9778), .B2(n9746), .A(n9745), .ZN(n9826) );
  MUX2_X1 U10713 ( .A(n9747), .B(n9826), .S(n9781), .Z(n9748) );
  OAI21_X1 U10714 ( .B1(n9829), .B2(n9753), .A(n9748), .ZN(P2_U3475) );
  INV_X1 U10715 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9751) );
  AOI21_X1 U10716 ( .B1(n9778), .B2(n9750), .A(n9749), .ZN(n9830) );
  MUX2_X1 U10717 ( .A(n9751), .B(n9830), .S(n9781), .Z(n9752) );
  OAI21_X1 U10718 ( .B1(n9834), .B2(n9753), .A(n9752), .ZN(P2_U3474) );
  NOR2_X1 U10719 ( .A1(n9754), .A2(n9766), .ZN(n9756) );
  AOI211_X1 U10720 ( .C1(n9771), .C2(n9757), .A(n9756), .B(n9755), .ZN(n10850)
         );
  OR2_X1 U10721 ( .A1(n10850), .A2(n7250), .ZN(n9758) );
  OAI21_X1 U10722 ( .B1(n9781), .B2(n9759), .A(n9758), .ZN(P2_U3473) );
  INV_X1 U10723 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9765) );
  NOR2_X1 U10724 ( .A1(n9760), .A2(n9773), .ZN(n9762) );
  AOI211_X1 U10725 ( .C1(n9778), .C2(n9763), .A(n9762), .B(n9761), .ZN(n10848)
         );
  OR2_X1 U10726 ( .A1(n10848), .A2(n7250), .ZN(n9764) );
  OAI21_X1 U10727 ( .B1(n9781), .B2(n9765), .A(n9764), .ZN(P2_U3472) );
  NOR2_X1 U10728 ( .A1(n9767), .A2(n9766), .ZN(n9769) );
  AOI211_X1 U10729 ( .C1(n9771), .C2(n9770), .A(n9769), .B(n9768), .ZN(n10832)
         );
  NAND2_X1 U10730 ( .A1(n7250), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n9772) );
  OAI21_X1 U10731 ( .B1(n10832), .B2(n7250), .A(n9772), .ZN(P2_U3471) );
  INV_X1 U10732 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9780) );
  NOR2_X1 U10733 ( .A1(n9774), .A2(n9773), .ZN(n9776) );
  AOI211_X1 U10734 ( .C1(n9778), .C2(n9777), .A(n9776), .B(n9775), .ZN(n10830)
         );
  OR2_X1 U10735 ( .A1(n10830), .A2(n7250), .ZN(n9779) );
  OAI21_X1 U10736 ( .B1(n9781), .B2(n9780), .A(n9779), .ZN(P2_U3470) );
  NOR2_X1 U10737 ( .A1(n7244), .A2(n9782), .ZN(n9785) );
  AOI21_X1 U10738 ( .B1(P2_REG0_REG_31__SCAN_IN), .B2(n7244), .A(n9785), .ZN(
        n9783) );
  OAI21_X1 U10739 ( .B1(n9784), .B2(n9833), .A(n9783), .ZN(P2_U3458) );
  AOI21_X1 U10740 ( .B1(P2_REG0_REG_30__SCAN_IN), .B2(n7244), .A(n9785), .ZN(
        n9786) );
  OAI21_X1 U10741 ( .B1(n9787), .B2(n9833), .A(n9786), .ZN(P2_U3457) );
  INV_X1 U10742 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9789) );
  MUX2_X1 U10743 ( .A(n9789), .B(n9788), .S(n10851), .Z(n9790) );
  OAI21_X1 U10744 ( .B1(n9791), .B2(n9833), .A(n9790), .ZN(P2_U3454) );
  MUX2_X1 U10745 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9792), .S(n10851), .Z(
        P2_U3453) );
  INV_X1 U10746 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9794) );
  MUX2_X1 U10747 ( .A(n9794), .B(n9793), .S(n10851), .Z(n9795) );
  OAI21_X1 U10748 ( .B1(n9796), .B2(n9833), .A(n9795), .ZN(P2_U3452) );
  MUX2_X1 U10749 ( .A(n9797), .B(P2_REG0_REG_24__SCAN_IN), .S(n7244), .Z(
        P2_U3451) );
  INV_X1 U10750 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9799) );
  MUX2_X1 U10751 ( .A(n9799), .B(n9798), .S(n10851), .Z(n9800) );
  OAI21_X1 U10752 ( .B1(n9801), .B2(n9833), .A(n9800), .ZN(P2_U3450) );
  INV_X1 U10753 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9803) );
  MUX2_X1 U10754 ( .A(n9803), .B(n9802), .S(n10851), .Z(n9804) );
  OAI21_X1 U10755 ( .B1(n9805), .B2(n9833), .A(n9804), .ZN(P2_U3449) );
  INV_X1 U10756 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9807) );
  MUX2_X1 U10757 ( .A(n9807), .B(n9806), .S(n10851), .Z(n9808) );
  OAI21_X1 U10758 ( .B1(n9809), .B2(n9833), .A(n9808), .ZN(P2_U3448) );
  INV_X1 U10759 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9811) );
  MUX2_X1 U10760 ( .A(n9811), .B(n9810), .S(n10851), .Z(n9812) );
  OAI21_X1 U10761 ( .B1(n9813), .B2(n9833), .A(n9812), .ZN(P2_U3447) );
  INV_X1 U10762 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9815) );
  MUX2_X1 U10763 ( .A(n9815), .B(n9814), .S(n10851), .Z(n9816) );
  OAI21_X1 U10764 ( .B1(n9817), .B2(n9833), .A(n9816), .ZN(P2_U3446) );
  INV_X1 U10765 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9819) );
  MUX2_X1 U10766 ( .A(n9819), .B(n9818), .S(n10851), .Z(n9820) );
  OAI21_X1 U10767 ( .B1(n9821), .B2(n9833), .A(n9820), .ZN(P2_U3444) );
  INV_X1 U10768 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9823) );
  MUX2_X1 U10769 ( .A(n9823), .B(n9822), .S(n10851), .Z(n9824) );
  OAI21_X1 U10770 ( .B1(n9825), .B2(n9833), .A(n9824), .ZN(P2_U3441) );
  INV_X1 U10771 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9827) );
  MUX2_X1 U10772 ( .A(n9827), .B(n9826), .S(n10851), .Z(n9828) );
  OAI21_X1 U10773 ( .B1(n9829), .B2(n9833), .A(n9828), .ZN(P2_U3438) );
  INV_X1 U10774 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9831) );
  MUX2_X1 U10775 ( .A(n9831), .B(n9830), .S(n10851), .Z(n9832) );
  OAI21_X1 U10776 ( .B1(n9834), .B2(n9833), .A(n9832), .ZN(P2_U3435) );
  INV_X1 U10777 ( .A(n9835), .ZN(n10479) );
  NOR4_X1 U10778 ( .A1(n6229), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n6352), .ZN(n9836) );
  AOI21_X1 U10779 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n9846), .A(n9836), .ZN(
        n9837) );
  OAI21_X1 U10780 ( .B1(n10479), .B2(n9856), .A(n9837), .ZN(P2_U3264) );
  AOI22_X1 U10781 ( .A1(n9838), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9846), .ZN(n9839) );
  OAI21_X1 U10782 ( .B1(n9840), .B2(n9856), .A(n9839), .ZN(P2_U3265) );
  INV_X1 U10783 ( .A(n9841), .ZN(n10480) );
  AOI22_X1 U10784 ( .A1(n9842), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n9846), .ZN(n9843) );
  OAI21_X1 U10785 ( .B1(n10480), .B2(n9856), .A(n9843), .ZN(P2_U3266) );
  INV_X1 U10786 ( .A(n9844), .ZN(n10484) );
  AOI21_X1 U10787 ( .B1(n9846), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n9845), .ZN(
        n9847) );
  OAI21_X1 U10788 ( .B1(n10484), .B2(n9856), .A(n9847), .ZN(P2_U3267) );
  NAND2_X1 U10789 ( .A1(n10486), .A2(n9848), .ZN(n9851) );
  INV_X1 U10790 ( .A(n9849), .ZN(n9850) );
  OAI211_X1 U10791 ( .C1(n9852), .C2(n9855), .A(n9851), .B(n9850), .ZN(
        P2_U3268) );
  INV_X1 U10792 ( .A(n9853), .ZN(n10491) );
  OAI222_X1 U10793 ( .A1(P2_U3151), .A2(n5156), .B1(n9856), .B2(n10491), .C1(
        n9855), .C2(n9854), .ZN(P2_U3269) );
  MUX2_X1 U10794 ( .A(n9857), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  NAND2_X1 U10795 ( .A1(n9858), .A2(n9859), .ZN(n9860) );
  XOR2_X1 U10796 ( .A(n9861), .B(n9860), .Z(n9868) );
  AOI21_X1 U10797 ( .B1(n10003), .B2(n10034), .A(n9862), .ZN(n9865) );
  NAND2_X1 U10798 ( .A1(n10015), .A2(n9863), .ZN(n9864) );
  OAI211_X1 U10799 ( .C1(n9925), .C2(n9991), .A(n9865), .B(n9864), .ZN(n9866)
         );
  AOI21_X1 U10800 ( .B1(n10427), .B2(n10023), .A(n9866), .ZN(n9867) );
  OAI21_X1 U10801 ( .B1(n9868), .B2(n10026), .A(n9867), .ZN(P1_U3215) );
  OR2_X1 U10802 ( .A1(n9870), .A2(n9869), .ZN(n9978) );
  NAND2_X1 U10803 ( .A1(n9978), .A2(n9977), .ZN(n9976) );
  NAND2_X1 U10804 ( .A1(n9870), .A2(n9869), .ZN(n9980) );
  NAND2_X1 U10805 ( .A1(n9871), .A2(n9941), .ZN(n9872) );
  AOI21_X1 U10806 ( .B1(n9976), .B2(n9980), .A(n9872), .ZN(n9944) );
  AND3_X1 U10807 ( .A1(n9976), .A2(n9980), .A3(n9872), .ZN(n9873) );
  OAI21_X1 U10808 ( .B1(n9944), .B2(n9873), .A(n10002), .ZN(n9878) );
  NOR2_X1 U10809 ( .A1(n10005), .A2(n10227), .ZN(n9876) );
  OAI22_X1 U10810 ( .A1(n10222), .A2(n9991), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9874), .ZN(n9875) );
  AOI211_X1 U10811 ( .C1(n10003), .C2(n10254), .A(n9876), .B(n9875), .ZN(n9877) );
  OAI211_X1 U10812 ( .C1(n10455), .C2(n10009), .A(n9878), .B(n9877), .ZN(
        P1_U3216) );
  INV_X1 U10813 ( .A(n9879), .ZN(n9957) );
  AOI21_X1 U10814 ( .B1(n9881), .B2(n9880), .A(n9957), .ZN(n9886) );
  NAND2_X1 U10815 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n10115)
         );
  OAI21_X1 U10816 ( .B1(n9991), .B2(n10302), .A(n10115), .ZN(n9882) );
  AOI21_X1 U10817 ( .B1(n10003), .B2(n10031), .A(n9882), .ZN(n9883) );
  OAI21_X1 U10818 ( .B1(n10005), .B2(n10290), .A(n9883), .ZN(n9884) );
  AOI21_X1 U10819 ( .B1(n10296), .B2(n10023), .A(n9884), .ZN(n9885) );
  OAI21_X1 U10820 ( .B1(n9886), .B2(n10026), .A(n9885), .ZN(P1_U3219) );
  INV_X1 U10821 ( .A(n10390), .ZN(n10263) );
  OAI21_X1 U10822 ( .B1(n9889), .B2(n9888), .A(n9887), .ZN(n9890) );
  NAND2_X1 U10823 ( .A1(n9890), .A2(n10002), .ZN(n9895) );
  OAI22_X1 U10824 ( .A1(n9991), .A2(n10377), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9891), .ZN(n9893) );
  NOR2_X1 U10825 ( .A1(n10005), .A2(n10258), .ZN(n9892) );
  AOI211_X1 U10826 ( .C1(n10003), .C2(n10388), .A(n9893), .B(n9892), .ZN(n9894) );
  OAI211_X1 U10827 ( .C1(n10263), .C2(n10009), .A(n9895), .B(n9894), .ZN(
        P1_U3223) );
  INV_X1 U10828 ( .A(n9896), .ZN(n9897) );
  AOI21_X1 U10829 ( .B1(n9899), .B2(n9898), .A(n9897), .ZN(n9908) );
  AOI21_X1 U10830 ( .B1(n10003), .B2(n10036), .A(n9900), .ZN(n9903) );
  NAND2_X1 U10831 ( .A1(n10015), .A2(n9901), .ZN(n9902) );
  OAI211_X1 U10832 ( .C1(n9904), .C2(n9991), .A(n9903), .B(n9902), .ZN(n9905)
         );
  AOI21_X1 U10833 ( .B1(n9906), .B2(n10023), .A(n9905), .ZN(n9907) );
  OAI21_X1 U10834 ( .B1(n9908), .B2(n10026), .A(n9907), .ZN(P1_U3224) );
  AOI21_X1 U10835 ( .B1(n9910), .B2(n9909), .A(n10000), .ZN(n9916) );
  OAI22_X1 U10836 ( .A1(n10208), .A2(n9991), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9911), .ZN(n9912) );
  AOI21_X1 U10837 ( .B1(n10003), .B2(n10205), .A(n9912), .ZN(n9913) );
  OAI21_X1 U10838 ( .B1(n10005), .B2(n10212), .A(n9913), .ZN(n9914) );
  AOI21_X1 U10839 ( .B1(n4961), .B2(n10023), .A(n9914), .ZN(n9915) );
  OAI21_X1 U10840 ( .B1(n9916), .B2(n10026), .A(n9915), .ZN(P1_U3225) );
  INV_X1 U10841 ( .A(n9917), .ZN(n9918) );
  AOI21_X1 U10842 ( .B1(n9920), .B2(n9919), .A(n9918), .ZN(n9928) );
  NAND2_X1 U10843 ( .A1(n10015), .A2(n9921), .ZN(n9924) );
  AOI21_X1 U10844 ( .B1(n10017), .B2(n9993), .A(n9922), .ZN(n9923) );
  OAI211_X1 U10845 ( .C1(n9925), .C2(n10020), .A(n9924), .B(n9923), .ZN(n9926)
         );
  AOI21_X1 U10846 ( .B1(n10422), .B2(n10023), .A(n9926), .ZN(n9927) );
  OAI21_X1 U10847 ( .B1(n9928), .B2(n10026), .A(n9927), .ZN(P1_U3226) );
  XNOR2_X1 U10848 ( .A(n9930), .B(n9929), .ZN(n9931) );
  XNOR2_X1 U10849 ( .A(n9932), .B(n9931), .ZN(n9940) );
  NAND2_X1 U10850 ( .A1(n10017), .A2(n10031), .ZN(n9934) );
  OAI211_X1 U10851 ( .C1(n10020), .C2(n9935), .A(n9934), .B(n9933), .ZN(n9937)
         );
  NOR2_X1 U10852 ( .A1(n10470), .A2(n10009), .ZN(n9936) );
  AOI211_X1 U10853 ( .C1(n9938), .C2(n10015), .A(n9937), .B(n9936), .ZN(n9939)
         );
  OAI21_X1 U10854 ( .B1(n9940), .B2(n10026), .A(n9939), .ZN(P1_U3228) );
  INV_X1 U10855 ( .A(n9941), .ZN(n9943) );
  NOR3_X1 U10856 ( .A1(n9944), .A2(n9943), .A3(n9942), .ZN(n9946) );
  OAI21_X1 U10857 ( .B1(n9946), .B2(n9945), .A(n10002), .ZN(n9952) );
  AOI22_X1 U10858 ( .A1(n10030), .A2(n10017), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9947) );
  OAI21_X1 U10859 ( .B1(n9948), .B2(n10020), .A(n9947), .ZN(n9949) );
  AOI21_X1 U10860 ( .B1(n9950), .B2(n10015), .A(n9949), .ZN(n9951) );
  OAI211_X1 U10861 ( .C1(n9953), .C2(n10009), .A(n9952), .B(n9951), .ZN(
        P1_U3229) );
  INV_X1 U10862 ( .A(n10273), .ZN(n10397) );
  INV_X1 U10863 ( .A(n9954), .ZN(n9956) );
  NOR3_X1 U10864 ( .A1(n9957), .A2(n9956), .A3(n9955), .ZN(n9960) );
  INV_X1 U10865 ( .A(n9958), .ZN(n9959) );
  OAI21_X1 U10866 ( .B1(n9960), .B2(n9959), .A(n10002), .ZN(n9964) );
  AOI22_X1 U10867 ( .A1(n10281), .A2(n10017), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9961) );
  OAI21_X1 U10868 ( .B1(n10396), .B2(n10020), .A(n9961), .ZN(n9962) );
  AOI21_X1 U10869 ( .B1(n10275), .B2(n10015), .A(n9962), .ZN(n9963) );
  OAI211_X1 U10870 ( .C1(n10397), .C2(n10009), .A(n9964), .B(n9963), .ZN(
        P1_U3233) );
  AOI21_X1 U10871 ( .B1(n9966), .B2(n9965), .A(n10026), .ZN(n9968) );
  NAND2_X1 U10872 ( .A1(n9968), .A2(n9967), .ZN(n9974) );
  AOI21_X1 U10873 ( .B1(n10003), .B2(n10035), .A(n9969), .ZN(n9970) );
  OAI21_X1 U10874 ( .B1(n10021), .B2(n9991), .A(n9970), .ZN(n9971) );
  AOI21_X1 U10875 ( .B1(n9972), .B2(n10015), .A(n9971), .ZN(n9973) );
  OAI211_X1 U10876 ( .C1(n9975), .C2(n10009), .A(n9974), .B(n9973), .ZN(
        P1_U3234) );
  INV_X1 U10877 ( .A(n9976), .ZN(n9981) );
  AOI21_X1 U10878 ( .B1(n9978), .B2(n9980), .A(n9977), .ZN(n9979) );
  AOI21_X1 U10879 ( .B1(n9981), .B2(n9980), .A(n9979), .ZN(n9986) );
  AOI22_X1 U10880 ( .A1(n10245), .A2(n10017), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9983) );
  NAND2_X1 U10881 ( .A1(n10003), .A2(n10281), .ZN(n9982) );
  OAI211_X1 U10882 ( .C1(n10005), .C2(n10240), .A(n9983), .B(n9982), .ZN(n9984) );
  AOI21_X1 U10883 ( .B1(n10383), .B2(n10023), .A(n9984), .ZN(n9985) );
  OAI21_X1 U10884 ( .B1(n9986), .B2(n10026), .A(n9985), .ZN(P1_U3235) );
  XOR2_X1 U10885 ( .A(n9988), .B(n9987), .Z(n9989) );
  XNOR2_X1 U10886 ( .A(n9990), .B(n9989), .ZN(n9997) );
  NAND2_X1 U10887 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10094)
         );
  OAI21_X1 U10888 ( .B1(n9991), .B2(n10396), .A(n10094), .ZN(n9992) );
  AOI21_X1 U10889 ( .B1(n10003), .B2(n9993), .A(n9992), .ZN(n9994) );
  OAI21_X1 U10890 ( .B1(n10005), .B2(n10327), .A(n9994), .ZN(n9995) );
  AOI21_X1 U10891 ( .B1(n10324), .B2(n10023), .A(n9995), .ZN(n9996) );
  OAI21_X1 U10892 ( .B1(n9997), .B2(n10026), .A(n9996), .ZN(P1_U3238) );
  OAI21_X1 U10893 ( .B1(n10000), .B2(n9999), .A(n9998), .ZN(n10001) );
  NAND3_X1 U10894 ( .A1(n5016), .A2(n10002), .A3(n10001), .ZN(n10008) );
  AOI22_X1 U10895 ( .A1(n10030), .A2(n10003), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10004) );
  OAI21_X1 U10896 ( .B1(n10005), .B2(n10192), .A(n10004), .ZN(n10006) );
  AOI21_X1 U10897 ( .B1(n10017), .B2(n10188), .A(n10006), .ZN(n10007) );
  OAI211_X1 U10898 ( .C1(n5242), .C2(n10009), .A(n10008), .B(n10007), .ZN(
        P1_U3240) );
  NAND2_X1 U10899 ( .A1(n10010), .A2(n10011), .ZN(n10012) );
  XOR2_X1 U10900 ( .A(n10013), .B(n10012), .Z(n10027) );
  NAND2_X1 U10901 ( .A1(n10015), .A2(n10014), .ZN(n10019) );
  AOI21_X1 U10902 ( .B1(n10017), .B2(n10032), .A(n10016), .ZN(n10018) );
  OAI211_X1 U10903 ( .C1(n10021), .C2(n10020), .A(n10019), .B(n10018), .ZN(
        n10022) );
  AOI21_X1 U10904 ( .B1(n10024), .B2(n10023), .A(n10022), .ZN(n10025) );
  OAI21_X1 U10905 ( .B1(n10027), .B2(n10026), .A(n10025), .ZN(P1_U3241) );
  MUX2_X1 U10906 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n10028), .S(n10852), .Z(
        P1_U3585) );
  MUX2_X1 U10907 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n10138), .S(n10852), .Z(
        P1_U3584) );
  MUX2_X1 U10908 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n10029), .S(n10852), .Z(
        P1_U3583) );
  MUX2_X1 U10909 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n10345), .S(n10852), .Z(
        P1_U3582) );
  MUX2_X1 U10910 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n10030), .S(n10852), .Z(
        P1_U3579) );
  MUX2_X1 U10911 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n10205), .S(n10852), .Z(
        P1_U3578) );
  MUX2_X1 U10912 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n10245), .S(n10852), .Z(
        P1_U3577) );
  MUX2_X1 U10913 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n10254), .S(n10852), .Z(
        P1_U3576) );
  MUX2_X1 U10914 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n10281), .S(n10852), .Z(
        P1_U3575) );
  MUX2_X1 U10915 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n10031), .S(n10852), .Z(
        P1_U3572) );
  MUX2_X1 U10916 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n10032), .S(n10852), .Z(
        P1_U3570) );
  MUX2_X1 U10917 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n10033), .S(n10852), .Z(
        P1_U3569) );
  MUX2_X1 U10918 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n10034), .S(n10852), .Z(
        P1_U3567) );
  MUX2_X1 U10919 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n10035), .S(n10852), .Z(
        P1_U3566) );
  MUX2_X1 U10920 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n10036), .S(n10852), .Z(
        P1_U3565) );
  MUX2_X1 U10921 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n10037), .S(n10852), .Z(
        P1_U3564) );
  MUX2_X1 U10922 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n10038), .S(n10852), .Z(
        P1_U3561) );
  MUX2_X1 U10923 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n10039), .S(n10852), .Z(
        P1_U3560) );
  MUX2_X1 U10924 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n10040), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10925 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n10041), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10926 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n10042), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10927 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n10043), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10928 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n10044), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U10929 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6960), .S(P1_U3973), .Z(
        P1_U3554) );
  OAI211_X1 U10930 ( .C1(n10047), .C2(n10046), .A(n10072), .B(n10045), .ZN(
        n10055) );
  OAI211_X1 U10931 ( .C1(n10050), .C2(n10049), .A(n10120), .B(n10048), .ZN(
        n10054) );
  AOI22_X1 U10932 ( .A1(n10560), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n10053) );
  NAND2_X1 U10933 ( .A1(n10076), .A2(n10051), .ZN(n10052) );
  NAND4_X1 U10934 ( .A1(n10055), .A2(n10054), .A3(n10053), .A4(n10052), .ZN(
        P1_U3244) );
  NOR2_X1 U10935 ( .A1(n10117), .A2(n10061), .ZN(n10056) );
  AOI211_X1 U10936 ( .C1(n10560), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n10057), .B(
        n10056), .ZN(n10069) );
  OAI211_X1 U10937 ( .C1(n10060), .C2(n10059), .A(n10072), .B(n10058), .ZN(
        n10068) );
  MUX2_X1 U10938 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n7331), .S(n10061), .Z(
        n10064) );
  NAND3_X1 U10939 ( .A1(n10064), .A2(n10063), .A3(n10062), .ZN(n10065) );
  NAND3_X1 U10940 ( .A1(n10120), .A2(n10066), .A3(n10065), .ZN(n10067) );
  NAND3_X1 U10941 ( .A1(n10069), .A2(n10068), .A3(n10067), .ZN(P1_U3246) );
  INV_X1 U10942 ( .A(n10070), .ZN(n10071) );
  OAI211_X1 U10943 ( .C1(n10074), .C2(n10073), .A(n10072), .B(n10071), .ZN(
        n10087) );
  AOI21_X1 U10944 ( .B1(n10560), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10075), .ZN(
        n10086) );
  NAND2_X1 U10945 ( .A1(n10076), .A2(n10078), .ZN(n10085) );
  INV_X1 U10946 ( .A(n10077), .ZN(n10080) );
  MUX2_X1 U10947 ( .A(n7443), .B(P1_REG1_REG_5__SCAN_IN), .S(n10078), .Z(
        n10079) );
  NAND3_X1 U10948 ( .A1(n10081), .A2(n10080), .A3(n10079), .ZN(n10082) );
  NAND3_X1 U10949 ( .A1(n10120), .A2(n10083), .A3(n10082), .ZN(n10084) );
  NAND4_X1 U10950 ( .A1(n10087), .A2(n10086), .A3(n10085), .A4(n10084), .ZN(
        P1_U3248) );
  XNOR2_X1 U10951 ( .A(n10111), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n10092) );
  INV_X1 U10952 ( .A(n10088), .ZN(n10089) );
  OAI21_X1 U10953 ( .B1(n10096), .B2(P1_REG1_REG_17__SCAN_IN), .A(n10089), 
        .ZN(n10091) );
  NOR2_X1 U10954 ( .A1(n10092), .A2(n10091), .ZN(n10110) );
  AOI211_X1 U10955 ( .C1(n10092), .C2(n10091), .A(n10110), .B(n10090), .ZN(
        n10093) );
  INV_X1 U10956 ( .A(n10093), .ZN(n10104) );
  INV_X1 U10957 ( .A(n10094), .ZN(n10102) );
  OAI21_X1 U10958 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n10096), .A(n10095), 
        .ZN(n10100) );
  INV_X1 U10959 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n10098) );
  NOR2_X1 U10960 ( .A1(n10111), .A2(n10098), .ZN(n10097) );
  AOI21_X1 U10961 ( .B1(n10111), .B2(n10098), .A(n10097), .ZN(n10099) );
  NOR2_X1 U10962 ( .A1(n10100), .A2(n10099), .ZN(n10107) );
  AOI211_X1 U10963 ( .C1(n10100), .C2(n10099), .A(n10107), .B(n10122), .ZN(
        n10101) );
  AOI211_X1 U10964 ( .C1(n10560), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n10102), 
        .B(n10101), .ZN(n10103) );
  OAI211_X1 U10965 ( .C1(n10117), .C2(n10105), .A(n10104), .B(n10103), .ZN(
        P1_U3261) );
  INV_X1 U10966 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n10106) );
  MUX2_X1 U10967 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n10106), .S(n4966), .Z(
        n10109) );
  AOI21_X1 U10968 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n10111), .A(n10107), 
        .ZN(n10108) );
  XOR2_X1 U10969 ( .A(n10109), .B(n10108), .Z(n10123) );
  AOI21_X1 U10970 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n10111), .A(n10110), 
        .ZN(n10113) );
  INV_X1 U10971 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10407) );
  XNOR2_X1 U10972 ( .A(n4966), .B(n10407), .ZN(n10112) );
  XNOR2_X1 U10973 ( .A(n10113), .B(n10112), .ZN(n10119) );
  NAND2_X1 U10974 ( .A1(n10560), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n10114) );
  OAI211_X1 U10975 ( .C1(n10117), .C2(n10116), .A(n10115), .B(n10114), .ZN(
        n10118) );
  AOI21_X1 U10976 ( .B1(n10120), .B2(n10119), .A(n10118), .ZN(n10121) );
  OAI21_X1 U10977 ( .B1(n10123), .B2(n10122), .A(n10121), .ZN(P1_U3262) );
  NAND2_X1 U10978 ( .A1(n10152), .A2(n10147), .ZN(n10146) );
  INV_X1 U10979 ( .A(n10146), .ZN(n10131) );
  NAND2_X1 U10980 ( .A1(n10131), .A2(n10439), .ZN(n10130) );
  XNOR2_X1 U10981 ( .A(n10435), .B(n10130), .ZN(n10337) );
  NAND2_X1 U10982 ( .A1(n10337), .A2(n10178), .ZN(n10129) );
  AND2_X1 U10983 ( .A1(n10124), .A2(P1_B_REG_SCAN_IN), .ZN(n10125) );
  NOR2_X1 U10984 ( .A1(n10315), .A2(n10125), .ZN(n10139) );
  INV_X1 U10985 ( .A(n10139), .ZN(n10126) );
  NOR2_X1 U10986 ( .A1(n10335), .A2(n10340), .ZN(n10133) );
  AOI21_X1 U10987 ( .B1(n10335), .B2(P1_REG2_REG_31__SCAN_IN), .A(n10133), 
        .ZN(n10128) );
  OAI211_X1 U10988 ( .C1(n10435), .C2(n10325), .A(n10129), .B(n10128), .ZN(
        P1_U3263) );
  OAI211_X1 U10989 ( .C1(n10131), .C2(n10439), .A(n10292), .B(n10130), .ZN(
        n10341) );
  NOR2_X1 U10990 ( .A1(n10439), .A2(n10325), .ZN(n10132) );
  AOI211_X1 U10991 ( .C1(n10335), .C2(P1_REG2_REG_30__SCAN_IN), .A(n10133), 
        .B(n10132), .ZN(n10134) );
  OAI21_X1 U10992 ( .B1(n10341), .B2(n10264), .A(n10134), .ZN(P1_U3264) );
  XOR2_X1 U10993 ( .A(n10137), .B(n10143), .Z(n10140) );
  NAND2_X1 U10994 ( .A1(n10142), .A2(n10141), .ZN(n10145) );
  XNOR2_X1 U10995 ( .A(n10145), .B(n10144), .ZN(n10344) );
  OAI211_X1 U10996 ( .C1(n10152), .C2(n10147), .A(n10292), .B(n10146), .ZN(
        n10348) );
  NOR2_X1 U10997 ( .A1(n10348), .A2(n10264), .ZN(n10154) );
  INV_X1 U10998 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n10148) );
  OAI22_X1 U10999 ( .A1(n10149), .A2(n10326), .B1(n10148), .B2(n10328), .ZN(
        n10150) );
  AOI21_X1 U11000 ( .B1(n10345), .B2(n10159), .A(n10150), .ZN(n10151) );
  OAI21_X1 U11001 ( .B1(n10152), .B2(n10325), .A(n10151), .ZN(n10153) );
  AOI211_X1 U11002 ( .C1(n10344), .C2(n10321), .A(n10154), .B(n10153), .ZN(
        n10155) );
  OAI21_X1 U11003 ( .B1(n10350), .B2(n10335), .A(n10155), .ZN(P1_U3356) );
  NOR2_X1 U11004 ( .A1(n10156), .A2(n10293), .ZN(n10164) );
  INV_X1 U11005 ( .A(n10157), .ZN(n10162) );
  AOI22_X1 U11006 ( .A1(n10158), .A2(n10274), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n10335), .ZN(n10161) );
  NAND2_X1 U11007 ( .A1(n10188), .A2(n10159), .ZN(n10160) );
  OAI211_X1 U11008 ( .C1(n10162), .C2(n10325), .A(n10161), .B(n10160), .ZN(
        n10163) );
  AOI211_X1 U11009 ( .C1(n10165), .C2(n10328), .A(n10164), .B(n10163), .ZN(
        n10166) );
  OAI21_X1 U11010 ( .B1(n10167), .B2(n10307), .A(n10166), .ZN(P1_U3265) );
  OAI211_X1 U11011 ( .C1(n10171), .C2(n10170), .A(n10169), .B(n10312), .ZN(
        n10175) );
  OAI22_X1 U11012 ( .A1(n10172), .A2(n10315), .B1(n10208), .B2(n10395), .ZN(
        n10173) );
  INV_X1 U11013 ( .A(n10173), .ZN(n10174) );
  NAND2_X1 U11014 ( .A1(n10175), .A2(n10174), .ZN(n10354) );
  AOI21_X1 U11015 ( .B1(n10177), .B2(n4976), .A(n5240), .ZN(n10355) );
  NAND2_X1 U11016 ( .A1(n10355), .A2(n10178), .ZN(n10181) );
  AOI22_X1 U11017 ( .A1(n10179), .A2(n10274), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10335), .ZN(n10180) );
  OAI211_X1 U11018 ( .C1(n6149), .C2(n10325), .A(n10181), .B(n10180), .ZN(
        n10182) );
  AOI21_X1 U11019 ( .B1(n10328), .B2(n10354), .A(n10182), .ZN(n10183) );
  OAI21_X1 U11020 ( .B1(n10353), .B2(n10307), .A(n10183), .ZN(P1_U3266) );
  AND2_X1 U11021 ( .A1(n10184), .A2(n10185), .ZN(n10187) );
  OAI21_X1 U11022 ( .B1(n10187), .B2(n10190), .A(n10186), .ZN(n10189) );
  AOI22_X1 U11023 ( .A1(n10189), .A2(n10312), .B1(n10282), .B2(n10188), .ZN(
        n10359) );
  XNOR2_X1 U11024 ( .A(n10191), .B(n10190), .ZN(n10362) );
  NAND2_X1 U11025 ( .A1(n10362), .A2(n10321), .ZN(n10200) );
  INV_X1 U11026 ( .A(n10192), .ZN(n10193) );
  AOI22_X1 U11027 ( .A1(n10193), .A2(n10274), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n10335), .ZN(n10194) );
  OAI21_X1 U11028 ( .B1(n10360), .B2(n10278), .A(n10194), .ZN(n10197) );
  INV_X1 U11029 ( .A(n10195), .ZN(n10209) );
  OAI211_X1 U11030 ( .C1(n5242), .C2(n10209), .A(n10292), .B(n4976), .ZN(
        n10358) );
  NOR2_X1 U11031 ( .A1(n10358), .A2(n10264), .ZN(n10196) );
  AOI211_X1 U11032 ( .C1(n10297), .C2(n10198), .A(n10197), .B(n10196), .ZN(
        n10199) );
  OAI211_X1 U11033 ( .C1(n10335), .C2(n10359), .A(n10200), .B(n10199), .ZN(
        P1_U3267) );
  XNOR2_X1 U11034 ( .A(n10202), .B(n10201), .ZN(n10367) );
  INV_X1 U11035 ( .A(n10367), .ZN(n10218) );
  OAI211_X1 U11036 ( .C1(n10204), .C2(n10203), .A(n10184), .B(n10312), .ZN(
        n10207) );
  NAND2_X1 U11037 ( .A1(n10205), .A2(n10389), .ZN(n10206) );
  OAI211_X1 U11038 ( .C1(n10208), .C2(n10315), .A(n10207), .B(n10206), .ZN(
        n10365) );
  INV_X1 U11039 ( .A(n4961), .ZN(n10450) );
  AOI211_X1 U11040 ( .C1(n4961), .C2(n10210), .A(n10803), .B(n10209), .ZN(
        n10366) );
  NAND2_X1 U11041 ( .A1(n10366), .A2(n10286), .ZN(n10215) );
  INV_X1 U11042 ( .A(n10212), .ZN(n10213) );
  AOI22_X1 U11043 ( .A1(n10213), .A2(n10274), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10335), .ZN(n10214) );
  OAI211_X1 U11044 ( .C1(n10450), .C2(n10325), .A(n10215), .B(n10214), .ZN(
        n10216) );
  AOI21_X1 U11045 ( .B1(n10328), .B2(n10365), .A(n10216), .ZN(n10217) );
  OAI21_X1 U11046 ( .B1(n10218), .B2(n10307), .A(n10217), .ZN(P1_U3268) );
  OAI21_X1 U11047 ( .B1(n10221), .B2(n10220), .A(n10219), .ZN(n10224) );
  NOR2_X1 U11048 ( .A1(n10222), .A2(n10315), .ZN(n10223) );
  AOI21_X1 U11049 ( .B1(n10224), .B2(n10312), .A(n10223), .ZN(n10376) );
  XNOR2_X1 U11050 ( .A(n10226), .B(n10225), .ZN(n10379) );
  NAND2_X1 U11051 ( .A1(n10379), .A2(n10321), .ZN(n10236) );
  INV_X1 U11052 ( .A(n10227), .ZN(n10228) );
  AOI22_X1 U11053 ( .A1(n10228), .A2(n10274), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10335), .ZN(n10229) );
  OAI21_X1 U11054 ( .B1(n10377), .B2(n10278), .A(n10229), .ZN(n10233) );
  INV_X1 U11055 ( .A(n10230), .ZN(n10239) );
  OAI211_X1 U11056 ( .C1(n10455), .C2(n10239), .A(n10231), .B(n10292), .ZN(
        n10375) );
  NOR2_X1 U11057 ( .A1(n10375), .A2(n10264), .ZN(n10232) );
  AOI211_X1 U11058 ( .C1(n10297), .C2(n10234), .A(n10233), .B(n10232), .ZN(
        n10235) );
  OAI211_X1 U11059 ( .C1(n10335), .C2(n10376), .A(n10236), .B(n10235), .ZN(
        P1_U3270) );
  XNOR2_X1 U11060 ( .A(n10237), .B(n5514), .ZN(n10386) );
  AOI211_X1 U11061 ( .C1(n10383), .C2(n10262), .A(n10803), .B(n10239), .ZN(
        n10382) );
  INV_X1 U11062 ( .A(n10383), .ZN(n10243) );
  INV_X1 U11063 ( .A(n10240), .ZN(n10241) );
  AOI22_X1 U11064 ( .A1(n10241), .A2(n10274), .B1(n10335), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n10242) );
  OAI21_X1 U11065 ( .B1(n10243), .B2(n10325), .A(n10242), .ZN(n10248) );
  XNOR2_X1 U11066 ( .A(n5514), .B(n10244), .ZN(n10246) );
  AOI222_X1 U11067 ( .A1(n10312), .A2(n10246), .B1(n10245), .B2(n10282), .C1(
        n10281), .C2(n10389), .ZN(n10385) );
  NOR2_X1 U11068 ( .A1(n10385), .A2(n10335), .ZN(n10247) );
  AOI211_X1 U11069 ( .C1(n10382), .C2(n10331), .A(n10248), .B(n10247), .ZN(
        n10249) );
  OAI21_X1 U11070 ( .B1(n10307), .B2(n10386), .A(n10249), .ZN(P1_U3271) );
  NAND2_X1 U11071 ( .A1(n10251), .A2(n10250), .ZN(n10253) );
  XNOR2_X1 U11072 ( .A(n10253), .B(n10252), .ZN(n10255) );
  AOI22_X1 U11073 ( .A1(n10255), .A2(n10312), .B1(n10282), .B2(n10254), .ZN(
        n10393) );
  XNOR2_X1 U11074 ( .A(n10257), .B(n10256), .ZN(n10387) );
  NAND2_X1 U11075 ( .A1(n10387), .A2(n10321), .ZN(n10268) );
  INV_X1 U11076 ( .A(n10258), .ZN(n10259) );
  AOI22_X1 U11077 ( .A1(n10335), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n10259), 
        .B2(n10274), .ZN(n10260) );
  OAI21_X1 U11078 ( .B1(n10278), .B2(n10302), .A(n10260), .ZN(n10266) );
  INV_X1 U11079 ( .A(n10261), .ZN(n10272) );
  OAI211_X1 U11080 ( .C1(n10263), .C2(n10272), .A(n10292), .B(n10262), .ZN(
        n10391) );
  NOR2_X1 U11081 ( .A1(n10391), .A2(n10264), .ZN(n10265) );
  AOI211_X1 U11082 ( .C1(n10297), .C2(n10390), .A(n10266), .B(n10265), .ZN(
        n10267) );
  OAI211_X1 U11083 ( .C1(n10335), .C2(n10393), .A(n10268), .B(n10267), .ZN(
        P1_U3272) );
  INV_X1 U11084 ( .A(n10269), .ZN(n10270) );
  AOI21_X1 U11085 ( .B1(n10279), .B2(n10271), .A(n10270), .ZN(n10402) );
  AOI211_X1 U11086 ( .C1(n10273), .C2(n10291), .A(n10803), .B(n10272), .ZN(
        n10399) );
  NAND2_X1 U11087 ( .A1(n10273), .A2(n10297), .ZN(n10277) );
  AOI22_X1 U11088 ( .A1(n10335), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n10275), 
        .B2(n10274), .ZN(n10276) );
  OAI211_X1 U11089 ( .C1(n10396), .C2(n10278), .A(n10277), .B(n10276), .ZN(
        n10285) );
  XNOR2_X1 U11090 ( .A(n10280), .B(n10279), .ZN(n10283) );
  AOI22_X1 U11091 ( .A1(n10283), .A2(n10312), .B1(n10282), .B2(n10281), .ZN(
        n10401) );
  NOR2_X1 U11092 ( .A1(n10401), .A2(n10335), .ZN(n10284) );
  AOI211_X1 U11093 ( .C1(n10399), .C2(n10286), .A(n10285), .B(n10284), .ZN(
        n10287) );
  OAI21_X1 U11094 ( .B1(n10402), .B2(n10307), .A(n10287), .ZN(P1_U3273) );
  OAI21_X1 U11095 ( .B1(n10289), .B2(n5952), .A(n10288), .ZN(n10405) );
  OAI22_X1 U11096 ( .A1(n10328), .A2(n10106), .B1(n10290), .B2(n10326), .ZN(
        n10295) );
  OAI211_X1 U11097 ( .C1(n10462), .C2(n10322), .A(n10292), .B(n10291), .ZN(
        n10403) );
  NOR2_X1 U11098 ( .A1(n10403), .A2(n10293), .ZN(n10294) );
  AOI211_X1 U11099 ( .C1(n10297), .C2(n10296), .A(n10295), .B(n10294), .ZN(
        n10306) );
  OAI21_X1 U11100 ( .B1(n10300), .B2(n10299), .A(n10298), .ZN(n10304) );
  OAI22_X1 U11101 ( .A1(n10302), .A2(n10315), .B1(n10301), .B2(n10395), .ZN(
        n10303) );
  AOI21_X1 U11102 ( .B1(n10304), .B2(n10312), .A(n10303), .ZN(n10404) );
  OR2_X1 U11103 ( .A1(n10404), .A2(n10335), .ZN(n10305) );
  OAI211_X1 U11104 ( .C1(n10405), .C2(n10307), .A(n10306), .B(n10305), .ZN(
        P1_U3274) );
  NAND2_X1 U11105 ( .A1(n10309), .A2(n10308), .ZN(n10311) );
  INV_X1 U11106 ( .A(n10320), .ZN(n10310) );
  XNOR2_X1 U11107 ( .A(n10311), .B(n10310), .ZN(n10313) );
  NAND2_X1 U11108 ( .A1(n10313), .A2(n10312), .ZN(n10318) );
  OAI22_X1 U11109 ( .A1(n10396), .A2(n10315), .B1(n10314), .B2(n10395), .ZN(
        n10316) );
  INV_X1 U11110 ( .A(n10316), .ZN(n10317) );
  NAND2_X1 U11111 ( .A1(n10318), .A2(n10317), .ZN(n10409) );
  INV_X1 U11112 ( .A(n10409), .ZN(n10334) );
  XNOR2_X1 U11113 ( .A(n10319), .B(n10320), .ZN(n10411) );
  NAND2_X1 U11114 ( .A1(n10411), .A2(n10321), .ZN(n10333) );
  AOI211_X1 U11115 ( .C1(n10324), .C2(n10323), .A(n10803), .B(n10322), .ZN(
        n10410) );
  NOR2_X1 U11116 ( .A1(n5235), .A2(n10325), .ZN(n10330) );
  OAI22_X1 U11117 ( .A1(n10328), .A2(n10098), .B1(n10327), .B2(n10326), .ZN(
        n10329) );
  AOI211_X1 U11118 ( .C1(n10410), .C2(n10331), .A(n10330), .B(n10329), .ZN(
        n10332) );
  OAI211_X1 U11119 ( .C1(n10335), .C2(n10334), .A(n10333), .B(n10332), .ZN(
        P1_U3275) );
  INV_X1 U11120 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10338) );
  INV_X1 U11121 ( .A(n10340), .ZN(n10336) );
  AOI21_X1 U11122 ( .B1(n10337), .B2(n10292), .A(n10336), .ZN(n10432) );
  MUX2_X1 U11123 ( .A(n10338), .B(n10432), .S(n10842), .Z(n10339) );
  OAI21_X1 U11124 ( .B1(n10435), .B2(n10419), .A(n10339), .ZN(P1_U3553) );
  INV_X1 U11125 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10342) );
  AND2_X1 U11126 ( .A1(n10341), .A2(n10340), .ZN(n10436) );
  MUX2_X1 U11127 ( .A(n10342), .B(n10436), .S(n10842), .Z(n10343) );
  OAI21_X1 U11128 ( .B1(n10439), .B2(n10419), .A(n10343), .ZN(P1_U3552) );
  NAND2_X1 U11129 ( .A1(n10344), .A2(n10838), .ZN(n10352) );
  AOI22_X1 U11130 ( .A1(n10346), .A2(n10428), .B1(n10389), .B2(n10345), .ZN(
        n10347) );
  NAND2_X1 U11131 ( .A1(n10352), .A2(n10351), .ZN(n10440) );
  MUX2_X1 U11132 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10440), .S(n10842), .Z(
        P1_U3551) );
  MUX2_X1 U11133 ( .A(n10356), .B(n10441), .S(n10842), .Z(n10357) );
  OAI21_X1 U11134 ( .B1(n6149), .B2(n10419), .A(n10357), .ZN(P1_U3549) );
  OAI211_X1 U11135 ( .C1(n10360), .C2(n10395), .A(n10359), .B(n10358), .ZN(
        n10361) );
  AOI21_X1 U11136 ( .B1(n10362), .B2(n10838), .A(n10361), .ZN(n10444) );
  MUX2_X1 U11137 ( .A(n10363), .B(n10444), .S(n10842), .Z(n10364) );
  OAI21_X1 U11138 ( .B1(n5242), .B2(n10419), .A(n10364), .ZN(P1_U3548) );
  AOI211_X1 U11139 ( .C1(n10367), .C2(n10838), .A(n10366), .B(n10365), .ZN(
        n10447) );
  MUX2_X1 U11140 ( .A(n10368), .B(n10447), .S(n10842), .Z(n10369) );
  OAI21_X1 U11141 ( .B1(n10450), .B2(n10419), .A(n10369), .ZN(P1_U3547) );
  AOI211_X1 U11142 ( .C1(n10428), .C2(n10372), .A(n10371), .B(n10370), .ZN(
        n10373) );
  OAI21_X1 U11143 ( .B1(n10374), .B2(n10425), .A(n10373), .ZN(n10451) );
  MUX2_X1 U11144 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10451), .S(n10842), .Z(
        P1_U3546) );
  OAI211_X1 U11145 ( .C1(n10377), .C2(n10395), .A(n10376), .B(n10375), .ZN(
        n10378) );
  AOI21_X1 U11146 ( .B1(n10379), .B2(n10838), .A(n10378), .ZN(n10452) );
  MUX2_X1 U11147 ( .A(n10380), .B(n10452), .S(n10842), .Z(n10381) );
  OAI21_X1 U11148 ( .B1(n10455), .B2(n10419), .A(n10381), .ZN(P1_U3545) );
  AOI21_X1 U11149 ( .B1(n10428), .B2(n10383), .A(n10382), .ZN(n10384) );
  OAI211_X1 U11150 ( .C1(n10386), .C2(n10425), .A(n10385), .B(n10384), .ZN(
        n10456) );
  MUX2_X1 U11151 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10456), .S(n10842), .Z(
        P1_U3544) );
  NAND2_X1 U11152 ( .A1(n10387), .A2(n10838), .ZN(n10394) );
  AOI22_X1 U11153 ( .A1(n10390), .A2(n10428), .B1(n10389), .B2(n10388), .ZN(
        n10392) );
  NAND4_X1 U11154 ( .A1(n10394), .A2(n10393), .A3(n10392), .A4(n10391), .ZN(
        n10457) );
  MUX2_X1 U11155 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10457), .S(n10842), .Z(
        P1_U3543) );
  OAI22_X1 U11156 ( .A1(n10397), .A2(n10835), .B1(n10396), .B2(n10395), .ZN(
        n10398) );
  NOR2_X1 U11157 ( .A1(n10399), .A2(n10398), .ZN(n10400) );
  OAI211_X1 U11158 ( .C1(n10402), .C2(n10425), .A(n10401), .B(n10400), .ZN(
        n10458) );
  MUX2_X1 U11159 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10458), .S(n10842), .Z(
        P1_U3542) );
  OAI211_X1 U11160 ( .C1(n10405), .C2(n10425), .A(n10404), .B(n10403), .ZN(
        n10406) );
  INV_X1 U11161 ( .A(n10406), .ZN(n10459) );
  MUX2_X1 U11162 ( .A(n10407), .B(n10459), .S(n10842), .Z(n10408) );
  OAI21_X1 U11163 ( .B1(n10462), .B2(n10419), .A(n10408), .ZN(P1_U3541) );
  AOI211_X1 U11164 ( .C1(n10411), .C2(n10838), .A(n10410), .B(n10409), .ZN(
        n10463) );
  MUX2_X1 U11165 ( .A(n10412), .B(n10463), .S(n10842), .Z(n10413) );
  OAI21_X1 U11166 ( .B1(n5235), .B2(n10419), .A(n10413), .ZN(P1_U3540) );
  INV_X1 U11167 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10417) );
  AOI211_X1 U11168 ( .C1(n10416), .C2(n10838), .A(n10415), .B(n10414), .ZN(
        n10466) );
  MUX2_X1 U11169 ( .A(n10417), .B(n10466), .S(n10842), .Z(n10418) );
  OAI21_X1 U11170 ( .B1(n10470), .B2(n10419), .A(n10418), .ZN(P1_U3539) );
  AOI211_X1 U11171 ( .C1(n10428), .C2(n10422), .A(n10421), .B(n10420), .ZN(
        n10423) );
  OAI21_X1 U11172 ( .B1(n10425), .B2(n10424), .A(n10423), .ZN(n10471) );
  MUX2_X1 U11173 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10471), .S(n10842), .Z(
        P1_U3538) );
  AOI21_X1 U11174 ( .B1(n10428), .B2(n10427), .A(n10426), .ZN(n10429) );
  OAI211_X1 U11175 ( .C1(n10793), .C2(n10431), .A(n10430), .B(n10429), .ZN(
        n10472) );
  MUX2_X1 U11176 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10472), .S(n10842), .Z(
        P1_U3536) );
  INV_X1 U11177 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10433) );
  MUX2_X1 U11178 ( .A(n10433), .B(n10432), .S(n10846), .Z(n10434) );
  OAI21_X1 U11179 ( .B1(n10435), .B2(n10469), .A(n10434), .ZN(P1_U3521) );
  INV_X1 U11180 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10437) );
  MUX2_X1 U11181 ( .A(n10437), .B(n10436), .S(n10846), .Z(n10438) );
  OAI21_X1 U11182 ( .B1(n10439), .B2(n10469), .A(n10438), .ZN(P1_U3520) );
  MUX2_X1 U11183 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10440), .S(n10846), .Z(
        P1_U3519) );
  INV_X1 U11184 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10442) );
  MUX2_X1 U11185 ( .A(n10442), .B(n10441), .S(n10846), .Z(n10443) );
  OAI21_X1 U11186 ( .B1(n6149), .B2(n10469), .A(n10443), .ZN(P1_U3517) );
  INV_X1 U11187 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10445) );
  MUX2_X1 U11188 ( .A(n10445), .B(n10444), .S(n10846), .Z(n10446) );
  OAI21_X1 U11189 ( .B1(n5242), .B2(n10469), .A(n10446), .ZN(P1_U3516) );
  INV_X1 U11190 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10448) );
  MUX2_X1 U11191 ( .A(n10448), .B(n10447), .S(n10846), .Z(n10449) );
  OAI21_X1 U11192 ( .B1(n10450), .B2(n10469), .A(n10449), .ZN(P1_U3515) );
  MUX2_X1 U11193 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10451), .S(n10846), .Z(
        P1_U3514) );
  INV_X1 U11194 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10453) );
  MUX2_X1 U11195 ( .A(n10453), .B(n10452), .S(n10846), .Z(n10454) );
  OAI21_X1 U11196 ( .B1(n10455), .B2(n10469), .A(n10454), .ZN(P1_U3513) );
  MUX2_X1 U11197 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10456), .S(n10846), .Z(
        P1_U3512) );
  MUX2_X1 U11198 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10457), .S(n10846), .Z(
        P1_U3511) );
  MUX2_X1 U11199 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10458), .S(n10846), .Z(
        P1_U3510) );
  INV_X1 U11200 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10460) );
  MUX2_X1 U11201 ( .A(n10460), .B(n10459), .S(n10846), .Z(n10461) );
  OAI21_X1 U11202 ( .B1(n10462), .B2(n10469), .A(n10461), .ZN(P1_U3509) );
  INV_X1 U11203 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10464) );
  MUX2_X1 U11204 ( .A(n10464), .B(n10463), .S(n10846), .Z(n10465) );
  OAI21_X1 U11205 ( .B1(n5235), .B2(n10469), .A(n10465), .ZN(P1_U3507) );
  INV_X1 U11206 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n10467) );
  MUX2_X1 U11207 ( .A(n10467), .B(n10466), .S(n10846), .Z(n10468) );
  OAI21_X1 U11208 ( .B1(n10470), .B2(n10469), .A(n10468), .ZN(P1_U3504) );
  MUX2_X1 U11209 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10471), .S(n10846), .Z(
        P1_U3501) );
  MUX2_X1 U11210 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10472), .S(n10846), .Z(
        P1_U3495) );
  MUX2_X1 U11211 ( .A(n10473), .B(P1_D_REG_0__SCAN_IN), .S(n10497), .Z(
        P1_U3439) );
  NOR4_X1 U11212 ( .A1(n10475), .A2(P1_IR_REG_30__SCAN_IN), .A3(n10474), .A4(
        P1_U3086), .ZN(n10476) );
  AOI21_X1 U11213 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n10477), .A(n10476), 
        .ZN(n10478) );
  OAI21_X1 U11214 ( .B1(n10479), .B2(n10492), .A(n10478), .ZN(P1_U3324) );
  OAI222_X1 U11215 ( .A1(n10494), .A2(n10482), .B1(P1_U3086), .B2(n10481), 
        .C1(n10492), .C2(n10480), .ZN(P1_U3326) );
  OAI222_X1 U11216 ( .A1(n10485), .A2(P1_U3086), .B1(n10492), .B2(n10484), 
        .C1(n10483), .C2(n10494), .ZN(P1_U3327) );
  INV_X1 U11217 ( .A(n10486), .ZN(n10488) );
  OAI222_X1 U11218 ( .A1(n10489), .A2(P1_U3086), .B1(n10492), .B2(n10488), 
        .C1(n10487), .C2(n10494), .ZN(P1_U3328) );
  OAI222_X1 U11219 ( .A1(n10494), .A2(n10493), .B1(n10492), .B2(n10491), .C1(
        n10490), .C2(P1_U3086), .ZN(P1_U3329) );
  INV_X1 U11220 ( .A(n10495), .ZN(n10496) );
  MUX2_X1 U11221 ( .A(n10496), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AND2_X1 U11222 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10497), .ZN(P1_U3323) );
  AND2_X1 U11223 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10497), .ZN(P1_U3322) );
  AND2_X1 U11224 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10497), .ZN(P1_U3321) );
  AND2_X1 U11225 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10497), .ZN(P1_U3320) );
  AND2_X1 U11226 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10497), .ZN(P1_U3319) );
  AND2_X1 U11227 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10497), .ZN(P1_U3318) );
  AND2_X1 U11228 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10497), .ZN(P1_U3317) );
  AND2_X1 U11229 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10497), .ZN(P1_U3316) );
  AND2_X1 U11230 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10497), .ZN(P1_U3315) );
  AND2_X1 U11231 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10497), .ZN(P1_U3314) );
  AND2_X1 U11232 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10497), .ZN(P1_U3313) );
  AND2_X1 U11233 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10497), .ZN(P1_U3312) );
  AND2_X1 U11234 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10497), .ZN(P1_U3311) );
  AND2_X1 U11235 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10497), .ZN(P1_U3310) );
  AND2_X1 U11236 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10497), .ZN(P1_U3309) );
  AND2_X1 U11237 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10497), .ZN(P1_U3308) );
  AND2_X1 U11238 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10497), .ZN(P1_U3307) );
  AND2_X1 U11239 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10497), .ZN(P1_U3306) );
  AND2_X1 U11240 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10497), .ZN(P1_U3305) );
  AND2_X1 U11241 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10497), .ZN(P1_U3304) );
  AND2_X1 U11242 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10497), .ZN(P1_U3303) );
  AND2_X1 U11243 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10497), .ZN(P1_U3302) );
  AND2_X1 U11244 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10497), .ZN(P1_U3301) );
  AND2_X1 U11245 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10497), .ZN(P1_U3300) );
  AND2_X1 U11246 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10497), .ZN(P1_U3299) );
  AND2_X1 U11247 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10497), .ZN(P1_U3298) );
  AND2_X1 U11248 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10497), .ZN(P1_U3297) );
  AND2_X1 U11249 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10497), .ZN(P1_U3296) );
  AND2_X1 U11250 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10497), .ZN(P1_U3295) );
  AND2_X1 U11251 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10497), .ZN(P1_U3294) );
  XOR2_X1 U11252 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI222_X1 U11253 ( .A1(n10588), .A2(n10501), .B1(n10588), .B2(n10500), .C1(
        n10499), .C2(n10498), .ZN(ADD_1068_U5) );
  AOI21_X1 U11254 ( .B1(n10504), .B2(n10503), .A(n10502), .ZN(ADD_1068_U54) );
  AOI21_X1 U11255 ( .B1(n10507), .B2(n10506), .A(n10505), .ZN(ADD_1068_U53) );
  OAI21_X1 U11256 ( .B1(n10510), .B2(n10509), .A(n10508), .ZN(ADD_1068_U52) );
  OAI21_X1 U11257 ( .B1(n10513), .B2(n10512), .A(n10511), .ZN(ADD_1068_U51) );
  OAI21_X1 U11258 ( .B1(n10516), .B2(n10515), .A(n10514), .ZN(ADD_1068_U50) );
  OAI21_X1 U11259 ( .B1(n10519), .B2(n10518), .A(n10517), .ZN(ADD_1068_U49) );
  OAI21_X1 U11260 ( .B1(n10522), .B2(n10521), .A(n10520), .ZN(ADD_1068_U48) );
  OAI21_X1 U11261 ( .B1(n10525), .B2(n10524), .A(n10523), .ZN(ADD_1068_U47) );
  OAI21_X1 U11262 ( .B1(n10528), .B2(n10527), .A(n10526), .ZN(ADD_1068_U63) );
  OAI21_X1 U11263 ( .B1(n10531), .B2(n10530), .A(n10529), .ZN(ADD_1068_U62) );
  OAI21_X1 U11264 ( .B1(n10534), .B2(n10533), .A(n10532), .ZN(ADD_1068_U61) );
  OAI21_X1 U11265 ( .B1(n10537), .B2(n10536), .A(n10535), .ZN(ADD_1068_U60) );
  OAI21_X1 U11266 ( .B1(n10540), .B2(n10539), .A(n10538), .ZN(ADD_1068_U59) );
  OAI21_X1 U11267 ( .B1(n10543), .B2(n10542), .A(n10541), .ZN(ADD_1068_U58) );
  OAI21_X1 U11268 ( .B1(n10546), .B2(n10545), .A(n10544), .ZN(ADD_1068_U57) );
  OAI21_X1 U11269 ( .B1(n10549), .B2(n10548), .A(n10547), .ZN(ADD_1068_U56) );
  OAI21_X1 U11270 ( .B1(n10552), .B2(n10551), .A(n10550), .ZN(ADD_1068_U55) );
  INV_X1 U11271 ( .A(n10553), .ZN(n10556) );
  OAI22_X1 U11272 ( .A1(n10556), .A2(n6957), .B1(n10555), .B2(n10554), .ZN(
        n10558) );
  XOR2_X1 U11273 ( .A(n10558), .B(n10557), .Z(n10562) );
  AOI22_X1 U11274 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n10560), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n10561) );
  OAI21_X1 U11275 ( .B1(n10563), .B2(n10562), .A(n10561), .ZN(P1_U3243) );
  AOI22_X1 U11276 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(n10737), .B1(n10757), .B2(
        P2_ADDR_REG_0__SCAN_IN), .ZN(n10569) );
  INV_X1 U11277 ( .A(n10564), .ZN(n10567) );
  OAI21_X1 U11278 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n10565), .A(n10583), .ZN(
        n10566) );
  OAI21_X1 U11279 ( .B1(n10567), .B2(n10772), .A(n10566), .ZN(n10568) );
  OAI211_X1 U11280 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10570), .A(n10569), .B(
        n10568), .ZN(P2_U3182) );
  INV_X1 U11281 ( .A(n10572), .ZN(n10573) );
  AOI21_X1 U11282 ( .B1(n10575), .B2(n10574), .A(n10573), .ZN(n10581) );
  OAI21_X1 U11283 ( .B1(n5276), .B2(P2_REG1_REG_1__SCAN_IN), .A(n10577), .ZN(
        n10579) );
  AOI22_X1 U11284 ( .A1(n10745), .A2(n10579), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(P2_U3151), .ZN(n10580) );
  OAI21_X1 U11285 ( .B1(n10581), .B2(n10747), .A(n10580), .ZN(n10582) );
  AOI21_X1 U11286 ( .B1(n6245), .B2(n10737), .A(n10582), .ZN(n10587) );
  XOR2_X1 U11287 ( .A(n10584), .B(n10583), .Z(n10585) );
  NAND2_X1 U11288 ( .A1(n10585), .A2(n10772), .ZN(n10586) );
  OAI211_X1 U11289 ( .C1(n10588), .C2(n10605), .A(n10587), .B(n10586), .ZN(
        P2_U3183) );
  INV_X1 U11290 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10606) );
  AOI21_X1 U11291 ( .B1(n10591), .B2(n10590), .A(n10589), .ZN(n10597) );
  XOR2_X1 U11292 ( .A(n10593), .B(n10592), .Z(n10595) );
  AOI21_X1 U11293 ( .B1(n10745), .B2(n10595), .A(n10594), .ZN(n10596) );
  OAI21_X1 U11294 ( .B1(n10597), .B2(n10747), .A(n10596), .ZN(n10598) );
  AOI21_X1 U11295 ( .B1(n10599), .B2(n10737), .A(n10598), .ZN(n10604) );
  OAI211_X1 U11296 ( .C1(n10602), .C2(n10601), .A(n10600), .B(n10772), .ZN(
        n10603) );
  OAI211_X1 U11297 ( .C1(n10606), .C2(n10605), .A(n10604), .B(n10603), .ZN(
        P2_U3186) );
  OAI21_X1 U11298 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(n10608), .A(n10607), .ZN(
        n10609) );
  AOI22_X1 U11299 ( .A1(n10737), .A2(n10610), .B1(n10745), .B2(n10609), .ZN(
        n10622) );
  AOI21_X1 U11300 ( .B1(n10613), .B2(n10612), .A(n10611), .ZN(n10614) );
  NOR2_X1 U11301 ( .A1(n10614), .A2(n10747), .ZN(n10615) );
  AOI211_X1 U11302 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n10757), .A(n10616), .B(
        n10615), .ZN(n10621) );
  OAI211_X1 U11303 ( .C1(n10619), .C2(n10618), .A(n10617), .B(n10772), .ZN(
        n10620) );
  NAND3_X1 U11304 ( .A1(n10622), .A2(n10621), .A3(n10620), .ZN(P2_U3187) );
  AOI22_X1 U11305 ( .A1(n10623), .A2(n10737), .B1(n10757), .B2(
        P2_ADDR_REG_10__SCAN_IN), .ZN(n10640) );
  INV_X1 U11306 ( .A(n10624), .ZN(n10626) );
  NAND2_X1 U11307 ( .A1(n10626), .A2(n10625), .ZN(n10627) );
  XNOR2_X1 U11308 ( .A(n10628), .B(n10627), .ZN(n10633) );
  OAI21_X1 U11309 ( .B1(n10631), .B2(n10630), .A(n10629), .ZN(n10632) );
  AOI22_X1 U11310 ( .A1(n10633), .A2(n10772), .B1(n10745), .B2(n10632), .ZN(
        n10639) );
  NAND2_X1 U11311 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3151), .ZN(n10638)
         );
  AOI21_X1 U11312 ( .B1(n5039), .B2(n10635), .A(n10634), .ZN(n10636) );
  OR2_X1 U11313 ( .A1(n10636), .A2(n10747), .ZN(n10637) );
  NAND4_X1 U11314 ( .A1(n10640), .A2(n10639), .A3(n10638), .A4(n10637), .ZN(
        P2_U3192) );
  AOI22_X1 U11315 ( .A1(n10641), .A2(n10737), .B1(n10757), .B2(
        P2_ADDR_REG_11__SCAN_IN), .ZN(n10656) );
  OAI21_X1 U11316 ( .B1(n10644), .B2(n10643), .A(n10642), .ZN(n10648) );
  OAI21_X1 U11317 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n10646), .A(n10645), 
        .ZN(n10647) );
  AOI22_X1 U11318 ( .A1(n10648), .A2(n10772), .B1(n10745), .B2(n10647), .ZN(
        n10655) );
  NAND2_X1 U11319 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3151), .ZN(n10654)
         );
  AOI21_X1 U11320 ( .B1(n10651), .B2(n10650), .A(n10649), .ZN(n10652) );
  OR2_X1 U11321 ( .A1(n10747), .A2(n10652), .ZN(n10653) );
  NAND4_X1 U11322 ( .A1(n10656), .A2(n10655), .A3(n10654), .A4(n10653), .ZN(
        P2_U3193) );
  AOI22_X1 U11323 ( .A1(n10657), .A2(n10737), .B1(n10757), .B2(
        P2_ADDR_REG_12__SCAN_IN), .ZN(n10672) );
  OAI21_X1 U11324 ( .B1(n10660), .B2(n10659), .A(n10658), .ZN(n10665) );
  OAI21_X1 U11325 ( .B1(n10663), .B2(n10662), .A(n10661), .ZN(n10664) );
  AOI22_X1 U11326 ( .A1(n10665), .A2(n10745), .B1(n10772), .B2(n10664), .ZN(
        n10671) );
  AOI21_X1 U11327 ( .B1(n5031), .B2(n10667), .A(n10666), .ZN(n10668) );
  OR2_X1 U11328 ( .A1(n10668), .A2(n10747), .ZN(n10669) );
  NAND4_X1 U11329 ( .A1(n10672), .A2(n10671), .A3(n10670), .A4(n10669), .ZN(
        P2_U3194) );
  AOI22_X1 U11330 ( .A1(n10673), .A2(n10737), .B1(n10757), .B2(
        P2_ADDR_REG_13__SCAN_IN), .ZN(n10688) );
  OAI21_X1 U11331 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n10675), .A(n10674), 
        .ZN(n10680) );
  OAI21_X1 U11332 ( .B1(n10678), .B2(n10677), .A(n10676), .ZN(n10679) );
  AOI22_X1 U11333 ( .A1(n10680), .A2(n10745), .B1(n10772), .B2(n10679), .ZN(
        n10687) );
  NAND2_X1 U11334 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3151), .ZN(n10686)
         );
  AOI21_X1 U11335 ( .B1(n10683), .B2(n10682), .A(n10681), .ZN(n10684) );
  OR2_X1 U11336 ( .A1(n10747), .A2(n10684), .ZN(n10685) );
  NAND4_X1 U11337 ( .A1(n10688), .A2(n10687), .A3(n10686), .A4(n10685), .ZN(
        P2_U3195) );
  AOI22_X1 U11338 ( .A1(n10689), .A2(n10737), .B1(n10757), .B2(
        P2_ADDR_REG_14__SCAN_IN), .ZN(n10704) );
  OAI21_X1 U11339 ( .B1(n10692), .B2(n10691), .A(n10690), .ZN(n10697) );
  OAI21_X1 U11340 ( .B1(n10695), .B2(n10694), .A(n10693), .ZN(n10696) );
  AOI22_X1 U11341 ( .A1(n10697), .A2(n10745), .B1(n10772), .B2(n10696), .ZN(
        n10703) );
  NAND2_X1 U11342 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3151), .ZN(n10702)
         );
  AOI21_X1 U11343 ( .B1(n5033), .B2(n10699), .A(n10698), .ZN(n10700) );
  OR2_X1 U11344 ( .A1(n10700), .A2(n10747), .ZN(n10701) );
  NAND4_X1 U11345 ( .A1(n10704), .A2(n10703), .A3(n10702), .A4(n10701), .ZN(
        P2_U3196) );
  AOI22_X1 U11346 ( .A1(n10705), .A2(n10737), .B1(n10757), .B2(
        P2_ADDR_REG_15__SCAN_IN), .ZN(n10720) );
  OAI21_X1 U11347 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n10707), .A(n10706), 
        .ZN(n10712) );
  OAI21_X1 U11348 ( .B1(n10710), .B2(n10709), .A(n10708), .ZN(n10711) );
  AOI22_X1 U11349 ( .A1(n10712), .A2(n10745), .B1(n10772), .B2(n10711), .ZN(
        n10719) );
  AOI21_X1 U11350 ( .B1(n10715), .B2(n10714), .A(n10713), .ZN(n10716) );
  OR2_X1 U11351 ( .A1(n10747), .A2(n10716), .ZN(n10717) );
  NAND4_X1 U11352 ( .A1(n10720), .A2(n10719), .A3(n10718), .A4(n10717), .ZN(
        P2_U3197) );
  AOI22_X1 U11353 ( .A1(n10721), .A2(n10737), .B1(n10757), .B2(
        P2_ADDR_REG_16__SCAN_IN), .ZN(n10736) );
  OAI21_X1 U11354 ( .B1(n10724), .B2(n10723), .A(n10722), .ZN(n10729) );
  OAI21_X1 U11355 ( .B1(n10727), .B2(n10726), .A(n10725), .ZN(n10728) );
  AOI22_X1 U11356 ( .A1(n10729), .A2(n10745), .B1(n10772), .B2(n10728), .ZN(
        n10735) );
  AOI21_X1 U11357 ( .B1(n4999), .B2(n10731), .A(n10730), .ZN(n10732) );
  OR2_X1 U11358 ( .A1(n10732), .A2(n10747), .ZN(n10733) );
  NAND4_X1 U11359 ( .A1(n10736), .A2(n10735), .A3(n10734), .A4(n10733), .ZN(
        P2_U3198) );
  AOI22_X1 U11360 ( .A1(n10738), .A2(n10737), .B1(n10757), .B2(
        P2_ADDR_REG_17__SCAN_IN), .ZN(n10752) );
  OAI21_X1 U11361 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n10740), .A(n10739), 
        .ZN(n10746) );
  OAI21_X1 U11362 ( .B1(n10743), .B2(n10742), .A(n10741), .ZN(n10744) );
  AOI22_X1 U11363 ( .A1(n10746), .A2(n10745), .B1(n10772), .B2(n10744), .ZN(
        n10751) );
  OAI21_X1 U11364 ( .B1(n4981), .B2(P2_REG2_REG_17__SCAN_IN), .A(n10759), .ZN(
        n10748) );
  NAND2_X1 U11365 ( .A1(n10748), .A2(n9468), .ZN(n10749) );
  NAND4_X1 U11366 ( .A1(n10752), .A2(n10751), .A3(n10750), .A4(n10749), .ZN(
        P2_U3199) );
  INV_X1 U11367 ( .A(n10762), .ZN(n10764) );
  NAND2_X1 U11368 ( .A1(n10764), .A2(n10763), .ZN(n10773) );
  OAI21_X1 U11369 ( .B1(n10773), .B2(n10766), .A(n10765), .ZN(n10768) );
  NAND3_X1 U11370 ( .A1(n10773), .A2(n10772), .A3(n10771), .ZN(n10774) );
  XOR2_X1 U11371 ( .A(n10776), .B(P1_RD_REG_SCAN_IN), .Z(U126) );
  INV_X1 U11372 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10777) );
  AOI22_X1 U11373 ( .A1(n10851), .A2(n10778), .B1(n10777), .B2(n7244), .ZN(
        P2_U3393) );
  INV_X1 U11374 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10779) );
  AOI22_X1 U11375 ( .A1(n10851), .A2(n10780), .B1(n10779), .B2(n7244), .ZN(
        P2_U3399) );
  INV_X1 U11376 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10781) );
  AOI22_X1 U11377 ( .A1(n10851), .A2(n10782), .B1(n10781), .B2(n7244), .ZN(
        P2_U3402) );
  OAI21_X1 U11378 ( .B1(n10784), .B2(n10835), .A(n10783), .ZN(n10786) );
  AOI211_X1 U11379 ( .C1(n10838), .C2(n10787), .A(n10786), .B(n10785), .ZN(
        n10790) );
  AOI22_X1 U11380 ( .A1(n10842), .A2(n10790), .B1(n10788), .B2(n10840), .ZN(
        P1_U3526) );
  INV_X1 U11381 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10789) );
  AOI22_X1 U11382 ( .A1(n10846), .A2(n10790), .B1(n10789), .B2(n10843), .ZN(
        P1_U3465) );
  INV_X1 U11383 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10791) );
  AOI22_X1 U11384 ( .A1(n10851), .A2(n10792), .B1(n10791), .B2(n7244), .ZN(
        P2_U3408) );
  INV_X1 U11385 ( .A(n10793), .ZN(n10799) );
  OAI21_X1 U11386 ( .B1(n10795), .B2(n10835), .A(n10794), .ZN(n10797) );
  AOI211_X1 U11387 ( .C1(n10799), .C2(n10798), .A(n10797), .B(n10796), .ZN(
        n10801) );
  AOI22_X1 U11388 ( .A1(n10842), .A2(n10801), .B1(n7441), .B2(n10840), .ZN(
        P1_U3528) );
  INV_X1 U11389 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10800) );
  AOI22_X1 U11390 ( .A1(n10846), .A2(n10801), .B1(n10800), .B2(n10843), .ZN(
        P1_U3471) );
  OAI22_X1 U11391 ( .A1(n10804), .A2(n10803), .B1(n10802), .B2(n10835), .ZN(
        n10806) );
  AOI211_X1 U11392 ( .C1(n10838), .C2(n10807), .A(n10806), .B(n10805), .ZN(
        n10809) );
  AOI22_X1 U11393 ( .A1(n10842), .A2(n10809), .B1(n7464), .B2(n10840), .ZN(
        P1_U3530) );
  INV_X1 U11394 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10808) );
  AOI22_X1 U11395 ( .A1(n10846), .A2(n10809), .B1(n10808), .B2(n10843), .ZN(
        P1_U3477) );
  INV_X1 U11396 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10810) );
  AOI22_X1 U11397 ( .A1(n10851), .A2(n10811), .B1(n10810), .B2(n7244), .ZN(
        P2_U3414) );
  OAI211_X1 U11398 ( .C1(n10814), .C2(n10835), .A(n10813), .B(n10812), .ZN(
        n10815) );
  AOI21_X1 U11399 ( .B1(n10838), .B2(n10816), .A(n10815), .ZN(n10818) );
  AOI22_X1 U11400 ( .A1(n10842), .A2(n10818), .B1(n7484), .B2(n10840), .ZN(
        P1_U3531) );
  INV_X1 U11401 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10817) );
  AOI22_X1 U11402 ( .A1(n10846), .A2(n10818), .B1(n10817), .B2(n10843), .ZN(
        P1_U3480) );
  OAI211_X1 U11403 ( .C1(n10821), .C2(n10835), .A(n10820), .B(n10819), .ZN(
        n10822) );
  AOI21_X1 U11404 ( .B1(n10823), .B2(n10838), .A(n10822), .ZN(n10826) );
  AOI22_X1 U11405 ( .A1(n10842), .A2(n10826), .B1(n10824), .B2(n10840), .ZN(
        P1_U3532) );
  INV_X1 U11406 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10825) );
  AOI22_X1 U11407 ( .A1(n10846), .A2(n10826), .B1(n10825), .B2(n10843), .ZN(
        P1_U3483) );
  INV_X1 U11408 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10827) );
  AOI22_X1 U11409 ( .A1(n10851), .A2(n10828), .B1(n10827), .B2(n7244), .ZN(
        P2_U3420) );
  INV_X1 U11410 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10829) );
  AOI22_X1 U11411 ( .A1(n10851), .A2(n10830), .B1(n10829), .B2(n7244), .ZN(
        P2_U3423) );
  INV_X1 U11412 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10831) );
  AOI22_X1 U11413 ( .A1(n10851), .A2(n10832), .B1(n10831), .B2(n7244), .ZN(
        P2_U3426) );
  OAI211_X1 U11414 ( .C1(n10836), .C2(n10835), .A(n10834), .B(n10833), .ZN(
        n10837) );
  AOI21_X1 U11415 ( .B1(n10839), .B2(n10838), .A(n10837), .ZN(n10845) );
  AOI22_X1 U11416 ( .A1(n10842), .A2(n10845), .B1(n10841), .B2(n10840), .ZN(
        P1_U3534) );
  INV_X1 U11417 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10844) );
  AOI22_X1 U11418 ( .A1(n10846), .A2(n10845), .B1(n10844), .B2(n10843), .ZN(
        P1_U3489) );
  INV_X1 U11419 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10847) );
  AOI22_X1 U11420 ( .A1(n10851), .A2(n10848), .B1(n10847), .B2(n7244), .ZN(
        P2_U3429) );
  INV_X1 U11421 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10849) );
  AOI22_X1 U11422 ( .A1(n10851), .A2(n10850), .B1(n10849), .B2(n7244), .ZN(
        P2_U3432) );
  XNOR2_X1 U11423 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  NAND2_X1 U6454 ( .A1(n5543), .A2(n5542), .ZN(n9119) );
  INV_X1 U5040 ( .A(n6966), .ZN(n6983) );
  CLKBUF_X1 U5046 ( .A(n9646), .Z(n4956) );
  NAND2_X1 U5081 ( .A1(n7262), .A2(n9369), .ZN(n9269) );
  CLKBUF_X1 U5089 ( .A(n6273), .Z(n6594) );
  CLKBUF_X2 U5232 ( .A(n6269), .Z(n6595) );
  OR2_X1 U5245 ( .A1(n6240), .A2(n6224), .ZN(n5354) );
  CLKBUF_X2 U6257 ( .A(n6959), .Z(n7165) );
  CLKBUF_X1 U6400 ( .A(n6115), .Z(n4966) );
endmodule

