

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, 
        keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, 
        keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, 
        keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, 
        keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, 
        keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, 
        keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, 
        keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, 
        keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, 
        keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, 
        keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2004, n2006, n2007, n2008, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597;

  INV_X2 U2247 ( .A(n2029), .ZN(n2743) );
  NAND2_X4 U2248 ( .A1(n2866), .A2(n2225), .ZN(n2355) );
  INV_X1 U2249 ( .A(n2004), .ZN(n2007) );
  INV_X1 U2250 ( .A(n2239), .ZN(n2225) );
  NAND4_X1 U2251 ( .A1(n2054), .A2(n2055), .A3(n2051), .A4(n2218), .ZN(n2573)
         );
  INV_X1 U2252 ( .A(n2004), .ZN(n2008) );
  INV_X1 U2253 ( .A(IR_REG_31__SCAN_IN), .ZN(n2869) );
  INV_X1 U2254 ( .A(n2224), .ZN(n2866) );
  XNOR2_X2 U2255 ( .A(n2222), .B(n2221), .ZN(n2224) );
  XNOR2_X2 U2256 ( .A(n2068), .B(IR_REG_29__SCAN_IN), .ZN(n2239) );
  MUX2_X1 U2257 ( .A(REG0_REG_28__SCAN_IN), .B(n2611), .S(n4431), .Z(n2612) );
  MUX2_X1 U2258 ( .A(REG1_REG_28__SCAN_IN), .B(n2611), .S(n4443), .Z(n2604) );
  INV_X4 U2259 ( .A(n2799), .ZN(n2810) );
  INV_X2 U2260 ( .A(n2829), .ZN(n2805) );
  INV_X1 U2261 ( .A(n2627), .ZN(n2166) );
  CLKBUF_X2 U2262 ( .A(n2627), .Z(n3813) );
  INV_X1 U2263 ( .A(n2254), .ZN(n3105) );
  INV_X4 U2264 ( .A(n2813), .ZN(n2829) );
  INV_X1 U2265 ( .A(n3569), .ZN(n3091) );
  NAND4_X1 U2266 ( .A1(n2272), .A2(n2271), .A3(n2270), .A4(n2269), .ZN(n3569)
         );
  NAND4_X1 U2267 ( .A1(n2244), .A2(n2243), .A3(n2242), .A4(n2241), .ZN(n2627)
         );
  INV_X4 U2268 ( .A(n2812), .ZN(n2628) );
  CLKBUF_X2 U2269 ( .A(n2248), .Z(n2006) );
  INV_X1 U2270 ( .A(n2248), .ZN(n2004) );
  NAND2_X2 U2271 ( .A1(n2233), .A2(n2232), .ZN(n2326) );
  NAND2_X1 U2272 ( .A1(n3470), .A2(n2780), .ZN(n3472) );
  NAND2_X1 U2273 ( .A1(n3490), .A2(n2012), .ZN(n2129) );
  NAND2_X1 U2274 ( .A1(n2761), .A2(n2012), .ZN(n2132) );
  OR2_X1 U2275 ( .A1(n3491), .A2(n3493), .ZN(n3490) );
  XNOR2_X1 U2276 ( .A(n3883), .B(n3882), .ZN(n4339) );
  AND2_X1 U2277 ( .A1(n3881), .A2(n3880), .ZN(n3883) );
  OR2_X1 U2278 ( .A1(n3866), .A2(n3865), .ZN(n3881) );
  AND2_X1 U2279 ( .A1(n2102), .A2(n2020), .ZN(n3866) );
  OR2_X1 U2280 ( .A1(n4117), .A2(n2444), .ZN(n2195) );
  AND2_X1 U2281 ( .A1(n4115), .A2(n4114), .ZN(n4117) );
  AND2_X1 U2282 ( .A1(n3862), .A2(n3861), .ZN(n3863) );
  OR2_X1 U2283 ( .A1(n3307), .A2(n3306), .ZN(n3862) );
  AND2_X1 U2284 ( .A1(n2021), .A2(n2093), .ZN(n3307) );
  NAND2_X1 U2285 ( .A1(n4317), .A2(n3297), .ZN(n3852) );
  NAND2_X1 U2286 ( .A1(n3949), .A2(n3907), .ZN(n3908) );
  AND2_X1 U2287 ( .A1(n2103), .A2(n2026), .ZN(n4304) );
  AOI21_X1 U2288 ( .B1(n2135), .B2(n2139), .A(n2023), .ZN(n2134) );
  OR2_X1 U2289 ( .A1(n3202), .A2(n3201), .ZN(n2137) );
  NAND2_X2 U2290 ( .A1(n3675), .A2(n2533), .ZN(n3755) );
  XNOR2_X1 U2291 ( .A(n2934), .B(n2923), .ZN(n2935) );
  NAND2_X1 U2292 ( .A1(n2285), .A2(n2284), .ZN(n3812) );
  NAND3_X1 U2293 ( .A1(n2238), .A2(n2237), .A3(n2236), .ZN(n3814) );
  AND2_X2 U2294 ( .A1(n2628), .A2(n4424), .ZN(n2799) );
  OR2_X1 U2295 ( .A1(n2355), .A2(n2887), .ZN(n2241) );
  INV_X1 U2296 ( .A(n2624), .ZN(n3047) );
  NAND2_X2 U2297 ( .A1(n2584), .A2(n2583), .ZN(n2615) );
  XNOR2_X1 U2298 ( .A(n2578), .B(IR_REG_24__SCAN_IN), .ZN(n2584) );
  MUX2_X1 U2299 ( .A(IR_REG_31__SCAN_IN), .B(n2523), .S(IR_REG_21__SCAN_IN), 
        .Z(n2526) );
  XNOR2_X1 U2300 ( .A(n2531), .B(n2575), .ZN(n2623) );
  NAND2_X1 U2301 ( .A1(n2581), .A2(n2019), .ZN(n2601) );
  XNOR2_X1 U2302 ( .A(n2527), .B(IR_REG_19__SCAN_IN), .ZN(n4277) );
  OR2_X1 U2303 ( .A1(n2576), .A2(n2869), .ZN(n2531) );
  OR2_X1 U2304 ( .A1(n2574), .A2(n2188), .ZN(n2860) );
  NOR2_X1 U2305 ( .A1(n2382), .A2(n2186), .ZN(n2428) );
  NOR2_X1 U2306 ( .A1(n2052), .A2(n2261), .ZN(n2051) );
  OAI211_X1 U2307 ( .C1(IR_REG_31__SCAN_IN), .C2(IR_REG_1__SCAN_IN), .A(n2155), 
        .B(n2246), .ZN(n2886) );
  INV_X1 U2308 ( .A(n2383), .ZN(n2055) );
  NOR2_X1 U2309 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2210)
         );
  NOR2_X1 U2310 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2208)
         );
  NOR2_X1 U2311 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2209)
         );
  NOR2_X1 U2312 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2207)
         );
  INV_X1 U2313 ( .A(IR_REG_13__SCAN_IN), .ZN(n2385) );
  NOR2_X2 U2314 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2245)
         );
  INV_X1 U2315 ( .A(IR_REG_3__SCAN_IN), .ZN(n2273) );
  INV_X1 U2316 ( .A(IR_REG_25__SCAN_IN), .ZN(n2219) );
  AND2_X4 U2317 ( .A1(n2224), .A2(n2225), .ZN(n2280) );
  AND2_X1 U2318 ( .A1(n2224), .A2(n2239), .ZN(n2248) );
  OAI21_X2 U2319 ( .B1(n3431), .B2(n3427), .A(n3428), .ZN(n3439) );
  NOR2_X1 U2320 ( .A1(n2175), .A2(n2483), .ZN(n2174) );
  INV_X1 U2321 ( .A(n2202), .ZN(n2175) );
  NAND2_X1 U2322 ( .A1(n2530), .A2(n2606), .ZN(n2624) );
  NOR2_X1 U2323 ( .A1(n3223), .A2(n2136), .ZN(n2135) );
  INV_X1 U2324 ( .A(n2137), .ZN(n2136) );
  AOI21_X1 U2325 ( .B1(n3814), .B2(n2829), .A(n2617), .ZN(n2625) );
  NOR2_X1 U2326 ( .A1(n2812), .A2(n2616), .ZN(n2617) );
  NAND2_X1 U2327 ( .A1(n2239), .A2(REG3_REG_1__SCAN_IN), .ZN(n2240) );
  NAND2_X1 U2328 ( .A1(n2153), .A2(n2524), .ZN(n2152) );
  INV_X1 U2329 ( .A(IR_REG_21__SCAN_IN), .ZN(n2524) );
  INV_X1 U2330 ( .A(n2521), .ZN(n2153) );
  AND2_X1 U2331 ( .A1(n3202), .A2(n3201), .ZN(n2139) );
  AOI21_X1 U2332 ( .B1(n3281), .B2(n3282), .A(n2683), .ZN(n3481) );
  OR2_X1 U2333 ( .A1(n2485), .A2(n2484), .ZN(n2494) );
  NOR2_X1 U2334 ( .A1(n2789), .A2(n2788), .ZN(n2790) );
  NAND2_X2 U2335 ( .A1(n2615), .A2(n2624), .ZN(n2812) );
  NAND2_X1 U2336 ( .A1(n2882), .A2(IR_REG_28__SCAN_IN), .ZN(n2232) );
  NAND2_X1 U2337 ( .A1(n2158), .A2(n2157), .ZN(n3874) );
  INV_X1 U2338 ( .A(n3859), .ZN(n2157) );
  AOI21_X1 U2339 ( .B1(n2170), .B2(n2171), .A(n2169), .ZN(n2168) );
  NOR2_X1 U2340 ( .A1(n3960), .A2(n3984), .ZN(n2169) );
  NAND2_X1 U2341 ( .A1(n2468), .A2(REG3_REG_23__SCAN_IN), .ZN(n2485) );
  AOI21_X1 U2342 ( .B1(n4069), .B2(n2454), .A(n2453), .ZN(n4049) );
  OR2_X1 U2343 ( .A1(n4101), .A2(n4081), .ZN(n2454) );
  NOR2_X1 U2344 ( .A1(n4054), .A2(n3765), .ZN(n2453) );
  AND2_X1 U2345 ( .A1(n2821), .A2(n2873), .ZN(n3042) );
  AND2_X1 U2346 ( .A1(n2623), .A2(n3788), .ZN(n2607) );
  NAND2_X1 U2347 ( .A1(n2607), .A2(n2606), .ZN(n4424) );
  OR2_X1 U2348 ( .A1(n4070), .A2(n2551), .ZN(n3719) );
  INV_X1 U2349 ( .A(n3085), .ZN(n2179) );
  AND2_X1 U2350 ( .A1(n3091), .A2(n3158), .ZN(n2291) );
  NAND2_X1 U2351 ( .A1(n2520), .A2(n2519), .ZN(n2521) );
  INV_X1 U2352 ( .A(n3811), .ZN(n2665) );
  NAND2_X1 U2353 ( .A1(n2060), .A2(n3400), .ZN(n2058) );
  AND2_X1 U2354 ( .A1(n2061), .A2(n3713), .ZN(n2060) );
  INV_X1 U2355 ( .A(n3715), .ZN(n2061) );
  AOI21_X1 U2356 ( .B1(n3751), .B2(n2363), .A(n2018), .ZN(n2183) );
  INV_X1 U2357 ( .A(n3484), .ZN(n2695) );
  AND2_X1 U2358 ( .A1(n3109), .A2(n2636), .ZN(n2076) );
  INV_X1 U2359 ( .A(n3103), .ZN(n3109) );
  AND2_X1 U2360 ( .A1(n3814), .A2(n3015), .ZN(n2965) );
  NAND2_X1 U2361 ( .A1(n3755), .A2(n2965), .ZN(n2967) );
  INV_X1 U2362 ( .A(IR_REG_26__SCAN_IN), .ZN(n2192) );
  INV_X1 U2363 ( .A(IR_REG_27__SCAN_IN), .ZN(n2220) );
  NAND2_X1 U2364 ( .A1(n2024), .A2(n2213), .ZN(n2186) );
  INV_X1 U2365 ( .A(IR_REG_6__SCAN_IN), .ZN(n2310) );
  INV_X1 U2366 ( .A(IR_REG_2__SCAN_IN), .ZN(n2211) );
  AOI21_X1 U2367 ( .B1(n3597), .B2(n3599), .A(n3598), .ZN(n3492) );
  XNOR2_X1 U2368 ( .A(n2633), .B(n2634), .ZN(n3020) );
  INV_X1 U2369 ( .A(n2671), .ZN(n2141) );
  NAND2_X1 U2370 ( .A1(n3200), .A2(n2135), .ZN(n2133) );
  OR2_X1 U2371 ( .A1(n2615), .A2(n2618), .ZN(n2196) );
  INV_X1 U2372 ( .A(n3575), .ZN(n3576) );
  NOR2_X1 U2373 ( .A1(n3589), .A2(n2131), .ZN(n2130) );
  INV_X1 U2374 ( .A(n3502), .ZN(n2131) );
  OAI22_X1 U2375 ( .A1(n2665), .A2(n2810), .B1(n2805), .B2(n2664), .ZN(n3201)
         );
  AND2_X1 U2376 ( .A1(n2822), .A2(n3042), .ZN(n2833) );
  OR2_X1 U2377 ( .A1(n2355), .A2(n2942), .ZN(n2235) );
  NAND2_X1 U2378 ( .A1(n2083), .A2(n2885), .ZN(n2906) );
  NAND2_X1 U2379 ( .A1(n2935), .A2(n2161), .ZN(n2159) );
  NOR2_X1 U2380 ( .A1(n2936), .A2(n2294), .ZN(n2161) );
  NAND2_X1 U2381 ( .A1(n2164), .A2(n2163), .ZN(n2162) );
  INV_X1 U2382 ( .A(n2936), .ZN(n2163) );
  INV_X1 U2383 ( .A(n2165), .ZN(n2164) );
  NAND2_X1 U2384 ( .A1(n3839), .A2(n2913), .ZN(n2929) );
  OAI21_X1 U2385 ( .B1(n2953), .B2(n2952), .A(n2954), .ZN(n3000) );
  NAND2_X1 U2386 ( .A1(n3291), .A2(n2034), .ZN(n3293) );
  NOR2_X1 U2387 ( .A1(n3301), .A2(n2104), .ZN(n3302) );
  AND2_X1 U2388 ( .A1(n4279), .A2(REG1_REG_9__SCAN_IN), .ZN(n2104) );
  AND2_X1 U2389 ( .A1(n3874), .A2(n3873), .ZN(n3875) );
  NAND2_X1 U2390 ( .A1(n2072), .A2(n2070), .ZN(n2069) );
  NOR2_X1 U2391 ( .A1(n3907), .A2(n3915), .ZN(n2072) );
  INV_X1 U2392 ( .A(n2071), .ZN(n2070) );
  INV_X1 U2393 ( .A(n2174), .ZN(n2173) );
  AOI21_X1 U2394 ( .B1(n2174), .B2(n2172), .A(n2039), .ZN(n2171) );
  INV_X1 U2395 ( .A(n2475), .ZN(n2172) );
  NAND2_X1 U2396 ( .A1(n2474), .A2(n4014), .ZN(n2475) );
  AND2_X1 U2397 ( .A1(n2455), .A2(REG3_REG_21__SCAN_IN), .ZN(n2461) );
  NAND2_X1 U2398 ( .A1(n4130), .A2(n3497), .ZN(n2194) );
  AND2_X1 U2399 ( .A1(n2445), .A2(n4105), .ZN(n2193) );
  OR2_X1 U2400 ( .A1(n2436), .A2(n2205), .ZN(n2447) );
  AND4_X1 U2401 ( .A1(n2427), .A2(n2426), .A3(n2425), .A4(n2424), .ZN(n4134)
         );
  NOR2_X1 U2402 ( .A1(n3624), .A2(n3463), .ZN(n2079) );
  INV_X1 U2403 ( .A(n3638), .ZN(n2048) );
  NAND2_X1 U2404 ( .A1(n2185), .A2(n2184), .ZN(n3335) );
  AOI21_X1 U2405 ( .B1(n2065), .B2(n2064), .A(n2063), .ZN(n2062) );
  INV_X1 U2406 ( .A(n3700), .ZN(n2064) );
  OAI21_X1 U2407 ( .B1(n3129), .B2(n2539), .A(n3696), .ZN(n3192) );
  OAI21_X1 U2408 ( .B1(n3118), .B2(n2537), .A(n3687), .ZN(n3152) );
  OR2_X1 U2409 ( .A1(n2530), .A2(n4425), .ZN(n2835) );
  NAND2_X1 U2410 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2279) );
  INV_X1 U2411 ( .A(n3567), .ZN(n3069) );
  AOI21_X1 U2412 ( .B1(n2049), .B2(n4126), .A(n3919), .ZN(n4175) );
  XNOR2_X1 U2413 ( .A(n2050), .B(n2032), .ZN(n2049) );
  NOR2_X1 U2414 ( .A1(n3983), .A2(n2071), .ZN(n3938) );
  AND2_X1 U2415 ( .A1(n3938), .A2(n2811), .ZN(n3922) );
  NOR2_X1 U2416 ( .A1(n3365), .A2(n2078), .ZN(n4150) );
  NAND2_X1 U2417 ( .A1(n2730), .A2(n2079), .ZN(n2078) );
  INV_X1 U2418 ( .A(n3444), .ZN(n3366) );
  NOR2_X1 U2419 ( .A1(n3343), .A2(n3432), .ZN(n3367) );
  NAND2_X1 U2420 ( .A1(n2582), .A2(n2857), .ZN(n2872) );
  OR2_X1 U2421 ( .A1(n2573), .A2(n2189), .ZN(n2562) );
  NAND2_X1 U2422 ( .A1(n2220), .A2(n2192), .ZN(n2189) );
  INV_X1 U2423 ( .A(n2186), .ZN(n2054) );
  NOR2_X1 U2424 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_21__SCAN_IN), .ZN(n2216)
         );
  NOR2_X1 U2425 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2215)
         );
  NAND2_X1 U2426 ( .A1(n2151), .A2(n2575), .ZN(n2150) );
  INV_X1 U2427 ( .A(n2152), .ZN(n2151) );
  INV_X1 U2428 ( .A(IR_REG_23__SCAN_IN), .ZN(n2586) );
  XNOR2_X1 U2429 ( .A(n2585), .B(n2586), .ZN(n2877) );
  XNOR2_X1 U2430 ( .A(n2529), .B(n2519), .ZN(n2606) );
  NAND2_X1 U2431 ( .A1(n2528), .A2(IR_REG_31__SCAN_IN), .ZN(n2529) );
  NAND2_X1 U2432 ( .A1(n2522), .A2(IR_REG_31__SCAN_IN), .ZN(n2527) );
  INV_X1 U2433 ( .A(IR_REG_16__SCAN_IN), .ZN(n4580) );
  NOR2_X1 U2434 ( .A1(n2341), .A2(IR_REG_9__SCAN_IN), .ZN(n2361) );
  NOR2_X1 U2435 ( .A1(n2384), .A2(IR_REG_5__SCAN_IN), .ZN(n2311) );
  NAND2_X1 U2436 ( .A1(n2142), .A2(n2145), .ZN(n3431) );
  AND2_X1 U2437 ( .A1(n2147), .A2(n2146), .ZN(n2145) );
  OR2_X1 U2438 ( .A1(n2692), .A2(n2697), .ZN(n2146) );
  AND2_X1 U2439 ( .A1(n2486), .A2(n2494), .ZN(n3986) );
  XNOR2_X1 U2440 ( .A(n3293), .B(n4388), .ZN(n4299) );
  NAND2_X1 U2441 ( .A1(n4299), .A2(REG2_REG_10__SCAN_IN), .ZN(n4298) );
  XNOR2_X1 U2442 ( .A(n3875), .B(n3882), .ZN(n4336) );
  NAND2_X1 U2443 ( .A1(n4347), .A2(n4348), .ZN(n4346) );
  NAND2_X1 U2444 ( .A1(n3886), .A2(n3887), .ZN(n2111) );
  NOR2_X1 U2445 ( .A1(n2108), .A2(n2106), .ZN(n2105) );
  INV_X1 U2446 ( .A(n2107), .ZN(n2106) );
  NOR2_X1 U2447 ( .A1(n4358), .A2(n3890), .ZN(n2108) );
  AOI21_X1 U2448 ( .B1(n4345), .B2(ADDR_REG_18__SCAN_IN), .A(n3888), .ZN(n2107) );
  NOR2_X1 U2449 ( .A1(n3886), .A2(n3887), .ZN(n3891) );
  OAI21_X1 U2450 ( .B1(n3922), .B2(n3921), .A(n2030), .ZN(n4174) );
  AND2_X1 U2451 ( .A1(n2173), .A2(n2016), .ZN(n2170) );
  OAI21_X1 U2452 ( .B1(n3914), .B2(n3913), .A(n3912), .ZN(n2050) );
  NAND2_X1 U2453 ( .A1(n3965), .A2(n3946), .ZN(n2071) );
  AND2_X1 U2454 ( .A1(n3178), .A2(n3193), .ZN(n2081) );
  INV_X1 U2455 ( .A(n2301), .ZN(n2177) );
  NAND2_X1 U2456 ( .A1(n2179), .A2(n2301), .ZN(n2178) );
  NOR2_X1 U2457 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2214)
         );
  INV_X1 U2458 ( .A(IR_REG_22__SCAN_IN), .ZN(n2575) );
  AND2_X1 U2459 ( .A1(n2123), .A2(n2033), .ZN(n2121) );
  NAND2_X1 U2460 ( .A1(n3607), .A2(n2124), .ZN(n2123) );
  INV_X1 U2461 ( .A(n2127), .ZN(n2124) );
  NOR2_X1 U2462 ( .A1(n2809), .A2(n2126), .ZN(n2120) );
  NAND2_X1 U2463 ( .A1(n2119), .A2(n2118), .ZN(n2117) );
  INV_X1 U2464 ( .A(n2809), .ZN(n2118) );
  NAND2_X1 U2465 ( .A1(n3451), .A2(n2121), .ZN(n2119) );
  INV_X1 U2466 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2316) );
  NOR2_X1 U2467 ( .A1(n2144), .A2(n2036), .ZN(n2143) );
  INV_X1 U2468 ( .A(n3480), .ZN(n2144) );
  OR2_X1 U2469 ( .A1(n2149), .A2(n2148), .ZN(n2147) );
  INV_X1 U2470 ( .A(n3386), .ZN(n2148) );
  AND2_X1 U2471 ( .A1(n2692), .A2(n2697), .ZN(n2149) );
  AND2_X1 U2472 ( .A1(n2733), .A2(n2732), .ZN(n2737) );
  NOR2_X1 U2473 ( .A1(n2365), .A2(n2364), .ZN(n2376) );
  NAND2_X1 U2474 ( .A1(n3481), .A2(n3480), .ZN(n3479) );
  INV_X1 U2475 ( .A(n3543), .ZN(n2113) );
  NAND2_X1 U2476 ( .A1(n2038), .A2(n2128), .ZN(n2127) );
  AND3_X1 U2477 ( .A1(n2162), .A2(n2159), .A3(n2042), .ZN(n2996) );
  OR2_X1 U2478 ( .A1(n4295), .A2(n4491), .ZN(n2103) );
  NAND2_X1 U2479 ( .A1(n2088), .A2(n2084), .ZN(n2093) );
  AND2_X1 U2480 ( .A1(n2089), .A2(n2086), .ZN(n2084) );
  NOR2_X1 U2481 ( .A1(n2087), .A2(n4502), .ZN(n2086) );
  INV_X1 U2482 ( .A(n2090), .ZN(n2087) );
  NAND2_X1 U2483 ( .A1(n4444), .A2(n2092), .ZN(n2090) );
  OR2_X1 U2484 ( .A1(n4302), .A2(n2091), .ZN(n2088) );
  NAND2_X1 U2485 ( .A1(n2156), .A2(n2094), .ZN(n2091) );
  NAND2_X1 U2486 ( .A1(n4307), .A2(n3295), .ZN(n3296) );
  NOR2_X1 U2487 ( .A1(n2101), .A2(n4501), .ZN(n2096) );
  OR2_X1 U2488 ( .A1(n3862), .A2(n4385), .ZN(n2097) );
  NAND2_X1 U2489 ( .A1(n3862), .A2(n2098), .ZN(n2095) );
  NOR2_X1 U2490 ( .A1(n2099), .A2(n4329), .ZN(n2098) );
  INV_X1 U2491 ( .A(n3861), .ZN(n2099) );
  OR2_X1 U2492 ( .A1(n4325), .A2(n3856), .ZN(n2158) );
  NAND2_X1 U2493 ( .A1(n4346), .A2(n2154), .ZN(n3877) );
  NAND2_X1 U2494 ( .A1(n4382), .A2(n4550), .ZN(n2154) );
  NOR2_X1 U2495 ( .A1(n3877), .A2(n3878), .ZN(n3894) );
  NOR2_X1 U2496 ( .A1(n2030), .A2(n4171), .ZN(n4168) );
  NOR2_X1 U2497 ( .A1(n4083), .A2(n4059), .ZN(n2082) );
  OAI21_X1 U2498 ( .B1(n3405), .B2(n2059), .A(n2057), .ZN(n2553) );
  INV_X1 U2499 ( .A(n2060), .ZN(n2059) );
  AND2_X1 U2500 ( .A1(n2552), .A2(n2058), .ZN(n2057) );
  NAND2_X1 U2501 ( .A1(n3404), .A2(n2060), .ZN(n4072) );
  OR2_X1 U2502 ( .A1(n2434), .A2(n2433), .ZN(n2436) );
  NAND2_X1 U2503 ( .A1(n3404), .A2(n3713), .ZN(n4142) );
  AND4_X1 U2504 ( .A1(n2440), .A2(n2439), .A3(n2438), .A4(n2437), .ZN(n4141)
         );
  AND2_X1 U2505 ( .A1(n3756), .A2(n4093), .ZN(n4158) );
  NAND2_X1 U2506 ( .A1(n3405), .A2(n3760), .ZN(n3404) );
  INV_X1 U2507 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3622) );
  OR2_X1 U2508 ( .A1(n2396), .A2(n3622), .ZN(n2407) );
  INV_X1 U2509 ( .A(n3805), .ZN(n3381) );
  NAND2_X1 U2510 ( .A1(n2047), .A2(n2013), .ZN(n3378) );
  AND2_X1 U2511 ( .A1(n2376), .A2(REG3_REG_13__SCAN_IN), .ZN(n2389) );
  NAND2_X1 U2512 ( .A1(n2546), .A2(n3708), .ZN(n3644) );
  AND2_X1 U2513 ( .A1(n3638), .A2(n3640), .ZN(n3747) );
  AOI21_X1 U2514 ( .B1(n2183), .B2(n2181), .A(n2037), .ZN(n2180) );
  INV_X1 U2515 ( .A(n2183), .ZN(n2182) );
  INV_X1 U2516 ( .A(n2363), .ZN(n2181) );
  AND2_X1 U2517 ( .A1(n3254), .A2(n3256), .ZN(n3751) );
  OR2_X1 U2518 ( .A1(n2317), .A2(n2316), .ZN(n2331) );
  NOR2_X1 U2519 ( .A1(n2331), .A2(n4461), .ZN(n2345) );
  INV_X1 U2520 ( .A(REG3_REG_9__SCAN_IN), .ZN(n4461) );
  NAND2_X1 U2521 ( .A1(n3192), .A2(n3699), .ZN(n2540) );
  INV_X1 U2522 ( .A(n3284), .ZN(n3178) );
  INV_X1 U2523 ( .A(n3482), .ZN(n3234) );
  INV_X1 U2524 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2302) );
  OR2_X1 U2525 ( .A1(n2303), .A2(n2302), .ZN(n2317) );
  INV_X1 U2526 ( .A(n4170), .ZN(n4139) );
  NAND2_X1 U2527 ( .A1(n2538), .A2(n3693), .ZN(n3129) );
  INV_X1 U2528 ( .A(n4133), .ZN(n4148) );
  OAI21_X1 U2529 ( .B1(n3152), .B2(n3148), .A(n3691), .ZN(n3089) );
  INV_X1 U2530 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2267) );
  INV_X1 U2531 ( .A(n4140), .ZN(n4129) );
  NAND2_X1 U2532 ( .A1(n2536), .A2(n3683), .ZN(n3118) );
  INV_X1 U2533 ( .A(n3117), .ZN(n3750) );
  AND2_X1 U2534 ( .A1(n2073), .A2(n2076), .ZN(n3159) );
  NOR2_X1 U2535 ( .A1(n3074), .A2(n3568), .ZN(n2073) );
  NAND2_X1 U2536 ( .A1(n2075), .A2(n2076), .ZN(n3116) );
  AND2_X1 U2537 ( .A1(n3683), .A2(n3680), .ZN(n3757) );
  INV_X1 U2538 ( .A(n3025), .ZN(n2974) );
  NAND2_X1 U2539 ( .A1(n3670), .A2(n2561), .ZN(n4126) );
  AND2_X1 U2540 ( .A1(n2607), .A2(n3790), .ZN(n4170) );
  OR2_X1 U2541 ( .A1(n4000), .A2(n3978), .ZN(n3983) );
  NAND2_X1 U2542 ( .A1(n4020), .A2(n4001), .ZN(n4000) );
  NOR2_X1 U2543 ( .A1(n4199), .A2(n4021), .ZN(n4020) );
  INV_X1 U2544 ( .A(n2082), .ZN(n4061) );
  NOR2_X1 U2545 ( .A1(n2326), .A2(n2452), .ZN(n4081) );
  OR2_X1 U2546 ( .A1(n4104), .A2(n4081), .ZN(n4083) );
  NOR2_X1 U2547 ( .A1(n4152), .A2(n4128), .ZN(n4106) );
  INV_X1 U2548 ( .A(n3497), .ZN(n4105) );
  NAND2_X1 U2549 ( .A1(n4150), .A2(n4149), .ZN(n4152) );
  OR2_X1 U2550 ( .A1(n3342), .A2(n3389), .ZN(n3343) );
  NAND2_X1 U2551 ( .A1(n3187), .A2(n2080), .ZN(n3342) );
  AND2_X1 U2552 ( .A1(n2081), .A2(n2687), .ZN(n2080) );
  NAND2_X1 U2553 ( .A1(n3187), .A2(n2081), .ZN(n3237) );
  NOR2_X1 U2554 ( .A1(n3136), .A2(n3225), .ZN(n3187) );
  AND2_X1 U2555 ( .A1(n3187), .A2(n3193), .ZN(n3188) );
  NOR2_X1 U2556 ( .A1(n3568), .A2(n3537), .ZN(n2074) );
  OR2_X1 U2557 ( .A1(n3161), .A2(n3205), .ZN(n3136) );
  INV_X1 U2558 ( .A(n4417), .ZN(n4411) );
  NOR2_X1 U2559 ( .A1(n3074), .A2(n3073), .ZN(n3110) );
  NAND2_X1 U2560 ( .A1(n2967), .A2(n2247), .ZN(n3065) );
  AND3_X1 U2561 ( .A1(n2600), .A2(n2599), .A3(n2598), .ZN(n2610) );
  INV_X1 U2562 ( .A(IR_REG_30__SCAN_IN), .ZN(n2221) );
  NAND2_X1 U2563 ( .A1(n2870), .A2(IR_REG_31__SCAN_IN), .ZN(n2222) );
  NAND2_X1 U2564 ( .A1(n2562), .A2(n2230), .ZN(n2883) );
  AND2_X1 U2565 ( .A1(n2019), .A2(n2231), .ZN(n2882) );
  AND2_X1 U2566 ( .A1(IR_REG_27__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2231)
         );
  INV_X1 U2567 ( .A(n2576), .ZN(n2525) );
  NAND2_X1 U2568 ( .A1(n2017), .A2(IR_REG_31__SCAN_IN), .ZN(n2523) );
  INV_X1 U2569 ( .A(IR_REG_17__SCAN_IN), .ZN(n2228) );
  INV_X1 U2570 ( .A(IR_REG_15__SCAN_IN), .ZN(n2403) );
  INV_X1 U2571 ( .A(IR_REG_8__SCAN_IN), .ZN(n2324) );
  OR2_X1 U2572 ( .A1(n2261), .A2(n2275), .ZN(n2384) );
  OR2_X1 U2573 ( .A1(n3200), .A2(n2139), .ZN(n2138) );
  CLKBUF_X1 U2574 ( .A(n3459), .Z(n3460) );
  AND2_X1 U2575 ( .A1(n3473), .A2(n3471), .ZN(n2780) );
  INV_X1 U2576 ( .A(n4053), .ZN(n4059) );
  OAI21_X1 U2577 ( .B1(n2761), .B2(n3490), .A(n2760), .ZN(n3508) );
  NAND2_X1 U2578 ( .A1(n2792), .A2(n3554), .ZN(n3515) );
  NAND2_X1 U2579 ( .A1(n2133), .A2(n2011), .ZN(n2140) );
  AND2_X1 U2580 ( .A1(n2833), .A2(n2830), .ZN(n3626) );
  INV_X1 U2581 ( .A(n2640), .ZN(n2638) );
  AND2_X1 U2582 ( .A1(n2633), .A2(n2634), .ZN(n2635) );
  AND2_X1 U2583 ( .A1(n2492), .A2(n2491), .ZN(n3960) );
  INV_X1 U2584 ( .A(n3623), .ZN(n3610) );
  AND2_X1 U2585 ( .A1(n2833), .A2(n2824), .ZN(n3632) );
  AND2_X1 U2586 ( .A1(n2843), .A2(n3010), .ZN(n3630) );
  OAI21_X1 U2587 ( .B1(n3941), .B2(n2398), .A(n2507), .ZN(n3962) );
  NAND2_X1 U2588 ( .A1(n2481), .A2(n2480), .ZN(n4017) );
  OAI21_X1 U2589 ( .B1(n4062), .B2(n2398), .A(n2460), .ZN(n4037) );
  OAI211_X1 U2590 ( .C1(n2355), .C2(n4085), .A(n2451), .B(n2450), .ZN(n4101)
         );
  OAI211_X1 U2591 ( .C1(n4108), .C2(n2398), .A(n2227), .B(n2226), .ZN(n4130)
         );
  INV_X1 U2592 ( .A(n4134), .ZN(n3803) );
  NOR2_X1 U2593 ( .A1(n2204), .A2(n2283), .ZN(n2284) );
  NAND4_X1 U2594 ( .A1(n2260), .A2(n2259), .A3(n2258), .A4(n2257), .ZN(n3567)
         );
  OR2_X1 U2595 ( .A1(n2398), .A2(n3018), .ZN(n2236) );
  NAND2_X1 U2596 ( .A1(n2280), .A2(REG0_REG_0__SCAN_IN), .ZN(n2237) );
  NAND2_X1 U2597 ( .A1(n3815), .A2(n3816), .ZN(n3830) );
  XNOR2_X1 U2598 ( .A(n2906), .B(n2896), .ZN(n2905) );
  AND2_X1 U2599 ( .A1(n2160), .A2(n2165), .ZN(n2937) );
  NAND2_X1 U2600 ( .A1(n2159), .A2(n2162), .ZN(n2950) );
  NAND2_X1 U2601 ( .A1(n2935), .A2(REG2_REG_6__SCAN_IN), .ZN(n2160) );
  NAND2_X1 U2602 ( .A1(n2931), .A2(n2930), .ZN(n2953) );
  XNOR2_X1 U2603 ( .A(n3000), .B(n3001), .ZN(n2955) );
  XNOR2_X1 U2604 ( .A(n3302), .B(n4388), .ZN(n4295) );
  INV_X1 U2605 ( .A(n2103), .ZN(n4294) );
  NAND2_X1 U2606 ( .A1(n4298), .A2(n3294), .ZN(n4308) );
  XNOR2_X1 U2607 ( .A(n3296), .B(n2156), .ZN(n4318) );
  NAND2_X1 U2608 ( .A1(n4318), .A2(REG2_REG_12__SCAN_IN), .ZN(n4317) );
  INV_X1 U2609 ( .A(n2158), .ZN(n3858) );
  NAND2_X1 U2610 ( .A1(n4335), .A2(n3876), .ZN(n4347) );
  AND2_X1 U2611 ( .A1(n2881), .A2(n2879), .ZN(n4345) );
  AND2_X1 U2612 ( .A1(n2945), .A2(n3796), .ZN(n4355) );
  OAI21_X1 U2613 ( .B1(n4007), .B2(n2173), .A(n2171), .ZN(n3972) );
  NAND2_X1 U2614 ( .A1(n4007), .A2(n2475), .ZN(n2176) );
  NAND2_X1 U2615 ( .A1(n2082), .A2(n3590), .ZN(n4199) );
  INV_X1 U2616 ( .A(n2195), .ZN(n4091) );
  INV_X1 U2617 ( .A(n2079), .ZN(n2077) );
  NAND2_X1 U2618 ( .A1(n3335), .A2(n2363), .ZN(n3267) );
  OR2_X2 U2619 ( .A1(n3011), .A2(n2835), .ZN(n4153) );
  INV_X1 U2620 ( .A(n4277), .ZN(n3900) );
  AND2_X2 U2621 ( .A1(n2610), .A2(n2822), .ZN(n4443) );
  AND2_X1 U2622 ( .A1(n4175), .A2(n4176), .ZN(n2200) );
  OR2_X1 U2623 ( .A1(n4174), .A2(n4424), .ZN(n4176) );
  AND2_X2 U2624 ( .A1(n2610), .A2(n3043), .ZN(n4431) );
  NAND2_X1 U2625 ( .A1(n2188), .A2(n2187), .ZN(n2870) );
  NOR2_X1 U2626 ( .A1(n2190), .A2(IR_REG_29__SCAN_IN), .ZN(n2187) );
  OR2_X1 U2627 ( .A1(n2223), .A2(n2869), .ZN(n2068) );
  INV_X1 U2628 ( .A(n2601), .ZN(n2857) );
  NAND2_X1 U2629 ( .A1(n2577), .A2(IR_REG_31__SCAN_IN), .ZN(n2578) );
  AND2_X1 U2630 ( .A1(n2877), .A2(STATE_REG_SCAN_IN), .ZN(n4380) );
  XNOR2_X1 U2631 ( .A(n2373), .B(IR_REG_11__SCAN_IN), .ZN(n4386) );
  NOR2_X1 U2632 ( .A1(n2342), .A2(n2361), .ZN(n4279) );
  AND2_X1 U2633 ( .A1(n2286), .A2(n2263), .ZN(n4285) );
  OR2_X1 U2634 ( .A1(n2245), .A2(n2869), .ZN(n2253) );
  NAND2_X1 U2635 ( .A1(n2109), .A2(n2022), .ZN(U3258) );
  OR2_X1 U2636 ( .A1(n2110), .A2(n3891), .ZN(n2109) );
  NAND2_X1 U2637 ( .A1(n2111), .A2(n4353), .ZN(n2110) );
  OR2_X1 U2638 ( .A1(n3928), .A2(n4271), .ZN(n2613) );
  INV_X1 U2639 ( .A(n2326), .ZN(n2467) );
  AND4_X1 U2640 ( .A1(n2054), .A2(n2056), .A3(n2055), .A4(n2218), .ZN(n2010)
         );
  AND2_X1 U2641 ( .A1(n2134), .A2(n2046), .ZN(n2011) );
  INV_X1 U2642 ( .A(n4444), .ZN(n2156) );
  AND2_X1 U2643 ( .A1(n2760), .A2(n2043), .ZN(n2012) );
  NAND2_X1 U2644 ( .A1(n2056), .A2(n2055), .ZN(n2382) );
  AND2_X1 U2645 ( .A1(n3641), .A2(n3639), .ZN(n2013) );
  OR2_X1 U2646 ( .A1(n2382), .A2(IR_REG_14__SCAN_IN), .ZN(n2014) );
  AND2_X1 U2647 ( .A1(n2041), .A2(n3544), .ZN(n2015) );
  OR2_X1 U2648 ( .A1(n3997), .A2(n3978), .ZN(n2016) );
  OR2_X1 U2649 ( .A1(n2522), .A2(n2521), .ZN(n2017) );
  NAND2_X1 U2650 ( .A1(n2176), .A2(n2202), .ZN(n3991) );
  NAND4_X1 U2651 ( .A1(n2252), .A2(n2251), .A3(n2250), .A4(n2249), .ZN(n2254)
         );
  NAND2_X1 U2652 ( .A1(n2122), .A2(n2127), .ZN(n3606) );
  AND2_X1 U2653 ( .A1(n3807), .A2(n3432), .ZN(n2018) );
  OR2_X1 U2654 ( .A1(n2573), .A2(IR_REG_26__SCAN_IN), .ZN(n2019) );
  OR2_X1 U2655 ( .A1(n3863), .A2(n4385), .ZN(n2020) );
  NAND2_X2 U2656 ( .A1(n2615), .A2(n3047), .ZN(n2813) );
  OR2_X1 U2657 ( .A1(n3304), .A2(n2156), .ZN(n2021) );
  AND2_X1 U2658 ( .A1(n3889), .A2(n2105), .ZN(n2022) );
  INV_X1 U2659 ( .A(n2126), .ZN(n2125) );
  AND2_X1 U2660 ( .A1(n2670), .A2(n2141), .ZN(n2023) );
  AND2_X1 U2661 ( .A1(n4580), .A2(n2403), .ZN(n2024) );
  NAND3_X1 U2662 ( .A1(n2132), .A2(n2129), .A3(n2130), .ZN(n3470) );
  AND2_X1 U2663 ( .A1(n2171), .A2(n2016), .ZN(n2025) );
  OR2_X1 U2664 ( .A1(n3302), .A2(n4388), .ZN(n2026) );
  AND2_X1 U2665 ( .A1(n2116), .A2(n2121), .ZN(n2027) );
  XNOR2_X1 U2666 ( .A(n2631), .B(n2743), .ZN(n2633) );
  NAND2_X1 U2667 ( .A1(n3811), .A2(n3205), .ZN(n2028) );
  AND2_X1 U2668 ( .A1(n2624), .A2(n2826), .ZN(n2029) );
  OAI22_X1 U2669 ( .A1(n3354), .A2(n2388), .B1(n2705), .B2(n3366), .ZN(n3312)
         );
  OR2_X1 U2670 ( .A1(n3983), .A2(n2069), .ZN(n2030) );
  OR2_X1 U2671 ( .A1(n3983), .A2(n2800), .ZN(n2031) );
  INV_X1 U2672 ( .A(IR_REG_19__SCAN_IN), .ZN(n2520) );
  XOR2_X1 U2673 ( .A(n3740), .B(n3921), .Z(n2032) );
  NAND2_X1 U2674 ( .A1(n2112), .A2(n2738), .ZN(n3545) );
  NAND2_X1 U2675 ( .A1(n2114), .A2(n2015), .ZN(n3597) );
  NAND2_X1 U2676 ( .A1(n3479), .A2(n2692), .ZN(n3384) );
  OR2_X1 U2677 ( .A1(n2804), .A2(n2803), .ZN(n2033) );
  INV_X1 U2678 ( .A(IR_REG_20__SCAN_IN), .ZN(n2519) );
  AND2_X1 U2679 ( .A1(n3716), .A2(n3713), .ZN(n3760) );
  INV_X1 U2680 ( .A(IR_REG_28__SCAN_IN), .ZN(n2191) );
  OR2_X1 U2681 ( .A1(n3292), .A2(n3180), .ZN(n2034) );
  NOR2_X1 U2682 ( .A1(n3962), .A2(n3939), .ZN(n2035) );
  NOR2_X1 U2683 ( .A1(n3386), .A2(n3385), .ZN(n2036) );
  AOI21_X1 U2684 ( .B1(n3644), .B2(n3747), .A(n2048), .ZN(n2047) );
  AND2_X1 U2685 ( .A1(n3361), .A2(n3259), .ZN(n2037) );
  INV_X1 U2686 ( .A(n2094), .ZN(n2092) );
  NAND2_X1 U2687 ( .A1(n4386), .A2(REG1_REG_11__SCAN_IN), .ZN(n2094) );
  NOR2_X1 U2688 ( .A1(n2795), .A2(n2794), .ZN(n2038) );
  NOR2_X1 U2689 ( .A1(n4017), .A2(n2482), .ZN(n2039) );
  INV_X1 U2690 ( .A(IR_REG_14__SCAN_IN), .ZN(n2213) );
  AND2_X1 U2691 ( .A1(n3525), .A2(n3543), .ZN(n2040) );
  OR2_X1 U2692 ( .A1(n2738), .A2(n2113), .ZN(n2041) );
  NAND2_X1 U2693 ( .A1(n4280), .A2(REG2_REG_7__SCAN_IN), .ZN(n2042) );
  INV_X1 U2694 ( .A(n2066), .ZN(n2065) );
  NAND2_X1 U2695 ( .A1(n2067), .A2(n3705), .ZN(n2066) );
  AND2_X1 U2696 ( .A1(n3044), .A2(n4153), .ZN(n4377) );
  OAI21_X1 U2697 ( .B1(n2522), .B2(n2150), .A(IR_REG_31__SCAN_IN), .ZN(n2585)
         );
  NAND2_X1 U2698 ( .A1(n2526), .A2(n2525), .ZN(n3788) );
  INV_X1 U2699 ( .A(n3788), .ZN(n2530) );
  INV_X1 U2700 ( .A(n2398), .ZN(n2449) );
  INV_X1 U2701 ( .A(n4014), .ZN(n4021) );
  NAND2_X1 U2702 ( .A1(n2330), .A2(n2329), .ZN(n3182) );
  NAND2_X1 U2703 ( .A1(n3534), .A2(n2663), .ZN(n3200) );
  NAND2_X1 U2704 ( .A1(n2140), .A2(n3271), .ZN(n3281) );
  NAND2_X1 U2705 ( .A1(n2133), .A2(n2134), .ZN(n3270) );
  NAND2_X1 U2706 ( .A1(n2138), .A2(n2137), .ZN(n3222) );
  OR2_X1 U2707 ( .A1(n2768), .A2(n2767), .ZN(n2043) );
  OR2_X1 U2708 ( .A1(n3365), .A2(n3463), .ZN(n2044) );
  INV_X1 U2709 ( .A(n3702), .ZN(n2063) );
  OR2_X1 U2710 ( .A1(n3365), .A2(n2077), .ZN(n2045) );
  AND2_X1 U2711 ( .A1(n2428), .A2(n2228), .ZN(n2441) );
  AND2_X1 U2712 ( .A1(n2945), .A2(n2984), .ZN(n4353) );
  INV_X1 U2713 ( .A(n3074), .ZN(n2075) );
  OR2_X1 U2714 ( .A1(n2677), .A2(n2676), .ZN(n2046) );
  INV_X1 U2715 ( .A(n3590), .ZN(n4042) );
  INV_X1 U2716 ( .A(n3965), .ZN(n2800) );
  INV_X1 U2717 ( .A(n2101), .ZN(n2100) );
  NOR2_X1 U2718 ( .A1(n3861), .A2(n4385), .ZN(n2101) );
  INV_X1 U2719 ( .A(n3885), .ZN(n4382) );
  NOR2_X1 U2720 ( .A1(n2261), .A2(n2212), .ZN(n2056) );
  NAND2_X1 U2721 ( .A1(n2053), .A2(n2219), .ZN(n2052) );
  INV_X1 U2722 ( .A(n2212), .ZN(n2053) );
  OAI21_X1 U2723 ( .B1(n3173), .B2(n2066), .A(n2062), .ZN(n3337) );
  OAI21_X1 U2724 ( .B1(n3173), .B2(n3172), .A(n3700), .ZN(n3232) );
  NAND2_X1 U2725 ( .A1(n3700), .A2(n3172), .ZN(n2067) );
  NAND3_X1 U2726 ( .A1(n2076), .A2(n2075), .A3(n2074), .ZN(n3161) );
  NAND2_X1 U2727 ( .A1(n3367), .A2(n3366), .ZN(n3365) );
  NAND2_X1 U2728 ( .A1(n4106), .A2(n4105), .ZN(n4104) );
  NAND2_X1 U2729 ( .A1(n2905), .A2(REG1_REG_3__SCAN_IN), .ZN(n2908) );
  NAND2_X1 U2730 ( .A1(n3825), .A2(n3826), .ZN(n2083) );
  NAND2_X1 U2731 ( .A1(n2089), .A2(n2085), .ZN(n4314) );
  AND2_X1 U2732 ( .A1(n2088), .A2(n2090), .ZN(n2085) );
  NOR2_X1 U2733 ( .A1(n4302), .A2(n2092), .ZN(n3304) );
  NAND2_X1 U2734 ( .A1(n4302), .A2(n4444), .ZN(n2089) );
  INV_X1 U2735 ( .A(n2093), .ZN(n4313) );
  NAND3_X1 U2736 ( .A1(n2097), .A2(n2100), .A3(n2095), .ZN(n4323) );
  NAND3_X1 U2737 ( .A1(n2097), .A2(n2096), .A3(n2095), .ZN(n2102) );
  INV_X1 U2738 ( .A(n2102), .ZN(n4322) );
  NAND3_X1 U2739 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .A3(
        IR_REG_1__SCAN_IN), .ZN(n2155) );
  NAND3_X1 U2740 ( .A1(n2736), .A2(n3521), .A3(n3525), .ZN(n2112) );
  NAND3_X1 U2741 ( .A1(n2736), .A2(n3521), .A3(n2040), .ZN(n2114) );
  NAND2_X1 U2742 ( .A1(n2115), .A2(n2117), .ZN(n2818) );
  NAND3_X1 U2743 ( .A1(n2792), .A2(n2120), .A3(n3554), .ZN(n2115) );
  NAND3_X1 U2744 ( .A1(n2792), .A2(n3554), .A3(n2125), .ZN(n2116) );
  NAND3_X1 U2745 ( .A1(n2792), .A2(n3554), .A3(n2128), .ZN(n2122) );
  NAND2_X1 U2746 ( .A1(n3607), .A2(n2128), .ZN(n2126) );
  INV_X1 U2747 ( .A(n3513), .ZN(n2128) );
  NAND3_X1 U2748 ( .A1(n2132), .A2(n3502), .A3(n2129), .ZN(n3588) );
  NAND2_X1 U2749 ( .A1(n3481), .A2(n2143), .ZN(n2142) );
  NOR2_X1 U2750 ( .A1(n2522), .A2(n2152), .ZN(n2576) );
  MUX2_X1 U2751 ( .A(n2887), .B(REG2_REG_1__SCAN_IN), .S(n2886), .Z(n3815) );
  NAND2_X1 U2752 ( .A1(n2934), .A2(n4281), .ZN(n2165) );
  NAND2_X1 U2753 ( .A1(n2166), .A2(n3025), .ZN(n2533) );
  OAI22_X1 U2754 ( .A1(n3759), .A2(n2963), .B1(n4140), .B2(n2166), .ZN(n4368)
         );
  OAI22_X1 U2755 ( .A1(n3610), .A2(n2166), .B1(n3069), .B2(n3612), .ZN(n3033)
         );
  NAND2_X1 U2756 ( .A1(n4007), .A2(n2025), .ZN(n2167) );
  NAND2_X1 U2757 ( .A1(n2167), .A2(n2168), .ZN(n3954) );
  NAND2_X1 U2758 ( .A1(n3139), .A2(n3748), .ZN(n3140) );
  OAI22_X2 U2759 ( .A1(n3084), .A2(n2178), .B1(n2177), .B2(n2300), .ZN(n3139)
         );
  NAND2_X1 U2760 ( .A1(n3140), .A2(n2315), .ZN(n3186) );
  XNOR2_X1 U2761 ( .A(n3906), .B(n3905), .ZN(n3936) );
  OAI21_X2 U2762 ( .B1(n3937), .B2(n2035), .A(n2508), .ZN(n3906) );
  OAI21_X1 U2763 ( .B1(n3334), .B2(n2182), .A(n2180), .ZN(n3354) );
  INV_X1 U2764 ( .A(n3751), .ZN(n2184) );
  INV_X1 U2765 ( .A(n3334), .ZN(n2185) );
  NOR2_X1 U2766 ( .A1(n2573), .A2(n2190), .ZN(n2223) );
  INV_X1 U2767 ( .A(n2573), .ZN(n2188) );
  NAND3_X1 U2768 ( .A1(n2220), .A2(n2192), .A3(n2191), .ZN(n2190) );
  OAI21_X2 U2769 ( .B1(n3182), .B2(n2343), .A(n2344), .ZN(n3240) );
  NAND3_X1 U2770 ( .A1(n2967), .A2(n2535), .A3(n2247), .ZN(n3063) );
  AOI21_X2 U2771 ( .B1(n2195), .B2(n2194), .A(n2193), .ZN(n4069) );
  XNOR2_X2 U2772 ( .A(n2253), .B(IR_REG_2__SCAN_IN), .ZN(n4286) );
  NAND2_X1 U2773 ( .A1(n2615), .A2(n4380), .ZN(n3011) );
  NAND2_X1 U2774 ( .A1(n3029), .A2(n2641), .ZN(n3056) );
  NOR2_X1 U2775 ( .A1(n3597), .A2(n3599), .ZN(n3491) );
  NAND2_X1 U2776 ( .A1(n2245), .A2(n2211), .ZN(n2261) );
  NAND2_X2 U2777 ( .A1(n2866), .A2(n2239), .ZN(n2398) );
  NAND2_X2 U2778 ( .A1(n4030), .A2(n2203), .ZN(n4007) );
  INV_X1 U2779 ( .A(n4049), .ZN(n4050) );
  NOR2_X2 U2780 ( .A1(n3019), .A2(n2635), .ZN(n3030) );
  NOR2_X1 U2781 ( .A1(n3021), .A2(n3020), .ZN(n3019) );
  OAI21_X1 U2782 ( .B1(n4024), .B2(n2398), .A(n2473), .ZN(n4036) );
  OR2_X1 U2783 ( .A1(n2813), .A2(n2974), .ZN(n2197) );
  AND2_X1 U2784 ( .A1(n2648), .A2(n2647), .ZN(n2198) );
  NAND2_X1 U2785 ( .A1(n4037), .A2(n4059), .ZN(n2199) );
  AND2_X1 U2786 ( .A1(n4076), .A2(n4053), .ZN(n2201) );
  OAI22_X1 U2787 ( .A1(n3240), .A2(n2352), .B1(n2541), .B2(n2687), .ZN(n3334)
         );
  OR2_X1 U2788 ( .A1(n2474), .A2(n4014), .ZN(n2202) );
  OR2_X1 U2789 ( .A1(n4015), .A2(n3590), .ZN(n2203) );
  INV_X1 U2790 ( .A(n4424), .ZN(n2619) );
  NOR2_X1 U2791 ( .A1(n2398), .A2(n3570), .ZN(n2204) );
  AND4_X1 U2792 ( .A1(n2217), .A2(n2216), .A3(n2215), .A4(n2214), .ZN(n2218)
         );
  INV_X1 U2793 ( .A(n4036), .ZN(n2474) );
  NAND2_X1 U2794 ( .A1(n3025), .A2(n2628), .ZN(n2629) );
  OR2_X1 U2795 ( .A1(n2623), .A2(n4277), .ZN(n2826) );
  AND2_X1 U2796 ( .A1(n3741), .A2(n3955), .ZN(n3654) );
  NAND2_X1 U2797 ( .A1(n3154), .A2(n3568), .ZN(n3684) );
  NAND2_X1 U2798 ( .A1(n2288), .A2(n3117), .ZN(n3085) );
  INV_X1 U2799 ( .A(IR_REG_4__SCAN_IN), .ZN(n2274) );
  INV_X1 U2800 ( .A(n2787), .ZN(n2788) );
  INV_X1 U2801 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2406) );
  INV_X1 U2802 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2364) );
  INV_X1 U2803 ( .A(IR_REG_18__SCAN_IN), .ZN(n2229) );
  NOR2_X1 U2804 ( .A1(n2601), .A2(n2860), .ZN(n2583) );
  AND2_X1 U2805 ( .A1(n2808), .A2(n2807), .ZN(n2809) );
  NAND2_X1 U2806 ( .A1(n2625), .A2(n2029), .ZN(n2626) );
  NOR2_X1 U2807 ( .A1(n2494), .A2(n4539), .ZN(n2502) );
  NOR2_X1 U2808 ( .A1(n2447), .A2(n2446), .ZN(n2455) );
  INV_X1 U2809 ( .A(n4384), .ZN(n3882) );
  AND2_X1 U2810 ( .A1(n2502), .A2(REG3_REG_27__SCAN_IN), .ZN(n2509) );
  AND2_X1 U2811 ( .A1(n4141), .A2(n4118), .ZN(n2444) );
  NAND2_X1 U2812 ( .A1(n2422), .A2(REG3_REG_17__SCAN_IN), .ZN(n2434) );
  NOR2_X1 U2813 ( .A1(n2407), .A2(n2406), .ZN(n2422) );
  NAND2_X1 U2814 ( .A1(n2389), .A2(REG3_REG_14__SCAN_IN), .ZN(n2396) );
  OR2_X1 U2815 ( .A1(n2353), .A2(n3388), .ZN(n2365) );
  NAND2_X1 U2816 ( .A1(n2292), .A2(REG3_REG_6__SCAN_IN), .ZN(n2303) );
  NAND2_X1 U2817 ( .A1(n3678), .A2(n3681), .ZN(n2535) );
  INV_X1 U2818 ( .A(n3527), .ZN(n2730) );
  AND2_X1 U2819 ( .A1(n2530), .A2(n4276), .ZN(n2878) );
  NAND2_X1 U2820 ( .A1(n2345), .A2(REG3_REG_10__SCAN_IN), .ZN(n2353) );
  OR2_X1 U2821 ( .A1(n3576), .A2(n2759), .ZN(n2760) );
  NOR2_X1 U2822 ( .A1(n2279), .A2(n2267), .ZN(n2292) );
  NAND2_X1 U2823 ( .A1(n3472), .A2(n2790), .ZN(n3553) );
  INV_X1 U2824 ( .A(n3626), .ZN(n3612) );
  OR2_X1 U2825 ( .A1(n3930), .A2(n2398), .ZN(n2517) );
  AND2_X1 U2826 ( .A1(n2461), .A2(REG3_REG_22__SCAN_IN), .ZN(n2468) );
  AOI21_X1 U2827 ( .B1(n3004), .B2(n3003), .A(n3002), .ZN(n3006) );
  INV_X1 U2828 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3388) );
  AND2_X1 U2829 ( .A1(n2881), .A2(n2880), .ZN(n2945) );
  OR2_X1 U2830 ( .A1(n2509), .A2(n2503), .ZN(n3941) );
  INV_X1 U2831 ( .A(n4017), .ZN(n3982) );
  OR2_X1 U2832 ( .A1(n3747), .A2(n2419), .ZN(n3396) );
  OR2_X1 U2833 ( .A1(n2419), .A2(n2418), .ZN(n3397) );
  NAND2_X1 U2834 ( .A1(n2878), .A2(n2982), .ZN(n4133) );
  OR2_X1 U2835 ( .A1(n2872), .A2(D_REG_0__SCAN_IN), .ZN(n2603) );
  INV_X1 U2836 ( .A(n4126), .ZN(n4143) );
  NAND2_X1 U2837 ( .A1(n2532), .A2(n3900), .ZN(n4080) );
  INV_X1 U2838 ( .A(n2584), .ZN(n2602) );
  OR3_X1 U2839 ( .A1(n2338), .A2(IR_REG_8__SCAN_IN), .A3(IR_REG_7__SCAN_IN), 
        .ZN(n2341) );
  NAND2_X1 U2840 ( .A1(n2845), .A2(n2844), .ZN(n2846) );
  AND2_X1 U2841 ( .A1(n2833), .A2(n2832), .ZN(n3623) );
  AOI21_X1 U2842 ( .B1(n3056), .B2(n3055), .A(n2198), .ZN(n3564) );
  NAND2_X1 U2843 ( .A1(n2836), .A2(n4153), .ZN(n3625) );
  AND2_X1 U2844 ( .A1(n2517), .A2(n2516), .ZN(n3918) );
  AND2_X1 U2845 ( .A1(n2945), .A2(n4287), .ZN(n4330) );
  AOI21_X1 U2846 ( .B1(n4049), .B2(n2199), .A(n2201), .ZN(n4032) );
  OR2_X1 U2847 ( .A1(n2413), .A2(n2412), .ZN(n4147) );
  INV_X1 U2848 ( .A(n4107), .ZN(n4362) );
  AND2_X1 U2849 ( .A1(n2603), .A2(n2875), .ZN(n2822) );
  NAND2_X1 U2850 ( .A1(n4080), .A2(n4425), .ZN(n4417) );
  INV_X1 U2851 ( .A(n2822), .ZN(n3043) );
  INV_X1 U2852 ( .A(n3011), .ZN(n3041) );
  INV_X1 U2853 ( .A(n2606), .ZN(n3790) );
  NOR2_X1 U2854 ( .A1(n2850), .A2(n2615), .ZN(n2897) );
  NOR2_X1 U2855 ( .A1(n2847), .A2(n2846), .ZN(n2848) );
  INV_X1 U2856 ( .A(n3632), .ZN(n3617) );
  INV_X1 U2857 ( .A(n3918), .ZN(n3949) );
  INV_X1 U2858 ( .A(n3960), .ZN(n3997) );
  INV_X1 U2859 ( .A(n4141), .ZN(n3802) );
  INV_X1 U2860 ( .A(n4285), .ZN(n2896) );
  INV_X1 U2861 ( .A(n4330), .ZN(n4358) );
  INV_X1 U2862 ( .A(n4353), .ZN(n4321) );
  NAND2_X1 U2863 ( .A1(n4375), .A2(n3142), .ZN(n4137) );
  OR2_X1 U2864 ( .A1(n3135), .A2(n4424), .ZN(n4107) );
  OR2_X1 U2865 ( .A1(n3928), .A2(n4223), .ZN(n2608) );
  NAND2_X1 U2866 ( .A1(n4443), .A2(n2619), .ZN(n4223) );
  INV_X1 U2867 ( .A(n4443), .ZN(n4441) );
  NAND2_X1 U2868 ( .A1(n4431), .A2(n2619), .ZN(n4271) );
  AND3_X1 U2869 ( .A1(n4422), .A2(n4421), .A3(n4420), .ZN(n4440) );
  INV_X1 U2870 ( .A(n4431), .ZN(n4429) );
  NAND2_X1 U2871 ( .A1(n2872), .A2(n3041), .ZN(n4378) );
  AND2_X1 U2872 ( .A1(n2405), .A2(n2414), .ZN(n4278) );
  AND2_X1 U2873 ( .A1(n2323), .A2(n2314), .ZN(n4280) );
  INV_X1 U2874 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2433) );
  INV_X1 U2875 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2205) );
  NAND2_X1 U2876 ( .A1(n2436), .A2(n2205), .ZN(n2206) );
  NAND2_X1 U2877 ( .A1(n2447), .A2(n2206), .ZN(n4108) );
  NAND4_X1 U2878 ( .A1(n2210), .A2(n2209), .A3(n2208), .A4(n2207), .ZN(n2383)
         );
  NAND3_X1 U2879 ( .A1(n2274), .A2(n2273), .A3(n2385), .ZN(n2212) );
  NOR2_X1 U2880 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2217)
         );
  AOI22_X1 U2881 ( .A1(n2006), .A2(REG1_REG_19__SCAN_IN), .B1(n2280), .B2(
        REG0_REG_19__SCAN_IN), .ZN(n2227) );
  INV_X1 U2882 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4109) );
  OR2_X1 U2883 ( .A1(n2355), .A2(n4109), .ZN(n2226) );
  INV_X1 U2884 ( .A(n4130), .ZN(n2445) );
  NAND2_X1 U2885 ( .A1(n2441), .A2(n2229), .ZN(n2522) );
  NAND2_X1 U2886 ( .A1(n2220), .A2(n2869), .ZN(n2230) );
  NAND2_X1 U2887 ( .A1(n2883), .A2(n2191), .ZN(n2233) );
  MUX2_X1 U2888 ( .A(DATAI_19_), .B(n4277), .S(n2326), .Z(n3497) );
  INV_X1 U2889 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2942) );
  NAND2_X1 U2890 ( .A1(n2007), .A2(REG1_REG_0__SCAN_IN), .ZN(n2234) );
  AND2_X1 U2891 ( .A1(n2235), .A2(n2234), .ZN(n2238) );
  INV_X1 U2892 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3018) );
  MUX2_X1 U2893 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(n2326), .Z(n3015) );
  NAND2_X1 U2894 ( .A1(n2007), .A2(REG1_REG_1__SCAN_IN), .ZN(n2244) );
  OR2_X1 U2895 ( .A1(n2240), .A2(n2224), .ZN(n2243) );
  NAND2_X1 U2896 ( .A1(n2280), .A2(REG0_REG_1__SCAN_IN), .ZN(n2242) );
  INV_X1 U2897 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2887) );
  INV_X1 U2898 ( .A(n2245), .ZN(n2246) );
  INV_X1 U2899 ( .A(n2886), .ZN(n3820) );
  MUX2_X1 U2900 ( .A(DATAI_1_), .B(n3820), .S(n2326), .Z(n3025) );
  NAND2_X1 U2901 ( .A1(n3813), .A2(n2974), .ZN(n3675) );
  NAND2_X1 U2902 ( .A1(n3813), .A2(n3025), .ZN(n2247) );
  INV_X1 U2903 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3036) );
  OR2_X1 U2904 ( .A1(n2398), .A2(n3036), .ZN(n2252) );
  NAND2_X1 U2905 ( .A1(n2008), .A2(REG1_REG_2__SCAN_IN), .ZN(n2251) );
  INV_X1 U2906 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2888) );
  OR2_X1 U2907 ( .A1(n2355), .A2(n2888), .ZN(n2250) );
  NAND2_X1 U2908 ( .A1(n2280), .A2(REG0_REG_2__SCAN_IN), .ZN(n2249) );
  MUX2_X1 U2909 ( .A(DATAI_2_), .B(n4286), .S(n2326), .Z(n3073) );
  NAND2_X1 U2910 ( .A1(n3105), .A2(n3073), .ZN(n3678) );
  INV_X1 U2911 ( .A(n3073), .ZN(n2636) );
  NAND2_X1 U2912 ( .A1(n2254), .A2(n2636), .ZN(n3681) );
  NAND2_X1 U2913 ( .A1(n3105), .A2(n2636), .ZN(n2255) );
  NAND2_X1 U2914 ( .A1(n3063), .A2(n2255), .ZN(n3101) );
  NAND2_X1 U2915 ( .A1(n2006), .A2(REG1_REG_3__SCAN_IN), .ZN(n2260) );
  NAND2_X1 U2916 ( .A1(n2280), .A2(REG0_REG_3__SCAN_IN), .ZN(n2259) );
  OR2_X1 U2917 ( .A1(n2398), .A2(REG3_REG_3__SCAN_IN), .ZN(n2258) );
  INV_X1 U2918 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2256) );
  OR2_X1 U2919 ( .A1(n2355), .A2(n2256), .ZN(n2257) );
  NAND2_X1 U2920 ( .A1(n2261), .A2(IR_REG_31__SCAN_IN), .ZN(n2262) );
  NAND2_X1 U2921 ( .A1(n2262), .A2(n2273), .ZN(n2286) );
  OR2_X1 U2922 ( .A1(n2262), .A2(n2273), .ZN(n2263) );
  MUX2_X1 U2923 ( .A(DATAI_3_), .B(n4285), .S(n2326), .Z(n3103) );
  NAND2_X1 U2924 ( .A1(n3567), .A2(n3103), .ZN(n2264) );
  NAND2_X1 U2925 ( .A1(n3101), .A2(n2264), .ZN(n2266) );
  NAND2_X1 U2926 ( .A1(n3069), .A2(n3109), .ZN(n2265) );
  NAND2_X1 U2927 ( .A1(n2266), .A2(n2265), .ZN(n3084) );
  NAND2_X1 U2928 ( .A1(n2280), .A2(REG0_REG_5__SCAN_IN), .ZN(n2272) );
  NAND2_X1 U2929 ( .A1(n2008), .A2(REG1_REG_5__SCAN_IN), .ZN(n2271) );
  AND2_X1 U2930 ( .A1(n2279), .A2(n2267), .ZN(n2268) );
  OR2_X1 U2931 ( .A1(n2268), .A2(n2292), .ZN(n3538) );
  OR2_X1 U2932 ( .A1(n2398), .A2(n3538), .ZN(n2270) );
  INV_X1 U2933 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3157) );
  OR2_X1 U2934 ( .A1(n2355), .A2(n3157), .ZN(n2269) );
  INV_X1 U2935 ( .A(DATAI_5_), .ZN(n2278) );
  NAND2_X1 U2936 ( .A1(n2274), .A2(n2273), .ZN(n2275) );
  NAND2_X1 U2937 ( .A1(n2384), .A2(IR_REG_31__SCAN_IN), .ZN(n2277) );
  INV_X1 U2938 ( .A(IR_REG_5__SCAN_IN), .ZN(n2276) );
  XNOR2_X1 U2939 ( .A(n2277), .B(n2276), .ZN(n4282) );
  MUX2_X1 U2940 ( .A(n2278), .B(n4282), .S(n2326), .Z(n3158) );
  INV_X1 U2941 ( .A(n2291), .ZN(n2288) );
  INV_X1 U2942 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2921) );
  OR2_X1 U2943 ( .A1(n2355), .A2(n2921), .ZN(n2285) );
  OAI21_X1 U2944 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        n2279), .ZN(n3570) );
  NAND2_X1 U2945 ( .A1(n2280), .A2(REG0_REG_4__SCAN_IN), .ZN(n2282) );
  NAND2_X1 U2946 ( .A1(n2006), .A2(REG1_REG_4__SCAN_IN), .ZN(n2281) );
  NAND2_X1 U2947 ( .A1(n2282), .A2(n2281), .ZN(n2283) );
  INV_X1 U2948 ( .A(n3812), .ZN(n3154) );
  NAND2_X1 U2949 ( .A1(n2286), .A2(IR_REG_31__SCAN_IN), .ZN(n2287) );
  XNOR2_X1 U2950 ( .A(n2287), .B(IR_REG_4__SCAN_IN), .ZN(n4284) );
  MUX2_X1 U2951 ( .A(DATAI_4_), .B(n4284), .S(n2326), .Z(n3568) );
  INV_X1 U2952 ( .A(n3568), .ZN(n2652) );
  NAND2_X1 U2953 ( .A1(n3812), .A2(n2652), .ZN(n3687) );
  NAND2_X1 U2954 ( .A1(n3684), .A2(n3687), .ZN(n3117) );
  NAND2_X1 U2955 ( .A1(n3812), .A2(n3568), .ZN(n3149) );
  INV_X1 U2956 ( .A(n3158), .ZN(n3537) );
  NAND2_X1 U2957 ( .A1(n3569), .A2(n3537), .ZN(n2289) );
  AND2_X1 U2958 ( .A1(n3149), .A2(n2289), .ZN(n2290) );
  OR2_X1 U2959 ( .A1(n2291), .A2(n2290), .ZN(n3086) );
  NAND2_X1 U2960 ( .A1(n2280), .A2(REG0_REG_6__SCAN_IN), .ZN(n2298) );
  NAND2_X1 U2961 ( .A1(n2007), .A2(REG1_REG_6__SCAN_IN), .ZN(n2297) );
  OR2_X1 U2962 ( .A1(n2292), .A2(REG3_REG_6__SCAN_IN), .ZN(n2293) );
  NAND2_X1 U2963 ( .A1(n2303), .A2(n2293), .ZN(n3208) );
  OR2_X1 U2964 ( .A1(n2398), .A2(n3208), .ZN(n2296) );
  INV_X1 U2965 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2294) );
  OR2_X1 U2966 ( .A1(n2355), .A2(n2294), .ZN(n2295) );
  NAND4_X1 U2967 ( .A1(n2298), .A2(n2297), .A3(n2296), .A4(n2295), .ZN(n3811)
         );
  OR2_X1 U2968 ( .A1(n2311), .A2(n2869), .ZN(n2299) );
  XNOR2_X1 U2969 ( .A(n2299), .B(IR_REG_6__SCAN_IN), .ZN(n4281) );
  MUX2_X1 U2970 ( .A(DATAI_6_), .B(n4281), .S(n2326), .Z(n3205) );
  AND2_X1 U2971 ( .A1(n3086), .A2(n2028), .ZN(n2300) );
  INV_X1 U2972 ( .A(n3205), .ZN(n2664) );
  NAND2_X1 U2973 ( .A1(n2665), .A2(n2664), .ZN(n2301) );
  NAND2_X1 U2974 ( .A1(n2280), .A2(REG0_REG_7__SCAN_IN), .ZN(n2309) );
  NAND2_X1 U2975 ( .A1(n2008), .A2(REG1_REG_7__SCAN_IN), .ZN(n2308) );
  NAND2_X1 U2976 ( .A1(n2303), .A2(n2302), .ZN(n2304) );
  NAND2_X1 U2977 ( .A1(n2317), .A2(n2304), .ZN(n3228) );
  OR2_X1 U2978 ( .A1(n2398), .A2(n3228), .ZN(n2307) );
  INV_X1 U2979 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2305) );
  OR2_X1 U2980 ( .A1(n2355), .A2(n2305), .ZN(n2306) );
  NAND4_X1 U2981 ( .A1(n2309), .A2(n2308), .A3(n2307), .A4(n2306), .ZN(n3810)
         );
  INV_X1 U2982 ( .A(n3810), .ZN(n2668) );
  NAND2_X1 U2983 ( .A1(n2311), .A2(n2310), .ZN(n2338) );
  NAND2_X1 U2984 ( .A1(n2338), .A2(IR_REG_31__SCAN_IN), .ZN(n2313) );
  INV_X1 U2985 ( .A(IR_REG_7__SCAN_IN), .ZN(n2312) );
  NAND2_X1 U2986 ( .A1(n2313), .A2(n2312), .ZN(n2323) );
  OR2_X1 U2987 ( .A1(n2313), .A2(n2312), .ZN(n2314) );
  MUX2_X1 U2988 ( .A(DATAI_7_), .B(n4280), .S(n2326), .Z(n3225) );
  NAND2_X1 U2989 ( .A1(n2668), .A2(n3225), .ZN(n3694) );
  INV_X1 U2990 ( .A(n3225), .ZN(n3130) );
  NAND2_X1 U2991 ( .A1(n3810), .A2(n3130), .ZN(n3696) );
  NAND2_X1 U2992 ( .A1(n3694), .A2(n3696), .ZN(n3748) );
  NAND2_X1 U2993 ( .A1(n3810), .A2(n3225), .ZN(n2315) );
  NAND2_X1 U2994 ( .A1(n2280), .A2(REG0_REG_8__SCAN_IN), .ZN(n2322) );
  NAND2_X1 U2995 ( .A1(n2006), .A2(REG1_REG_8__SCAN_IN), .ZN(n2321) );
  NAND2_X1 U2996 ( .A1(n2317), .A2(n2316), .ZN(n2318) );
  NAND2_X1 U2997 ( .A1(n2331), .A2(n2318), .ZN(n3277) );
  OR2_X1 U2998 ( .A1(n2398), .A2(n3277), .ZN(n2320) );
  INV_X1 U2999 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3190) );
  OR2_X1 U3000 ( .A1(n2355), .A2(n3190), .ZN(n2319) );
  NAND4_X1 U3001 ( .A1(n2322), .A2(n2321), .A3(n2320), .A4(n2319), .ZN(n3809)
         );
  INV_X1 U3002 ( .A(n3809), .ZN(n3131) );
  INV_X1 U3003 ( .A(DATAI_8_), .ZN(n2327) );
  NAND2_X1 U3004 ( .A1(n2323), .A2(IR_REG_31__SCAN_IN), .ZN(n2325) );
  XNOR2_X1 U3005 ( .A(n2325), .B(n2324), .ZN(n3001) );
  MUX2_X1 U3006 ( .A(n2327), .B(n3001), .S(n2326), .Z(n3193) );
  NAND2_X1 U3007 ( .A1(n3131), .A2(n3193), .ZN(n2328) );
  NAND2_X1 U3008 ( .A1(n3186), .A2(n2328), .ZN(n2330) );
  INV_X1 U3009 ( .A(n3193), .ZN(n3274) );
  NAND2_X1 U3010 ( .A1(n3809), .A2(n3274), .ZN(n2329) );
  NAND2_X1 U3011 ( .A1(n2280), .A2(REG0_REG_9__SCAN_IN), .ZN(n2337) );
  NAND2_X1 U3012 ( .A1(n2008), .A2(REG1_REG_9__SCAN_IN), .ZN(n2336) );
  INV_X1 U3013 ( .A(n2345), .ZN(n2333) );
  NAND2_X1 U3014 ( .A1(n2331), .A2(n4461), .ZN(n2332) );
  NAND2_X1 U3015 ( .A1(n2333), .A2(n2332), .ZN(n3287) );
  OR2_X1 U3016 ( .A1(n2398), .A2(n3287), .ZN(n2335) );
  INV_X1 U3017 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3180) );
  OR2_X1 U3018 ( .A1(n2355), .A2(n3180), .ZN(n2334) );
  NAND4_X1 U3019 ( .A1(n2337), .A2(n2336), .A3(n2335), .A4(n2334), .ZN(n3482)
         );
  NAND2_X1 U3020 ( .A1(n2341), .A2(IR_REG_31__SCAN_IN), .ZN(n2339) );
  MUX2_X1 U3021 ( .A(IR_REG_31__SCAN_IN), .B(n2339), .S(IR_REG_9__SCAN_IN), 
        .Z(n2340) );
  INV_X1 U3022 ( .A(n2340), .ZN(n2342) );
  MUX2_X1 U3023 ( .A(DATAI_9_), .B(n4279), .S(n2326), .Z(n3284) );
  AND2_X1 U3024 ( .A1(n3482), .A2(n3284), .ZN(n2343) );
  NAND2_X1 U3025 ( .A1(n3234), .A2(n3178), .ZN(n2344) );
  NAND2_X1 U3026 ( .A1(n2280), .A2(REG0_REG_10__SCAN_IN), .ZN(n2350) );
  NAND2_X1 U3027 ( .A1(n2007), .A2(REG1_REG_10__SCAN_IN), .ZN(n2349) );
  OR2_X1 U3028 ( .A1(n2345), .A2(REG3_REG_10__SCAN_IN), .ZN(n2346) );
  NAND2_X1 U3029 ( .A1(n2353), .A2(n2346), .ZN(n3485) );
  OR2_X1 U3030 ( .A1(n2398), .A2(n3485), .ZN(n2348) );
  INV_X1 U3031 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3239) );
  OR2_X1 U3032 ( .A1(n2355), .A2(n3239), .ZN(n2347) );
  NAND4_X1 U3033 ( .A1(n2350), .A2(n2349), .A3(n2348), .A4(n2347), .ZN(n3808)
         );
  OR2_X1 U3034 ( .A1(n2361), .A2(n2869), .ZN(n2351) );
  XNOR2_X1 U3035 ( .A(n2351), .B(IR_REG_10__SCAN_IN), .ZN(n3303) );
  MUX2_X1 U3036 ( .A(DATAI_10_), .B(n3303), .S(n2326), .Z(n3483) );
  NOR2_X1 U3037 ( .A1(n3808), .A2(n3483), .ZN(n2352) );
  INV_X1 U3038 ( .A(n3808), .ZN(n2541) );
  INV_X1 U3039 ( .A(n3483), .ZN(n2687) );
  NAND2_X1 U3040 ( .A1(n2280), .A2(REG0_REG_11__SCAN_IN), .ZN(n2359) );
  NAND2_X1 U3041 ( .A1(n2007), .A2(REG1_REG_11__SCAN_IN), .ZN(n2358) );
  NAND2_X1 U3042 ( .A1(n2353), .A2(n3388), .ZN(n2354) );
  NAND2_X1 U3043 ( .A1(n2365), .A2(n2354), .ZN(n3392) );
  OR2_X1 U3044 ( .A1(n2398), .A2(n3392), .ZN(n2357) );
  INV_X1 U3045 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3346) );
  OR2_X1 U3046 ( .A1(n2355), .A2(n3346), .ZN(n2356) );
  NAND4_X1 U3047 ( .A1(n2359), .A2(n2358), .A3(n2357), .A4(n2356), .ZN(n3484)
         );
  INV_X1 U3048 ( .A(IR_REG_10__SCAN_IN), .ZN(n2360) );
  NAND2_X1 U3049 ( .A1(n2361), .A2(n2360), .ZN(n2362) );
  NAND2_X1 U3050 ( .A1(n2362), .A2(IR_REG_31__SCAN_IN), .ZN(n2373) );
  MUX2_X1 U3051 ( .A(DATAI_11_), .B(n4386), .S(n2326), .Z(n3389) );
  NAND2_X1 U3052 ( .A1(n2695), .A2(n3389), .ZN(n3254) );
  INV_X1 U3053 ( .A(n3389), .ZN(n3344) );
  NAND2_X1 U3054 ( .A1(n3484), .A2(n3344), .ZN(n3256) );
  NAND2_X1 U3055 ( .A1(n2695), .A2(n3344), .ZN(n2363) );
  NAND2_X1 U3056 ( .A1(n2280), .A2(REG0_REG_12__SCAN_IN), .ZN(n2371) );
  NAND2_X1 U3057 ( .A1(n2006), .A2(REG1_REG_12__SCAN_IN), .ZN(n2370) );
  INV_X1 U3058 ( .A(n2376), .ZN(n2367) );
  NAND2_X1 U3059 ( .A1(n2365), .A2(n2364), .ZN(n2366) );
  NAND2_X1 U3060 ( .A1(n2367), .A2(n2366), .ZN(n3435) );
  OR2_X1 U3061 ( .A1(n2398), .A2(n3435), .ZN(n2369) );
  INV_X1 U3062 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3264) );
  OR2_X1 U3063 ( .A1(n2355), .A2(n3264), .ZN(n2368) );
  NAND4_X1 U3064 ( .A1(n2371), .A2(n2370), .A3(n2369), .A4(n2368), .ZN(n3807)
         );
  INV_X1 U3065 ( .A(IR_REG_11__SCAN_IN), .ZN(n2372) );
  NAND2_X1 U3066 ( .A1(n2373), .A2(n2372), .ZN(n2374) );
  NAND2_X1 U3067 ( .A1(n2374), .A2(IR_REG_31__SCAN_IN), .ZN(n2375) );
  XNOR2_X1 U3068 ( .A(n2375), .B(IR_REG_12__SCAN_IN), .ZN(n4444) );
  MUX2_X1 U3069 ( .A(DATAI_12_), .B(n4444), .S(n2326), .Z(n3432) );
  INV_X1 U3070 ( .A(n3807), .ZN(n3361) );
  INV_X1 U3071 ( .A(n3432), .ZN(n3259) );
  NAND2_X1 U3072 ( .A1(n2008), .A2(REG1_REG_13__SCAN_IN), .ZN(n2381) );
  NAND2_X1 U3073 ( .A1(n2280), .A2(REG0_REG_13__SCAN_IN), .ZN(n2380) );
  NOR2_X1 U3074 ( .A1(n2376), .A2(REG3_REG_13__SCAN_IN), .ZN(n2377) );
  OR2_X1 U3075 ( .A1(n2389), .A2(n2377), .ZN(n3447) );
  OR2_X1 U3076 ( .A1(n2398), .A2(n3447), .ZN(n2379) );
  INV_X1 U3077 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3850) );
  OR2_X1 U3078 ( .A1(n2355), .A2(n3850), .ZN(n2378) );
  NAND4_X1 U3079 ( .A1(n2381), .A2(n2380), .A3(n2379), .A4(n2378), .ZN(n3806)
         );
  OAI21_X1 U3080 ( .B1(n2384), .B2(n2383), .A(IR_REG_31__SCAN_IN), .ZN(n2386)
         );
  MUX2_X1 U3081 ( .A(n2386), .B(IR_REG_31__SCAN_IN), .S(n2385), .Z(n2387) );
  AND2_X1 U3082 ( .A1(n2382), .A2(n2387), .ZN(n3853) );
  MUX2_X1 U3083 ( .A(DATAI_13_), .B(n3853), .S(n2326), .Z(n3444) );
  NOR2_X1 U3084 ( .A1(n3806), .A2(n3444), .ZN(n2388) );
  INV_X1 U3085 ( .A(n3806), .ZN(n2705) );
  NAND2_X1 U3086 ( .A1(n2280), .A2(REG0_REG_14__SCAN_IN), .ZN(n2394) );
  NAND2_X1 U3087 ( .A1(n2008), .A2(REG1_REG_14__SCAN_IN), .ZN(n2393) );
  OR2_X1 U3088 ( .A1(n2389), .A2(REG3_REG_14__SCAN_IN), .ZN(n2390) );
  NAND2_X1 U3089 ( .A1(n2396), .A2(n2390), .ZN(n3466) );
  OR2_X1 U3090 ( .A1(n2398), .A2(n3466), .ZN(n2392) );
  INV_X1 U3091 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3320) );
  OR2_X1 U3092 ( .A1(n2355), .A2(n3320), .ZN(n2391) );
  NAND4_X1 U3093 ( .A1(n2394), .A2(n2393), .A3(n2392), .A4(n2391), .ZN(n3805)
         );
  NAND2_X1 U3094 ( .A1(n2382), .A2(IR_REG_31__SCAN_IN), .ZN(n2395) );
  XNOR2_X1 U3095 ( .A(n2395), .B(IR_REG_14__SCAN_IN), .ZN(n4329) );
  MUX2_X1 U3096 ( .A(DATAI_14_), .B(n4329), .S(n2326), .Z(n3463) );
  NAND2_X1 U3097 ( .A1(n3381), .A2(n3463), .ZN(n3638) );
  INV_X1 U3098 ( .A(n3463), .ZN(n3318) );
  NAND2_X1 U3099 ( .A1(n3805), .A2(n3318), .ZN(n3640) );
  NAND2_X1 U3100 ( .A1(n2280), .A2(REG0_REG_15__SCAN_IN), .ZN(n2402) );
  NAND2_X1 U3101 ( .A1(n2006), .A2(REG1_REG_15__SCAN_IN), .ZN(n2401) );
  NAND2_X1 U3102 ( .A1(n2396), .A2(n3622), .ZN(n2397) );
  NAND2_X1 U3103 ( .A1(n2407), .A2(n2397), .ZN(n3629) );
  OR2_X1 U3104 ( .A1(n2398), .A2(n3629), .ZN(n2400) );
  INV_X1 U3105 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3376) );
  OR2_X1 U3106 ( .A1(n2355), .A2(n3376), .ZN(n2399) );
  NAND4_X1 U3107 ( .A1(n2402), .A2(n2401), .A3(n2400), .A4(n2399), .ZN(n3804)
         );
  NAND2_X1 U3108 ( .A1(n2014), .A2(IR_REG_31__SCAN_IN), .ZN(n2404) );
  OR2_X1 U3109 ( .A1(n2404), .A2(n2403), .ZN(n2405) );
  NAND2_X1 U3110 ( .A1(n2404), .A2(n2403), .ZN(n2414) );
  MUX2_X1 U3111 ( .A(DATAI_15_), .B(n4278), .S(n2326), .Z(n3624) );
  AND2_X1 U3112 ( .A1(n3804), .A2(n3624), .ZN(n2419) );
  AND2_X1 U3113 ( .A1(n2407), .A2(n2406), .ZN(n2408) );
  OR2_X1 U3114 ( .A1(n2408), .A2(n2422), .ZN(n3530) );
  INV_X1 U3115 ( .A(REG2_REG_16__SCAN_IN), .ZN(n3402) );
  OR2_X1 U3116 ( .A1(n2355), .A2(n3402), .ZN(n2409) );
  OAI21_X1 U3117 ( .B1(n2398), .B2(n3530), .A(n2409), .ZN(n2413) );
  NAND2_X1 U3118 ( .A1(n2280), .A2(REG0_REG_16__SCAN_IN), .ZN(n2411) );
  NAND2_X1 U3119 ( .A1(n2007), .A2(REG1_REG_16__SCAN_IN), .ZN(n2410) );
  NAND2_X1 U3120 ( .A1(n2411), .A2(n2410), .ZN(n2412) );
  INV_X1 U3121 ( .A(n4147), .ZN(n2416) );
  NAND2_X1 U3122 ( .A1(n2414), .A2(IR_REG_31__SCAN_IN), .ZN(n2415) );
  XNOR2_X1 U3123 ( .A(n2415), .B(n4580), .ZN(n4384) );
  MUX2_X1 U3124 ( .A(DATAI_16_), .B(n3882), .S(n2326), .Z(n3527) );
  NAND2_X1 U3125 ( .A1(n2416), .A2(n3527), .ZN(n3716) );
  NAND2_X1 U3126 ( .A1(n4147), .A2(n2730), .ZN(n3713) );
  INV_X1 U3127 ( .A(n3760), .ZN(n3400) );
  NAND2_X1 U3128 ( .A1(n3381), .A2(n3318), .ZN(n3372) );
  INV_X1 U3129 ( .A(n3804), .ZN(n3408) );
  INV_X1 U3130 ( .A(n3624), .ZN(n3375) );
  NAND2_X1 U3131 ( .A1(n3408), .A2(n3375), .ZN(n2417) );
  AND2_X1 U3132 ( .A1(n3372), .A2(n2417), .ZN(n2418) );
  AND2_X1 U3133 ( .A1(n3400), .A2(n3397), .ZN(n2420) );
  OAI21_X1 U3134 ( .B1(n3312), .B2(n3396), .A(n2420), .ZN(n3399) );
  NAND2_X1 U3135 ( .A1(n4147), .A2(n3527), .ZN(n2421) );
  NAND2_X1 U3136 ( .A1(n3399), .A2(n2421), .ZN(n4159) );
  NAND2_X1 U3137 ( .A1(n2280), .A2(REG0_REG_17__SCAN_IN), .ZN(n2427) );
  NAND2_X1 U3138 ( .A1(n2008), .A2(REG1_REG_17__SCAN_IN), .ZN(n2426) );
  OR2_X1 U3139 ( .A1(n2422), .A2(REG3_REG_17__SCAN_IN), .ZN(n2423) );
  NAND2_X1 U3140 ( .A1(n2434), .A2(n2423), .ZN(n4154) );
  OR2_X1 U3141 ( .A1(n4154), .A2(n2398), .ZN(n2425) );
  INV_X1 U3142 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4550) );
  OR2_X1 U3143 ( .A1(n2355), .A2(n4550), .ZN(n2424) );
  INV_X1 U3144 ( .A(DATAI_17_), .ZN(n2430) );
  OR2_X1 U3145 ( .A1(n2428), .A2(n2869), .ZN(n2429) );
  XNOR2_X1 U3146 ( .A(n2429), .B(IR_REG_17__SCAN_IN), .ZN(n3885) );
  MUX2_X1 U3147 ( .A(n2430), .B(n4382), .S(n2326), .Z(n4149) );
  NAND2_X1 U31480 ( .A1(n4134), .A2(n4149), .ZN(n2432) );
  INV_X1 U31490 ( .A(n4149), .ZN(n3547) );
  AND2_X1 U3150 ( .A1(n3803), .A2(n3547), .ZN(n2431) );
  AOI21_X1 U3151 ( .B1(n4159), .B2(n2432), .A(n2431), .ZN(n4115) );
  NAND2_X1 U3152 ( .A1(n2434), .A2(n2433), .ZN(n2435) );
  NAND2_X1 U3153 ( .A1(n2436), .A2(n2435), .ZN(n4120) );
  OR2_X1 U3154 ( .A1(n4120), .A2(n2398), .ZN(n2440) );
  NAND2_X1 U3155 ( .A1(n2280), .A2(REG0_REG_18__SCAN_IN), .ZN(n2439) );
  NAND2_X1 U3156 ( .A1(n2007), .A2(REG1_REG_18__SCAN_IN), .ZN(n2438) );
  INV_X1 U3157 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4121) );
  OR2_X1 U3158 ( .A1(n2355), .A2(n4121), .ZN(n2437) );
  INV_X1 U3159 ( .A(n2441), .ZN(n2442) );
  NAND2_X1 U3160 ( .A1(n2442), .A2(IR_REG_31__SCAN_IN), .ZN(n2443) );
  XNOR2_X1 U3161 ( .A(n2443), .B(IR_REG_18__SCAN_IN), .ZN(n3895) );
  MUX2_X1 U3162 ( .A(DATAI_18_), .B(n3895), .S(n2326), .Z(n4128) );
  NAND2_X1 U3163 ( .A1(n4141), .A2(n4128), .ZN(n4095) );
  INV_X1 U3164 ( .A(n4128), .ZN(n4118) );
  NAND2_X1 U3165 ( .A1(n3802), .A2(n4118), .ZN(n4096) );
  NAND2_X1 U3166 ( .A1(n4095), .A2(n4096), .ZN(n4114) );
  INV_X1 U3167 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4085) );
  INV_X1 U3168 ( .A(REG3_REG_20__SCAN_IN), .ZN(n2446) );
  AND2_X1 U3169 ( .A1(n2447), .A2(n2446), .ZN(n2448) );
  NOR2_X1 U3170 ( .A1(n2455), .A2(n2448), .ZN(n3581) );
  NAND2_X1 U3171 ( .A1(n3581), .A2(n2449), .ZN(n2451) );
  AOI22_X1 U3172 ( .A1(n2006), .A2(REG1_REG_20__SCAN_IN), .B1(n2280), .B2(
        REG0_REG_20__SCAN_IN), .ZN(n2450) );
  INV_X1 U3173 ( .A(DATAI_20_), .ZN(n2452) );
  INV_X1 U3174 ( .A(n4101), .ZN(n4054) );
  INV_X1 U3175 ( .A(n4081), .ZN(n3765) );
  NOR2_X1 U3176 ( .A1(n2455), .A2(REG3_REG_21__SCAN_IN), .ZN(n2456) );
  OR2_X1 U3177 ( .A1(n2461), .A2(n2456), .ZN(n4062) );
  INV_X1 U3178 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4063) );
  NAND2_X1 U3179 ( .A1(n2280), .A2(REG0_REG_21__SCAN_IN), .ZN(n2458) );
  NAND2_X1 U3180 ( .A1(n2007), .A2(REG1_REG_21__SCAN_IN), .ZN(n2457) );
  OAI211_X1 U3181 ( .C1(n4063), .C2(n2355), .A(n2458), .B(n2457), .ZN(n2459)
         );
  INV_X1 U3182 ( .A(n2459), .ZN(n2460) );
  NAND2_X1 U3183 ( .A1(n2467), .A2(DATAI_21_), .ZN(n4053) );
  INV_X1 U3184 ( .A(n4037), .ZN(n4076) );
  NOR2_X1 U3185 ( .A1(n2461), .A2(REG3_REG_22__SCAN_IN), .ZN(n2462) );
  OR2_X1 U3186 ( .A1(n2468), .A2(n2462), .ZN(n4043) );
  INV_X1 U3187 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4044) );
  NAND2_X1 U3188 ( .A1(n2008), .A2(REG1_REG_22__SCAN_IN), .ZN(n2464) );
  NAND2_X1 U3189 ( .A1(n2280), .A2(REG0_REG_22__SCAN_IN), .ZN(n2463) );
  OAI211_X1 U3190 ( .C1(n2355), .C2(n4044), .A(n2464), .B(n2463), .ZN(n2465)
         );
  INV_X1 U3191 ( .A(n2465), .ZN(n2466) );
  OAI21_X1 U3192 ( .B1(n4043), .B2(n2398), .A(n2466), .ZN(n4056) );
  NAND2_X1 U3193 ( .A1(n2467), .A2(DATAI_22_), .ZN(n3590) );
  OR2_X1 U3194 ( .A1(n4056), .A2(n3590), .ZN(n4011) );
  NAND2_X1 U3195 ( .A1(n4056), .A2(n3590), .ZN(n2554) );
  NAND2_X1 U3196 ( .A1(n4011), .A2(n2554), .ZN(n4031) );
  NAND2_X1 U3197 ( .A1(n4032), .A2(n4031), .ZN(n4030) );
  INV_X1 U3198 ( .A(n4056), .ZN(n4015) );
  OR2_X1 U3199 ( .A1(n2468), .A2(REG3_REG_23__SCAN_IN), .ZN(n2469) );
  NAND2_X1 U3200 ( .A1(n2485), .A2(n2469), .ZN(n4024) );
  INV_X1 U3201 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4025) );
  NAND2_X1 U3202 ( .A1(n2006), .A2(REG1_REG_23__SCAN_IN), .ZN(n2471) );
  NAND2_X1 U3203 ( .A1(n2280), .A2(REG0_REG_23__SCAN_IN), .ZN(n2470) );
  OAI211_X1 U3204 ( .C1(n4025), .C2(n2355), .A(n2471), .B(n2470), .ZN(n2472)
         );
  INV_X1 U3205 ( .A(n2472), .ZN(n2473) );
  NAND2_X1 U3206 ( .A1(n2467), .A2(DATAI_23_), .ZN(n4014) );
  XNOR2_X1 U3207 ( .A(n2485), .B(REG3_REG_24__SCAN_IN), .ZN(n4002) );
  NAND2_X1 U3208 ( .A1(n4002), .A2(n2449), .ZN(n2481) );
  INV_X1 U3209 ( .A(REG2_REG_24__SCAN_IN), .ZN(n2478) );
  NAND2_X1 U32100 ( .A1(n2280), .A2(REG0_REG_24__SCAN_IN), .ZN(n2477) );
  NAND2_X1 U32110 ( .A1(n2008), .A2(REG1_REG_24__SCAN_IN), .ZN(n2476) );
  OAI211_X1 U32120 ( .C1(n2478), .C2(n2355), .A(n2477), .B(n2476), .ZN(n2479)
         );
  INV_X1 U32130 ( .A(n2479), .ZN(n2480) );
  NAND2_X1 U32140 ( .A1(n2467), .A2(DATAI_24_), .ZN(n4001) );
  NOR2_X1 U32150 ( .A1(n3982), .A2(n4001), .ZN(n2483) );
  INV_X1 U32160 ( .A(n4001), .ZN(n2482) );
  INV_X1 U32170 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3557) );
  INV_X1 U32180 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3516) );
  OAI21_X1 U32190 ( .B1(n2485), .B2(n3557), .A(n3516), .ZN(n2486) );
  NAND2_X1 U32200 ( .A1(REG3_REG_24__SCAN_IN), .A2(REG3_REG_25__SCAN_IN), .ZN(
        n2484) );
  NAND2_X1 U32210 ( .A1(n3986), .A2(n2449), .ZN(n2492) );
  INV_X1 U32220 ( .A(REG2_REG_25__SCAN_IN), .ZN(n2489) );
  NAND2_X1 U32230 ( .A1(n2006), .A2(REG1_REG_25__SCAN_IN), .ZN(n2488) );
  NAND2_X1 U32240 ( .A1(n2280), .A2(REG0_REG_25__SCAN_IN), .ZN(n2487) );
  OAI211_X1 U32250 ( .C1(n2489), .C2(n2355), .A(n2488), .B(n2487), .ZN(n2490)
         );
  INV_X1 U32260 ( .A(n2490), .ZN(n2491) );
  INV_X1 U32270 ( .A(DATAI_25_), .ZN(n2493) );
  NOR2_X1 U32280 ( .A1(n2326), .A2(n2493), .ZN(n3978) );
  INV_X1 U32290 ( .A(n3978), .ZN(n3984) );
  INV_X1 U32300 ( .A(REG3_REG_26__SCAN_IN), .ZN(n4539) );
  AND2_X1 U32310 ( .A1(n2494), .A2(n4539), .ZN(n2495) );
  OR2_X1 U32320 ( .A1(n2495), .A2(n2502), .ZN(n3609) );
  INV_X1 U32330 ( .A(REG2_REG_26__SCAN_IN), .ZN(n2498) );
  NAND2_X1 U32340 ( .A1(n2280), .A2(REG0_REG_26__SCAN_IN), .ZN(n2497) );
  NAND2_X1 U32350 ( .A1(n2008), .A2(REG1_REG_26__SCAN_IN), .ZN(n2496) );
  OAI211_X1 U32360 ( .C1(n2498), .C2(n2355), .A(n2497), .B(n2496), .ZN(n2499)
         );
  INV_X1 U32370 ( .A(n2499), .ZN(n2500) );
  OAI21_X1 U32380 ( .B1(n3609), .B2(n2398), .A(n2500), .ZN(n3979) );
  INV_X1 U32390 ( .A(n3979), .ZN(n3947) );
  NAND2_X1 U32400 ( .A1(n2467), .A2(DATAI_26_), .ZN(n3965) );
  NOR2_X1 U32410 ( .A1(n3947), .A2(n3965), .ZN(n2501) );
  OAI22_X1 U32420 ( .A1(n3954), .A2(n2501), .B1(n2800), .B2(n3979), .ZN(n3937)
         );
  NOR2_X1 U32430 ( .A1(n2502), .A2(REG3_REG_27__SCAN_IN), .ZN(n2503) );
  INV_X1 U32440 ( .A(REG2_REG_27__SCAN_IN), .ZN(n3940) );
  NAND2_X1 U32450 ( .A1(n2006), .A2(REG1_REG_27__SCAN_IN), .ZN(n2505) );
  NAND2_X1 U32460 ( .A1(n2280), .A2(REG0_REG_27__SCAN_IN), .ZN(n2504) );
  OAI211_X1 U32470 ( .C1(n3940), .C2(n2355), .A(n2505), .B(n2504), .ZN(n2506)
         );
  INV_X1 U32480 ( .A(n2506), .ZN(n2507) );
  NAND2_X1 U32490 ( .A1(n2467), .A2(DATAI_27_), .ZN(n3946) );
  INV_X1 U32500 ( .A(n3946), .ZN(n3939) );
  NAND2_X1 U32510 ( .A1(n3962), .A2(n3939), .ZN(n2508) );
  NAND2_X1 U32520 ( .A1(n2509), .A2(REG3_REG_28__SCAN_IN), .ZN(n3920) );
  INV_X1 U32530 ( .A(n2509), .ZN(n2511) );
  INV_X1 U32540 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2510) );
  NAND2_X1 U32550 ( .A1(n2511), .A2(n2510), .ZN(n2512) );
  NAND2_X1 U32560 ( .A1(n3920), .A2(n2512), .ZN(n3930) );
  INV_X1 U32570 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3929) );
  NAND2_X1 U32580 ( .A1(n2007), .A2(REG1_REG_28__SCAN_IN), .ZN(n2514) );
  NAND2_X1 U32590 ( .A1(n2280), .A2(REG0_REG_28__SCAN_IN), .ZN(n2513) );
  OAI211_X1 U32600 ( .C1(n3929), .C2(n2355), .A(n2514), .B(n2513), .ZN(n2515)
         );
  INV_X1 U32610 ( .A(n2515), .ZN(n2516) );
  INV_X1 U32620 ( .A(DATAI_28_), .ZN(n2518) );
  NOR2_X1 U32630 ( .A1(n2326), .A2(n2518), .ZN(n3907) );
  INV_X1 U32640 ( .A(n3907), .ZN(n2811) );
  NAND2_X1 U32650 ( .A1(n3949), .A2(n2811), .ZN(n3911) );
  NAND2_X1 U32660 ( .A1(n3918), .A2(n3907), .ZN(n3912) );
  NAND2_X1 U32670 ( .A1(n3911), .A2(n3912), .ZN(n3905) );
  NAND2_X1 U32680 ( .A1(n2527), .A2(n2520), .ZN(n2528) );
  XNOR2_X1 U32690 ( .A(n3047), .B(n2623), .ZN(n2532) );
  AND2_X1 U32700 ( .A1(n2606), .A2(n4277), .ZN(n4367) );
  NAND2_X1 U32710 ( .A1(n4367), .A2(n2623), .ZN(n4425) );
  INV_X1 U32720 ( .A(n3814), .ZN(n3023) );
  NAND2_X1 U32730 ( .A1(n3023), .A2(n3015), .ZN(n3674) );
  OR2_X1 U32740 ( .A1(n3755), .A2(n3674), .ZN(n2534) );
  NAND2_X1 U32750 ( .A1(n2534), .A2(n2533), .ZN(n3067) );
  INV_X1 U32760 ( .A(n2535), .ZN(n3749) );
  NAND2_X1 U32770 ( .A1(n3067), .A2(n3749), .ZN(n3066) );
  NAND2_X1 U32780 ( .A1(n3066), .A2(n3678), .ZN(n3102) );
  NAND2_X1 U32790 ( .A1(n3069), .A2(n3103), .ZN(n3683) );
  NAND2_X1 U32800 ( .A1(n3567), .A2(n3109), .ZN(n3680) );
  NAND2_X1 U32810 ( .A1(n3102), .A2(n3757), .ZN(n2536) );
  INV_X1 U32820 ( .A(n3684), .ZN(n2537) );
  AND2_X1 U32830 ( .A1(n3569), .A2(n3158), .ZN(n3148) );
  NAND2_X1 U32840 ( .A1(n3091), .A2(n3537), .ZN(n3691) );
  NAND2_X1 U32850 ( .A1(n3811), .A2(n2664), .ZN(n3689) );
  NAND2_X1 U32860 ( .A1(n3089), .A2(n3689), .ZN(n2538) );
  NAND2_X1 U32870 ( .A1(n2665), .A2(n3205), .ZN(n3693) );
  INV_X1 U32880 ( .A(n3694), .ZN(n2539) );
  NAND2_X1 U32890 ( .A1(n3131), .A2(n3274), .ZN(n3699) );
  NAND2_X1 U32900 ( .A1(n3809), .A2(n3193), .ZN(n3695) );
  NAND2_X1 U32910 ( .A1(n2540), .A2(n3695), .ZN(n3173) );
  AND2_X1 U32920 ( .A1(n3482), .A2(n3178), .ZN(n3172) );
  NAND2_X1 U32930 ( .A1(n3234), .A2(n3284), .ZN(n3700) );
  NAND2_X1 U32940 ( .A1(n3808), .A2(n2687), .ZN(n3705) );
  NAND2_X1 U32950 ( .A1(n2541), .A2(n3483), .ZN(n3702) );
  NAND2_X1 U32960 ( .A1(n3807), .A2(n3259), .ZN(n3355) );
  NAND2_X1 U32970 ( .A1(n3806), .A2(n3366), .ZN(n3351) );
  NAND2_X1 U32980 ( .A1(n3355), .A2(n3351), .ZN(n2543) );
  INV_X1 U32990 ( .A(n3256), .ZN(n2542) );
  NOR2_X1 U33000 ( .A1(n2543), .A2(n2542), .ZN(n3706) );
  NAND2_X1 U33010 ( .A1(n3337), .A2(n3706), .ZN(n2546) );
  NAND2_X1 U33020 ( .A1(n3361), .A2(n3432), .ZN(n3357) );
  NAND2_X1 U33030 ( .A1(n3254), .A2(n3357), .ZN(n2545) );
  INV_X1 U33040 ( .A(n2543), .ZN(n2544) );
  NOR2_X1 U33050 ( .A1(n3806), .A2(n3366), .ZN(n3352) );
  AOI21_X1 U33060 ( .B1(n2545), .B2(n2544), .A(n3352), .ZN(n3708) );
  NAND2_X1 U33070 ( .A1(n3408), .A2(n3624), .ZN(n3641) );
  NAND2_X1 U33080 ( .A1(n3804), .A2(n3375), .ZN(n3639) );
  NAND2_X1 U33090 ( .A1(n3378), .A2(n3639), .ZN(n3405) );
  NAND2_X1 U33100 ( .A1(n4130), .A2(n4105), .ZN(n3766) );
  NAND2_X1 U33110 ( .A1(n3766), .A2(n4096), .ZN(n2547) );
  AND2_X1 U33120 ( .A1(n3803), .A2(n4149), .ZN(n4092) );
  OR2_X1 U33130 ( .A1(n2547), .A2(n4092), .ZN(n3715) );
  INV_X1 U33140 ( .A(n2547), .ZN(n2549) );
  NAND2_X1 U33150 ( .A1(n4134), .A2(n3547), .ZN(n4093) );
  NAND2_X1 U33160 ( .A1(n4095), .A2(n4093), .ZN(n2548) );
  NAND2_X1 U33170 ( .A1(n2549), .A2(n2548), .ZN(n2550) );
  OR2_X1 U33180 ( .A1(n4130), .A2(n4105), .ZN(n3767) );
  NAND2_X1 U33190 ( .A1(n2550), .A2(n3767), .ZN(n4070) );
  NOR2_X1 U33200 ( .A1(n4101), .A2(n3765), .ZN(n2551) );
  INV_X1 U33210 ( .A(n3719), .ZN(n2552) );
  NAND2_X1 U33220 ( .A1(n4101), .A2(n3765), .ZN(n3718) );
  NAND2_X1 U33230 ( .A1(n2553), .A2(n3718), .ZN(n4051) );
  OR2_X1 U33240 ( .A1(n4037), .A2(n4053), .ZN(n4009) );
  AND2_X1 U33250 ( .A1(n4011), .A2(n4009), .ZN(n3722) );
  NAND2_X1 U33260 ( .A1(n4051), .A2(n3722), .ZN(n2557) );
  NAND2_X1 U33270 ( .A1(n4036), .A2(n4014), .ZN(n3764) );
  AND2_X1 U33280 ( .A1(n3764), .A2(n2554), .ZN(n3726) );
  AND2_X1 U33290 ( .A1(n4037), .A2(n4053), .ZN(n4008) );
  NAND2_X1 U33300 ( .A1(n4011), .A2(n4008), .ZN(n2555) );
  NAND2_X1 U33310 ( .A1(n3726), .A2(n2555), .ZN(n3648) );
  INV_X1 U33320 ( .A(n3648), .ZN(n2556) );
  NAND2_X1 U33330 ( .A1(n2557), .A2(n2556), .ZN(n3993) );
  OR2_X1 U33340 ( .A1(n4017), .A2(n4001), .ZN(n3783) );
  OR2_X1 U33350 ( .A1(n4036), .A2(n4014), .ZN(n3992) );
  NAND2_X1 U33360 ( .A1(n3783), .A2(n3992), .ZN(n3724) );
  INV_X1 U33370 ( .A(n3724), .ZN(n2558) );
  NAND2_X1 U33380 ( .A1(n3993), .A2(n2558), .ZN(n3974) );
  OR2_X1 U33390 ( .A1(n3979), .A2(n3965), .ZN(n3741) );
  NAND2_X1 U33400 ( .A1(n3960), .A2(n3978), .ZN(n3955) );
  INV_X1 U33410 ( .A(n3654), .ZN(n3723) );
  NAND2_X1 U33420 ( .A1(n3997), .A2(n3984), .ZN(n3743) );
  NAND2_X1 U33430 ( .A1(n4017), .A2(n4001), .ZN(n3973) );
  AND2_X1 U33440 ( .A1(n3743), .A2(n3973), .ZN(n3650) );
  INV_X1 U33450 ( .A(n3650), .ZN(n3956) );
  NAND2_X1 U33460 ( .A1(n3956), .A2(n3654), .ZN(n2559) );
  AND2_X1 U33470 ( .A1(n3979), .A2(n3965), .ZN(n3664) );
  INV_X1 U33480 ( .A(n3664), .ZN(n3742) );
  NAND2_X1 U33490 ( .A1(n2559), .A2(n3742), .ZN(n3728) );
  INV_X1 U33500 ( .A(n3728), .ZN(n2560) );
  OAI21_X1 U33510 ( .B1(n3974), .B2(n3723), .A(n2560), .ZN(n3944) );
  XNOR2_X1 U33520 ( .A(n3962), .B(n3946), .ZN(n3945) );
  NOR2_X1 U3353 ( .A1(n3944), .A2(n3945), .ZN(n3943) );
  OR2_X1 U33540 ( .A1(n3962), .A2(n3946), .ZN(n3653) );
  INV_X1 U3355 ( .A(n3653), .ZN(n3659) );
  NOR2_X1 U3356 ( .A1(n3943), .A2(n3659), .ZN(n3914) );
  XNOR2_X1 U3357 ( .A(n3914), .B(n3905), .ZN(n2571) );
  NAND2_X1 U3358 ( .A1(n2530), .A2(n3790), .ZN(n3670) );
  INV_X1 U3359 ( .A(n2623), .ZN(n4276) );
  NAND2_X1 U3360 ( .A1(n4276), .A2(n4277), .ZN(n2561) );
  INV_X1 U3361 ( .A(n3962), .ZN(n3673) );
  NAND2_X1 U3362 ( .A1(n2562), .A2(IR_REG_31__SCAN_IN), .ZN(n2563) );
  XNOR2_X1 U3363 ( .A(n2563), .B(n2191), .ZN(n4287) );
  INV_X1 U3364 ( .A(n4287), .ZN(n2982) );
  OR2_X1 U3365 ( .A1(n3920), .A2(n2398), .ZN(n2568) );
  INV_X1 U3366 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3923) );
  NAND2_X1 U3367 ( .A1(n2280), .A2(REG0_REG_29__SCAN_IN), .ZN(n2565) );
  NAND2_X1 U3368 ( .A1(n2008), .A2(REG1_REG_29__SCAN_IN), .ZN(n2564) );
  OAI211_X1 U3369 ( .C1(n3923), .C2(n2355), .A(n2565), .B(n2564), .ZN(n2566)
         );
  INV_X1 U3370 ( .A(n2566), .ZN(n2567) );
  NAND2_X1 U3371 ( .A1(n2568), .A2(n2567), .ZN(n3740) );
  NAND2_X1 U3372 ( .A1(n2878), .A2(n4287), .ZN(n4140) );
  AOI22_X1 U3373 ( .A1(n3740), .A2(n4129), .B1(n3907), .B2(n4170), .ZN(n2569)
         );
  OAI21_X1 U3374 ( .B1(n3673), .B2(n4133), .A(n2569), .ZN(n2570) );
  AOI21_X1 U3375 ( .B1(n2571), .B2(n4126), .A(n2570), .ZN(n3931) );
  OAI21_X1 U3376 ( .B1(n3936), .B2(n4411), .A(n3931), .ZN(n2611) );
  NOR2_X1 U3377 ( .A1(n2010), .A2(n2869), .ZN(n2572) );
  MUX2_X1 U3378 ( .A(n2869), .B(n2572), .S(IR_REG_25__SCAN_IN), .Z(n2574) );
  NAND2_X1 U3379 ( .A1(n2860), .A2(B_REG_SCAN_IN), .ZN(n2579) );
  NAND2_X1 U3380 ( .A1(n2585), .A2(n2586), .ZN(n2577) );
  MUX2_X1 U3381 ( .A(n2579), .B(B_REG_SCAN_IN), .S(n2584), .Z(n2582) );
  NAND2_X1 U3382 ( .A1(n2573), .A2(IR_REG_31__SCAN_IN), .ZN(n2580) );
  MUX2_X1 U3383 ( .A(IR_REG_31__SCAN_IN), .B(n2580), .S(IR_REG_26__SCAN_IN), 
        .Z(n2581) );
  NAND2_X1 U3384 ( .A1(n2601), .A2(n2860), .ZN(n2873) );
  OAI21_X1 U3385 ( .B1(n2872), .B2(D_REG_1__SCAN_IN), .A(n2873), .ZN(n2600) );
  NAND2_X1 U3386 ( .A1(n2606), .A2(n3900), .ZN(n2587) );
  NAND2_X1 U3387 ( .A1(n2878), .A2(n2587), .ZN(n3040) );
  NAND2_X1 U3388 ( .A1(n3040), .A2(n2835), .ZN(n2588) );
  NOR2_X1 U3389 ( .A1(n3011), .A2(n2588), .ZN(n2599) );
  NOR4_X1 U3390 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_19__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2592) );
  NOR4_X1 U3391 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_17__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2591) );
  NOR4_X1 U3392 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_28__SCAN_IN), .ZN(n2590) );
  NOR4_X1 U3393 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_23__SCAN_IN), .ZN(n2589) );
  NAND4_X1 U3394 ( .A1(n2592), .A2(n2591), .A3(n2590), .A4(n2589), .ZN(n2597)
         );
  NOR2_X1 U3395 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_15__SCAN_IN), .ZN(n4575)
         );
  NOR4_X1 U3396 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_31__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2595) );
  NOR4_X1 U3397 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_10__SCAN_IN), .ZN(n2594) );
  NOR4_X1 U3398 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_6__SCAN_IN), .ZN(n2593) );
  NAND4_X1 U3399 ( .A1(n4575), .A2(n2595), .A3(n2594), .A4(n2593), .ZN(n2596)
         );
  NOR2_X1 U3400 ( .A1(n2597), .A2(n2596), .ZN(n2819) );
  OR2_X1 U3401 ( .A1(n2872), .A2(n2819), .ZN(n2598) );
  NAND2_X1 U3402 ( .A1(n2602), .A2(n2601), .ZN(n2875) );
  INV_X1 U3403 ( .A(n2604), .ZN(n2609) );
  NAND2_X1 U3404 ( .A1(n2974), .A2(n2616), .ZN(n3074) );
  INV_X1 U3405 ( .A(n3922), .ZN(n2605) );
  OAI21_X1 U3406 ( .B1(n3938), .B2(n2811), .A(n2605), .ZN(n3928) );
  NAND2_X1 U3407 ( .A1(n2609), .A2(n2608), .ZN(U3546) );
  INV_X1 U3408 ( .A(n2612), .ZN(n2614) );
  NAND2_X1 U3409 ( .A1(n2614), .A2(n2613), .ZN(U3514) );
  INV_X2 U3410 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3411 ( .A(n3015), .ZN(n2616) );
  INV_X1 U3412 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2618) );
  NAND2_X1 U3413 ( .A1(n2625), .A2(n2196), .ZN(n2979) );
  NAND2_X1 U3414 ( .A1(n2799), .A2(n3814), .ZN(n2622) );
  INV_X1 U3415 ( .A(n2615), .ZN(n2620) );
  AOI22_X1 U3416 ( .A1(n2829), .A2(n3015), .B1(n2620), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2621) );
  NAND2_X1 U3417 ( .A1(n2622), .A2(n2621), .ZN(n2978) );
  NAND2_X1 U3418 ( .A1(n2979), .A2(n2978), .ZN(n2977) );
  AND2_X1 U3419 ( .A1(n2977), .A2(n2626), .ZN(n3021) );
  NAND2_X1 U3420 ( .A1(n2627), .A2(n2829), .ZN(n2630) );
  NAND2_X1 U3421 ( .A1(n2630), .A2(n2629), .ZN(n2631) );
  NAND2_X1 U3422 ( .A1(n3813), .A2(n2799), .ZN(n2632) );
  NAND2_X1 U3423 ( .A1(n2632), .A2(n2197), .ZN(n2634) );
  OAI22_X1 U3424 ( .A1(n2810), .A2(n3105), .B1(n2805), .B2(n2636), .ZN(n2640)
         );
  OAI22_X1 U3425 ( .A1(n3105), .A2(n2813), .B1(n2812), .B2(n2636), .ZN(n2637)
         );
  XNOR2_X1 U3426 ( .A(n2637), .B(n2743), .ZN(n2639) );
  XNOR2_X1 U3427 ( .A(n2638), .B(n2639), .ZN(n3031) );
  NAND2_X1 U3428 ( .A1(n3030), .A2(n3031), .ZN(n3029) );
  OR2_X1 U3429 ( .A1(n2640), .A2(n2639), .ZN(n2641) );
  OAI22_X1 U3430 ( .A1(n3069), .A2(n2810), .B1(n2805), .B2(n3109), .ZN(n2646)
         );
  NAND2_X1 U3431 ( .A1(n3567), .A2(n2829), .ZN(n2643) );
  NAND2_X1 U3432 ( .A1(n2628), .A2(n3103), .ZN(n2642) );
  NAND2_X1 U3433 ( .A1(n2643), .A2(n2642), .ZN(n2644) );
  XNOR2_X1 U3434 ( .A(n2644), .B(n2743), .ZN(n2645) );
  XOR2_X1 U3435 ( .A(n2646), .B(n2645), .Z(n3055) );
  INV_X1 U3436 ( .A(n2645), .ZN(n2648) );
  INV_X1 U3437 ( .A(n2646), .ZN(n2647) );
  NAND2_X1 U3438 ( .A1(n3812), .A2(n2829), .ZN(n2650) );
  NAND2_X1 U3439 ( .A1(n2628), .A2(n3568), .ZN(n2649) );
  NAND2_X1 U3440 ( .A1(n2650), .A2(n2649), .ZN(n2651) );
  XNOR2_X1 U3441 ( .A(n2651), .B(n2743), .ZN(n2654) );
  NOR2_X1 U3442 ( .A1(n2805), .A2(n2652), .ZN(n2653) );
  AOI21_X1 U3443 ( .B1(n2799), .B2(n3812), .A(n2653), .ZN(n2655) );
  XNOR2_X1 U3444 ( .A(n2654), .B(n2655), .ZN(n3563) );
  NAND2_X1 U3445 ( .A1(n3564), .A2(n3563), .ZN(n3562) );
  INV_X1 U3446 ( .A(n2655), .ZN(n2656) );
  NAND2_X1 U3447 ( .A1(n2654), .A2(n2656), .ZN(n2657) );
  NAND2_X1 U3448 ( .A1(n3562), .A2(n2657), .ZN(n3536) );
  OAI22_X1 U3449 ( .A1(n3091), .A2(n2813), .B1(n2812), .B2(n3158), .ZN(n2658)
         );
  XNOR2_X1 U3450 ( .A(n2658), .B(n2743), .ZN(n2660) );
  NOR2_X1 U3451 ( .A1(n2805), .A2(n3158), .ZN(n2659) );
  AOI21_X1 U3452 ( .B1(n2799), .B2(n3569), .A(n2659), .ZN(n2661) );
  XNOR2_X1 U3453 ( .A(n2660), .B(n2661), .ZN(n3535) );
  NAND2_X1 U3454 ( .A1(n3536), .A2(n3535), .ZN(n3534) );
  INV_X1 U3455 ( .A(n2661), .ZN(n2662) );
  NAND2_X1 U3456 ( .A1(n2660), .A2(n2662), .ZN(n2663) );
  OAI22_X1 U3457 ( .A1(n2665), .A2(n2805), .B1(n2812), .B2(n2664), .ZN(n2666)
         );
  XNOR2_X1 U34580 ( .A(n2666), .B(n2743), .ZN(n3202) );
  NOR2_X1 U34590 ( .A1(n2805), .A2(n3130), .ZN(n2667) );
  AOI21_X1 U3460 ( .B1(n2799), .B2(n3810), .A(n2667), .ZN(n2671) );
  OAI22_X1 U3461 ( .A1(n2668), .A2(n2805), .B1(n2812), .B2(n3130), .ZN(n2669)
         );
  XNOR2_X1 U3462 ( .A(n2669), .B(n2743), .ZN(n2670) );
  XOR2_X1 U3463 ( .A(n2671), .B(n2670), .Z(n3223) );
  NAND2_X1 U3464 ( .A1(n3809), .A2(n2829), .ZN(n2673) );
  NAND2_X1 U3465 ( .A1(n3274), .A2(n2628), .ZN(n2672) );
  NAND2_X1 U3466 ( .A1(n2673), .A2(n2672), .ZN(n2674) );
  XNOR2_X1 U34670 ( .A(n2674), .B(n2029), .ZN(n2677) );
  NOR2_X1 U3468 ( .A1(n2805), .A2(n3193), .ZN(n2675) );
  AOI21_X1 U34690 ( .B1(n2799), .B2(n3809), .A(n2675), .ZN(n2676) );
  NAND2_X1 U3470 ( .A1(n2677), .A2(n2676), .ZN(n3271) );
  OAI22_X1 U34710 ( .A1(n3234), .A2(n2810), .B1(n2805), .B2(n3178), .ZN(n2681)
         );
  NAND2_X1 U3472 ( .A1(n3482), .A2(n2829), .ZN(n2679) );
  NAND2_X1 U34730 ( .A1(n2628), .A2(n3284), .ZN(n2678) );
  NAND2_X1 U3474 ( .A1(n2679), .A2(n2678), .ZN(n2680) );
  XNOR2_X1 U34750 ( .A(n2680), .B(n2743), .ZN(n2682) );
  XOR2_X1 U3476 ( .A(n2681), .B(n2682), .Z(n3282) );
  NOR2_X1 U34770 ( .A1(n2682), .A2(n2681), .ZN(n2683) );
  NAND2_X1 U3478 ( .A1(n3808), .A2(n2829), .ZN(n2685) );
  NAND2_X1 U34790 ( .A1(n2628), .A2(n3483), .ZN(n2684) );
  NAND2_X1 U3480 ( .A1(n2685), .A2(n2684), .ZN(n2686) );
  XNOR2_X1 U34810 ( .A(n2686), .B(n2743), .ZN(n2691) );
  NOR2_X1 U3482 ( .A1(n2805), .A2(n2687), .ZN(n2688) );
  AOI21_X1 U34830 ( .B1(n2799), .B2(n3808), .A(n2688), .ZN(n2689) );
  XNOR2_X1 U3484 ( .A(n2691), .B(n2689), .ZN(n3480) );
  INV_X1 U34850 ( .A(n2689), .ZN(n2690) );
  NAND2_X1 U3486 ( .A1(n2691), .A2(n2690), .ZN(n2692) );
  NAND2_X1 U34870 ( .A1(n2799), .A2(n3484), .ZN(n2694) );
  NAND2_X1 U3488 ( .A1(n2829), .A2(n3389), .ZN(n2693) );
  NAND2_X1 U34890 ( .A1(n2694), .A2(n2693), .ZN(n3385) );
  INV_X1 U3490 ( .A(n3385), .ZN(n2697) );
  OAI22_X1 U34910 ( .A1(n2695), .A2(n2805), .B1(n2812), .B2(n3344), .ZN(n2696)
         );
  XNOR2_X1 U3492 ( .A(n2696), .B(n2743), .ZN(n3386) );
  NAND2_X1 U34930 ( .A1(n3807), .A2(n2829), .ZN(n2699) );
  NAND2_X1 U3494 ( .A1(n2628), .A2(n3432), .ZN(n2698) );
  NAND2_X1 U34950 ( .A1(n2699), .A2(n2698), .ZN(n2700) );
  XNOR2_X1 U3496 ( .A(n2700), .B(n2029), .ZN(n2703) );
  NOR2_X1 U34970 ( .A1(n2805), .A2(n3259), .ZN(n2701) );
  AOI21_X1 U3498 ( .B1(n2799), .B2(n3807), .A(n2701), .ZN(n2702) );
  NOR2_X1 U34990 ( .A1(n2703), .A2(n2702), .ZN(n3427) );
  NAND2_X1 U3500 ( .A1(n2703), .A2(n2702), .ZN(n3428) );
  OAI22_X1 U35010 ( .A1(n2705), .A2(n2813), .B1(n2812), .B2(n3366), .ZN(n2704)
         );
  XOR2_X1 U3502 ( .A(n2743), .B(n2704), .Z(n3441) );
  NAND2_X1 U35030 ( .A1(n3439), .A2(n3441), .ZN(n2708) );
  OAI22_X1 U3504 ( .A1(n2705), .A2(n2810), .B1(n2805), .B2(n3366), .ZN(n3440)
         );
  INV_X1 U35050 ( .A(n3439), .ZN(n2707) );
  INV_X1 U35060 ( .A(n3441), .ZN(n2706) );
  AOI22_X2 U35070 ( .A1(n2708), .A2(n3440), .B1(n2707), .B2(n2706), .ZN(n3459)
         );
  NAND2_X1 U35080 ( .A1(n3805), .A2(n2829), .ZN(n2710) );
  NAND2_X1 U35090 ( .A1(n2628), .A2(n3463), .ZN(n2709) );
  NAND2_X1 U35100 ( .A1(n2710), .A2(n2709), .ZN(n2711) );
  XNOR2_X1 U35110 ( .A(n2711), .B(n2743), .ZN(n2717) );
  NAND2_X1 U35120 ( .A1(n2799), .A2(n3805), .ZN(n2713) );
  NAND2_X1 U35130 ( .A1(n2829), .A2(n3463), .ZN(n2712) );
  NAND2_X1 U35140 ( .A1(n2713), .A2(n2712), .ZN(n2718) );
  NAND2_X1 U35150 ( .A1(n2717), .A2(n2718), .ZN(n3457) );
  OAI22_X1 U35160 ( .A1(n3408), .A2(n2805), .B1(n2812), .B2(n3375), .ZN(n2714)
         );
  XOR2_X1 U35170 ( .A(n2743), .B(n2714), .Z(n2716) );
  AND2_X1 U35180 ( .A1(n3457), .A2(n2716), .ZN(n2715) );
  NAND2_X1 U35190 ( .A1(n3459), .A2(n2715), .ZN(n3523) );
  INV_X1 U35200 ( .A(n2716), .ZN(n2724) );
  INV_X1 U35210 ( .A(n2717), .ZN(n2720) );
  INV_X1 U35220 ( .A(n2718), .ZN(n2719) );
  NAND2_X1 U35230 ( .A1(n2720), .A2(n2719), .ZN(n3458) );
  OR2_X1 U35240 ( .A1(n2724), .A2(n3458), .ZN(n3522) );
  NAND2_X1 U35250 ( .A1(n2799), .A2(n3804), .ZN(n2722) );
  NAND2_X1 U35260 ( .A1(n2829), .A2(n3624), .ZN(n2721) );
  NAND2_X1 U35270 ( .A1(n2722), .A2(n2721), .ZN(n3620) );
  AND2_X1 U35280 ( .A1(n3522), .A2(n3620), .ZN(n2723) );
  NAND2_X1 U35290 ( .A1(n3523), .A2(n2723), .ZN(n2736) );
  NAND2_X1 U35300 ( .A1(n3459), .A2(n3457), .ZN(n2726) );
  AND2_X1 U35310 ( .A1(n3458), .A2(n2724), .ZN(n2725) );
  NAND2_X1 U35320 ( .A1(n2726), .A2(n2725), .ZN(n3521) );
  NAND2_X1 U35330 ( .A1(n4147), .A2(n2829), .ZN(n2728) );
  NAND2_X1 U35340 ( .A1(n2628), .A2(n3527), .ZN(n2727) );
  NAND2_X1 U35350 ( .A1(n2728), .A2(n2727), .ZN(n2729) );
  XNOR2_X1 U35360 ( .A(n2729), .B(n2029), .ZN(n2733) );
  INV_X1 U35370 ( .A(n2733), .ZN(n2735) );
  NOR2_X1 U35380 ( .A1(n2805), .A2(n2730), .ZN(n2731) );
  AOI21_X1 U35390 ( .B1(n2799), .B2(n4147), .A(n2731), .ZN(n2732) );
  INV_X1 U35400 ( .A(n2732), .ZN(n2734) );
  AOI21_X1 U35410 ( .B1(n2735), .B2(n2734), .A(n2737), .ZN(n3525) );
  INV_X1 U35420 ( .A(n2737), .ZN(n2738) );
  OAI22_X1 U35430 ( .A1(n4134), .A2(n2805), .B1(n2812), .B2(n4149), .ZN(n2739)
         );
  XNOR2_X1 U35440 ( .A(n2739), .B(n2743), .ZN(n2741) );
  OAI22_X1 U35450 ( .A1(n4134), .A2(n2810), .B1(n2805), .B2(n4149), .ZN(n2740)
         );
  NAND2_X1 U35460 ( .A1(n2741), .A2(n2740), .ZN(n3543) );
  OR2_X1 U35470 ( .A1(n2741), .A2(n2740), .ZN(n3544) );
  AOI22_X1 U35480 ( .A1(n3802), .A2(n2799), .B1(n2829), .B2(n4128), .ZN(n3599)
         );
  OAI22_X1 U35490 ( .A1(n4141), .A2(n2805), .B1(n2812), .B2(n4118), .ZN(n2742)
         );
  XOR2_X1 U35500 ( .A(n2743), .B(n2742), .Z(n3598) );
  NAND2_X1 U35510 ( .A1(n4101), .A2(n2829), .ZN(n2745) );
  NAND2_X1 U35520 ( .A1(n2628), .A2(n4081), .ZN(n2744) );
  NAND2_X1 U35530 ( .A1(n2745), .A2(n2744), .ZN(n2746) );
  XNOR2_X1 U35540 ( .A(n2746), .B(n2743), .ZN(n2755) );
  NAND2_X1 U35550 ( .A1(n4101), .A2(n2799), .ZN(n2748) );
  NAND2_X1 U35560 ( .A1(n2829), .A2(n4081), .ZN(n2747) );
  NAND2_X1 U35570 ( .A1(n2748), .A2(n2747), .ZN(n2756) );
  NAND2_X1 U35580 ( .A1(n2755), .A2(n2756), .ZN(n3575) );
  OR2_X1 U35590 ( .A1(n3492), .A2(n3576), .ZN(n2761) );
  NAND2_X1 U35600 ( .A1(n4130), .A2(n2829), .ZN(n2750) );
  NAND2_X1 U35610 ( .A1(n2628), .A2(n3497), .ZN(n2749) );
  NAND2_X1 U35620 ( .A1(n2750), .A2(n2749), .ZN(n2751) );
  XNOR2_X1 U35630 ( .A(n2751), .B(n2029), .ZN(n2754) );
  NOR2_X1 U35640 ( .A1(n2805), .A2(n4105), .ZN(n2752) );
  AOI21_X1 U35650 ( .B1(n4130), .B2(n2799), .A(n2752), .ZN(n2753) );
  NAND2_X1 U35660 ( .A1(n2754), .A2(n2753), .ZN(n3503) );
  OAI21_X1 U35670 ( .B1(n2754), .B2(n2753), .A(n3503), .ZN(n3493) );
  INV_X1 U35680 ( .A(n2755), .ZN(n2758) );
  INV_X1 U35690 ( .A(n2756), .ZN(n2757) );
  NAND2_X1 U35700 ( .A1(n2758), .A2(n2757), .ZN(n3505) );
  AND2_X1 U35710 ( .A1(n3503), .A2(n3505), .ZN(n2759) );
  NAND2_X1 U35720 ( .A1(n4037), .A2(n2829), .ZN(n2763) );
  NAND2_X1 U35730 ( .A1(n2628), .A2(n4059), .ZN(n2762) );
  NAND2_X1 U35740 ( .A1(n2763), .A2(n2762), .ZN(n2764) );
  XNOR2_X1 U35750 ( .A(n2764), .B(n2743), .ZN(n2768) );
  NAND2_X1 U35760 ( .A1(n4037), .A2(n2799), .ZN(n2766) );
  NAND2_X1 U35770 ( .A1(n2829), .A2(n4059), .ZN(n2765) );
  NAND2_X1 U35780 ( .A1(n2766), .A2(n2765), .ZN(n2767) );
  NAND2_X1 U35790 ( .A1(n2768), .A2(n2767), .ZN(n3502) );
  NAND2_X1 U35800 ( .A1(n4056), .A2(n2829), .ZN(n2770) );
  NAND2_X1 U35810 ( .A1(n2628), .A2(n4042), .ZN(n2769) );
  NAND2_X1 U3582 ( .A1(n2770), .A2(n2769), .ZN(n2771) );
  XNOR2_X1 U3583 ( .A(n2771), .B(n2743), .ZN(n2776) );
  OAI22_X1 U3584 ( .A1(n4015), .A2(n2810), .B1(n2805), .B2(n3590), .ZN(n2777)
         );
  XNOR2_X1 U3585 ( .A(n2776), .B(n2777), .ZN(n3589) );
  NAND2_X1 U3586 ( .A1(n4036), .A2(n2829), .ZN(n2773) );
  NAND2_X1 U3587 ( .A1(n2628), .A2(n4021), .ZN(n2772) );
  NAND2_X1 U3588 ( .A1(n2773), .A2(n2772), .ZN(n2774) );
  XNOR2_X1 U3589 ( .A(n2774), .B(n2743), .ZN(n2783) );
  NOR2_X1 U3590 ( .A1(n2805), .A2(n4014), .ZN(n2775) );
  AOI21_X1 U3591 ( .B1(n4036), .B2(n2799), .A(n2775), .ZN(n2781) );
  XNOR2_X1 U3592 ( .A(n2783), .B(n2781), .ZN(n3473) );
  INV_X1 U3593 ( .A(n2776), .ZN(n2779) );
  INV_X1 U3594 ( .A(n2777), .ZN(n2778) );
  NAND2_X1 U3595 ( .A1(n2779), .A2(n2778), .ZN(n3471) );
  INV_X1 U3596 ( .A(n2781), .ZN(n2782) );
  NAND2_X1 U3597 ( .A1(n2783), .A2(n2782), .ZN(n2786) );
  NAND2_X1 U3598 ( .A1(n3472), .A2(n2786), .ZN(n2785) );
  NOR2_X1 U3599 ( .A1(n2805), .A2(n4001), .ZN(n2784) );
  AOI21_X1 U3600 ( .B1(n4017), .B2(n2799), .A(n2784), .ZN(n2787) );
  NAND2_X2 U3601 ( .A1(n2785), .A2(n2788), .ZN(n3554) );
  INV_X1 U3602 ( .A(n2786), .ZN(n2789) );
  OAI22_X1 U3603 ( .A1(n3982), .A2(n2813), .B1(n2812), .B2(n4001), .ZN(n2791)
         );
  XNOR2_X1 U3604 ( .A(n2791), .B(n2743), .ZN(n3556) );
  NAND2_X1 U3605 ( .A1(n3553), .A2(n3556), .ZN(n2792) );
  OAI22_X1 U3606 ( .A1(n3960), .A2(n2805), .B1(n2812), .B2(n3984), .ZN(n2793)
         );
  XNOR2_X1 U3607 ( .A(n2793), .B(n2743), .ZN(n2795) );
  OAI22_X1 U3608 ( .A1(n3960), .A2(n2810), .B1(n2805), .B2(n3984), .ZN(n2794)
         );
  AND2_X1 U3609 ( .A1(n2795), .A2(n2794), .ZN(n3513) );
  NAND2_X1 U3610 ( .A1(n3979), .A2(n2829), .ZN(n2797) );
  NAND2_X1 U3611 ( .A1(n2628), .A2(n2800), .ZN(n2796) );
  NAND2_X1 U3612 ( .A1(n2797), .A2(n2796), .ZN(n2798) );
  XNOR2_X1 U3613 ( .A(n2798), .B(n2743), .ZN(n2804) );
  NAND2_X1 U3614 ( .A1(n3979), .A2(n2799), .ZN(n2802) );
  NAND2_X1 U3615 ( .A1(n2829), .A2(n2800), .ZN(n2801) );
  NAND2_X1 U3616 ( .A1(n2802), .A2(n2801), .ZN(n2803) );
  NAND2_X1 U3617 ( .A1(n2804), .A2(n2803), .ZN(n3607) );
  OAI22_X1 U3618 ( .A1(n3673), .A2(n2810), .B1(n3946), .B2(n2805), .ZN(n2807)
         );
  OAI22_X1 U3619 ( .A1(n3673), .A2(n2813), .B1(n3946), .B2(n2812), .ZN(n2806)
         );
  XNOR2_X1 U3620 ( .A(n2806), .B(n2743), .ZN(n2808) );
  XOR2_X1 U3621 ( .A(n2807), .B(n2808), .Z(n3451) );
  OAI22_X1 U3622 ( .A1(n3918), .A2(n2810), .B1(n2805), .B2(n2811), .ZN(n2816)
         );
  OAI22_X1 U3623 ( .A1(n3918), .A2(n2813), .B1(n2812), .B2(n2811), .ZN(n2814)
         );
  XNOR2_X1 U3624 ( .A(n2814), .B(n2743), .ZN(n2815) );
  XOR2_X1 U3625 ( .A(n2816), .B(n2815), .Z(n2817) );
  XNOR2_X1 U3626 ( .A(n2818), .B(n2817), .ZN(n2825) );
  AND2_X1 U3627 ( .A1(n2819), .A2(D_REG_1__SCAN_IN), .ZN(n2820) );
  OR2_X1 U3628 ( .A1(n2872), .A2(n2820), .ZN(n2821) );
  AOI21_X1 U3629 ( .B1(n4277), .B2(n2607), .A(n2878), .ZN(n2823) );
  NAND2_X1 U3630 ( .A1(n4139), .A2(n2823), .ZN(n2837) );
  NOR2_X1 U3631 ( .A1(n2837), .A2(n3011), .ZN(n2824) );
  NAND2_X1 U3632 ( .A1(n2825), .A2(n3632), .ZN(n2849) );
  INV_X1 U3633 ( .A(n2826), .ZN(n2827) );
  AND2_X1 U3634 ( .A1(n4380), .A2(n2827), .ZN(n2828) );
  NAND2_X1 U3635 ( .A1(n2829), .A2(n2828), .ZN(n2841) );
  NOR2_X1 U3636 ( .A1(n2841), .A2(n2982), .ZN(n2830) );
  AOI22_X1 U3637 ( .A1(n3740), .A2(n3626), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n2831) );
  INV_X1 U3638 ( .A(n2831), .ZN(n2847) );
  NOR2_X1 U3639 ( .A1(n2841), .A2(n4287), .ZN(n2832) );
  INV_X1 U3640 ( .A(n2833), .ZN(n2842) );
  NAND2_X1 U3641 ( .A1(n3041), .A2(n4170), .ZN(n2834) );
  OR2_X1 U3642 ( .A1(n2842), .A2(n2834), .ZN(n2836) );
  AOI22_X1 U3643 ( .A1(n3962), .A2(n3623), .B1(n3907), .B2(n3625), .ZN(n2845)
         );
  NAND2_X1 U3644 ( .A1(n2837), .A2(n4139), .ZN(n2838) );
  NAND2_X1 U3645 ( .A1(n2842), .A2(n2838), .ZN(n2839) );
  NAND2_X1 U3646 ( .A1(n2839), .A2(n3040), .ZN(n3012) );
  NAND2_X1 U3647 ( .A1(n2615), .A2(n2877), .ZN(n2840) );
  OAI21_X1 U3648 ( .B1(n3012), .B2(n2840), .A(STATE_REG_SCAN_IN), .ZN(n2843)
         );
  INV_X1 U3649 ( .A(n2841), .ZN(n3797) );
  NAND2_X1 U3650 ( .A1(n2842), .A2(n3797), .ZN(n3010) );
  OR2_X1 U3651 ( .A1(n3930), .A2(n3630), .ZN(n2844) );
  NAND2_X1 U3652 ( .A1(n2849), .A2(n2848), .ZN(U3217) );
  INV_X1 U3653 ( .A(n4380), .ZN(n2850) );
  INV_X1 U3654 ( .A(DATAI_1_), .ZN(n2851) );
  MUX2_X1 U3655 ( .A(n2886), .B(n2851), .S(U3149), .Z(n2852) );
  INV_X1 U3656 ( .A(n2852), .ZN(U3351) );
  INV_X1 U3657 ( .A(DATAI_13_), .ZN(n2854) );
  NAND2_X1 U3658 ( .A1(n3853), .A2(STATE_REG_SCAN_IN), .ZN(n2853) );
  OAI21_X1 U3659 ( .B1(STATE_REG_SCAN_IN), .B2(n2854), .A(n2853), .ZN(U3339)
         );
  MUX2_X1 U3660 ( .A(n2327), .B(n3001), .S(STATE_REG_SCAN_IN), .Z(n2855) );
  INV_X1 U3661 ( .A(n2855), .ZN(U3344) );
  INV_X1 U3662 ( .A(DATAI_18_), .ZN(n4450) );
  NAND2_X1 U3663 ( .A1(n3895), .A2(STATE_REG_SCAN_IN), .ZN(n2856) );
  OAI21_X1 U3664 ( .B1(STATE_REG_SCAN_IN), .B2(n4450), .A(n2856), .ZN(U3334)
         );
  INV_X1 U3665 ( .A(DATAI_26_), .ZN(n2859) );
  NAND2_X1 U3666 ( .A1(n2857), .A2(STATE_REG_SCAN_IN), .ZN(n2858) );
  OAI21_X1 U3667 ( .B1(STATE_REG_SCAN_IN), .B2(n2859), .A(n2858), .ZN(U3326)
         );
  INV_X1 U3668 ( .A(n2860), .ZN(n2861) );
  NAND2_X1 U3669 ( .A1(n2861), .A2(STATE_REG_SCAN_IN), .ZN(n2862) );
  OAI21_X1 U3670 ( .B1(STATE_REG_SCAN_IN), .B2(n2493), .A(n2862), .ZN(U3327)
         );
  NAND2_X1 U3671 ( .A1(n3790), .A2(STATE_REG_SCAN_IN), .ZN(n2863) );
  OAI21_X1 U3672 ( .B1(STATE_REG_SCAN_IN), .B2(n2452), .A(n2863), .ZN(U3332)
         );
  INV_X1 U3673 ( .A(DATAI_21_), .ZN(n2865) );
  NAND2_X1 U3674 ( .A1(n2530), .A2(STATE_REG_SCAN_IN), .ZN(n2864) );
  OAI21_X1 U3675 ( .B1(STATE_REG_SCAN_IN), .B2(n2865), .A(n2864), .ZN(U3331)
         );
  INV_X1 U3676 ( .A(DATAI_30_), .ZN(n2868) );
  NAND2_X1 U3677 ( .A1(n2866), .A2(STATE_REG_SCAN_IN), .ZN(n2867) );
  OAI21_X1 U3678 ( .B1(STATE_REG_SCAN_IN), .B2(n2868), .A(n2867), .ZN(U3322)
         );
  INV_X1 U3679 ( .A(DATAI_31_), .ZN(n4446) );
  OR4_X1 U3680 ( .A1(n2870), .A2(IR_REG_30__SCAN_IN), .A3(n2869), .A4(U3149), 
        .ZN(n2871) );
  OAI21_X1 U3681 ( .B1(STATE_REG_SCAN_IN), .B2(n4446), .A(n2871), .ZN(U3321)
         );
  INV_X1 U3682 ( .A(D_REG_1__SCAN_IN), .ZN(n4472) );
  INV_X1 U3683 ( .A(n2873), .ZN(n2874) );
  AOI22_X1 U3684 ( .A1(n4378), .A2(n4472), .B1(n2874), .B2(n4380), .ZN(U3459)
         );
  INV_X1 U3685 ( .A(D_REG_0__SCAN_IN), .ZN(n4578) );
  INV_X1 U3686 ( .A(n2875), .ZN(n2876) );
  AOI22_X1 U3687 ( .A1(n4378), .A2(n4578), .B1(n2876), .B2(n4380), .ZN(U3458)
         );
  OR2_X1 U3688 ( .A1(n2877), .A2(U3149), .ZN(n3800) );
  NAND2_X1 U3689 ( .A1(n3011), .A2(n3800), .ZN(n2881) );
  AOI21_X1 U3690 ( .B1(n2878), .B2(n2877), .A(n2326), .ZN(n2880) );
  INV_X1 U3691 ( .A(n2880), .ZN(n2879) );
  NOR2_X1 U3692 ( .A1(n4345), .A2(n2897), .ZN(U3148) );
  NOR2_X1 U3693 ( .A1(n2883), .A2(n2882), .ZN(n4275) );
  INV_X1 U3694 ( .A(n4275), .ZN(n2984) );
  XNOR2_X1 U3695 ( .A(n2886), .B(REG1_REG_1__SCAN_IN), .ZN(n3819) );
  AND2_X1 U3696 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3818)
         );
  NAND2_X1 U3697 ( .A1(n3819), .A2(n3818), .ZN(n3817) );
  NAND2_X1 U3698 ( .A1(n3820), .A2(REG1_REG_1__SCAN_IN), .ZN(n2884) );
  NAND2_X1 U3699 ( .A1(n3817), .A2(n2884), .ZN(n3825) );
  INV_X1 U3700 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3080) );
  XNOR2_X1 U3701 ( .A(n4286), .B(n3080), .ZN(n3826) );
  NAND2_X1 U3702 ( .A1(n4286), .A2(REG1_REG_2__SCAN_IN), .ZN(n2885) );
  XOR2_X1 U3703 ( .A(n2905), .B(REG1_REG_3__SCAN_IN), .Z(n2893) );
  AND2_X1 U3704 ( .A1(n2982), .A2(n4275), .ZN(n3796) );
  AND2_X1 U3705 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3816)
         );
  NAND2_X1 U3706 ( .A1(n3820), .A2(REG2_REG_1__SCAN_IN), .ZN(n3829) );
  NAND2_X1 U3707 ( .A1(n3830), .A2(n3829), .ZN(n2890) );
  MUX2_X1 U3708 ( .A(REG2_REG_2__SCAN_IN), .B(n2888), .S(n4286), .Z(n2889) );
  NAND2_X1 U3709 ( .A1(n2890), .A2(n2889), .ZN(n3832) );
  NAND2_X1 U3710 ( .A1(n4286), .A2(REG2_REG_2__SCAN_IN), .ZN(n2891) );
  NAND2_X1 U3711 ( .A1(n3832), .A2(n2891), .ZN(n2915) );
  XNOR2_X1 U3712 ( .A(n2915), .B(n2896), .ZN(n2914) );
  XOR2_X1 U3713 ( .A(REG2_REG_3__SCAN_IN), .B(n2914), .Z(n2892) );
  AOI22_X1 U3714 ( .A1(n4353), .A2(n2893), .B1(n4355), .B2(n2892), .ZN(n2895)
         );
  INV_X1 U3715 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4462) );
  NOR2_X1 U3716 ( .A1(STATE_REG_SCAN_IN), .A2(n4462), .ZN(n3057) );
  AOI21_X1 U3717 ( .B1(n4345), .B2(ADDR_REG_3__SCAN_IN), .A(n3057), .ZN(n2894)
         );
  OAI211_X1 U3718 ( .C1(n2896), .C2(n4358), .A(n2895), .B(n2894), .ZN(U3243)
         );
  INV_X1 U3719 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n4561) );
  NAND2_X1 U3720 ( .A1(n4147), .A2(U4043), .ZN(n2898) );
  OAI21_X1 U3721 ( .B1(n2897), .B2(n4561), .A(n2898), .ZN(U3566) );
  INV_X1 U3722 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n4566) );
  NAND2_X1 U3723 ( .A1(n3567), .A2(U4043), .ZN(n2899) );
  OAI21_X1 U3724 ( .B1(n2897), .B2(n4566), .A(n2899), .ZN(U3553) );
  INV_X1 U3725 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n4563) );
  NAND2_X1 U3726 ( .A1(n3482), .A2(U4043), .ZN(n2900) );
  OAI21_X1 U3727 ( .B1(n2897), .B2(n4563), .A(n2900), .ZN(U3559) );
  INV_X1 U3728 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n4533) );
  NAND2_X1 U3729 ( .A1(n4130), .A2(U4043), .ZN(n2901) );
  OAI21_X1 U3730 ( .B1(U4043), .B2(n4533), .A(n2901), .ZN(U3569) );
  INV_X1 U3731 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n4564) );
  NAND2_X1 U3732 ( .A1(n3569), .A2(U4043), .ZN(n2902) );
  OAI21_X1 U3733 ( .B1(U4043), .B2(n4564), .A(n2902), .ZN(U3555) );
  INV_X1 U3734 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n4560) );
  NAND2_X1 U3735 ( .A1(n4101), .A2(U4043), .ZN(n2903) );
  OAI21_X1 U3736 ( .B1(U4043), .B2(n4560), .A(n2903), .ZN(U3570) );
  INV_X1 U3737 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n4565) );
  NAND2_X1 U3738 ( .A1(n3484), .A2(U4043), .ZN(n2904) );
  OAI21_X1 U3739 ( .B1(n2897), .B2(n4565), .A(n2904), .ZN(U3561) );
  NAND2_X1 U3740 ( .A1(n2906), .A2(n4285), .ZN(n2907) );
  NAND2_X1 U3741 ( .A1(n2908), .A2(n2907), .ZN(n2909) );
  INV_X1 U3742 ( .A(n4284), .ZN(n2919) );
  XNOR2_X1 U3743 ( .A(n2909), .B(n2919), .ZN(n2987) );
  NAND2_X1 U3744 ( .A1(n2987), .A2(REG1_REG_4__SCAN_IN), .ZN(n2911) );
  NAND2_X1 U3745 ( .A1(n2909), .A2(n4284), .ZN(n2910) );
  NAND2_X1 U3746 ( .A1(n2911), .A2(n2910), .ZN(n3840) );
  INV_X1 U3747 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2912) );
  MUX2_X1 U3748 ( .A(n2912), .B(REG1_REG_5__SCAN_IN), .S(n4282), .Z(n3841) );
  NAND2_X1 U3749 ( .A1(n3840), .A2(n3841), .ZN(n3839) );
  OR2_X1 U3750 ( .A1(n4282), .A2(n2912), .ZN(n2913) );
  INV_X1 U3751 ( .A(n4281), .ZN(n2923) );
  XNOR2_X1 U3752 ( .A(n2929), .B(n2923), .ZN(n2928) );
  XNOR2_X1 U3753 ( .A(n2928), .B(REG1_REG_6__SCAN_IN), .ZN(n2927) );
  NAND2_X1 U3754 ( .A1(n2914), .A2(REG2_REG_3__SCAN_IN), .ZN(n2917) );
  NAND2_X1 U3755 ( .A1(n2915), .A2(n4285), .ZN(n2916) );
  NAND2_X1 U3756 ( .A1(n2917), .A2(n2916), .ZN(n2918) );
  XNOR2_X1 U3757 ( .A(n2918), .B(n4284), .ZN(n2988) );
  INV_X1 U3758 ( .A(n2918), .ZN(n2920) );
  OAI22_X1 U3759 ( .A1(n2988), .A2(n2921), .B1(n2920), .B2(n2919), .ZN(n3843)
         );
  MUX2_X1 U3760 ( .A(n3157), .B(REG2_REG_5__SCAN_IN), .S(n4282), .Z(n3844) );
  NAND2_X1 U3761 ( .A1(n3843), .A2(n3844), .ZN(n3842) );
  OAI21_X1 U3762 ( .B1(n4282), .B2(n3157), .A(n3842), .ZN(n2934) );
  XOR2_X1 U3763 ( .A(REG2_REG_6__SCAN_IN), .B(n2935), .Z(n2925) );
  AND2_X1 U3764 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3204) );
  AOI21_X1 U3765 ( .B1(n4345), .B2(ADDR_REG_6__SCAN_IN), .A(n3204), .ZN(n2922)
         );
  OAI21_X1 U3766 ( .B1(n4358), .B2(n2923), .A(n2922), .ZN(n2924) );
  AOI21_X1 U3767 ( .B1(n4355), .B2(n2925), .A(n2924), .ZN(n2926) );
  OAI21_X1 U3768 ( .B1(n2927), .B2(n4321), .A(n2926), .ZN(U3246) );
  INV_X1 U3769 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4437) );
  MUX2_X1 U3770 ( .A(n4437), .B(REG1_REG_7__SCAN_IN), .S(n4280), .Z(n2932) );
  NAND2_X1 U3771 ( .A1(n2928), .A2(REG1_REG_6__SCAN_IN), .ZN(n2931) );
  NAND2_X1 U3772 ( .A1(n2929), .A2(n4281), .ZN(n2930) );
  XOR2_X1 U3773 ( .A(n2932), .B(n2953), .Z(n2941) );
  AND2_X1 U3774 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3224) );
  AOI21_X1 U3775 ( .B1(n4345), .B2(ADDR_REG_7__SCAN_IN), .A(n3224), .ZN(n2933)
         );
  INV_X1 U3776 ( .A(n2933), .ZN(n2939) );
  MUX2_X1 U3777 ( .A(n2305), .B(REG2_REG_7__SCAN_IN), .S(n4280), .Z(n2936) );
  INV_X1 U3778 ( .A(n4355), .ZN(n4324) );
  AOI211_X1 U3779 ( .C1(n2937), .C2(n2936), .A(n4324), .B(n2950), .ZN(n2938)
         );
  AOI211_X1 U3780 ( .C1(n4330), .C2(n4280), .A(n2939), .B(n2938), .ZN(n2940)
         );
  OAI21_X1 U3781 ( .B1(n4321), .B2(n2941), .A(n2940), .ZN(U3247) );
  AOI21_X1 U3782 ( .B1(n4275), .B2(n2942), .A(n4287), .ZN(n2986) );
  NOR2_X1 U3783 ( .A1(n4275), .A2(REG1_REG_0__SCAN_IN), .ZN(n2943) );
  OAI21_X1 U3784 ( .B1(IR_REG_0__SCAN_IN), .B2(n2943), .A(n2986), .ZN(n2944)
         );
  OAI211_X1 U3785 ( .C1(n2986), .C2(IR_REG_0__SCAN_IN), .A(n2945), .B(n2944), 
        .ZN(n2946) );
  OAI21_X1 U3786 ( .B1(STATE_REG_SCAN_IN), .B2(n3018), .A(n2946), .ZN(n2948)
         );
  INV_X1 U3787 ( .A(IR_REG_0__SCAN_IN), .ZN(n4390) );
  NOR3_X1 U3788 ( .A1(n4321), .A2(REG1_REG_0__SCAN_IN), .A3(n4390), .ZN(n2947)
         );
  AOI211_X1 U3789 ( .C1(n4345), .C2(ADDR_REG_0__SCAN_IN), .A(n2948), .B(n2947), 
        .ZN(n2949) );
  INV_X1 U3790 ( .A(n2949), .ZN(U3240) );
  XNOR2_X1 U3791 ( .A(n2996), .B(n3001), .ZN(n2997) );
  XNOR2_X1 U3792 ( .A(n2997), .B(REG2_REG_8__SCAN_IN), .ZN(n2959) );
  AND2_X1 U3793 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3273) );
  AOI21_X1 U3794 ( .B1(n4345), .B2(ADDR_REG_8__SCAN_IN), .A(n3273), .ZN(n2951)
         );
  OAI21_X1 U3795 ( .B1(n4358), .B2(n3001), .A(n2951), .ZN(n2958) );
  INV_X1 U3796 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2956) );
  AND2_X1 U3797 ( .A1(n4280), .A2(REG1_REG_7__SCAN_IN), .ZN(n2952) );
  OR2_X1 U3798 ( .A1(n4280), .A2(REG1_REG_7__SCAN_IN), .ZN(n2954) );
  NOR2_X1 U3799 ( .A1(n2955), .A2(n2956), .ZN(n3002) );
  AOI211_X1 U3800 ( .C1(n2956), .C2(n2955), .A(n4321), .B(n3002), .ZN(n2957)
         );
  AOI211_X1 U3801 ( .C1(n4355), .C2(n2959), .A(n2958), .B(n2957), .ZN(n2960)
         );
  INV_X1 U3802 ( .A(n2960), .ZN(U3248) );
  INV_X1 U3803 ( .A(n4425), .ZN(n4402) );
  NAND2_X1 U3804 ( .A1(n3814), .A2(n2616), .ZN(n3676) );
  AND2_X1 U3805 ( .A1(n3674), .A2(n3676), .ZN(n3759) );
  INV_X1 U3806 ( .A(n3759), .ZN(n4372) );
  INV_X1 U3807 ( .A(n2607), .ZN(n2961) );
  NOR2_X1 U3808 ( .A1(n2616), .A2(n2961), .ZN(n4370) );
  INV_X1 U3809 ( .A(n4080), .ZN(n2962) );
  NOR2_X1 U3810 ( .A1(n2962), .A2(n4126), .ZN(n2963) );
  AOI211_X1 U3811 ( .C1(n4402), .C2(n4372), .A(n4370), .B(n4368), .ZN(n4392)
         );
  NAND2_X1 U3812 ( .A1(n4441), .A2(REG1_REG_0__SCAN_IN), .ZN(n2964) );
  OAI21_X1 U3813 ( .B1(n4392), .B2(n4441), .A(n2964), .ZN(U3518) );
  OR2_X1 U3814 ( .A1(n3755), .A2(n2965), .ZN(n2966) );
  NAND2_X1 U3815 ( .A1(n2967), .A2(n2966), .ZN(n3049) );
  NAND2_X1 U3816 ( .A1(n3814), .A2(n4148), .ZN(n2969) );
  NAND2_X1 U3817 ( .A1(n2254), .A2(n4129), .ZN(n2968) );
  OAI211_X1 U3818 ( .C1(n4139), .C2(n2974), .A(n2969), .B(n2968), .ZN(n2970)
         );
  INV_X1 U3819 ( .A(n2970), .ZN(n2973) );
  XNOR2_X1 U3820 ( .A(n3755), .B(n3674), .ZN(n2971) );
  NAND2_X1 U3821 ( .A1(n2971), .A2(n4126), .ZN(n2972) );
  OAI211_X1 U3822 ( .C1(n3049), .C2(n4080), .A(n2973), .B(n2972), .ZN(n3045)
         );
  OAI21_X1 U3823 ( .B1(n2616), .B2(n2974), .A(n3074), .ZN(n3053) );
  OAI22_X1 U3824 ( .A1(n3049), .A2(n4425), .B1(n4424), .B2(n3053), .ZN(n2975)
         );
  NOR2_X1 U3825 ( .A1(n3045), .A2(n2975), .ZN(n4394) );
  NAND2_X1 U3826 ( .A1(n4441), .A2(REG1_REG_1__SCAN_IN), .ZN(n2976) );
  OAI21_X1 U3827 ( .B1(n4394), .B2(n4441), .A(n2976), .ZN(U3519) );
  INV_X1 U3828 ( .A(n2977), .ZN(n2981) );
  NOR2_X1 U3829 ( .A1(n2979), .A2(n2978), .ZN(n2980) );
  NOR2_X1 U3830 ( .A1(n2981), .A2(n2980), .ZN(n3014) );
  NAND2_X1 U3831 ( .A1(n3014), .A2(n2984), .ZN(n2983) );
  OAI211_X1 U3832 ( .C1(n3816), .C2(n2984), .A(n2983), .B(n2982), .ZN(n2985)
         );
  OAI211_X1 U3833 ( .C1(IR_REG_0__SCAN_IN), .C2(n2986), .A(n2985), .B(U4043), 
        .ZN(n3836) );
  XOR2_X1 U3834 ( .A(n2987), .B(REG1_REG_4__SCAN_IN), .Z(n2994) );
  NAND2_X1 U3835 ( .A1(n4345), .A2(ADDR_REG_4__SCAN_IN), .ZN(n2992) );
  NAND2_X1 U3836 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3565) );
  XNOR2_X1 U3837 ( .A(n2988), .B(REG2_REG_4__SCAN_IN), .ZN(n2989) );
  NAND2_X1 U3838 ( .A1(n4355), .A2(n2989), .ZN(n2991) );
  NAND2_X1 U3839 ( .A1(n4330), .A2(n4284), .ZN(n2990) );
  NAND4_X1 U3840 ( .A1(n2992), .A2(n3565), .A3(n2991), .A4(n2990), .ZN(n2993)
         );
  AOI21_X1 U3841 ( .B1(n4353), .B2(n2994), .A(n2993), .ZN(n2995) );
  NAND2_X1 U3842 ( .A1(n3836), .A2(n2995), .ZN(U3244) );
  INV_X1 U3843 ( .A(n4279), .ZN(n3292) );
  OAI22_X1 U3844 ( .A1(n2997), .A2(n3190), .B1(n2996), .B2(n3001), .ZN(n2999)
         );
  MUX2_X1 U3845 ( .A(REG2_REG_9__SCAN_IN), .B(n3180), .S(n4279), .Z(n2998) );
  NAND2_X1 U3846 ( .A1(n2999), .A2(n2998), .ZN(n3291) );
  OAI211_X1 U3847 ( .C1(n2999), .C2(n2998), .A(n3291), .B(n4355), .ZN(n3009)
         );
  NOR2_X1 U3848 ( .A1(STATE_REG_SCAN_IN), .A2(n4461), .ZN(n3283) );
  INV_X1 U3849 ( .A(n3000), .ZN(n3004) );
  INV_X1 U3850 ( .A(n3001), .ZN(n3003) );
  MUX2_X1 U3851 ( .A(n4439), .B(REG1_REG_9__SCAN_IN), .S(n4279), .Z(n3005) );
  NOR2_X1 U3852 ( .A1(n3006), .A2(n3005), .ZN(n3301) );
  AOI211_X1 U3853 ( .C1(n3006), .C2(n3005), .A(n3301), .B(n4321), .ZN(n3007)
         );
  AOI211_X1 U3854 ( .C1(n4345), .C2(ADDR_REG_9__SCAN_IN), .A(n3283), .B(n3007), 
        .ZN(n3008) );
  OAI211_X1 U3855 ( .C1(n4358), .C2(n3292), .A(n3009), .B(n3008), .ZN(U3249)
         );
  INV_X1 U3856 ( .A(n3010), .ZN(n3013) );
  NOR3_X1 U3857 ( .A1(n3013), .A2(n3012), .A3(n3011), .ZN(n3037) );
  AOI22_X1 U3858 ( .A1(n3014), .A2(n3632), .B1(n3626), .B2(n3813), .ZN(n3017)
         );
  NAND2_X1 U3859 ( .A1(n3625), .A2(n3015), .ZN(n3016) );
  OAI211_X1 U3860 ( .C1(n3037), .C2(n3018), .A(n3017), .B(n3016), .ZN(U3229)
         );
  INV_X1 U3861 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3028) );
  AOI211_X1 U3862 ( .C1(n3021), .C2(n3020), .A(n3617), .B(n3019), .ZN(n3022)
         );
  INV_X1 U3863 ( .A(n3022), .ZN(n3027) );
  OAI22_X1 U3864 ( .A1(n3023), .A2(n3610), .B1(n3612), .B2(n3105), .ZN(n3024)
         );
  AOI21_X1 U3865 ( .B1(n3025), .B2(n3625), .A(n3024), .ZN(n3026) );
  OAI211_X1 U3866 ( .C1(n3037), .C2(n3028), .A(n3027), .B(n3026), .ZN(U3219)
         );
  OAI21_X1 U3867 ( .B1(n3031), .B2(n3030), .A(n3029), .ZN(n3032) );
  NAND2_X1 U3868 ( .A1(n3032), .A2(n3632), .ZN(n3035) );
  AOI21_X1 U3869 ( .B1(n3073), .B2(n3625), .A(n3033), .ZN(n3034) );
  OAI211_X1 U3870 ( .C1(n3037), .C2(n3036), .A(n3035), .B(n3034), .ZN(U3234)
         );
  INV_X1 U3871 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n4535) );
  NAND2_X1 U3872 ( .A1(n3979), .A2(U4043), .ZN(n3038) );
  OAI21_X1 U3873 ( .B1(n2897), .B2(n4535), .A(n3038), .ZN(U3576) );
  INV_X1 U3874 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n4558) );
  NAND2_X1 U3875 ( .A1(n3740), .A2(U4043), .ZN(n3039) );
  OAI21_X1 U3876 ( .B1(U4043), .B2(n4558), .A(n3039), .ZN(U3579) );
  NAND4_X1 U3877 ( .A1(n3043), .A2(n3042), .A3(n3041), .A4(n3040), .ZN(n3044)
         );
  NAND2_X1 U3878 ( .A1(n4375), .A2(n3900), .ZN(n3135) );
  MUX2_X1 U3880 ( .A(REG2_REG_1__SCAN_IN), .B(n3045), .S(n4375), .Z(n3046) );
  INV_X1 U3881 ( .A(n3046), .ZN(n3052) );
  NAND2_X1 U3882 ( .A1(n3047), .A2(n4277), .ZN(n3141) );
  INV_X1 U3883 ( .A(n3141), .ZN(n3048) );
  NAND2_X1 U3884 ( .A1(n4375), .A2(n3048), .ZN(n4090) );
  INV_X1 U3885 ( .A(n4090), .ZN(n4373) );
  INV_X1 U3886 ( .A(n3049), .ZN(n3050) );
  INV_X1 U3887 ( .A(n4153), .ZN(n4371) );
  AOI22_X1 U3888 ( .A1(n4373), .A2(n3050), .B1(REG3_REG_1__SCAN_IN), .B2(n4371), .ZN(n3051) );
  OAI211_X1 U3889 ( .C1(n4107), .C2(n3053), .A(n3052), .B(n3051), .ZN(U3289)
         );
  INV_X1 U3890 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n4559) );
  NAND2_X1 U3891 ( .A1(n3962), .A2(U4043), .ZN(n3054) );
  OAI21_X1 U3892 ( .B1(U4043), .B2(n4559), .A(n3054), .ZN(U3577) );
  XNOR2_X1 U3893 ( .A(n3056), .B(n3055), .ZN(n3061) );
  AOI21_X1 U3894 ( .B1(n3623), .B2(n2254), .A(n3057), .ZN(n3059) );
  AOI22_X1 U3895 ( .A1(n3626), .A2(n3812), .B1(n3625), .B2(n3103), .ZN(n3058)
         );
  OAI211_X1 U3896 ( .C1(n3630), .C2(REG3_REG_3__SCAN_IN), .A(n3059), .B(n3058), 
        .ZN(n3060) );
  AOI21_X1 U3897 ( .B1(n3061), .B2(n3632), .A(n3060), .ZN(n3062) );
  INV_X1 U3898 ( .A(n3062), .ZN(U3215) );
  INV_X1 U3899 ( .A(n3063), .ZN(n3064) );
  AOI21_X1 U3900 ( .B1(n3749), .B2(n3065), .A(n3064), .ZN(n4359) );
  OAI21_X1 U3901 ( .B1(n3749), .B2(n3067), .A(n3066), .ZN(n3072) );
  AOI22_X1 U3902 ( .A1(n3813), .A2(n4148), .B1(n3073), .B2(n4170), .ZN(n3068)
         );
  OAI21_X1 U3903 ( .B1(n3069), .B2(n4140), .A(n3068), .ZN(n3071) );
  NOR2_X1 U3904 ( .A1(n4359), .A2(n4080), .ZN(n3070) );
  AOI211_X1 U3905 ( .C1(n4126), .C2(n3072), .A(n3071), .B(n3070), .ZN(n4366)
         );
  OAI21_X1 U3906 ( .B1(n4359), .B2(n4425), .A(n4366), .ZN(n3082) );
  INV_X1 U3907 ( .A(n3110), .ZN(n3076) );
  NAND2_X1 U3908 ( .A1(n3074), .A2(n3073), .ZN(n3075) );
  NAND2_X1 U3909 ( .A1(n3076), .A2(n3075), .ZN(n4360) );
  INV_X1 U3910 ( .A(REG0_REG_2__SCAN_IN), .ZN(n3077) );
  OAI22_X1 U3911 ( .A1(n4271), .A2(n4360), .B1(n4431), .B2(n3077), .ZN(n3078)
         );
  AOI21_X1 U3912 ( .B1(n3082), .B2(n4431), .A(n3078), .ZN(n3079) );
  INV_X1 U3913 ( .A(n3079), .ZN(U3471) );
  OAI22_X1 U3914 ( .A1(n4223), .A2(n4360), .B1(n4443), .B2(n3080), .ZN(n3081)
         );
  AOI21_X1 U3915 ( .B1(n3082), .B2(n4443), .A(n3081), .ZN(n3083) );
  INV_X1 U3916 ( .A(n3083), .ZN(U3520) );
  AND2_X1 U3917 ( .A1(n3693), .A2(n3689), .ZN(n3746) );
  OR2_X1 U3918 ( .A1(n3084), .A2(n3085), .ZN(n3087) );
  NAND2_X1 U3919 ( .A1(n3087), .A2(n3086), .ZN(n3088) );
  XOR2_X1 U3920 ( .A(n3746), .B(n3088), .Z(n3166) );
  XNOR2_X1 U3921 ( .A(n3089), .B(n3746), .ZN(n3093) );
  AOI22_X1 U3922 ( .A1(n3810), .A2(n4129), .B1(n3205), .B2(n4170), .ZN(n3090)
         );
  OAI21_X1 U3923 ( .B1(n3091), .B2(n4133), .A(n3090), .ZN(n3092) );
  AOI21_X1 U3924 ( .B1(n3093), .B2(n4126), .A(n3092), .ZN(n3171) );
  OAI21_X1 U3925 ( .B1(n3166), .B2(n4411), .A(n3171), .ZN(n3099) );
  NAND2_X1 U3926 ( .A1(n3161), .A2(n3205), .ZN(n3094) );
  NAND2_X1 U3927 ( .A1(n3136), .A2(n3094), .ZN(n3165) );
  INV_X1 U3928 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3095) );
  OAI22_X1 U3929 ( .A1(n3165), .A2(n4223), .B1(n4443), .B2(n3095), .ZN(n3096)
         );
  AOI21_X1 U3930 ( .B1(n3099), .B2(n4443), .A(n3096), .ZN(n3097) );
  INV_X1 U3931 ( .A(n3097), .ZN(U3524) );
  INV_X1 U3932 ( .A(REG0_REG_6__SCAN_IN), .ZN(n4576) );
  OAI22_X1 U3933 ( .A1(n3165), .A2(n4271), .B1(n4431), .B2(n4576), .ZN(n3098)
         );
  AOI21_X1 U3934 ( .B1(n3099), .B2(n4431), .A(n3098), .ZN(n3100) );
  INV_X1 U3935 ( .A(n3100), .ZN(U3479) );
  XNOR2_X1 U3936 ( .A(n3101), .B(n3757), .ZN(n4396) );
  XNOR2_X1 U3937 ( .A(n3102), .B(n3757), .ZN(n3107) );
  AOI22_X1 U3938 ( .A1(n3812), .A2(n4129), .B1(n4170), .B2(n3103), .ZN(n3104)
         );
  OAI21_X1 U3939 ( .B1(n3105), .B2(n4133), .A(n3104), .ZN(n3106) );
  AOI21_X1 U3940 ( .B1(n3107), .B2(n4126), .A(n3106), .ZN(n3108) );
  OAI21_X1 U3941 ( .B1(n4396), .B2(n4080), .A(n3108), .ZN(n4398) );
  INV_X1 U3942 ( .A(n4398), .ZN(n3115) );
  INV_X1 U3943 ( .A(n4396), .ZN(n3113) );
  OAI21_X1 U3944 ( .B1(n3110), .B2(n3109), .A(n3116), .ZN(n4395) );
  AOI22_X1 U3945 ( .A1(n4377), .A2(REG2_REG_3__SCAN_IN), .B1(n4371), .B2(n4462), .ZN(n3111) );
  OAI21_X1 U3946 ( .B1(n4107), .B2(n4395), .A(n3111), .ZN(n3112) );
  AOI21_X1 U3947 ( .B1(n3113), .B2(n4373), .A(n3112), .ZN(n3114) );
  OAI21_X1 U3948 ( .B1(n3115), .B2(n4377), .A(n3114), .ZN(U3287) );
  AOI211_X1 U3949 ( .C1(n3568), .C2(n3116), .A(n4424), .B(n3159), .ZN(n4401)
         );
  NOR2_X1 U3950 ( .A1(n4153), .A2(n3570), .ZN(n3125) );
  XNOR2_X1 U3951 ( .A(n3118), .B(n3750), .ZN(n3123) );
  OR2_X1 U3952 ( .A1(n3084), .A2(n3750), .ZN(n3150) );
  NAND2_X1 U3953 ( .A1(n3084), .A2(n3750), .ZN(n3119) );
  NAND2_X1 U3954 ( .A1(n3150), .A2(n3119), .ZN(n3126) );
  AOI22_X1 U3955 ( .A1(n3567), .A2(n4148), .B1(n3568), .B2(n4170), .ZN(n3121)
         );
  NAND2_X1 U3956 ( .A1(n3569), .A2(n4129), .ZN(n3120) );
  OAI211_X1 U3957 ( .C1(n3126), .C2(n4080), .A(n3121), .B(n3120), .ZN(n3122)
         );
  AOI21_X1 U3958 ( .B1(n3123), .B2(n4126), .A(n3122), .ZN(n3124) );
  INV_X1 U3959 ( .A(n3124), .ZN(n4400) );
  AOI211_X1 U3960 ( .C1(n4401), .C2(n3900), .A(n3125), .B(n4400), .ZN(n3128)
         );
  INV_X1 U3961 ( .A(n3126), .ZN(n4403) );
  AOI22_X1 U3962 ( .A1(n4403), .A2(n4373), .B1(REG2_REG_4__SCAN_IN), .B2(n4377), .ZN(n3127) );
  OAI21_X1 U3963 ( .B1(n3128), .B2(n4377), .A(n3127), .ZN(U3286) );
  XNOR2_X1 U3964 ( .A(n3748), .B(n3129), .ZN(n3134) );
  OAI22_X1 U3965 ( .A1(n3131), .A2(n4140), .B1(n4139), .B2(n3130), .ZN(n3132)
         );
  AOI21_X1 U3966 ( .B1(n4148), .B2(n3811), .A(n3132), .ZN(n3133) );
  OAI21_X1 U3967 ( .B1(n3134), .B2(n4143), .A(n3133), .ZN(n4413) );
  INV_X1 U3968 ( .A(n4413), .ZN(n3147) );
  INV_X1 U3969 ( .A(n3135), .ZN(n4123) );
  NAND2_X1 U3970 ( .A1(n3136), .A2(n3225), .ZN(n3137) );
  NAND2_X1 U3971 ( .A1(n3137), .A2(n2619), .ZN(n3138) );
  NOR2_X1 U3972 ( .A1(n3187), .A2(n3138), .ZN(n4414) );
  OAI22_X1 U3973 ( .A1(n4375), .A2(n2305), .B1(n3228), .B2(n4153), .ZN(n3145)
         );
  NOR2_X1 U3974 ( .A1(n3139), .A2(n3748), .ZN(n4412) );
  INV_X1 U3975 ( .A(n3140), .ZN(n3143) );
  NAND2_X1 U3976 ( .A1(n4080), .A2(n3141), .ZN(n3142) );
  NOR3_X1 U3977 ( .A1(n4412), .A2(n3143), .A3(n4137), .ZN(n3144) );
  AOI211_X1 U3978 ( .C1(n4123), .C2(n4414), .A(n3145), .B(n3144), .ZN(n3146)
         );
  OAI21_X1 U3979 ( .B1(n4377), .B2(n3147), .A(n3146), .ZN(U3283) );
  INV_X1 U3980 ( .A(n3148), .ZN(n3686) );
  AND2_X1 U3981 ( .A1(n3686), .A2(n3691), .ZN(n3745) );
  NAND2_X1 U3982 ( .A1(n3150), .A2(n3149), .ZN(n3151) );
  XOR2_X1 U3983 ( .A(n3745), .B(n3151), .Z(n4406) );
  XOR2_X1 U3984 ( .A(n3745), .B(n3152), .Z(n3156) );
  AOI22_X1 U3985 ( .A1(n3811), .A2(n4129), .B1(n4170), .B2(n3537), .ZN(n3153)
         );
  OAI21_X1 U3986 ( .B1(n3154), .B2(n4133), .A(n3153), .ZN(n3155) );
  AOI21_X1 U3987 ( .B1(n3156), .B2(n4126), .A(n3155), .ZN(n4405) );
  MUX2_X1 U3988 ( .A(n4405), .B(n3157), .S(n4377), .Z(n3164) );
  OR2_X1 U3989 ( .A1(n3159), .A2(n3158), .ZN(n3160) );
  AND2_X1 U3990 ( .A1(n3161), .A2(n3160), .ZN(n4409) );
  INV_X1 U3991 ( .A(n3538), .ZN(n3162) );
  AOI22_X1 U3992 ( .A1(n4362), .A2(n4409), .B1(n3162), .B2(n4371), .ZN(n3163)
         );
  OAI211_X1 U3993 ( .C1(n4137), .C2(n4406), .A(n3164), .B(n3163), .ZN(U3285)
         );
  INV_X1 U3994 ( .A(n3165), .ZN(n3169) );
  OAI22_X1 U3995 ( .A1(n4375), .A2(n2294), .B1(n3208), .B2(n4153), .ZN(n3168)
         );
  NOR2_X1 U3996 ( .A1(n3166), .A2(n4137), .ZN(n3167) );
  AOI211_X1 U3997 ( .C1(n3169), .C2(n4362), .A(n3168), .B(n3167), .ZN(n3170)
         );
  OAI21_X1 U3998 ( .B1(n4377), .B2(n3171), .A(n3170), .ZN(U3284) );
  INV_X1 U3999 ( .A(n3172), .ZN(n3703) );
  NAND2_X1 U4000 ( .A1(n3703), .A2(n3700), .ZN(n3774) );
  XNOR2_X1 U4001 ( .A(n3173), .B(n3774), .ZN(n3177) );
  NAND2_X1 U4002 ( .A1(n3809), .A2(n4148), .ZN(n3175) );
  NAND2_X1 U4003 ( .A1(n3808), .A2(n4129), .ZN(n3174) );
  OAI211_X1 U4004 ( .C1(n4139), .C2(n3178), .A(n3175), .B(n3174), .ZN(n3176)
         );
  AOI21_X1 U4005 ( .B1(n3177), .B2(n4126), .A(n3176), .ZN(n4421) );
  OR2_X1 U4006 ( .A1(n3188), .A2(n3178), .ZN(n3179) );
  AND2_X1 U4007 ( .A1(n3237), .A2(n3179), .ZN(n4419) );
  OAI22_X1 U4009 ( .A1(n4375), .A2(n3180), .B1(n3287), .B2(n4153), .ZN(n3181)
         );
  AOI21_X1 U4010 ( .B1(n4419), .B2(n4362), .A(n3181), .ZN(n3185) );
  INV_X1 U4011 ( .A(n3774), .ZN(n3183) );
  XNOR2_X1 U4012 ( .A(n3182), .B(n3183), .ZN(n4418) );
  INV_X1 U4013 ( .A(n4137), .ZN(n4160) );
  NAND2_X1 U4014 ( .A1(n4418), .A2(n4160), .ZN(n3184) );
  OAI211_X1 U4015 ( .C1(n4421), .C2(n4377), .A(n3185), .B(n3184), .ZN(U3281)
         );
  NAND2_X1 U4016 ( .A1(n3699), .A2(n3695), .ZN(n3773) );
  XOR2_X1 U4017 ( .A(n3186), .B(n3773), .Z(n3213) );
  INV_X1 U4018 ( .A(n3213), .ZN(n3199) );
  INV_X1 U4019 ( .A(n3187), .ZN(n3189) );
  AOI21_X1 U4020 ( .B1(n3274), .B2(n3189), .A(n3188), .ZN(n3219) );
  OAI22_X1 U4021 ( .A1(n4375), .A2(n3190), .B1(n3277), .B2(n4153), .ZN(n3191)
         );
  AOI21_X1 U4022 ( .B1(n3219), .B2(n4362), .A(n3191), .ZN(n3198) );
  XOR2_X1 U4023 ( .A(n3773), .B(n3192), .Z(n3196) );
  OAI22_X1 U4024 ( .A1(n3234), .A2(n4140), .B1(n3193), .B2(n4139), .ZN(n3194)
         );
  AOI21_X1 U4025 ( .B1(n4148), .B2(n3810), .A(n3194), .ZN(n3195) );
  OAI21_X1 U4026 ( .B1(n3196), .B2(n4143), .A(n3195), .ZN(n3212) );
  NAND2_X1 U4027 ( .A1(n3212), .A2(n4375), .ZN(n3197) );
  OAI211_X1 U4028 ( .C1(n3199), .C2(n4137), .A(n3198), .B(n3197), .ZN(U3282)
         );
  XNOR2_X1 U4029 ( .A(n3202), .B(n3201), .ZN(n3203) );
  XNOR2_X1 U4030 ( .A(n3200), .B(n3203), .ZN(n3210) );
  AOI21_X1 U4031 ( .B1(n3623), .B2(n3569), .A(n3204), .ZN(n3207) );
  AOI22_X1 U4032 ( .A1(n3626), .A2(n3810), .B1(n3625), .B2(n3205), .ZN(n3206)
         );
  OAI211_X1 U4033 ( .C1(n3630), .C2(n3208), .A(n3207), .B(n3206), .ZN(n3209)
         );
  AOI21_X1 U4034 ( .B1(n3210), .B2(n3632), .A(n3209), .ZN(n3211) );
  INV_X1 U4035 ( .A(n3211), .ZN(U3236) );
  AOI21_X1 U4036 ( .B1(n3213), .B2(n4417), .A(n3212), .ZN(n3221) );
  INV_X1 U4037 ( .A(n4271), .ZN(n3216) );
  INV_X1 U4038 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3214) );
  NOR2_X1 U4039 ( .A1(n4431), .A2(n3214), .ZN(n3215) );
  AOI21_X1 U4040 ( .B1(n3219), .B2(n3216), .A(n3215), .ZN(n3217) );
  OAI21_X1 U4041 ( .B1(n3221), .B2(n4429), .A(n3217), .ZN(U3483) );
  INV_X1 U4042 ( .A(n4223), .ZN(n3218) );
  AOI22_X1 U40430 ( .A1(n3219), .A2(n3218), .B1(n4441), .B2(
        REG1_REG_8__SCAN_IN), .ZN(n3220) );
  OAI21_X1 U4044 ( .B1(n3221), .B2(n4441), .A(n3220), .ZN(U3526) );
  XOR2_X1 U4045 ( .A(n3222), .B(n3223), .Z(n3230) );
  AOI21_X1 U4046 ( .B1(n3626), .B2(n3809), .A(n3224), .ZN(n3227) );
  AOI22_X1 U4047 ( .A1(n3623), .A2(n3811), .B1(n3625), .B2(n3225), .ZN(n3226)
         );
  OAI211_X1 U4048 ( .C1(n3630), .C2(n3228), .A(n3227), .B(n3226), .ZN(n3229)
         );
  AOI21_X1 U4049 ( .B1(n3230), .B2(n3632), .A(n3229), .ZN(n3231) );
  INV_X1 U4050 ( .A(n3231), .ZN(U3210) );
  NAND2_X1 U4051 ( .A1(n3702), .A2(n3705), .ZN(n3771) );
  XOR2_X1 U4052 ( .A(n3771), .B(n3232), .Z(n3236) );
  AOI22_X1 U4053 ( .A1(n3484), .A2(n4129), .B1(n4170), .B2(n3483), .ZN(n3233)
         );
  OAI21_X1 U4054 ( .B1(n3234), .B2(n4133), .A(n3233), .ZN(n3235) );
  AOI21_X1 U4055 ( .B1(n3236), .B2(n4126), .A(n3235), .ZN(n3245) );
  NAND2_X1 U4056 ( .A1(n3237), .A2(n3483), .ZN(n3238) );
  NAND2_X1 U4057 ( .A1(n3342), .A2(n3238), .ZN(n3250) );
  INV_X1 U4058 ( .A(n3250), .ZN(n3243) );
  OAI22_X1 U4059 ( .A1(n4375), .A2(n3239), .B1(n3485), .B2(n4153), .ZN(n3242)
         );
  XOR2_X1 U4060 ( .A(n3771), .B(n3240), .Z(n3246) );
  NOR2_X1 U4061 ( .A1(n3246), .A2(n4137), .ZN(n3241) );
  AOI211_X1 U4062 ( .C1(n3243), .C2(n4362), .A(n3242), .B(n3241), .ZN(n3244)
         );
  OAI21_X1 U4063 ( .B1(n4377), .B2(n3245), .A(n3244), .ZN(U3280) );
  OAI21_X1 U4064 ( .B1(n3246), .B2(n4411), .A(n3245), .ZN(n3252) );
  INV_X1 U4065 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3247) );
  OAI22_X1 U4066 ( .A1(n3250), .A2(n4271), .B1(n4431), .B2(n3247), .ZN(n3248)
         );
  AOI21_X1 U4067 ( .B1(n3252), .B2(n4431), .A(n3248), .ZN(n3249) );
  INV_X1 U4068 ( .A(n3249), .ZN(U3487) );
  INV_X1 U4069 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4491) );
  OAI22_X1 U4070 ( .A1(n3250), .A2(n4223), .B1(n4443), .B2(n4491), .ZN(n3251)
         );
  AOI21_X1 U4071 ( .B1(n3252), .B2(n4443), .A(n3251), .ZN(n3253) );
  INV_X1 U4072 ( .A(n3253), .ZN(U3528) );
  INV_X1 U4073 ( .A(n3254), .ZN(n3255) );
  AOI21_X1 U4074 ( .B1(n3337), .B2(n3256), .A(n3255), .ZN(n3358) );
  NAND2_X1 U4075 ( .A1(n3357), .A2(n3355), .ZN(n3772) );
  XNOR2_X1 U4076 ( .A(n3358), .B(n3772), .ZN(n3261) );
  NAND2_X1 U4077 ( .A1(n3484), .A2(n4148), .ZN(n3258) );
  NAND2_X1 U4078 ( .A1(n3806), .A2(n4129), .ZN(n3257) );
  OAI211_X1 U4079 ( .C1(n4139), .C2(n3259), .A(n3258), .B(n3257), .ZN(n3260)
         );
  AOI21_X1 U4080 ( .B1(n3261), .B2(n4126), .A(n3260), .ZN(n3326) );
  INV_X1 U4081 ( .A(n3367), .ZN(n3263) );
  NAND2_X1 U4082 ( .A1(n3343), .A2(n3432), .ZN(n3262) );
  NAND2_X1 U4083 ( .A1(n3263), .A2(n3262), .ZN(n3333) );
  INV_X1 U4084 ( .A(n3333), .ZN(n3266) );
  OAI22_X1 U4085 ( .A1(n4375), .A2(n3264), .B1(n3435), .B2(n4153), .ZN(n3265)
         );
  AOI21_X1 U4086 ( .B1(n3266), .B2(n4362), .A(n3265), .ZN(n3269) );
  XNOR2_X1 U4087 ( .A(n3267), .B(n3772), .ZN(n3325) );
  NAND2_X1 U4088 ( .A1(n3325), .A2(n4160), .ZN(n3268) );
  OAI211_X1 U4089 ( .C1(n3326), .C2(n4377), .A(n3269), .B(n3268), .ZN(U3278)
         );
  NAND2_X1 U4090 ( .A1(n2046), .A2(n3271), .ZN(n3272) );
  XNOR2_X1 U4091 ( .A(n3270), .B(n3272), .ZN(n3279) );
  AOI21_X1 U4092 ( .B1(n3623), .B2(n3810), .A(n3273), .ZN(n3276) );
  AOI22_X1 U4093 ( .A1(n3626), .A2(n3482), .B1(n3625), .B2(n3274), .ZN(n3275)
         );
  OAI211_X1 U4094 ( .C1(n3630), .C2(n3277), .A(n3276), .B(n3275), .ZN(n3278)
         );
  AOI21_X1 U4095 ( .B1(n3279), .B2(n3632), .A(n3278), .ZN(n3280) );
  INV_X1 U4096 ( .A(n3280), .ZN(U3218) );
  XNOR2_X1 U4097 ( .A(n3281), .B(n3282), .ZN(n3289) );
  AOI21_X1 U4098 ( .B1(n3623), .B2(n3809), .A(n3283), .ZN(n3286) );
  AOI22_X1 U4099 ( .A1(n3626), .A2(n3808), .B1(n3625), .B2(n3284), .ZN(n3285)
         );
  OAI211_X1 U4100 ( .C1(n3630), .C2(n3287), .A(n3286), .B(n3285), .ZN(n3288)
         );
  AOI21_X1 U4101 ( .B1(n3289), .B2(n3632), .A(n3288), .ZN(n3290) );
  INV_X1 U4102 ( .A(n3290), .ZN(U3228) );
  INV_X1 U4103 ( .A(n3853), .ZN(n3311) );
  NAND2_X1 U4104 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4386), .ZN(n3295) );
  INV_X1 U4105 ( .A(n4386), .ZN(n4312) );
  AOI22_X1 U4106 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4386), .B1(n4312), .B2(
        n3346), .ZN(n4309) );
  NAND2_X1 U4107 ( .A1(n3303), .A2(n3293), .ZN(n3294) );
  INV_X1 U4108 ( .A(n3303), .ZN(n4388) );
  NAND2_X1 U4109 ( .A1(n4309), .A2(n4308), .ZN(n4307) );
  NAND2_X1 U4110 ( .A1(n4444), .A2(n3296), .ZN(n3297) );
  NOR2_X1 U4111 ( .A1(n3311), .A2(n3850), .ZN(n3298) );
  AOI21_X1 U4112 ( .B1(n3850), .B2(n3311), .A(n3298), .ZN(n3300) );
  AOI21_X1 U4113 ( .B1(n3300), .B2(n3852), .A(n4324), .ZN(n3299) );
  OAI21_X1 U4114 ( .B1(n3852), .B2(n3300), .A(n3299), .ZN(n3310) );
  INV_X1 U4115 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4572) );
  NOR2_X1 U4116 ( .A1(STATE_REG_SCAN_IN), .A2(n4572), .ZN(n3443) );
  INV_X1 U4117 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4577) );
  AOI22_X1 U4118 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4312), .B1(n4386), .B2(
        n4577), .ZN(n4303) );
  NOR2_X1 U4119 ( .A1(n4304), .A2(n4303), .ZN(n4302) );
  INV_X1 U4120 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4502) );
  NAND2_X1 U4121 ( .A1(n3853), .A2(REG1_REG_13__SCAN_IN), .ZN(n3861) );
  OAI21_X1 U4122 ( .B1(n3853), .B2(REG1_REG_13__SCAN_IN), .A(n3861), .ZN(n3306) );
  INV_X1 U4123 ( .A(n3862), .ZN(n3305) );
  AOI211_X1 U4124 ( .C1(n3307), .C2(n3306), .A(n3305), .B(n4321), .ZN(n3308)
         );
  AOI211_X1 U4125 ( .C1(n4345), .C2(ADDR_REG_13__SCAN_IN), .A(n3443), .B(n3308), .ZN(n3309) );
  OAI211_X1 U4126 ( .C1(n4358), .C2(n3311), .A(n3310), .B(n3309), .ZN(U3253)
         );
  INV_X1 U4127 ( .A(n3312), .ZN(n3314) );
  INV_X1 U4128 ( .A(n3747), .ZN(n3313) );
  OR2_X1 U4129 ( .A1(n3312), .A2(n3747), .ZN(n3373) );
  OAI21_X1 U4130 ( .B1(n3314), .B2(n3313), .A(n3373), .ZN(n3412) );
  INV_X1 U4131 ( .A(n3412), .ZN(n3324) );
  XOR2_X1 U4132 ( .A(n3747), .B(n3644), .Z(n3317) );
  OAI22_X1 U4133 ( .A1(n3408), .A2(n4140), .B1(n4139), .B2(n3318), .ZN(n3315)
         );
  AOI21_X1 U4134 ( .B1(n4148), .B2(n3806), .A(n3315), .ZN(n3316) );
  OAI21_X1 U4135 ( .B1(n3317), .B2(n4143), .A(n3316), .ZN(n3411) );
  INV_X1 U4136 ( .A(n3365), .ZN(n3319) );
  OAI21_X1 U4137 ( .B1(n3319), .B2(n3318), .A(n2044), .ZN(n3417) );
  NOR2_X1 U4138 ( .A1(n3417), .A2(n4107), .ZN(n3322) );
  OAI22_X1 U4139 ( .A1(n4375), .A2(n3320), .B1(n3466), .B2(n4153), .ZN(n3321)
         );
  AOI211_X1 U4140 ( .C1(n3411), .C2(n4375), .A(n3322), .B(n3321), .ZN(n3323)
         );
  OAI21_X1 U4141 ( .B1(n3324), .B2(n4137), .A(n3323), .ZN(U3276) );
  NAND2_X1 U4142 ( .A1(n3325), .A2(n4417), .ZN(n3327) );
  NAND2_X1 U4143 ( .A1(n3327), .A2(n3326), .ZN(n3330) );
  MUX2_X1 U4144 ( .A(REG0_REG_12__SCAN_IN), .B(n3330), .S(n4431), .Z(n3328) );
  INV_X1 U4145 ( .A(n3328), .ZN(n3329) );
  OAI21_X1 U4146 ( .B1(n3333), .B2(n4271), .A(n3329), .ZN(U3491) );
  MUX2_X1 U4147 ( .A(REG1_REG_12__SCAN_IN), .B(n3330), .S(n4443), .Z(n3331) );
  INV_X1 U4148 ( .A(n3331), .ZN(n3332) );
  OAI21_X1 U4149 ( .B1(n4223), .B2(n3333), .A(n3332), .ZN(U3530) );
  INV_X1 U4150 ( .A(n3335), .ZN(n3336) );
  AOI21_X1 U4151 ( .B1(n3751), .B2(n3334), .A(n3336), .ZN(n4426) );
  XOR2_X1 U4152 ( .A(n3751), .B(n3337), .Z(n3341) );
  OAI22_X1 U4153 ( .A1(n3361), .A2(n4140), .B1(n4139), .B2(n3344), .ZN(n3339)
         );
  NOR2_X1 U4154 ( .A1(n4426), .A2(n4080), .ZN(n3338) );
  AOI211_X1 U4155 ( .C1(n4148), .C2(n3808), .A(n3339), .B(n3338), .ZN(n3340)
         );
  OAI21_X1 U4156 ( .B1(n4143), .B2(n3341), .A(n3340), .ZN(n4428) );
  NAND2_X1 U4157 ( .A1(n4428), .A2(n4375), .ZN(n3350) );
  INV_X1 U4158 ( .A(n3342), .ZN(n3345) );
  OAI21_X1 U4159 ( .B1(n3345), .B2(n3344), .A(n3343), .ZN(n4423) );
  INV_X1 U4160 ( .A(n4423), .ZN(n3348) );
  OAI22_X1 U4161 ( .A1(n4375), .A2(n3346), .B1(n3392), .B2(n4153), .ZN(n3347)
         );
  AOI21_X1 U4162 ( .B1(n3348), .B2(n4362), .A(n3347), .ZN(n3349) );
  OAI211_X1 U4163 ( .C1(n4426), .C2(n4090), .A(n3350), .B(n3349), .ZN(U3279)
         );
  INV_X1 U4164 ( .A(n3351), .ZN(n3353) );
  OR2_X1 U4165 ( .A1(n3353), .A2(n3352), .ZN(n3768) );
  XOR2_X1 U4166 ( .A(n3768), .B(n3354), .Z(n3418) );
  INV_X1 U4167 ( .A(n3355), .ZN(n3356) );
  AOI21_X1 U4168 ( .B1(n3358), .B2(n3357), .A(n3356), .ZN(n3359) );
  XOR2_X1 U4169 ( .A(n3768), .B(n3359), .Z(n3363) );
  AOI22_X1 U4170 ( .A1(n3805), .A2(n4129), .B1(n4170), .B2(n3444), .ZN(n3360)
         );
  OAI21_X1 U4171 ( .B1(n3361), .B2(n4133), .A(n3360), .ZN(n3362) );
  AOI21_X1 U4172 ( .B1(n3363), .B2(n4126), .A(n3362), .ZN(n3364) );
  OAI21_X1 U4173 ( .B1(n3418), .B2(n4080), .A(n3364), .ZN(n3419) );
  NAND2_X1 U4174 ( .A1(n3419), .A2(n4375), .ZN(n3371) );
  OAI21_X1 U4175 ( .B1(n3367), .B2(n3366), .A(n3365), .ZN(n3426) );
  INV_X1 U4176 ( .A(n3426), .ZN(n3369) );
  OAI22_X1 U4177 ( .A1(n4375), .A2(n3850), .B1(n3447), .B2(n4153), .ZN(n3368)
         );
  AOI21_X1 U4178 ( .B1(n3369), .B2(n4362), .A(n3368), .ZN(n3370) );
  OAI211_X1 U4179 ( .C1(n3418), .C2(n4090), .A(n3371), .B(n3370), .ZN(U3277)
         );
  NAND2_X1 U4180 ( .A1(n3373), .A2(n3372), .ZN(n3374) );
  XNOR2_X1 U4181 ( .A(n3374), .B(n2013), .ZN(n4231) );
  XNOR2_X1 U4182 ( .A(n2044), .B(n3375), .ZN(n4229) );
  OAI22_X1 U4183 ( .A1(n4375), .A2(n3376), .B1(n3629), .B2(n4153), .ZN(n3377)
         );
  AOI21_X1 U4184 ( .B1(n4229), .B2(n4362), .A(n3377), .ZN(n3383) );
  OAI211_X1 U4185 ( .C1(n2047), .C2(n2013), .A(n4126), .B(n3378), .ZN(n3380)
         );
  AOI22_X1 U4186 ( .A1(n4147), .A2(n4129), .B1(n4170), .B2(n3624), .ZN(n3379)
         );
  OAI211_X1 U4187 ( .C1(n3381), .C2(n4133), .A(n3380), .B(n3379), .ZN(n4228)
         );
  NAND2_X1 U4188 ( .A1(n4228), .A2(n4375), .ZN(n3382) );
  OAI211_X1 U4189 ( .C1(n4231), .C2(n4137), .A(n3383), .B(n3382), .ZN(U3275)
         );
  XNOR2_X1 U4190 ( .A(n3386), .B(n3385), .ZN(n3387) );
  XNOR2_X1 U4191 ( .A(n3384), .B(n3387), .ZN(n3394) );
  NOR2_X1 U4192 ( .A1(STATE_REG_SCAN_IN), .A2(n3388), .ZN(n4305) );
  AOI21_X1 U4193 ( .B1(n3626), .B2(n3807), .A(n4305), .ZN(n3391) );
  AOI22_X1 U4194 ( .A1(n3623), .A2(n3808), .B1(n3625), .B2(n3389), .ZN(n3390)
         );
  OAI211_X1 U4195 ( .C1(n3630), .C2(n3392), .A(n3391), .B(n3390), .ZN(n3393)
         );
  AOI21_X1 U4196 ( .B1(n3394), .B2(n3632), .A(n3393), .ZN(n3395) );
  INV_X1 U4197 ( .A(n3395), .ZN(U3233) );
  OR2_X1 U4198 ( .A1(n3312), .A2(n3396), .ZN(n3398) );
  AND2_X1 U4199 ( .A1(n3398), .A2(n3397), .ZN(n3401) );
  OAI21_X1 U4200 ( .B1(n3401), .B2(n3400), .A(n3399), .ZN(n4227) );
  AOI21_X1 U4201 ( .B1(n3527), .B2(n2045), .A(n4150), .ZN(n4225) );
  OAI22_X1 U4202 ( .A1(n4375), .A2(n3402), .B1(n3530), .B2(n4153), .ZN(n3403)
         );
  AOI21_X1 U4203 ( .B1(n4225), .B2(n4362), .A(n3403), .ZN(n3410) );
  OAI211_X1 U4204 ( .C1(n3405), .C2(n3760), .A(n3404), .B(n4126), .ZN(n3407)
         );
  AOI22_X1 U4205 ( .A1(n3803), .A2(n4129), .B1(n4170), .B2(n3527), .ZN(n3406)
         );
  OAI211_X1 U4206 ( .C1(n3408), .C2(n4133), .A(n3407), .B(n3406), .ZN(n4224)
         );
  NAND2_X1 U4207 ( .A1(n4224), .A2(n4375), .ZN(n3409) );
  OAI211_X1 U4208 ( .C1(n4227), .C2(n4137), .A(n3410), .B(n3409), .ZN(U3274)
         );
  INV_X1 U4209 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3413) );
  AOI21_X1 U4210 ( .B1(n3412), .B2(n4417), .A(n3411), .ZN(n3415) );
  MUX2_X1 U4211 ( .A(n3413), .B(n3415), .S(n4431), .Z(n3414) );
  OAI21_X1 U4212 ( .B1(n3417), .B2(n4271), .A(n3414), .ZN(U3495) );
  INV_X1 U4213 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4501) );
  MUX2_X1 U4214 ( .A(n4501), .B(n3415), .S(n4443), .Z(n3416) );
  OAI21_X1 U4215 ( .B1(n4223), .B2(n3417), .A(n3416), .ZN(U3532) );
  INV_X1 U4216 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3421) );
  INV_X1 U4217 ( .A(n3418), .ZN(n3420) );
  AOI21_X1 U4218 ( .B1(n4402), .B2(n3420), .A(n3419), .ZN(n3423) );
  MUX2_X1 U4219 ( .A(n3421), .B(n3423), .S(n4443), .Z(n3422) );
  OAI21_X1 U4220 ( .B1(n4223), .B2(n3426), .A(n3422), .ZN(U3531) );
  INV_X1 U4221 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3424) );
  MUX2_X1 U4222 ( .A(n3424), .B(n3423), .S(n4431), .Z(n3425) );
  OAI21_X1 U4223 ( .B1(n3426), .B2(n4271), .A(n3425), .ZN(U3493) );
  INV_X1 U4224 ( .A(n3427), .ZN(n3429) );
  NAND2_X1 U4225 ( .A1(n3429), .A2(n3428), .ZN(n3430) );
  XNOR2_X1 U4226 ( .A(n3431), .B(n3430), .ZN(n3437) );
  AND2_X1 U4227 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4315) );
  AOI21_X1 U4228 ( .B1(n3623), .B2(n3484), .A(n4315), .ZN(n3434) );
  AOI22_X1 U4229 ( .A1(n3626), .A2(n3806), .B1(n3625), .B2(n3432), .ZN(n3433)
         );
  OAI211_X1 U4230 ( .C1(n3630), .C2(n3435), .A(n3434), .B(n3433), .ZN(n3436)
         );
  AOI21_X1 U4231 ( .B1(n3437), .B2(n3632), .A(n3436), .ZN(n3438) );
  INV_X1 U4232 ( .A(n3438), .ZN(U3221) );
  XNOR2_X1 U4233 ( .A(n3441), .B(n3440), .ZN(n3442) );
  XNOR2_X1 U4234 ( .A(n3439), .B(n3442), .ZN(n3449) );
  AOI21_X1 U4235 ( .B1(n3623), .B2(n3807), .A(n3443), .ZN(n3446) );
  AOI22_X1 U4236 ( .A1(n3626), .A2(n3805), .B1(n3625), .B2(n3444), .ZN(n3445)
         );
  OAI211_X1 U4237 ( .C1(n3630), .C2(n3447), .A(n3446), .B(n3445), .ZN(n3448)
         );
  AOI21_X1 U4238 ( .B1(n3449), .B2(n3632), .A(n3448), .ZN(n3450) );
  INV_X1 U4239 ( .A(n3450), .ZN(U3231) );
  XNOR2_X1 U4240 ( .A(n2027), .B(n3451), .ZN(n3456) );
  NOR2_X1 U4241 ( .A1(n3941), .A2(n3630), .ZN(n3454) );
  INV_X1 U4242 ( .A(n3625), .ZN(n3611) );
  AOI22_X1 U4243 ( .A1(n3979), .A2(n3623), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3452) );
  OAI21_X1 U4244 ( .B1(n3611), .B2(n3946), .A(n3452), .ZN(n3453) );
  AOI211_X1 U4245 ( .C1(n3626), .C2(n3949), .A(n3454), .B(n3453), .ZN(n3455)
         );
  OAI21_X1 U4246 ( .B1(n3456), .B2(n3617), .A(n3455), .ZN(U3211) );
  NAND2_X1 U4247 ( .A1(n3458), .A2(n3457), .ZN(n3461) );
  XOR2_X1 U4248 ( .A(n3461), .B(n3460), .Z(n3468) );
  NAND2_X1 U4249 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4331) );
  INV_X1 U4250 ( .A(n4331), .ZN(n3462) );
  AOI21_X1 U4251 ( .B1(n3623), .B2(n3806), .A(n3462), .ZN(n3465) );
  AOI22_X1 U4252 ( .A1(n3626), .A2(n3804), .B1(n3625), .B2(n3463), .ZN(n3464)
         );
  OAI211_X1 U4253 ( .C1(n3630), .C2(n3466), .A(n3465), .B(n3464), .ZN(n3467)
         );
  AOI21_X1 U4254 ( .B1(n3468), .B2(n3632), .A(n3467), .ZN(n3469) );
  INV_X1 U4255 ( .A(n3469), .ZN(U3212) );
  AND2_X1 U4256 ( .A1(n3470), .A2(n3471), .ZN(n3474) );
  OAI211_X1 U4257 ( .C1(n3474), .C2(n3473), .A(n3632), .B(n3472), .ZN(n3478)
         );
  NOR2_X1 U4258 ( .A1(n4015), .A2(n3610), .ZN(n3476) );
  OAI22_X1 U4259 ( .A1(n3982), .A2(n3612), .B1(n3611), .B2(n4014), .ZN(n3475)
         );
  AOI211_X1 U4260 ( .C1(REG3_REG_23__SCAN_IN), .C2(U3149), .A(n3476), .B(n3475), .ZN(n3477) );
  OAI211_X1 U4261 ( .C1(n3630), .C2(n4024), .A(n3478), .B(n3477), .ZN(U3213)
         );
  OAI211_X1 U4262 ( .C1(n3481), .C2(n3480), .A(n3479), .B(n3632), .ZN(n3489)
         );
  AND2_X1 U4263 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4296) );
  AOI21_X1 U4264 ( .B1(n3623), .B2(n3482), .A(n4296), .ZN(n3488) );
  AOI22_X1 U4265 ( .A1(n3626), .A2(n3484), .B1(n3625), .B2(n3483), .ZN(n3487)
         );
  OR2_X1 U4266 ( .A1(n3630), .A2(n3485), .ZN(n3486) );
  NAND4_X1 U4267 ( .A1(n3489), .A2(n3488), .A3(n3487), .A4(n3486), .ZN(U3214)
         );
  OR2_X1 U4268 ( .A1(n3492), .A2(n3490), .ZN(n3504) );
  OR2_X1 U4269 ( .A1(n3492), .A2(n3491), .ZN(n3494) );
  NAND2_X1 U4270 ( .A1(n3494), .A2(n3493), .ZN(n3495) );
  AOI21_X1 U4271 ( .B1(n3504), .B2(n3495), .A(n3617), .ZN(n3501) );
  NAND2_X1 U4272 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3899) );
  INV_X1 U4273 ( .A(n3899), .ZN(n3496) );
  AOI21_X1 U4274 ( .B1(n3626), .B2(n4101), .A(n3496), .ZN(n3499) );
  AOI22_X1 U4275 ( .A1(n3623), .A2(n3802), .B1(n3625), .B2(n3497), .ZN(n3498)
         );
  OAI211_X1 U4276 ( .C1(n3630), .C2(n4108), .A(n3499), .B(n3498), .ZN(n3500)
         );
  OR2_X1 U4277 ( .A1(n3501), .A2(n3500), .ZN(U3216) );
  NAND2_X1 U4278 ( .A1(n2043), .A2(n3502), .ZN(n3507) );
  NAND2_X1 U4279 ( .A1(n3504), .A2(n3503), .ZN(n3577) );
  INV_X1 U4280 ( .A(n3505), .ZN(n3579) );
  OAI211_X1 U4281 ( .C1(n3577), .C2(n3579), .A(n3575), .B(n3507), .ZN(n3506)
         );
  OAI211_X1 U4282 ( .C1(n3508), .C2(n3507), .A(n3632), .B(n3506), .ZN(n3512)
         );
  AOI22_X1 U4283 ( .A1(n4056), .A2(n3626), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3511) );
  AOI22_X1 U4284 ( .A1(n3623), .A2(n4101), .B1(n3625), .B2(n4059), .ZN(n3510)
         );
  OR2_X1 U4285 ( .A1(n3630), .A2(n4062), .ZN(n3509) );
  NAND4_X1 U4286 ( .A1(n3512), .A2(n3511), .A3(n3510), .A4(n3509), .ZN(U3220)
         );
  NOR2_X1 U4287 ( .A1(n2038), .A2(n3513), .ZN(n3514) );
  XNOR2_X1 U4288 ( .A(n3515), .B(n3514), .ZN(n3520) );
  INV_X1 U4289 ( .A(n3630), .ZN(n3615) );
  OAI22_X1 U4290 ( .A1(n3982), .A2(n3610), .B1(n3611), .B2(n3984), .ZN(n3518)
         );
  OAI22_X1 U4291 ( .A1(n3947), .A2(n3612), .B1(STATE_REG_SCAN_IN), .B2(n3516), 
        .ZN(n3517) );
  AOI211_X1 U4292 ( .C1(n3986), .C2(n3615), .A(n3518), .B(n3517), .ZN(n3519)
         );
  OAI21_X1 U4293 ( .B1(n3520), .B2(n3617), .A(n3519), .ZN(U3222) );
  INV_X1 U4294 ( .A(n3521), .ZN(n3524) );
  AND2_X1 U4295 ( .A1(n3523), .A2(n3522), .ZN(n3619) );
  OAI21_X1 U4296 ( .B1(n3524), .B2(n3620), .A(n3619), .ZN(n3526) );
  XNOR2_X1 U4297 ( .A(n3526), .B(n3525), .ZN(n3532) );
  AND2_X1 U4298 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n4334) );
  AOI21_X1 U4299 ( .B1(n3623), .B2(n3804), .A(n4334), .ZN(n3529) );
  AOI22_X1 U4300 ( .A1(n3626), .A2(n3803), .B1(n3625), .B2(n3527), .ZN(n3528)
         );
  OAI211_X1 U4301 ( .C1(n3630), .C2(n3530), .A(n3529), .B(n3528), .ZN(n3531)
         );
  AOI21_X1 U4302 ( .B1(n3532), .B2(n3632), .A(n3531), .ZN(n3533) );
  INV_X1 U4303 ( .A(n3533), .ZN(U3223) );
  OAI211_X1 U4304 ( .C1(n3536), .C2(n3535), .A(n3534), .B(n3632), .ZN(n3542)
         );
  AND2_X1 U4305 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3838) );
  AOI21_X1 U4306 ( .B1(n3626), .B2(n3811), .A(n3838), .ZN(n3541) );
  AOI22_X1 U4307 ( .A1(n3623), .A2(n3812), .B1(n3625), .B2(n3537), .ZN(n3540)
         );
  OR2_X1 U4308 ( .A1(n3630), .A2(n3538), .ZN(n3539) );
  NAND4_X1 U4309 ( .A1(n3542), .A2(n3541), .A3(n3540), .A4(n3539), .ZN(U3224)
         );
  NAND2_X1 U4310 ( .A1(n3544), .A2(n3543), .ZN(n3546) );
  XOR2_X1 U4311 ( .A(n3546), .B(n3545), .Z(n3551) );
  AND2_X1 U4312 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4344) );
  AOI21_X1 U4313 ( .B1(n3626), .B2(n3802), .A(n4344), .ZN(n3549) );
  AOI22_X1 U4314 ( .A1(n3623), .A2(n4147), .B1(n3625), .B2(n3547), .ZN(n3548)
         );
  OAI211_X1 U4315 ( .C1(n3630), .C2(n4154), .A(n3549), .B(n3548), .ZN(n3550)
         );
  AOI21_X1 U4316 ( .B1(n3551), .B2(n3632), .A(n3550), .ZN(n3552) );
  INV_X1 U4317 ( .A(n3552), .ZN(U3225) );
  NAND2_X1 U4318 ( .A1(n3554), .A2(n3553), .ZN(n3555) );
  XOR2_X1 U4319 ( .A(n3556), .B(n3555), .Z(n3561) );
  OAI22_X1 U4320 ( .A1(n2474), .A2(n3610), .B1(n3611), .B2(n4001), .ZN(n3559)
         );
  OAI22_X1 U4321 ( .A1(n3960), .A2(n3612), .B1(STATE_REG_SCAN_IN), .B2(n3557), 
        .ZN(n3558) );
  AOI211_X1 U4322 ( .C1(n4002), .C2(n3615), .A(n3559), .B(n3558), .ZN(n3560)
         );
  OAI21_X1 U4323 ( .B1(n3561), .B2(n3617), .A(n3560), .ZN(U3226) );
  OAI211_X1 U4324 ( .C1(n3564), .C2(n3563), .A(n3562), .B(n3632), .ZN(n3574)
         );
  INV_X1 U4325 ( .A(n3565), .ZN(n3566) );
  AOI21_X1 U4326 ( .B1(n3623), .B2(n3567), .A(n3566), .ZN(n3573) );
  AOI22_X1 U4327 ( .A1(n3626), .A2(n3569), .B1(n3625), .B2(n3568), .ZN(n3572)
         );
  OR2_X1 U4328 ( .A1(n3630), .A2(n3570), .ZN(n3571) );
  NAND4_X1 U4329 ( .A1(n3574), .A2(n3573), .A3(n3572), .A4(n3571), .ZN(U3227)
         );
  NAND2_X1 U4330 ( .A1(n3577), .A2(n3575), .ZN(n3580) );
  NOR2_X1 U4331 ( .A1(n3579), .A2(n3576), .ZN(n3578) );
  OAI22_X1 U4332 ( .A1(n3580), .A2(n3579), .B1(n3578), .B2(n3577), .ZN(n3585)
         );
  INV_X1 U4333 ( .A(n3581), .ZN(n4084) );
  AOI22_X1 U4334 ( .A1(n3626), .A2(n4037), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n3583) );
  AOI22_X1 U4335 ( .A1(n3623), .A2(n4130), .B1(n3625), .B2(n4081), .ZN(n3582)
         );
  OAI211_X1 U4336 ( .C1(n3630), .C2(n4084), .A(n3583), .B(n3582), .ZN(n3584)
         );
  AOI21_X1 U4337 ( .B1(n3585), .B2(n3632), .A(n3584), .ZN(n3586) );
  INV_X1 U4338 ( .A(n3586), .ZN(U3230) );
  INV_X1 U4339 ( .A(n3470), .ZN(n3587) );
  AOI21_X1 U4340 ( .B1(n3589), .B2(n3588), .A(n3587), .ZN(n3596) );
  INV_X1 U4341 ( .A(n4043), .ZN(n3594) );
  OAI22_X1 U4342 ( .A1(n4076), .A2(n3610), .B1(n3611), .B2(n3590), .ZN(n3593)
         );
  INV_X1 U4343 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3591) );
  OAI22_X1 U4344 ( .A1(n2474), .A2(n3612), .B1(STATE_REG_SCAN_IN), .B2(n3591), 
        .ZN(n3592) );
  AOI211_X1 U4345 ( .C1(n3594), .C2(n3615), .A(n3593), .B(n3592), .ZN(n3595)
         );
  OAI21_X1 U4346 ( .B1(n3596), .B2(n3617), .A(n3595), .ZN(U3232) );
  XOR2_X1 U4347 ( .A(n3599), .B(n3598), .Z(n3600) );
  XNOR2_X1 U4348 ( .A(n3597), .B(n3600), .ZN(n3604) );
  AND2_X1 U4349 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n3888) );
  AOI21_X1 U4350 ( .B1(n3626), .B2(n4130), .A(n3888), .ZN(n3602) );
  AOI22_X1 U4351 ( .A1(n3623), .A2(n3803), .B1(n3625), .B2(n4128), .ZN(n3601)
         );
  OAI211_X1 U4352 ( .C1(n3630), .C2(n4120), .A(n3602), .B(n3601), .ZN(n3603)
         );
  AOI21_X1 U4353 ( .B1(n3604), .B2(n3632), .A(n3603), .ZN(n3605) );
  INV_X1 U4354 ( .A(n3605), .ZN(U3235) );
  NAND2_X1 U4355 ( .A1(n2033), .A2(n3607), .ZN(n3608) );
  XNOR2_X1 U4356 ( .A(n3606), .B(n3608), .ZN(n3618) );
  INV_X1 U4357 ( .A(n3609), .ZN(n3967) );
  OAI22_X1 U4358 ( .A1(n3960), .A2(n3610), .B1(STATE_REG_SCAN_IN), .B2(n4539), 
        .ZN(n3614) );
  OAI22_X1 U4359 ( .A1(n3673), .A2(n3612), .B1(n3611), .B2(n3965), .ZN(n3613)
         );
  AOI211_X1 U4360 ( .C1(n3967), .C2(n3615), .A(n3614), .B(n3613), .ZN(n3616)
         );
  OAI21_X1 U4361 ( .B1(n3618), .B2(n3617), .A(n3616), .ZN(U3237) );
  NAND2_X1 U4362 ( .A1(n3521), .A2(n3619), .ZN(n3621) );
  XNOR2_X1 U4363 ( .A(n3621), .B(n3620), .ZN(n3633) );
  NOR2_X1 U4364 ( .A1(STATE_REG_SCAN_IN), .A2(n3622), .ZN(n3868) );
  AOI21_X1 U4365 ( .B1(n3623), .B2(n3805), .A(n3868), .ZN(n3628) );
  AOI22_X1 U4366 ( .A1(n3626), .A2(n4147), .B1(n3625), .B2(n3624), .ZN(n3627)
         );
  OAI211_X1 U4367 ( .C1(n3630), .C2(n3629), .A(n3628), .B(n3627), .ZN(n3631)
         );
  AOI21_X1 U4368 ( .B1(n3633), .B2(n3632), .A(n3631), .ZN(n3634) );
  INV_X1 U4369 ( .A(n3634), .ZN(U3238) );
  NAND2_X1 U4370 ( .A1(n2467), .A2(DATAI_30_), .ZN(n4163) );
  INV_X1 U4371 ( .A(REG2_REG_31__SCAN_IN), .ZN(n3637) );
  NAND2_X1 U4372 ( .A1(n2007), .A2(REG1_REG_31__SCAN_IN), .ZN(n3636) );
  NAND2_X1 U4373 ( .A1(n2280), .A2(REG0_REG_31__SCAN_IN), .ZN(n3635) );
  OAI211_X1 U4374 ( .C1(n2355), .C2(n3637), .A(n3636), .B(n3635), .ZN(n4165)
         );
  NAND2_X1 U4375 ( .A1(n3638), .A2(n3641), .ZN(n3707) );
  INV_X1 U4376 ( .A(n3639), .ZN(n3643) );
  INV_X1 U4377 ( .A(n3640), .ZN(n3642) );
  OAI21_X1 U4378 ( .B1(n3643), .B2(n3642), .A(n3641), .ZN(n3712) );
  OAI21_X1 U4379 ( .B1(n3644), .B2(n3707), .A(n3712), .ZN(n3646) );
  INV_X1 U4380 ( .A(n3713), .ZN(n3645) );
  AOI211_X1 U4381 ( .C1(n3646), .C2(n3716), .A(n3645), .B(n3715), .ZN(n3647)
         );
  OAI21_X1 U4382 ( .B1(n3647), .B2(n3719), .A(n3718), .ZN(n3649) );
  AOI21_X1 U4383 ( .B1(n3722), .B2(n3649), .A(n3648), .ZN(n3651) );
  OAI21_X1 U4384 ( .B1(n3651), .B2(n3724), .A(n3650), .ZN(n3652) );
  NAND4_X1 U4385 ( .A1(n3654), .A2(n3912), .A3(n3653), .A4(n3652), .ZN(n3667)
         );
  INV_X1 U4386 ( .A(n3740), .ZN(n3661) );
  NAND2_X1 U4387 ( .A1(n2467), .A2(DATAI_29_), .ZN(n3921) );
  INV_X1 U4388 ( .A(n3921), .ZN(n3915) );
  NAND2_X1 U4389 ( .A1(n2467), .A2(DATAI_31_), .ZN(n3734) );
  NAND2_X1 U4390 ( .A1(n4165), .A2(n3734), .ZN(n3737) );
  INV_X1 U4391 ( .A(REG2_REG_30__SCAN_IN), .ZN(n3657) );
  NAND2_X1 U4392 ( .A1(n2007), .A2(REG1_REG_30__SCAN_IN), .ZN(n3656) );
  NAND2_X1 U4393 ( .A1(n2280), .A2(REG0_REG_30__SCAN_IN), .ZN(n3655) );
  OAI211_X1 U4394 ( .C1(n2355), .C2(n3657), .A(n3656), .B(n3655), .ZN(n3916)
         );
  OR2_X1 U4395 ( .A1(n3916), .A2(n4163), .ZN(n3658) );
  NAND2_X1 U4396 ( .A1(n3737), .A2(n3658), .ZN(n3770) );
  AOI21_X1 U4397 ( .B1(n3661), .B2(n3915), .A(n3770), .ZN(n3662) );
  INV_X1 U4398 ( .A(n3662), .ZN(n3666) );
  INV_X1 U4399 ( .A(n3912), .ZN(n3660) );
  NOR2_X1 U4400 ( .A1(n3660), .A2(n3659), .ZN(n3663) );
  OAI21_X1 U4401 ( .B1(n3661), .B2(n3915), .A(n3911), .ZN(n3727) );
  OAI21_X1 U4402 ( .B1(n3663), .B2(n3727), .A(n3662), .ZN(n3731) );
  NOR3_X1 U4403 ( .A1(n3664), .A2(n3945), .A3(n3727), .ZN(n3665) );
  OAI22_X1 U4404 ( .A1(n3667), .A2(n3666), .B1(n3731), .B2(n3665), .ZN(n3668)
         );
  OAI21_X1 U4405 ( .B1(n4163), .B2(n4165), .A(n3668), .ZN(n3672) );
  AND2_X1 U4406 ( .A1(n3916), .A2(n4163), .ZN(n3733) );
  INV_X1 U4407 ( .A(n4165), .ZN(n3669) );
  INV_X1 U4408 ( .A(n3734), .ZN(n4166) );
  OAI21_X1 U4409 ( .B1(n3733), .B2(n3669), .A(n4166), .ZN(n3671) );
  AOI21_X1 U4410 ( .B1(n3672), .B2(n3671), .A(n3670), .ZN(n3794) );
  NOR2_X1 U4411 ( .A1(n3673), .A2(n3939), .ZN(n3730) );
  INV_X1 U4412 ( .A(n3674), .ZN(n3677) );
  OAI211_X1 U4413 ( .C1(n3677), .C2(n2530), .A(n3676), .B(n3675), .ZN(n3679)
         );
  NAND3_X1 U4414 ( .A1(n3679), .A2(n3678), .A3(n2533), .ZN(n3682) );
  NAND3_X1 U4415 ( .A1(n3682), .A2(n3681), .A3(n3680), .ZN(n3685) );
  NAND3_X1 U4416 ( .A1(n3685), .A2(n3684), .A3(n3683), .ZN(n3688) );
  NAND3_X1 U4417 ( .A1(n3688), .A2(n3687), .A3(n3686), .ZN(n3692) );
  INV_X1 U4418 ( .A(n3689), .ZN(n3690) );
  AOI21_X1 U4419 ( .B1(n3692), .B2(n3691), .A(n3690), .ZN(n3698) );
  NAND2_X1 U4420 ( .A1(n3694), .A2(n3693), .ZN(n3697) );
  OAI211_X1 U4421 ( .C1(n3698), .C2(n3697), .A(n3696), .B(n3695), .ZN(n3701)
         );
  NAND3_X1 U4422 ( .A1(n3701), .A2(n3700), .A3(n3699), .ZN(n3704) );
  AOI21_X1 U4423 ( .B1(n3704), .B2(n3703), .A(n2063), .ZN(n3711) );
  NAND2_X1 U4424 ( .A1(n3706), .A2(n3705), .ZN(n3710) );
  INV_X1 U4425 ( .A(n3707), .ZN(n3709) );
  OAI211_X1 U4426 ( .C1(n3711), .C2(n3710), .A(n3709), .B(n3708), .ZN(n3714)
         );
  NAND3_X1 U4427 ( .A1(n3714), .A2(n3713), .A3(n3712), .ZN(n3717) );
  AOI21_X1 U4428 ( .B1(n3717), .B2(n3716), .A(n3715), .ZN(n3720) );
  INV_X1 U4429 ( .A(n4008), .ZN(n3744) );
  OAI211_X1 U4430 ( .C1(n3720), .C2(n3719), .A(n3744), .B(n3718), .ZN(n3721)
         );
  NAND2_X1 U4431 ( .A1(n3722), .A2(n3721), .ZN(n3725) );
  AOI211_X1 U4432 ( .C1(n3726), .C2(n3725), .A(n3724), .B(n3723), .ZN(n3729)
         );
  NOR4_X1 U4433 ( .A1(n3730), .A2(n3729), .A3(n3728), .A4(n3727), .ZN(n3732)
         );
  OR2_X1 U4434 ( .A1(n3732), .A2(n3731), .ZN(n3739) );
  INV_X1 U4435 ( .A(n3733), .ZN(n3736) );
  OR2_X1 U4436 ( .A1(n4165), .A2(n3734), .ZN(n3735) );
  NAND2_X1 U4437 ( .A1(n3736), .A2(n3735), .ZN(n3769) );
  NAND2_X1 U4438 ( .A1(n3769), .A2(n3737), .ZN(n3738) );
  NAND2_X1 U4439 ( .A1(n3739), .A2(n3738), .ZN(n3792) );
  INV_X1 U4440 ( .A(n3905), .ZN(n3787) );
  NAND2_X1 U4441 ( .A1(n3742), .A2(n3741), .ZN(n3958) );
  NAND2_X1 U4442 ( .A1(n3743), .A2(n3955), .ZN(n3975) );
  NAND2_X1 U4443 ( .A1(n3744), .A2(n4009), .ZN(n4052) );
  INV_X1 U4444 ( .A(n4114), .ZN(n4124) );
  NAND4_X1 U4445 ( .A1(n4124), .A2(n3747), .A3(n3746), .A4(n3745), .ZN(n3754)
         );
  INV_X1 U4446 ( .A(n3748), .ZN(n3752) );
  NAND4_X1 U4447 ( .A1(n3752), .A2(n3751), .A3(n3750), .A4(n3749), .ZN(n3753)
         );
  OR2_X1 U4448 ( .A1(n3754), .A2(n3753), .ZN(n3763) );
  INV_X1 U4449 ( .A(n3755), .ZN(n3758) );
  INV_X1 U4450 ( .A(n4092), .ZN(n3756) );
  NAND4_X1 U4451 ( .A1(n3758), .A2(n4158), .A3(n2013), .A4(n3757), .ZN(n3762)
         );
  NAND2_X1 U4452 ( .A1(n3760), .A2(n3759), .ZN(n3761) );
  NOR4_X1 U4453 ( .A1(n4052), .A2(n3763), .A3(n3762), .A4(n3761), .ZN(n3782)
         );
  NAND2_X1 U4454 ( .A1(n3992), .A2(n3764), .ZN(n4012) );
  INV_X1 U4455 ( .A(n4012), .ZN(n3781) );
  XNOR2_X1 U4456 ( .A(n4101), .B(n3765), .ZN(n4068) );
  INV_X1 U4457 ( .A(n4068), .ZN(n4073) );
  NAND2_X1 U4458 ( .A1(n3767), .A2(n3766), .ZN(n4099) );
  NOR2_X1 U4459 ( .A1(n4099), .A2(n3768), .ZN(n3778) );
  NOR2_X1 U4460 ( .A1(n3770), .A2(n3769), .ZN(n3777) );
  NOR2_X1 U4461 ( .A1(n3772), .A2(n3771), .ZN(n3776) );
  NOR2_X1 U4462 ( .A1(n3774), .A2(n3773), .ZN(n3775) );
  NAND4_X1 U4463 ( .A1(n3778), .A2(n3777), .A3(n3776), .A4(n3775), .ZN(n3779)
         );
  NOR2_X1 U4464 ( .A1(n4031), .A2(n3779), .ZN(n3780) );
  NAND4_X1 U4465 ( .A1(n3782), .A2(n3781), .A3(n4073), .A4(n3780), .ZN(n3784)
         );
  NAND2_X1 U4466 ( .A1(n3783), .A2(n3973), .ZN(n3994) );
  NOR4_X1 U4467 ( .A1(n3958), .A2(n3975), .A3(n3784), .A4(n3994), .ZN(n3786)
         );
  INV_X1 U4468 ( .A(n3945), .ZN(n3785) );
  NAND4_X1 U4469 ( .A1(n3787), .A2(n2032), .A3(n3786), .A4(n3785), .ZN(n3789)
         );
  AND2_X1 U4470 ( .A1(n3789), .A2(n3788), .ZN(n3791) );
  MUX2_X1 U4471 ( .A(n3792), .B(n3791), .S(n3790), .Z(n3793) );
  NOR2_X1 U4472 ( .A1(n3794), .A2(n3793), .ZN(n3795) );
  XNOR2_X1 U4473 ( .A(n3795), .B(n4277), .ZN(n3801) );
  NAND2_X1 U4474 ( .A1(n3797), .A2(n3796), .ZN(n3798) );
  OAI211_X1 U4475 ( .C1(n4276), .C2(n3800), .A(n3798), .B(B_REG_SCAN_IN), .ZN(
        n3799) );
  OAI21_X1 U4476 ( .B1(n3801), .B2(n3800), .A(n3799), .ZN(U3239) );
  MUX2_X1 U4477 ( .A(DATAO_REG_31__SCAN_IN), .B(n4165), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4478 ( .A(DATAO_REG_30__SCAN_IN), .B(n3916), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4479 ( .A(DATAO_REG_28__SCAN_IN), .B(n3949), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4480 ( .A(DATAO_REG_25__SCAN_IN), .B(n3997), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4481 ( .A(DATAO_REG_24__SCAN_IN), .B(n4017), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U4482 ( .A(DATAO_REG_23__SCAN_IN), .B(n4036), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U4483 ( .A(DATAO_REG_22__SCAN_IN), .B(n4056), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4484 ( .A(DATAO_REG_21__SCAN_IN), .B(n4037), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U4485 ( .A(DATAO_REG_18__SCAN_IN), .B(n3802), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4486 ( .A(DATAO_REG_17__SCAN_IN), .B(n3803), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4487 ( .A(DATAO_REG_15__SCAN_IN), .B(n3804), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U4488 ( .A(DATAO_REG_14__SCAN_IN), .B(n3805), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4489 ( .A(DATAO_REG_13__SCAN_IN), .B(n3806), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4490 ( .A(DATAO_REG_12__SCAN_IN), .B(n3807), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4491 ( .A(DATAO_REG_10__SCAN_IN), .B(n3808), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U4492 ( .A(DATAO_REG_8__SCAN_IN), .B(n3809), .S(U4043), .Z(U3558) );
  MUX2_X1 U4493 ( .A(DATAO_REG_7__SCAN_IN), .B(n3810), .S(U4043), .Z(U3557) );
  MUX2_X1 U4494 ( .A(DATAO_REG_6__SCAN_IN), .B(n3811), .S(U4043), .Z(U3556) );
  MUX2_X1 U4495 ( .A(DATAO_REG_4__SCAN_IN), .B(n3812), .S(U4043), .Z(U3554) );
  MUX2_X1 U4496 ( .A(DATAO_REG_2__SCAN_IN), .B(n2254), .S(U4043), .Z(U3552) );
  MUX2_X1 U4497 ( .A(DATAO_REG_1__SCAN_IN), .B(n3813), .S(U4043), .Z(U3551) );
  MUX2_X1 U4498 ( .A(DATAO_REG_0__SCAN_IN), .B(n3814), .S(U4043), .Z(U3550) );
  OAI211_X1 U4499 ( .C1(n3816), .C2(n3815), .A(n4355), .B(n3830), .ZN(n3824)
         );
  OAI211_X1 U4500 ( .C1(n3819), .C2(n3818), .A(n4353), .B(n3817), .ZN(n3823)
         );
  AOI22_X1 U4501 ( .A1(n4345), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3822) );
  NAND2_X1 U4502 ( .A1(n4330), .A2(n3820), .ZN(n3821) );
  NAND4_X1 U4503 ( .A1(n3824), .A2(n3823), .A3(n3822), .A4(n3821), .ZN(U3241)
         );
  AOI22_X1 U4504 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4345), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3835) );
  XOR2_X1 U4505 ( .A(n3826), .B(n3825), .Z(n3827) );
  AOI22_X1 U4506 ( .A1(n4286), .A2(n4330), .B1(n4353), .B2(n3827), .ZN(n3834)
         );
  MUX2_X1 U4507 ( .A(n2888), .B(REG2_REG_2__SCAN_IN), .S(n4286), .Z(n3828) );
  NAND3_X1 U4508 ( .A1(n3830), .A2(n3829), .A3(n3828), .ZN(n3831) );
  NAND3_X1 U4509 ( .A1(n4355), .A2(n3832), .A3(n3831), .ZN(n3833) );
  NAND4_X1 U4510 ( .A1(n3836), .A2(n3835), .A3(n3834), .A4(n3833), .ZN(U3242)
         );
  NOR2_X1 U4511 ( .A1(n4358), .A2(n4282), .ZN(n3837) );
  AOI211_X1 U4512 ( .C1(n4345), .C2(ADDR_REG_5__SCAN_IN), .A(n3838), .B(n3837), 
        .ZN(n3847) );
  OAI211_X1 U4513 ( .C1(n3841), .C2(n3840), .A(n4353), .B(n3839), .ZN(n3846)
         );
  OAI211_X1 U4514 ( .C1(n3844), .C2(n3843), .A(n4355), .B(n3842), .ZN(n3845)
         );
  NAND3_X1 U4515 ( .A1(n3847), .A2(n3846), .A3(n3845), .ZN(U3245) );
  INV_X1 U4516 ( .A(n4278), .ZN(n3871) );
  NAND2_X1 U4517 ( .A1(n3871), .A2(REG2_REG_15__SCAN_IN), .ZN(n3849) );
  NAND2_X1 U4518 ( .A1(n4278), .A2(n3376), .ZN(n3848) );
  AND2_X1 U4519 ( .A1(n3849), .A2(n3848), .ZN(n3859) );
  INV_X1 U4520 ( .A(n4329), .ZN(n4385) );
  INV_X1 U4521 ( .A(n3852), .ZN(n3851) );
  NOR2_X1 U4522 ( .A1(n3851), .A2(n3850), .ZN(n3854) );
  OAI22_X1 U4523 ( .A1(n3854), .A2(n3853), .B1(REG2_REG_13__SCAN_IN), .B2(
        n3852), .ZN(n3855) );
  NOR2_X1 U4524 ( .A1(n4385), .A2(n3855), .ZN(n3856) );
  XOR2_X1 U4525 ( .A(n4329), .B(n3855), .Z(n4326) );
  NOR2_X1 U4526 ( .A1(n3320), .A2(n4326), .ZN(n4325) );
  INV_X1 U4527 ( .A(n3874), .ZN(n3857) );
  AOI21_X1 U4528 ( .B1(n3859), .B2(n3858), .A(n3857), .ZN(n3860) );
  NAND2_X1 U4529 ( .A1(n4355), .A2(n3860), .ZN(n3870) );
  NAND2_X1 U4530 ( .A1(n4278), .A2(REG1_REG_15__SCAN_IN), .ZN(n3880) );
  OAI21_X1 U4531 ( .B1(n4278), .B2(REG1_REG_15__SCAN_IN), .A(n3880), .ZN(n3865) );
  INV_X1 U4532 ( .A(n3881), .ZN(n3864) );
  AOI211_X1 U4533 ( .C1(n3866), .C2(n3865), .A(n3864), .B(n4321), .ZN(n3867)
         );
  AOI211_X1 U4534 ( .C1(n4345), .C2(ADDR_REG_15__SCAN_IN), .A(n3868), .B(n3867), .ZN(n3869) );
  OAI211_X1 U4535 ( .C1(n3871), .C2(n4358), .A(n3870), .B(n3869), .ZN(U3255)
         );
  INV_X1 U4536 ( .A(n3895), .ZN(n3890) );
  XNOR2_X1 U4537 ( .A(n3895), .B(REG2_REG_18__SCAN_IN), .ZN(n3878) );
  NOR2_X1 U4538 ( .A1(n3885), .A2(REG2_REG_17__SCAN_IN), .ZN(n3872) );
  AOI21_X1 U4539 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3885), .A(n3872), .ZN(n4348) );
  NAND2_X1 U4540 ( .A1(n4278), .A2(REG2_REG_15__SCAN_IN), .ZN(n3873) );
  NAND2_X1 U4541 ( .A1(n3875), .A2(n4384), .ZN(n3876) );
  NAND2_X1 U4542 ( .A1(n4336), .A2(n3402), .ZN(n4335) );
  AOI21_X1 U4543 ( .B1(n3878), .B2(n3877), .A(n3894), .ZN(n3879) );
  NAND2_X1 U4544 ( .A1(n4355), .A2(n3879), .ZN(n3889) );
  XNOR2_X1 U4545 ( .A(n3895), .B(REG1_REG_18__SCAN_IN), .ZN(n3887) );
  INV_X1 U4546 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4551) );
  AOI22_X1 U4547 ( .A1(n3885), .A2(REG1_REG_17__SCAN_IN), .B1(n4551), .B2(
        n4382), .ZN(n4351) );
  NAND2_X1 U4548 ( .A1(n3883), .A2(n4384), .ZN(n3884) );
  INV_X1 U4549 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4338) );
  NAND2_X1 U4550 ( .A1(n4339), .A2(n4338), .ZN(n4337) );
  NAND2_X1 U4551 ( .A1(n3884), .A2(n4337), .ZN(n4350) );
  NAND2_X1 U4552 ( .A1(n4351), .A2(n4350), .ZN(n4349) );
  OAI21_X1 U4553 ( .B1(n3885), .B2(REG1_REG_17__SCAN_IN), .A(n4349), .ZN(n3886) );
  AOI21_X1 U4554 ( .B1(n3895), .B2(REG1_REG_18__SCAN_IN), .A(n3891), .ZN(n3893) );
  XNOR2_X1 U4555 ( .A(n4277), .B(REG1_REG_19__SCAN_IN), .ZN(n3892) );
  XNOR2_X1 U4556 ( .A(n3893), .B(n3892), .ZN(n3904) );
  AOI21_X1 U4557 ( .B1(n3895), .B2(REG2_REG_18__SCAN_IN), .A(n3894), .ZN(n3897) );
  MUX2_X1 U4558 ( .A(REG2_REG_19__SCAN_IN), .B(n4109), .S(n4277), .Z(n3896) );
  XNOR2_X1 U4559 ( .A(n3897), .B(n3896), .ZN(n3902) );
  NAND2_X1 U4560 ( .A1(n4345), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3898) );
  OAI211_X1 U4561 ( .C1(n4358), .C2(n3900), .A(n3899), .B(n3898), .ZN(n3901)
         );
  AOI21_X1 U4562 ( .B1(n3902), .B2(n4355), .A(n3901), .ZN(n3903) );
  OAI21_X1 U4563 ( .B1(n3904), .B2(n4321), .A(n3903), .ZN(U3259) );
  NAND2_X1 U4564 ( .A1(n3906), .A2(n3905), .ZN(n3909) );
  NAND2_X1 U4565 ( .A1(n3909), .A2(n3908), .ZN(n3910) );
  XNOR2_X1 U4566 ( .A(n3910), .B(n2032), .ZN(n4173) );
  INV_X1 U4567 ( .A(n4173), .ZN(n3927) );
  INV_X1 U4568 ( .A(n3911), .ZN(n3913) );
  AOI21_X1 U4569 ( .B1(B_REG_SCAN_IN), .B2(n4275), .A(n4140), .ZN(n4164) );
  AOI22_X1 U4570 ( .A1(n3916), .A2(n4164), .B1(n4170), .B2(n3915), .ZN(n3917)
         );
  OAI21_X1 U4571 ( .B1(n3918), .B2(n4133), .A(n3917), .ZN(n3919) );
  OAI21_X1 U4572 ( .B1(n3920), .B2(n4153), .A(n4175), .ZN(n3925) );
  OAI22_X1 U4573 ( .A1(n4174), .A2(n4107), .B1(n3923), .B2(n4375), .ZN(n3924)
         );
  AOI21_X1 U4574 ( .B1(n3925), .B2(n4375), .A(n3924), .ZN(n3926) );
  OAI21_X1 U4575 ( .B1(n3927), .B2(n4137), .A(n3926), .ZN(U3354) );
  INV_X1 U4576 ( .A(n3928), .ZN(n3934) );
  OAI22_X1 U4577 ( .A1(n3930), .A2(n4153), .B1(n3929), .B2(n4375), .ZN(n3933)
         );
  NOR2_X1 U4578 ( .A1(n3931), .A2(n4377), .ZN(n3932) );
  AOI211_X1 U4579 ( .C1(n4362), .C2(n3934), .A(n3933), .B(n3932), .ZN(n3935)
         );
  OAI21_X1 U4580 ( .B1(n3936), .B2(n4137), .A(n3935), .ZN(U3262) );
  XOR2_X1 U4581 ( .A(n3945), .B(n3937), .Z(n4181) );
  AOI21_X1 U4582 ( .B1(n3939), .B2(n2031), .A(n3938), .ZN(n4179) );
  OAI22_X1 U4583 ( .A1(n3941), .A2(n4153), .B1(n3940), .B2(n4375), .ZN(n3942)
         );
  AOI21_X1 U4584 ( .B1(n4179), .B2(n4362), .A(n3942), .ZN(n3953) );
  AOI21_X1 U4585 ( .B1(n3945), .B2(n3944), .A(n3943), .ZN(n3951) );
  OAI22_X1 U4586 ( .A1(n3947), .A2(n4133), .B1(n3946), .B2(n4139), .ZN(n3948)
         );
  AOI21_X1 U4587 ( .B1(n3949), .B2(n4129), .A(n3948), .ZN(n3950) );
  OAI21_X1 U4588 ( .B1(n3951), .B2(n4143), .A(n3950), .ZN(n4178) );
  NAND2_X1 U4589 ( .A1(n4178), .A2(n4375), .ZN(n3952) );
  OAI211_X1 U4590 ( .C1(n4181), .C2(n4137), .A(n3953), .B(n3952), .ZN(U3263)
         );
  XOR2_X1 U4591 ( .A(n3958), .B(n3954), .Z(n4183) );
  INV_X1 U4592 ( .A(n4183), .ZN(n3971) );
  INV_X1 U4593 ( .A(n3974), .ZN(n3957) );
  OAI21_X1 U4594 ( .B1(n3957), .B2(n3956), .A(n3955), .ZN(n3959) );
  XNOR2_X1 U4595 ( .A(n3959), .B(n3958), .ZN(n3964) );
  OAI22_X1 U4596 ( .A1(n3960), .A2(n4133), .B1(n3965), .B2(n4139), .ZN(n3961)
         );
  AOI21_X1 U4597 ( .B1(n3962), .B2(n4129), .A(n3961), .ZN(n3963) );
  OAI21_X1 U4598 ( .B1(n3964), .B2(n4143), .A(n3963), .ZN(n4182) );
  INV_X1 U4599 ( .A(n3983), .ZN(n3966) );
  OAI21_X1 U4600 ( .B1(n3966), .B2(n3965), .A(n2031), .ZN(n4242) );
  AOI22_X1 U4601 ( .A1(n3967), .A2(n4371), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4377), .ZN(n3968) );
  OAI21_X1 U4602 ( .B1(n4242), .B2(n4107), .A(n3968), .ZN(n3969) );
  AOI21_X1 U4603 ( .B1(n4182), .B2(n4375), .A(n3969), .ZN(n3970) );
  OAI21_X1 U4604 ( .B1(n3971), .B2(n4137), .A(n3970), .ZN(U3264) );
  XNOR2_X1 U4605 ( .A(n3972), .B(n3975), .ZN(n4187) );
  INV_X1 U4606 ( .A(n4187), .ZN(n3990) );
  NAND2_X1 U4607 ( .A1(n3974), .A2(n3973), .ZN(n3976) );
  XNOR2_X1 U4608 ( .A(n3976), .B(n3975), .ZN(n3977) );
  NAND2_X1 U4609 ( .A1(n3977), .A2(n4126), .ZN(n3981) );
  AOI22_X1 U4610 ( .A1(n3979), .A2(n4129), .B1(n4170), .B2(n3978), .ZN(n3980)
         );
  OAI211_X1 U4611 ( .C1(n3982), .C2(n4133), .A(n3981), .B(n3980), .ZN(n4186)
         );
  INV_X1 U4612 ( .A(n4000), .ZN(n3985) );
  OAI21_X1 U4613 ( .B1(n3985), .B2(n3984), .A(n3983), .ZN(n4246) );
  AOI22_X1 U4614 ( .A1(n3986), .A2(n4371), .B1(n4377), .B2(
        REG2_REG_25__SCAN_IN), .ZN(n3987) );
  OAI21_X1 U4615 ( .B1(n4246), .B2(n4107), .A(n3987), .ZN(n3988) );
  AOI21_X1 U4616 ( .B1(n4186), .B2(n4375), .A(n3988), .ZN(n3989) );
  OAI21_X1 U4617 ( .B1(n3990), .B2(n4137), .A(n3989), .ZN(U3265) );
  XOR2_X1 U4618 ( .A(n3994), .B(n3991), .Z(n4191) );
  INV_X1 U4619 ( .A(n4191), .ZN(n4006) );
  NAND2_X1 U4620 ( .A1(n3993), .A2(n3992), .ZN(n3995) );
  XNOR2_X1 U4621 ( .A(n3995), .B(n3994), .ZN(n3999) );
  OAI22_X1 U4622 ( .A1(n2474), .A2(n4133), .B1(n4139), .B2(n4001), .ZN(n3996)
         );
  AOI21_X1 U4623 ( .B1(n4129), .B2(n3997), .A(n3996), .ZN(n3998) );
  OAI21_X1 U4624 ( .B1(n3999), .B2(n4143), .A(n3998), .ZN(n4190) );
  OAI21_X1 U4625 ( .B1(n4020), .B2(n4001), .A(n4000), .ZN(n4249) );
  AOI22_X1 U4626 ( .A1(n4002), .A2(n4371), .B1(n4377), .B2(
        REG2_REG_24__SCAN_IN), .ZN(n4003) );
  OAI21_X1 U4627 ( .B1(n4249), .B2(n4107), .A(n4003), .ZN(n4004) );
  AOI21_X1 U4628 ( .B1(n4190), .B2(n4375), .A(n4004), .ZN(n4005) );
  OAI21_X1 U4629 ( .B1(n4006), .B2(n4137), .A(n4005), .ZN(U3266) );
  XOR2_X1 U4630 ( .A(n4012), .B(n4007), .Z(n4195) );
  INV_X1 U4631 ( .A(n4195), .ZN(n4029) );
  OR2_X1 U4632 ( .A1(n4051), .A2(n4008), .ZN(n4010) );
  NAND2_X1 U4633 ( .A1(n4010), .A2(n4009), .ZN(n4034) );
  INV_X1 U4634 ( .A(n4031), .ZN(n4035) );
  NAND2_X1 U4635 ( .A1(n4034), .A2(n4035), .ZN(n4033) );
  NAND2_X1 U4636 ( .A1(n4033), .A2(n4011), .ZN(n4013) );
  XNOR2_X1 U4637 ( .A(n4013), .B(n4012), .ZN(n4019) );
  OAI22_X1 U4638 ( .A1(n4015), .A2(n4133), .B1(n4139), .B2(n4014), .ZN(n4016)
         );
  AOI21_X1 U4639 ( .B1(n4129), .B2(n4017), .A(n4016), .ZN(n4018) );
  OAI21_X1 U4640 ( .B1(n4019), .B2(n4143), .A(n4018), .ZN(n4194) );
  INV_X1 U4641 ( .A(n4020), .ZN(n4023) );
  NAND2_X1 U4642 ( .A1(n4199), .A2(n4021), .ZN(n4022) );
  NAND2_X1 U4643 ( .A1(n4023), .A2(n4022), .ZN(n4253) );
  NOR2_X1 U4644 ( .A1(n4253), .A2(n4107), .ZN(n4027) );
  OAI22_X1 U4645 ( .A1(n4025), .A2(n4375), .B1(n4024), .B2(n4153), .ZN(n4026)
         );
  AOI211_X1 U4646 ( .C1(n4194), .C2(n4375), .A(n4027), .B(n4026), .ZN(n4028)
         );
  OAI21_X1 U4647 ( .B1(n4029), .B2(n4137), .A(n4028), .ZN(U3267) );
  OAI21_X1 U4648 ( .B1(n4032), .B2(n4031), .A(n4030), .ZN(n4202) );
  OAI21_X1 U4649 ( .B1(n4035), .B2(n4034), .A(n4033), .ZN(n4041) );
  NAND2_X1 U4650 ( .A1(n4036), .A2(n4129), .ZN(n4039) );
  AOI22_X1 U4651 ( .A1(n4037), .A2(n4148), .B1(n4042), .B2(n4170), .ZN(n4038)
         );
  NAND2_X1 U4652 ( .A1(n4039), .A2(n4038), .ZN(n4040) );
  AOI21_X1 U4653 ( .B1(n4041), .B2(n4126), .A(n4040), .ZN(n4201) );
  INV_X1 U4654 ( .A(n4201), .ZN(n4047) );
  NAND2_X1 U4655 ( .A1(n4061), .A2(n4042), .ZN(n4198) );
  AND3_X1 U4656 ( .A1(n4199), .A2(n4362), .A3(n4198), .ZN(n4046) );
  OAI22_X1 U4657 ( .A1(n4375), .A2(n4044), .B1(n4043), .B2(n4153), .ZN(n4045)
         );
  AOI211_X1 U4658 ( .C1(n4047), .C2(n4375), .A(n4046), .B(n4045), .ZN(n4048)
         );
  OAI21_X1 U4659 ( .B1(n4202), .B2(n4137), .A(n4048), .ZN(U3268) );
  XOR2_X1 U4660 ( .A(n4052), .B(n4050), .Z(n4204) );
  INV_X1 U4661 ( .A(n4204), .ZN(n4067) );
  XOR2_X1 U4662 ( .A(n4052), .B(n4051), .Z(n4058) );
  OAI22_X1 U4663 ( .A1(n4054), .A2(n4133), .B1(n4053), .B2(n4139), .ZN(n4055)
         );
  AOI21_X1 U4664 ( .B1(n4129), .B2(n4056), .A(n4055), .ZN(n4057) );
  OAI21_X1 U4665 ( .B1(n4058), .B2(n4143), .A(n4057), .ZN(n4203) );
  NAND2_X1 U4666 ( .A1(n4083), .A2(n4059), .ZN(n4060) );
  NAND2_X1 U4667 ( .A1(n4061), .A2(n4060), .ZN(n4258) );
  NOR2_X1 U4668 ( .A1(n4258), .A2(n4107), .ZN(n4065) );
  OAI22_X1 U4669 ( .A1(n4375), .A2(n4063), .B1(n4062), .B2(n4153), .ZN(n4064)
         );
  AOI211_X1 U4670 ( .C1(n4203), .C2(n4375), .A(n4065), .B(n4064), .ZN(n4066)
         );
  OAI21_X1 U4671 ( .B1(n4067), .B2(n4137), .A(n4066), .ZN(U3269) );
  XNOR2_X1 U4672 ( .A(n4069), .B(n4068), .ZN(n4206) );
  INV_X1 U4673 ( .A(n4070), .ZN(n4071) );
  NAND2_X1 U4674 ( .A1(n4072), .A2(n4071), .ZN(n4074) );
  XNOR2_X1 U4675 ( .A(n4074), .B(n4073), .ZN(n4078) );
  AOI22_X1 U4676 ( .A1(n4130), .A2(n4148), .B1(n4081), .B2(n4170), .ZN(n4075)
         );
  OAI21_X1 U4677 ( .B1(n4076), .B2(n4140), .A(n4075), .ZN(n4077) );
  AOI21_X1 U4678 ( .B1(n4078), .B2(n4126), .A(n4077), .ZN(n4079) );
  OAI21_X1 U4679 ( .B1(n4206), .B2(n4080), .A(n4079), .ZN(n4207) );
  NAND2_X1 U4680 ( .A1(n4207), .A2(n4375), .ZN(n4089) );
  NAND2_X1 U4681 ( .A1(n4104), .A2(n4081), .ZN(n4082) );
  NAND2_X1 U4682 ( .A1(n4083), .A2(n4082), .ZN(n4262) );
  INV_X1 U4683 ( .A(n4262), .ZN(n4087) );
  OAI22_X1 U4684 ( .A1(n4375), .A2(n4085), .B1(n4084), .B2(n4153), .ZN(n4086)
         );
  AOI21_X1 U4685 ( .B1(n4087), .B2(n4362), .A(n4086), .ZN(n4088) );
  OAI211_X1 U4686 ( .C1(n4206), .C2(n4090), .A(n4089), .B(n4088), .ZN(U3270)
         );
  XOR2_X1 U4687 ( .A(n4099), .B(n4091), .Z(n4211) );
  INV_X1 U4688 ( .A(n4211), .ZN(n4113) );
  OR2_X1 U4689 ( .A1(n4142), .A2(n4092), .ZN(n4094) );
  NAND2_X1 U4690 ( .A1(n4094), .A2(n4093), .ZN(n4125) );
  INV_X1 U4691 ( .A(n4095), .ZN(n4097) );
  OAI21_X1 U4692 ( .B1(n4125), .B2(n4097), .A(n4096), .ZN(n4098) );
  XOR2_X1 U4693 ( .A(n4099), .B(n4098), .Z(n4103) );
  OAI22_X1 U4694 ( .A1(n4141), .A2(n4133), .B1(n4105), .B2(n4139), .ZN(n4100)
         );
  AOI21_X1 U4695 ( .B1(n4101), .B2(n4129), .A(n4100), .ZN(n4102) );
  OAI21_X1 U4696 ( .B1(n4103), .B2(n4143), .A(n4102), .ZN(n4210) );
  OAI21_X1 U4697 ( .B1(n4106), .B2(n4105), .A(n4104), .ZN(n4266) );
  NOR2_X1 U4698 ( .A1(n4266), .A2(n4107), .ZN(n4111) );
  OAI22_X1 U4699 ( .A1(n4375), .A2(n4109), .B1(n4108), .B2(n4153), .ZN(n4110)
         );
  AOI211_X1 U4700 ( .C1(n4210), .C2(n4375), .A(n4111), .B(n4110), .ZN(n4112)
         );
  OAI21_X1 U4701 ( .B1(n4113), .B2(n4137), .A(n4112), .ZN(U3271) );
  NOR2_X1 U4702 ( .A1(n4115), .A2(n4114), .ZN(n4116) );
  OR2_X1 U4703 ( .A1(n4117), .A2(n4116), .ZN(n4214) );
  INV_X1 U4704 ( .A(n4214), .ZN(n4138) );
  XNOR2_X1 U4705 ( .A(n4152), .B(n4118), .ZN(n4119) );
  AND2_X1 U4706 ( .A1(n4119), .A2(n2619), .ZN(n4215) );
  OAI22_X1 U4707 ( .A1(n4375), .A2(n4121), .B1(n4120), .B2(n4153), .ZN(n4122)
         );
  AOI21_X1 U4708 ( .B1(n4215), .B2(n4123), .A(n4122), .ZN(n4136) );
  XNOR2_X1 U4709 ( .A(n4125), .B(n4124), .ZN(n4127) );
  NAND2_X1 U4710 ( .A1(n4127), .A2(n4126), .ZN(n4132) );
  AOI22_X1 U4711 ( .A1(n4130), .A2(n4129), .B1(n4170), .B2(n4128), .ZN(n4131)
         );
  OAI211_X1 U4712 ( .C1(n4134), .C2(n4133), .A(n4132), .B(n4131), .ZN(n4216)
         );
  NAND2_X1 U4713 ( .A1(n4216), .A2(n4375), .ZN(n4135) );
  OAI211_X1 U4714 ( .C1(n4138), .C2(n4137), .A(n4136), .B(n4135), .ZN(U3272)
         );
  OAI22_X1 U4715 ( .A1(n4141), .A2(n4140), .B1(n4149), .B2(n4139), .ZN(n4146)
         );
  XNOR2_X1 U4716 ( .A(n4142), .B(n4158), .ZN(n4144) );
  NOR2_X1 U4717 ( .A1(n4144), .A2(n4143), .ZN(n4145) );
  AOI211_X1 U4718 ( .C1(n4148), .C2(n4147), .A(n4146), .B(n4145), .ZN(n4219)
         );
  OR2_X1 U4719 ( .A1(n4150), .A2(n4149), .ZN(n4151) );
  NAND2_X1 U4720 ( .A1(n4152), .A2(n4151), .ZN(n4272) );
  INV_X1 U4721 ( .A(n4272), .ZN(n4157) );
  OAI22_X1 U4722 ( .A1(n4375), .A2(n4550), .B1(n4154), .B2(n4153), .ZN(n4156)
         );
  AOI21_X1 U4723 ( .B1(n4157), .B2(n4362), .A(n4156), .ZN(n4162) );
  XNOR2_X1 U4724 ( .A(n4159), .B(n4158), .ZN(n4221) );
  NAND2_X1 U4725 ( .A1(n4221), .A2(n4160), .ZN(n4161) );
  OAI211_X1 U4726 ( .C1(n4219), .C2(n4377), .A(n4162), .B(n4161), .ZN(U3273)
         );
  INV_X1 U4727 ( .A(n4163), .ZN(n4171) );
  XNOR2_X1 U4728 ( .A(n4168), .B(n4166), .ZN(n4288) );
  INV_X1 U4729 ( .A(n4288), .ZN(n4234) );
  INV_X1 U4730 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4507) );
  AND2_X1 U4731 ( .A1(n4165), .A2(n4164), .ZN(n4169) );
  AOI21_X1 U4732 ( .B1(n4166), .B2(n4170), .A(n4169), .ZN(n4290) );
  MUX2_X1 U4733 ( .A(n4507), .B(n4290), .S(n4443), .Z(n4167) );
  OAI21_X1 U4734 ( .B1(n4234), .B2(n4223), .A(n4167), .ZN(U3549) );
  AOI21_X1 U4735 ( .B1(n4171), .B2(n2030), .A(n4168), .ZN(n4291) );
  INV_X1 U4736 ( .A(n4291), .ZN(n4236) );
  INV_X1 U4737 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4505) );
  AOI21_X1 U4738 ( .B1(n4171), .B2(n4170), .A(n4169), .ZN(n4293) );
  MUX2_X1 U4739 ( .A(n4505), .B(n4293), .S(n4443), .Z(n4172) );
  OAI21_X1 U4740 ( .B1(n4236), .B2(n4223), .A(n4172), .ZN(U3548) );
  NAND2_X1 U4741 ( .A1(n4173), .A2(n4417), .ZN(n4177) );
  NAND2_X1 U4742 ( .A1(n4177), .A2(n2200), .ZN(n4237) );
  MUX2_X1 U4743 ( .A(REG1_REG_29__SCAN_IN), .B(n4237), .S(n4443), .Z(U3547) );
  AOI21_X1 U4744 ( .B1(n2619), .B2(n4179), .A(n4178), .ZN(n4180) );
  OAI21_X1 U4745 ( .B1(n4181), .B2(n4411), .A(n4180), .ZN(n4238) );
  MUX2_X1 U4746 ( .A(REG1_REG_27__SCAN_IN), .B(n4238), .S(n4443), .Z(U3545) );
  INV_X1 U4747 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4184) );
  AOI21_X1 U4748 ( .B1(n4183), .B2(n4417), .A(n4182), .ZN(n4239) );
  MUX2_X1 U4749 ( .A(n4184), .B(n4239), .S(n4443), .Z(n4185) );
  OAI21_X1 U4750 ( .B1(n4223), .B2(n4242), .A(n4185), .ZN(U3544) );
  INV_X1 U4751 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4188) );
  AOI21_X1 U4752 ( .B1(n4187), .B2(n4417), .A(n4186), .ZN(n4243) );
  MUX2_X1 U4753 ( .A(n4188), .B(n4243), .S(n4443), .Z(n4189) );
  OAI21_X1 U4754 ( .B1(n4223), .B2(n4246), .A(n4189), .ZN(U3543) );
  INV_X1 U4755 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4192) );
  AOI21_X1 U4756 ( .B1(n4191), .B2(n4417), .A(n4190), .ZN(n4247) );
  MUX2_X1 U4757 ( .A(n4192), .B(n4247), .S(n4443), .Z(n4193) );
  OAI21_X1 U4758 ( .B1(n4223), .B2(n4249), .A(n4193), .ZN(U3542) );
  INV_X1 U4759 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4196) );
  AOI21_X1 U4760 ( .B1(n4195), .B2(n4417), .A(n4194), .ZN(n4250) );
  MUX2_X1 U4761 ( .A(n4196), .B(n4250), .S(n4443), .Z(n4197) );
  OAI21_X1 U4762 ( .B1(n4223), .B2(n4253), .A(n4197), .ZN(U3541) );
  NAND3_X1 U4763 ( .A1(n4199), .A2(n2619), .A3(n4198), .ZN(n4200) );
  OAI211_X1 U4764 ( .C1(n4202), .C2(n4411), .A(n4201), .B(n4200), .ZN(n4254)
         );
  MUX2_X1 U4765 ( .A(REG1_REG_22__SCAN_IN), .B(n4254), .S(n4443), .Z(U3540) );
  INV_X1 U4766 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4553) );
  AOI21_X1 U4767 ( .B1(n4204), .B2(n4417), .A(n4203), .ZN(n4255) );
  MUX2_X1 U4768 ( .A(n4553), .B(n4255), .S(n4443), .Z(n4205) );
  OAI21_X1 U4769 ( .B1(n4223), .B2(n4258), .A(n4205), .ZN(U3539) );
  INV_X1 U4770 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4552) );
  INV_X1 U4771 ( .A(n4206), .ZN(n4208) );
  AOI21_X1 U4772 ( .B1(n4402), .B2(n4208), .A(n4207), .ZN(n4259) );
  MUX2_X1 U4773 ( .A(n4552), .B(n4259), .S(n4443), .Z(n4209) );
  OAI21_X1 U4774 ( .B1(n4223), .B2(n4262), .A(n4209), .ZN(U3538) );
  INV_X1 U4775 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4212) );
  AOI21_X1 U4776 ( .B1(n4211), .B2(n4417), .A(n4210), .ZN(n4263) );
  MUX2_X1 U4777 ( .A(n4212), .B(n4263), .S(n4443), .Z(n4213) );
  OAI21_X1 U4778 ( .B1(n4223), .B2(n4266), .A(n4213), .ZN(U3537) );
  NAND2_X1 U4779 ( .A1(n4214), .A2(n4417), .ZN(n4218) );
  NOR2_X1 U4780 ( .A1(n4216), .A2(n4215), .ZN(n4217) );
  NAND2_X1 U4781 ( .A1(n4218), .A2(n4217), .ZN(n4267) );
  MUX2_X1 U4782 ( .A(n4267), .B(REG1_REG_18__SCAN_IN), .S(n4441), .Z(U3536) );
  INV_X1 U4783 ( .A(n4219), .ZN(n4220) );
  AOI21_X1 U4784 ( .B1(n4221), .B2(n4417), .A(n4220), .ZN(n4268) );
  MUX2_X1 U4785 ( .A(n4551), .B(n4268), .S(n4443), .Z(n4222) );
  OAI21_X1 U4786 ( .B1(n4223), .B2(n4272), .A(n4222), .ZN(U3535) );
  AOI21_X1 U4787 ( .B1(n2619), .B2(n4225), .A(n4224), .ZN(n4226) );
  OAI21_X1 U4788 ( .B1(n4227), .B2(n4411), .A(n4226), .ZN(n4273) );
  MUX2_X1 U4789 ( .A(REG1_REG_16__SCAN_IN), .B(n4273), .S(n4443), .Z(U3534) );
  AOI21_X1 U4790 ( .B1(n2619), .B2(n4229), .A(n4228), .ZN(n4230) );
  OAI21_X1 U4791 ( .B1(n4231), .B2(n4411), .A(n4230), .ZN(n4274) );
  MUX2_X1 U4792 ( .A(REG1_REG_15__SCAN_IN), .B(n4274), .S(n4443), .Z(U3533) );
  INV_X1 U4793 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4232) );
  MUX2_X1 U4794 ( .A(n4232), .B(n4290), .S(n4431), .Z(n4233) );
  OAI21_X1 U4795 ( .B1(n4234), .B2(n4271), .A(n4233), .ZN(U3517) );
  INV_X1 U4796 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4488) );
  MUX2_X1 U4797 ( .A(n4488), .B(n4293), .S(n4431), .Z(n4235) );
  OAI21_X1 U4798 ( .B1(n4236), .B2(n4271), .A(n4235), .ZN(U3516) );
  MUX2_X1 U4799 ( .A(REG0_REG_29__SCAN_IN), .B(n4237), .S(n4431), .Z(U3515) );
  MUX2_X1 U4800 ( .A(REG0_REG_27__SCAN_IN), .B(n4238), .S(n4431), .Z(U3513) );
  INV_X1 U4801 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4240) );
  MUX2_X1 U4802 ( .A(n4240), .B(n4239), .S(n4431), .Z(n4241) );
  OAI21_X1 U4803 ( .B1(n4242), .B2(n4271), .A(n4241), .ZN(U3512) );
  INV_X1 U4804 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4244) );
  MUX2_X1 U4805 ( .A(n4244), .B(n4243), .S(n4431), .Z(n4245) );
  OAI21_X1 U4806 ( .B1(n4246), .B2(n4271), .A(n4245), .ZN(U3511) );
  INV_X1 U4807 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4489) );
  MUX2_X1 U4808 ( .A(n4489), .B(n4247), .S(n4431), .Z(n4248) );
  OAI21_X1 U4809 ( .B1(n4249), .B2(n4271), .A(n4248), .ZN(U3510) );
  INV_X1 U4810 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4251) );
  MUX2_X1 U4811 ( .A(n4251), .B(n4250), .S(n4431), .Z(n4252) );
  OAI21_X1 U4812 ( .B1(n4253), .B2(n4271), .A(n4252), .ZN(U3509) );
  MUX2_X1 U4813 ( .A(REG0_REG_22__SCAN_IN), .B(n4254), .S(n4431), .Z(U3508) );
  INV_X1 U4814 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4256) );
  MUX2_X1 U4815 ( .A(n4256), .B(n4255), .S(n4431), .Z(n4257) );
  OAI21_X1 U4816 ( .B1(n4258), .B2(n4271), .A(n4257), .ZN(U3507) );
  INV_X1 U4817 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4260) );
  MUX2_X1 U4818 ( .A(n4260), .B(n4259), .S(n4431), .Z(n4261) );
  OAI21_X1 U4819 ( .B1(n4262), .B2(n4271), .A(n4261), .ZN(U3506) );
  INV_X1 U4820 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4264) );
  MUX2_X1 U4821 ( .A(n4264), .B(n4263), .S(n4431), .Z(n4265) );
  OAI21_X1 U4822 ( .B1(n4266), .B2(n4271), .A(n4265), .ZN(U3505) );
  MUX2_X1 U4823 ( .A(n4267), .B(REG0_REG_18__SCAN_IN), .S(n4429), .Z(U3503) );
  INV_X1 U4824 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4269) );
  MUX2_X1 U4825 ( .A(n4269), .B(n4268), .S(n4431), .Z(n4270) );
  OAI21_X1 U4826 ( .B1(n4272), .B2(n4271), .A(n4270), .ZN(U3501) );
  MUX2_X1 U4827 ( .A(REG0_REG_16__SCAN_IN), .B(n4273), .S(n4431), .Z(U3499) );
  MUX2_X1 U4828 ( .A(REG0_REG_15__SCAN_IN), .B(n4274), .S(n4431), .Z(U3497) );
  MUX2_X1 U4829 ( .A(DATAI_29_), .B(n2239), .S(STATE_REG_SCAN_IN), .Z(U3323)
         );
  MUX2_X1 U4830 ( .A(DATAI_27_), .B(n4275), .S(STATE_REG_SCAN_IN), .Z(U3325)
         );
  MUX2_X1 U4831 ( .A(DATAI_24_), .B(n2584), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U4832 ( .A(DATAI_22_), .B(n4276), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U4833 ( .A(DATAI_19_), .B(n4277), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U4834 ( .A(n4278), .B(DATAI_15_), .S(U3149), .Z(U3337) );
  MUX2_X1 U4835 ( .A(n4279), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U4836 ( .A(n4280), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U4837 ( .A(n4281), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  INV_X1 U4838 ( .A(n4282), .ZN(n4283) );
  MUX2_X1 U4839 ( .A(DATAI_5_), .B(n4283), .S(STATE_REG_SCAN_IN), .Z(U3347) );
  MUX2_X1 U4840 ( .A(DATAI_4_), .B(n4284), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4841 ( .A(n4285), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4842 ( .A(n4286), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  AOI22_X1 U4843 ( .A1(STATE_REG_SCAN_IN), .A2(n4287), .B1(n2518), .B2(U3149), 
        .ZN(U3324) );
  AOI22_X1 U4844 ( .A1(n4288), .A2(n4362), .B1(n4377), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n4289) );
  OAI21_X1 U4845 ( .B1(n4377), .B2(n4290), .A(n4289), .ZN(U3260) );
  AOI22_X1 U4846 ( .A1(n4291), .A2(n4362), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4377), .ZN(n4292) );
  OAI21_X1 U4847 ( .B1(n4377), .B2(n4293), .A(n4292), .ZN(U3261) );
  AOI211_X1 U4848 ( .C1(n4491), .C2(n4295), .A(n4294), .B(n4321), .ZN(n4297)
         );
  AOI211_X1 U4849 ( .C1(n4345), .C2(ADDR_REG_10__SCAN_IN), .A(n4297), .B(n4296), .ZN(n4301) );
  OAI211_X1 U4850 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4299), .A(n4355), .B(n4298), .ZN(n4300) );
  OAI211_X1 U4851 ( .C1(n4358), .C2(n4388), .A(n4301), .B(n4300), .ZN(U3250)
         );
  AOI211_X1 U4852 ( .C1(n4304), .C2(n4303), .A(n4302), .B(n4321), .ZN(n4306)
         );
  AOI211_X1 U4853 ( .C1(n4345), .C2(ADDR_REG_11__SCAN_IN), .A(n4306), .B(n4305), .ZN(n4311) );
  OAI211_X1 U4854 ( .C1(n4309), .C2(n4308), .A(n4355), .B(n4307), .ZN(n4310)
         );
  OAI211_X1 U4855 ( .C1(n4358), .C2(n4312), .A(n4311), .B(n4310), .ZN(U3251)
         );
  AOI211_X1 U4856 ( .C1(n4502), .C2(n4314), .A(n4313), .B(n4321), .ZN(n4316)
         );
  AOI211_X1 U4857 ( .C1(n4345), .C2(ADDR_REG_12__SCAN_IN), .A(n4316), .B(n4315), .ZN(n4320) );
  OAI211_X1 U4858 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4318), .A(n4355), .B(n4317), .ZN(n4319) );
  OAI211_X1 U4859 ( .C1(n4358), .C2(n2156), .A(n4320), .B(n4319), .ZN(U3252)
         );
  INV_X1 U4860 ( .A(n4345), .ZN(n4333) );
  INV_X1 U4861 ( .A(ADDR_REG_14__SCAN_IN), .ZN(n4562) );
  AOI211_X1 U4862 ( .C1(n4501), .C2(n4323), .A(n4322), .B(n4321), .ZN(n4328)
         );
  AOI211_X1 U4863 ( .C1(n3320), .C2(n4326), .A(n4325), .B(n4324), .ZN(n4327)
         );
  AOI211_X1 U4864 ( .C1(n4330), .C2(n4329), .A(n4328), .B(n4327), .ZN(n4332)
         );
  OAI211_X1 U4865 ( .C1(n4333), .C2(n4562), .A(n4332), .B(n4331), .ZN(U3254)
         );
  AOI21_X1 U4866 ( .B1(n4345), .B2(ADDR_REG_16__SCAN_IN), .A(n4334), .ZN(n4343) );
  OAI21_X1 U4867 ( .B1(n4336), .B2(n3402), .A(n4335), .ZN(n4341) );
  OAI21_X1 U4868 ( .B1(n4339), .B2(n4338), .A(n4337), .ZN(n4340) );
  AOI22_X1 U4869 ( .A1(n4355), .A2(n4341), .B1(n4353), .B2(n4340), .ZN(n4342)
         );
  OAI211_X1 U4870 ( .C1(n4384), .C2(n4358), .A(n4343), .B(n4342), .ZN(U3256)
         );
  AOI21_X1 U4871 ( .B1(n4345), .B2(ADDR_REG_17__SCAN_IN), .A(n4344), .ZN(n4357) );
  OAI21_X1 U4872 ( .B1(n4348), .B2(n4347), .A(n4346), .ZN(n4354) );
  OAI21_X1 U4873 ( .B1(n4351), .B2(n4350), .A(n4349), .ZN(n4352) );
  AOI22_X1 U4874 ( .A1(n4355), .A2(n4354), .B1(n4353), .B2(n4352), .ZN(n4356)
         );
  OAI211_X1 U4875 ( .C1(n4382), .C2(n4358), .A(n4357), .B(n4356), .ZN(U3257)
         );
  AOI22_X1 U4876 ( .A1(REG2_REG_2__SCAN_IN), .A2(n4377), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4371), .ZN(n4365) );
  INV_X1 U4877 ( .A(n4359), .ZN(n4363) );
  INV_X1 U4878 ( .A(n4360), .ZN(n4361) );
  AOI22_X1 U4879 ( .A1(n4363), .A2(n4373), .B1(n4362), .B2(n4361), .ZN(n4364)
         );
  OAI211_X1 U4880 ( .C1(n4377), .C2(n4366), .A(n4365), .B(n4364), .ZN(U3288)
         );
  INV_X1 U4881 ( .A(n4367), .ZN(n4369) );
  AOI21_X1 U4882 ( .B1(n4370), .B2(n4369), .A(n4368), .ZN(n4376) );
  AOI22_X1 U4883 ( .A1(n4373), .A2(n4372), .B1(REG3_REG_0__SCAN_IN), .B2(n4371), .ZN(n4374) );
  OAI221_X1 U4884 ( .B1(n4377), .B2(n4376), .C1(n4375), .C2(n2942), .A(n4374), 
        .ZN(U3290) );
  INV_X1 U4885 ( .A(n4378), .ZN(n4379) );
  INV_X1 U4886 ( .A(D_REG_31__SCAN_IN), .ZN(n4483) );
  NOR2_X1 U4887 ( .A1(n4379), .A2(n4483), .ZN(U3291) );
  AND2_X1 U4888 ( .A1(D_REG_30__SCAN_IN), .A2(n4378), .ZN(U3292) );
  AND2_X1 U4889 ( .A1(D_REG_29__SCAN_IN), .A2(n4378), .ZN(U3293) );
  AND2_X1 U4890 ( .A1(D_REG_28__SCAN_IN), .A2(n4378), .ZN(U3294) );
  AND2_X1 U4891 ( .A1(D_REG_27__SCAN_IN), .A2(n4378), .ZN(U3295) );
  AND2_X1 U4892 ( .A1(D_REG_26__SCAN_IN), .A2(n4378), .ZN(U3296) );
  AND2_X1 U4893 ( .A1(D_REG_25__SCAN_IN), .A2(n4378), .ZN(U3297) );
  AND2_X1 U4894 ( .A1(D_REG_24__SCAN_IN), .A2(n4378), .ZN(U3298) );
  AND2_X1 U4895 ( .A1(D_REG_23__SCAN_IN), .A2(n4378), .ZN(U3299) );
  AND2_X1 U4896 ( .A1(D_REG_22__SCAN_IN), .A2(n4378), .ZN(U3300) );
  AND2_X1 U4897 ( .A1(D_REG_21__SCAN_IN), .A2(n4378), .ZN(U3301) );
  AND2_X1 U4898 ( .A1(D_REG_20__SCAN_IN), .A2(n4378), .ZN(U3302) );
  AND2_X1 U4899 ( .A1(D_REG_19__SCAN_IN), .A2(n4378), .ZN(U3303) );
  AND2_X1 U4900 ( .A1(D_REG_18__SCAN_IN), .A2(n4378), .ZN(U3304) );
  AND2_X1 U4901 ( .A1(D_REG_17__SCAN_IN), .A2(n4378), .ZN(U3305) );
  INV_X1 U4902 ( .A(D_REG_16__SCAN_IN), .ZN(n4475) );
  NOR2_X1 U4903 ( .A1(n4379), .A2(n4475), .ZN(U3306) );
  INV_X1 U4904 ( .A(D_REG_15__SCAN_IN), .ZN(n4474) );
  NOR2_X1 U4905 ( .A1(n4379), .A2(n4474), .ZN(U3307) );
  AND2_X1 U4906 ( .A1(D_REG_14__SCAN_IN), .A2(n4378), .ZN(U3308) );
  AND2_X1 U4907 ( .A1(D_REG_13__SCAN_IN), .A2(n4378), .ZN(U3309) );
  AND2_X1 U4908 ( .A1(D_REG_12__SCAN_IN), .A2(n4378), .ZN(U3310) );
  AND2_X1 U4909 ( .A1(D_REG_11__SCAN_IN), .A2(n4378), .ZN(U3311) );
  AND2_X1 U4910 ( .A1(D_REG_10__SCAN_IN), .A2(n4378), .ZN(U3312) );
  AND2_X1 U4911 ( .A1(D_REG_9__SCAN_IN), .A2(n4378), .ZN(U3313) );
  AND2_X1 U4912 ( .A1(D_REG_8__SCAN_IN), .A2(n4378), .ZN(U3314) );
  AND2_X1 U4913 ( .A1(D_REG_7__SCAN_IN), .A2(n4378), .ZN(U3315) );
  AND2_X1 U4914 ( .A1(D_REG_6__SCAN_IN), .A2(n4378), .ZN(U3316) );
  AND2_X1 U4915 ( .A1(D_REG_5__SCAN_IN), .A2(n4378), .ZN(U3317) );
  INV_X1 U4916 ( .A(D_REG_4__SCAN_IN), .ZN(n4582) );
  NOR2_X1 U4917 ( .A1(n4379), .A2(n4582), .ZN(U3318) );
  AND2_X1 U4918 ( .A1(D_REG_3__SCAN_IN), .A2(n4378), .ZN(U3319) );
  INV_X1 U4919 ( .A(D_REG_2__SCAN_IN), .ZN(n4470) );
  NOR2_X1 U4920 ( .A1(n4379), .A2(n4470), .ZN(U3320) );
  INV_X1 U4921 ( .A(DATAI_23_), .ZN(n4381) );
  AOI21_X1 U4922 ( .B1(U3149), .B2(n4381), .A(n4380), .ZN(U3329) );
  AOI22_X1 U4923 ( .A1(STATE_REG_SCAN_IN), .A2(n4382), .B1(n2430), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U4924 ( .A(DATAI_16_), .ZN(n4383) );
  AOI22_X1 U4925 ( .A1(STATE_REG_SCAN_IN), .A2(n4384), .B1(n4383), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U4926 ( .A(DATAI_14_), .ZN(n4452) );
  AOI22_X1 U4927 ( .A1(STATE_REG_SCAN_IN), .A2(n4385), .B1(n4452), .B2(U3149), 
        .ZN(U3338) );
  OAI22_X1 U4928 ( .A1(U3149), .A2(n4386), .B1(DATAI_11_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4387) );
  INV_X1 U4929 ( .A(n4387), .ZN(U3341) );
  INV_X1 U4930 ( .A(DATAI_10_), .ZN(n4453) );
  AOI22_X1 U4931 ( .A1(STATE_REG_SCAN_IN), .A2(n4388), .B1(n4453), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U4932 ( .A(DATAI_0_), .ZN(n4389) );
  AOI22_X1 U4933 ( .A1(STATE_REG_SCAN_IN), .A2(n4390), .B1(n4389), .B2(U3149), 
        .ZN(U3352) );
  INV_X1 U4934 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4391) );
  AOI22_X1 U4935 ( .A1(n4431), .A2(n4392), .B1(n4391), .B2(n4429), .ZN(U3467)
         );
  INV_X1 U4936 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4393) );
  AOI22_X1 U4937 ( .A1(n4431), .A2(n4394), .B1(n4393), .B2(n4429), .ZN(U3469)
         );
  OAI22_X1 U4938 ( .A1(n4396), .A2(n4425), .B1(n4424), .B2(n4395), .ZN(n4397)
         );
  NOR2_X1 U4939 ( .A1(n4398), .A2(n4397), .ZN(n4433) );
  INV_X1 U4940 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4399) );
  AOI22_X1 U4941 ( .A1(n4431), .A2(n4433), .B1(n4399), .B2(n4429), .ZN(U3473)
         );
  AOI211_X1 U4942 ( .C1(n4403), .C2(n4402), .A(n4401), .B(n4400), .ZN(n4435)
         );
  INV_X1 U4943 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4404) );
  AOI22_X1 U4944 ( .A1(n4431), .A2(n4435), .B1(n4404), .B2(n4429), .ZN(U3475)
         );
  INV_X1 U4945 ( .A(n4405), .ZN(n4408) );
  NOR2_X1 U4946 ( .A1(n4406), .A2(n4411), .ZN(n4407) );
  AOI211_X1 U4947 ( .C1(n2619), .C2(n4409), .A(n4408), .B(n4407), .ZN(n4436)
         );
  INV_X1 U4948 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4410) );
  AOI22_X1 U4949 ( .A1(n4431), .A2(n4436), .B1(n4410), .B2(n4429), .ZN(U3477)
         );
  NOR2_X1 U4950 ( .A1(n4412), .A2(n4411), .ZN(n4415) );
  AOI211_X1 U4951 ( .C1(n4415), .C2(n3140), .A(n4414), .B(n4413), .ZN(n4438)
         );
  INV_X1 U4952 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4416) );
  AOI22_X1 U4953 ( .A1(n4431), .A2(n4438), .B1(n4416), .B2(n4429), .ZN(U3481)
         );
  NAND2_X1 U4954 ( .A1(n4418), .A2(n4417), .ZN(n4422) );
  NAND2_X1 U4955 ( .A1(n4419), .A2(n2619), .ZN(n4420) );
  INV_X1 U4956 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4486) );
  AOI22_X1 U4957 ( .A1(n4431), .A2(n4440), .B1(n4486), .B2(n4429), .ZN(U3485)
         );
  OAI22_X1 U4958 ( .A1(n4426), .A2(n4425), .B1(n4424), .B2(n4423), .ZN(n4427)
         );
  NOR2_X1 U4959 ( .A1(n4428), .A2(n4427), .ZN(n4442) );
  INV_X1 U4960 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4430) );
  AOI22_X1 U4961 ( .A1(n4431), .A2(n4442), .B1(n4430), .B2(n4429), .ZN(U3489)
         );
  INV_X1 U4962 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4432) );
  AOI22_X1 U4963 ( .A1(n4443), .A2(n4433), .B1(n4432), .B2(n4441), .ZN(U3521)
         );
  INV_X1 U4964 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4434) );
  AOI22_X1 U4965 ( .A1(n4443), .A2(n4435), .B1(n4434), .B2(n4441), .ZN(U3522)
         );
  AOI22_X1 U4966 ( .A1(n4443), .A2(n4436), .B1(n2912), .B2(n4441), .ZN(U3523)
         );
  AOI22_X1 U4967 ( .A1(n4443), .A2(n4438), .B1(n4437), .B2(n4441), .ZN(U3525)
         );
  INV_X1 U4968 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4439) );
  AOI22_X1 U4969 ( .A1(n4443), .A2(n4440), .B1(n4439), .B2(n4441), .ZN(U3527)
         );
  AOI22_X1 U4970 ( .A1(n4443), .A2(n4442), .B1(n4577), .B2(n4441), .ZN(U3529)
         );
  AOI22_X1 U4971 ( .A1(STATE_REG_SCAN_IN), .A2(n4444), .B1(DATAI_12_), .B2(
        U3149), .ZN(n4597) );
  INV_X1 U4972 ( .A(DATAI_24_), .ZN(n4447) );
  AOI22_X1 U4973 ( .A1(n4447), .A2(keyinput17), .B1(keyinput2), .B2(n4446), 
        .ZN(n4445) );
  OAI221_X1 U4974 ( .B1(n4447), .B2(keyinput17), .C1(n4446), .C2(keyinput2), 
        .A(n4445), .ZN(n4457) );
  INV_X1 U4975 ( .A(DATAI_19_), .ZN(n4570) );
  INV_X1 U4976 ( .A(DATAI_22_), .ZN(n4571) );
  AOI22_X1 U4977 ( .A1(n4570), .A2(keyinput16), .B1(n4571), .B2(keyinput33), 
        .ZN(n4448) );
  OAI221_X1 U4978 ( .B1(n4570), .B2(keyinput16), .C1(n4571), .C2(keyinput33), 
        .A(n4448), .ZN(n4456) );
  AOI22_X1 U4979 ( .A1(n4450), .A2(keyinput1), .B1(n2430), .B2(keyinput48), 
        .ZN(n4449) );
  OAI221_X1 U4980 ( .B1(n4450), .B2(keyinput1), .C1(n2430), .C2(keyinput48), 
        .A(n4449), .ZN(n4455) );
  AOI22_X1 U4981 ( .A1(n4453), .A2(keyinput62), .B1(n4452), .B2(keyinput59), 
        .ZN(n4451) );
  OAI221_X1 U4982 ( .B1(n4453), .B2(keyinput62), .C1(n4452), .C2(keyinput59), 
        .A(n4451), .ZN(n4454) );
  NOR4_X1 U4983 ( .A1(n4457), .A2(n4456), .A3(n4455), .A4(n4454), .ZN(n4499)
         );
  INV_X1 U4984 ( .A(IR_REG_1__SCAN_IN), .ZN(n4573) );
  AOI22_X1 U4985 ( .A1(n4572), .A2(keyinput29), .B1(n4573), .B2(keyinput11), 
        .ZN(n4458) );
  OAI221_X1 U4986 ( .B1(n4572), .B2(keyinput29), .C1(n4573), .C2(keyinput11), 
        .A(n4458), .ZN(n4468) );
  AOI22_X1 U4987 ( .A1(U3149), .A2(keyinput61), .B1(keyinput22), .B2(n2278), 
        .ZN(n4459) );
  OAI221_X1 U4988 ( .B1(U3149), .B2(keyinput61), .C1(n2278), .C2(keyinput22), 
        .A(n4459), .ZN(n4467) );
  AOI22_X1 U4989 ( .A1(n4462), .A2(keyinput39), .B1(n4461), .B2(keyinput20), 
        .ZN(n4460) );
  OAI221_X1 U4990 ( .B1(n4462), .B2(keyinput39), .C1(n4461), .C2(keyinput20), 
        .A(n4460), .ZN(n4466) );
  XOR2_X1 U4991 ( .A(n2324), .B(keyinput8), .Z(n4464) );
  XNOR2_X1 U4992 ( .A(IR_REG_4__SCAN_IN), .B(keyinput6), .ZN(n4463) );
  NAND2_X1 U4993 ( .A1(n4464), .A2(n4463), .ZN(n4465) );
  NOR4_X1 U4994 ( .A1(n4468), .A2(n4467), .A3(n4466), .A4(n4465), .ZN(n4498)
         );
  AOI22_X1 U4995 ( .A1(n4470), .A2(keyinput31), .B1(keyinput38), .B2(n4582), 
        .ZN(n4469) );
  OAI221_X1 U4996 ( .B1(n4470), .B2(keyinput31), .C1(n4582), .C2(keyinput38), 
        .A(n4469), .ZN(n4481) );
  AOI22_X1 U4997 ( .A1(n4578), .A2(keyinput21), .B1(n4472), .B2(keyinput32), 
        .ZN(n4471) );
  OAI221_X1 U4998 ( .B1(n4578), .B2(keyinput21), .C1(n4472), .C2(keyinput32), 
        .A(n4471), .ZN(n4480) );
  AOI22_X1 U4999 ( .A1(n4475), .A2(keyinput15), .B1(keyinput60), .B2(n4474), 
        .ZN(n4473) );
  OAI221_X1 U5000 ( .B1(n4475), .B2(keyinput15), .C1(n4474), .C2(keyinput60), 
        .A(n4473), .ZN(n4479) );
  XOR2_X1 U5001 ( .A(n2520), .B(keyinput40), .Z(n4477) );
  XNOR2_X1 U5002 ( .A(IR_REG_16__SCAN_IN), .B(keyinput50), .ZN(n4476) );
  NAND2_X1 U5003 ( .A1(n4477), .A2(n4476), .ZN(n4478) );
  NOR4_X1 U5004 ( .A1(n4481), .A2(n4480), .A3(n4479), .A4(n4478), .ZN(n4497)
         );
  AOI22_X1 U5005 ( .A1(n4576), .A2(keyinput42), .B1(n4483), .B2(keyinput56), 
        .ZN(n4482) );
  OAI221_X1 U5006 ( .B1(n4576), .B2(keyinput42), .C1(n4483), .C2(keyinput56), 
        .A(n4482), .ZN(n4495) );
  INV_X1 U5007 ( .A(REG0_REG_18__SCAN_IN), .ZN(n4485) );
  AOI22_X1 U5008 ( .A1(n4486), .A2(keyinput54), .B1(keyinput26), .B2(n4485), 
        .ZN(n4484) );
  OAI221_X1 U5009 ( .B1(n4486), .B2(keyinput54), .C1(n4485), .C2(keyinput26), 
        .A(n4484), .ZN(n4494) );
  AOI22_X1 U5010 ( .A1(n4489), .A2(keyinput36), .B1(keyinput10), .B2(n4488), 
        .ZN(n4487) );
  OAI221_X1 U5011 ( .B1(n4489), .B2(keyinput36), .C1(n4488), .C2(keyinput10), 
        .A(n4487), .ZN(n4493) );
  AOI22_X1 U5012 ( .A1(n4577), .A2(keyinput3), .B1(keyinput58), .B2(n4491), 
        .ZN(n4490) );
  OAI221_X1 U5013 ( .B1(n4577), .B2(keyinput3), .C1(n4491), .C2(keyinput58), 
        .A(n4490), .ZN(n4492) );
  NOR4_X1 U5014 ( .A1(n4495), .A2(n4494), .A3(n4493), .A4(n4492), .ZN(n4496)
         );
  NAND4_X1 U5015 ( .A1(n4499), .A2(n4498), .A3(n4497), .A4(n4496), .ZN(n4549)
         );
  AOI22_X1 U5016 ( .A1(n4502), .A2(keyinput25), .B1(n4501), .B2(keyinput24), 
        .ZN(n4500) );
  OAI221_X1 U5017 ( .B1(n4502), .B2(keyinput25), .C1(n4501), .C2(keyinput24), 
        .A(n4500), .ZN(n4511) );
  AOI22_X1 U5018 ( .A1(n4551), .A2(keyinput9), .B1(n4552), .B2(keyinput45), 
        .ZN(n4503) );
  OAI221_X1 U5019 ( .B1(n4551), .B2(keyinput9), .C1(n4552), .C2(keyinput45), 
        .A(n4503), .ZN(n4510) );
  AOI22_X1 U5020 ( .A1(n4553), .A2(keyinput34), .B1(keyinput5), .B2(n4505), 
        .ZN(n4504) );
  OAI221_X1 U5021 ( .B1(n4553), .B2(keyinput34), .C1(n4505), .C2(keyinput5), 
        .A(n4504), .ZN(n4509) );
  AOI22_X1 U5022 ( .A1(n2256), .A2(keyinput37), .B1(keyinput47), .B2(n4507), 
        .ZN(n4506) );
  OAI221_X1 U5023 ( .B1(n2256), .B2(keyinput37), .C1(n4507), .C2(keyinput47), 
        .A(n4506), .ZN(n4508) );
  NOR4_X1 U5024 ( .A1(n4511), .A2(n4510), .A3(n4509), .A4(n4508), .ZN(n4547)
         );
  AOI22_X1 U5025 ( .A1(n2294), .A2(keyinput35), .B1(keyinput18), .B2(n3157), 
        .ZN(n4512) );
  OAI221_X1 U5026 ( .B1(n2294), .B2(keyinput35), .C1(n3157), .C2(keyinput18), 
        .A(n4512), .ZN(n4520) );
  AOI22_X1 U5027 ( .A1(n4550), .A2(keyinput46), .B1(keyinput55), .B2(n3264), 
        .ZN(n4513) );
  OAI221_X1 U5028 ( .B1(n4550), .B2(keyinput46), .C1(n3264), .C2(keyinput55), 
        .A(n4513), .ZN(n4519) );
  AOI22_X1 U5029 ( .A1(n2489), .A2(keyinput28), .B1(keyinput0), .B2(n4044), 
        .ZN(n4514) );
  OAI221_X1 U5030 ( .B1(n2489), .B2(keyinput28), .C1(n4044), .C2(keyinput0), 
        .A(n4514), .ZN(n4518) );
  INV_X1 U5031 ( .A(ADDR_REG_19__SCAN_IN), .ZN(n4516) );
  AOI22_X1 U5032 ( .A1(n4516), .A2(keyinput51), .B1(n2498), .B2(keyinput30), 
        .ZN(n4515) );
  OAI221_X1 U5033 ( .B1(n4516), .B2(keyinput51), .C1(n2498), .C2(keyinput30), 
        .A(n4515), .ZN(n4517) );
  NOR4_X1 U5034 ( .A1(n4520), .A2(n4519), .A3(n4518), .A4(n4517), .ZN(n4546)
         );
  INV_X1 U5035 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n4522) );
  AOI22_X1 U5036 ( .A1(n4522), .A2(keyinput19), .B1(n4562), .B2(keyinput63), 
        .ZN(n4521) );
  OAI221_X1 U5037 ( .B1(n4522), .B2(keyinput19), .C1(n4562), .C2(keyinput63), 
        .A(n4521), .ZN(n4531) );
  INV_X1 U5038 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n4525) );
  INV_X1 U5039 ( .A(ADDR_REG_12__SCAN_IN), .ZN(n4524) );
  AOI22_X1 U5040 ( .A1(n4525), .A2(keyinput23), .B1(n4524), .B2(keyinput44), 
        .ZN(n4523) );
  OAI221_X1 U5041 ( .B1(n4525), .B2(keyinput23), .C1(n4524), .C2(keyinput44), 
        .A(n4523), .ZN(n4530) );
  AOI22_X1 U5042 ( .A1(n4566), .A2(keyinput13), .B1(keyinput12), .B2(n4564), 
        .ZN(n4526) );
  OAI221_X1 U5043 ( .B1(n4566), .B2(keyinput13), .C1(n4564), .C2(keyinput12), 
        .A(n4526), .ZN(n4529) );
  AOI22_X1 U5044 ( .A1(n4565), .A2(keyinput7), .B1(keyinput27), .B2(n4563), 
        .ZN(n4527) );
  OAI221_X1 U5045 ( .B1(n4565), .B2(keyinput7), .C1(n4563), .C2(keyinput27), 
        .A(n4527), .ZN(n4528) );
  NOR4_X1 U5046 ( .A1(n4531), .A2(n4530), .A3(n4529), .A4(n4528), .ZN(n4545)
         );
  AOI22_X1 U5047 ( .A1(n4533), .A2(keyinput14), .B1(n4561), .B2(keyinput49), 
        .ZN(n4532) );
  OAI221_X1 U5048 ( .B1(n4533), .B2(keyinput14), .C1(n4561), .C2(keyinput49), 
        .A(n4532), .ZN(n4543) );
  AOI22_X1 U5049 ( .A1(n4535), .A2(keyinput43), .B1(n4560), .B2(keyinput57), 
        .ZN(n4534) );
  OAI221_X1 U5050 ( .B1(n4535), .B2(keyinput43), .C1(n4560), .C2(keyinput57), 
        .A(n4534), .ZN(n4542) );
  AOI22_X1 U5051 ( .A1(n4559), .A2(keyinput41), .B1(keyinput52), .B2(n4558), 
        .ZN(n4536) );
  OAI221_X1 U5052 ( .B1(n4559), .B2(keyinput41), .C1(n4558), .C2(keyinput52), 
        .A(n4536), .ZN(n4541) );
  INV_X1 U5053 ( .A(B_REG_SCAN_IN), .ZN(n4538) );
  AOI22_X1 U5054 ( .A1(n4539), .A2(keyinput53), .B1(n4538), .B2(keyinput4), 
        .ZN(n4537) );
  OAI221_X1 U5055 ( .B1(n4539), .B2(keyinput53), .C1(n4538), .C2(keyinput4), 
        .A(n4537), .ZN(n4540) );
  NOR4_X1 U5056 ( .A1(n4543), .A2(n4542), .A3(n4541), .A4(n4540), .ZN(n4544)
         );
  NAND4_X1 U5057 ( .A1(n4547), .A2(n4546), .A3(n4545), .A4(n4544), .ZN(n4548)
         );
  NOR2_X1 U5058 ( .A1(n4549), .A2(n4548), .ZN(n4595) );
  NAND4_X1 U5059 ( .A1(REG2_REG_12__SCAN_IN), .A2(REG2_REG_5__SCAN_IN), .A3(
        n4550), .A4(n2294), .ZN(n4557) );
  NAND4_X1 U5060 ( .A1(REG2_REG_26__SCAN_IN), .A2(REG2_REG_22__SCAN_IN), .A3(
        ADDR_REG_19__SCAN_IN), .A4(n2489), .ZN(n4556) );
  NAND4_X1 U5061 ( .A1(REG1_REG_14__SCAN_IN), .A2(REG1_REG_12__SCAN_IN), .A3(
        n4552), .A4(n4551), .ZN(n4555) );
  NAND4_X1 U5062 ( .A1(REG2_REG_3__SCAN_IN), .A2(REG1_REG_30__SCAN_IN), .A3(
        REG1_REG_31__SCAN_IN), .A4(n4553), .ZN(n4554) );
  NOR4_X1 U5063 ( .A1(n4557), .A2(n4556), .A3(n4555), .A4(n4554), .ZN(n4593)
         );
  NOR4_X1 U5064 ( .A1(B_REG_SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .A3(n4559), 
        .A4(n4558), .ZN(n4592) );
  NAND4_X1 U5065 ( .A1(DATAO_REG_19__SCAN_IN), .A2(DATAO_REG_26__SCAN_IN), 
        .A3(n4561), .A4(n4560), .ZN(n4569) );
  NAND3_X1 U5066 ( .A1(ADDR_REG_13__SCAN_IN), .A2(ADDR_REG_12__SCAN_IN), .A3(
        n4562), .ZN(n4568) );
  NAND4_X1 U5067 ( .A1(n4566), .A2(n4565), .A3(n4564), .A4(n4563), .ZN(n4567)
         );
  NOR4_X1 U5068 ( .A1(ADDR_REG_5__SCAN_IN), .A2(n4569), .A3(n4568), .A4(n4567), 
        .ZN(n4591) );
  NAND4_X1 U5069 ( .A1(IR_REG_4__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .A3(
        REG3_REG_3__SCAN_IN), .A4(n2324), .ZN(n4589) );
  NAND4_X1 U5070 ( .A1(n4572), .A2(n4571), .A3(n4570), .A4(n2278), .ZN(n4588)
         );
  NOR4_X1 U5071 ( .A1(DATAI_14_), .A2(DATAI_10_), .A3(DATAI_24_), .A4(
        DATAI_31_), .ZN(n4574) );
  NAND4_X1 U5072 ( .A1(n4575), .A2(STATE_REG_SCAN_IN), .A3(n4574), .A4(n4573), 
        .ZN(n4587) );
  NOR4_X1 U5073 ( .A1(D_REG_31__SCAN_IN), .A2(REG1_REG_10__SCAN_IN), .A3(n4577), .A4(n4576), .ZN(n4585) );
  NOR4_X1 U5074 ( .A1(D_REG_1__SCAN_IN), .A2(REG0_REG_24__SCAN_IN), .A3(
        REG0_REG_30__SCAN_IN), .A4(n4578), .ZN(n4584) );
  NOR4_X1 U5075 ( .A1(DATAI_17_), .A2(REG0_REG_9__SCAN_IN), .A3(
        REG0_REG_18__SCAN_IN), .A4(DATAI_18_), .ZN(n4579) );
  NAND2_X1 U5076 ( .A1(n2520), .A2(n4579), .ZN(n4581) );
  NOR4_X1 U5077 ( .A1(n4582), .A2(n4581), .A3(n4580), .A4(D_REG_2__SCAN_IN), 
        .ZN(n4583) );
  NAND3_X1 U5078 ( .A1(n4585), .A2(n4584), .A3(n4583), .ZN(n4586) );
  NOR4_X1 U5079 ( .A1(n4589), .A2(n4588), .A3(n4587), .A4(n4586), .ZN(n4590)
         );
  NAND4_X1 U5080 ( .A1(n4593), .A2(n4592), .A3(n4591), .A4(n4590), .ZN(n4594)
         );
  XNOR2_X1 U5081 ( .A(n4595), .B(n4594), .ZN(n4596) );
  XNOR2_X1 U5082 ( .A(n4597), .B(n4596), .ZN(U3340) );
  CLKBUF_X2 U2246 ( .A(n2897), .Z(U4043) );
  INV_X2 U3879 ( .A(n4377), .ZN(n4375) );
endmodule

