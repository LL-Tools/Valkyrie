

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983;

  MUX2_X1 U7283 ( .A(n10412), .B(n9377), .S(n15886), .Z(n9374) );
  AND2_X1 U7284 ( .A1(n7362), .A2(n7363), .ZN(n10026) );
  NAND2_X1 U7285 ( .A1(n13501), .A2(n13499), .ZN(n13788) );
  NAND2_X1 U7286 ( .A1(n14595), .A2(n14166), .ZN(n9193) );
  AND2_X1 U7287 ( .A1(n13858), .A2(n8659), .ZN(n8660) );
  AND2_X1 U7288 ( .A1(n8658), .A2(n8657), .ZN(n13858) );
  CLKBUF_X2 U7289 ( .A(n9437), .Z(n9954) );
  INV_X1 U7290 ( .A(n12251), .ZN(n6548) );
  NAND4_X1 U7291 ( .A1(n9616), .A2(n9615), .A3(n9614), .A4(n9613), .ZN(n14954)
         );
  OAI21_X1 U7292 ( .B1(n9409), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9402) );
  AND2_X1 U7293 ( .A1(n8737), .A2(n8736), .ZN(n6600) );
  NAND4_X2 U7294 ( .A1(n8895), .A2(n8894), .A3(n8893), .A4(n8892), .ZN(n12775)
         );
  NAND2_X1 U7295 ( .A1(n10626), .A2(n9260), .ZN(n9169) );
  XNOR2_X1 U7296 ( .A(n6984), .B(n8782), .ZN(n10637) );
  INV_X2 U7297 ( .A(n10481), .ZN(n8129) );
  XNOR2_X1 U7298 ( .A(n9435), .B(P1_IR_REG_22__SCAN_IN), .ZN(n15553) );
  AND4_X1 U7299 ( .A1(n8847), .A2(n8773), .A3(n8772), .A4(n8771), .ZN(n8777)
         );
  NOR2_X1 U7300 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n8774) );
  NOR2_X1 U7301 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n8770) );
  CLKBUF_X2 U7302 ( .A(n12821), .Z(n6542) );
  OR2_X1 U7303 ( .A1(n13774), .A2(n7676), .ZN(n7363) );
  INV_X1 U7304 ( .A(n13965), .ZN(n8154) );
  INV_X2 U7305 ( .A(n9437), .ZN(n9923) );
  INV_X1 U7306 ( .A(n13514), .ZN(n13519) );
  AND2_X1 U7307 ( .A1(n14323), .A2(n7914), .ZN(n10015) );
  OAI21_X1 U7308 ( .B1(n14450), .B2(n7124), .A(n7122), .ZN(n14425) );
  NAND2_X1 U7309 ( .A1(n8853), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8948) );
  NAND2_X2 U7310 ( .A1(n10626), .A2(n8129), .ZN(n8902) );
  INV_X2 U7311 ( .A(n7327), .ZN(n9123) );
  NOR2_X1 U7312 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n8768) );
  NOR2_X1 U7313 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n8769) );
  NOR2_X1 U7314 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n8776) );
  INV_X1 U7315 ( .A(n9931), .ZN(n9677) );
  INV_X1 U7316 ( .A(n9934), .ZN(n9914) );
  OAI21_X1 U7317 ( .B1(n14836), .B2(n7173), .A(n7171), .ZN(n7883) );
  AOI21_X2 U7318 ( .B1(n9078), .B2(n6600), .A(n8743), .ZN(n8744) );
  INV_X2 U7319 ( .A(n12695), .ZN(n13261) );
  INV_X1 U7320 ( .A(n10063), .ZN(n8418) );
  INV_X1 U7321 ( .A(n8891), .ZN(n9283) );
  AND2_X1 U7322 ( .A1(n14323), .A2(n6729), .ZN(n12753) );
  OAI211_X1 U7323 ( .C1(n12919), .C2(n10014), .A(n10016), .B(n10836), .ZN(
        n12997) );
  INV_X1 U7324 ( .A(n8902), .ZN(n12733) );
  AND2_X1 U7325 ( .A1(n10019), .A2(n13176), .ZN(n7421) );
  OAI21_X1 U7326 ( .B1(n7850), .B2(n7849), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6983) );
  AND3_X1 U7327 ( .A1(n8775), .A2(n7836), .A3(n8812), .ZN(n7834) );
  AND2_X1 U7328 ( .A1(n9768), .A2(n9767), .ZN(n15466) );
  INV_X1 U7329 ( .A(n9608), .ZN(n9987) );
  OR2_X1 U7330 ( .A1(n15396), .A2(n15395), .ZN(n7961) );
  XNOR2_X1 U7331 ( .A(n9395), .B(n9420), .ZN(n9984) );
  NAND2_X1 U7333 ( .A1(n7421), .A2(n7422), .ZN(n10023) );
  XNOR2_X1 U7334 ( .A(n6983), .B(n8793), .ZN(n9282) );
  AND2_X1 U7335 ( .A1(n9957), .A2(n9973), .ZN(n9411) );
  NAND2_X1 U7336 ( .A1(n9801), .A2(n9800), .ZN(n15455) );
  XNOR2_X1 U7337 ( .A(n8810), .B(n8809), .ZN(n10983) );
  AOI21_X1 U7338 ( .B1(n7367), .B2(n15959), .A(n7365), .ZN(n7364) );
  OAI21_X1 U7339 ( .B1(n10023), .B2(n15890), .A(n7350), .ZN(n10022) );
  OAI21_X1 U7340 ( .B1(n10023), .B2(n15885), .A(n7423), .ZN(n10024) );
  INV_X1 U7341 ( .A(n15716), .ZN(n15367) );
  INV_X2 U7342 ( .A(n15714), .ZN(n6546) );
  AND4_X2 U7343 ( .A1(n6881), .A2(n6933), .A3(n6931), .A4(n6932), .ZN(n6535)
         );
  AND2_X1 U7345 ( .A1(n15184), .A2(n13067), .ZN(n6536) );
  AND4_X1 U7346 ( .A1(n9548), .A2(n9547), .A3(n9546), .A4(n9545), .ZN(n6537)
         );
  AND4_X1 U7347 ( .A1(n9530), .A2(n9529), .A3(n9528), .A4(n9527), .ZN(n6538)
         );
  INV_X1 U7348 ( .A(n6537), .ZN(n6539) );
  NOR2_X2 U7349 ( .A1(n10026), .A2(n13557), .ZN(n10025) );
  NAND3_X2 U7350 ( .A1(n6612), .A2(n8126), .A3(n8125), .ZN(n15906) );
  XNOR2_X1 U7351 ( .A(n15684), .B(n14954), .ZN(n15671) );
  NAND2_X2 U7352 ( .A1(n11806), .A2(n11807), .ZN(n13239) );
  NOR2_X2 U7353 ( .A1(n15491), .A2(n7989), .ZN(n7987) );
  AND2_X2 U7354 ( .A1(n11790), .A2(n11098), .ZN(n11095) );
  NOR2_X2 U7355 ( .A1(n7541), .A2(n10058), .ZN(n11308) );
  NAND2_X2 U7356 ( .A1(n8475), .A2(n8474), .ZN(n13805) );
  INV_X1 U7357 ( .A(n6538), .ZN(n6540) );
  OR2_X1 U7358 ( .A1(n13476), .A2(n13890), .ZN(n8652) );
  OAI211_X2 U7359 ( .C1(n8442), .C2(n13671), .A(n8380), .B(n8379), .ZN(n13890)
         );
  AOI21_X2 U7360 ( .B1(n15211), .B2(n6638), .A(n7457), .ZN(n15139) );
  OAI211_X2 U7361 ( .C1(n8891), .C2(n7438), .A(n7437), .B(n8907), .ZN(n14243)
         );
  XNOR2_X2 U7362 ( .A(n12775), .B(n6553), .ZN(n12961) );
  INV_X2 U7363 ( .A(n13803), .ZN(n13776) );
  NAND2_X2 U7364 ( .A1(n7262), .A2(n7260), .ZN(n13803) );
  CLKBUF_X1 U7365 ( .A(n12821), .Z(n6541) );
  INV_X1 U7366 ( .A(n12777), .ZN(n12821) );
  NAND2_X1 U7367 ( .A1(n11777), .A2(n15905), .ZN(n13411) );
  INV_X2 U7368 ( .A(n6550), .ZN(n12433) );
  INV_X4 U7369 ( .A(n12413), .ZN(n6549) );
  NAND4_X2 U7370 ( .A1(n8859), .A2(n8858), .A3(n8857), .A4(n8856), .ZN(n14239)
         );
  XNOR2_X2 U7371 ( .A(n8705), .B(SI_5_), .ZN(n8865) );
  AND2_X1 U7372 ( .A1(n9923), .A2(n15733), .ZN(n6543) );
  XNOR2_X2 U7373 ( .A(n13150), .B(n7291), .ZN(n14164) );
  NAND2_X2 U7374 ( .A1(n14078), .A2(n13146), .ZN(n13150) );
  XNOR2_X2 U7375 ( .A(n9077), .B(n9076), .ZN(n10784) );
  NOR2_X2 U7376 ( .A1(n15677), .A2(n15684), .ZN(n11587) );
  NAND2_X2 U7377 ( .A1(n9607), .A2(n9606), .ZN(n15684) );
  NOR3_X2 U7378 ( .A1(n15823), .A2(n15822), .A3(n15827), .ZN(n15824) );
  NAND2_X2 U7379 ( .A1(n9959), .A2(n9411), .ZN(n9477) );
  NAND2_X1 U7382 ( .A1(n9425), .A2(n9426), .ZN(n9509) );
  NAND2_X2 U7383 ( .A1(n7084), .A2(n8253), .ZN(n11391) );
  OAI21_X2 U7384 ( .B1(n9434), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9435) );
  XNOR2_X2 U7385 ( .A(n9423), .B(n9422), .ZN(n9426) );
  AND2_X1 U7386 ( .A1(n7837), .A2(n7839), .ZN(n13203) );
  MUX2_X1 U7387 ( .A(n9378), .B(n9377), .S(n15893), .Z(n9380) );
  NAND2_X1 U7388 ( .A1(n7216), .A2(n7214), .ZN(n15389) );
  NAND2_X1 U7389 ( .A1(n15247), .A2(n13059), .ZN(n15235) );
  OAI21_X2 U7390 ( .B1(n14425), .B2(n7868), .A(n7866), .ZN(n14378) );
  NAND2_X1 U7391 ( .A1(n13057), .A2(n13056), .ZN(n15247) );
  NAND2_X1 U7392 ( .A1(n15280), .A2(n15282), .ZN(n15281) );
  OAI21_X1 U7393 ( .B1(n14595), .B2(n14166), .A(n9193), .ZN(n14379) );
  OAI21_X1 U7394 ( .B1(n14808), .B2(n7187), .A(n7185), .ZN(n7190) );
  AND2_X1 U7395 ( .A1(n6905), .A2(n6720), .ZN(n6904) );
  NAND2_X1 U7396 ( .A1(n12018), .A2(n12644), .ZN(n13010) );
  AND2_X1 U7397 ( .A1(n13048), .A2(n13047), .ZN(n15345) );
  INV_X2 U7398 ( .A(n13790), .ZN(n13338) );
  BUF_X1 U7399 ( .A(n14815), .Z(n7298) );
  NAND4_X1 U7400 ( .A1(n8520), .A2(n8519), .A3(n8518), .A4(n8517), .ZN(n13790)
         );
  NAND2_X1 U7401 ( .A1(n15691), .A2(n15694), .ZN(n15690) );
  OR2_X1 U7402 ( .A1(n8806), .A2(n10928), .ZN(n8808) );
  NAND2_X1 U7403 ( .A1(n11269), .A2(n11268), .ZN(n13354) );
  NAND2_X2 U7404 ( .A1(n12430), .A2(n12435), .ZN(n15708) );
  INV_X1 U7405 ( .A(n14239), .ZN(n12800) );
  NAND2_X2 U7406 ( .A1(n13411), .A2(n13415), .ZN(n11594) );
  NOR2_X1 U7407 ( .A1(n15906), .A2(n11211), .ZN(n15904) );
  NAND4_X1 U7408 ( .A1(n8844), .A2(n8843), .A3(n8842), .A4(n8841), .ZN(n14242)
         );
  NOR2_X2 U7409 ( .A1(n6599), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8377) );
  NAND2_X1 U7410 ( .A1(n15864), .A2(n10843), .ZN(n15843) );
  INV_X1 U7411 ( .A(n9931), .ZN(n9501) );
  INV_X4 U7412 ( .A(n13166), .ZN(n7818) );
  CLKBUF_X2 U7413 ( .A(n9488), .Z(n12583) );
  NAND2_X1 U7414 ( .A1(n9427), .A2(n9426), .ZN(n9990) );
  OR2_X1 U7415 ( .A1(n6603), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n9314) );
  OAI21_X1 U7416 ( .B1(n13688), .B2(n6799), .A(n13667), .ZN(n6798) );
  NAND2_X1 U7417 ( .A1(n7837), .A2(n6637), .ZN(n13201) );
  AOI21_X1 U7418 ( .B1(n6842), .B2(n15763), .A(n15157), .ZN(n15414) );
  NAND2_X1 U7419 ( .A1(n14100), .A2(n14099), .ZN(n14098) );
  AND2_X1 U7420 ( .A1(n7550), .A2(n7549), .ZN(n7548) );
  OR2_X1 U7421 ( .A1(n13689), .A2(n7551), .ZN(n7550) );
  INV_X1 U7422 ( .A(n13689), .ZN(n6547) );
  AND2_X1 U7423 ( .A1(n12692), .A2(n6639), .ZN(n12694) );
  NAND2_X1 U7424 ( .A1(n6536), .A2(n15171), .ZN(n15170) );
  AOI21_X1 U7425 ( .B1(n7683), .B2(n7681), .A(n7680), .ZN(n12701) );
  OR2_X1 U7426 ( .A1(n15148), .A2(n15135), .ZN(n15130) );
  AND2_X1 U7427 ( .A1(n13150), .A2(n13149), .ZN(n14053) );
  OAI21_X1 U7428 ( .B1(n14396), .B2(n7006), .A(n7004), .ZN(n14334) );
  AOI21_X1 U7429 ( .B1(n6834), .B2(n7709), .A(n6610), .ZN(n15186) );
  AOI21_X1 U7430 ( .B1(n7172), .B2(n7175), .A(n7886), .ZN(n7171) );
  NOR2_X1 U7431 ( .A1(n14377), .A2(n9194), .ZN(n14350) );
  AOI211_X1 U7432 ( .C1(n14615), .C2(n10017), .A(n14614), .B(n14613), .ZN(
        n14710) );
  NAND2_X1 U7433 ( .A1(n15235), .A2(n7228), .ZN(n6834) );
  AOI21_X1 U7434 ( .B1(n7005), .B2(n7007), .A(n6656), .ZN(n7004) );
  NAND2_X1 U7435 ( .A1(n15263), .A2(n7951), .ZN(n7949) );
  AOI21_X1 U7436 ( .B1(n14046), .B2(n13119), .A(n13118), .ZN(n14124) );
  XOR2_X1 U7437 ( .A(n14219), .B(n14576), .Z(n14303) );
  INV_X1 U7438 ( .A(n7007), .ZN(n7006) );
  OR2_X1 U7439 ( .A1(n14750), .A2(n14751), .ZN(n7270) );
  NAND2_X1 U7440 ( .A1(n15321), .A2(n13018), .ZN(n15297) );
  AOI22_X1 U7441 ( .A1(n12735), .A2(n12734), .B1(n12733), .B2(
        P1_DATAO_REG_31__SCAN_IN), .ZN(n14570) );
  OR2_X1 U7442 ( .A1(n15218), .A2(n15428), .ZN(n15203) );
  AOI211_X1 U7443 ( .C1(n14615), .C2(n14444), .A(n14635), .B(n14443), .ZN(
        n14614) );
  OR2_X1 U7444 ( .A1(n14075), .A2(n13140), .ZN(n13142) );
  NAND2_X1 U7445 ( .A1(n14139), .A2(n13138), .ZN(n7347) );
  AND2_X1 U7446 ( .A1(n7707), .A2(n15201), .ZN(n7709) );
  INV_X1 U7447 ( .A(n7190), .ZN(n14750) );
  NAND2_X1 U7448 ( .A1(n8453), .A2(n8452), .ZN(n13923) );
  OR2_X1 U7449 ( .A1(n14181), .A2(n13135), .ZN(n14138) );
  NAND2_X1 U7450 ( .A1(n7117), .A2(n7114), .ZN(n14477) );
  OAI21_X1 U7451 ( .B1(n13342), .B2(n12673), .A(n7326), .ZN(n13288) );
  NAND2_X1 U7452 ( .A1(n9666), .A2(n9665), .ZN(n14893) );
  OR2_X1 U7453 ( .A1(n13831), .A2(n13849), .ZN(n13487) );
  NAND2_X1 U7454 ( .A1(n13010), .A2(n13009), .ZN(n15369) );
  NAND2_X1 U7455 ( .A1(n9822), .A2(n9821), .ZN(n15443) );
  NAND2_X1 U7456 ( .A1(n13012), .A2(n13011), .ZN(n15320) );
  NAND2_X1 U7457 ( .A1(n8436), .A2(n8435), .ZN(n13831) );
  INV_X1 U7458 ( .A(n13012), .ZN(n15334) );
  NAND2_X1 U7459 ( .A1(n9185), .A2(n9184), .ZN(n14595) );
  NAND2_X1 U7460 ( .A1(n9399), .A2(n9398), .ZN(n15447) );
  NAND2_X1 U7461 ( .A1(n7985), .A2(n7988), .ZN(n15346) );
  NAND2_X1 U7462 ( .A1(n9142), .A2(n9141), .ZN(n14610) );
  NAND2_X1 U7463 ( .A1(n9171), .A2(n9170), .ZN(n14600) );
  AND2_X1 U7464 ( .A1(n15244), .A2(n12529), .ZN(n15282) );
  XNOR2_X1 U7465 ( .A(n9155), .B(n9154), .ZN(n11109) );
  XNOR2_X1 U7466 ( .A(n9183), .B(n9182), .ZN(n11458) );
  AOI21_X1 U7467 ( .B1(n11901), .B2(n11900), .A(n11899), .ZN(n11908) );
  INV_X1 U7468 ( .A(n15345), .ZN(n15341) );
  OR2_X1 U7469 ( .A1(n12482), .A2(n12483), .ZN(n12484) );
  NAND2_X1 U7470 ( .A1(n7572), .A2(n9151), .ZN(n9155) );
  NAND2_X1 U7471 ( .A1(n9733), .A2(n9732), .ZN(n15479) );
  NAND2_X1 U7472 ( .A1(n7609), .A2(n8434), .ZN(n8461) );
  NAND2_X1 U7473 ( .A1(n9083), .A2(n9082), .ZN(n14500) );
  NAND2_X1 U7474 ( .A1(n7210), .A2(n8402), .ZN(n8433) );
  AND2_X1 U7475 ( .A1(n9689), .A2(n9688), .ZN(n14815) );
  NAND2_X1 U7476 ( .A1(n8357), .A2(n8356), .ZN(n13465) );
  NAND2_X1 U7477 ( .A1(n9009), .A2(n9008), .ZN(n14658) );
  NAND2_X1 U7478 ( .A1(n7490), .A2(n7491), .ZN(n9166) );
  NAND2_X1 U7479 ( .A1(n8390), .A2(n8389), .ZN(n14017) );
  NAND2_X1 U7480 ( .A1(n9670), .A2(n9669), .ZN(n14891) );
  NAND2_X1 U7481 ( .A1(n6928), .A2(n11317), .ZN(n10146) );
  XNOR2_X1 U7482 ( .A(n9093), .B(n9092), .ZN(n10708) );
  NAND2_X1 U7483 ( .A1(n6796), .A2(n8752), .ZN(n8806) );
  OAI21_X1 U7484 ( .B1(n7342), .B2(n9056), .A(n9057), .ZN(n9075) );
  NAND2_X1 U7485 ( .A1(n6879), .A2(n9645), .ZN(n12475) );
  AND2_X1 U7486 ( .A1(n13407), .A2(n13454), .ZN(n13453) );
  AND2_X1 U7487 ( .A1(n13440), .A2(n13439), .ZN(n13539) );
  AND2_X1 U7488 ( .A1(n6926), .A2(n11145), .ZN(n10056) );
  NOR2_X1 U7489 ( .A1(n6926), .A2(n11145), .ZN(n6925) );
  NOR2_X1 U7490 ( .A1(n15973), .A2(n15948), .ZN(n13942) );
  NAND2_X1 U7491 ( .A1(n6832), .A2(n8716), .ZN(n8719) );
  NOR2_X1 U7492 ( .A1(n7476), .A2(n7474), .ZN(n7473) );
  OAI21_X1 U7493 ( .B1(n6832), .B2(n7104), .A(n7102), .ZN(n7105) );
  INV_X1 U7494 ( .A(n15880), .ZN(n12799) );
  NAND2_X1 U7495 ( .A1(n8954), .A2(n8713), .ZN(n7056) );
  NAND4_X1 U7496 ( .A1(n8104), .A2(n8832), .A3(n8831), .A4(n8830), .ZN(n14241)
         );
  XNOR2_X1 U7497 ( .A(n8921), .B(n8922), .ZN(n10220) );
  NOR2_X2 U7498 ( .A1(n6982), .A2(n6981), .ZN(n11326) );
  NAND2_X1 U7499 ( .A1(n6698), .A2(n8850), .ZN(n12784) );
  NAND2_X1 U7500 ( .A1(n6917), .A2(n7277), .ZN(n11777) );
  INV_X2 U7501 ( .A(n8889), .ZN(n12737) );
  NAND4_X1 U7502 ( .A1(n8171), .A2(n8170), .A3(n8169), .A4(n8168), .ZN(n13589)
         );
  NAND4_X1 U7503 ( .A1(n8159), .A2(n8158), .A3(n8157), .A4(n8156), .ZN(n13590)
         );
  OAI21_X1 U7504 ( .B1(n15732), .B2(n9954), .A(n9463), .ZN(n9464) );
  NAND2_X1 U7505 ( .A1(n8798), .A2(n8799), .ZN(n8889) );
  INV_X2 U7506 ( .A(n9169), .ZN(n12734) );
  NAND2_X1 U7507 ( .A1(n6701), .A2(n6565), .ZN(n7503) );
  OAI211_X2 U7508 ( .C1(n8176), .C2(SI_2_), .A(n7777), .B(n7776), .ZN(n13965)
         );
  INV_X1 U7509 ( .A(n10842), .ZN(n10843) );
  AND4_X1 U7510 ( .A1(n9569), .A2(n9568), .A3(n9567), .A4(n9566), .ZN(n12418)
         );
  OAI211_X1 U7511 ( .C1(n13372), .C2(n10519), .A(n7385), .B(n7384), .ZN(n11778) );
  INV_X2 U7512 ( .A(n13372), .ZN(n13369) );
  NAND4_X1 U7513 ( .A1(n9493), .A2(n9492), .A3(n9491), .A4(n9490), .ZN(n15638)
         );
  NAND2_X1 U7514 ( .A1(n13084), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8797) );
  XNOR2_X1 U7515 ( .A(n8710), .B(SI_7_), .ZN(n8936) );
  AOI21_X1 U7516 ( .B1(n8708), .B2(n7396), .A(n6673), .ZN(n7100) );
  INV_X1 U7517 ( .A(n8122), .ZN(n14036) );
  OR2_X2 U7518 ( .A1(n11066), .A2(n12622), .ZN(n15733) );
  INV_X1 U7519 ( .A(n11064), .ZN(n12438) );
  NAND2_X2 U7520 ( .A1(n12767), .A2(n10856), .ZN(n13166) );
  NAND4_X1 U7521 ( .A1(n9471), .A2(n9470), .A3(n9469), .A4(n9468), .ZN(n14958)
         );
  NAND2_X2 U7522 ( .A1(n10063), .A2(n8129), .ZN(n13372) );
  NAND2_X2 U7523 ( .A1(n10063), .A2(n10481), .ZN(n8176) );
  CLKBUF_X2 U7524 ( .A(n9608), .Z(n9927) );
  NAND2_X2 U7525 ( .A1(n13570), .A2(n8665), .ZN(n13514) );
  BUF_X2 U7526 ( .A(n12584), .Z(n12579) );
  CLKBUF_X1 U7527 ( .A(n9494), .Z(n12615) );
  AND2_X1 U7528 ( .A1(n8707), .A2(n8919), .ZN(n8708) );
  NAND2_X1 U7529 ( .A1(n8588), .A2(n8587), .ZN(n12123) );
  AND2_X1 U7530 ( .A1(n8120), .A2(n8119), .ZN(n8122) );
  INV_X2 U7531 ( .A(n9779), .ZN(n12614) );
  NAND2_X1 U7532 ( .A1(n8781), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6984) );
  AND2_X1 U7533 ( .A1(n9410), .A2(n9409), .ZN(n9959) );
  BUF_X2 U7534 ( .A(n15553), .Z(n6809) );
  XNOR2_X1 U7535 ( .A(n9273), .B(n9329), .ZN(n12409) );
  NAND2_X2 U7536 ( .A1(n8136), .A2(n8135), .ZN(n13717) );
  XNOR2_X1 U7537 ( .A(n8818), .B(n8817), .ZN(n12987) );
  INV_X2 U7538 ( .A(n15550), .ZN(n10985) );
  NAND2_X1 U7539 ( .A1(n7841), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9273) );
  NAND2_X1 U7540 ( .A1(n8135), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8133) );
  XNOR2_X1 U7541 ( .A(n8620), .B(n8619), .ZN(n11213) );
  CLKBUF_X1 U7543 ( .A(n15649), .Z(n7374) );
  XNOR2_X1 U7544 ( .A(n8404), .B(n7302), .ZN(n13745) );
  NAND2_X1 U7545 ( .A1(n6711), .A2(n6882), .ZN(n8135) );
  MUX2_X1 U7546 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8134), .S(
        P3_IR_REG_27__SCAN_IN), .Z(n8136) );
  XNOR2_X1 U7547 ( .A(n9438), .B(P1_IR_REG_19__SCAN_IN), .ZN(n15112) );
  NAND2_X1 U7548 ( .A1(n9314), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7148) );
  NOR2_X1 U7549 ( .A1(n8387), .A2(n8578), .ZN(n8584) );
  AND2_X1 U7550 ( .A1(n8814), .A2(n6633), .ZN(n9323) );
  NAND2_X1 U7551 ( .A1(n8119), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8116) );
  NAND2_X1 U7552 ( .A1(n7227), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9423) );
  XNOR2_X1 U7553 ( .A(n7571), .B(n8189), .ZN(n11697) );
  NAND2_X1 U7554 ( .A1(n6535), .A2(n8106), .ZN(n8387) );
  AND2_X1 U7555 ( .A1(n6633), .A2(n8816), .ZN(n7840) );
  AND2_X1 U7556 ( .A1(n8000), .A2(n7879), .ZN(n9414) );
  XNOR2_X1 U7557 ( .A(n6921), .B(n10321), .ZN(n10523) );
  NAND3_X1 U7558 ( .A1(n8833), .A2(n7834), .A3(n7833), .ZN(n9303) );
  AND3_X1 U7559 ( .A1(n8113), .A2(n7313), .A3(n6733), .ZN(n6918) );
  INV_X1 U7560 ( .A(n8276), .ZN(n8106) );
  AND2_X1 U7561 ( .A1(n9550), .A2(n7761), .ZN(n7760) );
  NAND2_X1 U7562 ( .A1(n8898), .A2(n8897), .ZN(n14250) );
  AND2_X2 U7563 ( .A1(n9388), .A2(n9456), .ZN(n9550) );
  AND2_X1 U7564 ( .A1(n8774), .A2(n8776), .ZN(n7833) );
  AND4_X1 U7565 ( .A1(n8112), .A2(n8111), .A3(n8110), .A4(n8109), .ZN(n8113)
         );
  AND2_X2 U7566 ( .A1(n8847), .A2(n7051), .ZN(n8833) );
  NOR2_X2 U7567 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9456) );
  INV_X1 U7568 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8304) );
  NOR2_X1 U7569 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n9388) );
  NOR2_X1 U7570 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n9381) );
  NOR2_X1 U7571 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n9382) );
  INV_X4 U7572 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X4 U7573 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7574 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n8115) );
  NOR2_X1 U7575 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n6932) );
  INV_X1 U7576 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9643) );
  INV_X1 U7577 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n7836) );
  NOR2_X1 U7578 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), .ZN(
        n8108) );
  NOR2_X1 U7579 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n9384) );
  INV_X4 U7580 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X1 U7581 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8181) );
  NOR2_X2 U7582 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n8151) );
  NOR2_X1 U7583 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n9406) );
  NAND2_X1 U7584 ( .A1(n9414), .A2(n9401), .ZN(n9409) );
  NOR2_X2 U7585 ( .A1(n14558), .A2(n14653), .ZN(n6791) );
  AND2_X1 U7586 ( .A1(n12997), .A2(n10018), .ZN(n10019) );
  INV_X1 U7587 ( .A(n6549), .ZN(n6550) );
  INV_X1 U7588 ( .A(n6549), .ZN(n6551) );
  NAND2_X2 U7589 ( .A1(n9475), .A2(n8129), .ZN(n9779) );
  OAI211_X1 U7590 ( .C1(n10626), .C2(n14250), .A(n8904), .B(n8903), .ZN(n12778) );
  NOR2_X1 U7591 ( .A1(n9291), .A2(n9290), .ZN(n6554) );
  INV_X4 U7592 ( .A(n12806), .ZN(n12777) );
  OR2_X1 U7593 ( .A1(n12778), .A2(n11158), .ZN(n11706) );
  AND2_X4 U7594 ( .A1(n8121), .A2(n8122), .ZN(n8199) );
  OAI21_X1 U7595 ( .B1(n7062), .B2(n9193), .A(n6690), .ZN(n7414) );
  MUX2_X1 U7596 ( .A(n14873), .B(n14815), .S(n12624), .Z(n12492) );
  AND2_X1 U7597 ( .A1(n7972), .A2(n8733), .ZN(n7971) );
  NAND2_X1 U7598 ( .A1(n8729), .A2(n7973), .ZN(n7972) );
  NAND2_X1 U7599 ( .A1(n8719), .A2(n7574), .ZN(n7970) );
  NOR2_X1 U7600 ( .A1(n7974), .A2(n7104), .ZN(n7574) );
  INV_X1 U7601 ( .A(n8729), .ZN(n7974) );
  NAND4_X1 U7602 ( .A1(n8108), .A2(n8107), .A3(n8304), .A4(n10272), .ZN(n8386)
         );
  NOR2_X1 U7603 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), .ZN(
        n8107) );
  NAND2_X1 U7604 ( .A1(n8151), .A2(n8251), .ZN(n8276) );
  XNOR2_X1 U7605 ( .A(n11326), .B(n13166), .ZN(n11039) );
  INV_X1 U7606 ( .A(n8931), .ZN(n9266) );
  INV_X1 U7607 ( .A(n9053), .ZN(n7845) );
  XNOR2_X1 U7608 ( .A(n12627), .B(n15118), .ZN(n12653) );
  NOR2_X1 U7609 ( .A1(n15425), .A2(n14939), .ZN(n7980) );
  NAND2_X1 U7610 ( .A1(n6831), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9890) );
  NAND2_X1 U7611 ( .A1(n7165), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9395) );
  NAND2_X1 U7612 ( .A1(n9205), .A2(n8765), .ZN(n9210) );
  AND2_X1 U7613 ( .A1(n9550), .A2(n9405), .ZN(n7879) );
  NAND2_X1 U7614 ( .A1(n11844), .A2(n7926), .ZN(n7290) );
  INV_X1 U7615 ( .A(n11848), .ZN(n7926) );
  NAND2_X1 U7616 ( .A1(n14027), .A2(n13561), .ZN(n11599) );
  OR2_X1 U7617 ( .A1(n13348), .A2(n12672), .ZN(n7326) );
  OAI21_X1 U7618 ( .B1(n7414), .B2(n7411), .A(n7412), .ZN(n14335) );
  AOI21_X1 U7619 ( .B1(n7415), .B2(n7062), .A(n7413), .ZN(n7412) );
  INV_X1 U7620 ( .A(n14337), .ZN(n7413) );
  XNOR2_X1 U7621 ( .A(n15150), .B(n14914), .ZN(n15141) );
  NAND2_X1 U7622 ( .A1(n15139), .A2(n15141), .ZN(n7301) );
  NAND2_X1 U7623 ( .A1(n7954), .A2(n7953), .ZN(n15212) );
  OR2_X1 U7624 ( .A1(n15443), .A2(n14942), .ZN(n7953) );
  NAND2_X1 U7625 ( .A1(n7949), .A2(n7948), .ZN(n7954) );
  AND2_X1 U7626 ( .A1(n7950), .A2(n15227), .ZN(n7948) );
  OAI21_X1 U7627 ( .B1(n15597), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n15596), .ZN(
        n15605) );
  INV_X1 U7628 ( .A(n12492), .ZN(n7726) );
  INV_X1 U7629 ( .A(n12488), .ZN(n7728) );
  INV_X1 U7630 ( .A(n12489), .ZN(n7722) );
  INV_X1 U7631 ( .A(n12811), .ZN(n7136) );
  AND2_X1 U7632 ( .A1(n12494), .A2(n15345), .ZN(n7724) );
  AND2_X1 U7633 ( .A1(n13533), .A2(n8018), .ZN(n8017) );
  NAND2_X1 U7634 ( .A1(n7162), .A2(n12890), .ZN(n12894) );
  NAND2_X1 U7635 ( .A1(n12891), .A2(n8060), .ZN(n8059) );
  INV_X1 U7636 ( .A(n12893), .ZN(n8060) );
  NAND2_X1 U7637 ( .A1(n13490), .A2(n8004), .ZN(n8011) );
  NAND2_X1 U7638 ( .A1(n6808), .A2(n6807), .ZN(n12557) );
  INV_X1 U7639 ( .A(n12555), .ZN(n6807) );
  INV_X1 U7640 ( .A(n12556), .ZN(n6808) );
  NAND2_X1 U7641 ( .A1(n6702), .A2(n13478), .ZN(n7811) );
  NAND2_X1 U7642 ( .A1(n12386), .A2(n13474), .ZN(n7814) );
  INV_X1 U7643 ( .A(n8273), .ZN(n7602) );
  INV_X1 U7644 ( .A(n7601), .ZN(n7600) );
  OAI21_X1 U7645 ( .B1(n8271), .B2(n7602), .A(n8287), .ZN(n7601) );
  OAI21_X1 U7646 ( .B1(n10537), .B2(n6681), .A(n7248), .ZN(n7287) );
  NAND2_X1 U7647 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(n7249), .ZN(n7248) );
  INV_X1 U7648 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7249) );
  NAND2_X1 U7649 ( .A1(n7570), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7569) );
  NAND2_X1 U7650 ( .A1(n11687), .A2(n10053), .ZN(n10054) );
  NAND2_X1 U7651 ( .A1(n7097), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7093) );
  AOI21_X1 U7652 ( .B1(n7409), .B2(n7408), .A(n6674), .ZN(n7407) );
  NAND3_X1 U7653 ( .A1(n7409), .A2(n6920), .A3(n7672), .ZN(n7406) );
  OR2_X1 U7654 ( .A1(n13912), .A2(n13776), .ZN(n13501) );
  NAND2_X1 U7655 ( .A1(n6908), .A2(n6906), .ZN(n6903) );
  AND2_X1 U7656 ( .A1(n6907), .A2(n8651), .ZN(n6906) );
  OR3_X1 U7657 ( .A1(n11128), .A2(n13735), .A3(n11213), .ZN(n8630) );
  OR2_X1 U7658 ( .A1(n13990), .A2(n13826), .ZN(n13495) );
  NAND2_X1 U7659 ( .A1(n6909), .A2(n7386), .ZN(n13833) );
  AOI21_X1 U7660 ( .B1(n8662), .B2(n7387), .A(n6661), .ZN(n7386) );
  NAND2_X1 U7661 ( .A1(n6904), .A2(n6903), .ZN(n6909) );
  INV_X1 U7662 ( .A(n8661), .ZN(n7387) );
  NOR2_X1 U7663 ( .A1(P3_IR_REG_26__SCAN_IN), .A2(P3_IR_REG_25__SCAN_IN), .ZN(
        n8105) );
  NAND2_X1 U7664 ( .A1(n8114), .A2(n8113), .ZN(n8578) );
  AND2_X1 U7665 ( .A1(n7944), .A2(n7943), .ZN(n7942) );
  NOR2_X1 U7666 ( .A1(n7039), .A2(P3_IR_REG_19__SCAN_IN), .ZN(n7038) );
  NOR2_X1 U7667 ( .A1(n8276), .A2(n8386), .ZN(n7941) );
  INV_X1 U7668 ( .A(n8319), .ZN(n7226) );
  NAND2_X1 U7669 ( .A1(n14570), .A2(n12953), .ZN(n8050) );
  NAND2_X1 U7670 ( .A1(n14420), .A2(n14225), .ZN(n7876) );
  AND2_X1 U7671 ( .A1(n9052), .A2(n6709), .ZN(n7848) );
  NAND2_X1 U7672 ( .A1(n11109), .A2(n12734), .ZN(n7587) );
  INV_X1 U7673 ( .A(n14226), .ZN(n9361) );
  INV_X1 U7674 ( .A(n7439), .ZN(n7001) );
  NAND2_X1 U7675 ( .A1(n14454), .A2(n9359), .ZN(n7441) );
  OR2_X1 U7676 ( .A1(n14615), .A2(n14227), .ZN(n12978) );
  NOR2_X1 U7677 ( .A1(n6578), .A2(n9357), .ZN(n7744) );
  INV_X1 U7678 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8793) );
  INV_X1 U7679 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8771) );
  NOR2_X1 U7680 ( .A1(n6563), .A2(n14743), .ZN(n7906) );
  INV_X1 U7681 ( .A(n9427), .ZN(n9425) );
  NAND2_X1 U7682 ( .A1(n7540), .A2(n7539), .ZN(n15046) );
  NAND2_X1 U7683 ( .A1(n15044), .A2(n15043), .ZN(n7539) );
  OR2_X1 U7684 ( .A1(n9944), .A2(n9943), .ZN(n9985) );
  INV_X1 U7685 ( .A(n13068), .ZN(n7691) );
  NAND2_X1 U7686 ( .A1(n7194), .A2(n13050), .ZN(n7193) );
  INV_X1 U7687 ( .A(n13046), .ZN(n7194) );
  INV_X1 U7688 ( .A(n14946), .ZN(n14831) );
  NAND2_X1 U7689 ( .A1(n14815), .A2(n12486), .ZN(n7989) );
  OR2_X1 U7690 ( .A1(n15638), .A2(n15743), .ZN(n12426) );
  OR2_X1 U7691 ( .A1(n13013), .A2(n15370), .ZN(n13017) );
  OR2_X1 U7692 ( .A1(n13014), .A2(n15317), .ZN(n13013) );
  NAND2_X1 U7693 ( .A1(n15553), .A2(n15112), .ZN(n12412) );
  INV_X1 U7694 ( .A(n12590), .ZN(n7489) );
  INV_X1 U7695 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9389) );
  NOR2_X1 U7696 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n9390) );
  AOI21_X1 U7697 ( .B1(n9209), .B2(n7511), .A(n6763), .ZN(n7510) );
  NAND2_X1 U7698 ( .A1(n7499), .A2(n7500), .ZN(n9151) );
  AND2_X1 U7699 ( .A1(n9079), .A2(n10781), .ZN(n9057) );
  NAND2_X1 U7700 ( .A1(n13288), .A2(n12674), .ZN(n7036) );
  INV_X1 U7701 ( .A(n7930), .ZN(n7929) );
  AOI22_X1 U7702 ( .A1(n11843), .A2(n11842), .B1(n11841), .B2(n13585), .ZN(
        n11844) );
  NAND2_X1 U7703 ( .A1(n11781), .A2(n11780), .ZN(n11782) );
  AND3_X1 U7704 ( .A1(n13558), .A2(n7231), .A3(n7230), .ZN(n13560) );
  NOR2_X1 U7705 ( .A1(n13556), .A2(n7312), .ZN(n7231) );
  INV_X1 U7706 ( .A(n11128), .ZN(n13570) );
  INV_X1 U7707 ( .A(n13377), .ZN(n8667) );
  INV_X1 U7708 ( .A(n13376), .ZN(n8668) );
  INV_X1 U7709 ( .A(n8199), .ZN(n8442) );
  OR2_X1 U7710 ( .A1(n10052), .A2(n10523), .ZN(n7570) );
  NAND2_X1 U7711 ( .A1(n11682), .A2(n7095), .ZN(n7097) );
  NOR2_X1 U7712 ( .A1(n10530), .A2(n7096), .ZN(n7095) );
  INV_X1 U7713 ( .A(n10072), .ZN(n7096) );
  OR2_X1 U7714 ( .A1(n10054), .A2(n10530), .ZN(n7557) );
  NAND3_X1 U7715 ( .A1(n13633), .A2(n10134), .A3(n10135), .ZN(n13649) );
  XNOR2_X1 U7716 ( .A(n13676), .B(n7380), .ZN(n13651) );
  NAND2_X1 U7717 ( .A1(n11925), .A2(n8248), .ZN(n13442) );
  AND2_X1 U7718 ( .A1(n13443), .A2(n13442), .ZN(n13538) );
  INV_X1 U7719 ( .A(n13585), .ZN(n11925) );
  INV_X1 U7720 ( .A(n13745), .ZN(n13735) );
  NOR2_X1 U7721 ( .A1(n11271), .A2(n15948), .ZN(n11275) );
  AOI21_X1 U7722 ( .B1(n10041), .B2(n13557), .A(n6884), .ZN(n13362) );
  INV_X1 U7723 ( .A(n13523), .ZN(n6884) );
  NOR2_X1 U7724 ( .A1(n13824), .A2(n7420), .ZN(n7419) );
  OR2_X1 U7725 ( .A1(n13514), .A2(n8673), .ZN(n15914) );
  INV_X1 U7726 ( .A(n15914), .ZN(n13889) );
  INV_X1 U7727 ( .A(n11271), .ZN(n13567) );
  INV_X1 U7728 ( .A(n8386), .ZN(n8114) );
  AND2_X1 U7729 ( .A1(n8105), .A2(n8030), .ZN(n7313) );
  INV_X1 U7730 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8030) );
  NAND2_X1 U7731 ( .A1(n7229), .A2(n7613), .ZN(n8563) );
  AOI21_X1 U7732 ( .B1(n7615), .B2(n7614), .A(n6781), .ZN(n7613) );
  OR2_X1 U7733 ( .A1(n8523), .A2(n7616), .ZN(n7229) );
  AOI21_X1 U7734 ( .B1(n7620), .B2(n8522), .A(n6782), .ZN(n7619) );
  AND2_X1 U7735 ( .A1(n7209), .A2(n7607), .ZN(n7208) );
  AOI21_X1 U7736 ( .B1(n7610), .B2(n7612), .A(n7608), .ZN(n7607) );
  INV_X1 U7737 ( .A(n11227), .ZN(n7828) );
  NAND2_X1 U7738 ( .A1(n8789), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9113) );
  INV_X1 U7739 ( .A(n9099), .ZN(n8789) );
  INV_X1 U7740 ( .A(n14508), .ZN(n13148) );
  NOR2_X1 U7741 ( .A1(n10838), .A2(n10837), .ZN(n10847) );
  AND2_X1 U7742 ( .A1(n9224), .A2(n9223), .ZN(n14101) );
  AND2_X1 U7743 ( .A1(n9192), .A2(n9191), .ZN(n14166) );
  AND2_X1 U7744 ( .A1(n9164), .A2(n9163), .ZN(n14165) );
  AND2_X1 U7745 ( .A1(n9135), .A2(n9134), .ZN(n12884) );
  AND3_X1 U7746 ( .A1(n9091), .A2(n9090), .A3(n9089), .ZN(n14116) );
  INV_X1 U7747 ( .A(n8798), .ZN(n6986) );
  NAND2_X1 U7748 ( .A1(n7044), .A2(n7043), .ZN(n12337) );
  AOI21_X1 U7749 ( .B1(n7045), .B2(n7047), .A(n6780), .ZN(n7043) );
  NAND2_X1 U7750 ( .A1(n7063), .A2(n7466), .ZN(n9205) );
  INV_X1 U7751 ( .A(n9202), .ZN(n7064) );
  INV_X1 U7752 ( .A(n7869), .ZN(n7868) );
  AOI21_X1 U7753 ( .B1(n7869), .B2(n7867), .A(n6676), .ZN(n7866) );
  NOR2_X1 U7754 ( .A1(n14398), .A2(n7870), .ZN(n7869) );
  NAND2_X1 U7755 ( .A1(n14425), .A2(n7874), .ZN(n7871) );
  INV_X1 U7756 ( .A(n7441), .ZN(n7440) );
  INV_X1 U7757 ( .A(n9051), .ZN(n9050) );
  NOR2_X2 U7758 ( .A1(n11557), .A2(n12799), .ZN(n11790) );
  BUF_X1 U7759 ( .A(n10626), .Z(n7327) );
  OAI21_X1 U7760 ( .B1(n14318), .B2(n7576), .A(n7580), .ZN(n10020) );
  INV_X1 U7761 ( .A(n7575), .ZN(n7580) );
  OAI21_X1 U7762 ( .B1(n7582), .B2(n7576), .A(n12983), .ZN(n7575) );
  NAND2_X1 U7763 ( .A1(n14391), .A2(n9363), .ZN(n14396) );
  AND2_X1 U7764 ( .A1(n9311), .A2(n9317), .ZN(n15852) );
  INV_X1 U7765 ( .A(n8833), .ZN(n8860) );
  NAND2_X1 U7766 ( .A1(n7880), .A2(n6646), .ZN(n7169) );
  OAI21_X1 U7767 ( .B1(n15743), .B2(n9954), .A(n9499), .ZN(n9500) );
  AND2_X1 U7768 ( .A1(n7884), .A2(n7882), .ZN(n7881) );
  NAND2_X1 U7769 ( .A1(n9832), .A2(n6564), .ZN(n7882) );
  NAND2_X1 U7771 ( .A1(n9425), .A2(n9424), .ZN(n9594) );
  NAND2_X1 U7772 ( .A1(n9427), .A2(n9424), .ZN(n9608) );
  AND2_X1 U7773 ( .A1(n7526), .A2(n10575), .ZN(n7514) );
  INV_X1 U7774 ( .A(n14993), .ZN(n7526) );
  OR2_X1 U7775 ( .A1(n7522), .A2(n14993), .ZN(n7521) );
  AOI21_X1 U7776 ( .B1(n10575), .B2(n14978), .A(n7523), .ZN(n7522) );
  INV_X1 U7777 ( .A(n14994), .ZN(n7523) );
  NAND2_X1 U7778 ( .A1(n12617), .A2(n12616), .ZN(n12627) );
  NAND2_X1 U7779 ( .A1(n15170), .A2(n7690), .ZN(n7219) );
  NOR2_X1 U7780 ( .A1(n15141), .A2(n7218), .ZN(n7217) );
  INV_X1 U7781 ( .A(n13070), .ZN(n7218) );
  AOI21_X1 U7782 ( .B1(n7979), .B2(n7976), .A(n6666), .ZN(n7975) );
  INV_X1 U7783 ( .A(n7982), .ZN(n7976) );
  AND2_X1 U7784 ( .A1(n9891), .A2(n6615), .ZN(n15174) );
  NAND2_X1 U7785 ( .A1(n15199), .A2(n7982), .ZN(n7981) );
  AOI21_X1 U7786 ( .B1(n7951), .B2(n15266), .A(n6663), .ZN(n7950) );
  OR2_X1 U7787 ( .A1(n15455), .A2(n14944), .ZN(n7956) );
  OR2_X1 U7788 ( .A1(n15263), .A2(n15266), .ZN(n7957) );
  NOR2_X1 U7789 ( .A1(n8089), .A2(n6647), .ZN(n7451) );
  INV_X1 U7790 ( .A(n9494), .ZN(n9799) );
  INV_X1 U7791 ( .A(n9475), .ZN(n9798) );
  NAND2_X1 U7792 ( .A1(n9475), .A2(n10481), .ZN(n9494) );
  NAND2_X2 U7793 ( .A1(n9984), .A2(n15649), .ZN(n9475) );
  NOR2_X1 U7794 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n9386) );
  XNOR2_X1 U7795 ( .A(n9976), .B(P1_IR_REG_23__SCAN_IN), .ZN(n10187) );
  XNOR2_X1 U7796 ( .A(n9415), .B(P1_IR_REG_20__SCAN_IN), .ZN(n12622) );
  OR2_X1 U7797 ( .A1(n9414), .A2(n9394), .ZN(n9415) );
  NAND3_X1 U7798 ( .A1(n7946), .A2(n8695), .A3(SI_1_), .ZN(n7945) );
  INV_X1 U7799 ( .A(n9456), .ZN(n9496) );
  AOI21_X1 U7800 ( .B1(n15978), .B2(n15977), .A(n10567), .ZN(n10569) );
  NAND2_X1 U7801 ( .A1(n10942), .A2(n10941), .ZN(n10951) );
  XNOR2_X1 U7802 ( .A(n11717), .B(n10960), .ZN(n10961) );
  NAND2_X1 U7803 ( .A1(n9213), .A2(n9212), .ZN(n14327) );
  NAND2_X1 U7804 ( .A1(n9286), .A2(n9287), .ZN(n7061) );
  NAND2_X1 U7805 ( .A1(n14682), .A2(n15893), .ZN(n7110) );
  NAND2_X1 U7806 ( .A1(n6659), .A2(n7301), .ZN(n15404) );
  NAND2_X1 U7807 ( .A1(n12134), .A2(n12133), .ZN(n12271) );
  INV_X1 U7808 ( .A(n7637), .ZN(n7266) );
  NAND2_X1 U7809 ( .A1(n15613), .A2(n7640), .ZN(n7638) );
  INV_X1 U7810 ( .A(n7639), .ZN(n7636) );
  INV_X1 U7811 ( .A(n12802), .ZN(n8081) );
  INV_X1 U7812 ( .A(n12801), .ZN(n8083) );
  NOR2_X1 U7813 ( .A1(n8083), .A2(n8081), .ZN(n8080) );
  AND2_X1 U7814 ( .A1(n8082), .A2(n8079), .ZN(n8077) );
  NAND2_X1 U7815 ( .A1(n8083), .A2(n8081), .ZN(n8079) );
  NAND2_X1 U7816 ( .A1(n8077), .A2(n8080), .ZN(n8075) );
  AOI21_X1 U7817 ( .B1(n8080), .B2(n8079), .A(n8082), .ZN(n8078) );
  NAND2_X1 U7818 ( .A1(n8072), .A2(n8071), .ZN(n8070) );
  NAND2_X1 U7819 ( .A1(n12804), .A2(n8079), .ZN(n8071) );
  INV_X1 U7820 ( .A(n8077), .ZN(n8072) );
  NAND2_X1 U7821 ( .A1(n7727), .A2(n7726), .ZN(n7725) );
  NAND2_X1 U7822 ( .A1(n7721), .A2(n7720), .ZN(n7719) );
  INV_X1 U7823 ( .A(n12491), .ZN(n7727) );
  AOI21_X1 U7824 ( .B1(n12813), .B2(n12814), .A(n8035), .ZN(n8034) );
  INV_X1 U7825 ( .A(n12812), .ZN(n8035) );
  NOR2_X1 U7826 ( .A1(n12813), .A2(n12814), .ZN(n8033) );
  AND2_X1 U7827 ( .A1(n8015), .A2(n8022), .ZN(n8014) );
  NAND2_X1 U7828 ( .A1(n6694), .A2(n13519), .ZN(n8022) );
  NAND2_X1 U7829 ( .A1(n8017), .A2(n6583), .ZN(n8015) );
  OAI21_X1 U7830 ( .B1(n13417), .B2(n6942), .A(n6649), .ZN(n6941) );
  NAND2_X1 U7831 ( .A1(n6916), .A2(n6943), .ZN(n6942) );
  NAND2_X1 U7832 ( .A1(n12883), .A2(n6800), .ZN(n8065) );
  AND2_X1 U7833 ( .A1(n12882), .A2(n8067), .ZN(n6800) );
  NOR2_X1 U7834 ( .A1(n12886), .A2(n12885), .ZN(n8066) );
  NAND2_X1 U7835 ( .A1(n7752), .A2(n12542), .ZN(n7756) );
  INV_X1 U7836 ( .A(n12896), .ZN(n7339) );
  NAND2_X1 U7837 ( .A1(n8058), .A2(n12896), .ZN(n8057) );
  NAND2_X1 U7838 ( .A1(n8061), .A2(n8059), .ZN(n8058) );
  INV_X1 U7839 ( .A(n12895), .ZN(n6792) );
  NAND2_X1 U7840 ( .A1(n7161), .A2(n7160), .ZN(n7340) );
  INV_X1 U7841 ( .A(n8061), .ZN(n7160) );
  INV_X1 U7842 ( .A(n8026), .ZN(n8025) );
  AOI21_X1 U7843 ( .B1(n8028), .B2(n8029), .A(n13477), .ZN(n8026) );
  AND2_X1 U7844 ( .A1(n8012), .A2(n8011), .ZN(n8001) );
  NAND2_X1 U7845 ( .A1(n13490), .A2(n8003), .ZN(n8012) );
  NAND2_X1 U7846 ( .A1(n13832), .A2(n13486), .ZN(n8003) );
  NOR2_X1 U7847 ( .A1(n7306), .A2(n13536), .ZN(n7305) );
  NOR2_X1 U7848 ( .A1(n7308), .A2(n13958), .ZN(n7307) );
  NOR2_X1 U7849 ( .A1(n12966), .A2(n6956), .ZN(n12970) );
  AOI21_X1 U7850 ( .B1(n7501), .B2(n7504), .A(n6692), .ZN(n7498) );
  AOI21_X1 U7851 ( .B1(n8005), .B2(n6643), .A(n7333), .ZN(n13513) );
  INV_X1 U7852 ( .A(n8645), .ZN(n7402) );
  NAND2_X1 U7853 ( .A1(n15479), .A2(n14830), .ZN(n12632) );
  OR2_X1 U7854 ( .A1(n8806), .A2(n7496), .ZN(n7490) );
  NOR2_X1 U7855 ( .A1(n6566), .A2(n7498), .ZN(n7496) );
  AOI21_X1 U7856 ( .B1(n7503), .B2(n7504), .A(n11214), .ZN(n7500) );
  NAND2_X1 U7857 ( .A1(n9260), .A2(n10755), .ZN(n7341) );
  OAI21_X1 U7858 ( .B1(n10481), .B2(n7317), .A(n7316), .ZN(n8710) );
  NAND2_X1 U7859 ( .A1(n9260), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7316) );
  INV_X1 U7860 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7654) );
  INV_X1 U7861 ( .A(n12231), .ZN(n7031) );
  NAND2_X1 U7862 ( .A1(n15906), .A2(n11211), .ZN(n13410) );
  NAND2_X1 U7863 ( .A1(n11373), .A2(n10070), .ZN(n7066) );
  NAND2_X1 U7864 ( .A1(n7082), .A2(n7081), .ZN(n10077) );
  AOI21_X1 U7865 ( .B1(n7083), .B2(n7627), .A(n6748), .ZN(n7081) );
  AND2_X1 U7866 ( .A1(n13656), .A2(n13655), .ZN(n13657) );
  OAI22_X1 U7867 ( .A1(n13681), .A2(n6811), .B1(n6812), .B2(n6810), .ZN(n13716) );
  INV_X1 U7868 ( .A(n6815), .ZN(n6810) );
  NAND2_X1 U7869 ( .A1(n7378), .A2(n6815), .ZN(n6811) );
  INV_X1 U7870 ( .A(n6813), .ZN(n6812) );
  NOR2_X1 U7871 ( .A1(n8527), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n6849) );
  AND2_X1 U7872 ( .A1(n7361), .A2(n7259), .ZN(n8511) );
  INV_X1 U7873 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n7259) );
  OR2_X1 U7874 ( .A1(n13788), .A2(n8493), .ZN(n7782) );
  NOR2_X1 U7875 ( .A1(n8637), .A2(n7669), .ZN(n7668) );
  INV_X1 U7876 ( .A(n8634), .ZN(n7669) );
  NAND2_X1 U7877 ( .A1(n6894), .A2(n11509), .ZN(n6891) );
  NAND2_X1 U7878 ( .A1(n6914), .A2(n6912), .ZN(n8635) );
  NAND2_X1 U7879 ( .A1(n13959), .A2(n6915), .ZN(n6914) );
  NOR2_X1 U7880 ( .A1(n6916), .A2(n6561), .ZN(n6915) );
  INV_X1 U7881 ( .A(n13412), .ZN(n8665) );
  INV_X1 U7882 ( .A(n11213), .ZN(n11596) );
  AND2_X1 U7883 ( .A1(n13908), .A2(n13790), .ZN(n7685) );
  NAND2_X1 U7884 ( .A1(n7418), .A2(n6662), .ZN(n6920) );
  NAND2_X1 U7885 ( .A1(n7674), .A2(n13826), .ZN(n7673) );
  INV_X1 U7886 ( .A(n13990), .ZN(n7674) );
  AND2_X1 U7887 ( .A1(n7809), .A2(n6713), .ZN(n7808) );
  NAND2_X1 U7888 ( .A1(n7811), .A2(n7813), .ZN(n7809) );
  INV_X1 U7889 ( .A(n7811), .ZN(n7810) );
  NAND2_X1 U7890 ( .A1(n8646), .A2(n7401), .ZN(n7400) );
  AND2_X1 U7891 ( .A1(n13459), .A2(n8315), .ZN(n7788) );
  OR2_X1 U7892 ( .A1(n12245), .A2(n13580), .ZN(n13459) );
  AOI21_X1 U7893 ( .B1(n7591), .B2(n7593), .A(n6747), .ZN(n7589) );
  AND2_X1 U7894 ( .A1(n7595), .A2(n8234), .ZN(n7594) );
  NAND2_X1 U7895 ( .A1(n8224), .A2(n8223), .ZN(n7595) );
  NOR2_X1 U7896 ( .A1(n13089), .A2(n7822), .ZN(n7821) );
  INV_X1 U7897 ( .A(n12183), .ZN(n7822) );
  OR2_X1 U7898 ( .A1(n8860), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n8923) );
  INV_X1 U7899 ( .A(n7467), .ZN(n7468) );
  AND2_X1 U7900 ( .A1(n7876), .A2(n14424), .ZN(n7874) );
  NOR2_X1 U7901 ( .A1(n9129), .A2(n8821), .ZN(n7325) );
  NOR2_X1 U7902 ( .A1(n7847), .A2(n6560), .ZN(n7113) );
  NOR2_X1 U7903 ( .A1(n7847), .A2(n6560), .ZN(n7116) );
  AND2_X1 U7904 ( .A1(n6571), .A2(n7918), .ZN(n7917) );
  INV_X1 U7905 ( .A(n7848), .ZN(n7119) );
  NAND2_X1 U7906 ( .A1(n7859), .A2(n14235), .ZN(n7858) );
  OR2_X1 U7907 ( .A1(n11363), .A2(n8985), .ZN(n7857) );
  AND2_X1 U7908 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n8853) );
  AND2_X1 U7909 ( .A1(n10967), .A2(n10968), .ZN(n8910) );
  NOR2_X1 U7910 ( .A1(n6567), .A2(n7445), .ZN(n7444) );
  INV_X1 U7911 ( .A(n9369), .ZN(n7445) );
  NOR2_X1 U7912 ( .A1(n7433), .A2(n14369), .ZN(n7432) );
  INV_X1 U7913 ( .A(n14365), .ZN(n7433) );
  OAI21_X1 U7914 ( .B1(n7002), .B2(n7001), .A(n12977), .ZN(n7000) );
  NAND3_X1 U7915 ( .A1(n9315), .A2(n7843), .A3(n7842), .ZN(n9302) );
  INV_X1 U7916 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7843) );
  INV_X1 U7917 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n7842) );
  INV_X1 U7918 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8815) );
  NOR2_X1 U7919 ( .A1(n9735), .A2(n9417), .ZN(n6830) );
  NAND2_X1 U7920 ( .A1(n11064), .A2(n9477), .ZN(n9437) );
  INV_X1 U7921 ( .A(n9466), .ZN(n9934) );
  AND2_X1 U7922 ( .A1(n7887), .A2(n14863), .ZN(n7177) );
  NAND2_X1 U7923 ( .A1(n7176), .A2(n14863), .ZN(n7175) );
  INV_X1 U7924 ( .A(n7889), .ZN(n7176) );
  NAND2_X1 U7925 ( .A1(n15394), .A2(n15400), .ZN(n7998) );
  NOR2_X1 U7926 ( .A1(n15185), .A2(n7983), .ZN(n7982) );
  INV_X1 U7927 ( .A(n13024), .ZN(n7983) );
  INV_X1 U7928 ( .A(n14942), .ZN(n13060) );
  OR2_X1 U7929 ( .A1(n15461), .A2(n14838), .ZN(n15244) );
  NAND2_X1 U7930 ( .A1(n7967), .A2(n12498), .ZN(n13051) );
  NAND2_X1 U7931 ( .A1(n13051), .A2(n12632), .ZN(n13012) );
  OR2_X1 U7932 ( .A1(n15486), .A2(n14923), .ZN(n13048) );
  NAND2_X1 U7933 ( .A1(n15486), .A2(n14923), .ZN(n13047) );
  NAND2_X1 U7934 ( .A1(n9977), .A2(n11065), .ZN(n11064) );
  NOR2_X1 U7935 ( .A1(n7513), .A2(n9233), .ZN(n7511) );
  INV_X1 U7936 ( .A(n8744), .ZN(n7476) );
  NAND2_X1 U7937 ( .A1(n8748), .A2(n8749), .ZN(n7471) );
  INV_X1 U7938 ( .A(n9004), .ZN(n7383) );
  NAND2_X1 U7939 ( .A1(n7237), .A2(P1_ADDR_REG_1__SCAN_IN), .ZN(n7234) );
  NAND2_X1 U7940 ( .A1(n7236), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n10532) );
  INV_X1 U7941 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7236) );
  INV_X1 U7942 ( .A(n7287), .ZN(n10539) );
  NAND2_X1 U7943 ( .A1(n10948), .A2(n10947), .ZN(n10954) );
  OAI21_X1 U7944 ( .B1(n12129), .B2(n12128), .A(n12127), .ZN(n12274) );
  OR2_X1 U7945 ( .A1(n12325), .A2(n7031), .ZN(n7030) );
  INV_X1 U7946 ( .A(n7028), .ZN(n7027) );
  OAI21_X1 U7947 ( .B1(n12325), .B2(n7029), .A(n12327), .ZN(n7028) );
  OR2_X1 U7948 ( .A1(n12228), .A2(n7031), .ZN(n7029) );
  XNOR2_X1 U7949 ( .A(n12695), .B(n12178), .ZN(n11841) );
  AND2_X1 U7950 ( .A1(n7937), .A2(n7035), .ZN(n7034) );
  AND2_X1 U7951 ( .A1(n13272), .A2(n12688), .ZN(n7937) );
  NAND2_X1 U7952 ( .A1(n7938), .A2(n13251), .ZN(n7035) );
  INV_X1 U7953 ( .A(n13410), .ZN(n13409) );
  NAND2_X1 U7954 ( .A1(n7274), .A2(n7273), .ZN(n13248) );
  NAND2_X1 U7955 ( .A1(n7290), .A2(n12036), .ZN(n7289) );
  NAND2_X1 U7956 ( .A1(n8529), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8128) );
  AND2_X1 U7957 ( .A1(n11381), .A2(n10091), .ZN(n8087) );
  NOR2_X1 U7958 ( .A1(n11240), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10049) );
  NAND2_X1 U7959 ( .A1(n11377), .A2(n11378), .ZN(n11376) );
  NAND2_X1 U7960 ( .A1(n7567), .A2(n11683), .ZN(n11687) );
  NAND2_X1 U7961 ( .A1(n7066), .A2(n10523), .ZN(n11679) );
  NAND2_X1 U7962 ( .A1(n6570), .A2(n7557), .ZN(n11635) );
  OR2_X1 U7963 ( .A1(n7093), .A2(n7092), .ZN(n11638) );
  INV_X1 U7964 ( .A(n11615), .ZN(n7092) );
  NAND2_X1 U7965 ( .A1(n7093), .A2(n11615), .ZN(n10073) );
  AND2_X1 U7966 ( .A1(n10076), .A2(n7632), .ZN(n7631) );
  OR2_X1 U7967 ( .A1(n7629), .A2(n7628), .ZN(n11304) );
  NAND2_X1 U7968 ( .A1(n7630), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7629) );
  INV_X1 U7969 ( .A(n10149), .ZN(n7628) );
  OAI21_X1 U7970 ( .B1(n11312), .B2(n11311), .A(n11310), .ZN(n11309) );
  NAND2_X1 U7971 ( .A1(n13649), .A2(n13648), .ZN(n13676) );
  NOR2_X1 U7972 ( .A1(n13651), .A2(n13650), .ZN(n13677) );
  NOR2_X1 U7973 ( .A1(n7352), .A2(n13723), .ZN(n13702) );
  AND2_X1 U7974 ( .A1(n13701), .A2(n13700), .ZN(n7352) );
  INV_X1 U7975 ( .A(n7555), .ZN(n7552) );
  INV_X1 U7976 ( .A(n13737), .ZN(n7553) );
  OR2_X1 U7977 ( .A1(n13689), .A2(n7555), .ZN(n7554) );
  NAND2_X1 U7978 ( .A1(n6898), .A2(n6896), .ZN(n12700) );
  AOI21_X1 U7979 ( .B1(n6899), .B2(n6901), .A(n6897), .ZN(n6896) );
  NAND2_X1 U7980 ( .A1(n13781), .A2(n6899), .ZN(n6898) );
  INV_X1 U7981 ( .A(n13510), .ZN(n6897) );
  NAND2_X1 U7982 ( .A1(n6849), .A2(n6848), .ZN(n8554) );
  INV_X1 U7983 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n6848) );
  INV_X1 U7984 ( .A(n7679), .ZN(n7681) );
  INV_X1 U7985 ( .A(n6849), .ZN(n8539) );
  INV_X1 U7986 ( .A(n7782), .ZN(n7781) );
  NAND2_X1 U7987 ( .A1(n13802), .A2(n13551), .ZN(n7410) );
  AND2_X1 U7988 ( .A1(n8428), .A2(n8427), .ZN(n13848) );
  NAND2_X1 U7989 ( .A1(n6697), .A2(n6903), .ZN(n13860) );
  NAND2_X1 U7990 ( .A1(n8377), .A2(n6850), .ZN(n8421) );
  AND2_X1 U7991 ( .A1(n8376), .A2(n10245), .ZN(n6850) );
  AND2_X1 U7992 ( .A1(n8377), .A2(n8376), .ZN(n8391) );
  NAND2_X1 U7993 ( .A1(n8326), .A2(n10403), .ZN(n8360) );
  INV_X1 U7994 ( .A(n13581), .ZN(n12237) );
  NAND2_X1 U7995 ( .A1(n13432), .A2(n13430), .ZN(n6894) );
  AND2_X1 U7996 ( .A1(n13428), .A2(n13430), .ZN(n7773) );
  INV_X1 U7997 ( .A(n13588), .ZN(n11820) );
  OAI211_X1 U7998 ( .C1(n10063), .C2(n6902), .A(n8178), .B(n8177), .ZN(n12081)
         );
  XNOR2_X1 U7999 ( .A(n13591), .B(n8154), .ZN(n13951) );
  NAND2_X1 U8000 ( .A1(n8631), .A2(n8630), .ZN(n12708) );
  OR2_X1 U8001 ( .A1(n10039), .A2(n8625), .ZN(n8676) );
  INV_X1 U8002 ( .A(n13575), .ZN(n12703) );
  NAND2_X1 U8003 ( .A1(n8570), .A2(n8569), .ZN(n13902) );
  NAND2_X1 U8004 ( .A1(n6920), .A2(n7672), .ZN(n13802) );
  NAND2_X1 U8005 ( .A1(n8476), .A2(n13495), .ZN(n13800) );
  INV_X1 U8006 ( .A(SI_22_), .ZN(n8763) );
  NAND2_X1 U8007 ( .A1(n12047), .A2(n6887), .ZN(n6886) );
  OR2_X1 U8008 ( .A1(n13465), .A2(n13579), .ZN(n13462) );
  NAND2_X1 U8009 ( .A1(n12086), .A2(n12088), .ZN(n7789) );
  OR2_X1 U8010 ( .A1(n13514), .A2(n8672), .ZN(n15916) );
  NAND2_X1 U8011 ( .A1(n12046), .A2(n13407), .ZN(n12086) );
  OR2_X1 U8012 ( .A1(n7798), .A2(n8270), .ZN(n7795) );
  AOI21_X1 U8013 ( .B1(n11757), .B2(n13442), .A(n7799), .ZN(n7798) );
  INV_X1 U8014 ( .A(n13447), .ZN(n7799) );
  NOR2_X1 U8015 ( .A1(n11875), .A2(n8233), .ZN(n11758) );
  INV_X1 U8016 ( .A(n13960), .ZN(n15911) );
  INV_X1 U8017 ( .A(n15916), .ZN(n13886) );
  OAI21_X1 U8018 ( .B1(n8563), .B2(n8562), .A(n8564), .ZN(n8566) );
  MUX2_X1 U8019 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8118), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n8120) );
  NOR2_X1 U8020 ( .A1(n8534), .A2(n7621), .ZN(n7620) );
  INV_X1 U8021 ( .A(n8521), .ZN(n7621) );
  NOR2_X1 U8022 ( .A1(n8276), .A2(n7779), .ZN(n7778) );
  INV_X1 U8023 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8579) );
  NAND2_X1 U8024 ( .A1(n8507), .A2(n8506), .ZN(n8523) );
  OR2_X1 U8025 ( .A1(n8505), .A2(n11770), .ZN(n8506) );
  OAI21_X1 U8026 ( .B1(n8610), .B2(P3_IR_REG_23__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8583) );
  AND2_X1 U8027 ( .A1(n8619), .A2(n8621), .ZN(n7944) );
  INV_X1 U8028 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8619) );
  AND3_X1 U8029 ( .A1(n7941), .A2(n6535), .A3(n7038), .ZN(n8617) );
  INV_X1 U8030 ( .A(n7039), .ZN(n7037) );
  AOI21_X1 U8031 ( .B1(n7198), .B2(n8382), .A(n8398), .ZN(n7196) );
  AOI21_X1 U8032 ( .B1(n7224), .B2(n7226), .A(n7222), .ZN(n7221) );
  INV_X1 U8033 ( .A(n8337), .ZN(n7222) );
  INV_X1 U8034 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n10272) );
  AOI21_X1 U8035 ( .B1(n7204), .B2(n7206), .A(n7202), .ZN(n7201) );
  INV_X1 U8036 ( .A(n7598), .ZN(n7202) );
  XNOR2_X1 U8037 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n8287) );
  NAND2_X1 U8038 ( .A1(n7203), .A2(n8250), .ZN(n8272) );
  NAND2_X1 U8039 ( .A1(n7590), .A2(n7589), .ZN(n7203) );
  XNOR2_X1 U8040 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n8271) );
  OR2_X1 U8041 ( .A1(n8257), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n8274) );
  XNOR2_X1 U8042 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n8234) );
  NAND2_X1 U8043 ( .A1(n7191), .A2(n8194), .ZN(n8208) );
  NAND2_X1 U8044 ( .A1(n8908), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8144) );
  INV_X1 U8045 ( .A(n11244), .ZN(n6977) );
  INV_X1 U8046 ( .A(n13103), .ZN(n7824) );
  NAND2_X1 U8047 ( .A1(n10857), .A2(n10858), .ZN(n7820) );
  NAND2_X1 U8048 ( .A1(n7292), .A2(n14508), .ZN(n7816) );
  NAND2_X1 U8049 ( .A1(n7818), .A2(n12770), .ZN(n7817) );
  AOI21_X1 U8050 ( .B1(n6970), .B2(n6972), .A(n6968), .ZN(n6967) );
  INV_X1 U8051 ( .A(n14172), .ZN(n6968) );
  INV_X1 U8052 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9112) );
  INV_X1 U8053 ( .A(n11039), .ZN(n11042) );
  OR2_X1 U8054 ( .A1(n13135), .A2(n13134), .ZN(n14139) );
  AND2_X1 U8055 ( .A1(n14066), .A2(n14064), .ZN(n13134) );
  AND2_X1 U8056 ( .A1(n12763), .A2(n12988), .ZN(n10625) );
  AND2_X1 U8057 ( .A1(n6962), .A2(n11110), .ZN(n8048) );
  XNOR2_X1 U8058 ( .A(n6963), .B(n12987), .ZN(n6962) );
  NOR3_X1 U8059 ( .A1(n12982), .A2(n6964), .A3(n6611), .ZN(n6963) );
  NAND2_X1 U8060 ( .A1(n8049), .A2(n8051), .ZN(n8045) );
  NAND2_X1 U8061 ( .A1(n8048), .A2(n8043), .ZN(n7144) );
  NAND2_X1 U8062 ( .A1(n8044), .A2(n15844), .ZN(n8043) );
  AND2_X1 U8063 ( .A1(n9178), .A2(n9177), .ZN(n14059) );
  AND3_X1 U8064 ( .A1(n9117), .A2(n9116), .A3(n9115), .ZN(n14183) );
  AND3_X1 U8065 ( .A1(n9103), .A2(n9102), .A3(n9101), .ZN(n14205) );
  AND4_X1 U8066 ( .A1(n9073), .A2(n9072), .A3(n9071), .A4(n9070), .ZN(n14203)
         );
  AND4_X1 U8067 ( .A1(n9031), .A2(n9030), .A3(n9029), .A4(n9028), .ZN(n14091)
         );
  AND4_X1 U8068 ( .A1(n9000), .A2(n8999), .A3(n8998), .A4(n8997), .ZN(n12817)
         );
  AND4_X1 U8069 ( .A1(n8953), .A2(n8952), .A3(n8951), .A4(n8950), .ZN(n12809)
         );
  OR2_X1 U8070 ( .A1(n8931), .A2(n10641), .ZN(n8892) );
  OR2_X1 U8071 ( .A1(n10695), .A2(n10694), .ZN(n10806) );
  OR2_X1 U8072 ( .A1(n11010), .A2(n11009), .ZN(n11537) );
  INV_X1 U8073 ( .A(n7046), .ZN(n7045) );
  OAI21_X1 U8074 ( .B1(n12192), .B2(n7047), .A(n11983), .ZN(n7046) );
  XNOR2_X1 U8075 ( .A(n14295), .B(n14294), .ZN(n14298) );
  AND2_X1 U8076 ( .A1(n9217), .A2(n9225), .ZN(n14326) );
  NAND2_X1 U8077 ( .A1(n9193), .A2(n14379), .ZN(n7416) );
  INV_X1 U8078 ( .A(n7414), .ZN(n7415) );
  NAND2_X1 U8079 ( .A1(n7873), .A2(n7876), .ZN(n7872) );
  NAND2_X1 U8080 ( .A1(n9165), .A2(n7877), .ZN(n7873) );
  AOI21_X1 U8081 ( .B1(n7125), .B2(n7123), .A(n6691), .ZN(n7122) );
  INV_X1 U8082 ( .A(n7125), .ZN(n7124) );
  INV_X1 U8083 ( .A(n9136), .ZN(n7123) );
  NAND2_X1 U8084 ( .A1(n7845), .A2(n7121), .ZN(n7120) );
  NAND2_X1 U8085 ( .A1(n7119), .A2(n7121), .ZN(n7118) );
  NAND2_X1 U8086 ( .A1(n9053), .A2(n7848), .ZN(n7846) );
  INV_X1 U8087 ( .A(n7106), .ZN(n9052) );
  OAI21_X1 U8088 ( .B1(n9051), .B2(n14528), .A(n12958), .ZN(n7106) );
  OR2_X1 U8089 ( .A1(n7854), .A2(n8985), .ZN(n7853) );
  INV_X1 U8090 ( .A(n7852), .ZN(n7851) );
  OAI21_X1 U8091 ( .B1(n7855), .B2(n7854), .A(n12975), .ZN(n7852) );
  AND2_X1 U8092 ( .A1(n12973), .A2(n7435), .ZN(n7434) );
  OR2_X1 U8093 ( .A1(n12971), .A2(n7436), .ZN(n7435) );
  INV_X1 U8094 ( .A(n9351), .ZN(n7436) );
  NAND2_X1 U8095 ( .A1(n11362), .A2(n12971), .ZN(n11361) );
  OR2_X1 U8096 ( .A1(n14240), .A2(n15873), .ZN(n11796) );
  NAND2_X1 U8097 ( .A1(n8886), .A2(n8887), .ZN(n12795) );
  NAND2_X1 U8098 ( .A1(n8839), .A2(n6628), .ZN(n6981) );
  AND2_X1 U8099 ( .A1(n12734), .A2(n10212), .ZN(n6982) );
  NAND2_X1 U8100 ( .A1(n9278), .A2(n9277), .ZN(n14556) );
  NAND2_X1 U8101 ( .A1(n8784), .A2(n8783), .ZN(n14585) );
  AND2_X1 U8102 ( .A1(n14354), .A2(n9367), .ZN(n7007) );
  NAND2_X1 U8103 ( .A1(n14396), .A2(n7432), .ZN(n14366) );
  NAND2_X1 U8104 ( .A1(n14423), .A2(n6667), .ZN(n14391) );
  NOR2_X1 U8105 ( .A1(n7441), .A2(n7003), .ZN(n7002) );
  INV_X1 U8106 ( .A(n8092), .ZN(n7003) );
  AOI21_X1 U8107 ( .B1(n7440), .B2(n6960), .A(n6655), .ZN(n7439) );
  NAND2_X1 U8108 ( .A1(n14487), .A2(n8092), .ZN(n14464) );
  NAND2_X1 U8109 ( .A1(n14464), .A2(n14476), .ZN(n14463) );
  AND2_X1 U8110 ( .A1(n14634), .A2(n14116), .ZN(n9358) );
  NAND2_X1 U8111 ( .A1(n9354), .A2(n9353), .ZN(n14537) );
  OR2_X1 U8112 ( .A1(n14653), .A2(n7107), .ZN(n9353) );
  NAND2_X1 U8113 ( .A1(n14551), .A2(n6648), .ZN(n9354) );
  NAND2_X1 U8114 ( .A1(n7376), .A2(n7375), .ZN(n8781) );
  INV_X1 U8115 ( .A(n7850), .ZN(n7375) );
  INV_X1 U8116 ( .A(n7443), .ZN(n7376) );
  OR2_X1 U8117 ( .A1(n8796), .A2(n8780), .ZN(n8794) );
  NOR2_X1 U8118 ( .A1(n7443), .A2(n7442), .ZN(n8796) );
  OR3_X1 U8119 ( .A1(n9303), .A2(n9302), .A3(n9301), .ZN(n9307) );
  OR2_X1 U8120 ( .A1(n8927), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n8939) );
  INV_X1 U8121 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8908) );
  OR2_X1 U8122 ( .A1(n14908), .A2(n6559), .ZN(n7908) );
  INV_X1 U8123 ( .A(n14807), .ZN(n7186) );
  INV_X1 U8124 ( .A(n7303), .ZN(n9802) );
  OR2_X1 U8125 ( .A1(n7897), .A2(n7893), .ZN(n7892) );
  INV_X1 U8126 ( .A(n7899), .ZN(n7893) );
  AND2_X1 U8127 ( .A1(n14902), .A2(n7898), .ZN(n7897) );
  NAND2_X1 U8128 ( .A1(n14837), .A2(n7900), .ZN(n7898) );
  NOR2_X1 U8129 ( .A1(n7906), .A2(n7183), .ZN(n7904) );
  INV_X1 U8130 ( .A(n7906), .ZN(n7902) );
  NOR2_X1 U8131 ( .A1(n12002), .A2(n7168), .ZN(n7167) );
  INV_X1 U8132 ( .A(n11115), .ZN(n7168) );
  NAND2_X1 U8133 ( .A1(n7299), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9611) );
  INV_X1 U8134 ( .A(n9592), .ZN(n7299) );
  NOR2_X1 U8135 ( .A1(n14860), .A2(n6564), .ZN(n14796) );
  NAND2_X1 U8136 ( .A1(n6830), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9787) );
  NAND2_X1 U8137 ( .A1(n14760), .A2(n9868), .ZN(n7184) );
  NAND2_X1 U8138 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n9543) );
  NAND2_X1 U8139 ( .A1(n10989), .A2(n10990), .ZN(n11028) );
  NOR2_X1 U8140 ( .A1(n7189), .A2(n14872), .ZN(n7188) );
  INV_X1 U8141 ( .A(n9703), .ZN(n7189) );
  NAND2_X1 U8142 ( .A1(n14796), .A2(n14797), .ZN(n14795) );
  AND2_X1 U8143 ( .A1(n9664), .A2(n9663), .ZN(n9665) );
  OR2_X1 U8144 ( .A1(n9659), .A2(n9660), .ZN(n9664) );
  OR2_X1 U8145 ( .A1(n9722), .A2(n9721), .ZN(n7269) );
  NAND2_X1 U8146 ( .A1(n7293), .A2(n12573), .ZN(n12575) );
  AND2_X1 U8147 ( .A1(n6829), .A2(n9911), .ZN(n13069) );
  OR2_X1 U8148 ( .A1(n15161), .A2(n9907), .ZN(n6829) );
  INV_X1 U8149 ( .A(n10597), .ZN(n6863) );
  INV_X1 U8150 ( .A(n10598), .ZN(n6862) );
  NOR2_X1 U8151 ( .A1(n10762), .A2(n7538), .ZN(n15015) );
  AND2_X1 U8152 ( .A1(n10768), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7538) );
  OR2_X1 U8153 ( .A1(n10765), .A2(n10764), .ZN(n6875) );
  AND2_X1 U8154 ( .A1(n15037), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10912) );
  NAND2_X1 U8155 ( .A1(n6877), .A2(n6752), .ZN(n7540) );
  NOR2_X1 U8156 ( .A1(n15658), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n15657) );
  OR2_X1 U8157 ( .A1(n7998), .A2(n15150), .ZN(n7997) );
  INV_X1 U8158 ( .A(n7301), .ZN(n15140) );
  AND2_X1 U8159 ( .A1(n9945), .A2(n9985), .ZN(n15132) );
  NAND2_X1 U8160 ( .A1(n9904), .A2(n9903), .ZN(n15163) );
  NOR2_X1 U8161 ( .A1(n7977), .A2(n7461), .ZN(n7459) );
  INV_X1 U8162 ( .A(n7979), .ZN(n7977) );
  INV_X1 U8163 ( .A(n7980), .ZN(n7978) );
  NOR2_X1 U8164 ( .A1(n15171), .A2(n7980), .ZN(n7979) );
  NAND2_X1 U8165 ( .A1(n15211), .A2(n7460), .ZN(n15199) );
  INV_X1 U8166 ( .A(n15233), .ZN(n7712) );
  NAND2_X1 U8167 ( .A1(n15233), .A2(n7713), .ZN(n15215) );
  INV_X1 U8168 ( .A(n7708), .ZN(n7713) );
  OR2_X1 U8169 ( .A1(n9823), .A2(n14801), .ZN(n9835) );
  NOR2_X1 U8170 ( .A1(n15245), .A2(n7952), .ZN(n7951) );
  INV_X1 U8171 ( .A(n7956), .ZN(n7952) );
  AOI21_X1 U8172 ( .B1(n6867), .B2(n6865), .A(n6645), .ZN(n6864) );
  INV_X1 U8173 ( .A(n6867), .ZN(n6866) );
  INV_X1 U8174 ( .A(n13019), .ZN(n6865) );
  AOI21_X1 U8175 ( .B1(n7702), .B2(n7704), .A(n6660), .ZN(n7701) );
  OAI211_X1 U8176 ( .C1(n15339), .C2(n7195), .A(n7193), .B(n7702), .ZN(n6833)
         );
  AND2_X1 U8177 ( .A1(n15330), .A2(n15307), .ZN(n15299) );
  NOR2_X2 U8178 ( .A1(n15346), .A2(n15479), .ZN(n15330) );
  NAND2_X1 U8179 ( .A1(n11951), .A2(n11950), .ZN(n12017) );
  NAND2_X1 U8180 ( .A1(n10510), .A2(n12614), .ZN(n6879) );
  INV_X1 U8181 ( .A(n8089), .ZN(n7450) );
  AOI21_X1 U8182 ( .B1(n11347), .B2(n11346), .A(n11345), .ZN(n11578) );
  OR2_X1 U8183 ( .A1(n12414), .A2(n14955), .ZN(n11573) );
  INV_X1 U8184 ( .A(n15708), .ZN(n11194) );
  NAND2_X1 U8185 ( .A1(n7689), .A2(n12434), .ZN(n7688) );
  INV_X1 U8186 ( .A(n15223), .ZN(n15437) );
  INV_X1 U8187 ( .A(n15733), .ZN(n15678) );
  OR2_X1 U8188 ( .A1(n9977), .A2(n6809), .ZN(n11066) );
  NOR2_X1 U8189 ( .A1(n7483), .A2(n12613), .ZN(n7480) );
  AOI21_X1 U8190 ( .B1(n7488), .B2(n7486), .A(n6764), .ZN(n7485) );
  INV_X1 U8191 ( .A(n9261), .ZN(n7486) );
  INV_X1 U8192 ( .A(n7485), .ZN(n7483) );
  NOR2_X1 U8193 ( .A1(n7488), .A2(n12613), .ZN(n7482) );
  INV_X1 U8194 ( .A(n12613), .ZN(n7484) );
  NOR2_X1 U8195 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n7761) );
  INV_X1 U8196 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9392) );
  INV_X1 U8197 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9413) );
  INV_X1 U8198 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9412) );
  NAND2_X1 U8199 ( .A1(n7573), .A2(n8758), .ZN(n7572) );
  NAND2_X1 U8200 ( .A1(n6839), .A2(n6600), .ZN(n6838) );
  OR2_X1 U8201 ( .A1(n9685), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n9708) );
  OR2_X1 U8202 ( .A1(n9625), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n9626) );
  NAND2_X1 U8203 ( .A1(n9456), .A2(n6880), .ZN(n9514) );
  INV_X1 U8204 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6880) );
  NAND2_X1 U8205 ( .A1(n7531), .A2(n9394), .ZN(n7530) );
  INV_X1 U8206 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7531) );
  OR2_X1 U8207 ( .A1(n10537), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n7663) );
  NAND2_X1 U8208 ( .A1(n10537), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n10538) );
  NAND2_X1 U8209 ( .A1(n7257), .A2(n7356), .ZN(n7239) );
  NAND2_X1 U8210 ( .A1(n15581), .A2(n15580), .ZN(n15590) );
  OR2_X1 U8211 ( .A1(n15578), .A2(n15577), .ZN(n15581) );
  INV_X1 U8212 ( .A(n15949), .ZN(n11829) );
  INV_X1 U8213 ( .A(n13576), .ZN(n13775) );
  NAND2_X1 U8214 ( .A1(n8538), .A2(n8537), .ZN(n13229) );
  NAND2_X1 U8215 ( .A1(n12037), .A2(n12036), .ZN(n12225) );
  AND3_X1 U8216 ( .A1(n8165), .A2(n8164), .A3(n8163), .ZN(n13243) );
  INV_X1 U8217 ( .A(n13349), .ZN(n13319) );
  NAND2_X1 U8218 ( .A1(n7013), .A2(n6665), .ZN(n7011) );
  INV_X1 U8219 ( .A(n13334), .ZN(n7013) );
  INV_X1 U8220 ( .A(n13262), .ZN(n7018) );
  NAND2_X1 U8221 ( .A1(n13334), .A2(n6620), .ZN(n7012) );
  AND2_X1 U8222 ( .A1(n7014), .A2(n13325), .ZN(n7010) );
  OAI21_X1 U8223 ( .B1(n13262), .B2(n7016), .A(n7015), .ZN(n7014) );
  NAND2_X1 U8224 ( .A1(n13262), .A2(n7019), .ZN(n7015) );
  AND2_X1 U8225 ( .A1(n7017), .A2(n7019), .ZN(n7016) );
  NAND2_X1 U8226 ( .A1(n10063), .A2(n6580), .ZN(n7385) );
  OR2_X1 U8227 ( .A1(n10063), .A2(n11295), .ZN(n7384) );
  NAND2_X1 U8228 ( .A1(n7276), .A2(n7275), .ZN(n11605) );
  NAND2_X1 U8229 ( .A1(n13415), .A2(n12695), .ZN(n7275) );
  NAND2_X1 U8230 ( .A1(n11594), .A2(n13261), .ZN(n7276) );
  AND2_X1 U8231 ( .A1(n8445), .A2(n8444), .ZN(n13849) );
  AOI21_X1 U8232 ( .B1(n13221), .B2(n13220), .A(n13219), .ZN(n13280) );
  INV_X1 U8233 ( .A(n13300), .ZN(n7280) );
  NOR2_X1 U8234 ( .A1(n6573), .A2(n13360), .ZN(n7933) );
  NOR2_X1 U8235 ( .A1(n12693), .A2(n13812), .ZN(n7935) );
  AOI21_X1 U8236 ( .B1(n12693), .B2(n13497), .A(n13214), .ZN(n7936) );
  NAND2_X1 U8237 ( .A1(n8497), .A2(n8496), .ZN(n13912) );
  AND2_X1 U8238 ( .A1(n13240), .A2(n13238), .ZN(n11806) );
  AND2_X1 U8239 ( .A1(n8412), .A2(n8411), .ZN(n13864) );
  XNOR2_X1 U8240 ( .A(n13221), .B(n13212), .ZN(n13317) );
  NAND2_X1 U8241 ( .A1(n11593), .A2(n13889), .ZN(n13352) );
  AND2_X1 U8242 ( .A1(n11276), .A2(n11275), .ZN(n13357) );
  NAND2_X1 U8243 ( .A1(n13528), .A2(n13565), .ZN(n7332) );
  AOI21_X1 U8244 ( .B1(n6934), .B2(n7230), .A(n13556), .ZN(n13528) );
  INV_X1 U8245 ( .A(n13571), .ZN(n7804) );
  NAND4_X1 U8246 ( .A1(n8546), .A2(n8545), .A3(n8544), .A4(n8543), .ZN(n13768)
         );
  NOR2_X1 U8247 ( .A1(n6751), .A2(n7261), .ZN(n7260) );
  NAND2_X1 U8248 ( .A1(n13795), .A2(n8529), .ZN(n7262) );
  NAND2_X1 U8249 ( .A1(n8502), .A2(n8503), .ZN(n7261) );
  INV_X1 U8250 ( .A(n13848), .ZN(n13887) );
  NOR2_X1 U8251 ( .A1(n6547), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n6799) );
  NAND2_X1 U8252 ( .A1(n7554), .A2(n6569), .ZN(n13734) );
  AND2_X1 U8253 ( .A1(n6826), .A2(n6772), .ZN(n13732) );
  OAI21_X1 U8254 ( .B1(n13740), .B2(n6576), .A(n13748), .ZN(n6826) );
  AND2_X1 U8255 ( .A1(n10086), .A2(n7288), .ZN(n13754) );
  NAND2_X1 U8256 ( .A1(n8551), .A2(n8550), .ZN(n13269) );
  NAND2_X1 U8257 ( .A1(n8406), .A2(n8405), .ZN(n13853) );
  AND2_X1 U8258 ( .A1(n11213), .A2(n13735), .ZN(n15896) );
  NAND2_X1 U8259 ( .A1(n11275), .A2(n15896), .ZN(n15923) );
  NAND2_X1 U8260 ( .A1(n15960), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n7366) );
  XNOR2_X1 U8261 ( .A(n13362), .B(n8577), .ZN(n13901) );
  NAND2_X1 U8262 ( .A1(n15960), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n7426) );
  NAND2_X1 U8263 ( .A1(n13779), .A2(n13505), .ZN(n13765) );
  AOI21_X1 U8264 ( .B1(n7430), .B2(n13960), .A(n7427), .ZN(n13975) );
  NAND2_X1 U8265 ( .A1(n7429), .A2(n7428), .ZN(n7427) );
  XNOR2_X1 U8266 ( .A(n13767), .B(n13766), .ZN(n7430) );
  NAND2_X1 U8267 ( .A1(n13790), .A2(n13889), .ZN(n7428) );
  INV_X1 U8268 ( .A(n14013), .ZN(n14018) );
  NAND2_X1 U8269 ( .A1(n13141), .A2(n6607), .ZN(n7343) );
  OR2_X1 U8270 ( .A1(n13140), .A2(n14076), .ZN(n13141) );
  OR2_X1 U8271 ( .A1(n14054), .A2(n14058), .ZN(n8095) );
  NAND2_X1 U8272 ( .A1(n14164), .A2(n6794), .ZN(n6793) );
  AND2_X1 U8273 ( .A1(n11015), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14194) );
  NAND2_X1 U8274 ( .A1(n14190), .A2(n14191), .ZN(n7258) );
  INV_X1 U8275 ( .A(n14161), .ZN(n14213) );
  NAND2_X1 U8276 ( .A1(n10844), .A2(n15843), .ZN(n14211) );
  OR2_X1 U8277 ( .A1(n14311), .A2(n8961), .ZN(n9231) );
  NAND2_X1 U8278 ( .A1(n8805), .A2(n8804), .ZN(n14221) );
  NAND2_X1 U8279 ( .A1(n9201), .A2(n9200), .ZN(n14222) );
  OR2_X1 U8280 ( .A1(n14357), .A2(n8961), .ZN(n9201) );
  INV_X1 U8281 ( .A(n14059), .ZN(n14224) );
  NAND2_X1 U8282 ( .A1(n9150), .A2(n9149), .ZN(n14226) );
  INV_X1 U8283 ( .A(n12884), .ZN(n14228) );
  INV_X1 U8284 ( .A(n14091), .ZN(n9355) );
  OAI211_X1 U8285 ( .C1(n14250), .C2(n10641), .A(n10642), .B(n7052), .ZN(
        n14254) );
  NAND2_X1 U8286 ( .A1(n14250), .A2(n10641), .ZN(n7052) );
  NAND2_X1 U8287 ( .A1(n14264), .A2(n14265), .ZN(n14281) );
  NAND2_X1 U8288 ( .A1(n14274), .A2(n6806), .ZN(n15816) );
  OR2_X1 U8289 ( .A1(n14277), .A2(n8828), .ZN(n6806) );
  OR2_X1 U8290 ( .A1(n15834), .A2(n15833), .ZN(n15835) );
  OR2_X1 U8291 ( .A1(n14298), .A2(n15832), .ZN(n7048) );
  NAND2_X1 U8292 ( .A1(n14298), .A2(n15811), .ZN(n7337) );
  NAND2_X1 U8293 ( .A1(n10012), .A2(n10013), .ZN(n7422) );
  NAND2_X1 U8294 ( .A1(n9025), .A2(n9024), .ZN(n14648) );
  OR2_X1 U8295 ( .A1(n6626), .A2(n9169), .ZN(n7008) );
  NOR2_X1 U8296 ( .A1(n12721), .A2(n9292), .ZN(n9377) );
  XNOR2_X1 U8297 ( .A(n7772), .B(n12984), .ZN(n12723) );
  OAI21_X1 U8298 ( .B1(n10021), .B2(n12983), .A(n10020), .ZN(n12994) );
  NAND2_X1 U8299 ( .A1(n14581), .A2(n7111), .ZN(n14682) );
  AND2_X1 U8300 ( .A1(n14580), .A2(n6705), .ZN(n7111) );
  NAND2_X1 U8301 ( .A1(n9319), .A2(n9318), .ZN(n15860) );
  INV_X1 U8302 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n12407) );
  OR2_X1 U8303 ( .A1(n9494), .A2(n10487), .ZN(n7163) );
  OR2_X1 U8304 ( .A1(n9779), .A2(n10594), .ZN(n7164) );
  NAND2_X1 U8305 ( .A1(n9886), .A2(n9885), .ZN(n14822) );
  NAND2_X1 U8306 ( .A1(n9534), .A2(n9533), .ZN(n15756) );
  INV_X1 U8307 ( .A(n15163), .ZN(n15410) );
  NAND2_X1 U8308 ( .A1(n7179), .A2(n7178), .ZN(n14909) );
  OR2_X1 U8309 ( .A1(n7181), .A2(n6696), .ZN(n7178) );
  INV_X1 U8310 ( .A(n15634), .ZN(n14910) );
  INV_X1 U8311 ( .A(n14917), .ZN(n7372) );
  OR2_X1 U8312 ( .A1(n9998), .A2(n15517), .ZN(n14928) );
  AND2_X1 U8313 ( .A1(n15632), .A2(n15757), .ZN(n14930) );
  OAI21_X1 U8314 ( .B1(n12604), .B2(n7733), .A(n7732), .ZN(n12662) );
  NAND2_X1 U8315 ( .A1(n7741), .A2(n7734), .ZN(n7733) );
  NAND2_X1 U8316 ( .A1(n7731), .A2(n7741), .ZN(n7732) );
  INV_X1 U8317 ( .A(n7737), .ZN(n7734) );
  XNOR2_X1 U8318 ( .A(n7469), .B(n15314), .ZN(n12657) );
  NAND2_X1 U8319 ( .A1(n9930), .A2(n9929), .ZN(n14936) );
  NAND2_X1 U8320 ( .A1(n9897), .A2(n9896), .ZN(n14938) );
  NAND2_X1 U8321 ( .A1(n9876), .A2(n9875), .ZN(n14939) );
  NAND2_X1 U8322 ( .A1(n9859), .A2(n9858), .ZN(n14940) );
  OR2_X1 U8323 ( .A1(n14765), .A2(n9907), .ZN(n9859) );
  NAND2_X1 U8324 ( .A1(n9841), .A2(n9840), .ZN(n14941) );
  NAND2_X1 U8325 ( .A1(n9433), .A2(n9432), .ZN(n14943) );
  NAND2_X1 U8326 ( .A1(n9810), .A2(n9809), .ZN(n14944) );
  OR2_X1 U8327 ( .A1(n9608), .A2(n9457), .ZN(n9462) );
  OR2_X1 U8328 ( .A1(n9608), .A2(n15648), .ZN(n9469) );
  OR2_X1 U8329 ( .A1(n9594), .A2(n11296), .ZN(n9468) );
  NOR2_X1 U8330 ( .A1(n7519), .A2(n7525), .ZN(n7518) );
  INV_X1 U8331 ( .A(n10576), .ZN(n7519) );
  NOR2_X1 U8332 ( .A1(n15657), .A2(n6871), .ZN(n15066) );
  NAND2_X1 U8333 ( .A1(n6873), .A2(n6872), .ZN(n6871) );
  INV_X1 U8334 ( .A(n15049), .ZN(n6872) );
  INV_X1 U8335 ( .A(n15047), .ZN(n6873) );
  OAI22_X1 U8336 ( .A1(n15109), .A2(n15661), .B1(n15111), .B2(n15107), .ZN(
        n7534) );
  INV_X1 U8337 ( .A(n7536), .ZN(n7535) );
  OAI21_X1 U8338 ( .B1(n15110), .B2(n15111), .A(n15659), .ZN(n7536) );
  INV_X1 U8339 ( .A(n12627), .ZN(n15379) );
  OAI211_X1 U8340 ( .C1(n15140), .C2(n7965), .A(n7964), .B(n7963), .ZN(n7962)
         );
  NAND2_X1 U8341 ( .A1(n15387), .A2(n7966), .ZN(n7965) );
  INV_X1 U8342 ( .A(n13030), .ZN(n7964) );
  NAND2_X1 U8343 ( .A1(n15140), .A2(n13031), .ZN(n7963) );
  AND2_X1 U8344 ( .A1(n7219), .A2(n7217), .ZN(n15144) );
  NAND2_X1 U8345 ( .A1(n9870), .A2(n9869), .ZN(n15425) );
  NAND2_X1 U8346 ( .A1(n9850), .A2(n9849), .ZN(n15428) );
  NAND2_X1 U8347 ( .A1(n9629), .A2(n9628), .ZN(n14778) );
  OR2_X1 U8348 ( .A1(n9494), .A2(n10214), .ZN(n7462) );
  NOR2_X1 U8349 ( .A1(n6546), .A2(n15709), .ZN(n15295) );
  NAND2_X1 U8350 ( .A1(n6689), .A2(n6876), .ZN(n15524) );
  OR2_X1 U8351 ( .A1(n15403), .A2(n15760), .ZN(n6876) );
  INV_X1 U8352 ( .A(n15401), .ZN(n7455) );
  INV_X1 U8353 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n15545) );
  INV_X1 U8354 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10931) );
  NAND2_X1 U8355 ( .A1(n10570), .A2(n10571), .ZN(n7232) );
  NAND2_X1 U8356 ( .A1(n7232), .A2(n10677), .ZN(n7667) );
  INV_X1 U8357 ( .A(n10961), .ZN(n7651) );
  INV_X1 U8358 ( .A(n7239), .ZN(n7238) );
  INV_X1 U8359 ( .A(n12279), .ZN(n7664) );
  OR2_X1 U8360 ( .A1(n7256), .A2(n7255), .ZN(n15575) );
  INV_X1 U8361 ( .A(n15565), .ZN(n7256) );
  NAND2_X1 U8362 ( .A1(n7643), .A2(n7641), .ZN(n7635) );
  NAND2_X1 U8363 ( .A1(n7642), .A2(n7641), .ZN(n7634) );
  NOR2_X1 U8364 ( .A1(n7241), .A2(n7240), .ZN(n15618) );
  INV_X1 U8365 ( .A(n7267), .ZN(n7241) );
  NAND2_X1 U8366 ( .A1(n12792), .A2(n12794), .ZN(n8053) );
  AND2_X1 U8367 ( .A1(n12432), .A2(n12431), .ZN(n8103) );
  NAND2_X1 U8368 ( .A1(n12428), .A2(n12433), .ZN(n12432) );
  AND2_X1 U8369 ( .A1(n12430), .A2(n12426), .ZN(n12447) );
  NAND2_X1 U8370 ( .A1(n8069), .A2(n8073), .ZN(n7141) );
  INV_X1 U8371 ( .A(n8074), .ZN(n8073) );
  OAI21_X1 U8372 ( .B1(n8078), .B2(n8076), .A(n8075), .ZN(n8074) );
  NAND2_X1 U8373 ( .A1(n12460), .A2(n12462), .ZN(n7770) );
  OR2_X1 U8374 ( .A1(n12460), .A2(n12462), .ZN(n7769) );
  NAND2_X1 U8375 ( .A1(n7141), .A2(n12811), .ZN(n7140) );
  INV_X1 U8376 ( .A(n12810), .ZN(n7139) );
  INV_X1 U8377 ( .A(n7141), .ZN(n7137) );
  AND2_X1 U8378 ( .A1(n12488), .A2(n12489), .ZN(n7721) );
  NAND2_X1 U8379 ( .A1(n12479), .A2(n12476), .ZN(n7750) );
  INV_X1 U8380 ( .A(n7720), .ZN(n7716) );
  MUX2_X1 U8381 ( .A(n14203), .B(n12850), .S(n12777), .Z(n12861) );
  INV_X1 U8382 ( .A(n12503), .ZN(n12504) );
  OAI21_X1 U8383 ( .B1(n15341), .B2(n12502), .A(n12501), .ZN(n12503) );
  NAND2_X1 U8384 ( .A1(n13429), .A2(n13514), .ZN(n8020) );
  NAND2_X1 U8385 ( .A1(n13426), .A2(n13519), .ZN(n8021) );
  AOI21_X1 U8386 ( .B1(n8179), .B2(n13514), .A(n8019), .ZN(n8018) );
  NOR2_X1 U8387 ( .A1(n13425), .A2(n13514), .ZN(n8019) );
  NAND2_X1 U8388 ( .A1(n13418), .A2(n13514), .ZN(n6943) );
  OAI21_X1 U8389 ( .B1(n8034), .B2(n8033), .A(n12823), .ZN(n12842) );
  AOI21_X1 U8390 ( .B1(n6940), .B2(n13435), .A(n6939), .ZN(n13436) );
  AND2_X1 U8391 ( .A1(n13434), .A2(n13514), .ZN(n6939) );
  NAND2_X1 U8392 ( .A1(n8014), .A2(n6941), .ZN(n6940) );
  NOR2_X1 U8393 ( .A1(n8066), .A2(n8064), .ZN(n8063) );
  NAND2_X1 U8394 ( .A1(n12544), .A2(n12540), .ZN(n7757) );
  AND2_X1 U8395 ( .A1(n12892), .A2(n12893), .ZN(n8061) );
  NAND2_X1 U8396 ( .A1(n6952), .A2(n6950), .ZN(n6949) );
  NAND2_X1 U8397 ( .A1(n6951), .A2(n13514), .ZN(n6950) );
  INV_X1 U8398 ( .A(n13452), .ZN(n6951) );
  INV_X1 U8399 ( .A(n13545), .ZN(n6946) );
  NAND2_X1 U8400 ( .A1(n13458), .A2(n13519), .ZN(n6945) );
  AOI21_X1 U8401 ( .B1(n6948), .B2(n6947), .A(n6944), .ZN(n13464) );
  NAND2_X1 U8402 ( .A1(n13456), .A2(n13519), .ZN(n6947) );
  NAND2_X1 U8403 ( .A1(n6946), .A2(n6945), .ZN(n6944) );
  NAND2_X1 U8404 ( .A1(n6949), .A2(n13457), .ZN(n6948) );
  OR2_X1 U8405 ( .A1(n8056), .A2(n6792), .ZN(n12898) );
  AND2_X1 U8406 ( .A1(n8059), .A2(n7339), .ZN(n7338) );
  AND2_X1 U8407 ( .A1(n12901), .A2(n8039), .ZN(n8038) );
  NAND2_X1 U8408 ( .A1(n12899), .A2(n12902), .ZN(n8037) );
  NAND2_X1 U8409 ( .A1(n7767), .A2(n12551), .ZN(n7766) );
  INV_X1 U8410 ( .A(n13532), .ZN(n7308) );
  NOR2_X1 U8411 ( .A1(n8023), .A2(n8659), .ZN(n6955) );
  AND2_X1 U8412 ( .A1(n8027), .A2(n8024), .ZN(n8023) );
  NAND2_X1 U8413 ( .A1(n8025), .A2(n8656), .ZN(n8024) );
  OR2_X1 U8414 ( .A1(n13479), .A2(n13478), .ZN(n8027) );
  INV_X1 U8415 ( .A(n8011), .ZN(n8002) );
  NAND2_X1 U8416 ( .A1(n13824), .A2(n8001), .ZN(n8009) );
  AOI21_X1 U8417 ( .B1(n8006), .B2(n13498), .A(n13788), .ZN(n8005) );
  OAI21_X1 U8418 ( .B1(n8008), .B2(n8010), .A(n8013), .ZN(n8006) );
  AND2_X1 U8419 ( .A1(n7408), .A2(n13496), .ZN(n8013) );
  NOR2_X1 U8420 ( .A1(n13489), .A2(n8002), .ZN(n8010) );
  NAND2_X1 U8421 ( .A1(n7334), .A2(n13780), .ZN(n7333) );
  INV_X1 U8422 ( .A(n13504), .ZN(n7334) );
  NAND2_X1 U8423 ( .A1(n7158), .A2(n7150), .ZN(n7149) );
  AND2_X1 U8424 ( .A1(n7157), .A2(n12906), .ZN(n7150) );
  NAND2_X1 U8425 ( .A1(n7159), .A2(n7152), .ZN(n7151) );
  AND2_X1 U8426 ( .A1(n7157), .A2(n12903), .ZN(n7152) );
  NAND2_X1 U8427 ( .A1(n12559), .A2(n7764), .ZN(n7296) );
  INV_X1 U8428 ( .A(n9152), .ZN(n7495) );
  INV_X1 U8429 ( .A(n8721), .ZN(n7973) );
  OAI21_X1 U8430 ( .B1(n10481), .B2(P2_DATAO_REG_12__SCAN_IN), .A(n7264), .ZN(
        n8723) );
  NAND2_X1 U8431 ( .A1(n9260), .A2(n10707), .ZN(n7264) );
  AND2_X1 U8432 ( .A1(n7305), .A2(n13533), .ZN(n13540) );
  NOR2_X1 U8433 ( .A1(n13877), .A2(n7403), .ZN(n7311) );
  INV_X1 U8434 ( .A(n11624), .ZN(n6820) );
  OAI21_X1 U8435 ( .B1(n13680), .B2(n6814), .A(n13714), .ZN(n6813) );
  NAND2_X1 U8436 ( .A1(n13713), .A2(n13712), .ZN(n6815) );
  NAND2_X1 U8437 ( .A1(n7679), .A2(n7684), .ZN(n7678) );
  NOR2_X1 U8438 ( .A1(n13780), .A2(n7680), .ZN(n7677) );
  OR2_X1 U8439 ( .A1(n13269), .A2(n12703), .ZN(n13524) );
  AOI21_X1 U8440 ( .B1(n7788), .B2(n13542), .A(n7786), .ZN(n7785) );
  NAND2_X1 U8441 ( .A1(n8649), .A2(n13460), .ZN(n7786) );
  NOR2_X1 U8442 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n8251) );
  NOR2_X1 U8443 ( .A1(n14516), .A2(n14501), .ZN(n6961) );
  NOR2_X1 U8444 ( .A1(n9216), .A2(n9215), .ZN(n7323) );
  NAND2_X1 U8445 ( .A1(n7057), .A2(n7058), .ZN(n7467) );
  AOI21_X1 U8446 ( .B1(n7059), .B2(n6597), .A(n6765), .ZN(n7058) );
  NAND2_X1 U8447 ( .A1(n7490), .A2(n6582), .ZN(n7057) );
  NOR2_X1 U8448 ( .A1(n9835), .A2(n14886), .ZN(n6831) );
  AND2_X1 U8449 ( .A1(n13051), .A2(n6707), .ZN(n7705) );
  INV_X1 U8450 ( .A(n9232), .ZN(n9235) );
  AND2_X1 U8451 ( .A1(n7494), .A2(n7492), .ZN(n7491) );
  NAND2_X1 U8452 ( .A1(n6566), .A2(n7493), .ZN(n7492) );
  AOI21_X1 U8453 ( .B1(n7498), .B2(n7502), .A(n7495), .ZN(n7494) );
  INV_X1 U8454 ( .A(n7503), .ZN(n7493) );
  OAI21_X1 U8455 ( .B1(n8706), .B2(n7345), .A(n7344), .ZN(n8709) );
  NAND2_X1 U8456 ( .A1(n8706), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7344) );
  NAND2_X1 U8457 ( .A1(n8837), .A2(n8698), .ZN(n8701) );
  NOR2_X1 U8458 ( .A1(n8884), .A2(n8699), .ZN(n8700) );
  OAI21_X1 U8459 ( .B1(n8706), .B2(n7358), .A(n7357), .ZN(n8702) );
  NAND2_X1 U8460 ( .A1(n8706), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7357) );
  CLKBUF_X1 U8461 ( .A(n10250), .Z(n10365) );
  AND2_X1 U8462 ( .A1(n10759), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n10273) );
  INV_X1 U8463 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10533) );
  NAND2_X1 U8464 ( .A1(n8031), .A2(n13557), .ZN(n7312) );
  NAND2_X1 U8465 ( .A1(n13520), .A2(n13519), .ZN(n8032) );
  NAND2_X1 U8466 ( .A1(n13717), .A2(n15961), .ZN(n7379) );
  NAND2_X1 U8467 ( .A1(n6820), .A2(n6819), .ZN(n6817) );
  INV_X1 U8468 ( .A(n11625), .ZN(n6819) );
  AND2_X1 U8469 ( .A1(n10509), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n6927) );
  INV_X1 U8470 ( .A(n10147), .ZN(n7545) );
  INV_X1 U8471 ( .A(n10146), .ZN(n7541) );
  NAND2_X1 U8472 ( .A1(n7556), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7555) );
  INV_X1 U8473 ( .A(n13505), .ZN(n6901) );
  INV_X1 U8474 ( .A(n6900), .ZN(n6899) );
  OAI21_X1 U8475 ( .B1(n13780), .B2(n6901), .A(n13509), .ZN(n6900) );
  NAND2_X1 U8476 ( .A1(n13766), .A2(n7682), .ZN(n7679) );
  INV_X1 U8477 ( .A(n7685), .ZN(n7682) );
  NOR2_X1 U8478 ( .A1(n13780), .A2(n7405), .ZN(n7404) );
  INV_X1 U8479 ( .A(n7407), .ZN(n7405) );
  NAND2_X1 U8480 ( .A1(n7398), .A2(n8651), .ZN(n6905) );
  NOR2_X1 U8481 ( .A1(n8636), .A2(n7393), .ZN(n7388) );
  NOR2_X1 U8482 ( .A1(n7394), .A2(n7393), .ZN(n7391) );
  INV_X1 U8483 ( .A(n7668), .ZN(n7394) );
  INV_X1 U8484 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n7368) );
  INV_X1 U8485 ( .A(n12081), .ZN(n11811) );
  AND2_X1 U8486 ( .A1(n13524), .A2(n13523), .ZN(n13557) );
  OR2_X1 U8487 ( .A1(n13977), .A2(n13775), .ZN(n13509) );
  OR2_X1 U8488 ( .A1(n13923), .A2(n13836), .ZN(n13491) );
  NAND2_X1 U8489 ( .A1(n7807), .A2(n7811), .ZN(n13870) );
  NAND2_X1 U8490 ( .A1(n8381), .A2(n7812), .ZN(n7807) );
  NAND2_X1 U8491 ( .A1(n6623), .A2(n7787), .ZN(n7784) );
  INV_X1 U8492 ( .A(n7788), .ZN(n7787) );
  AND2_X1 U8493 ( .A1(n6623), .A2(n6888), .ZN(n6887) );
  NAND2_X1 U8494 ( .A1(n6889), .A2(n13407), .ZN(n6888) );
  NAND2_X1 U8495 ( .A1(n6887), .A2(n13408), .ZN(n6885) );
  INV_X1 U8496 ( .A(n7620), .ZN(n7614) );
  INV_X1 U8497 ( .A(n7611), .ZN(n7610) );
  OAI21_X1 U8498 ( .B1(n8432), .B2(n7612), .A(n8460), .ZN(n7611) );
  INV_X1 U8499 ( .A(n8434), .ZN(n7612) );
  INV_X1 U8500 ( .A(n8465), .ZN(n7608) );
  AND2_X1 U8501 ( .A1(n7610), .A2(n7212), .ZN(n7211) );
  NAND2_X1 U8502 ( .A1(n8413), .A2(n8402), .ZN(n7212) );
  NAND2_X1 U8503 ( .A1(n7211), .A2(n7213), .ZN(n7209) );
  INV_X1 U8504 ( .A(n8402), .ZN(n7213) );
  NAND2_X1 U8505 ( .A1(n8403), .A2(n7040), .ZN(n7039) );
  INV_X1 U8506 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7040) );
  INV_X1 U8507 ( .A(n10273), .ZN(n8400) );
  INV_X1 U8508 ( .A(n7225), .ZN(n7224) );
  OAI21_X1 U8509 ( .B1(n8317), .B2(n7226), .A(n8334), .ZN(n7225) );
  INV_X1 U8510 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n8726) );
  INV_X1 U8511 ( .A(n8250), .ZN(n7206) );
  AOI21_X1 U8512 ( .B1(n7600), .B2(n7602), .A(n6686), .ZN(n7598) );
  INV_X1 U8513 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n8289) );
  INV_X1 U8514 ( .A(n7205), .ZN(n7204) );
  OAI21_X1 U8515 ( .B1(n7589), .B2(n7206), .A(n7600), .ZN(n7205) );
  NAND2_X1 U8516 ( .A1(n8143), .A2(n8152), .ZN(n7604) );
  INV_X1 U8517 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9067) );
  INV_X1 U8518 ( .A(n12984), .ZN(n6965) );
  NOR2_X1 U8519 ( .A1(n14576), .A2(n13180), .ZN(n7914) );
  NAND2_X1 U8520 ( .A1(n7323), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n9250) );
  INV_X1 U8521 ( .A(n7323), .ZN(n9225) );
  NAND2_X1 U8522 ( .A1(n7467), .A2(n11935), .ZN(n7466) );
  INV_X1 U8523 ( .A(n7872), .ZN(n7870) );
  INV_X1 U8524 ( .A(n7874), .ZN(n7867) );
  NOR2_X1 U8525 ( .A1(n6670), .A2(n7127), .ZN(n7125) );
  NOR2_X1 U8526 ( .A1(n9068), .A2(n9067), .ZN(n7324) );
  NAND2_X1 U8527 ( .A1(n14529), .A2(n12959), .ZN(n9051) );
  NAND2_X1 U8528 ( .A1(n7108), .A2(n7107), .ZN(n14528) );
  NOR2_X1 U8529 ( .A1(n6568), .A2(n9352), .ZN(n6987) );
  INV_X1 U8530 ( .A(n12159), .ZN(n7854) );
  INV_X1 U8531 ( .A(n7858), .ZN(n7856) );
  OR2_X1 U8532 ( .A1(n11558), .A2(n12795), .ZN(n11557) );
  NOR2_X1 U8533 ( .A1(n11706), .A2(n12784), .ZN(n10965) );
  INV_X1 U8534 ( .A(n7432), .ZN(n7005) );
  NAND2_X1 U8535 ( .A1(n7587), .A2(n7586), .ZN(n9364) );
  AND2_X1 U8536 ( .A1(n14165), .A2(n9156), .ZN(n7586) );
  NOR2_X1 U8537 ( .A1(n14620), .A2(n7916), .ZN(n7915) );
  INV_X1 U8538 ( .A(n7917), .ZN(n7916) );
  XNOR2_X1 U8539 ( .A(n14668), .B(n14236), .ZN(n12969) );
  INV_X1 U8540 ( .A(n10977), .ZN(n12965) );
  NAND3_X1 U8541 ( .A1(n8811), .A2(n8813), .A3(n8779), .ZN(n7850) );
  INV_X1 U8542 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8761) );
  NOR2_X1 U8543 ( .A1(n9787), .A2(n9418), .ZN(n7303) );
  NOR2_X1 U8544 ( .A1(n9671), .A2(n10915), .ZN(n7304) );
  INV_X1 U8545 ( .A(n7177), .ZN(n7172) );
  INV_X1 U8546 ( .A(n7175), .ZN(n7173) );
  INV_X1 U8547 ( .A(n7885), .ZN(n7884) );
  OAI21_X1 U8548 ( .B1(n14797), .B2(n7886), .A(n14882), .ZN(n7885) );
  NOR2_X1 U8549 ( .A1(n12572), .A2(n12569), .ZN(n7763) );
  INV_X1 U8550 ( .A(n12569), .ZN(n7762) );
  INV_X1 U8551 ( .A(n9426), .ZN(n9424) );
  NOR2_X1 U8552 ( .A1(n7710), .A2(n15227), .ZN(n7228) );
  NAND2_X1 U8553 ( .A1(n7995), .A2(n14805), .ZN(n7994) );
  NOR2_X1 U8554 ( .A1(n15298), .A2(n15461), .ZN(n7265) );
  NAND2_X1 U8555 ( .A1(n13062), .A2(n13061), .ZN(n7708) );
  INV_X1 U8556 ( .A(n6831), .ZN(n9852) );
  NOR2_X1 U8557 ( .A1(n15447), .A2(n15455), .ZN(n7995) );
  NOR2_X1 U8558 ( .A1(n13021), .A2(n6868), .ZN(n6867) );
  INV_X1 U8559 ( .A(n13020), .ZN(n6868) );
  INV_X1 U8560 ( .A(n13050), .ZN(n7195) );
  AND2_X1 U8561 ( .A1(n7706), .A2(n7703), .ZN(n7702) );
  NAND2_X1 U8562 ( .A1(n7705), .A2(n13012), .ZN(n7703) );
  AND2_X1 U8563 ( .A1(n15296), .A2(n15293), .ZN(n7706) );
  INV_X1 U8564 ( .A(n7705), .ZN(n7704) );
  NOR2_X1 U8565 ( .A1(n15368), .A2(n14949), .ZN(n13044) );
  INV_X1 U8566 ( .A(n13047), .ZN(n13045) );
  AND2_X1 U8567 ( .A1(n11342), .A2(n12417), .ZN(n7991) );
  NAND2_X1 U8568 ( .A1(n11191), .A2(n8084), .ZN(n11337) );
  NOR2_X2 U8569 ( .A1(n15203), .A2(n15425), .ZN(n15191) );
  INV_X1 U8570 ( .A(n7265), .ZN(n15285) );
  INV_X1 U8571 ( .A(n15328), .ZN(n13011) );
  NOR2_X1 U8572 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n9385) );
  NAND2_X1 U8573 ( .A1(n6565), .A2(n6668), .ZN(n7504) );
  INV_X1 U8574 ( .A(n9076), .ZN(n6837) );
  NAND2_X1 U8575 ( .A1(n6841), .A2(n6840), .ZN(n6839) );
  INV_X1 U8576 ( .A(n9078), .ZN(n6840) );
  NAND2_X1 U8577 ( .A1(n6795), .A2(n8742), .ZN(n9074) );
  OR2_X1 U8578 ( .A1(n9708), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n9724) );
  NOR2_X1 U8579 ( .A1(n7969), .A2(n9055), .ZN(n7968) );
  INV_X1 U8580 ( .A(n7971), .ZN(n7969) );
  INV_X1 U8581 ( .A(n7103), .ZN(n7102) );
  OAI21_X1 U8582 ( .B1(n8716), .B2(n7104), .A(n8721), .ZN(n7103) );
  OR2_X1 U8583 ( .A1(n9604), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9625) );
  INV_X1 U8584 ( .A(n8936), .ZN(n7099) );
  NAND2_X1 U8585 ( .A1(n8865), .A2(n8704), .ZN(n8919) );
  NAND2_X1 U8586 ( .A1(n8701), .A2(n8700), .ZN(n8864) );
  NAND2_X1 U8587 ( .A1(n7315), .A2(n7314), .ZN(n7660) );
  NAND2_X1 U8588 ( .A1(n10956), .A2(n10955), .ZN(n11717) );
  OR2_X1 U8589 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n10954), .ZN(n10955) );
  NAND2_X1 U8590 ( .A1(n12277), .A2(n12276), .ZN(n12291) );
  OR2_X1 U8591 ( .A1(n12274), .A2(n12273), .ZN(n12277) );
  INV_X1 U8592 ( .A(n7653), .ZN(n7254) );
  INV_X1 U8593 ( .A(n15572), .ZN(n7253) );
  NOR2_X1 U8594 ( .A1(n13259), .A2(n7022), .ZN(n7021) );
  INV_X1 U8595 ( .A(n13335), .ZN(n7022) );
  INV_X1 U8596 ( .A(n7021), .ZN(n7017) );
  INV_X1 U8597 ( .A(n7020), .ZN(n7019) );
  OAI22_X1 U8598 ( .A1(n13259), .A2(n7024), .B1(n13768), .B2(n13258), .ZN(
        n7020) );
  INV_X1 U8599 ( .A(n11839), .ZN(n12172) );
  XNOR2_X1 U8600 ( .A(n12695), .B(n13243), .ZN(n11808) );
  NAND2_X1 U8601 ( .A1(n12229), .A2(n12228), .ZN(n12353) );
  AOI21_X1 U8602 ( .B1(n7034), .B2(n7939), .A(n6619), .ZN(n7032) );
  OR2_X1 U8603 ( .A1(n8421), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8423) );
  INV_X1 U8604 ( .A(n13527), .ZN(n8031) );
  AND4_X1 U8605 ( .A1(n13381), .A2(n13380), .A3(n13379), .A4(n13378), .ZN(
        n13758) );
  NAND2_X1 U8606 ( .A1(n8572), .A2(n11531), .ZN(n8159) );
  AND2_X1 U8607 ( .A1(n8138), .A2(n8139), .ZN(n6917) );
  OR2_X1 U8608 ( .A1(n13376), .A2(n8137), .ZN(n8138) );
  OR2_X1 U8609 ( .A1(n13377), .A2(n11280), .ZN(n8139) );
  OR2_X1 U8610 ( .A1(n11288), .A2(n15961), .ZN(n11290) );
  AOI21_X1 U8611 ( .B1(n11382), .B2(n11381), .A(n11380), .ZN(n13600) );
  XNOR2_X1 U8612 ( .A(n11697), .B(n11506), .ZN(n11683) );
  NAND2_X1 U8613 ( .A1(n7568), .A2(n11684), .ZN(n13594) );
  INV_X1 U8614 ( .A(n7569), .ZN(n7568) );
  NAND2_X1 U8615 ( .A1(n6785), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n13595) );
  OAI21_X1 U8616 ( .B1(n13600), .B2(n13599), .A(n8094), .ZN(n13598) );
  NAND2_X1 U8617 ( .A1(n6822), .A2(n11645), .ZN(n6821) );
  NAND2_X1 U8618 ( .A1(n6818), .A2(n6817), .ZN(n11623) );
  NAND2_X1 U8619 ( .A1(n11618), .A2(n10074), .ZN(n7075) );
  AOI21_X1 U8620 ( .B1(n11137), .B2(n10163), .A(n10162), .ZN(n11312) );
  AOI21_X1 U8621 ( .B1(n7626), .B2(n6581), .A(n6786), .ZN(n7083) );
  NAND2_X1 U8622 ( .A1(n7541), .A2(n7545), .ZN(n7543) );
  NAND2_X1 U8623 ( .A1(n11308), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n11307) );
  NAND2_X1 U8624 ( .A1(n7566), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7565) );
  NAND2_X1 U8625 ( .A1(n7087), .A2(n7091), .ZN(n10083) );
  INV_X1 U8626 ( .A(n10082), .ZN(n7087) );
  NAND3_X1 U8627 ( .A1(n13631), .A2(n13630), .A3(n13629), .ZN(n13633) );
  NAND2_X1 U8628 ( .A1(n13615), .A2(n10081), .ZN(n10082) );
  NAND2_X1 U8629 ( .A1(n10082), .A2(n10744), .ZN(n10085) );
  NAND2_X1 U8630 ( .A1(n6746), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n13637) );
  NAND2_X1 U8631 ( .A1(n13643), .A2(n7380), .ZN(n13663) );
  NAND2_X1 U8632 ( .A1(n7558), .A2(n13678), .ZN(n7561) );
  OR2_X1 U8633 ( .A1(n13657), .A2(n13678), .ZN(n13672) );
  NAND2_X1 U8634 ( .A1(n13658), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n13674) );
  NAND2_X1 U8635 ( .A1(n13658), .A2(n6777), .ZN(n7067) );
  NAND2_X1 U8636 ( .A1(n7069), .A2(n7071), .ZN(n7068) );
  INV_X1 U8637 ( .A(n13672), .ZN(n7069) );
  NAND2_X1 U8638 ( .A1(n13665), .A2(n13664), .ZN(n7559) );
  NAND2_X1 U8639 ( .A1(n13691), .A2(n7378), .ZN(n13715) );
  AND2_X1 U8640 ( .A1(n13722), .A2(n13725), .ZN(n6825) );
  NOR2_X1 U8641 ( .A1(n13719), .A2(n13718), .ZN(n13740) );
  OAI21_X1 U8642 ( .B1(n13800), .B2(n7782), .A(n7780), .ZN(n13781) );
  AOI21_X1 U8643 ( .B1(n7781), .B2(n13551), .A(n13503), .ZN(n7780) );
  INV_X1 U8644 ( .A(n7683), .ZN(n13773) );
  NAND2_X1 U8645 ( .A1(n8454), .A2(n13274), .ZN(n8469) );
  OR2_X1 U8646 ( .A1(n13998), .A2(n13849), .ZN(n8088) );
  INV_X1 U8647 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n8437) );
  AND2_X1 U8648 ( .A1(n8438), .A2(n8437), .ZN(n8454) );
  NOR2_X1 U8649 ( .A1(n8423), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8438) );
  NAND2_X1 U8650 ( .A1(n13882), .A2(n8651), .ZN(n13859) );
  INV_X1 U8651 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n8376) );
  NOR2_X1 U8652 ( .A1(n8309), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8326) );
  OAI21_X1 U8653 ( .B1(n11758), .B2(n7792), .A(n7790), .ZN(n12047) );
  AOI21_X1 U8654 ( .B1(n7793), .B2(n7797), .A(n7791), .ZN(n7790) );
  INV_X1 U8655 ( .A(n7793), .ZN(n7792) );
  AND2_X1 U8656 ( .A1(n7795), .A2(n13455), .ZN(n7793) );
  NAND2_X1 U8657 ( .A1(n12047), .A2(n13453), .ZN(n12046) );
  NAND2_X1 U8658 ( .A1(n6845), .A2(n6844), .ZN(n8309) );
  INV_X1 U8659 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n6844) );
  INV_X1 U8660 ( .A(n8293), .ZN(n6845) );
  NAND2_X1 U8661 ( .A1(n6847), .A2(n6846), .ZN(n8293) );
  INV_X1 U8662 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n6846) );
  INV_X1 U8663 ( .A(n8280), .ZN(n6847) );
  INV_X1 U8664 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8262) );
  NAND2_X1 U8665 ( .A1(n7670), .A2(n8638), .ZN(n11759) );
  NAND2_X1 U8666 ( .A1(n8635), .A2(n7668), .ZN(n7392) );
  INV_X1 U8667 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n8240) );
  AND2_X1 U8668 ( .A1(n8241), .A2(n8240), .ZN(n8263) );
  NAND2_X1 U8669 ( .A1(n6892), .A2(n6890), .ZN(n11876) );
  NAND2_X1 U8670 ( .A1(n6891), .A2(n8215), .ZN(n6890) );
  INV_X1 U8671 ( .A(n13539), .ZN(n13437) );
  INV_X1 U8672 ( .A(n13587), .ZN(n11880) );
  NOR2_X1 U8673 ( .A1(n8197), .A2(n6852), .ZN(n8241) );
  NAND2_X1 U8674 ( .A1(n7368), .A2(n6853), .ZN(n6852) );
  INV_X1 U8675 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n6853) );
  NAND2_X1 U8676 ( .A1(n6851), .A2(n7368), .ZN(n8216) );
  INV_X1 U8677 ( .A(n8197), .ZN(n6851) );
  INV_X1 U8678 ( .A(n13586), .ZN(n11840) );
  NAND2_X1 U8679 ( .A1(n8635), .A2(n8634), .ZN(n11491) );
  NAND2_X1 U8680 ( .A1(n8181), .A2(n8180), .ZN(n8197) );
  INV_X1 U8681 ( .A(n8633), .ZN(n6911) );
  AOI21_X1 U8682 ( .B1(n8633), .B2(n6916), .A(n6561), .ZN(n6910) );
  NAND2_X1 U8683 ( .A1(n13959), .A2(n13958), .ZN(n13957) );
  OR2_X1 U8684 ( .A1(n13372), .A2(n10515), .ZN(n7777) );
  INV_X1 U8685 ( .A(n13590), .ZN(n13955) );
  INV_X1 U8686 ( .A(n11777), .ZN(n13954) );
  AND4_X1 U8687 ( .A1(n13381), .A2(n8671), .A3(n8670), .A4(n8669), .ZN(n13385)
         );
  INV_X1 U8688 ( .A(n13768), .ZN(n10028) );
  INV_X1 U8689 ( .A(n13557), .ZN(n13521) );
  NAND2_X1 U8690 ( .A1(n13781), .A2(n13780), .ZN(n13779) );
  NOR2_X1 U8691 ( .A1(n13773), .A2(n7685), .ZN(n13767) );
  NAND2_X1 U8692 ( .A1(n13768), .A2(n13886), .ZN(n7429) );
  AND2_X1 U8693 ( .A1(n13491), .A2(n13492), .ZN(n13824) );
  INV_X1 U8694 ( .A(n13833), .ZN(n8663) );
  AOI21_X1 U8695 ( .B1(n7808), .B2(n7810), .A(n6693), .ZN(n7806) );
  AND3_X1 U8696 ( .A1(n8346), .A2(n8345), .A3(n8344), .ZN(n13344) );
  NAND2_X1 U8697 ( .A1(n7400), .A2(n8647), .ZN(n12314) );
  NAND2_X1 U8698 ( .A1(n7400), .A2(n6907), .ZN(n12316) );
  NAND2_X1 U8699 ( .A1(n7789), .A2(n7788), .ZN(n12313) );
  INV_X1 U8700 ( .A(n8578), .ZN(n6882) );
  XNOR2_X1 U8701 ( .A(n8505), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n8504) );
  XNOR2_X1 U8702 ( .A(n8612), .B(n8611), .ZN(n11259) );
  INV_X1 U8703 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8611) );
  AND2_X1 U8704 ( .A1(n8494), .A2(n8480), .ZN(n8481) );
  NAND2_X1 U8705 ( .A1(n8433), .A2(n8432), .ZN(n7609) );
  OR2_X1 U8706 ( .A1(n8447), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8449) );
  AOI21_X1 U8707 ( .B1(n8383), .B2(n7199), .A(n6762), .ZN(n7198) );
  INV_X1 U8708 ( .A(n8370), .ZN(n7199) );
  NAND2_X1 U8709 ( .A1(n7223), .A2(n8319), .ZN(n8348) );
  OR2_X1 U8710 ( .A1(n8338), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n8353) );
  XNOR2_X1 U8711 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8300) );
  INV_X1 U8712 ( .A(n7594), .ZN(n7593) );
  AOI21_X1 U8713 ( .B1(n7594), .B2(n7592), .A(n6685), .ZN(n7591) );
  INV_X1 U8714 ( .A(n8223), .ZN(n7592) );
  AND2_X1 U8715 ( .A1(n10493), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8224) );
  OR2_X1 U8716 ( .A1(n8205), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n8226) );
  INV_X1 U8717 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n8209) );
  XNOR2_X1 U8718 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n8207) );
  OR2_X1 U8719 ( .A1(n8253), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n8188) );
  NAND2_X1 U8720 ( .A1(n8175), .A2(n8174), .ZN(n8193) );
  XNOR2_X1 U8721 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n8192) );
  XNOR2_X1 U8722 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8172) );
  NAND2_X1 U8723 ( .A1(n10595), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8152) );
  INV_X1 U8724 ( .A(n8144), .ZN(n7605) );
  INV_X1 U8725 ( .A(n8143), .ZN(n7606) );
  AND2_X1 U8726 ( .A1(n13168), .A2(n13167), .ZN(n13171) );
  AND2_X1 U8727 ( .A1(n13108), .A2(n13107), .ZN(n14107) );
  NAND2_X1 U8728 ( .A1(n13165), .A2(n13164), .ZN(n7839) );
  INV_X1 U8729 ( .A(n13125), .ZN(n7826) );
  NAND2_X1 U8730 ( .A1(n7347), .A2(n7346), .ZN(n14076) );
  INV_X1 U8731 ( .A(n13139), .ZN(n7346) );
  AND2_X1 U8732 ( .A1(n13147), .A2(n14163), .ZN(n6794) );
  NAND2_X1 U8733 ( .A1(n7321), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9044) );
  INV_X1 U8734 ( .A(n9042), .ZN(n7321) );
  NAND2_X1 U8735 ( .A1(n6980), .A2(n13102), .ZN(n14087) );
  NAND2_X1 U8736 ( .A1(n8788), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9011) );
  INV_X1 U8737 ( .A(n8994), .ZN(n8788) );
  NAND2_X1 U8738 ( .A1(n7322), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n9042) );
  INV_X1 U8739 ( .A(n9011), .ZN(n7322) );
  AOI21_X1 U8740 ( .B1(n7821), .B2(n6971), .A(n6640), .ZN(n6970) );
  INV_X1 U8741 ( .A(n12144), .ZN(n6971) );
  INV_X1 U8742 ( .A(n7821), .ZN(n6972) );
  NAND3_X1 U8743 ( .A1(n7815), .A2(n7820), .A3(n7819), .ZN(n10881) );
  NAND2_X1 U8744 ( .A1(n14124), .A2(n14123), .ZN(n14122) );
  OR2_X1 U8745 ( .A1(n10839), .A2(n10638), .ZN(n14204) );
  NAND2_X1 U8746 ( .A1(n11229), .A2(n11230), .ZN(n11245) );
  AND2_X1 U8747 ( .A1(n12927), .A2(n12942), .ZN(n12928) );
  AND2_X1 U8748 ( .A1(n9271), .A2(n9270), .ZN(n12924) );
  AOI21_X1 U8749 ( .B1(n10682), .B2(n10681), .A(n6805), .ZN(n10713) );
  AND2_X1 U8750 ( .A1(n10689), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6805) );
  AOI21_X1 U8751 ( .B1(n6594), .B2(n15833), .A(n7055), .ZN(n7054) );
  OR2_X1 U8752 ( .A1(n9080), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n9094) );
  NAND2_X1 U8753 ( .A1(n7041), .A2(n11655), .ZN(n11980) );
  NAND2_X1 U8754 ( .A1(n11652), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7041) );
  AOI21_X1 U8755 ( .B1(n11973), .B2(P2_REG1_REG_15__SCAN_IN), .A(n6631), .ZN(
        n12194) );
  INV_X1 U8756 ( .A(n11985), .ZN(n7047) );
  OR2_X1 U8757 ( .A1(n12337), .A2(n14289), .ZN(n14292) );
  NAND2_X1 U8758 ( .A1(n9265), .A2(n9264), .ZN(n12926) );
  AOI22_X1 U8759 ( .A1(n14218), .A2(n14192), .B1(n12741), .B2(n14216), .ZN(
        n9287) );
  INV_X1 U8760 ( .A(n7864), .ZN(n7863) );
  OAI21_X1 U8761 ( .B1(n14303), .B2(n7865), .A(n6672), .ZN(n7864) );
  NOR2_X1 U8762 ( .A1(n14303), .A2(n7862), .ZN(n7861) );
  INV_X1 U8763 ( .A(n12957), .ZN(n7862) );
  INV_X1 U8764 ( .A(n14204), .ZN(n14193) );
  OAI21_X1 U8765 ( .B1(n14346), .B2(n14221), .A(n14335), .ZN(n14320) );
  AND2_X1 U8766 ( .A1(n7865), .A2(n12957), .ZN(n14319) );
  NOR2_X1 U8767 ( .A1(n14378), .A2(n14379), .ZN(n14377) );
  NOR3_X1 U8768 ( .A1(n14605), .A2(n14600), .A3(n14595), .ZN(n7911) );
  NOR2_X1 U8769 ( .A1(n14600), .A2(n14605), .ZN(n7910) );
  NAND2_X1 U8770 ( .A1(n7325), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n9157) );
  OR2_X1 U8771 ( .A1(n9157), .A2(n14081), .ZN(n9172) );
  NAND2_X1 U8772 ( .A1(n8790), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9129) );
  INV_X1 U8773 ( .A(n7325), .ZN(n9144) );
  NAND2_X1 U8774 ( .A1(n7845), .A2(n7113), .ZN(n7117) );
  AOI21_X1 U8775 ( .B1(n6621), .B2(n9104), .A(n6560), .ZN(n7115) );
  NAND2_X1 U8776 ( .A1(n14522), .A2(n6571), .ZN(n8097) );
  NAND2_X1 U8777 ( .A1(n7324), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9099) );
  INV_X1 U8778 ( .A(n7324), .ZN(n9087) );
  NAND2_X1 U8779 ( .A1(n14522), .A2(n14634), .ZN(n14506) );
  NAND2_X1 U8780 ( .A1(n14653), .A2(n14152), .ZN(n14529) );
  OAI211_X1 U8781 ( .C1(n6991), .C2(n11362), .A(n6990), .B(n6989), .ZN(n14551)
         );
  NAND2_X1 U8782 ( .A1(n6680), .A2(n6995), .ZN(n6990) );
  OR2_X1 U8783 ( .A1(n6994), .A2(n9352), .ZN(n6991) );
  NAND2_X1 U8784 ( .A1(n6988), .A2(n6987), .ZN(n6989) );
  NAND2_X1 U8785 ( .A1(n6993), .A2(n6992), .ZN(n12157) );
  NOR2_X1 U8786 ( .A1(n12818), .A2(n7923), .ZN(n7921) );
  NAND2_X1 U8787 ( .A1(n7857), .A2(n7858), .ZN(n12061) );
  INV_X1 U8788 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8978) );
  AND2_X1 U8789 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n8785) );
  NAND2_X1 U8790 ( .A1(n11095), .A2(n6572), .ZN(n11751) );
  NAND2_X1 U8791 ( .A1(n11095), .A2(n12808), .ZN(n11753) );
  NAND2_X1 U8792 ( .A1(n10965), .A2(n11326), .ZN(n11558) );
  NAND2_X1 U8793 ( .A1(n9336), .A2(n11150), .ZN(n11151) );
  NAND2_X1 U8794 ( .A1(n15844), .A2(n12988), .ZN(n12764) );
  NOR2_X1 U8795 ( .A1(n14309), .A2(n7578), .ZN(n7582) );
  NAND2_X1 U8796 ( .A1(n6567), .A2(n9371), .ZN(n7577) );
  NAND2_X1 U8797 ( .A1(n7583), .A2(n9371), .ZN(n7446) );
  NAND2_X1 U8798 ( .A1(n7583), .A2(n7582), .ZN(n14574) );
  AND2_X1 U8799 ( .A1(n9366), .A2(n14395), .ZN(n14365) );
  OR2_X1 U8800 ( .A1(n12979), .A2(n14393), .ZN(n14395) );
  NAND2_X1 U8801 ( .A1(n6999), .A2(n7001), .ZN(n6997) );
  INV_X1 U8802 ( .A(n7000), .ZN(n6999) );
  INV_X1 U8803 ( .A(n14500), .ZN(n14634) );
  INV_X1 U8804 ( .A(n10836), .ZN(n14635) );
  AOI21_X1 U8805 ( .B1(n7744), .B2(n9356), .A(n6675), .ZN(n7743) );
  AND2_X1 U8806 ( .A1(n12959), .A2(n12958), .ZN(n14536) );
  OAI21_X1 U8807 ( .B1(n11548), .B2(n11394), .A(n9348), .ZN(n11396) );
  INV_X1 U8808 ( .A(n12784), .ZN(n15867) );
  AND3_X1 U8809 ( .A1(n10832), .A2(n15864), .A3(n10834), .ZN(n11092) );
  INV_X1 U8810 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9329) );
  INV_X1 U8811 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8816) );
  AND2_X1 U8812 ( .A1(n9109), .A2(n9332), .ZN(n12341) );
  OR2_X1 U8813 ( .A1(n9036), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n9019) );
  AND2_X1 U8814 ( .A1(n7833), .A2(n7832), .ZN(n7835) );
  AND2_X1 U8815 ( .A1(n8775), .A2(n7836), .ZN(n7832) );
  NAND2_X1 U8816 ( .A1(n8811), .A2(n8833), .ZN(n8973) );
  AND2_X1 U8817 ( .A1(n8878), .A2(n8877), .ZN(n10651) );
  OAI21_X1 U8818 ( .B1(n15631), .B2(n9954), .A(n9517), .ZN(n9518) );
  AND2_X1 U8819 ( .A1(n7899), .A2(n7900), .ZN(n7895) );
  INV_X1 U8820 ( .A(n9936), .ZN(n9952) );
  INV_X1 U8821 ( .A(n6830), .ZN(n9749) );
  NAND2_X1 U8822 ( .A1(n6828), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9646) );
  INV_X1 U8823 ( .A(n9611), .ZN(n6828) );
  OR2_X1 U8824 ( .A1(n9646), .A2(n10766), .ZN(n9648) );
  NAND2_X1 U8825 ( .A1(n10184), .A2(n10183), .ZN(n10182) );
  NAND2_X1 U8826 ( .A1(n7303), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9804) );
  NAND2_X1 U8827 ( .A1(n7170), .A2(n7175), .ZN(n14860) );
  NAND2_X1 U8828 ( .A1(n14836), .A2(n7177), .ZN(n7170) );
  NOR2_X1 U8829 ( .A1(n7891), .A2(n7888), .ZN(n7887) );
  INV_X1 U8830 ( .A(n7895), .ZN(n7888) );
  INV_X1 U8831 ( .A(n14788), .ZN(n7891) );
  AOI21_X1 U8832 ( .B1(n7890), .B2(n14788), .A(n6683), .ZN(n7889) );
  INV_X1 U8833 ( .A(n7892), .ZN(n7890) );
  NAND2_X1 U8834 ( .A1(n7304), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9694) );
  INV_X1 U8835 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9445) );
  OR2_X1 U8836 ( .A1(n9694), .A2(n9445), .ZN(n9735) );
  NAND2_X1 U8837 ( .A1(n6827), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9671) );
  INV_X1 U8838 ( .A(n9648), .ZN(n6827) );
  INV_X1 U8839 ( .A(n7304), .ZN(n9692) );
  AOI22_X1 U8840 ( .A1(n11057), .A2(n6543), .B1(n11171), .B2(n9931), .ZN(n9483) );
  OR2_X1 U8841 ( .A1(n9778), .A2(n9777), .ZN(n7900) );
  NAND2_X1 U8842 ( .A1(n11028), .A2(n9559), .ZN(n7880) );
  INV_X1 U8843 ( .A(n7181), .ZN(n7180) );
  NAND2_X1 U8844 ( .A1(n7182), .A2(n6559), .ZN(n7181) );
  NAND2_X1 U8845 ( .A1(n14817), .A2(n7183), .ZN(n7182) );
  NAND2_X1 U8846 ( .A1(n12653), .A2(n6657), .ZN(n7736) );
  NOR2_X1 U8847 ( .A1(n12605), .A2(n12606), .ZN(n7740) );
  NAND2_X1 U8848 ( .A1(n7735), .A2(n7737), .ZN(n7730) );
  NOR2_X1 U8849 ( .A1(n7739), .A2(n7738), .ZN(n7737) );
  INV_X1 U8850 ( .A(n12603), .ZN(n7738) );
  INV_X1 U8851 ( .A(n12602), .ZN(n7739) );
  AND2_X1 U8852 ( .A1(n12651), .A2(n15387), .ZN(n7470) );
  AND4_X1 U8853 ( .A1(n9740), .A2(n9739), .A3(n9738), .A4(n9737), .ZN(n14830)
         );
  AND4_X1 U8854 ( .A1(n9451), .A2(n9450), .A3(n9449), .A4(n9448), .ZN(n14754)
         );
  AND4_X1 U8855 ( .A1(n9699), .A2(n9698), .A3(n9697), .A4(n9696), .ZN(n14873)
         );
  NAND2_X1 U8856 ( .A1(n9987), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9513) );
  NOR2_X1 U8857 ( .A1(n14963), .A2(n7527), .ZN(n14962) );
  NAND2_X1 U8858 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n7527) );
  AND2_X1 U8859 ( .A1(n10588), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7525) );
  INV_X1 U8860 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10766) );
  AND2_X1 U8861 ( .A1(n6875), .A2(n6714), .ZN(n15027) );
  OR2_X1 U8862 ( .A1(n11465), .A2(n6878), .ZN(n6877) );
  OR2_X1 U8863 ( .A1(n11440), .A2(n11438), .ZN(n6878) );
  NOR2_X1 U8864 ( .A1(n11467), .A2(n11466), .ZN(n11465) );
  OR2_X1 U8865 ( .A1(n11446), .A2(n11447), .ZN(n11484) );
  XNOR2_X1 U8866 ( .A(n15046), .B(n15660), .ZN(n15658) );
  INV_X1 U8867 ( .A(n15046), .ZN(n15045) );
  OR2_X1 U8868 ( .A1(n15058), .A2(n15059), .ZN(n15072) );
  OR2_X1 U8869 ( .A1(n9765), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n9780) );
  NOR2_X1 U8870 ( .A1(n13029), .A2(n15128), .ZN(n7966) );
  NAND2_X1 U8871 ( .A1(n9905), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n9944) );
  NAND2_X1 U8872 ( .A1(n7219), .A2(n13070), .ZN(n15142) );
  NAND2_X1 U8873 ( .A1(n7309), .A2(n7265), .ZN(n15218) );
  NOR2_X1 U8874 ( .A1(n7994), .A2(n15437), .ZN(n7309) );
  OR2_X1 U8875 ( .A1(n9804), .A2(n14866), .ZN(n9823) );
  NOR2_X1 U8876 ( .A1(n15285), .A2(n7993), .ZN(n15254) );
  INV_X1 U8877 ( .A(n7995), .ZN(n7993) );
  NOR2_X1 U8878 ( .A1(n15285), .A2(n15455), .ZN(n15270) );
  AND3_X1 U8879 ( .A1(n9791), .A2(n9790), .A3(n9789), .ZN(n14838) );
  INV_X1 U8880 ( .A(n13015), .ZN(n15318) );
  NAND2_X1 U8881 ( .A1(n7192), .A2(n13050), .ZN(n15335) );
  NAND2_X1 U8882 ( .A1(n15339), .A2(n13046), .ZN(n7192) );
  NAND2_X1 U8883 ( .A1(n15335), .A2(n15334), .ZN(n15333) );
  AND4_X1 U8884 ( .A1(n9716), .A2(n9715), .A3(n9714), .A4(n9713), .ZN(n14923)
         );
  NOR2_X1 U8885 ( .A1(n15486), .A2(n7986), .ZN(n7985) );
  NAND2_X1 U8886 ( .A1(n7988), .A2(n7987), .ZN(n15361) );
  NOR2_X1 U8887 ( .A1(n12211), .A2(n7989), .ZN(n15360) );
  NAND2_X1 U8888 ( .A1(n12017), .A2(n12016), .ZN(n12018) );
  NOR2_X1 U8889 ( .A1(n12211), .A2(n14891), .ZN(n12026) );
  INV_X1 U8890 ( .A(n7451), .ZN(n7447) );
  INV_X1 U8891 ( .A(n11569), .ZN(n7449) );
  NAND2_X1 U8892 ( .A1(n9416), .A2(n6671), .ZN(n9592) );
  NAND2_X1 U8893 ( .A1(n9416), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9564) );
  AND2_X1 U8894 ( .A1(n7991), .A2(n11425), .ZN(n11586) );
  INV_X1 U8895 ( .A(n12459), .ZN(n11342) );
  NAND2_X1 U8896 ( .A1(n11425), .A2(n11342), .ZN(n11353) );
  INV_X1 U8897 ( .A(n14922), .ZN(n15637) );
  INV_X1 U8898 ( .A(n7689), .ZN(n12427) );
  NAND2_X1 U8899 ( .A1(n15732), .A2(n11298), .ZN(n11175) );
  NAND3_X1 U8900 ( .A1(n6678), .A2(n7984), .A3(n9498), .ZN(n11186) );
  OR2_X1 U8901 ( .A1(n6626), .A2(n9779), .ZN(n7984) );
  NAND2_X1 U8902 ( .A1(n12426), .A2(n12434), .ZN(n12634) );
  NAND2_X1 U8903 ( .A1(n15678), .A2(n15112), .ZN(n11063) );
  INV_X1 U8904 ( .A(n14913), .ZN(n15636) );
  NAND2_X1 U8905 ( .A1(n9962), .A2(n10227), .ZN(n11059) );
  NAND2_X1 U8906 ( .A1(n7215), .A2(n6605), .ZN(n7214) );
  NAND2_X1 U8907 ( .A1(n15170), .A2(n6632), .ZN(n7216) );
  INV_X1 U8908 ( .A(n7217), .ZN(n7215) );
  NAND2_X1 U8909 ( .A1(n15402), .A2(n15763), .ZN(n7692) );
  INV_X1 U8910 ( .A(n14815), .ZN(n15497) );
  OR2_X1 U8911 ( .A1(n12618), .A2(n15314), .ZN(n15770) );
  OR2_X1 U8912 ( .A1(n11301), .A2(n15112), .ZN(n15745) );
  AND2_X1 U8913 ( .A1(n9477), .A2(n10228), .ZN(n10224) );
  XNOR2_X1 U8914 ( .A(n12611), .B(n12607), .ZN(n13195) );
  NAND2_X1 U8915 ( .A1(n12591), .A2(n12590), .ZN(n12611) );
  OAI21_X1 U8916 ( .B1(n9210), .B2(n7508), .A(n7505), .ZN(n9244) );
  AOI21_X1 U8917 ( .B1(n7507), .B2(n7506), .A(n6767), .ZN(n7505) );
  INV_X1 U8918 ( .A(n7511), .ZN(n7506) );
  XNOR2_X1 U8919 ( .A(n9397), .B(n9396), .ZN(n15649) );
  XNOR2_X1 U8920 ( .A(n9242), .B(n9236), .ZN(n12267) );
  NAND2_X1 U8921 ( .A1(n7509), .A2(n7510), .ZN(n9242) );
  NAND2_X1 U8922 ( .A1(n9210), .A2(n7511), .ZN(n7509) );
  AND2_X1 U8923 ( .A1(n9205), .A2(n9204), .ZN(n11769) );
  AND2_X1 U8924 ( .A1(n6642), .A2(n7065), .ZN(n9107) );
  NAND2_X1 U8925 ( .A1(n7475), .A2(n8744), .ZN(n9093) );
  NAND2_X1 U8926 ( .A1(n7342), .A2(n7477), .ZN(n7475) );
  NAND2_X1 U8927 ( .A1(n9063), .A2(n9075), .ZN(n9077) );
  XNOR2_X1 U8928 ( .A(n9035), .B(n9034), .ZN(n10678) );
  AND2_X1 U8929 ( .A1(n9572), .A2(n9571), .ZN(n9586) );
  AOI21_X1 U8930 ( .B1(n8706), .B2(n8908), .A(n9473), .ZN(n7947) );
  NAND2_X1 U8931 ( .A1(n10532), .A2(n7234), .ZN(n10552) );
  NAND2_X1 U8932 ( .A1(n10543), .A2(n10544), .ZN(n10566) );
  NAND2_X1 U8933 ( .A1(n7667), .A2(n10934), .ZN(n10939) );
  NAND2_X1 U8934 ( .A1(n11730), .A2(n11729), .ZN(n12129) );
  OR2_X1 U8935 ( .A1(n11727), .A2(n11726), .ZN(n11730) );
  AND2_X1 U8936 ( .A1(n7646), .A2(n12126), .ZN(n12131) );
  INV_X1 U8937 ( .A(n7641), .ZN(n7640) );
  OR2_X1 U8938 ( .A1(n7640), .A2(n15613), .ZN(n7639) );
  NAND2_X1 U8939 ( .A1(n15604), .A2(n7645), .ZN(n7641) );
  NAND2_X1 U8940 ( .A1(n8592), .A2(n8609), .ZN(n11260) );
  AND4_X1 U8941 ( .A1(n8332), .A2(n8331), .A3(n8330), .A4(n8329), .ZN(n12332)
         );
  NAND2_X1 U8942 ( .A1(n7026), .A2(n6644), .ZN(n12671) );
  NAND2_X1 U8943 ( .A1(n7027), .A2(n7030), .ZN(n7025) );
  OAI21_X1 U8944 ( .B1(n12229), .B2(n7030), .A(n7027), .ZN(n12329) );
  INV_X1 U8945 ( .A(n7290), .ZN(n7925) );
  AND2_X1 U8946 ( .A1(n8239), .A2(n8238), .ZN(n12178) );
  XNOR2_X1 U8947 ( .A(n11841), .B(n13585), .ZN(n12175) );
  NAND2_X1 U8948 ( .A1(n11601), .A2(n11605), .ZN(n11781) );
  INV_X1 U8949 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n13274) );
  OAI21_X1 U8950 ( .B1(n7274), .B2(n7939), .A(n7034), .ZN(n13271) );
  NAND2_X1 U8951 ( .A1(n8510), .A2(n8509), .ZN(n13908) );
  NAND2_X1 U8952 ( .A1(n7036), .A2(n12676), .ZN(n13301) );
  NAND2_X1 U8953 ( .A1(n11845), .A2(n11844), .ZN(n11847) );
  NAND2_X1 U8954 ( .A1(n13248), .A2(n7938), .ZN(n13311) );
  NAND2_X1 U8955 ( .A1(n13248), .A2(n12685), .ZN(n13310) );
  NAND2_X1 U8956 ( .A1(n8325), .A2(n8324), .ZN(n12245) );
  AND2_X1 U8957 ( .A1(n8397), .A2(n8396), .ZN(n13865) );
  INV_X1 U8958 ( .A(n12332), .ZN(n13580) );
  NAND4_X1 U8959 ( .A1(n8187), .A2(n8186), .A3(n8185), .A4(n8184), .ZN(n13588)
         );
  NAND4_X1 U8960 ( .A1(n8150), .A2(n8149), .A3(n8148), .A4(n8147), .ZN(n13591)
         );
  NAND2_X1 U8961 ( .A1(n8572), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8150) );
  OAI21_X1 U8962 ( .B1(n13717), .B2(n11240), .A(n7329), .ZN(n11216) );
  NAND2_X1 U8963 ( .A1(n13717), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n7329) );
  INV_X1 U8964 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n11217) );
  NAND2_X1 U8965 ( .A1(n13722), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11218) );
  NAND2_X1 U8966 ( .A1(n11290), .A2(n10069), .ZN(n11374) );
  NAND2_X1 U8967 ( .A1(n6821), .A2(n10107), .ZN(n11647) );
  NAND2_X1 U8968 ( .A1(n11615), .A2(n7097), .ZN(n11636) );
  NAND2_X1 U8969 ( .A1(n7557), .A2(n11610), .ZN(n11633) );
  NAND2_X1 U8970 ( .A1(n7072), .A2(n7080), .ZN(n11139) );
  OAI21_X1 U8971 ( .B1(n11618), .B2(n7077), .A(n7074), .ZN(n7073) );
  INV_X1 U8972 ( .A(n7076), .ZN(n7074) );
  AND2_X1 U8973 ( .A1(n10167), .A2(n7080), .ZN(n11140) );
  NAND2_X1 U8974 ( .A1(n10170), .A2(n10076), .ZN(n7625) );
  NAND2_X1 U8975 ( .A1(n10170), .A2(n7631), .ZN(n7630) );
  OAI21_X1 U8976 ( .B1(n10075), .B2(n7627), .A(n7083), .ZN(n10151) );
  NOR2_X1 U8977 ( .A1(n10152), .A2(n10126), .ZN(n11966) );
  NAND2_X1 U8978 ( .A1(n6593), .A2(n10125), .ZN(n6824) );
  NAND2_X1 U8979 ( .A1(n11965), .A2(n6593), .ZN(n6823) );
  NAND2_X1 U8980 ( .A1(n13620), .A2(n13619), .ZN(n13631) );
  NOR2_X1 U8981 ( .A1(n7565), .A2(n10062), .ZN(n13625) );
  NAND2_X1 U8982 ( .A1(n7564), .A2(n7566), .ZN(n13626) );
  OAI21_X1 U8983 ( .B1(n10082), .B2(n7089), .A(n7088), .ZN(n13656) );
  NOR2_X1 U8984 ( .A1(n7090), .A2(n7091), .ZN(n7089) );
  NAND2_X1 U8985 ( .A1(n7090), .A2(n6558), .ZN(n7088) );
  NAND2_X1 U8986 ( .A1(n10131), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7090) );
  AND3_X1 U8987 ( .A1(n7561), .A2(n13663), .A3(P3_REG2_REG_15__SCAN_IN), .ZN(
        n13666) );
  NOR2_X1 U8988 ( .A1(n13677), .A2(n7328), .ZN(n13681) );
  AND2_X1 U8989 ( .A1(n13679), .A2(n13678), .ZN(n7328) );
  NAND2_X1 U8990 ( .A1(n13681), .A2(n13680), .ZN(n13691) );
  NAND2_X1 U8991 ( .A1(n7068), .A2(n7067), .ZN(n13698) );
  OR2_X1 U8992 ( .A1(n13737), .A2(n13733), .ZN(n7549) );
  NAND2_X1 U8993 ( .A1(n7553), .A2(n7552), .ZN(n7551) );
  AND2_X1 U8994 ( .A1(n13737), .A2(n13733), .ZN(n7547) );
  INV_X1 U8995 ( .A(n13753), .ZN(n7622) );
  NAND2_X1 U8996 ( .A1(n8540), .A2(n8554), .ZN(n13225) );
  AOI21_X1 U8997 ( .B1(n12749), .B2(n12708), .A(n12707), .ZN(n12751) );
  NAND2_X1 U8998 ( .A1(n8513), .A2(n8499), .ZN(n13795) );
  AND2_X1 U8999 ( .A1(n7783), .A2(n13500), .ZN(n13794) );
  NAND2_X1 U9000 ( .A1(n7783), .A2(n7781), .ZN(n13792) );
  NAND2_X1 U9001 ( .A1(n13800), .A2(n7408), .ZN(n7783) );
  AND2_X1 U9002 ( .A1(n7410), .A2(n6616), .ZN(n13789) );
  NAND2_X1 U9003 ( .A1(n7410), .A2(n7409), .ZN(n13787) );
  NAND2_X1 U9004 ( .A1(n13860), .A2(n8661), .ZN(n13846) );
  NAND2_X1 U9005 ( .A1(n8420), .A2(n8419), .ZN(n13874) );
  OAI21_X1 U9006 ( .B1(n11758), .B2(n11757), .A(n13442), .ZN(n11918) );
  NAND2_X1 U9007 ( .A1(n8232), .A2(n8231), .ZN(n15949) );
  AOI22_X1 U9008 ( .A1(n8568), .A2(n10502), .B1(n8418), .B2(n11145), .ZN(n8231) );
  INV_X1 U9009 ( .A(n13880), .ZN(n13852) );
  AND2_X1 U9010 ( .A1(n6893), .A2(n6894), .ZN(n11510) );
  AND2_X1 U9011 ( .A1(n7774), .A2(n7773), .ZN(n6895) );
  AOI21_X1 U9012 ( .B1(n11523), .B2(n11524), .A(n13426), .ZN(n11500) );
  NAND2_X1 U9013 ( .A1(n7775), .A2(n7774), .ZN(n11499) );
  INV_X2 U9014 ( .A(n15903), .ZN(n15921) );
  INV_X1 U9015 ( .A(n15923), .ZN(n15901) );
  INV_X1 U9016 ( .A(n13942), .ZN(n13940) );
  NAND2_X1 U9017 ( .A1(n13371), .A2(n13370), .ZN(n13968) );
  XNOR2_X1 U9018 ( .A(n10041), .B(n13521), .ZN(n13192) );
  INV_X1 U9019 ( .A(n13229), .ZN(n12746) );
  NAND2_X1 U9020 ( .A1(n8485), .A2(n8484), .ZN(n13984) );
  NAND2_X1 U9021 ( .A1(n8468), .A2(n8467), .ZN(n13990) );
  INV_X1 U9022 ( .A(n13831), .ZN(n13998) );
  OAI21_X1 U9023 ( .B1(n8381), .B2(n12386), .A(n13474), .ZN(n13878) );
  NAND2_X1 U9024 ( .A1(n8375), .A2(n8374), .ZN(n13476) );
  NAND2_X1 U9025 ( .A1(n8342), .A2(n8341), .ZN(n13356) );
  AND2_X1 U9026 ( .A1(n7789), .A2(n8315), .ZN(n12244) );
  NAND2_X1 U9027 ( .A1(n8646), .A2(n8645), .ZN(n12242) );
  NAND2_X1 U9028 ( .A1(n7794), .A2(n7795), .ZN(n11893) );
  NAND2_X1 U9029 ( .A1(n11758), .A2(n7796), .ZN(n7794) );
  NAND2_X1 U9030 ( .A1(n8597), .A2(n8596), .ZN(n14024) );
  OR2_X1 U9031 ( .A1(n10783), .A2(P3_D_REG_1__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U9032 ( .A1(n6548), .A2(P3_D_REG_0__SCAN_IN), .ZN(n7369) );
  AND2_X1 U9033 ( .A1(n11259), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14026) );
  NAND4_X1 U9034 ( .A1(n6918), .A2(n8106), .A3(n6535), .A4(n8114), .ZN(n8119)
         );
  INV_X1 U9035 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n6919) );
  NAND2_X1 U9036 ( .A1(n13365), .A2(n7597), .ZN(n13373) );
  OR2_X1 U9037 ( .A1(n13008), .A2(n13007), .ZN(n7597) );
  OR2_X1 U9038 ( .A1(n8566), .A2(n8565), .ZN(n8567) );
  NAND2_X1 U9039 ( .A1(n7617), .A2(n7619), .ZN(n8548) );
  NAND2_X1 U9040 ( .A1(n8523), .A2(n7620), .ZN(n7617) );
  OR2_X1 U9041 ( .A1(n8523), .A2(n8522), .ZN(n7618) );
  INV_X1 U9042 ( .A(SI_23_), .ZN(n11414) );
  XNOR2_X1 U9043 ( .A(n8616), .B(n7943), .ZN(n11128) );
  NAND2_X1 U9044 ( .A1(n8617), .A2(n7944), .ZN(n8615) );
  INV_X1 U9045 ( .A(SI_21_), .ZN(n11453) );
  NAND2_X1 U9046 ( .A1(n7351), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8622) );
  NAND2_X1 U9047 ( .A1(n8617), .A2(n8619), .ZN(n7351) );
  NAND2_X1 U9048 ( .A1(n8618), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8620) );
  INV_X1 U9049 ( .A(SI_19_), .ZN(n10929) );
  INV_X1 U9050 ( .A(SI_17_), .ZN(n10871) );
  INV_X1 U9051 ( .A(SI_16_), .ZN(n10824) );
  XNOR2_X1 U9052 ( .A(n8384), .B(n8382), .ZN(n10822) );
  NAND2_X1 U9053 ( .A1(n8371), .A2(n8370), .ZN(n8384) );
  INV_X1 U9054 ( .A(SI_15_), .ZN(n10754) );
  INV_X1 U9055 ( .A(SI_12_), .ZN(n10617) );
  NAND2_X1 U9056 ( .A1(n7599), .A2(n8273), .ZN(n8288) );
  NAND2_X1 U9057 ( .A1(n8272), .A2(n8271), .ZN(n7599) );
  NAND2_X1 U9058 ( .A1(n8253), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6921) );
  INV_X1 U9059 ( .A(n7085), .ZN(n7084) );
  NAND2_X1 U9060 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n7086) );
  NAND2_X1 U9061 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n7355) );
  INV_X1 U9062 ( .A(n6976), .ZN(n6975) );
  NOR2_X1 U9063 ( .A1(n6977), .A2(n11668), .ZN(n6976) );
  AOI21_X1 U9064 ( .B1(n14090), .B2(n7823), .A(n6579), .ZN(n6979) );
  NAND2_X1 U9065 ( .A1(n12184), .A2(n12183), .ZN(n13088) );
  NAND2_X1 U9066 ( .A1(n7820), .A2(n7819), .ZN(n10862) );
  NAND2_X1 U9067 ( .A1(n7816), .A2(n7817), .ZN(n10863) );
  INV_X1 U9068 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n14081) );
  NAND2_X1 U9069 ( .A1(n14130), .A2(n13157), .ZN(n14100) );
  NAND2_X1 U9070 ( .A1(n12734), .A2(n10216), .ZN(n7844) );
  INV_X1 U9071 ( .A(n12795), .ZN(n15873) );
  NAND2_X1 U9072 ( .A1(n7830), .A2(n7831), .ZN(n11228) );
  OR2_X1 U9073 ( .A1(n11038), .A2(n11037), .ZN(n7831) );
  NAND2_X1 U9074 ( .A1(n12143), .A2(n12144), .ZN(n12184) );
  INV_X1 U9075 ( .A(n7347), .ZN(n14140) );
  NAND2_X1 U9076 ( .A1(n14087), .A2(n13103), .ZN(n14151) );
  INV_X1 U9077 ( .A(n13149), .ZN(n7291) );
  AND2_X1 U9078 ( .A1(n10847), .A2(n10840), .ZN(n14161) );
  INV_X1 U9079 ( .A(n14196), .ZN(n14206) );
  NAND2_X1 U9080 ( .A1(n14122), .A2(n13125), .ZN(n14182) );
  NAND2_X1 U9081 ( .A1(n11245), .A2(n11244), .ZN(n11669) );
  AND2_X1 U9082 ( .A1(n10625), .A2(n10638), .ZN(n14192) );
  NAND2_X1 U9083 ( .A1(n8046), .A2(n8045), .ZN(n8040) );
  NAND2_X1 U9084 ( .A1(n8044), .A2(n8052), .ZN(n8046) );
  INV_X1 U9085 ( .A(n12954), .ZN(n8052) );
  NAND2_X1 U9086 ( .A1(n8045), .A2(n12955), .ZN(n8041) );
  INV_X1 U9087 ( .A(n12993), .ZN(n8047) );
  INV_X1 U9088 ( .A(n14166), .ZN(n14223) );
  INV_X1 U9089 ( .A(n14165), .ZN(n14225) );
  OR2_X1 U9090 ( .A1(n8891), .A2(n8869), .ZN(n8874) );
  OR2_X1 U9091 ( .A1(n8961), .A2(n14248), .ZN(n8893) );
  NAND2_X1 U9092 ( .A1(n10644), .A2(n14254), .ZN(n14264) );
  NOR2_X1 U9093 ( .A1(n14259), .A2(n14258), .ZN(n14276) );
  NAND2_X1 U9094 ( .A1(n15816), .A2(n15817), .ZN(n15814) );
  AND2_X1 U9095 ( .A1(n8928), .A2(n8939), .ZN(n10730) );
  OAI22_X1 U9096 ( .A1(n10726), .A2(n10725), .B1(n10624), .B2(n10623), .ZN(
        n10682) );
  AND2_X1 U9097 ( .A1(n15835), .A2(n10808), .ZN(n10812) );
  OAI22_X1 U9098 ( .A1(n10897), .A2(n10896), .B1(n10895), .B2(n10894), .ZN(
        n10898) );
  XNOR2_X1 U9099 ( .A(n11654), .B(n11656), .ZN(n11652) );
  XNOR2_X1 U9100 ( .A(n11980), .B(n11661), .ZN(n11978) );
  NAND2_X1 U9101 ( .A1(n12191), .A2(n12192), .ZN(n12190) );
  OAI22_X1 U9102 ( .A1(n12194), .A2(n12193), .B1(n11975), .B2(n14632), .ZN(
        n12343) );
  NAND2_X1 U9103 ( .A1(n7042), .A2(n7045), .ZN(n12336) );
  OR2_X1 U9104 ( .A1(n12191), .A2(n7047), .ZN(n7042) );
  OR2_X1 U9105 ( .A1(n12340), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n14293) );
  OAI211_X1 U9106 ( .C1(n12755), .C2(n7913), .A(n12754), .B(n10836), .ZN(
        n14572) );
  INV_X1 U9107 ( .A(n12926), .ZN(n12925) );
  INV_X1 U9108 ( .A(n14585), .ZN(n14346) );
  OAI21_X1 U9109 ( .B1(n14378), .B2(n7062), .A(n7415), .ZN(n14336) );
  NAND2_X1 U9110 ( .A1(n7871), .A2(n7872), .ZN(n14387) );
  AND2_X1 U9111 ( .A1(n7875), .A2(n7877), .ZN(n14412) );
  NAND2_X1 U9112 ( .A1(n14425), .A2(n14424), .ZN(n7875) );
  AND2_X1 U9113 ( .A1(n7126), .A2(n7129), .ZN(n14440) );
  NAND2_X1 U9114 ( .A1(n14450), .A2(n9136), .ZN(n7126) );
  NAND2_X1 U9115 ( .A1(n14463), .A2(n7440), .ZN(n14453) );
  AND3_X1 U9116 ( .A1(n7120), .A2(n7118), .A3(n6621), .ZN(n14483) );
  NAND2_X1 U9117 ( .A1(n7846), .A2(n6556), .ZN(n14502) );
  NAND2_X1 U9118 ( .A1(n9052), .A2(n9053), .ZN(n14512) );
  OAI21_X1 U9119 ( .B1(n11362), .B2(n7436), .A(n7434), .ZN(n12059) );
  NAND2_X1 U9120 ( .A1(n11361), .A2(n9351), .ZN(n12057) );
  NAND2_X1 U9121 ( .A1(n14366), .A2(n7007), .ZN(n14353) );
  AND2_X1 U9122 ( .A1(n14366), .A2(n9367), .ZN(n14355) );
  NAND2_X1 U9123 ( .A1(n6998), .A2(n7439), .ZN(n14438) );
  NAND2_X1 U9124 ( .A1(n14487), .A2(n7002), .ZN(n6998) );
  OR2_X1 U9125 ( .A1(n14537), .A2(n9356), .ZN(n7745) );
  INV_X1 U9126 ( .A(n15857), .ZN(n15858) );
  AND2_X1 U9127 ( .A1(n10833), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15864) );
  INV_X1 U9128 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n13078) );
  INV_X1 U9129 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8795) );
  INV_X1 U9130 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n12221) );
  XNOR2_X1 U9131 ( .A(n9310), .B(n8779), .ZN(n12223) );
  XNOR2_X1 U9132 ( .A(n9308), .B(P2_IR_REG_24__SCAN_IN), .ZN(n11768) );
  INV_X1 U9133 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11770) );
  INV_X1 U9134 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11132) );
  INV_X1 U9135 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10891) );
  INV_X1 U9136 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10760) );
  INV_X1 U9137 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10711) );
  INV_X1 U9138 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10755) );
  INV_X1 U9139 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10785) );
  INV_X1 U9140 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10707) );
  INV_X1 U9141 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10620) );
  INV_X1 U9142 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10493) );
  NOR2_X1 U9143 ( .A1(n10481), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13080) );
  INV_X1 U9144 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10498) );
  INV_X1 U9145 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10213) );
  XNOR2_X1 U9146 ( .A(n8835), .B(n8834), .ZN(n14277) );
  OAI211_X1 U9147 ( .C1(n8848), .C2(n7051), .A(n8860), .B(n7050), .ZN(n14262)
         );
  NAND2_X1 U9148 ( .A1(n7051), .A2(n8780), .ZN(n7050) );
  INV_X1 U9149 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10595) );
  NAND2_X1 U9150 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n8896) );
  OR2_X1 U9151 ( .A1(n10187), .A2(P1_U3086), .ZN(n10047) );
  NAND2_X1 U9152 ( .A1(n7169), .A2(n11115), .ZN(n12001) );
  NAND2_X1 U9153 ( .A1(n7905), .A2(n6563), .ZN(n14744) );
  INV_X1 U9154 ( .A(n7188), .ZN(n7187) );
  AOI21_X1 U9155 ( .B1(n7186), .B2(n7188), .A(n6687), .ZN(n7185) );
  NAND3_X1 U9156 ( .A1(n7878), .A2(n9507), .A3(n9524), .ZN(n15642) );
  NAND2_X1 U9157 ( .A1(n14789), .A2(n14788), .ZN(n14787) );
  NAND2_X1 U9158 ( .A1(n7894), .A2(n7892), .ZN(n14789) );
  NAND2_X1 U9159 ( .A1(n14836), .A2(n7895), .ZN(n7894) );
  NAND2_X1 U9160 ( .A1(n7903), .A2(n7901), .ZN(n9983) );
  NAND2_X1 U9161 ( .A1(n6704), .A2(n7902), .ZN(n7901) );
  NAND2_X1 U9162 ( .A1(n11999), .A2(n9603), .ZN(n11866) );
  NAND2_X1 U9163 ( .A1(n10182), .A2(n7359), .ZN(n12725) );
  NAND2_X1 U9164 ( .A1(n7360), .A2(n10789), .ZN(n7359) );
  INV_X1 U9165 ( .A(n10183), .ZN(n7360) );
  INV_X1 U9166 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n14801) );
  NAND2_X1 U9167 ( .A1(n14808), .A2(n14807), .ZN(n14806) );
  INV_X1 U9168 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14866) );
  NAND2_X1 U9169 ( .A1(n7174), .A2(n7889), .ZN(n14862) );
  NAND2_X1 U9170 ( .A1(n14836), .A2(n7887), .ZN(n7174) );
  AND2_X1 U9171 ( .A1(n14806), .A2(n7188), .ZN(n14870) );
  NAND2_X1 U9172 ( .A1(n14806), .A2(n9703), .ZN(n14871) );
  NAND2_X1 U9173 ( .A1(n14795), .A2(n9832), .ZN(n14881) );
  NAND2_X1 U9174 ( .A1(n7896), .A2(n7900), .ZN(n14903) );
  OR2_X1 U9175 ( .A1(n14836), .A2(n14837), .ZN(n7896) );
  NAND2_X1 U9176 ( .A1(n7880), .A2(n9562), .ZN(n11117) );
  NAND2_X1 U9177 ( .A1(n9723), .A2(n12614), .ZN(n9733) );
  INV_X1 U9178 ( .A(n13025), .ZN(n14935) );
  INV_X1 U9179 ( .A(n13069), .ZN(n14937) );
  OAI21_X1 U9180 ( .B1(n15229), .B2(n9907), .A(n9828), .ZN(n14942) );
  INV_X1 U9181 ( .A(n14838), .ZN(n14945) );
  NAND2_X1 U9182 ( .A1(n9773), .A2(n9772), .ZN(n14946) );
  INV_X1 U9183 ( .A(n14754), .ZN(n14949) );
  NAND2_X1 U9184 ( .A1(n9513), .A2(n6617), .ZN(n14957) );
  NAND2_X1 U9185 ( .A1(n7524), .A2(n10575), .ZN(n14995) );
  NOR2_X1 U9186 ( .A1(n7516), .A2(n7515), .ZN(n10577) );
  NAND2_X1 U9187 ( .A1(n7521), .A2(n7517), .ZN(n7516) );
  INV_X1 U9188 ( .A(n7520), .ZN(n7515) );
  INV_X1 U9189 ( .A(n7525), .ZN(n7517) );
  NAND2_X1 U9190 ( .A1(n6861), .A2(n6859), .ZN(n10762) );
  NAND2_X1 U9191 ( .A1(n6862), .A2(n6860), .ZN(n6859) );
  INV_X1 U9192 ( .A(n10599), .ZN(n6860) );
  AND2_X1 U9193 ( .A1(n15015), .A2(n15014), .ZN(n15016) );
  NOR2_X1 U9194 ( .A1(n15016), .A2(n7537), .ZN(n10765) );
  NOR2_X1 U9195 ( .A1(n10771), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7537) );
  INV_X1 U9196 ( .A(n6875), .ZN(n15030) );
  NOR2_X1 U9197 ( .A1(n15027), .A2(n6874), .ZN(n11437) );
  OR2_X1 U9198 ( .A1(n10912), .A2(n10914), .ZN(n6874) );
  INV_X1 U9199 ( .A(n6877), .ZN(n11477) );
  INV_X1 U9200 ( .A(n7540), .ZN(n15042) );
  AND2_X1 U9201 ( .A1(n10190), .A2(n7686), .ZN(n15651) );
  AND2_X1 U9202 ( .A1(n15070), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6870) );
  INV_X1 U9203 ( .A(n15111), .ZN(n15665) );
  NOR2_X1 U9204 ( .A1(n7997), .A2(n15121), .ZN(n7996) );
  XNOR2_X1 U9205 ( .A(n7272), .B(n7271), .ZN(n15403) );
  INV_X1 U9206 ( .A(n15129), .ZN(n7271) );
  INV_X1 U9207 ( .A(n15128), .ZN(n7300) );
  XNOR2_X1 U9208 ( .A(n6843), .B(n7458), .ZN(n6842) );
  NAND2_X1 U9209 ( .A1(n15170), .A2(n13068), .ZN(n6843) );
  NAND2_X1 U9210 ( .A1(n7456), .A2(n7975), .ZN(n15155) );
  NAND2_X1 U9211 ( .A1(n15211), .A2(n7459), .ZN(n7456) );
  INV_X1 U9212 ( .A(n14822), .ZN(n15417) );
  NAND2_X1 U9213 ( .A1(n7981), .A2(n7979), .ZN(n15168) );
  NAND2_X1 U9214 ( .A1(n15199), .A2(n13024), .ZN(n15183) );
  NAND2_X1 U9215 ( .A1(n15215), .A2(n13064), .ZN(n15202) );
  AND2_X1 U9216 ( .A1(n15211), .A2(n13022), .ZN(n15200) );
  NOR2_X1 U9217 ( .A1(n7712), .A2(n7711), .ZN(n8099) );
  INV_X1 U9218 ( .A(n13061), .ZN(n7711) );
  NAND2_X1 U9219 ( .A1(n7949), .A2(n7950), .ZN(n15228) );
  NAND2_X1 U9220 ( .A1(n7957), .A2(n7951), .ZN(n15243) );
  NAND2_X1 U9221 ( .A1(n6869), .A2(n13020), .ZN(n15279) );
  NAND2_X1 U9222 ( .A1(n15297), .A2(n13019), .ZN(n6869) );
  OR2_X1 U9223 ( .A1(n7694), .A2(n7697), .ZN(n11581) );
  INV_X1 U9224 ( .A(n7695), .ZN(n7694) );
  AND2_X1 U9225 ( .A1(n7452), .A2(n7450), .ZN(n11948) );
  OR2_X1 U9226 ( .A1(n11578), .A2(n11577), .ZN(n7696) );
  AOI21_X1 U9227 ( .B1(n11194), .B2(n15707), .A(n12428), .ZN(n11424) );
  NOR2_X2 U9228 ( .A1(n6546), .A2(n11067), .ZN(n15716) );
  NAND2_X1 U9229 ( .A1(n15404), .A2(n15738), .ZN(n15406) );
  NAND2_X1 U9230 ( .A1(n10224), .A2(n10795), .ZN(n15729) );
  OAI22_X1 U9231 ( .A1(n7483), .A2(n7482), .B1(n12613), .B2(n7485), .ZN(n7481)
         );
  NAND2_X1 U9232 ( .A1(n15544), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9421) );
  INV_X1 U9233 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n12219) );
  INV_X1 U9234 ( .A(n9959), .ZN(n11774) );
  INV_X1 U9235 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11113) );
  NAND2_X1 U9236 ( .A1(n9434), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7268) );
  NAND2_X1 U9237 ( .A1(n9140), .A2(n7572), .ZN(n12408) );
  INV_X1 U9238 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10890) );
  INV_X1 U9239 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10759) );
  INV_X1 U9240 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10709) );
  INV_X1 U9241 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10787) );
  AND2_X1 U9242 ( .A1(n9687), .A2(n9708), .ZN(n11471) );
  XNOR2_X1 U9243 ( .A(n9627), .B(P1_IR_REG_10__SCAN_IN), .ZN(n15037) );
  INV_X1 U9244 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10514) );
  INV_X1 U9245 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10490) );
  NAND2_X1 U9246 ( .A1(n9514), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9515) );
  NAND2_X1 U9247 ( .A1(n7528), .A2(n9496), .ZN(n10488) );
  INV_X1 U9248 ( .A(n7529), .ZN(n7528) );
  OAI21_X1 U9249 ( .B1(n9455), .B2(n7531), .A(n7530), .ZN(n7529) );
  INV_X1 U9250 ( .A(P1_RD_REG_SCAN_IN), .ZN(n10207) );
  NAND2_X1 U9251 ( .A1(n7663), .A2(n10538), .ZN(n7662) );
  XNOR2_X1 U9252 ( .A(n10939), .B(P2_ADDR_REG_6__SCAN_IN), .ZN(n15554) );
  XNOR2_X1 U9253 ( .A(n10951), .B(n10943), .ZN(n15556) );
  NAND2_X1 U9254 ( .A1(n15558), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n11725) );
  NAND2_X1 U9255 ( .A1(n7665), .A2(n12289), .ZN(n15562) );
  XNOR2_X1 U9256 ( .A(n15568), .B(n12295), .ZN(n15560) );
  NAND2_X1 U9257 ( .A1(n15593), .A2(n15592), .ZN(n15596) );
  AND2_X1 U9258 ( .A1(n6636), .A2(n7656), .ZN(n15597) );
  NAND2_X1 U9259 ( .A1(n7009), .A2(n13270), .ZN(P3_U3160) );
  NAND2_X1 U9260 ( .A1(n6596), .A2(n13325), .ZN(n7934) );
  NAND2_X1 U9261 ( .A1(n13239), .A2(n11810), .ZN(n12078) );
  OAI21_X1 U9262 ( .B1(n13401), .B2(n13400), .A(n13399), .ZN(n7803) );
  AND2_X1 U9263 ( .A1(n13705), .A2(n13704), .ZN(n6797) );
  AND2_X1 U9264 ( .A1(n13732), .A2(n13731), .ZN(n6922) );
  OAI21_X1 U9265 ( .B1(n13901), .B2(n13894), .A(n6766), .ZN(n6883) );
  OAI211_X1 U9266 ( .C1(n13899), .C2(n15973), .A(n13904), .B(n6758), .ZN(
        P3_U3488) );
  NAND2_X1 U9267 ( .A1(n8690), .A2(n7366), .ZN(n7365) );
  OAI21_X1 U9268 ( .B1(n13975), .B2(n15960), .A(n7424), .ZN(P3_U3453) );
  INV_X1 U9269 ( .A(n7425), .ZN(n7424) );
  OAI21_X1 U9270 ( .B1(n13979), .B2(n14021), .A(n6759), .ZN(n7425) );
  AND2_X1 U9271 ( .A1(n7258), .A2(n7837), .ZN(n14199) );
  NAND2_X1 U9272 ( .A1(n7337), .A2(n14299), .ZN(n7336) );
  NAND2_X1 U9273 ( .A1(n15890), .A2(n10458), .ZN(n7350) );
  NAND2_X1 U9274 ( .A1(n7319), .A2(n11417), .ZN(n7318) );
  NAND2_X1 U9275 ( .A1(n15890), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n7109) );
  OAI21_X1 U9276 ( .B1(n12723), .B2(n14734), .A(n9374), .ZN(P2_U3496) );
  OR2_X1 U9277 ( .A1(n15886), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7423) );
  NAND2_X1 U9278 ( .A1(n7319), .A2(n11419), .ZN(n7320) );
  OAI21_X1 U9279 ( .B1(n7377), .B2(n15634), .A(n14823), .ZN(P1_U3225) );
  XNOR2_X1 U9280 ( .A(n14816), .B(n7907), .ZN(n7377) );
  NOR2_X1 U9281 ( .A1(n7372), .A2(n7371), .ZN(n7370) );
  NOR2_X1 U9282 ( .A1(n15410), .A2(n14918), .ZN(n7371) );
  OR2_X1 U9283 ( .A1(n12665), .A2(n12664), .ZN(n7295) );
  NAND2_X1 U9284 ( .A1(n7534), .A2(n15314), .ZN(n7533) );
  INV_X1 U9285 ( .A(n7962), .ZN(n15397) );
  NAND2_X1 U9286 ( .A1(n15789), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7958) );
  NAND2_X1 U9287 ( .A1(n15789), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7453) );
  NAND2_X1 U9288 ( .A1(n10934), .A2(n7666), .ZN(n10935) );
  INV_X1 U9289 ( .A(n7667), .ZN(n7666) );
  NAND2_X1 U9290 ( .A1(n7238), .A2(n11714), .ZN(n11715) );
  NAND2_X1 U9291 ( .A1(n7257), .A2(n11714), .ZN(n10963) );
  NAND2_X1 U9292 ( .A1(n15575), .A2(n7655), .ZN(n15584) );
  OR2_X1 U9293 ( .A1(n15576), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7655) );
  NAND2_X1 U9294 ( .A1(n7245), .A2(n7267), .ZN(n15614) );
  AND2_X1 U9295 ( .A1(n7633), .A2(n7266), .ZN(n7245) );
  OAI211_X1 U9296 ( .C1(n7244), .C2(n15618), .A(n7243), .B(n7242), .ZN(
        SUB_1596_U4) );
  NAND2_X1 U9297 ( .A1(n15617), .A2(n7247), .ZN(n7243) );
  NAND2_X1 U9298 ( .A1(n6584), .A2(n7267), .ZN(n7242) );
  INV_X1 U9299 ( .A(n11145), .ZN(n7077) );
  AND2_X1 U9300 ( .A1(n8007), .A2(n13498), .ZN(n6555) );
  OR2_X1 U9301 ( .A1(n12850), .A2(n14232), .ZN(n6556) );
  AND4_X1 U9302 ( .A1(n6960), .A2(n6586), .A3(n14536), .A4(n14550), .ZN(n6557)
         );
  NAND2_X1 U9303 ( .A1(n13810), .A2(n13805), .ZN(n7672) );
  OR2_X1 U9304 ( .A1(n7624), .A2(n7091), .ZN(n6558) );
  OR2_X1 U9305 ( .A1(n13984), .A2(n13497), .ZN(n13500) );
  INV_X1 U9306 ( .A(n8706), .ZN(n8712) );
  OR2_X1 U9307 ( .A1(n9902), .A2(n9901), .ZN(n6559) );
  AND2_X1 U9308 ( .A1(n14631), .A2(n14205), .ZN(n6560) );
  AND2_X1 U9309 ( .A1(n13590), .A2(n13243), .ZN(n6561) );
  AND2_X1 U9310 ( .A1(n15585), .A2(n15586), .ZN(n6562) );
  AND2_X1 U9311 ( .A1(n7908), .A2(n9920), .ZN(n6563) );
  AND2_X1 U9312 ( .A1(n9819), .A2(n9820), .ZN(n6564) );
  INV_X1 U9313 ( .A(n7627), .ZN(n7626) );
  OAI22_X1 U9314 ( .A1(n7631), .A2(n12154), .B1(n10076), .B2(n7632), .ZN(n7627) );
  INV_X1 U9315 ( .A(n7939), .ZN(n7938) );
  NAND2_X1 U9316 ( .A1(n7940), .A2(n12685), .ZN(n7939) );
  NAND2_X1 U9317 ( .A1(n8757), .A2(n10929), .ZN(n6565) );
  AND2_X1 U9318 ( .A1(n7500), .A2(n9153), .ZN(n6566) );
  NOR2_X1 U9319 ( .A1(n14582), .A2(n14101), .ZN(n6567) );
  NOR2_X1 U9320 ( .A1(n12816), .A2(n12817), .ZN(n6568) );
  OR2_X2 U9321 ( .A1(n13708), .A2(n13707), .ZN(n6569) );
  AND4_X1 U9322 ( .A1(n8984), .A2(n8983), .A3(n8982), .A4(n8981), .ZN(n12820)
         );
  AND2_X1 U9323 ( .A1(n11610), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n6570) );
  OAI21_X1 U9324 ( .B1(n7639), .B2(n7644), .A(n7638), .ZN(n7637) );
  XNOR2_X1 U9325 ( .A(n15163), .B(n13069), .ZN(n15156) );
  AND2_X1 U9326 ( .A1(n14634), .A2(n7919), .ZN(n6571) );
  AND2_X1 U9327 ( .A1(n12808), .A2(n7924), .ZN(n6572) );
  INV_X1 U9328 ( .A(n8749), .ZN(n7474) );
  OR2_X1 U9329 ( .A1(n12764), .A2(n12763), .ZN(n12806) );
  INV_X1 U9330 ( .A(n13551), .ZN(n7408) );
  NAND2_X1 U9331 ( .A1(n9039), .A2(n9038), .ZN(n14653) );
  INV_X1 U9332 ( .A(n14653), .ZN(n7108) );
  XOR2_X1 U9333 ( .A(n6745), .B(n7935), .Z(n6573) );
  OAI211_X1 U9334 ( .C1(n9262), .C2(n6768), .A(n7481), .B(n7479), .ZN(n12735)
         );
  AND4_X1 U9335 ( .A1(n9387), .A2(n9386), .A3(n9385), .A4(n9384), .ZN(n6574)
         );
  XNOR2_X1 U9336 ( .A(n7268), .B(n9413), .ZN(n11112) );
  AND2_X1 U9337 ( .A1(n7909), .A2(n14420), .ZN(n6575) );
  AND2_X1 U9338 ( .A1(n13719), .A2(n13718), .ZN(n6576) );
  AND2_X1 U9339 ( .A1(n12224), .A2(n13583), .ZN(n6577) );
  NOR2_X1 U9340 ( .A1(n12850), .A2(n14203), .ZN(n6578) );
  INV_X1 U9341 ( .A(n15400), .ZN(n15135) );
  AND2_X1 U9342 ( .A1(n9940), .A2(n9939), .ZN(n15400) );
  AND2_X1 U9343 ( .A1(n13105), .A2(n13104), .ZN(n6579) );
  INV_X1 U9344 ( .A(n13406), .ZN(n7791) );
  INV_X1 U9345 ( .A(n14576), .ZN(n14307) );
  NAND2_X1 U9346 ( .A1(n9239), .A2(n9238), .ZN(n14576) );
  AND2_X1 U9347 ( .A1(n10481), .A2(SI_1_), .ZN(n6580) );
  INV_X1 U9348 ( .A(n12818), .ZN(n12816) );
  NAND2_X1 U9349 ( .A1(n8992), .A2(n8991), .ZN(n12818) );
  NAND2_X1 U9350 ( .A1(n10166), .A2(n6749), .ZN(n6581) );
  AND2_X1 U9351 ( .A1(n7491), .A2(n7059), .ZN(n6582) );
  NAND2_X1 U9352 ( .A1(n13534), .A2(n6727), .ZN(n6583) );
  AND3_X1 U9353 ( .A1(n7266), .A2(n7633), .A3(n6725), .ZN(n6584) );
  NAND2_X1 U9354 ( .A1(n7635), .A2(n6629), .ZN(n15616) );
  NAND2_X1 U9355 ( .A1(n6614), .A2(n8050), .ZN(n8049) );
  INV_X1 U9356 ( .A(n8049), .ZN(n8044) );
  INV_X1 U9357 ( .A(n14615), .ZN(n7128) );
  AND2_X1 U9358 ( .A1(n7863), .A2(n6966), .ZN(n6585) );
  INV_X1 U9359 ( .A(n12899), .ZN(n8039) );
  AND2_X1 U9360 ( .A1(n9001), .A2(n12975), .ZN(n6586) );
  INV_X1 U9361 ( .A(n15671), .ZN(n15675) );
  INV_X1 U9362 ( .A(n15675), .ZN(n7700) );
  AND3_X1 U9363 ( .A1(n8028), .A2(n13869), .A3(n8656), .ZN(n6587) );
  OR2_X1 U9364 ( .A1(n15572), .A2(n6562), .ZN(n6588) );
  INV_X1 U9365 ( .A(n14222), .ZN(n7417) );
  AND3_X1 U9366 ( .A1(n6548), .A2(P3_B_REG_SCAN_IN), .A3(n12123), .ZN(n6589)
         );
  INV_X1 U9367 ( .A(n12560), .ZN(n7764) );
  NAND2_X1 U9368 ( .A1(n8868), .A2(n8917), .ZN(n12963) );
  NAND2_X1 U9369 ( .A1(n13525), .A2(n13524), .ZN(n6590) );
  NAND2_X1 U9370 ( .A1(n12732), .A2(n12731), .ZN(n12985) );
  INV_X1 U9371 ( .A(n12985), .ZN(n7913) );
  NOR2_X1 U9372 ( .A1(n8648), .A2(n7402), .ZN(n7401) );
  AND2_X1 U9373 ( .A1(n6699), .A2(n6885), .ZN(n6591) );
  INV_X1 U9374 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9422) );
  INV_X1 U9375 ( .A(n11964), .ZN(n7353) );
  AND2_X1 U9376 ( .A1(n8689), .A2(n8688), .ZN(n15960) );
  AND2_X1 U9377 ( .A1(n11095), .A2(n7922), .ZN(n6592) );
  INV_X1 U9378 ( .A(n11317), .ZN(n7632) );
  NAND2_X1 U9379 ( .A1(n10128), .A2(n7353), .ZN(n6593) );
  AND2_X1 U9380 ( .A1(n10811), .A2(n10808), .ZN(n6594) );
  XNOR2_X1 U9381 ( .A(n9208), .B(SI_25_), .ZN(n9209) );
  AND2_X1 U9382 ( .A1(n6773), .A2(n7775), .ZN(n6595) );
  AND2_X1 U9383 ( .A1(n8491), .A2(n8490), .ZN(n13497) );
  XOR2_X1 U9384 ( .A(n6745), .B(n7936), .Z(n6596) );
  AND2_X1 U9385 ( .A1(n9167), .A2(n8763), .ZN(n6597) );
  INV_X1 U9386 ( .A(n13678), .ZN(n7380) );
  INV_X1 U9387 ( .A(n10744), .ZN(n7091) );
  AND2_X1 U9388 ( .A1(n13664), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n6598) );
  OR2_X1 U9389 ( .A1(n8360), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n6599) );
  INV_X1 U9390 ( .A(n7771), .ZN(n15631) );
  NAND2_X1 U9391 ( .A1(n8526), .A2(n8525), .ZN(n13977) );
  INV_X1 U9392 ( .A(n11697), .ZN(n6902) );
  NAND2_X1 U9393 ( .A1(n9884), .A2(n9883), .ZN(n14816) );
  NAND2_X1 U9394 ( .A1(n15235), .A2(n15234), .ZN(n15233) );
  INV_X1 U9395 ( .A(n11326), .ZN(n12791) );
  OR2_X1 U9396 ( .A1(n9867), .A2(n14763), .ZN(n6601) );
  OR2_X1 U9397 ( .A1(n10602), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6602) );
  OR2_X1 U9398 ( .A1(n9303), .A2(n9301), .ZN(n6603) );
  INV_X1 U9399 ( .A(n7596), .ZN(n13974) );
  OAI21_X1 U9400 ( .B1(n13373), .B2(n13372), .A(n13375), .ZN(n7596) );
  AND2_X1 U9401 ( .A1(n15333), .A2(n13051), .ZN(n6604) );
  NAND2_X1 U9402 ( .A1(n15150), .A2(n14914), .ZN(n6605) );
  NAND2_X1 U9403 ( .A1(n14349), .A2(n7416), .ZN(n7062) );
  NOR2_X1 U9404 ( .A1(n13538), .A2(n11890), .ZN(n6606) );
  OR2_X1 U9405 ( .A1(n13142), .A2(n7826), .ZN(n6607) );
  AND2_X1 U9406 ( .A1(n13493), .A2(n13810), .ZN(n6608) );
  NAND2_X1 U9407 ( .A1(n13279), .A2(n13836), .ZN(n6609) );
  INV_X1 U9408 ( .A(n7576), .ZN(n7581) );
  NAND2_X1 U9409 ( .A1(n8124), .A2(n8122), .ZN(n8261) );
  INV_X1 U9410 ( .A(n7644), .ZN(n7642) );
  AND2_X1 U9411 ( .A1(n15428), .A2(n13065), .ZN(n6610) );
  XOR2_X1 U9412 ( .A(n12985), .B(n14216), .Z(n6611) );
  AND2_X1 U9413 ( .A1(n8128), .A2(n8127), .ZN(n6612) );
  NAND3_X1 U9414 ( .A1(n7941), .A2(n6535), .A3(n7037), .ZN(n6613) );
  OR3_X1 U9415 ( .A1(n14570), .A2(n12777), .A3(n14215), .ZN(n6614) );
  OR2_X1 U9416 ( .A1(n9890), .A2(n9889), .ZN(n6615) );
  XNOR2_X1 U9417 ( .A(n10487), .B(P1_DATAO_REG_1__SCAN_IN), .ZN(n8143) );
  NAND2_X1 U9418 ( .A1(n13984), .A2(n13812), .ZN(n6616) );
  AND3_X1 U9419 ( .A1(n9511), .A2(n9510), .A3(n9512), .ZN(n6617) );
  NOR2_X1 U9420 ( .A1(n14908), .A2(n7907), .ZN(n6618) );
  AND2_X1 U9421 ( .A1(n12690), .A2(n13836), .ZN(n6619) );
  AND2_X1 U9422 ( .A1(n13262), .A2(n7021), .ZN(n6620) );
  INV_X1 U9423 ( .A(n9352), .ZN(n6995) );
  AND2_X1 U9424 ( .A1(n14658), .A2(n14233), .ZN(n9352) );
  OR2_X1 U9425 ( .A1(n14500), .A2(n14116), .ZN(n6621) );
  AND2_X1 U9426 ( .A1(n6601), .A2(n14846), .ZN(n6622) );
  AND2_X1 U9427 ( .A1(n13469), .A2(n7785), .ZN(n6623) );
  AND2_X1 U9428 ( .A1(n7914), .A2(n12925), .ZN(n6624) );
  NAND2_X1 U9429 ( .A1(n8976), .A2(n8975), .ZN(n14663) );
  INV_X1 U9430 ( .A(n14663), .ZN(n7859) );
  INV_X1 U9431 ( .A(n9883), .ZN(n7183) );
  INV_X1 U9432 ( .A(n9934), .ZN(n10789) );
  INV_X1 U9433 ( .A(n14354), .ZN(n14349) );
  NOR2_X1 U9434 ( .A1(n15066), .A2(n6870), .ZN(n6625) );
  XNOR2_X1 U9435 ( .A(n8794), .B(P2_IR_REG_29__SCAN_IN), .ZN(n8799) );
  INV_X1 U9436 ( .A(n8799), .ZN(n6985) );
  XOR2_X1 U9437 ( .A(n8845), .B(n8846), .Z(n6626) );
  OR2_X1 U9438 ( .A1(n6569), .A2(n13737), .ZN(n6627) );
  OR2_X1 U9439 ( .A1(n7327), .A2(n14277), .ZN(n6628) );
  NAND2_X1 U9440 ( .A1(n10054), .A2(n10530), .ZN(n11610) );
  INV_X1 U9441 ( .A(n14631), .ZN(n7919) );
  AND2_X1 U9442 ( .A1(n7634), .A2(n15613), .ZN(n6629) );
  XNOR2_X1 U9443 ( .A(n13032), .B(n14934), .ZN(n15387) );
  AND3_X1 U9444 ( .A1(n15147), .A2(n15146), .A3(n15145), .ZN(n6630) );
  AND2_X1 U9445 ( .A1(n11974), .A2(n11979), .ZN(n6631) );
  AND2_X1 U9446 ( .A1(n7690), .A2(n6605), .ZN(n6632) );
  AND2_X1 U9447 ( .A1(n8813), .A2(n8815), .ZN(n6633) );
  NAND2_X1 U9448 ( .A1(n6881), .A2(n6933), .ZN(n6634) );
  INV_X1 U9449 ( .A(n8718), .ZN(n7104) );
  OR2_X1 U9450 ( .A1(n15605), .A2(n15604), .ZN(n6635) );
  INV_X1 U9451 ( .A(n12889), .ZN(n8064) );
  AND2_X1 U9452 ( .A1(n7251), .A2(n7250), .ZN(n6636) );
  AND2_X1 U9453 ( .A1(n13202), .A2(n7839), .ZN(n6637) );
  OR2_X1 U9454 ( .A1(n13949), .A2(n13582), .ZN(n13407) );
  AND2_X1 U9455 ( .A1(n7459), .A2(n15156), .ZN(n6638) );
  NAND2_X1 U9456 ( .A1(n13221), .A2(n12691), .ZN(n6639) );
  INV_X1 U9457 ( .A(n13251), .ZN(n7273) );
  AND4_X1 U9458 ( .A1(n9048), .A2(n9047), .A3(n9046), .A4(n9045), .ZN(n14152)
         );
  INV_X1 U9459 ( .A(n14152), .ZN(n7107) );
  INV_X1 U9460 ( .A(n13805), .ZN(n13826) );
  INV_X1 U9461 ( .A(n15368), .ZN(n15491) );
  AND2_X1 U9462 ( .A1(n13091), .A2(n13090), .ZN(n6640) );
  AND2_X1 U9463 ( .A1(n11667), .A2(n11666), .ZN(n6641) );
  AND2_X1 U9464 ( .A1(n7472), .A2(n7471), .ZN(n6642) );
  NAND2_X1 U9465 ( .A1(n9247), .A2(n9246), .ZN(n13180) );
  AND2_X1 U9466 ( .A1(n6954), .A2(n6953), .ZN(n6643) );
  AND2_X1 U9467 ( .A1(n13506), .A2(n13505), .ZN(n13780) );
  INV_X1 U9468 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7051) );
  AND2_X1 U9469 ( .A1(n7025), .A2(n12328), .ZN(n6644) );
  AND2_X1 U9470 ( .A1(n15461), .A2(n14945), .ZN(n6645) );
  INV_X1 U9471 ( .A(n6855), .ZN(n13530) );
  NAND2_X1 U9472 ( .A1(n13515), .A2(n13522), .ZN(n6855) );
  AND2_X1 U9473 ( .A1(n9562), .A2(n6779), .ZN(n6646) );
  NOR2_X1 U9474 ( .A1(n12475), .A2(n14953), .ZN(n6647) );
  OR2_X1 U9475 ( .A1(n7108), .A2(n14152), .ZN(n6648) );
  AND3_X1 U9476 ( .A1(n8016), .A2(n13533), .A3(n8018), .ZN(n6649) );
  OR2_X1 U9477 ( .A1(n13874), .A2(n13848), .ZN(n13843) );
  NAND2_X1 U9478 ( .A1(n14522), .A2(n7917), .ZN(n7920) );
  OR2_X1 U9479 ( .A1(n9475), .A2(n14977), .ZN(n6650) );
  INV_X1 U9480 ( .A(n9371), .ZN(n7578) );
  AND2_X1 U9481 ( .A1(n7981), .A2(n7978), .ZN(n6651) );
  AND2_X1 U9482 ( .A1(n8827), .A2(n8826), .ZN(n14184) );
  INV_X1 U9483 ( .A(n14184), .ZN(n14227) );
  INV_X1 U9484 ( .A(n7502), .ZN(n7501) );
  NAND2_X1 U9485 ( .A1(n7503), .A2(n11214), .ZN(n7502) );
  OR2_X1 U9486 ( .A1(n8469), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n6652) );
  OR2_X1 U9487 ( .A1(n13229), .A2(n13768), .ZN(n6653) );
  INV_X1 U9488 ( .A(n12552), .ZN(n7767) );
  AND2_X1 U9489 ( .A1(n13487), .A2(n13488), .ZN(n13832) );
  INV_X1 U9490 ( .A(n13832), .ZN(n8004) );
  NAND2_X1 U9491 ( .A1(n14500), .A2(n14116), .ZN(n6654) );
  AND2_X1 U9492 ( .A1(n9360), .A2(n12884), .ZN(n6655) );
  INV_X1 U9493 ( .A(n7797), .ZN(n7796) );
  NAND2_X1 U9494 ( .A1(n13448), .A2(n13442), .ZN(n7797) );
  INV_X1 U9495 ( .A(n7992), .ZN(n15231) );
  NOR2_X1 U9496 ( .A1(n15285), .A2(n7994), .ZN(n7992) );
  AND2_X1 U9497 ( .A1(n14590), .A2(n14222), .ZN(n6656) );
  OR2_X1 U9498 ( .A1(n12602), .A2(n12603), .ZN(n6657) );
  AND4_X1 U9499 ( .A1(n9383), .A2(n9382), .A3(n9381), .A4(n9643), .ZN(n6658)
         );
  OR2_X1 U9500 ( .A1(n15139), .A2(n15141), .ZN(n6659) );
  NAND2_X1 U9501 ( .A1(n7701), .A2(n6833), .ZN(n15280) );
  AND2_X1 U9502 ( .A1(n15466), .A2(n14946), .ZN(n6660) );
  AND2_X1 U9503 ( .A1(n13853), .A2(n13864), .ZN(n6661) );
  AND2_X1 U9504 ( .A1(n6609), .A2(n7673), .ZN(n6662) );
  AND2_X1 U9505 ( .A1(n15447), .A2(n14943), .ZN(n6663) );
  AND2_X1 U9506 ( .A1(n12593), .A2(n12592), .ZN(n15383) );
  INV_X1 U9507 ( .A(n15383), .ZN(n15121) );
  NAND2_X1 U9508 ( .A1(n9576), .A2(n9575), .ZN(n12416) );
  INV_X1 U9509 ( .A(n12416), .ZN(n12417) );
  NAND2_X1 U9510 ( .A1(n7559), .A2(n7560), .ZN(n6664) );
  AND2_X1 U9511 ( .A1(n7018), .A2(n7019), .ZN(n6665) );
  INV_X1 U9512 ( .A(n13453), .ZN(n6889) );
  INV_X1 U9513 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8817) );
  AND2_X1 U9514 ( .A1(n8867), .A2(n7844), .ZN(n15880) );
  AND2_X1 U9515 ( .A1(n14822), .A2(n14938), .ZN(n6666) );
  OR2_X1 U9516 ( .A1(n9362), .A2(n9361), .ZN(n6667) );
  OR2_X1 U9517 ( .A1(n8753), .A2(SI_18_), .ZN(n6668) );
  NAND2_X1 U9518 ( .A1(n12578), .A2(n12577), .ZN(n13032) );
  INV_X1 U9519 ( .A(n7684), .ZN(n7680) );
  OR2_X1 U9520 ( .A1(n13977), .A2(n13576), .ZN(n7684) );
  INV_X1 U9521 ( .A(n7847), .ZN(n7121) );
  NAND2_X1 U9522 ( .A1(n6556), .A2(n6654), .ZN(n7847) );
  AND2_X1 U9523 ( .A1(n13482), .A2(n13481), .ZN(n6669) );
  INV_X1 U9524 ( .A(n7813), .ZN(n7812) );
  NAND2_X1 U9525 ( .A1(n13478), .A2(n13474), .ZN(n7813) );
  AND2_X1 U9526 ( .A1(n7128), .A2(n14227), .ZN(n6670) );
  AND2_X1 U9527 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_REG3_REG_6__SCAN_IN), 
        .ZN(n6671) );
  OR2_X1 U9528 ( .A1(n14307), .A2(n14219), .ZN(n6672) );
  INV_X1 U9529 ( .A(n13951), .ZN(n13958) );
  INV_X1 U9530 ( .A(n13958), .ZN(n6916) );
  AND2_X1 U9531 ( .A1(n8709), .A2(SI_6_), .ZN(n6673) );
  INV_X1 U9532 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9610) );
  INV_X1 U9533 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9591) );
  INV_X1 U9534 ( .A(n8764), .ZN(n7059) );
  INV_X1 U9535 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10802) );
  INV_X1 U9536 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9394) );
  INV_X1 U9537 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9420) );
  NOR2_X1 U9538 ( .A1(n13912), .A2(n13803), .ZN(n6674) );
  NOR2_X1 U9539 ( .A1(n14643), .A2(n14232), .ZN(n6675) );
  NOR2_X1 U9540 ( .A1(n14600), .A2(n14059), .ZN(n6676) );
  AND2_X1 U9541 ( .A1(n7110), .A2(n7109), .ZN(n6677) );
  NAND2_X1 U9542 ( .A1(n7233), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n10551) );
  NAND2_X1 U9543 ( .A1(n9207), .A2(n9206), .ZN(n14590) );
  OR2_X1 U9544 ( .A1(n9475), .A2(n10582), .ZN(n6678) );
  INV_X1 U9545 ( .A(n7024), .ZN(n7023) );
  NAND2_X1 U9546 ( .A1(n13224), .A2(n13775), .ZN(n7024) );
  NAND2_X1 U9547 ( .A1(n7835), .A2(n8833), .ZN(n6679) );
  INV_X1 U9548 ( .A(n7461), .ZN(n7460) );
  NAND2_X1 U9549 ( .A1(n13023), .A2(n13022), .ZN(n7461) );
  INV_X1 U9550 ( .A(n7923), .ZN(n7922) );
  NAND2_X1 U9551 ( .A1(n6572), .A2(n7859), .ZN(n7923) );
  INV_X1 U9552 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7302) );
  AND2_X1 U9553 ( .A1(n12815), .A2(n14092), .ZN(n6680) );
  AND2_X1 U9554 ( .A1(n7661), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n6681) );
  AND2_X1 U9555 ( .A1(n7957), .A2(n7956), .ZN(n6682) );
  AND2_X1 U9556 ( .A1(n9815), .A2(n9817), .ZN(n6683) );
  NAND2_X1 U9557 ( .A1(n14576), .A2(n14219), .ZN(n6684) );
  AND2_X1 U9558 ( .A1(n7317), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n6685) );
  AND2_X1 U9559 ( .A1(n8289), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n6686) );
  NAND2_X1 U9560 ( .A1(n7719), .A2(n7725), .ZN(n7718) );
  INV_X1 U9561 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n8722) );
  OAI21_X1 U9562 ( .B1(n10074), .B2(n7077), .A(P3_REG1_REG_7__SCAN_IN), .ZN(
        n7076) );
  AND2_X1 U9563 ( .A1(n9706), .A2(n9707), .ZN(n6687) );
  AND2_X1 U9564 ( .A1(n9684), .A2(n9683), .ZN(n6688) );
  AND2_X1 U9565 ( .A1(n7692), .A2(n7455), .ZN(n6689) );
  NAND2_X1 U9566 ( .A1(n14590), .A2(n7417), .ZN(n6690) );
  AND2_X1 U9567 ( .A1(n7909), .A2(n7910), .ZN(n14370) );
  NAND2_X1 U9568 ( .A1(n7883), .A2(n7881), .ZN(n14760) );
  AND2_X1 U9569 ( .A1(n14615), .A2(n14184), .ZN(n6691) );
  NAND2_X1 U9570 ( .A1(n8758), .A2(n9153), .ZN(n6692) );
  NAND2_X1 U9571 ( .A1(n8431), .A2(n8430), .ZN(n6693) );
  INV_X1 U9572 ( .A(n7398), .ZN(n7397) );
  OAI21_X1 U9573 ( .B1(n7399), .B2(n7401), .A(n8650), .ZN(n7398) );
  INV_X1 U9574 ( .A(n9832), .ZN(n7886) );
  OR2_X1 U9575 ( .A1(n13438), .A2(n13431), .ZN(n6694) );
  AND3_X1 U9576 ( .A1(n13172), .A2(n13177), .A3(n14161), .ZN(n6695) );
  AND2_X1 U9577 ( .A1(n6622), .A2(n14817), .ZN(n6696) );
  AND2_X1 U9578 ( .A1(n6905), .A2(n8660), .ZN(n6697) );
  AND2_X1 U9579 ( .A1(n8849), .A2(n7008), .ZN(n6698) );
  AND2_X1 U9580 ( .A1(n7784), .A2(n8366), .ZN(n6699) );
  INV_X1 U9581 ( .A(n12804), .ZN(n8076) );
  AND2_X1 U9582 ( .A1(n7644), .A2(n15613), .ZN(n6700) );
  NAND2_X1 U9583 ( .A1(n8755), .A2(n8754), .ZN(n6701) );
  INV_X1 U9584 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7661) );
  MUX2_X1 U9585 ( .A(n14241), .B(n12791), .S(n6542), .Z(n12792) );
  NAND2_X1 U9586 ( .A1(n8656), .A2(n7814), .ZN(n6702) );
  AND2_X1 U9587 ( .A1(n12984), .A2(n14556), .ZN(n6703) );
  INV_X1 U9588 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8132) );
  NAND2_X1 U9589 ( .A1(n9938), .A2(n6618), .ZN(n6704) );
  AND2_X1 U9590 ( .A1(n13788), .A2(n6616), .ZN(n7409) );
  OR2_X1 U9591 ( .A1(n14582), .A2(n15879), .ZN(n6705) );
  NOR2_X1 U9592 ( .A1(n14150), .A2(n7824), .ZN(n7823) );
  AND3_X1 U9593 ( .A1(n7730), .A2(n7741), .A3(n12629), .ZN(n6706) );
  INV_X1 U9594 ( .A(n12574), .ZN(n7294) );
  NAND2_X1 U9595 ( .A1(n9922), .A2(n9921), .ZN(n15150) );
  OR2_X1 U9596 ( .A1(n15472), .A2(n13052), .ZN(n6707) );
  AND2_X1 U9597 ( .A1(n7418), .A2(n6609), .ZN(n6708) );
  OR2_X1 U9598 ( .A1(n14643), .A2(n14203), .ZN(n6709) );
  AND2_X1 U9599 ( .A1(n13557), .A2(n13520), .ZN(n6710) );
  AND3_X1 U9600 ( .A1(n6535), .A2(n8106), .A3(n7313), .ZN(n6711) );
  AND2_X1 U9601 ( .A1(n15565), .A2(n15564), .ZN(n6712) );
  INV_X1 U9602 ( .A(n15625), .ZN(n7247) );
  AND2_X1 U9603 ( .A1(n13483), .A2(n13480), .ZN(n6713) );
  NOR2_X1 U9604 ( .A1(n15028), .A2(n15029), .ZN(n6714) );
  NOR2_X1 U9605 ( .A1(n7736), .A2(n7740), .ZN(n7735) );
  INV_X1 U9606 ( .A(n7735), .ZN(n7731) );
  NAND2_X1 U9607 ( .A1(n13387), .A2(n13386), .ZN(n13559) );
  INV_X1 U9608 ( .A(n13559), .ZN(n7230) );
  NOR2_X1 U9609 ( .A1(n14454), .A2(n6959), .ZN(n6715) );
  AND2_X1 U9610 ( .A1(n9372), .A2(n9256), .ZN(n12983) );
  INV_X1 U9611 ( .A(n12983), .ZN(n6966) );
  AND2_X1 U9612 ( .A1(n10952), .A2(n7651), .ZN(n6716) );
  INV_X1 U9613 ( .A(n13064), .ZN(n7710) );
  AND2_X1 U9614 ( .A1(n14463), .A2(n9359), .ZN(n6717) );
  NAND2_X1 U9615 ( .A1(n15163), .A2(n14937), .ZN(n6718) );
  AND2_X1 U9616 ( .A1(n8782), .A2(n8793), .ZN(n6719) );
  AND2_X1 U9617 ( .A1(n8660), .A2(n8662), .ZN(n6720) );
  AND2_X1 U9618 ( .A1(n8215), .A2(n7773), .ZN(n6721) );
  OR2_X1 U9619 ( .A1(n9475), .A2(n10488), .ZN(n6722) );
  AND2_X1 U9620 ( .A1(n7280), .A2(n12676), .ZN(n6723) );
  AND2_X1 U9621 ( .A1(n9621), .A2(n9603), .ZN(n6724) );
  AND2_X1 U9622 ( .A1(n7247), .A2(n7246), .ZN(n6725) );
  OR2_X1 U9623 ( .A1(n7767), .A2(n12551), .ZN(n6726) );
  AND2_X1 U9624 ( .A1(n8021), .A2(n8020), .ZN(n6727) );
  OR2_X1 U9625 ( .A1(n7764), .A2(n12559), .ZN(n6728) );
  AND2_X1 U9626 ( .A1(n6624), .A2(n7913), .ZN(n6729) );
  AND2_X1 U9627 ( .A1(n13311), .A2(n12688), .ZN(n6730) );
  INV_X1 U9628 ( .A(n12908), .ZN(n7157) );
  AND2_X1 U9629 ( .A1(n13708), .A2(n13707), .ZN(n6731) );
  INV_X1 U9630 ( .A(n12956), .ZN(n7865) );
  OR2_X1 U9631 ( .A1(n6955), .A2(n6669), .ZN(n6732) );
  AND2_X1 U9632 ( .A1(n8132), .A2(n6919), .ZN(n6733) );
  NAND2_X1 U9633 ( .A1(n12951), .A2(n12950), .ZN(n6734) );
  AND2_X1 U9634 ( .A1(n15587), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n6735) );
  AND2_X1 U9635 ( .A1(n15163), .A2(n13069), .ZN(n6736) );
  AND2_X1 U9636 ( .A1(n6719), .A2(n8795), .ZN(n6737) );
  AND2_X1 U9637 ( .A1(n7422), .A2(n13176), .ZN(n6738) );
  AND2_X1 U9638 ( .A1(n6703), .A2(n6585), .ZN(n6739) );
  NAND2_X1 U9639 ( .A1(n8031), .A2(n13517), .ZN(n6740) );
  NAND2_X1 U9640 ( .A1(n12799), .A2(n12800), .ZN(n8917) );
  INV_X1 U9641 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9405) );
  AND2_X1 U9642 ( .A1(n7840), .A2(n8817), .ZN(n6741) );
  AND2_X1 U9643 ( .A1(n6588), .A2(n7254), .ZN(n6742) );
  AND2_X1 U9644 ( .A1(n6627), .A2(n13667), .ZN(n6743) );
  INV_X1 U9645 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n6931) );
  INV_X1 U9646 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9396) );
  INV_X1 U9647 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7345) );
  INV_X1 U9648 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8782) );
  INV_X1 U9649 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7317) );
  INV_X1 U9650 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10757) );
  OR2_X1 U9651 ( .A1(n13547), .A2(n7310), .ZN(n6744) );
  XOR2_X1 U9652 ( .A(n13211), .B(n13776), .Z(n6745) );
  INV_X1 U9653 ( .A(n14476), .ZN(n6960) );
  XNOR2_X1 U9654 ( .A(n8622), .B(n8621), .ZN(n13412) );
  NAND2_X1 U9655 ( .A1(n7625), .A2(n11317), .ZN(n10149) );
  NAND2_X1 U9656 ( .A1(n7169), .A2(n7167), .ZN(n11999) );
  INV_X1 U9657 ( .A(n15245), .ZN(n7955) );
  AND2_X1 U9658 ( .A1(n10083), .A2(n10085), .ZN(n6746) );
  NAND2_X1 U9659 ( .A1(n11740), .A2(n9350), .ZN(n11362) );
  NAND2_X1 U9660 ( .A1(n10075), .A2(n10166), .ZN(n10170) );
  NAND2_X1 U9661 ( .A1(n11845), .A2(n7925), .ZN(n12037) );
  OAI21_X1 U9662 ( .B1(n11363), .B2(n7853), .A(n7851), .ZN(n12158) );
  XNOR2_X1 U9663 ( .A(n8583), .B(P3_IR_REG_24__SCAN_IN), .ZN(n8592) );
  INV_X1 U9664 ( .A(n8592), .ZN(n7283) );
  NAND2_X1 U9665 ( .A1(n7857), .A2(n7855), .ZN(n12060) );
  INV_X1 U9666 ( .A(n13538), .ZN(n11757) );
  NAND2_X1 U9667 ( .A1(n6886), .A2(n6591), .ZN(n12383) );
  NAND2_X1 U9668 ( .A1(n12353), .A2(n12231), .ZN(n12326) );
  NAND2_X1 U9669 ( .A1(n7696), .A2(n11576), .ZN(n15670) );
  XOR2_X1 U9670 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .Z(n6747) );
  INV_X1 U9671 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7943) );
  AND2_X1 U9672 ( .A1(n10505), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n6748) );
  OR2_X1 U9673 ( .A1(n11317), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n6749) );
  AND2_X1 U9674 ( .A1(n11095), .A2(n7921), .ZN(n12068) );
  AND2_X1 U9675 ( .A1(n13957), .A2(n8633), .ZN(n6750) );
  INV_X1 U9676 ( .A(n7988), .ZN(n12211) );
  NAND2_X1 U9677 ( .A1(n7403), .A2(n8647), .ZN(n7399) );
  INV_X1 U9678 ( .A(n7399), .ZN(n6907) );
  AND2_X1 U9679 ( .A1(n8199), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n6751) );
  NOR2_X1 U9680 ( .A1(n11479), .A2(n11476), .ZN(n6752) );
  NAND2_X1 U9681 ( .A1(n6929), .A2(n6930), .ZN(n6753) );
  INV_X1 U9682 ( .A(n7488), .ZN(n7487) );
  NOR2_X1 U9683 ( .A1(n12610), .A2(n7489), .ZN(n7488) );
  OR2_X1 U9684 ( .A1(n15976), .A2(n13900), .ZN(n6754) );
  NOR2_X1 U9685 ( .A1(n11966), .A2(n11965), .ZN(n6755) );
  INV_X1 U9686 ( .A(n6791), .ZN(n14557) );
  AND2_X1 U9687 ( .A1(n13843), .A2(n13480), .ZN(n13869) );
  AND2_X1 U9688 ( .A1(n7543), .A2(n7542), .ZN(n6756) );
  OR2_X1 U9689 ( .A1(n9240), .A2(n12311), .ZN(n6757) );
  AND2_X1 U9690 ( .A1(n13462), .A2(n8649), .ZN(n13549) );
  INV_X1 U9691 ( .A(n13549), .ZN(n7403) );
  INV_X1 U9692 ( .A(n7513), .ZN(n7512) );
  NOR2_X1 U9693 ( .A1(n9208), .A2(SI_25_), .ZN(n7513) );
  AND2_X1 U9694 ( .A1(n13903), .A2(n6754), .ZN(n6758) );
  AND2_X1 U9695 ( .A1(n13978), .A2(n7426), .ZN(n6759) );
  NAND2_X1 U9696 ( .A1(n8814), .A2(n8813), .ZN(n6760) );
  NAND2_X1 U9697 ( .A1(n7941), .A2(n6535), .ZN(n6761) );
  AND2_X1 U9698 ( .A1(n10709), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n6762) );
  AND2_X1 U9699 ( .A1(n9235), .A2(SI_26_), .ZN(n6763) );
  AND2_X1 U9700 ( .A1(n12609), .A2(SI_30_), .ZN(n6764) );
  INV_X1 U9701 ( .A(n7508), .ZN(n7507) );
  NAND2_X1 U9702 ( .A1(n7510), .A2(n6757), .ZN(n7508) );
  NOR2_X1 U9703 ( .A1(n9181), .A2(SI_23_), .ZN(n6765) );
  AND2_X1 U9704 ( .A1(n8679), .A2(n8678), .ZN(n6766) );
  NOR2_X1 U9705 ( .A1(n9241), .A2(SI_27_), .ZN(n6767) );
  OR2_X1 U9706 ( .A1(n7487), .A2(n7484), .ZN(n6768) );
  AND2_X1 U9707 ( .A1(n7745), .A2(n7746), .ZN(n6769) );
  OR2_X1 U9708 ( .A1(n14307), .A2(n14171), .ZN(n6770) );
  AND2_X1 U9709 ( .A1(n15830), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6771) );
  NOR2_X1 U9710 ( .A1(n6825), .A2(n13721), .ZN(n6772) );
  NAND2_X1 U9711 ( .A1(n13402), .A2(n13478), .ZN(n13877) );
  AND2_X1 U9712 ( .A1(n7774), .A2(n13428), .ZN(n6773) );
  NAND2_X1 U9713 ( .A1(n10505), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6774) );
  AND2_X1 U9714 ( .A1(n7545), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n6775) );
  INV_X1 U9715 ( .A(n7129), .ZN(n7127) );
  NAND2_X1 U9716 ( .A1(n9360), .A2(n14228), .ZN(n7129) );
  NAND2_X1 U9717 ( .A1(n7094), .A2(n10530), .ZN(n11615) );
  INV_X1 U9718 ( .A(n12964), .ZN(n6958) );
  AND2_X2 U9719 ( .A1(n11092), .A2(n9376), .ZN(n15893) );
  AND2_X2 U9720 ( .A1(n11092), .A2(n9335), .ZN(n15886) );
  AND2_X2 U9721 ( .A1(n15520), .A2(n15519), .ZN(n15791) );
  AND2_X1 U9722 ( .A1(n15835), .A2(n6594), .ZN(n6776) );
  NAND2_X1 U9723 ( .A1(n6835), .A2(n6838), .ZN(n9723) );
  INV_X2 U9724 ( .A(n15973), .ZN(n15976) );
  AND2_X1 U9725 ( .A1(n10640), .A2(n10639), .ZN(n15811) );
  INV_X1 U9726 ( .A(n15479), .ZN(n7967) );
  NAND2_X1 U9727 ( .A1(n14243), .A2(n11158), .ZN(n11150) );
  INV_X1 U9728 ( .A(n11150), .ZN(n7292) );
  NAND2_X1 U9729 ( .A1(n8960), .A2(n8959), .ZN(n14668) );
  INV_X1 U9730 ( .A(n14668), .ZN(n7924) );
  INV_X1 U9731 ( .A(n14626), .ZN(n7918) );
  INV_X1 U9732 ( .A(n15486), .ZN(n7990) );
  NAND2_X1 U9733 ( .A1(n7075), .A2(n11145), .ZN(n10167) );
  NAND2_X1 U9734 ( .A1(n11256), .A2(n13567), .ZN(n13360) );
  NAND2_X1 U9735 ( .A1(n7878), .A2(n9507), .ZN(n15633) );
  INV_X1 U9736 ( .A(n7686), .ZN(n10189) );
  NAND2_X1 U9737 ( .A1(n10188), .A2(n9475), .ZN(n7686) );
  AND2_X1 U9738 ( .A1(n7071), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n6777) );
  OR2_X1 U9739 ( .A1(n9237), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6778) );
  INV_X1 U9740 ( .A(n10131), .ZN(n7624) );
  OAI21_X1 U9741 ( .B1(n15114), .B2(n15668), .A(n15113), .ZN(n7532) );
  NAND2_X1 U9742 ( .A1(n9581), .A2(n9582), .ZN(n6779) );
  AND2_X1 U9743 ( .A1(n12341), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6780) );
  INV_X1 U9744 ( .A(n13707), .ZN(n7556) );
  AND2_X1 U9745 ( .A1(n9237), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6781) );
  AND2_X1 U9746 ( .A1(n12219), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6782) );
  INV_X1 U9747 ( .A(n12430), .ZN(n12428) );
  INV_X1 U9748 ( .A(n7378), .ZN(n6814) );
  OR2_X1 U9749 ( .A1(n13693), .A2(n13692), .ZN(n7378) );
  AND2_X1 U9750 ( .A1(n11043), .A2(n7831), .ZN(n6783) );
  INV_X1 U9751 ( .A(n7616), .ZN(n7615) );
  NAND2_X1 U9752 ( .A1(n7619), .A2(n6778), .ZN(n7616) );
  OR2_X1 U9753 ( .A1(n13693), .A2(n13671), .ZN(n6784) );
  INV_X1 U9754 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7358) );
  XOR2_X1 U9755 ( .A(n7066), .B(n10523), .Z(n6785) );
  NAND2_X1 U9756 ( .A1(n11213), .A2(n13745), .ZN(n13529) );
  XOR2_X1 U9757 ( .A(n10505), .B(n12116), .Z(n6786) );
  INV_X1 U9758 ( .A(n12987), .ZN(n14299) );
  INV_X1 U9759 ( .A(n10903), .ZN(n7055) );
  AND2_X1 U9760 ( .A1(n7570), .A2(n11684), .ZN(n6787) );
  AND2_X1 U9761 ( .A1(n10596), .A2(n6602), .ZN(n6788) );
  AND2_X1 U9762 ( .A1(n9333), .A2(n9334), .ZN(n15844) );
  INV_X1 U9763 ( .A(n12955), .ZN(n8051) );
  NAND2_X1 U9764 ( .A1(n11134), .A2(n11110), .ZN(n9291) );
  AND2_X1 U9765 ( .A1(n7520), .A2(n7521), .ZN(n6789) );
  AND2_X1 U9766 ( .A1(n9276), .A2(n9314), .ZN(n12988) );
  INV_X1 U9767 ( .A(n12988), .ZN(n11110) );
  AND2_X1 U9768 ( .A1(n10934), .A2(n7232), .ZN(n6790) );
  INV_X1 U9769 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7585) );
  INV_X1 U9770 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7438) );
  INV_X1 U9771 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7356) );
  INV_X1 U9772 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n7246) );
  OR2_X1 U9773 ( .A1(n9169), .A2(n10594), .ZN(n8904) );
  NAND2_X1 U9774 ( .A1(n7912), .A2(n7911), .ZN(n14371) );
  NOR2_X2 U9775 ( .A1(n14428), .A2(n14610), .ZN(n7912) );
  NAND2_X1 U9776 ( .A1(n7138), .A2(n7135), .ZN(n12813) );
  OAI21_X1 U9777 ( .B1(n12900), .B2(n8038), .A(n8037), .ZN(n12904) );
  INV_X1 U9778 ( .A(n8065), .ZN(n8062) );
  NAND3_X1 U9779 ( .A1(n6793), .A2(n13153), .A3(n8095), .ZN(n14132) );
  NAND2_X1 U9780 ( .A1(n13201), .A2(n6695), .ZN(n13182) );
  NAND2_X1 U9781 ( .A1(n8735), .A2(SI_15_), .ZN(n6795) );
  NAND3_X1 U9782 ( .A1(n6642), .A2(n7065), .A3(n8751), .ZN(n6796) );
  OAI21_X1 U9783 ( .B1(n9260), .B2(P2_DATAO_REG_15__SCAN_IN), .A(n7341), .ZN(
        n8734) );
  OR2_X2 U9784 ( .A1(n9119), .A2(n9118), .ZN(n9121) );
  NAND2_X1 U9785 ( .A1(n6798), .A2(n6797), .ZN(P3_U3199) );
  AOI21_X1 U9786 ( .B1(n11635), .B2(n11610), .A(n11611), .ZN(n11613) );
  NAND2_X1 U9787 ( .A1(n11376), .A2(n10051), .ZN(n10052) );
  INV_X1 U9788 ( .A(n6928), .ZN(n10057) );
  NAND2_X1 U9789 ( .A1(n7544), .A2(n11964), .ZN(n6930) );
  NAND2_X1 U9790 ( .A1(n11143), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n10172) );
  NAND2_X1 U9791 ( .A1(n10060), .A2(n7091), .ZN(n7566) );
  OAI22_X1 U9792 ( .A1(n8151), .A2(n7086), .B1(P3_IR_REG_31__SCAN_IN), .B2(
        P3_IR_REG_2__SCAN_IN), .ZN(n7085) );
  AOI21_X1 U9793 ( .B1(n13608), .B2(n6930), .A(n13607), .ZN(n13610) );
  NAND2_X1 U9794 ( .A1(n6547), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n13709) );
  INV_X1 U9795 ( .A(n12894), .ZN(n7161) );
  NAND2_X1 U9796 ( .A1(n7137), .A2(n7136), .ZN(n7135) );
  NAND2_X1 U9797 ( .A1(n7140), .A2(n7139), .ZN(n7138) );
  NAND2_X1 U9798 ( .A1(n7340), .A2(n7338), .ZN(n12897) );
  NAND2_X1 U9799 ( .A1(n7158), .A2(n12906), .ZN(n7153) );
  NAND2_X1 U9800 ( .A1(n7156), .A2(n7155), .ZN(n12912) );
  OR2_X1 U9801 ( .A1(n12794), .A2(n12792), .ZN(n8055) );
  NAND2_X1 U9802 ( .A1(n7098), .A2(n8711), .ZN(n8954) );
  INV_X1 U9803 ( .A(n7718), .ZN(n7717) );
  NAND2_X1 U9804 ( .A1(n7105), .A2(n9002), .ZN(n9005) );
  NAND2_X1 U9805 ( .A1(n7278), .A2(n7383), .ZN(n9033) );
  OAI21_X1 U9806 ( .B1(n12490), .B2(n7718), .A(n7714), .ZN(n7723) );
  NAND2_X1 U9807 ( .A1(n12576), .A2(n7294), .ZN(n7293) );
  NAND3_X1 U9808 ( .A1(n6802), .A2(n6801), .A3(n6726), .ZN(n7765) );
  NAND2_X1 U9809 ( .A1(n12550), .A2(n12549), .ZN(n6801) );
  NAND2_X1 U9810 ( .A1(n12546), .A2(n12545), .ZN(n6802) );
  AOI22_X1 U9811 ( .A1(n14290), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n14288), 
        .B2(n14289), .ZN(n14291) );
  XNOR2_X1 U9812 ( .A(n14287), .B(n14289), .ZN(n14290) );
  OAI22_X1 U9813 ( .A1(n12570), .A2(n7763), .B1(n12571), .B2(n7762), .ZN(
        n12576) );
  OAI21_X1 U9814 ( .B1(n14297), .B2(n7336), .A(n7335), .ZN(n14301) );
  NAND2_X1 U9815 ( .A1(n7297), .A2(n7296), .ZN(n12563) );
  NAND3_X1 U9816 ( .A1(n12473), .A2(n12472), .A3(n6803), .ZN(n12477) );
  NAND2_X1 U9817 ( .A1(n6804), .A2(n7700), .ZN(n6803) );
  INV_X1 U9818 ( .A(n12474), .ZN(n6804) );
  NOR2_X1 U9819 ( .A1(n15824), .A2(n6771), .ZN(n10897) );
  NAND2_X1 U9820 ( .A1(n14296), .A2(n15815), .ZN(n7049) );
  NAND4_X1 U9821 ( .A1(n7778), .A2(n8114), .A3(n6535), .A4(n8113), .ZN(n8582)
         );
  NAND2_X1 U9822 ( .A1(n13716), .A2(n13725), .ZN(n13738) );
  NAND2_X1 U9823 ( .A1(n6816), .A2(n10114), .ZN(n11137) );
  NAND3_X1 U9824 ( .A1(n6818), .A2(n11135), .A3(n6817), .ZN(n6816) );
  NAND3_X1 U9825 ( .A1(n6821), .A2(n10107), .A3(n6820), .ZN(n6818) );
  INV_X1 U9826 ( .A(n11643), .ZN(n6822) );
  OAI21_X1 U9827 ( .B1(n10152), .B2(n6824), .A(n6823), .ZN(n13620) );
  XNOR2_X1 U9828 ( .A(n6832), .B(n8972), .ZN(n10510) );
  NAND2_X2 U9829 ( .A1(n7056), .A2(n8715), .ZN(n6832) );
  NAND2_X1 U9830 ( .A1(n9063), .A2(n6837), .ZN(n6836) );
  NAND3_X1 U9831 ( .A1(n6836), .A2(n9075), .A3(n9074), .ZN(n6835) );
  NAND2_X1 U9832 ( .A1(n7342), .A2(n9079), .ZN(n6841) );
  NOR3_X2 U9833 ( .A1(n8469), .A2(P3_REG3_REG_22__SCAN_IN), .A3(
        P3_REG3_REG_23__SCAN_IN), .ZN(n7361) );
  NAND2_X1 U9834 ( .A1(n6854), .A2(n6653), .ZN(n7362) );
  NAND2_X1 U9835 ( .A1(n7678), .A2(n6855), .ZN(n6854) );
  NAND2_X1 U9836 ( .A1(n7533), .A2(n6856), .ZN(P1_U3262) );
  AOI21_X1 U9837 ( .B1(n6857), .B2(n15112), .A(n7532), .ZN(n6856) );
  NAND2_X1 U9838 ( .A1(n6858), .A2(n7535), .ZN(n6857) );
  NAND2_X1 U9839 ( .A1(n15109), .A2(n15108), .ZN(n6858) );
  NAND3_X1 U9840 ( .A1(n10596), .A2(n6863), .A3(n6602), .ZN(n15002) );
  NAND4_X1 U9841 ( .A1(n10596), .A2(n6862), .A3(n6863), .A4(n6602), .ZN(n6861)
         );
  OAI21_X2 U9842 ( .B1(n15297), .B2(n6866), .A(n6864), .ZN(n15263) );
  NOR2_X2 U9843 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n6881) );
  INV_X1 U9844 ( .A(n6883), .ZN(n7675) );
  NAND3_X1 U9845 ( .A1(n6721), .A2(n7775), .A3(n7774), .ZN(n6892) );
  NAND2_X1 U9846 ( .A1(n6895), .A2(n7775), .ZN(n6893) );
  INV_X1 U9847 ( .A(n8646), .ZN(n6908) );
  OAI21_X1 U9848 ( .B1(n8646), .B2(n7399), .A(n7397), .ZN(n13882) );
  OAI21_X1 U9849 ( .B1(n13959), .B2(n6911), .A(n6910), .ZN(n11502) );
  INV_X1 U9850 ( .A(n6913), .ZN(n6912) );
  OAI21_X1 U9851 ( .B1(n8633), .B2(n6561), .A(n11501), .ZN(n6913) );
  NAND3_X1 U9852 ( .A1(n6917), .A2(n11778), .A3(n7277), .ZN(n13415) );
  NAND2_X1 U9853 ( .A1(n7404), .A2(n7406), .ZN(n7683) );
  NAND2_X1 U9854 ( .A1(n6923), .A2(n6922), .ZN(P3_U3200) );
  OAI21_X1 U9855 ( .B1(n13734), .B2(n6924), .A(n13667), .ZN(n6923) );
  AND2_X1 U9856 ( .A1(n13709), .A2(n6731), .ZN(n6924) );
  NOR2_X2 U9857 ( .A1(n10056), .A2(n6925), .ZN(n11143) );
  OR2_X2 U9858 ( .A1(n11613), .A2(n10055), .ZN(n6926) );
  OR2_X2 U9859 ( .A1(n10171), .A2(n6927), .ZN(n6928) );
  NAND2_X1 U9860 ( .A1(n10059), .A2(n7353), .ZN(n6929) );
  NAND3_X1 U9861 ( .A1(n6929), .A2(P3_REG2_REG_11__SCAN_IN), .A3(n6930), .ZN(
        n13608) );
  MUX2_X1 U9862 ( .A(n14042), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  MUX2_X1 U9863 ( .A(P3_IR_REG_0__SCAN_IN), .B(n14042), .S(n10063), .Z(n11277)
         );
  NOR2_X2 U9864 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n6933) );
  NAND2_X1 U9865 ( .A1(n6937), .A2(n6935), .ZN(n6934) );
  AOI21_X1 U9866 ( .B1(n6936), .B2(n6590), .A(n6740), .ZN(n6935) );
  OAI21_X1 U9867 ( .B1(n13518), .B2(n8032), .A(n13526), .ZN(n6936) );
  NAND2_X1 U9868 ( .A1(n6938), .A2(n6710), .ZN(n6937) );
  NAND2_X1 U9869 ( .A1(n13516), .A2(n13515), .ZN(n6938) );
  NAND4_X1 U9870 ( .A1(n13451), .A2(n13450), .A3(n13449), .A4(n13453), .ZN(
        n6952) );
  NAND2_X1 U9871 ( .A1(n6555), .A2(n6732), .ZN(n6953) );
  NAND3_X1 U9872 ( .A1(n13471), .A2(n6587), .A3(n6555), .ZN(n6954) );
  NAND3_X1 U9873 ( .A1(n8913), .A2(n6958), .A3(n10977), .ZN(n6956) );
  XNOR2_X1 U9874 ( .A(n11326), .B(n6957), .ZN(n10977) );
  INV_X1 U9875 ( .A(n14241), .ZN(n6957) );
  NAND4_X1 U9876 ( .A1(n12976), .A2(n12974), .A3(n6961), .A4(n6557), .ZN(n6959) );
  NAND4_X1 U9877 ( .A1(n6966), .A2(n12986), .A3(n14309), .A4(n6965), .ZN(n6964) );
  NAND2_X2 U9878 ( .A1(n14098), .A2(n7838), .ZN(n7837) );
  OAI21_X1 U9879 ( .B1(n12143), .B2(n6972), .A(n6970), .ZN(n14173) );
  NAND2_X1 U9880 ( .A1(n6969), .A2(n6967), .ZN(n13096) );
  NAND2_X1 U9881 ( .A1(n12143), .A2(n6970), .ZN(n6969) );
  OAI21_X1 U9882 ( .B1(n11229), .B2(n6975), .A(n6973), .ZN(n11901) );
  AOI21_X1 U9883 ( .B1(n6974), .B2(n6976), .A(n6641), .ZN(n6973) );
  INV_X1 U9884 ( .A(n11230), .ZN(n6974) );
  NAND2_X1 U9885 ( .A1(n14089), .A2(n7823), .ZN(n6978) );
  NAND2_X1 U9886 ( .A1(n6978), .A2(n6979), .ZN(n14046) );
  INV_X1 U9887 ( .A(n14089), .ZN(n6980) );
  NAND2_X2 U9888 ( .A1(n10637), .A2(n9282), .ZN(n10626) );
  OR2_X2 U9889 ( .A1(n8798), .A2(n6985), .ZN(n8961) );
  NAND2_X2 U9890 ( .A1(n6986), .A2(n6985), .ZN(n8931) );
  INV_X1 U9891 ( .A(n7434), .ZN(n6988) );
  AOI21_X1 U9892 ( .B1(n7434), .B2(n7436), .A(n6568), .ZN(n6992) );
  NAND2_X1 U9893 ( .A1(n11362), .A2(n7434), .ZN(n6993) );
  OR2_X1 U9894 ( .A1(n6568), .A2(n7436), .ZN(n6994) );
  NAND3_X1 U9895 ( .A1(n6997), .A2(n6996), .A3(n12978), .ZN(n14423) );
  NAND2_X1 U9896 ( .A1(n6999), .A2(n14487), .ZN(n6996) );
  AOI21_X1 U9897 ( .B1(n13334), .B2(n13335), .A(n7023), .ZN(n13260) );
  NAND3_X1 U9898 ( .A1(n7011), .A2(n7012), .A3(n7010), .ZN(n7009) );
  NAND2_X1 U9899 ( .A1(n12229), .A2(n7027), .ZN(n7026) );
  NAND2_X1 U9900 ( .A1(n7274), .A2(n7034), .ZN(n7033) );
  NAND2_X2 U9901 ( .A1(n7033), .A2(n7032), .ZN(n13221) );
  NAND2_X1 U9902 ( .A1(n7036), .A2(n6723), .ZN(n13302) );
  NAND4_X1 U9903 ( .A1(n7941), .A2(n6535), .A3(n7038), .A4(n7942), .ZN(n8610)
         );
  NAND3_X1 U9904 ( .A1(n7941), .A2(n6535), .A3(n8403), .ZN(n8415) );
  NAND2_X1 U9905 ( .A1(n12191), .A2(n7045), .ZN(n7044) );
  NAND3_X1 U9906 ( .A1(n7049), .A2(n12987), .A3(n7048), .ZN(n7335) );
  MUX2_X1 U9907 ( .A(n10645), .B(P2_REG2_REG_2__SCAN_IN), .S(n14262), .Z(
        n14265) );
  NAND2_X1 U9908 ( .A1(n7053), .A2(n7054), .ZN(n10905) );
  NAND2_X1 U9909 ( .A1(n15834), .A2(n6594), .ZN(n7053) );
  AOI21_X1 U9910 ( .B1(n6739), .B2(n7860), .A(n7061), .ZN(n7060) );
  NAND2_X1 U9911 ( .A1(n9288), .A2(n7060), .ZN(n12721) );
  NAND2_X1 U9912 ( .A1(n7860), .A2(n6585), .ZN(n10012) );
  AND2_X1 U9913 ( .A1(n8765), .A2(n7064), .ZN(n7063) );
  NAND2_X1 U9914 ( .A1(n7466), .A2(n8765), .ZN(n9203) );
  NAND3_X1 U9915 ( .A1(n9205), .A2(n12734), .A3(n9204), .ZN(n9207) );
  NAND2_X1 U9916 ( .A1(n7970), .A2(n7971), .ZN(n7342) );
  NAND3_X1 U9917 ( .A1(n7970), .A2(n7473), .A3(n7971), .ZN(n7065) );
  NAND2_X1 U9918 ( .A1(n11375), .A2(n11374), .ZN(n11373) );
  NAND3_X1 U9919 ( .A1(n7067), .A2(n7068), .A3(n6784), .ZN(n7070) );
  INV_X1 U9920 ( .A(n7070), .ZN(n13701) );
  AND2_X1 U9921 ( .A1(n7070), .A2(n13712), .ZN(n13723) );
  INV_X1 U9922 ( .A(n13673), .ZN(n7071) );
  NAND2_X1 U9923 ( .A1(n11618), .A2(n7078), .ZN(n7080) );
  INV_X1 U9924 ( .A(n7073), .ZN(n7072) );
  NOR2_X1 U9925 ( .A1(n7079), .A2(n11145), .ZN(n7078) );
  INV_X1 U9926 ( .A(n10074), .ZN(n7079) );
  NAND2_X1 U9927 ( .A1(n10075), .A2(n7083), .ZN(n7082) );
  NAND2_X1 U9928 ( .A1(n11682), .A2(n10072), .ZN(n7094) );
  NAND2_X1 U9929 ( .A1(n8937), .A2(n7099), .ZN(n7098) );
  NAND2_X1 U9930 ( .A1(n7101), .A2(n7100), .ZN(n8937) );
  NAND3_X1 U9931 ( .A1(n8701), .A2(n8708), .A3(n8700), .ZN(n7101) );
  NAND2_X1 U9932 ( .A1(n9474), .A2(n7947), .ZN(n8899) );
  OAI21_X2 U9933 ( .B1(n8694), .B2(n8899), .A(n7945), .ZN(n8845) );
  OR2_X1 U9934 ( .A1(n8706), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9474) );
  NAND2_X1 U9935 ( .A1(n8719), .A2(n8718), .ZN(n8988) );
  AOI21_X2 U9936 ( .B1(n7112), .B2(n14556), .A(n14322), .ZN(n14581) );
  XNOR2_X1 U9937 ( .A(n14320), .B(n14319), .ZN(n7112) );
  AOI21_X1 U9938 ( .B1(n7119), .B2(n7116), .A(n7115), .ZN(n7114) );
  NAND2_X1 U9939 ( .A1(n14477), .A2(n12864), .ZN(n14475) );
  NOR2_X4 U9940 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n8847) );
  NAND2_X1 U9941 ( .A1(n7132), .A2(n7130), .ZN(n12803) );
  NAND2_X1 U9942 ( .A1(n7131), .A2(n12798), .ZN(n7130) );
  INV_X1 U9943 ( .A(n7134), .ZN(n7131) );
  NAND2_X1 U9944 ( .A1(n7133), .A2(n12796), .ZN(n7132) );
  NAND2_X1 U9945 ( .A1(n7134), .A2(n12797), .ZN(n7133) );
  NAND2_X1 U9946 ( .A1(n8054), .A2(n8053), .ZN(n7134) );
  OAI211_X1 U9947 ( .C1(n7145), .C2(n7143), .A(n8047), .B(n7142), .ZN(n7263)
         );
  NAND3_X1 U9948 ( .A1(n7145), .A2(n8040), .A3(n7144), .ZN(n7142) );
  NAND3_X1 U9949 ( .A1(n8042), .A2(n8041), .A3(n7144), .ZN(n7143) );
  NAND2_X1 U9950 ( .A1(n7146), .A2(n6734), .ZN(n7145) );
  NAND2_X1 U9951 ( .A1(n7147), .A2(n12952), .ZN(n7146) );
  NAND3_X1 U9952 ( .A1(n12929), .A2(n12928), .A3(n12986), .ZN(n7147) );
  XNOR2_X2 U9953 ( .A(n7148), .B(P2_IR_REG_22__SCAN_IN), .ZN(n12763) );
  NAND2_X1 U9954 ( .A1(n7159), .A2(n12903), .ZN(n7154) );
  NAND2_X1 U9955 ( .A1(n12904), .A2(n12905), .ZN(n7159) );
  NAND3_X1 U9956 ( .A1(n7151), .A2(n7149), .A3(n12907), .ZN(n7156) );
  NAND3_X1 U9957 ( .A1(n7154), .A2(n7153), .A3(n12908), .ZN(n7155) );
  INV_X1 U9958 ( .A(n8036), .ZN(n7158) );
  OAI21_X1 U9959 ( .B1(n8062), .B2(n8066), .A(n8064), .ZN(n7162) );
  AND3_X2 U9960 ( .A1(n7164), .A2(n6722), .A3(n7163), .ZN(n15732) );
  NAND3_X1 U9961 ( .A1(n8000), .A2(n7999), .A3(n9550), .ZN(n7166) );
  NAND4_X1 U9962 ( .A1(n8000), .A2(n7999), .A3(n9550), .A4(n9396), .ZN(n7165)
         );
  NAND2_X1 U9963 ( .A1(n7166), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9397) );
  NAND3_X1 U9964 ( .A1(n14760), .A2(n7180), .A3(n9868), .ZN(n7179) );
  NAND2_X1 U9965 ( .A1(n7184), .A2(n6622), .ZN(n9884) );
  AND2_X1 U9966 ( .A1(n7184), .A2(n6601), .ZN(n14845) );
  NAND2_X1 U9967 ( .A1(n8208), .A2(n8207), .ZN(n8211) );
  NAND2_X1 U9968 ( .A1(n8193), .A2(n8192), .ZN(n7191) );
  OAI21_X1 U9969 ( .B1(n8371), .B2(n8382), .A(n7198), .ZN(n8399) );
  NAND2_X1 U9970 ( .A1(n7197), .A2(n7196), .ZN(n7588) );
  NAND2_X1 U9971 ( .A1(n8371), .A2(n7198), .ZN(n7197) );
  NAND2_X1 U9972 ( .A1(n7590), .A2(n7204), .ZN(n7200) );
  NAND2_X1 U9973 ( .A1(n7200), .A2(n7201), .ZN(n8301) );
  NAND2_X1 U9974 ( .A1(n8414), .A2(n7211), .ZN(n7207) );
  NAND2_X1 U9975 ( .A1(n7207), .A2(n7208), .ZN(n8478) );
  NAND2_X1 U9976 ( .A1(n8414), .A2(n8401), .ZN(n7210) );
  NAND2_X1 U9977 ( .A1(n8318), .A2(n7224), .ZN(n7220) );
  NAND2_X1 U9978 ( .A1(n7220), .A2(n7221), .ZN(n8369) );
  NAND2_X1 U9979 ( .A1(n8318), .A2(n8317), .ZN(n7223) );
  NAND3_X1 U9980 ( .A1(n7760), .A2(n7999), .A3(n8000), .ZN(n7227) );
  NAND4_X1 U9981 ( .A1(n7760), .A2(n8000), .A3(n7999), .A4(n9422), .ZN(n15544)
         );
  NAND2_X1 U9982 ( .A1(n7285), .A2(n10540), .ZN(n10542) );
  NAND3_X1 U9983 ( .A1(n7285), .A2(n10540), .A3(n7284), .ZN(n10544) );
  INV_X1 U9984 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7233) );
  INV_X1 U9985 ( .A(n10551), .ZN(n7235) );
  NAND3_X1 U9986 ( .A1(n7235), .A2(n10532), .A3(n7234), .ZN(n10554) );
  INV_X1 U9987 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n7237) );
  NAND2_X1 U9988 ( .A1(n7239), .A2(n11714), .ZN(n11721) );
  NAND2_X1 U9989 ( .A1(n15616), .A2(n15625), .ZN(n7244) );
  NAND3_X1 U9990 ( .A1(n7633), .A2(n7266), .A3(n7246), .ZN(n7240) );
  NAND3_X1 U9991 ( .A1(n7663), .A2(n7661), .A3(n10538), .ZN(n10547) );
  NAND2_X1 U9992 ( .A1(n6742), .A2(n7252), .ZN(n7250) );
  NAND3_X1 U9993 ( .A1(n15565), .A2(n7252), .A3(n15564), .ZN(n7251) );
  NAND2_X1 U9994 ( .A1(n15564), .A2(n15572), .ZN(n7255) );
  AOI21_X1 U9995 ( .B1(n7653), .B2(n7253), .A(n6735), .ZN(n7252) );
  NOR2_X1 U9996 ( .A1(n6712), .A2(n15572), .ZN(n15576) );
  INV_X1 U9997 ( .A(n15605), .ZN(n7643) );
  NAND2_X1 U9998 ( .A1(n10962), .A2(n10961), .ZN(n7257) );
  NOR2_X1 U9999 ( .A1(n6562), .A2(n7654), .ZN(n7653) );
  OAI211_X1 U10000 ( .C1(n11725), .C2(n7649), .A(n15839), .B(n7648), .ZN(n7646) );
  NAND2_X1 U10001 ( .A1(n7825), .A2(n7343), .ZN(n14078) );
  NAND2_X1 U10002 ( .A1(n7829), .A2(n7827), .ZN(n11229) );
  NAND2_X1 U10003 ( .A1(n7263), .A2(n12992), .ZN(P2_U3328) );
  INV_X1 U10004 ( .A(n12723), .ZN(n7279) );
  INV_X1 U10005 ( .A(n14685), .ZN(n7319) );
  OR2_X1 U10006 ( .A1(n11175), .A2(n11186), .ZN(n15718) );
  NOR2_X2 U10007 ( .A1(n12212), .A2(n14778), .ZN(n7988) );
  OAI21_X1 U10008 ( .B1(n15391), .B2(n15390), .A(n7960), .ZN(n15523) );
  NAND2_X1 U10009 ( .A1(n7643), .A2(n7636), .ZN(n7267) );
  NAND3_X1 U10010 ( .A1(n7687), .A2(n11195), .A3(n12430), .ZN(n11347) );
  NAND2_X1 U10011 ( .A1(n8547), .A2(n13522), .ZN(n10041) );
  NAND2_X1 U10012 ( .A1(n11940), .A2(n12641), .ZN(n12205) );
  NAND2_X1 U10013 ( .A1(n7693), .A2(n11578), .ZN(n7695) );
  XNOR2_X1 U10014 ( .A(n15389), .B(n15129), .ZN(n15402) );
  OAI211_X2 U10015 ( .C1(n9779), .C2(n10215), .A(n7462), .B(n6650), .ZN(n7771)
         );
  AOI21_X2 U10016 ( .B1(n10172), .B2(n10173), .A(n10174), .ZN(n10171) );
  NAND3_X1 U10017 ( .A1(n6743), .A2(n7546), .A3(n7548), .ZN(n7330) );
  NOR2_X1 U10018 ( .A1(n6736), .A2(n7691), .ZN(n7690) );
  NAND2_X1 U10019 ( .A1(n15524), .A2(n15791), .ZN(n7454) );
  NAND2_X1 U10020 ( .A1(n7708), .A2(n13064), .ZN(n7707) );
  OAI21_X1 U10021 ( .B1(SI_22_), .B2(n9166), .A(n9179), .ZN(n9833) );
  NAND2_X1 U10022 ( .A1(n15552), .A2(n9475), .ZN(n15223) );
  NAND2_X1 U10023 ( .A1(n8211), .A2(n8210), .ZN(n8225) );
  NAND2_X1 U10024 ( .A1(n8495), .A2(n8494), .ZN(n8505) );
  NAND2_X1 U10025 ( .A1(n7348), .A2(n8162), .ZN(n8173) );
  OAI21_X1 U10026 ( .B1(n8478), .B2(n8477), .A(n8479), .ZN(n8482) );
  NAND2_X1 U10027 ( .A1(n6653), .A2(n7677), .ZN(n7676) );
  AOI21_X1 U10028 ( .B1(n13269), .B2(n13575), .A(n10025), .ZN(n8664) );
  NAND2_X2 U10029 ( .A1(n7270), .A2(n7269), .ZN(n14824) );
  NAND2_X1 U10030 ( .A1(n8482), .A2(n8481), .ZN(n8495) );
  NAND2_X1 U10031 ( .A1(n8303), .A2(n8302), .ZN(n8318) );
  NAND2_X1 U10032 ( .A1(n7588), .A2(n8400), .ZN(n8414) );
  OAI22_X1 U10033 ( .A1(n15341), .A2(n15320), .B1(n12498), .B2(n15479), .ZN(
        n13014) );
  NAND2_X1 U10034 ( .A1(n7301), .A2(n7300), .ZN(n7272) );
  NAND2_X2 U10035 ( .A1(n15212), .A2(n15214), .ZN(n15211) );
  NAND2_X1 U10036 ( .A1(n6589), .A2(n7283), .ZN(n7282) );
  OAI22_X2 U10037 ( .A1(n13280), .A2(n13281), .B1(n13222), .B2(n13790), .ZN(
        n13334) );
  INV_X1 U10038 ( .A(n13250), .ZN(n7274) );
  AOI21_X1 U10039 ( .B1(n7281), .B2(n12036), .A(n6577), .ZN(n7381) );
  AND2_X1 U10040 ( .A1(n8141), .A2(n8140), .ZN(n7277) );
  NAND2_X1 U10041 ( .A1(n13302), .A2(n12679), .ZN(n13328) );
  OAI211_X1 U10042 ( .C1(n13239), .C2(n7928), .A(n7927), .B(n11860), .ZN(
        n11837) );
  NAND2_X1 U10043 ( .A1(n13326), .A2(n12682), .ZN(n13250) );
  INV_X1 U10044 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7284) );
  INV_X1 U10045 ( .A(n9005), .ZN(n7278) );
  NAND2_X1 U10046 ( .A1(n9414), .A2(n9412), .ZN(n9434) );
  AOI21_X1 U10047 ( .B1(n14958), .B2(n9936), .A(n9481), .ZN(n10184) );
  INV_X1 U10048 ( .A(n11845), .ZN(n7281) );
  NAND2_X1 U10049 ( .A1(n7289), .A2(n7381), .ZN(n12298) );
  INV_X1 U10050 ( .A(n11597), .ZN(n11598) );
  INV_X1 U10051 ( .A(n11577), .ZN(n7698) );
  NAND3_X1 U10052 ( .A1(n8591), .A2(n7282), .A3(n7369), .ZN(n14027) );
  OAI211_X1 U10053 ( .C1(n13528), .C2(n15917), .A(n13563), .B(n7332), .ZN(
        n7801) );
  NAND2_X1 U10054 ( .A1(n7287), .A2(n7286), .ZN(n7285) );
  INV_X1 U10055 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7286) );
  OR2_X1 U10056 ( .A1(n12869), .A2(n12868), .ZN(n12870) );
  NAND2_X1 U10057 ( .A1(n7931), .A2(n11810), .ZN(n7930) );
  NAND2_X1 U10058 ( .A1(n13328), .A2(n13327), .ZN(n13326) );
  NAND2_X1 U10059 ( .A1(n12671), .A2(n12670), .ZN(n13342) );
  BUF_X1 U10060 ( .A(n13717), .Z(n7288) );
  NAND2_X1 U10061 ( .A1(n12298), .A2(n12226), .ZN(n12229) );
  NAND2_X1 U10062 ( .A1(n11814), .A2(n11815), .ZN(n12077) );
  NAND3_X1 U10063 ( .A1(n13208), .A2(n13207), .A3(n6770), .ZN(P2_U3186) );
  NAND2_X1 U10064 ( .A1(n8068), .A2(n6737), .ZN(n13084) );
  NAND2_X1 U10065 ( .A1(n12663), .A2(n7295), .ZN(P1_U3242) );
  NAND3_X1 U10066 ( .A1(n12558), .A2(n12557), .A3(n6728), .ZN(n7297) );
  MUX2_X1 U10067 ( .A(n14950), .B(n15497), .S(n6549), .Z(n12491) );
  INV_X1 U10068 ( .A(n7361), .ZN(n8498) );
  OAI21_X1 U10069 ( .B1(n13899), .B2(n15903), .A(n7675), .ZN(P3_U3204) );
  NAND2_X1 U10070 ( .A1(n12131), .A2(n12132), .ZN(n12270) );
  NAND2_X2 U10071 ( .A1(n8820), .A2(n8819), .ZN(n14615) );
  NAND2_X1 U10072 ( .A1(n10020), .A2(n9372), .ZN(n7772) );
  NAND2_X1 U10073 ( .A1(n7279), .A2(n11417), .ZN(n9379) );
  INV_X1 U10074 ( .A(n15156), .ZN(n7458) );
  OAI21_X1 U10075 ( .B1(n7975), .B2(n7458), .A(n6718), .ZN(n7457) );
  NAND2_X1 U10076 ( .A1(n11576), .A2(n15671), .ZN(n7699) );
  OAI22_X1 U10077 ( .A1(n7698), .A2(n7699), .B1(n15684), .B2(n11579), .ZN(
        n7697) );
  NAND2_X1 U10078 ( .A1(n8864), .A2(n8703), .ZN(n8920) );
  AOI21_X1 U10079 ( .B1(n7801), .B2(n13564), .A(n7804), .ZN(n7800) );
  AOI21_X1 U10080 ( .B1(n7962), .B2(n15783), .A(n7961), .ZN(n7960) );
  NAND2_X1 U10081 ( .A1(n15523), .A2(n15791), .ZN(n7959) );
  OR4_X2 U10082 ( .A1(n13543), .A2(n6889), .A3(n13542), .A4(n13541), .ZN(
        n13546) );
  NAND3_X1 U10083 ( .A1(n13535), .A2(n13534), .A3(n7307), .ZN(n7306) );
  NAND3_X1 U10084 ( .A1(n13869), .A2(n13548), .A3(n7311), .ZN(n7310) );
  NAND2_X1 U10085 ( .A1(n15949), .A2(n13586), .ZN(n13439) );
  NAND2_X1 U10086 ( .A1(n11837), .A2(n11836), .ZN(n11845) );
  NAND2_X1 U10087 ( .A1(n7660), .A2(n10936), .ZN(n7657) );
  INV_X1 U10088 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n7314) );
  INV_X1 U10089 ( .A(n10541), .ZN(n7315) );
  NAND3_X1 U10090 ( .A1(n7695), .A2(n7382), .A3(n11580), .ZN(n11939) );
  NAND2_X1 U10091 ( .A1(n15186), .A2(n15185), .ZN(n15184) );
  NAND2_X1 U10092 ( .A1(n11165), .A2(n12440), .ZN(n7689) );
  NAND2_X1 U10093 ( .A1(n7688), .A2(n12426), .ZN(n15707) );
  NAND2_X1 U10094 ( .A1(n8706), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7584) );
  INV_X4 U10095 ( .A(n7395), .ZN(n8706) );
  NAND2_X2 U10096 ( .A1(n7465), .A2(n7463), .ZN(n7395) );
  NAND3_X1 U10097 ( .A1(n14578), .A2(n14577), .A3(n14579), .ZN(n7431) );
  NAND2_X1 U10098 ( .A1(n6677), .A2(n7318), .ZN(P2_U3525) );
  NAND2_X1 U10099 ( .A1(n14684), .A2(n7320), .ZN(P2_U3493) );
  NAND2_X1 U10100 ( .A1(n8791), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n9186) );
  NAND2_X1 U10101 ( .A1(n8792), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n9195) );
  INV_X1 U10102 ( .A(n8048), .ZN(n8042) );
  OAI21_X2 U10103 ( .B1(n13173), .B2(n8961), .A(n9255), .ZN(n14218) );
  NAND2_X1 U10104 ( .A1(n11782), .A2(n11783), .ZN(n11807) );
  NAND2_X1 U10105 ( .A1(n6711), .A2(n7671), .ZN(n8117) );
  NAND3_X1 U10106 ( .A1(n7331), .A2(n13756), .A3(n7330), .ZN(P3_U3201) );
  NAND2_X1 U10107 ( .A1(n13755), .A2(n13754), .ZN(n7331) );
  NAND2_X1 U10108 ( .A1(n11962), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n11961) );
  AOI21_X1 U10109 ( .B1(n13729), .B2(n13728), .A(n13727), .ZN(n13752) );
  INV_X1 U10110 ( .A(n10077), .ZN(n7354) );
  NAND2_X1 U10111 ( .A1(n7354), .A2(n7353), .ZN(n10078) );
  AND2_X2 U10112 ( .A1(n6658), .A2(n6574), .ZN(n8000) );
  AOI21_X2 U10113 ( .B1(n14893), .B2(n14892), .A(n6688), .ZN(n14808) );
  NAND2_X1 U10114 ( .A1(n8778), .A2(n8777), .ZN(n7443) );
  AOI21_X1 U10115 ( .B1(n15814), .B2(n10667), .A(n10666), .ZN(n10665) );
  NOR3_X1 U10116 ( .A1(n11002), .A2(n11001), .A3(n11004), .ZN(n11538) );
  NAND3_X1 U10117 ( .A1(n13141), .A2(n14123), .A3(n14124), .ZN(n7825) );
  NAND2_X1 U10118 ( .A1(n12724), .A2(n12725), .ZN(n9486) );
  XNOR2_X1 U10119 ( .A(n9483), .B(n9482), .ZN(n12724) );
  NAND2_X1 U10120 ( .A1(n12886), .A2(n12885), .ZN(n8067) );
  NAND2_X1 U10121 ( .A1(n7652), .A2(n10952), .ZN(n10962) );
  NAND2_X1 U10122 ( .A1(n12288), .A2(n12287), .ZN(n7665) );
  AOI21_X1 U10123 ( .B1(n12900), .B2(n8037), .A(n8038), .ZN(n8036) );
  NAND3_X1 U10124 ( .A1(n7604), .A2(n7603), .A3(n8160), .ZN(n7348) );
  NAND2_X1 U10125 ( .A1(n7618), .A2(n8521), .ZN(n8535) );
  INV_X1 U10126 ( .A(n13899), .ZN(n7367) );
  NAND2_X1 U10127 ( .A1(n8691), .A2(n7364), .ZN(P3_U3456) );
  NAND2_X1 U10128 ( .A1(n7349), .A2(n15386), .ZN(n15391) );
  NAND3_X1 U10129 ( .A1(n15389), .A2(n15384), .A3(n15387), .ZN(n7349) );
  INV_X1 U10130 ( .A(P2_RD_REG_SCAN_IN), .ZN(n10250) );
  INV_X1 U10131 ( .A(n9139), .ZN(n7573) );
  NAND2_X1 U10132 ( .A1(n7497), .A2(n7501), .ZN(n9137) );
  NAND2_X1 U10133 ( .A1(n8582), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8134) );
  XNOR2_X2 U10134 ( .A(n7355), .B(n8142), .ZN(n11295) );
  NAND3_X1 U10135 ( .A1(n12272), .A2(n7664), .A3(n12271), .ZN(n12288) );
  NAND2_X1 U10136 ( .A1(n9523), .A2(n9539), .ZN(n15635) );
  NAND2_X1 U10137 ( .A1(n8845), .A2(n8696), .ZN(n8837) );
  NAND2_X1 U10138 ( .A1(n10825), .A2(n10826), .ZN(n7878) );
  NAND2_X1 U10139 ( .A1(n11999), .A2(n6724), .ZN(n11868) );
  INV_X1 U10140 ( .A(n11112), .ZN(n9977) );
  NAND2_X1 U10141 ( .A1(n8263), .A2(n8262), .ZN(n8280) );
  NAND2_X1 U10142 ( .A1(n7373), .A2(n7370), .ZN(P1_U3240) );
  NAND2_X1 U10143 ( .A1(n14911), .A2(n14910), .ZN(n7373) );
  AOI21_X2 U10144 ( .B1(n14824), .B2(n9764), .A(n9763), .ZN(n14836) );
  AND2_X1 U10145 ( .A1(n11048), .A2(n11227), .ZN(n11049) );
  NAND2_X1 U10146 ( .A1(n9121), .A2(n8808), .ZN(n8810) );
  NAND2_X1 U10147 ( .A1(n13702), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n13729) );
  NOR2_X1 U10148 ( .A1(n13752), .A2(n13751), .ZN(n7623) );
  XNOR2_X1 U10149 ( .A(n7623), .B(n7622), .ZN(n13755) );
  NAND2_X1 U10150 ( .A1(n9033), .A2(n9032), .ZN(n9035) );
  NAND2_X1 U10151 ( .A1(n7959), .A2(n7958), .ZN(P1_U3525) );
  INV_X1 U10152 ( .A(n7987), .ZN(n7986) );
  NAND2_X1 U10153 ( .A1(n7454), .A2(n7453), .ZN(P1_U3524) );
  OAI21_X1 U10154 ( .B1(n13717), .B2(P3_REG2_REG_1__SCAN_IN), .A(n7379), .ZN(
        n10089) );
  XNOR2_X1 U10155 ( .A(n12695), .B(n13539), .ZN(n11839) );
  INV_X1 U10156 ( .A(n7697), .ZN(n7382) );
  NAND2_X1 U10157 ( .A1(n12637), .A2(n11572), .ZN(n11577) );
  NAND2_X4 U10158 ( .A1(n14038), .A2(n13717), .ZN(n10063) );
  NAND2_X1 U10159 ( .A1(n6606), .A2(n7388), .ZN(n7389) );
  NAND3_X1 U10160 ( .A1(n7390), .A2(n8641), .A3(n7389), .ZN(n8643) );
  NAND3_X1 U10161 ( .A1(n6606), .A2(n8635), .A3(n7391), .ZN(n7390) );
  NAND2_X1 U10162 ( .A1(n7392), .A2(n8636), .ZN(n7670) );
  INV_X1 U10163 ( .A(n8638), .ZN(n7393) );
  INV_X1 U10164 ( .A(n8846), .ZN(n8696) );
  XNOR2_X1 U10165 ( .A(n8697), .B(SI_2_), .ZN(n8846) );
  MUX2_X1 U10166 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n7395), .Z(n8697) );
  INV_X1 U10167 ( .A(n8703), .ZN(n7396) );
  NAND2_X1 U10168 ( .A1(n7406), .A2(n7407), .ZN(n13774) );
  INV_X1 U10169 ( .A(n14378), .ZN(n7411) );
  NAND2_X1 U10170 ( .A1(n13835), .A2(n7419), .ZN(n7418) );
  NAND2_X1 U10171 ( .A1(n13835), .A2(n8088), .ZN(n13823) );
  INV_X1 U10172 ( .A(n7418), .ZN(n13822) );
  INV_X1 U10173 ( .A(n8088), .ZN(n7420) );
  MUX2_X1 U10174 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n7431), .S(n15893), .Z(
        P2_U3526) );
  MUX2_X1 U10175 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n7431), .S(n15886), .Z(
        P2_U3494) );
  AND2_X1 U10176 ( .A1(n8906), .A2(n8905), .ZN(n7437) );
  NAND4_X1 U10177 ( .A1(n8811), .A2(n8813), .A3(n8779), .A4(n6719), .ZN(n7442)
         );
  NAND2_X1 U10178 ( .A1(n9370), .A2(n9369), .ZN(n14318) );
  NAND2_X1 U10179 ( .A1(n9370), .A2(n7444), .ZN(n7583) );
  NAND2_X1 U10180 ( .A1(n7446), .A2(n14309), .ZN(n14573) );
  NAND2_X1 U10181 ( .A1(n12202), .A2(n11949), .ZN(n11951) );
  OAI211_X2 U10182 ( .C1(n15676), .C2(n7447), .A(n7448), .B(n12208), .ZN(
        n12202) );
  NAND2_X1 U10183 ( .A1(n7452), .A2(n7451), .ZN(n12203) );
  NAND2_X1 U10184 ( .A1(n15676), .A2(n11569), .ZN(n7452) );
  NAND2_X1 U10185 ( .A1(n7451), .A2(n7449), .ZN(n7448) );
  OAI211_X2 U10186 ( .C1(n15369), .C2(n13013), .A(n13017), .B(n13016), .ZN(
        n15321) );
  INV_X1 U10187 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n15114) );
  INV_X1 U10188 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7464) );
  INV_X1 U10189 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n14302) );
  NAND4_X1 U10190 ( .A1(n10250), .A2(n7464), .A3(P2_ADDR_REG_19__SCAN_IN), 
        .A4(P1_ADDR_REG_19__SCAN_IN), .ZN(n7463) );
  NAND4_X1 U10191 ( .A1(n15114), .A2(n10207), .A3(n14302), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7465) );
  NAND2_X1 U10192 ( .A1(n7468), .A2(SI_24_), .ZN(n8765) );
  NAND3_X1 U10193 ( .A1(n7470), .A2(n12652), .A3(n12653), .ZN(n7469) );
  NAND3_X1 U10194 ( .A1(n7478), .A2(n8744), .A3(n8749), .ZN(n7472) );
  INV_X1 U10195 ( .A(n7478), .ZN(n7477) );
  NAND2_X1 U10196 ( .A1(n6600), .A2(n9079), .ZN(n7478) );
  NAND2_X1 U10197 ( .A1(n9262), .A2(n7480), .ZN(n7479) );
  NAND2_X1 U10198 ( .A1(n9262), .A2(n9261), .ZN(n12591) );
  NAND2_X1 U10199 ( .A1(n8806), .A2(n7503), .ZN(n7499) );
  OR2_X1 U10200 ( .A1(n8806), .A2(n7504), .ZN(n7497) );
  OAI21_X1 U10201 ( .B1(n9210), .B2(n9209), .A(n7512), .ZN(n9234) );
  NAND3_X1 U10202 ( .A1(n7521), .A2(n7520), .A3(n7518), .ZN(n10596) );
  NAND2_X1 U10203 ( .A1(n7514), .A2(n14982), .ZN(n7520) );
  OR2_X1 U10204 ( .A1(n14982), .A2(n14978), .ZN(n7524) );
  MUX2_X1 U10205 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9457), .S(n10488), .Z(
        n14963) );
  NAND3_X1 U10206 ( .A1(n7542), .A2(n6774), .A3(n7543), .ZN(n7544) );
  NAND2_X1 U10207 ( .A1(n11308), .A2(n6775), .ZN(n7542) );
  INV_X1 U10208 ( .A(n7544), .ZN(n10059) );
  NAND3_X1 U10209 ( .A1(n7554), .A2(n6569), .A3(n7547), .ZN(n7546) );
  NAND3_X1 U10210 ( .A1(n7561), .A2(n13663), .A3(n6598), .ZN(n7560) );
  INV_X1 U10211 ( .A(n13643), .ZN(n7558) );
  NAND3_X1 U10212 ( .A1(n7559), .A2(n7562), .A3(n7560), .ZN(n13687) );
  NAND2_X1 U10213 ( .A1(n7561), .A2(n13663), .ZN(n13644) );
  OR2_X1 U10214 ( .A1(n13693), .A2(n13686), .ZN(n7562) );
  NAND2_X1 U10215 ( .A1(n7563), .A2(n10130), .ZN(n13642) );
  NAND2_X1 U10216 ( .A1(n7565), .A2(n7564), .ZN(n7563) );
  INV_X1 U10217 ( .A(n10062), .ZN(n7564) );
  NAND2_X1 U10218 ( .A1(n7569), .A2(n11684), .ZN(n7567) );
  NAND2_X1 U10219 ( .A1(n8188), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7571) );
  OAI21_X2 U10220 ( .B1(n14309), .B2(n7577), .A(n6684), .ZN(n7576) );
  NAND2_X1 U10221 ( .A1(n7579), .A2(n7581), .ZN(n10021) );
  NAND2_X1 U10222 ( .A1(n14318), .A2(n7582), .ZN(n7579) );
  OAI21_X2 U10223 ( .B1(n8706), .B2(n7585), .A(n7584), .ZN(n8705) );
  INV_X1 U10224 ( .A(n14605), .ZN(n14420) );
  NAND2_X2 U10225 ( .A1(n7587), .A2(n9156), .ZN(n14605) );
  OAI21_X1 U10226 ( .B1(n8225), .B2(n7593), .A(n7591), .ZN(n8249) );
  NAND2_X1 U10227 ( .A1(n8225), .A2(n7591), .ZN(n7590) );
  OAI21_X1 U10228 ( .B1(n8225), .B2(n8224), .A(n8223), .ZN(n8235) );
  NAND2_X1 U10229 ( .A1(n8152), .A2(n8144), .ZN(n7603) );
  NAND2_X1 U10230 ( .A1(n8153), .A2(n8152), .ZN(n8161) );
  NAND2_X1 U10231 ( .A1(n7606), .A2(n7605), .ZN(n8153) );
  NAND2_X1 U10232 ( .A1(n13595), .A2(n11679), .ZN(n10071) );
  NAND2_X1 U10233 ( .A1(n11139), .A2(n10167), .ZN(n10075) );
  NAND2_X1 U10234 ( .A1(n10149), .A2(n7630), .ZN(n11306) );
  XNOR2_X1 U10235 ( .A(n13657), .B(n7380), .ZN(n13658) );
  NAND2_X1 U10236 ( .A1(n15605), .A2(n6700), .ZN(n7633) );
  NAND2_X1 U10237 ( .A1(n15605), .A2(n15604), .ZN(n15607) );
  OR2_X1 U10238 ( .A1(n15604), .A2(n7645), .ZN(n7644) );
  INV_X1 U10239 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n7645) );
  NAND2_X1 U10240 ( .A1(n11725), .A2(n11724), .ZN(n7650) );
  NAND2_X1 U10241 ( .A1(n11725), .A2(n7647), .ZN(n12126) );
  AND2_X1 U10242 ( .A1(n11724), .A2(n7649), .ZN(n7647) );
  OR2_X1 U10243 ( .A1(n11724), .A2(n7649), .ZN(n7648) );
  INV_X1 U10244 ( .A(n11735), .ZN(n7649) );
  NAND2_X1 U10245 ( .A1(n7650), .A2(n11735), .ZN(n12125) );
  NAND2_X1 U10246 ( .A1(n15556), .A2(n15557), .ZN(n7652) );
  NAND2_X1 U10247 ( .A1(n7652), .A2(n6716), .ZN(n11714) );
  INV_X1 U10248 ( .A(n6636), .ZN(n15593) );
  INV_X1 U10249 ( .A(n15592), .ZN(n7656) );
  NAND2_X1 U10250 ( .A1(n7657), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n7658) );
  NAND3_X1 U10251 ( .A1(n7660), .A2(n7659), .A3(n10936), .ZN(n10937) );
  NAND2_X1 U10252 ( .A1(n10937), .A2(n7658), .ZN(n10571) );
  INV_X1 U10253 ( .A(n10571), .ZN(n10568) );
  INV_X1 U10254 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7659) );
  NAND2_X1 U10255 ( .A1(n7662), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n10546) );
  NAND2_X1 U10256 ( .A1(n12272), .A2(n12271), .ZN(n12280) );
  NOR2_X1 U10257 ( .A1(n8578), .A2(P3_IR_REG_28__SCAN_IN), .ZN(n7671) );
  AOI21_X2 U10258 ( .B1(n8675), .B2(n13960), .A(n8674), .ZN(n13899) );
  NAND2_X1 U10259 ( .A1(n15707), .A2(n11194), .ZN(n7687) );
  INV_X1 U10260 ( .A(n7699), .ZN(n7693) );
  OR2_X1 U10261 ( .A1(n9608), .A2(n9487), .ZN(n9493) );
  AND2_X1 U10263 ( .A1(n7715), .A2(n7724), .ZN(n7714) );
  NAND2_X1 U10264 ( .A1(n7717), .A2(n7716), .ZN(n7715) );
  NAND2_X1 U10265 ( .A1(n7728), .A2(n7722), .ZN(n7720) );
  NAND2_X1 U10266 ( .A1(n7723), .A2(n12504), .ZN(n12514) );
  NAND2_X1 U10267 ( .A1(n12604), .A2(n7735), .ZN(n7729) );
  NAND2_X1 U10268 ( .A1(n7729), .A2(n6706), .ZN(n12660) );
  NAND3_X1 U10269 ( .A1(n12606), .A2(n12653), .A3(n12605), .ZN(n7741) );
  NAND2_X1 U10270 ( .A1(n14537), .A2(n7744), .ZN(n7742) );
  NAND2_X1 U10271 ( .A1(n7742), .A2(n7743), .ZN(n14498) );
  INV_X1 U10272 ( .A(n9357), .ZN(n7746) );
  NAND2_X1 U10273 ( .A1(n12477), .A2(n7750), .ZN(n7747) );
  OAI21_X1 U10274 ( .B1(n12477), .B2(n7751), .A(n7750), .ZN(n12482) );
  NAND2_X1 U10275 ( .A1(n7747), .A2(n7748), .ZN(n12481) );
  AOI21_X1 U10276 ( .B1(n7751), .B2(n7750), .A(n7749), .ZN(n7748) );
  INV_X1 U10277 ( .A(n12483), .ZN(n7749) );
  NOR2_X1 U10278 ( .A1(n12479), .A2(n12476), .ZN(n7751) );
  INV_X1 U10279 ( .A(n7756), .ZN(n7758) );
  NAND2_X1 U10280 ( .A1(n12543), .A2(n7759), .ZN(n7752) );
  NAND2_X1 U10281 ( .A1(n7754), .A2(n7753), .ZN(n12547) );
  NAND2_X1 U10282 ( .A1(n7758), .A2(n12544), .ZN(n7753) );
  NAND2_X1 U10283 ( .A1(n12541), .A2(n7755), .ZN(n7754) );
  NAND2_X1 U10284 ( .A1(n7756), .A2(n7757), .ZN(n7755) );
  INV_X1 U10285 ( .A(n12540), .ZN(n7759) );
  NAND2_X1 U10286 ( .A1(n12563), .A2(n12564), .ZN(n12562) );
  NAND2_X1 U10287 ( .A1(n7765), .A2(n7766), .ZN(n12556) );
  NAND2_X1 U10288 ( .A1(n7768), .A2(n7770), .ZN(n12469) );
  NAND3_X1 U10289 ( .A1(n12458), .A2(n12457), .A3(n7769), .ZN(n7768) );
  NAND3_X1 U10290 ( .A1(n9513), .A2(n7771), .A3(n6617), .ZN(n12430) );
  NAND2_X1 U10291 ( .A1(n15907), .A2(n8632), .ZN(n13959) );
  NAND2_X1 U10292 ( .A1(n8643), .A2(n8642), .ZN(n12049) );
  OR2_X1 U10293 ( .A1(n8653), .A2(n12384), .ZN(n8655) );
  OR2_X1 U10294 ( .A1(n8656), .A2(n13883), .ZN(n8658) );
  NAND2_X1 U10295 ( .A1(n12485), .A2(n12484), .ZN(n12490) );
  NAND2_X1 U10296 ( .A1(n8663), .A2(n8004), .ZN(n13835) );
  NAND2_X1 U10297 ( .A1(n11546), .A2(n12964), .ZN(n11548) );
  NAND2_X1 U10298 ( .A1(n14489), .A2(n14488), .ZN(n14487) );
  AOI21_X1 U10299 ( .B1(n14498), .B2(n14501), .A(n9358), .ZN(n14489) );
  NAND2_X1 U10300 ( .A1(n13426), .A2(n13534), .ZN(n7774) );
  NAND3_X1 U10301 ( .A1(n11523), .A2(n13534), .A3(n11524), .ZN(n7775) );
  OR2_X1 U10302 ( .A1(n10063), .A2(n10093), .ZN(n7776) );
  INV_X1 U10303 ( .A(n8105), .ZN(n7779) );
  NAND2_X1 U10304 ( .A1(n13398), .A2(n13564), .ZN(n7802) );
  OAI21_X1 U10305 ( .B1(n7803), .B2(n7802), .A(n7800), .ZN(P3_U3296) );
  NAND2_X1 U10306 ( .A1(n8381), .A2(n7808), .ZN(n7805) );
  NAND2_X1 U10307 ( .A1(n7805), .A2(n7806), .ZN(n13829) );
  NAND2_X1 U10308 ( .A1(n10860), .A2(n10859), .ZN(n7819) );
  AND2_X1 U10309 ( .A1(n7816), .A2(n7817), .ZN(n7815) );
  NAND2_X1 U10310 ( .A1(n10881), .A2(n7819), .ZN(n10882) );
  NAND2_X1 U10311 ( .A1(n11038), .A2(n7830), .ZN(n7829) );
  AOI21_X1 U10312 ( .B1(n7830), .B2(n11037), .A(n7828), .ZN(n7827) );
  AND2_X1 U10313 ( .A1(n11049), .A2(n11043), .ZN(n7830) );
  AND3_X2 U10314 ( .A1(n8774), .A2(n8776), .A3(n8775), .ZN(n8811) );
  NAND2_X1 U10315 ( .A1(n14098), .A2(n13161), .ZN(n14190) );
  NOR2_X1 U10316 ( .A1(n14191), .A2(n13160), .ZN(n7838) );
  NAND2_X1 U10317 ( .A1(n8814), .A2(n7840), .ZN(n9272) );
  NAND2_X1 U10318 ( .A1(n6741), .A2(n8814), .ZN(n7841) );
  INV_X1 U10319 ( .A(n9302), .ZN(n8767) );
  INV_X1 U10320 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9315) );
  NAND3_X1 U10321 ( .A1(n8778), .A2(n8782), .A3(n8777), .ZN(n7849) );
  NAND4_X1 U10322 ( .A1(n8778), .A2(n8777), .A3(n8811), .A4(n8813), .ZN(n9305)
         );
  NOR2_X1 U10323 ( .A1(n12973), .A2(n7856), .ZN(n7855) );
  NAND2_X1 U10324 ( .A1(n14320), .A2(n7861), .ZN(n7860) );
  NAND2_X1 U10325 ( .A1(n7860), .A2(n7863), .ZN(n10011) );
  AOI21_X1 U10326 ( .B1(n14320), .B2(n12957), .A(n12956), .ZN(n14304) );
  NAND2_X1 U10327 ( .A1(n14610), .A2(n9361), .ZN(n7877) );
  NAND2_X1 U10328 ( .A1(n8000), .A2(n9550), .ZN(n9404) );
  NAND2_X1 U10329 ( .A1(n9797), .A2(n9796), .ZN(n7899) );
  NAND2_X1 U10330 ( .A1(n9884), .A2(n7904), .ZN(n7903) );
  NAND2_X1 U10331 ( .A1(n14816), .A2(n6618), .ZN(n7905) );
  INV_X1 U10332 ( .A(n14817), .ZN(n7907) );
  OR2_X1 U10333 ( .A1(n8902), .A2(n10595), .ZN(n8903) );
  CLKBUF_X1 U10334 ( .A(n7912), .Z(n7909) );
  INV_X1 U10335 ( .A(n7909), .ZN(n14429) );
  NAND2_X1 U10336 ( .A1(n14323), .A2(n6624), .ZN(n12752) );
  AND2_X1 U10337 ( .A1(n14323), .A2(n14307), .ZN(n10014) );
  AND2_X2 U10338 ( .A1(n14522), .A2(n7915), .ZN(n14455) );
  INV_X1 U10339 ( .A(n7920), .ZN(n14467) );
  INV_X1 U10340 ( .A(n12077), .ZN(n7931) );
  NAND2_X1 U10341 ( .A1(n7930), .A2(n11815), .ZN(n7927) );
  INV_X1 U10342 ( .A(n11815), .ZN(n7928) );
  NAND2_X1 U10343 ( .A1(n12075), .A2(n11815), .ZN(n11859) );
  NAND2_X1 U10344 ( .A1(n13239), .A2(n7929), .ZN(n12075) );
  NAND2_X1 U10345 ( .A1(n12694), .A2(n7933), .ZN(n7932) );
  OAI211_X1 U10346 ( .C1(n12694), .C2(n7934), .A(n12699), .B(n7932), .ZN(
        P3_U3169) );
  XNOR2_X1 U10347 ( .A(n12694), .B(n12693), .ZN(n13232) );
  INV_X1 U10348 ( .A(n13309), .ZN(n7940) );
  NAND2_X1 U10349 ( .A1(n8712), .A2(n10487), .ZN(n7946) );
  NAND2_X1 U10350 ( .A1(n7970), .A2(n7968), .ZN(n9059) );
  INV_X1 U10351 ( .A(n11186), .ZN(n15743) );
  NAND3_X1 U10352 ( .A1(n11425), .A2(n12414), .A3(n7991), .ZN(n15677) );
  AND2_X2 U10353 ( .A1(n15717), .A2(n11431), .ZN(n11425) );
  NAND2_X1 U10354 ( .A1(n15159), .A2(n7996), .ZN(n15115) );
  NAND2_X1 U10355 ( .A1(n15159), .A2(n15407), .ZN(n15148) );
  NOR2_X2 U10356 ( .A1(n15148), .A2(n7998), .ZN(n15122) );
  NOR2_X2 U10357 ( .A1(n9400), .A2(n9393), .ZN(n7999) );
  NAND3_X1 U10358 ( .A1(n9406), .A2(n9390), .A3(n9389), .ZN(n9400) );
  INV_X1 U10359 ( .A(n11778), .ZN(n15905) );
  INV_X1 U10360 ( .A(n8008), .ZN(n8007) );
  NAND2_X1 U10361 ( .A1(n8009), .A2(n6608), .ZN(n8008) );
  INV_X1 U10362 ( .A(n13424), .ZN(n8016) );
  INV_X1 U10363 ( .A(n13473), .ZN(n8028) );
  INV_X1 U10364 ( .A(n13474), .ZN(n8029) );
  NAND2_X1 U10365 ( .A1(n9283), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8935) );
  NAND2_X1 U10366 ( .A1(n9283), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n9219) );
  NAND2_X1 U10367 ( .A1(n9283), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9227) );
  NAND3_X1 U10368 ( .A1(n12789), .A2(n12790), .A3(n8055), .ZN(n8054) );
  AOI21_X1 U10369 ( .B1(n12894), .B2(n8059), .A(n8057), .ZN(n8056) );
  NAND2_X1 U10370 ( .A1(n8065), .A2(n8063), .ZN(n12888) );
  INV_X1 U10371 ( .A(n8781), .ZN(n8068) );
  NAND2_X1 U10372 ( .A1(n12803), .A2(n8070), .ZN(n8069) );
  INV_X1 U10373 ( .A(n12805), .ZN(n8082) );
  INV_X1 U10374 ( .A(n12763), .ZN(n11134) );
  NAND2_X1 U10375 ( .A1(n10031), .A2(n10030), .ZN(n13188) );
  OR2_X1 U10376 ( .A1(n9522), .A2(n9521), .ZN(n9523) );
  NAND2_X1 U10377 ( .A1(n8918), .A2(n8917), .ZN(n11101) );
  NAND2_X1 U10378 ( .A1(n12440), .A2(n12443), .ZN(n11170) );
  NAND2_X1 U10379 ( .A1(n10012), .A2(n9281), .ZN(n9288) );
  BUF_X2 U10380 ( .A(n9465), .Z(n11057) );
  INV_X1 U10381 ( .A(n15150), .ZN(n15407) );
  INV_X1 U10382 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8189) );
  NAND2_X1 U10383 ( .A1(n8582), .A2(n8581), .ZN(n12251) );
  NAND2_X1 U10384 ( .A1(n11100), .A2(n8100), .ZN(n8968) );
  INV_X1 U10385 ( .A(n8121), .ZN(n8124) );
  NAND2_X2 U10386 ( .A1(n15690), .A2(n11567), .ZN(n15676) );
  OR2_X1 U10387 ( .A1(n8889), .A2(n8888), .ZN(n8895) );
  OR2_X1 U10388 ( .A1(n6540), .A2(n15756), .ZN(n8084) );
  AND2_X1 U10389 ( .A1(n12969), .A2(n11743), .ZN(n8085) );
  AND2_X1 U10390 ( .A1(n12513), .A2(n12512), .ZN(n8086) );
  INV_X1 U10391 ( .A(P3_U3897), .ZN(n13577) );
  AND2_X2 U10392 ( .A1(n10048), .A2(n14026), .ZN(P3_U3897) );
  NAND2_X2 U10393 ( .A1(n11093), .A2(n15843), .ZN(n15850) );
  NOR2_X1 U10394 ( .A1(n11580), .A2(n11568), .ZN(n8089) );
  NOR3_X1 U10395 ( .A1(n12827), .A2(n12826), .A3(n12825), .ZN(n8090) );
  OR2_X1 U10396 ( .A1(n12362), .A2(n12237), .ZN(n8091) );
  OR2_X1 U10397 ( .A1(n7919), .A2(n14205), .ZN(n8092) );
  AND2_X1 U10398 ( .A1(n9979), .A2(n14910), .ZN(n8093) );
  INV_X1 U10399 ( .A(n14620), .ZN(n9360) );
  INV_X1 U10400 ( .A(n15214), .ZN(n13062) );
  AND2_X1 U10401 ( .A1(n10841), .A2(n9289), .ZN(n15879) );
  INV_X1 U10402 ( .A(n15879), .ZN(n10017) );
  NAND2_X1 U10403 ( .A1(n8916), .A2(n8915), .ZN(n11797) );
  AND2_X1 U10404 ( .A1(n11691), .A2(n10100), .ZN(n8094) );
  OR2_X1 U10405 ( .A1(n12771), .A2(n12770), .ZN(n8096) );
  AND2_X1 U10406 ( .A1(n15387), .A2(n15388), .ZN(n8098) );
  NAND2_X1 U10407 ( .A1(n13953), .A2(n13419), .ZN(n11523) );
  INV_X1 U10408 ( .A(n11586), .ZN(n15701) );
  AND2_X1 U10409 ( .A1(n11399), .A2(n11745), .ZN(n8100) );
  INV_X1 U10410 ( .A(n13180), .ZN(n12919) );
  OR2_X1 U10411 ( .A1(n12994), .A2(n14734), .ZN(n8101) );
  OR2_X1 U10412 ( .A1(n12994), .A2(n14651), .ZN(n8102) );
  INV_X1 U10413 ( .A(n12641), .ZN(n12208) );
  INV_X1 U10414 ( .A(n12639), .ZN(n11580) );
  OR2_X1 U10415 ( .A1(n8889), .A2(n8828), .ZN(n8104) );
  INV_X1 U10416 ( .A(n12461), .ZN(n12462) );
  AND2_X1 U10417 ( .A1(n12467), .A2(n7700), .ZN(n12468) );
  MUX2_X1 U10418 ( .A(n14231), .B(n14500), .S(n12777), .Z(n12866) );
  NAND2_X1 U10419 ( .A1(n12839), .A2(n12838), .ZN(n12840) );
  NOR2_X1 U10420 ( .A1(n8090), .A2(n12840), .ZN(n12841) );
  AND2_X1 U10421 ( .A1(n12881), .A2(n12880), .ZN(n12882) );
  INV_X1 U10422 ( .A(n12891), .ZN(n12892) );
  INV_X1 U10423 ( .A(n12973), .ZN(n9001) );
  INV_X1 U10424 ( .A(n9118), .ZN(n8753) );
  INV_X1 U10425 ( .A(n13864), .ZN(n8429) );
  INV_X1 U10426 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9391) );
  INV_X1 U10427 ( .A(n13902), .ZN(n8576) );
  OAI21_X1 U10428 ( .B1(n13462), .B2(n13544), .A(n13472), .ZN(n8365) );
  INV_X1 U10429 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8403) );
  INV_X1 U10430 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8821) );
  NOR2_X1 U10431 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), 
        .ZN(n8766) );
  AND2_X1 U10432 ( .A1(n10484), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n10055) );
  INV_X1 U10433 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9026) );
  XNOR2_X1 U10434 ( .A(n14570), .B(n12938), .ZN(n12986) );
  NAND2_X1 U10435 ( .A1(n9279), .A2(n14556), .ZN(n9280) );
  AND2_X1 U10436 ( .A1(n9347), .A2(n11400), .ZN(n9348) );
  OR2_X1 U10437 ( .A1(n14241), .A2(n11326), .ZN(n11550) );
  INV_X1 U10438 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8779) );
  NOR2_X1 U10439 ( .A1(n13045), .A2(n13044), .ZN(n13046) );
  INV_X1 U10440 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n10239) );
  AND2_X1 U10441 ( .A1(n11718), .A2(n10959), .ZN(n11716) );
  INV_X1 U10442 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n10403) );
  NAND2_X1 U10443 ( .A1(n15903), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8678) );
  INV_X1 U10444 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n10245) );
  INV_X1 U10445 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8180) );
  OR2_X1 U10446 ( .A1(n10783), .A2(n8608), .ZN(n8681) );
  AND2_X1 U10447 ( .A1(n8644), .A2(n8091), .ZN(n8645) );
  INV_X1 U10448 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9237) );
  OR2_X1 U10449 ( .A1(n13151), .A2(n14223), .ZN(n13147) );
  INV_X1 U10450 ( .A(n12409), .ZN(n9290) );
  NAND2_X1 U10451 ( .A1(n8787), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8979) );
  OR2_X1 U10452 ( .A1(n9337), .A2(n15867), .ZN(n9338) );
  NAND2_X1 U10453 ( .A1(n15877), .A2(n11110), .ZN(n10842) );
  INV_X1 U10454 ( .A(n9816), .ZN(n9817) );
  OR2_X1 U10455 ( .A1(n9831), .A2(n9830), .ZN(n9832) );
  OR2_X1 U10456 ( .A1(n9594), .A2(n11068), .ZN(n9460) );
  INV_X1 U10457 ( .A(n14830), .ZN(n12498) );
  INV_X1 U10458 ( .A(n10795), .ZN(n10797) );
  AND2_X1 U10459 ( .A1(n10536), .A2(n10535), .ZN(n10549) );
  INV_X1 U10460 ( .A(n13214), .ZN(n12693) );
  OR2_X1 U10461 ( .A1(n11273), .A2(n11272), .ZN(n11592) );
  OR2_X1 U10462 ( .A1(n14024), .A2(n8682), .ZN(n11274) );
  AOI21_X1 U10463 ( .B1(n13818), .B2(n8572), .A(n8458), .ZN(n13836) );
  NAND2_X1 U10464 ( .A1(n11260), .A2(n14026), .ZN(n11271) );
  AND2_X1 U10465 ( .A1(n8681), .A2(n13567), .ZN(n8613) );
  INV_X1 U10466 ( .A(n13890), .ZN(n13475) );
  NAND2_X1 U10467 ( .A1(n10847), .A2(n10846), .ZN(n14196) );
  INV_X1 U10468 ( .A(n14194), .ZN(n14209) );
  INV_X1 U10469 ( .A(n8961), .ZN(n9218) );
  INV_X1 U10470 ( .A(n14192), .ZN(n14202) );
  NAND2_X1 U10471 ( .A1(n15850), .A2(n11097), .ZN(n14563) );
  OR2_X1 U10472 ( .A1(n12761), .A2(n12763), .ZN(n10841) );
  AND2_X1 U10473 ( .A1(n14648), .A2(n9355), .ZN(n9357) );
  INV_X1 U10474 ( .A(n14556), .ZN(n14534) );
  INV_X1 U10475 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n8812) );
  INV_X1 U10476 ( .A(n15635), .ZN(n9524) );
  INV_X1 U10477 ( .A(n11865), .ZN(n9621) );
  INV_X1 U10478 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14886) );
  INV_X1 U10479 ( .A(n14936), .ZN(n14914) );
  AND2_X1 U10480 ( .A1(n12654), .A2(n12628), .ZN(n12629) );
  INV_X1 U10481 ( .A(n9907), .ZN(n9986) );
  INV_X2 U10482 ( .A(n9990), .ZN(n12584) );
  INV_X1 U10483 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n15004) );
  INV_X1 U10484 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10915) );
  OR2_X1 U10485 ( .A1(n11463), .A2(n11464), .ZN(n11461) );
  OR2_X1 U10486 ( .A1(n12619), .A2(n10197), .ZN(n14913) );
  OR2_X1 U10487 ( .A1(n11063), .A2(n11062), .ZN(n15712) );
  AND2_X1 U10488 ( .A1(n15369), .A2(n15370), .ZN(n15371) );
  AND2_X1 U10489 ( .A1(n9957), .A2(n9958), .ZN(n9961) );
  INV_X1 U10490 ( .A(n8748), .ZN(n9092) );
  INV_X1 U10491 ( .A(n13360), .ZN(n13325) );
  INV_X1 U10492 ( .A(n13344), .ZN(n12672) );
  INV_X1 U10493 ( .A(n13748), .ZN(n13720) );
  INV_X1 U10494 ( .A(n13757), .ZN(n13667) );
  INV_X1 U10495 ( .A(n13746), .ZN(n13722) );
  AND2_X1 U10496 ( .A1(P3_U3897), .A2(n14038), .ZN(n13748) );
  NAND2_X1 U10497 ( .A1(n12706), .A2(n12705), .ZN(n12707) );
  NOR2_X1 U10498 ( .A1(n8676), .A2(n15896), .ZN(n11764) );
  AND2_X1 U10499 ( .A1(n11764), .A2(n15944), .ZN(n13880) );
  NAND2_X1 U10500 ( .A1(n8614), .A2(n8613), .ZN(n10039) );
  NOR2_X1 U10501 ( .A1(n12708), .A2(n15957), .ZN(n13933) );
  NAND2_X1 U10502 ( .A1(n8683), .A2(n13389), .ZN(n13960) );
  AND2_X1 U10503 ( .A1(n11128), .A2(n15896), .ZN(n15957) );
  NAND2_X1 U10504 ( .A1(n11128), .A2(n13412), .ZN(n15948) );
  NAND2_X1 U10505 ( .A1(n8595), .A2(n6548), .ZN(n10783) );
  INV_X1 U10506 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8621) );
  INV_X1 U10507 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8227) );
  OAI21_X1 U10508 ( .B1(n9314), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9316) );
  INV_X1 U10509 ( .A(n10807), .ZN(n15830) );
  NAND2_X1 U10510 ( .A1(n10640), .A2(n10635), .ZN(n15806) );
  INV_X1 U10511 ( .A(n15806), .ZN(n15831) );
  INV_X1 U10512 ( .A(n15825), .ZN(n15815) );
  INV_X1 U10513 ( .A(n14330), .ZN(n14567) );
  INV_X1 U10514 ( .A(n14563), .ZN(n14541) );
  INV_X1 U10515 ( .A(n15877), .ZN(n14673) );
  AND2_X1 U10516 ( .A1(n15844), .A2(n11134), .ZN(n15877) );
  AND2_X1 U10517 ( .A1(n11455), .A2(n10628), .ZN(n10833) );
  INV_X1 U10518 ( .A(n15646), .ZN(n14926) );
  INV_X1 U10519 ( .A(n15466), .ZN(n15303) );
  INV_X1 U10520 ( .A(n15742), .ZN(n15757) );
  INV_X1 U10521 ( .A(n14928), .ZN(n15641) );
  OR2_X1 U10522 ( .A1(n9999), .A2(P1_U3086), .ZN(n15517) );
  AND2_X1 U10523 ( .A1(n9951), .A2(n9950), .ZN(n13025) );
  INV_X1 U10524 ( .A(n15661), .ZN(n15108) );
  OR2_X1 U10525 ( .A1(n15654), .A2(n10197), .ZN(n15659) );
  OR2_X1 U10526 ( .A1(n15093), .A2(n15092), .ZN(n15105) );
  INV_X1 U10527 ( .A(n12414), .ZN(n15702) );
  NAND2_X2 U10528 ( .A1(n13035), .A2(n15712), .ZN(n15714) );
  OR2_X1 U10529 ( .A1(n11066), .A2(n9996), .ZN(n15742) );
  INV_X1 U10530 ( .A(n15763), .ZN(n15709) );
  AND2_X1 U10531 ( .A1(n15745), .A2(n15770), .ZN(n15760) );
  NAND2_X1 U10532 ( .A1(n12412), .A2(n12588), .ZN(n15763) );
  AND3_X1 U10533 ( .A1(n11063), .A2(n10799), .A3(n10798), .ZN(n15519) );
  NAND2_X1 U10534 ( .A1(n9961), .A2(n9960), .ZN(n10795) );
  AND2_X1 U10535 ( .A1(n9731), .A2(n9765), .ZN(n15053) );
  AND2_X1 U10536 ( .A1(n10140), .A2(n10139), .ZN(n15894) );
  INV_X1 U10537 ( .A(n13357), .ZN(n13333) );
  INV_X1 U10538 ( .A(n13497), .ZN(n13812) );
  INV_X1 U10539 ( .A(n13865), .ZN(n13578) );
  OR2_X1 U10540 ( .A1(n10138), .A2(n10066), .ZN(n13757) );
  OR2_X1 U10541 ( .A1(n15903), .A2(n15919), .ZN(n13894) );
  INV_X1 U10542 ( .A(n12748), .ZN(n11932) );
  AND2_X1 U10543 ( .A1(n8676), .A2(n15923), .ZN(n15903) );
  OR2_X1 U10544 ( .A1(n15973), .A2(n13933), .ZN(n13945) );
  OR2_X1 U10545 ( .A1(n10039), .A2(n10038), .ZN(n15973) );
  OR2_X1 U10546 ( .A1(n15960), .A2(n13933), .ZN(n14021) );
  INV_X2 U10547 ( .A(n15960), .ZN(n15959) );
  OR2_X1 U10548 ( .A1(n15960), .A2(n15948), .ZN(n14013) );
  NAND2_X1 U10549 ( .A1(n10783), .A2(n14026), .ZN(n10817) );
  INV_X1 U10550 ( .A(SI_24_), .ZN(n11935) );
  INV_X1 U10551 ( .A(SI_18_), .ZN(n10928) );
  INV_X1 U10552 ( .A(SI_13_), .ZN(n10743) );
  INV_X1 U10553 ( .A(n11650), .ZN(n10530) );
  XNOR2_X1 U10554 ( .A(n9316), .B(n9315), .ZN(n11455) );
  INV_X1 U10555 ( .A(n14595), .ZN(n14375) );
  INV_X1 U10556 ( .A(n14600), .ZN(n14403) );
  INV_X1 U10557 ( .A(n12924), .ZN(n14217) );
  NAND2_X1 U10558 ( .A1(n10640), .A2(n10633), .ZN(n15825) );
  INV_X1 U10559 ( .A(n15809), .ZN(n15840) );
  INV_X1 U10560 ( .A(n15850), .ZN(n14499) );
  NAND2_X1 U10561 ( .A1(n15850), .A2(n11094), .ZN(n14546) );
  INV_X1 U10562 ( .A(n15886), .ZN(n15885) );
  NOR2_X1 U10563 ( .A1(n15861), .A2(n15852), .ZN(n15857) );
  NAND2_X1 U10564 ( .A1(n9321), .A2(n9320), .ZN(n15863) );
  INV_X1 U10565 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n12286) );
  INV_X1 U10566 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11111) );
  INV_X1 U10567 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10703) );
  NAND2_X1 U10568 ( .A1(n10002), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15646) );
  INV_X1 U10569 ( .A(n15443), .ZN(n14805) );
  INV_X1 U10570 ( .A(n15447), .ZN(n15252) );
  OR2_X1 U10571 ( .A1(n9998), .A2(n9978), .ZN(n15634) );
  OR2_X1 U10572 ( .A1(n15654), .A2(n10200), .ZN(n15111) );
  OR2_X1 U10573 ( .A1(n15654), .A2(n10191), .ZN(n15661) );
  INV_X1 U10574 ( .A(n15720), .ZN(n15686) );
  OR2_X1 U10575 ( .A1(n6546), .A2(n11301), .ZN(n15374) );
  AND2_X2 U10576 ( .A1(n15519), .A2(n10800), .ZN(n15804) );
  NAND2_X1 U10577 ( .A1(n6630), .A2(n15409), .ZN(n15525) );
  AND4_X1 U10578 ( .A1(n15788), .A2(n15787), .A3(n15786), .A4(n15785), .ZN(
        n15803) );
  INV_X1 U10579 ( .A(n15791), .ZN(n15789) );
  INV_X1 U10580 ( .A(n10047), .ZN(n10228) );
  INV_X1 U10581 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n13003) );
  INV_X1 U10582 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11772) );
  INV_X1 U10583 ( .A(n12622), .ZN(n11065) );
  NAND2_X1 U10584 ( .A1(n10044), .A2(n10043), .ZN(P3_U3487) );
  AND2_X2 U10585 ( .A1(n11455), .A2(n10046), .ZN(P2_U3947) );
  NOR2_X1 U10586 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), 
        .ZN(n8112) );
  NOR2_X1 U10587 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), 
        .ZN(n8111) );
  NOR2_X1 U10588 ( .A1(P3_IR_REG_23__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), 
        .ZN(n8110) );
  NOR2_X1 U10589 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_22__SCAN_IN), 
        .ZN(n8109) );
  XNOR2_X2 U10590 ( .A(n8116), .B(n8115), .ZN(n8121) );
  NAND2_X1 U10591 ( .A1(n8117), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8118) );
  INV_X2 U10592 ( .A(n8261), .ZN(n8529) );
  NAND2_X1 U10593 ( .A1(n8199), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8127) );
  NAND2_X4 U10594 ( .A1(n8121), .A2(n14036), .ZN(n13376) );
  INV_X1 U10595 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n8123) );
  OR2_X1 U10596 ( .A1(n13376), .A2(n8123), .ZN(n8126) );
  NAND2_X4 U10597 ( .A1(n8124), .A2(n14036), .ZN(n13377) );
  INV_X1 U10598 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11240) );
  OR2_X1 U10599 ( .A1(n13377), .A2(n11240), .ZN(n8125) );
  CLKBUF_X3 U10600 ( .A(n8706), .Z(n10481) );
  NAND2_X1 U10601 ( .A1(n8129), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8130) );
  MUX2_X1 U10602 ( .A(n9474), .B(n8130), .S(n8908), .Z(n8131) );
  NAND2_X1 U10603 ( .A1(n10481), .A2(SI_0_), .ZN(n8909) );
  NAND2_X1 U10604 ( .A1(n8131), .A2(n8909), .ZN(n14042) );
  XNOR2_X2 U10605 ( .A(n8133), .B(n8132), .ZN(n14038) );
  INV_X1 U10606 ( .A(n11277), .ZN(n11211) );
  INV_X2 U10607 ( .A(n8261), .ZN(n8572) );
  NAND2_X1 U10608 ( .A1(n8572), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8141) );
  NAND2_X1 U10609 ( .A1(n8199), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8140) );
  INV_X1 U10610 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n11280) );
  INV_X1 U10611 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n8137) );
  INV_X1 U10612 ( .A(SI_1_), .ZN(n10518) );
  INV_X1 U10613 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n8142) );
  NAND2_X1 U10614 ( .A1(n8143), .A2(n8144), .ZN(n8145) );
  AND2_X1 U10615 ( .A1(n8145), .A2(n8153), .ZN(n10519) );
  NAND2_X1 U10616 ( .A1(n15904), .A2(n13411), .ZN(n11600) );
  NAND2_X1 U10617 ( .A1(n11600), .A2(n13415), .ZN(n13950) );
  NAND2_X1 U10618 ( .A1(n8199), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8149) );
  INV_X1 U10619 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10092) );
  OR2_X1 U10620 ( .A1(n13377), .A2(n10092), .ZN(n8148) );
  INV_X1 U10621 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n8146) );
  OR2_X1 U10622 ( .A1(n13376), .A2(n8146), .ZN(n8147) );
  NAND2_X1 U10623 ( .A1(n8151), .A2(n6931), .ZN(n8253) );
  INV_X1 U10624 ( .A(n11391), .ZN(n10093) );
  XNOR2_X1 U10625 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8160) );
  XNOR2_X1 U10626 ( .A(n8161), .B(n8160), .ZN(n10515) );
  NAND2_X1 U10627 ( .A1(n13950), .A2(n13951), .ZN(n13953) );
  INV_X1 U10628 ( .A(n13591), .ZN(n15915) );
  NAND2_X1 U10629 ( .A1(n15915), .A2(n8154), .ZN(n13419) );
  INV_X1 U10630 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n11531) );
  NAND2_X1 U10631 ( .A1(n8199), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8158) );
  INV_X1 U10632 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11529) );
  OR2_X1 U10633 ( .A1(n13377), .A2(n11529), .ZN(n8157) );
  INV_X1 U10634 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n8155) );
  OR2_X1 U10635 ( .A1(n13376), .A2(n8155), .ZN(n8156) );
  INV_X1 U10636 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10494) );
  NAND2_X1 U10637 ( .A1(n10494), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8162) );
  XNOR2_X1 U10638 ( .A(n8173), .B(n8172), .ZN(n10520) );
  OR2_X1 U10639 ( .A1(n13372), .A2(n10520), .ZN(n8165) );
  OR2_X1 U10640 ( .A1(n8176), .A2(SI_3_), .ZN(n8164) );
  NAND2_X1 U10641 ( .A1(n8418), .A2(n10523), .ZN(n8163) );
  NAND2_X1 U10642 ( .A1(n13955), .A2(n13243), .ZN(n13420) );
  INV_X1 U10643 ( .A(n13243), .ZN(n11530) );
  NAND2_X1 U10644 ( .A1(n13590), .A2(n11530), .ZN(n13427) );
  NAND2_X1 U10645 ( .A1(n13420), .A2(n13427), .ZN(n13531) );
  INV_X1 U10646 ( .A(n13531), .ZN(n11524) );
  INV_X1 U10647 ( .A(n13420), .ZN(n13426) );
  AND2_X1 U10648 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8166) );
  OR2_X1 U10649 ( .A1(n8166), .A2(n8181), .ZN(n12083) );
  NAND2_X1 U10650 ( .A1(n8572), .A2(n12083), .ZN(n8171) );
  NAND2_X1 U10651 ( .A1(n8199), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8170) );
  INV_X1 U10652 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11506) );
  OR2_X1 U10653 ( .A1(n13377), .A2(n11506), .ZN(n8169) );
  INV_X1 U10654 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n8167) );
  OR2_X1 U10655 ( .A1(n13376), .A2(n8167), .ZN(n8168) );
  INV_X1 U10656 ( .A(n13589), .ZN(n11855) );
  NAND2_X1 U10657 ( .A1(n8173), .A2(n8172), .ZN(n8175) );
  NAND2_X1 U10658 ( .A1(n10213), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8174) );
  XNOR2_X1 U10659 ( .A(n8193), .B(n8192), .ZN(n10524) );
  OR2_X1 U10660 ( .A1(n13372), .A2(n10524), .ZN(n8178) );
  OR2_X1 U10661 ( .A1(n8176), .A2(SI_4_), .ZN(n8177) );
  NAND2_X1 U10662 ( .A1(n11855), .A2(n11811), .ZN(n13428) );
  NAND2_X1 U10663 ( .A1(n13589), .A2(n12081), .ZN(n13425) );
  NAND2_X1 U10664 ( .A1(n13428), .A2(n13425), .ZN(n11501) );
  INV_X1 U10665 ( .A(n13428), .ZN(n8179) );
  OR2_X1 U10666 ( .A1(n8181), .A2(n8180), .ZN(n8182) );
  NAND2_X1 U10667 ( .A1(n8197), .A2(n8182), .ZN(n11854) );
  NAND2_X1 U10668 ( .A1(n8529), .A2(n11854), .ZN(n8187) );
  NAND2_X1 U10669 ( .A1(n8199), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8186) );
  INV_X1 U10670 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n8183) );
  OR2_X1 U10671 ( .A1(n13376), .A2(n8183), .ZN(n8185) );
  INV_X1 U10672 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11632) );
  OR2_X1 U10673 ( .A1(n13377), .A2(n11632), .ZN(n8184) );
  INV_X1 U10674 ( .A(n8188), .ZN(n8190) );
  NAND2_X1 U10675 ( .A1(n8190), .A2(n8189), .ZN(n8205) );
  NAND2_X1 U10676 ( .A1(n8205), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8191) );
  XNOR2_X1 U10677 ( .A(n8191), .B(P3_IR_REG_5__SCAN_IN), .ZN(n11650) );
  OR2_X1 U10678 ( .A1(n8176), .A2(SI_5_), .ZN(n8196) );
  NAND2_X1 U10679 ( .A1(n10498), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8194) );
  XNOR2_X1 U10680 ( .A(n8208), .B(n8207), .ZN(n10527) );
  OR2_X1 U10681 ( .A1(n13372), .A2(n10527), .ZN(n8195) );
  OAI211_X1 U10682 ( .C1(n11650), .C2(n10063), .A(n8196), .B(n8195), .ZN(
        n11495) );
  INV_X1 U10683 ( .A(n11495), .ZN(n11858) );
  NAND2_X1 U10684 ( .A1(n11820), .A2(n11858), .ZN(n13430) );
  NAND2_X1 U10685 ( .A1(n13588), .A2(n11495), .ZN(n13433) );
  NAND2_X1 U10686 ( .A1(n13430), .A2(n13433), .ZN(n13432) );
  NAND2_X1 U10687 ( .A1(n8197), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8198) );
  NAND2_X1 U10688 ( .A1(n8216), .A2(n8198), .ZN(n11804) );
  NAND2_X1 U10689 ( .A1(n8529), .A2(n11804), .ZN(n8204) );
  NAND2_X1 U10690 ( .A1(n8199), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8203) );
  INV_X1 U10691 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n8200) );
  OR2_X1 U10692 ( .A1(n13376), .A2(n8200), .ZN(n8202) );
  INV_X1 U10693 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11519) );
  OR2_X1 U10694 ( .A1(n13377), .A2(n11519), .ZN(n8201) );
  NAND4_X1 U10695 ( .A1(n8204), .A2(n8203), .A3(n8202), .A4(n8201), .ZN(n13587) );
  NAND2_X1 U10696 ( .A1(n8226), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8206) );
  XNOR2_X1 U10697 ( .A(n8206), .B(n8227), .ZN(n10484) );
  NAND2_X1 U10698 ( .A1(n8209), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8210) );
  XNOR2_X1 U10699 ( .A(n10493), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8212) );
  XNOR2_X1 U10700 ( .A(n8225), .B(n8212), .ZN(n10483) );
  OR2_X1 U10701 ( .A1(n13372), .A2(n10483), .ZN(n8214) );
  INV_X1 U10702 ( .A(SI_6_), .ZN(n10482) );
  OR2_X1 U10703 ( .A1(n8176), .A2(n10482), .ZN(n8213) );
  OAI211_X1 U10704 ( .C1(n10063), .C2(n10484), .A(n8214), .B(n8213), .ZN(
        n15943) );
  NAND2_X1 U10705 ( .A1(n11880), .A2(n15943), .ZN(n8215) );
  INV_X1 U10706 ( .A(n15943), .ZN(n11817) );
  NAND2_X1 U10707 ( .A1(n13587), .A2(n11817), .ZN(n13435) );
  NAND2_X1 U10708 ( .A1(n8215), .A2(n13435), .ZN(n13536) );
  INV_X1 U10709 ( .A(n13536), .ZN(n11509) );
  INV_X1 U10710 ( .A(n8215), .ZN(n13438) );
  NAND2_X1 U10711 ( .A1(n8199), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8222) );
  AND2_X1 U10712 ( .A1(n8216), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8217) );
  OR2_X1 U10713 ( .A1(n8217), .A2(n8241), .ZN(n11885) );
  NAND2_X1 U10714 ( .A1(n8529), .A2(n11885), .ZN(n8221) );
  INV_X1 U10715 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11887) );
  OR2_X1 U10716 ( .A1(n13377), .A2(n11887), .ZN(n8220) );
  INV_X1 U10717 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n8218) );
  OR2_X1 U10718 ( .A1(n13376), .A2(n8218), .ZN(n8219) );
  NAND4_X1 U10719 ( .A1(n8222), .A2(n8221), .A3(n8220), .A4(n8219), .ZN(n13586) );
  NAND2_X1 U10720 ( .A1(n7345), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8223) );
  XNOR2_X1 U10721 ( .A(n8235), .B(n8234), .ZN(n10501) );
  NAND2_X1 U10722 ( .A1(n10501), .A2(n13369), .ZN(n8232) );
  INV_X2 U10723 ( .A(n8176), .ZN(n8568) );
  INV_X1 U10724 ( .A(SI_7_), .ZN(n10502) );
  INV_X1 U10725 ( .A(n8226), .ZN(n8228) );
  NAND2_X1 U10726 ( .A1(n8228), .A2(n8227), .ZN(n8236) );
  NAND2_X1 U10727 ( .A1(n8236), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8230) );
  INV_X1 U10728 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8229) );
  XNOR2_X1 U10729 ( .A(n8230), .B(n8229), .ZN(n11145) );
  NAND2_X1 U10730 ( .A1(n11840), .A2(n11829), .ZN(n13440) );
  NOR2_X1 U10731 ( .A1(n11876), .A2(n13437), .ZN(n11875) );
  INV_X1 U10732 ( .A(n13440), .ZN(n8233) );
  XNOR2_X1 U10733 ( .A(n8249), .B(n6747), .ZN(n10506) );
  NAND2_X1 U10734 ( .A1(n10506), .A2(n13369), .ZN(n8239) );
  OAI21_X1 U10735 ( .B1(n8236), .B2(P3_IR_REG_7__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8237) );
  XNOR2_X1 U10736 ( .A(n8237), .B(P3_IR_REG_8__SCAN_IN), .ZN(n10115) );
  AOI22_X1 U10737 ( .A1(n8568), .A2(SI_8_), .B1(n10115), .B2(n8418), .ZN(n8238) );
  NOR2_X1 U10738 ( .A1(n8241), .A2(n8240), .ZN(n8242) );
  OR2_X1 U10739 ( .A1(n8263), .A2(n8242), .ZN(n12180) );
  NAND2_X1 U10740 ( .A1(n8572), .A2(n12180), .ZN(n8247) );
  NAND2_X1 U10741 ( .A1(n8199), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8246) );
  INV_X1 U10742 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11763) );
  OR2_X1 U10743 ( .A1(n13377), .A2(n11763), .ZN(n8245) );
  INV_X1 U10744 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n8243) );
  OR2_X1 U10745 ( .A1(n13376), .A2(n8243), .ZN(n8244) );
  NAND4_X1 U10746 ( .A1(n8247), .A2(n8246), .A3(n8245), .A4(n8244), .ZN(n13585) );
  NAND2_X1 U10747 ( .A1(n12178), .A2(n13585), .ZN(n13443) );
  INV_X1 U10748 ( .A(n12178), .ZN(n8248) );
  NAND2_X1 U10749 ( .A1(n10490), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8250) );
  XNOR2_X1 U10750 ( .A(n8272), .B(n8271), .ZN(n10499) );
  NAND2_X1 U10751 ( .A1(n10499), .A2(n13369), .ZN(n8260) );
  INV_X1 U10752 ( .A(SI_9_), .ZN(n10500) );
  INV_X1 U10753 ( .A(n8251), .ZN(n8252) );
  NOR2_X1 U10754 ( .A1(n6634), .A2(n8252), .ZN(n8255) );
  INV_X1 U10755 ( .A(n8253), .ZN(n8254) );
  NAND2_X1 U10756 ( .A1(n8255), .A2(n8254), .ZN(n8257) );
  NAND2_X1 U10757 ( .A1(n8257), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8256) );
  MUX2_X1 U10758 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8256), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n8258) );
  NAND2_X1 U10759 ( .A1(n8258), .A2(n8274), .ZN(n11317) );
  AOI22_X1 U10760 ( .A1(n8568), .A2(n10500), .B1(n8418), .B2(n11317), .ZN(
        n8259) );
  NAND2_X1 U10761 ( .A1(n8260), .A2(n8259), .ZN(n12156) );
  OR2_X1 U10762 ( .A1(n8263), .A2(n8262), .ZN(n8264) );
  NAND2_X1 U10763 ( .A1(n8280), .A2(n8264), .ZN(n11929) );
  NAND2_X1 U10764 ( .A1(n8529), .A2(n11929), .ZN(n8269) );
  NAND2_X1 U10765 ( .A1(n8199), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8268) );
  INV_X1 U10766 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n8265) );
  OR2_X1 U10767 ( .A1(n13376), .A2(n8265), .ZN(n8267) );
  INV_X1 U10768 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11928) );
  OR2_X1 U10769 ( .A1(n13377), .A2(n11928), .ZN(n8266) );
  NAND4_X1 U10770 ( .A1(n8269), .A2(n8268), .A3(n8267), .A4(n8266), .ZN(n13584) );
  NAND2_X1 U10771 ( .A1(n12156), .A2(n13584), .ZN(n13447) );
  OR2_X1 U10772 ( .A1(n12156), .A2(n13584), .ZN(n13448) );
  INV_X1 U10773 ( .A(n13448), .ZN(n8270) );
  NAND2_X1 U10774 ( .A1(n10514), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8273) );
  XNOR2_X1 U10775 ( .A(n8288), .B(n8287), .ZN(n10503) );
  NAND2_X1 U10776 ( .A1(n10503), .A2(n13369), .ZN(n8279) );
  INV_X1 U10777 ( .A(SI_10_), .ZN(n10504) );
  NAND2_X1 U10778 ( .A1(n8274), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8275) );
  MUX2_X1 U10779 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8275), .S(
        P3_IR_REG_10__SCAN_IN), .Z(n8277) );
  NAND2_X1 U10780 ( .A1(n8277), .A2(n8387), .ZN(n10505) );
  AOI22_X1 U10781 ( .A1(n8568), .A2(n10504), .B1(n8418), .B2(n10505), .ZN(
        n8278) );
  NAND2_X1 U10782 ( .A1(n8279), .A2(n8278), .ZN(n12119) );
  NAND2_X1 U10783 ( .A1(n8280), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8281) );
  NAND2_X1 U10784 ( .A1(n8293), .A2(n8281), .ZN(n12108) );
  NAND2_X1 U10785 ( .A1(n8529), .A2(n12108), .ZN(n8286) );
  NAND2_X1 U10786 ( .A1(n8199), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8285) );
  INV_X1 U10787 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n12110) );
  OR2_X1 U10788 ( .A1(n13377), .A2(n12110), .ZN(n8284) );
  INV_X1 U10789 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n8282) );
  OR2_X1 U10790 ( .A1(n13376), .A2(n8282), .ZN(n8283) );
  NAND4_X1 U10791 ( .A1(n8286), .A2(n8285), .A3(n8284), .A4(n8283), .ZN(n13583) );
  NAND2_X1 U10792 ( .A1(n12119), .A2(n13583), .ZN(n13455) );
  OR2_X1 U10793 ( .A1(n12119), .A2(n13583), .ZN(n13406) );
  XNOR2_X1 U10794 ( .A(n8301), .B(n8300), .ZN(n10531) );
  NAND2_X1 U10795 ( .A1(n10531), .A2(n13369), .ZN(n8292) );
  NAND2_X1 U10796 ( .A1(n8387), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8290) );
  XNOR2_X1 U10797 ( .A(n8290), .B(n8304), .ZN(n11964) );
  AOI22_X1 U10798 ( .A1(n8568), .A2(n10449), .B1(n8418), .B2(n11964), .ZN(
        n8291) );
  NAND2_X1 U10799 ( .A1(n8292), .A2(n8291), .ZN(n13949) );
  NAND2_X1 U10800 ( .A1(n8293), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8294) );
  NAND2_X1 U10801 ( .A1(n8309), .A2(n8294), .ZN(n12307) );
  NAND2_X1 U10802 ( .A1(n8572), .A2(n12307), .ZN(n8299) );
  NAND2_X1 U10803 ( .A1(n8199), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8298) );
  INV_X1 U10804 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n8295) );
  OR2_X1 U10805 ( .A1(n13376), .A2(n8295), .ZN(n8297) );
  INV_X1 U10806 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n12053) );
  OR2_X1 U10807 ( .A1(n13377), .A2(n12053), .ZN(n8296) );
  NAND4_X1 U10808 ( .A1(n8299), .A2(n8298), .A3(n8297), .A4(n8296), .ZN(n13582) );
  NAND2_X1 U10809 ( .A1(n13949), .A2(n13582), .ZN(n13454) );
  NAND2_X1 U10810 ( .A1(n8301), .A2(n8300), .ZN(n8303) );
  NAND2_X1 U10811 ( .A1(n8726), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8302) );
  XNOR2_X1 U10812 ( .A(n10707), .B(P2_DATAO_REG_12__SCAN_IN), .ZN(n8316) );
  XNOR2_X1 U10813 ( .A(n8318), .B(n8316), .ZN(n10615) );
  NAND2_X1 U10814 ( .A1(n10615), .A2(n13369), .ZN(n8308) );
  INV_X1 U10815 ( .A(n8387), .ZN(n8305) );
  NAND2_X1 U10816 ( .A1(n8305), .A2(n8304), .ZN(n8320) );
  NAND2_X1 U10817 ( .A1(n8320), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8306) );
  XNOR2_X1 U10818 ( .A(n8306), .B(P3_IR_REG_12__SCAN_IN), .ZN(n13614) );
  AOI22_X1 U10819 ( .A1(n8568), .A2(SI_12_), .B1(n8418), .B2(n13614), .ZN(
        n8307) );
  NAND2_X1 U10820 ( .A1(n8308), .A2(n8307), .ZN(n12264) );
  NAND2_X1 U10821 ( .A1(n8199), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8314) );
  AND2_X1 U10822 ( .A1(n8309), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8310) );
  OR2_X1 U10823 ( .A1(n8310), .A2(n8326), .ZN(n12359) );
  NAND2_X1 U10824 ( .A1(n8572), .A2(n12359), .ZN(n8313) );
  INV_X1 U10825 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12105) );
  OR2_X1 U10826 ( .A1(n13377), .A2(n12105), .ZN(n8312) );
  INV_X1 U10827 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n12095) );
  OR2_X1 U10828 ( .A1(n13376), .A2(n12095), .ZN(n8311) );
  NAND4_X1 U10829 ( .A1(n8314), .A2(n8313), .A3(n8312), .A4(n8311), .ZN(n13581) );
  OR2_X1 U10830 ( .A1(n12264), .A2(n12237), .ZN(n13457) );
  NAND2_X1 U10831 ( .A1(n12264), .A2(n12237), .ZN(n8315) );
  NAND2_X1 U10832 ( .A1(n13457), .A2(n8315), .ZN(n13542) );
  INV_X1 U10833 ( .A(n13542), .ZN(n12088) );
  INV_X1 U10834 ( .A(n8315), .ZN(n13458) );
  INV_X1 U10835 ( .A(n8316), .ZN(n8317) );
  NAND2_X1 U10836 ( .A1(n8722), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8319) );
  XNOR2_X1 U10837 ( .A(n8348), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8347) );
  XNOR2_X1 U10838 ( .A(n8347), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n10742) );
  NAND2_X1 U10839 ( .A1(n10742), .A2(n13369), .ZN(n8325) );
  INV_X1 U10840 ( .A(n8320), .ZN(n8322) );
  INV_X1 U10841 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8321) );
  NAND2_X1 U10842 ( .A1(n8322), .A2(n8321), .ZN(n8338) );
  NAND2_X1 U10843 ( .A1(n8338), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8323) );
  XNOR2_X1 U10844 ( .A(n8323), .B(n10272), .ZN(n10744) );
  AOI22_X1 U10845 ( .A1(n8568), .A2(n10743), .B1(n8418), .B2(n10744), .ZN(
        n8324) );
  OR2_X1 U10846 ( .A1(n8326), .A2(n10403), .ZN(n8327) );
  NAND2_X1 U10847 ( .A1(n8360), .A2(n8327), .ZN(n12255) );
  NAND2_X1 U10848 ( .A1(n8572), .A2(n12255), .ZN(n8332) );
  NAND2_X1 U10849 ( .A1(n8199), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8331) );
  INV_X1 U10850 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n13627) );
  OR2_X1 U10851 ( .A1(n13377), .A2(n13627), .ZN(n8330) );
  INV_X1 U10852 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n8328) );
  OR2_X1 U10853 ( .A1(n13376), .A2(n8328), .ZN(n8329) );
  NAND2_X1 U10854 ( .A1(n10785), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8335) );
  NAND2_X1 U10855 ( .A1(n10703), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n8333) );
  AND2_X1 U10856 ( .A1(n8335), .A2(n8333), .ZN(n8334) );
  NOR2_X1 U10857 ( .A1(n10703), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n8336) );
  AOI22_X1 U10858 ( .A1(n8336), .A2(n8335), .B1(P1_DATAO_REG_14__SCAN_IN), 
        .B2(n10787), .ZN(n8337) );
  XNOR2_X1 U10859 ( .A(n10755), .B(P2_DATAO_REG_15__SCAN_IN), .ZN(n8367) );
  XNOR2_X1 U10860 ( .A(n8369), .B(n8367), .ZN(n10752) );
  NAND2_X1 U10861 ( .A1(n10752), .A2(n13369), .ZN(n8342) );
  INV_X1 U10862 ( .A(n8353), .ZN(n8339) );
  INV_X1 U10863 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8354) );
  NAND2_X1 U10864 ( .A1(n8339), .A2(n8354), .ZN(n8372) );
  NAND2_X1 U10865 ( .A1(n8372), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8340) );
  XNOR2_X1 U10866 ( .A(n8340), .B(P3_IR_REG_15__SCAN_IN), .ZN(n13678) );
  AOI22_X1 U10867 ( .A1(n13678), .A2(n8418), .B1(n8568), .B2(SI_15_), .ZN(
        n8341) );
  AND2_X1 U10868 ( .A1(n6599), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8343) );
  OR2_X1 U10869 ( .A1(n8343), .A2(n8377), .ZN(n13355) );
  NAND2_X1 U10870 ( .A1(n13355), .A2(n8529), .ZN(n8346) );
  AOI22_X1 U10871 ( .A1(n8667), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n8199), .B2(
        P3_REG1_REG_15__SCAN_IN), .ZN(n8345) );
  NAND2_X1 U10872 ( .A1(n8668), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8344) );
  OR2_X1 U10873 ( .A1(n13356), .A2(n13344), .ZN(n13466) );
  NAND2_X1 U10874 ( .A1(n13356), .A2(n13344), .ZN(n13472) );
  NAND2_X1 U10875 ( .A1(n13466), .A2(n13472), .ZN(n13544) );
  INV_X1 U10876 ( .A(n13544), .ZN(n13469) );
  NAND2_X1 U10877 ( .A1(n8347), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8350) );
  INV_X1 U10878 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10705) );
  NAND2_X1 U10879 ( .A1(n8348), .A2(n10705), .ZN(n8349) );
  NAND2_X1 U10880 ( .A1(n8350), .A2(n8349), .ZN(n8352) );
  XNOR2_X1 U10881 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8351) );
  XNOR2_X1 U10882 ( .A(n8352), .B(n8351), .ZN(n10780) );
  NAND2_X1 U10883 ( .A1(n10780), .A2(n13369), .ZN(n8357) );
  INV_X1 U10884 ( .A(SI_14_), .ZN(n10781) );
  NAND2_X1 U10885 ( .A1(n8353), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8355) );
  XNOR2_X1 U10886 ( .A(n8355), .B(n8354), .ZN(n10782) );
  AOI22_X1 U10887 ( .A1(n8568), .A2(n10781), .B1(n8418), .B2(n10782), .ZN(
        n8356) );
  INV_X1 U10888 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n8364) );
  NAND2_X1 U10889 ( .A1(n8668), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8359) );
  NAND2_X1 U10890 ( .A1(n8667), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8358) );
  AND2_X1 U10891 ( .A1(n8359), .A2(n8358), .ZN(n8363) );
  NAND2_X1 U10892 ( .A1(n8360), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8361) );
  NAND2_X1 U10893 ( .A1(n6599), .A2(n8361), .ZN(n12366) );
  NAND2_X1 U10894 ( .A1(n12366), .A2(n8529), .ZN(n8362) );
  OAI211_X1 U10895 ( .C1(n8442), .C2(n8364), .A(n8363), .B(n8362), .ZN(n13579)
         );
  NAND2_X1 U10896 ( .A1(n13465), .A2(n13579), .ZN(n8649) );
  NAND2_X1 U10897 ( .A1(n12245), .A2(n13580), .ZN(n13460) );
  INV_X1 U10898 ( .A(n8365), .ZN(n8366) );
  INV_X1 U10899 ( .A(n12383), .ZN(n8381) );
  INV_X1 U10900 ( .A(n8367), .ZN(n8368) );
  NAND2_X1 U10901 ( .A1(n8369), .A2(n8368), .ZN(n8371) );
  NAND2_X1 U10902 ( .A1(n10757), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8370) );
  XNOR2_X1 U10903 ( .A(n10711), .B(P2_DATAO_REG_16__SCAN_IN), .ZN(n8382) );
  NAND2_X1 U10904 ( .A1(n10822), .A2(n13369), .ZN(n8375) );
  OAI21_X1 U10905 ( .B1(n8372), .B2(P3_IR_REG_15__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8373) );
  XNOR2_X1 U10906 ( .A(n8373), .B(P3_IR_REG_16__SCAN_IN), .ZN(n13693) );
  AOI22_X1 U10907 ( .A1(n13693), .A2(n8418), .B1(SI_16_), .B2(n8568), .ZN(
        n8374) );
  INV_X1 U10908 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13671) );
  NOR2_X1 U10909 ( .A1(n8377), .A2(n8376), .ZN(n8378) );
  OR2_X1 U10910 ( .A1(n8391), .A2(n8378), .ZN(n13295) );
  NAND2_X1 U10911 ( .A1(n13295), .A2(n8572), .ZN(n8380) );
  AOI22_X1 U10912 ( .A1(n8667), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n8668), .B2(
        P3_REG0_REG_16__SCAN_IN), .ZN(n8379) );
  XNOR2_X1 U10913 ( .A(n13476), .B(n13475), .ZN(n12386) );
  NAND2_X1 U10914 ( .A1(n13476), .A2(n13475), .ZN(n13474) );
  INV_X1 U10915 ( .A(n8382), .ZN(n8383) );
  NAND2_X1 U10916 ( .A1(n10760), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8385) );
  NAND2_X1 U10917 ( .A1(n8400), .A2(n8385), .ZN(n8398) );
  XNOR2_X1 U10918 ( .A(n8399), .B(n8398), .ZN(n10870) );
  NAND2_X1 U10919 ( .A1(n10870), .A2(n13369), .ZN(n8390) );
  NAND2_X1 U10920 ( .A1(n6761), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8388) );
  XNOR2_X1 U10921 ( .A(n8388), .B(P3_IR_REG_17__SCAN_IN), .ZN(n13700) );
  AOI22_X1 U10922 ( .A1(n8568), .A2(SI_17_), .B1(n8418), .B2(n13700), .ZN(
        n8389) );
  OR2_X1 U10923 ( .A1(n8391), .A2(n10245), .ZN(n8392) );
  NAND2_X1 U10924 ( .A1(n8421), .A2(n8392), .ZN(n13879) );
  NAND2_X1 U10925 ( .A1(n13879), .A2(n8529), .ZN(n8397) );
  INV_X1 U10926 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13891) );
  NAND2_X1 U10927 ( .A1(n8199), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8394) );
  NAND2_X1 U10928 ( .A1(n8668), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8393) );
  OAI211_X1 U10929 ( .C1(n13377), .C2(n13891), .A(n8394), .B(n8393), .ZN(n8395) );
  INV_X1 U10930 ( .A(n8395), .ZN(n8396) );
  OR2_X1 U10931 ( .A1(n14017), .A2(n13865), .ZN(n13402) );
  NAND2_X1 U10932 ( .A1(n14017), .A2(n13865), .ZN(n13478) );
  XNOR2_X1 U10933 ( .A(n10891), .B(P2_DATAO_REG_18__SCAN_IN), .ZN(n8413) );
  INV_X1 U10934 ( .A(n8413), .ZN(n8401) );
  NAND2_X1 U10935 ( .A1(n10890), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8402) );
  XNOR2_X1 U10936 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .ZN(n8432) );
  XNOR2_X1 U10937 ( .A(n8433), .B(n8432), .ZN(n10930) );
  NAND2_X1 U10938 ( .A1(n10930), .A2(n13369), .ZN(n8406) );
  NAND2_X1 U10939 ( .A1(n6613), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8404) );
  AOI22_X1 U10940 ( .A1(n8568), .A2(n10929), .B1(n8418), .B2(n13745), .ZN(
        n8405) );
  INV_X1 U10941 ( .A(n13853), .ZN(n14003) );
  AND2_X1 U10942 ( .A1(n8423), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8407) );
  OR2_X1 U10943 ( .A1(n8407), .A2(n8438), .ZN(n13850) );
  NAND2_X1 U10944 ( .A1(n13850), .A2(n8572), .ZN(n8412) );
  INV_X1 U10945 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n14007) );
  NAND2_X1 U10946 ( .A1(n8199), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8409) );
  NAND2_X1 U10947 ( .A1(n8667), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8408) );
  OAI211_X1 U10948 ( .C1(n13376), .C2(n14007), .A(n8409), .B(n8408), .ZN(n8410) );
  INV_X1 U10949 ( .A(n8410), .ZN(n8411) );
  NAND2_X1 U10950 ( .A1(n14003), .A2(n13864), .ZN(n13483) );
  XNOR2_X1 U10951 ( .A(n8414), .B(n8413), .ZN(n10926) );
  NAND2_X1 U10952 ( .A1(n10926), .A2(n13369), .ZN(n8420) );
  NAND2_X1 U10953 ( .A1(n8415), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8416) );
  MUX2_X1 U10954 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8416), .S(
        P3_IR_REG_18__SCAN_IN), .Z(n8417) );
  AND2_X1 U10955 ( .A1(n8417), .A2(n6613), .ZN(n13725) );
  AOI22_X1 U10956 ( .A1(n8568), .A2(SI_18_), .B1(n8418), .B2(n13725), .ZN(
        n8419) );
  NAND2_X1 U10957 ( .A1(n8421), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8422) );
  NAND2_X1 U10958 ( .A1(n8423), .A2(n8422), .ZN(n13866) );
  NAND2_X1 U10959 ( .A1(n13866), .A2(n8529), .ZN(n8428) );
  INV_X1 U10960 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13868) );
  NAND2_X1 U10961 ( .A1(n8668), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8425) );
  NAND2_X1 U10962 ( .A1(n8199), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8424) );
  OAI211_X1 U10963 ( .C1(n13377), .C2(n13868), .A(n8425), .B(n8424), .ZN(n8426) );
  INV_X1 U10964 ( .A(n8426), .ZN(n8427) );
  NAND2_X1 U10965 ( .A1(n13874), .A2(n13848), .ZN(n13480) );
  INV_X1 U10966 ( .A(n13843), .ZN(n13404) );
  OAI21_X1 U10967 ( .B1(n13404), .B2(n8429), .A(n13853), .ZN(n8431) );
  NAND2_X1 U10968 ( .A1(n13404), .A2(n8429), .ZN(n8430) );
  INV_X1 U10969 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10984) );
  NAND2_X1 U10970 ( .A1(n10984), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8434) );
  XNOR2_X1 U10971 ( .A(n8461), .B(P1_DATAO_REG_20__SCAN_IN), .ZN(n8447) );
  XNOR2_X1 U10972 ( .A(n8447), .B(n10931), .ZN(n11212) );
  NAND2_X1 U10973 ( .A1(n11212), .A2(n13369), .ZN(n8436) );
  INV_X1 U10974 ( .A(SI_20_), .ZN(n11214) );
  OR2_X1 U10975 ( .A1(n8176), .A2(n11214), .ZN(n8435) );
  NOR2_X1 U10976 ( .A1(n8438), .A2(n8437), .ZN(n8439) );
  OR2_X1 U10977 ( .A1(n8454), .A2(n8439), .ZN(n13830) );
  NAND2_X1 U10978 ( .A1(n13830), .A2(n8529), .ZN(n8445) );
  INV_X1 U10979 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n10291) );
  NAND2_X1 U10980 ( .A1(n8668), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8441) );
  NAND2_X1 U10981 ( .A1(n8667), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8440) );
  OAI211_X1 U10982 ( .C1(n10291), .C2(n8442), .A(n8441), .B(n8440), .ZN(n8443)
         );
  INV_X1 U10983 ( .A(n8443), .ZN(n8444) );
  NAND2_X1 U10984 ( .A1(n13831), .A2(n13849), .ZN(n13488) );
  NAND2_X1 U10985 ( .A1(n13829), .A2(n13832), .ZN(n8446) );
  NAND2_X1 U10986 ( .A1(n8446), .A2(n13487), .ZN(n13817) );
  NAND2_X1 U10987 ( .A1(n8461), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8448) );
  NAND2_X1 U10988 ( .A1(n8449), .A2(n8448), .ZN(n8451) );
  XNOR2_X1 U10989 ( .A(n11111), .B(P2_DATAO_REG_21__SCAN_IN), .ZN(n8450) );
  XNOR2_X1 U10990 ( .A(n8451), .B(n8450), .ZN(n11452) );
  NAND2_X1 U10991 ( .A1(n11452), .A2(n13369), .ZN(n8453) );
  OR2_X1 U10992 ( .A1(n8176), .A2(n11453), .ZN(n8452) );
  OR2_X1 U10993 ( .A1(n8454), .A2(n13274), .ZN(n8455) );
  NAND2_X1 U10994 ( .A1(n8469), .A2(n8455), .ZN(n13818) );
  INV_X1 U10995 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n13820) );
  NAND2_X1 U10996 ( .A1(n8668), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8457) );
  NAND2_X1 U10997 ( .A1(n8199), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8456) );
  OAI211_X1 U10998 ( .C1(n13377), .C2(n13820), .A(n8457), .B(n8456), .ZN(n8458) );
  NAND2_X1 U10999 ( .A1(n13923), .A2(n13836), .ZN(n13492) );
  NAND2_X1 U11000 ( .A1(n13817), .A2(n13492), .ZN(n8459) );
  NAND2_X1 U11001 ( .A1(n8459), .A2(n13491), .ZN(n13808) );
  AOI22_X1 U11002 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n12407), .B1(n11111), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8460) );
  NAND2_X1 U11003 ( .A1(n10931), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8462) );
  NAND2_X1 U11004 ( .A1(n8462), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8464) );
  NOR2_X1 U11005 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8463) );
  AOI22_X1 U11006 ( .A1(n8464), .A2(P1_DATAO_REG_21__SCAN_IN), .B1(n8463), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8465) );
  NAND2_X1 U11007 ( .A1(n11132), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8479) );
  NAND2_X1 U11008 ( .A1(n8761), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8466) );
  NAND2_X1 U11009 ( .A1(n8479), .A2(n8466), .ZN(n8477) );
  XNOR2_X1 U11010 ( .A(n8478), .B(n8477), .ZN(n11130) );
  NAND2_X1 U11011 ( .A1(n11130), .A2(n13369), .ZN(n8468) );
  OR2_X1 U11012 ( .A1(n8176), .A2(n8763), .ZN(n8467) );
  NAND2_X1 U11013 ( .A1(n8469), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8470) );
  NAND2_X1 U11014 ( .A1(n6652), .A2(n8470), .ZN(n13809) );
  NAND2_X1 U11015 ( .A1(n13809), .A2(n8529), .ZN(n8475) );
  INV_X1 U11016 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n13814) );
  NAND2_X1 U11017 ( .A1(n8668), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8472) );
  NAND2_X1 U11018 ( .A1(n8199), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8471) );
  OAI211_X1 U11019 ( .C1(n13377), .C2(n13814), .A(n8472), .B(n8471), .ZN(n8473) );
  INV_X1 U11020 ( .A(n8473), .ZN(n8474) );
  NAND2_X1 U11021 ( .A1(n13990), .A2(n13826), .ZN(n13494) );
  NAND2_X1 U11022 ( .A1(n13808), .A2(n13494), .ZN(n8476) );
  INV_X1 U11023 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11457) );
  NAND2_X1 U11024 ( .A1(n11457), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8494) );
  INV_X1 U11025 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11460) );
  NAND2_X1 U11026 ( .A1(n11460), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8480) );
  OR2_X1 U11027 ( .A1(n8482), .A2(n8481), .ZN(n8483) );
  NAND2_X1 U11028 ( .A1(n8495), .A2(n8483), .ZN(n11412) );
  NAND2_X1 U11029 ( .A1(n11412), .A2(n13369), .ZN(n8485) );
  OR2_X1 U11030 ( .A1(n8176), .A2(n11414), .ZN(n8484) );
  NAND2_X1 U11031 ( .A1(n6652), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8486) );
  NAND2_X1 U11032 ( .A1(n8486), .A2(n8498), .ZN(n13801) );
  NAND2_X1 U11033 ( .A1(n13801), .A2(n8572), .ZN(n8491) );
  INV_X1 U11034 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13983) );
  NAND2_X1 U11035 ( .A1(n8667), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8488) );
  NAND2_X1 U11036 ( .A1(n8199), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8487) );
  OAI211_X1 U11037 ( .C1(n13983), .C2(n13376), .A(n8488), .B(n8487), .ZN(n8489) );
  INV_X1 U11038 ( .A(n8489), .ZN(n8490) );
  NAND2_X1 U11039 ( .A1(n13984), .A2(n13497), .ZN(n8492) );
  NAND2_X1 U11040 ( .A1(n13500), .A2(n8492), .ZN(n13551) );
  INV_X1 U11041 ( .A(n13500), .ZN(n8493) );
  XNOR2_X1 U11042 ( .A(n8504), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n11934) );
  NAND2_X1 U11043 ( .A1(n11934), .A2(n13369), .ZN(n8497) );
  OR2_X1 U11044 ( .A1(n8176), .A2(n11935), .ZN(n8496) );
  NAND2_X1 U11045 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(n8498), .ZN(n8499) );
  INV_X1 U11046 ( .A(n8511), .ZN(n8513) );
  INV_X1 U11047 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n8500) );
  OR2_X1 U11048 ( .A1(n13376), .A2(n8500), .ZN(n8503) );
  INV_X1 U11049 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n8501) );
  OR2_X1 U11050 ( .A1(n13377), .A2(n8501), .ZN(n8502) );
  NAND2_X1 U11051 ( .A1(n13912), .A2(n13776), .ZN(n13499) );
  INV_X1 U11052 ( .A(n13788), .ZN(n13793) );
  NAND2_X1 U11053 ( .A1(n8504), .A2(n11772), .ZN(n8507) );
  INV_X1 U11054 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12103) );
  XNOR2_X1 U11055 ( .A(n12103), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8508) );
  XNOR2_X1 U11056 ( .A(n8523), .B(n8508), .ZN(n12120) );
  NAND2_X1 U11057 ( .A1(n12120), .A2(n13369), .ZN(n8510) );
  NAND2_X1 U11058 ( .A1(n8568), .A2(SI_25_), .ZN(n8509) );
  NAND2_X1 U11059 ( .A1(n8199), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8520) );
  INV_X1 U11060 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8512) );
  NAND2_X1 U11061 ( .A1(n8512), .A2(n8511), .ZN(n8527) );
  NAND2_X1 U11062 ( .A1(P3_REG3_REG_25__SCAN_IN), .A2(n8513), .ZN(n8514) );
  NAND2_X1 U11063 ( .A1(n8527), .A2(n8514), .ZN(n13782) );
  NAND2_X1 U11064 ( .A1(n8572), .A2(n13782), .ZN(n8519) );
  INV_X1 U11065 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n8515) );
  OR2_X1 U11066 ( .A1(n13377), .A2(n8515), .ZN(n8518) );
  INV_X1 U11067 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n8516) );
  OR2_X1 U11068 ( .A1(n13376), .A2(n8516), .ZN(n8517) );
  OR2_X1 U11069 ( .A1(n13908), .A2(n13338), .ZN(n13506) );
  NAND2_X1 U11070 ( .A1(n13908), .A2(n13338), .ZN(n13505) );
  NOR2_X1 U11071 ( .A1(n12103), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8522) );
  NAND2_X1 U11072 ( .A1(n12103), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8521) );
  XNOR2_X1 U11073 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .ZN(n8524) );
  XNOR2_X1 U11074 ( .A(n8535), .B(n8524), .ZN(n12248) );
  NAND2_X1 U11075 ( .A1(n12248), .A2(n13369), .ZN(n8526) );
  INV_X1 U11076 ( .A(SI_26_), .ZN(n12249) );
  OR2_X1 U11077 ( .A1(n8176), .A2(n12249), .ZN(n8525) );
  NAND2_X1 U11078 ( .A1(n8527), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8528) );
  NAND2_X1 U11079 ( .A1(n8539), .A2(n8528), .ZN(n13770) );
  NAND2_X1 U11080 ( .A1(n8529), .A2(n13770), .ZN(n8533) );
  NAND2_X1 U11081 ( .A1(n8199), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8532) );
  INV_X1 U11082 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13976) );
  OR2_X1 U11083 ( .A1(n13376), .A2(n13976), .ZN(n8531) );
  INV_X1 U11084 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n13769) );
  OR2_X1 U11085 ( .A1(n13377), .A2(n13769), .ZN(n8530) );
  NAND4_X1 U11086 ( .A1(n8533), .A2(n8532), .A3(n8531), .A4(n8530), .ZN(n13576) );
  NAND2_X1 U11087 ( .A1(n13977), .A2(n13775), .ZN(n13510) );
  AND2_X1 U11088 ( .A1(n12221), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8534) );
  XNOR2_X1 U11089 ( .A(n9237), .B(P2_DATAO_REG_27__SCAN_IN), .ZN(n8536) );
  XNOR2_X1 U11090 ( .A(n8548), .B(n8536), .ZN(n12310) );
  NAND2_X1 U11091 ( .A1(n12310), .A2(n13369), .ZN(n8538) );
  INV_X1 U11092 ( .A(SI_27_), .ZN(n12311) );
  OR2_X1 U11093 ( .A1(n8176), .A2(n12311), .ZN(n8537) );
  NAND2_X1 U11094 ( .A1(n8539), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8540) );
  NAND2_X1 U11095 ( .A1(n8529), .A2(n13225), .ZN(n8546) );
  NAND2_X1 U11096 ( .A1(n8199), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8545) );
  INV_X1 U11097 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n8541) );
  OR2_X1 U11098 ( .A1(n13377), .A2(n8541), .ZN(n8544) );
  INV_X1 U11099 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n8542) );
  OR2_X1 U11100 ( .A1(n13376), .A2(n8542), .ZN(n8543) );
  OR2_X1 U11101 ( .A1(n13229), .A2(n10028), .ZN(n13515) );
  NAND2_X1 U11102 ( .A1(n13229), .A2(n10028), .ZN(n13522) );
  NAND2_X1 U11103 ( .A1(n12700), .A2(n13530), .ZN(n8547) );
  XNOR2_X1 U11104 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .ZN(n8549) );
  XNOR2_X1 U11105 ( .A(n8563), .B(n8549), .ZN(n14037) );
  NAND2_X1 U11106 ( .A1(n14037), .A2(n13369), .ZN(n8551) );
  NAND2_X1 U11107 ( .A1(n8568), .A2(SI_28_), .ZN(n8550) );
  NAND2_X1 U11108 ( .A1(n8199), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8561) );
  INV_X1 U11109 ( .A(n8554), .ZN(n8553) );
  INV_X1 U11110 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n8552) );
  NAND2_X1 U11111 ( .A1(n8553), .A2(n8552), .ZN(n8677) );
  NAND2_X1 U11112 ( .A1(n8554), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8555) );
  NAND2_X1 U11113 ( .A1(n8677), .A2(n8555), .ZN(n13264) );
  NAND2_X1 U11114 ( .A1(n8572), .A2(n13264), .ZN(n8560) );
  INV_X1 U11115 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n8556) );
  OR2_X1 U11116 ( .A1(n13377), .A2(n8556), .ZN(n8559) );
  INV_X1 U11117 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n8557) );
  OR2_X1 U11118 ( .A1(n13376), .A2(n8557), .ZN(n8558) );
  NAND4_X1 U11119 ( .A1(n8561), .A2(n8560), .A3(n8559), .A4(n8558), .ZN(n13575) );
  NAND2_X1 U11120 ( .A1(n13269), .A2(n12703), .ZN(n13523) );
  AND2_X1 U11121 ( .A1(n12286), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8562) );
  INV_X1 U11122 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n13185) );
  NAND2_X1 U11123 ( .A1(n13185), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8564) );
  XNOR2_X1 U11124 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n8565) );
  NAND2_X1 U11125 ( .A1(n8566), .A2(n8565), .ZN(n13005) );
  NAND2_X1 U11126 ( .A1(n13005), .A2(n8567), .ZN(n14035) );
  OR2_X1 U11127 ( .A1(n14035), .A2(n13372), .ZN(n8570) );
  NAND2_X1 U11128 ( .A1(n8568), .A2(SI_29_), .ZN(n8569) );
  INV_X1 U11129 ( .A(n8677), .ZN(n8571) );
  NAND2_X1 U11130 ( .A1(n8572), .A2(n8571), .ZN(n13381) );
  NAND2_X1 U11131 ( .A1(n8667), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8575) );
  NAND2_X1 U11132 ( .A1(n8199), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8574) );
  NAND2_X1 U11133 ( .A1(n8668), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8573) );
  NAND4_X1 U11134 ( .A1(n13381), .A2(n8575), .A3(n8574), .A4(n8573), .ZN(
        n13574) );
  NAND2_X1 U11135 ( .A1(n8576), .A2(n13574), .ZN(n13517) );
  INV_X1 U11136 ( .A(n13574), .ZN(n13267) );
  NAND2_X1 U11137 ( .A1(n13902), .A2(n13267), .ZN(n13520) );
  NAND2_X1 U11138 ( .A1(n13517), .A2(n13520), .ZN(n13555) );
  INV_X1 U11139 ( .A(n13555), .ZN(n8577) );
  NAND2_X1 U11140 ( .A1(n8584), .A2(n8579), .ZN(n8587) );
  NAND2_X1 U11141 ( .A1(n8587), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8580) );
  MUX2_X1 U11142 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8580), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n8581) );
  INV_X1 U11143 ( .A(n8584), .ZN(n8585) );
  NAND2_X1 U11144 ( .A1(n8585), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8586) );
  MUX2_X1 U11145 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8586), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8588) );
  INV_X1 U11146 ( .A(n12123), .ZN(n8589) );
  OAI21_X1 U11147 ( .B1(P3_B_REG_SCAN_IN), .B2(n8589), .A(n6548), .ZN(n8590)
         );
  NAND2_X1 U11148 ( .A1(n8592), .A2(n8590), .ZN(n8591) );
  INV_X1 U11149 ( .A(P3_B_REG_SCAN_IN), .ZN(n8593) );
  XNOR2_X1 U11150 ( .A(n8592), .B(n8593), .ZN(n8594) );
  NAND2_X1 U11151 ( .A1(n8594), .A2(n12123), .ZN(n8595) );
  NAND2_X1 U11152 ( .A1(n12251), .A2(n12123), .ZN(n8596) );
  XNOR2_X1 U11153 ( .A(n14027), .B(n14024), .ZN(n8614) );
  NOR2_X1 U11154 ( .A1(P3_D_REG_8__SCAN_IN), .A2(P3_D_REG_25__SCAN_IN), .ZN(
        n8601) );
  NOR4_X1 U11155 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_2__SCAN_IN), .A3(
        P3_D_REG_11__SCAN_IN), .A4(P3_D_REG_17__SCAN_IN), .ZN(n8600) );
  NOR4_X1 U11156 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_10__SCAN_IN), .ZN(n8599) );
  NOR4_X1 U11157 ( .A1(P3_D_REG_22__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n8598) );
  NAND4_X1 U11158 ( .A1(n8601), .A2(n8600), .A3(n8599), .A4(n8598), .ZN(n8607)
         );
  NOR4_X1 U11159 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n8605) );
  NOR4_X1 U11160 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P3_D_REG_31__SCAN_IN), .A3(
        P3_D_REG_14__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n8604) );
  NOR4_X1 U11161 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8603) );
  NOR4_X1 U11162 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n8602) );
  NAND4_X1 U11163 ( .A1(n8605), .A2(n8604), .A3(n8603), .A4(n8602), .ZN(n8606)
         );
  NOR2_X1 U11164 ( .A1(n8607), .A2(n8606), .ZN(n8608) );
  NOR2_X1 U11165 ( .A1(n12251), .A2(n12123), .ZN(n8609) );
  NAND2_X1 U11166 ( .A1(n8610), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8612) );
  NAND2_X1 U11167 ( .A1(n8615), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8616) );
  INV_X1 U11168 ( .A(n8617), .ZN(n8618) );
  AND2_X1 U11169 ( .A1(n8630), .A2(n13514), .ZN(n8624) );
  MUX2_X1 U11170 ( .A(n13529), .B(n8630), .S(n13514), .Z(n10032) );
  NAND2_X1 U11171 ( .A1(n14024), .A2(n10032), .ZN(n8623) );
  OAI21_X1 U11172 ( .B1(n14024), .B2(n8624), .A(n8623), .ZN(n8625) );
  AND2_X1 U11173 ( .A1(n13412), .A2(n11213), .ZN(n8626) );
  XNOR2_X1 U11174 ( .A(n11128), .B(n8626), .ZN(n8628) );
  NAND2_X1 U11175 ( .A1(n13412), .A2(n13745), .ZN(n8627) );
  NAND2_X1 U11176 ( .A1(n8628), .A2(n8627), .ZN(n11262) );
  INV_X1 U11177 ( .A(n13529), .ZN(n13565) );
  AND2_X1 U11178 ( .A1(n15948), .A2(n13565), .ZN(n8629) );
  NAND2_X1 U11179 ( .A1(n11262), .A2(n8629), .ZN(n8631) );
  AND2_X1 U11180 ( .A1(n8665), .A2(n15896), .ZN(n11490) );
  NOR2_X1 U11181 ( .A1(n12708), .A2(n11490), .ZN(n15919) );
  NAND2_X1 U11182 ( .A1(n13495), .A2(n13494), .ZN(n13550) );
  INV_X1 U11183 ( .A(n13923), .ZN(n13279) );
  NAND2_X1 U11184 ( .A1(n15906), .A2(n11277), .ZN(n11604) );
  NAND2_X1 U11185 ( .A1(n11594), .A2(n11604), .ZN(n15907) );
  NAND2_X1 U11186 ( .A1(n13954), .A2(n15905), .ZN(n8632) );
  NAND2_X1 U11187 ( .A1(n15915), .A2(n13965), .ZN(n11525) );
  AND2_X1 U11188 ( .A1(n13531), .A2(n11525), .ZN(n8633) );
  NAND2_X1 U11189 ( .A1(n13589), .A2(n11811), .ZN(n8634) );
  NAND2_X1 U11190 ( .A1(n13587), .A2(n15943), .ZN(n11877) );
  NAND2_X1 U11191 ( .A1(n13432), .A2(n11877), .ZN(n8637) );
  NAND2_X1 U11192 ( .A1(n11820), .A2(n11495), .ZN(n11511) );
  NAND2_X1 U11193 ( .A1(n13536), .A2(n11511), .ZN(n11513) );
  AOI21_X1 U11194 ( .B1(n11513), .B2(n11877), .A(n13539), .ZN(n8636) );
  NAND2_X1 U11195 ( .A1(n13586), .A2(n11829), .ZN(n8638) );
  INV_X1 U11196 ( .A(n13584), .ZN(n12034) );
  NOR2_X1 U11197 ( .A1(n12156), .A2(n12034), .ZN(n11890) );
  NAND2_X1 U11198 ( .A1(n13406), .A2(n13455), .ZN(n13541) );
  NAND2_X1 U11199 ( .A1(n13448), .A2(n13447), .ZN(n11920) );
  NAND2_X1 U11200 ( .A1(n12178), .A2(n11925), .ZN(n11921) );
  NAND2_X1 U11201 ( .A1(n11920), .A2(n11921), .ZN(n11889) );
  INV_X1 U11202 ( .A(n11890), .ZN(n8639) );
  NAND2_X1 U11203 ( .A1(n11889), .A2(n8639), .ZN(n8640) );
  AND2_X1 U11204 ( .A1(n13541), .A2(n8640), .ZN(n8641) );
  INV_X1 U11205 ( .A(n13583), .ZN(n12304) );
  OR2_X1 U11206 ( .A1(n12119), .A2(n12304), .ZN(n8642) );
  INV_X1 U11207 ( .A(n13582), .ZN(n12357) );
  NAND2_X1 U11208 ( .A1(n13949), .A2(n12357), .ZN(n12087) );
  NAND3_X1 U11209 ( .A1(n12049), .A2(n13542), .A3(n12087), .ZN(n8646) );
  NAND3_X1 U11210 ( .A1(n13542), .A2(n13453), .A3(n12087), .ZN(n8644) );
  INV_X1 U11211 ( .A(n12264), .ZN(n12362) );
  NOR2_X1 U11212 ( .A1(n12245), .A2(n12332), .ZN(n8648) );
  NAND2_X1 U11213 ( .A1(n12245), .A2(n12332), .ZN(n8647) );
  INV_X1 U11214 ( .A(n13579), .ZN(n13351) );
  OR2_X1 U11215 ( .A1(n13465), .A2(n13351), .ZN(n8650) );
  AND2_X1 U11216 ( .A1(n13544), .A2(n8652), .ZN(n13881) );
  AND2_X1 U11217 ( .A1(n13881), .A2(n13877), .ZN(n8651) );
  INV_X1 U11218 ( .A(n13877), .ZN(n8656) );
  INV_X1 U11219 ( .A(n8652), .ZN(n8653) );
  NAND2_X1 U11220 ( .A1(n13356), .A2(n12672), .ZN(n12384) );
  NAND2_X1 U11221 ( .A1(n13476), .A2(n13890), .ZN(n8654) );
  AND2_X1 U11222 ( .A1(n8655), .A2(n8654), .ZN(n13883) );
  NAND2_X1 U11223 ( .A1(n14017), .A2(n13578), .ZN(n8657) );
  INV_X1 U11224 ( .A(n13869), .ZN(n8659) );
  OR2_X1 U11225 ( .A1(n13874), .A2(n13887), .ZN(n8661) );
  OR2_X1 U11226 ( .A1(n13853), .A2(n13864), .ZN(n8662) );
  NAND2_X2 U11227 ( .A1(n13509), .A2(n13510), .ZN(n13766) );
  XNOR2_X1 U11228 ( .A(n8664), .B(n13555), .ZN(n8675) );
  NAND2_X1 U11229 ( .A1(n13570), .A2(n13735), .ZN(n8683) );
  NAND2_X1 U11230 ( .A1(n8665), .A2(n11596), .ZN(n13389) );
  INV_X1 U11231 ( .A(n14038), .ZN(n13566) );
  INV_X1 U11232 ( .A(n7288), .ZN(n13736) );
  NAND2_X1 U11233 ( .A1(n13566), .A2(n13736), .ZN(n10066) );
  AND2_X1 U11234 ( .A1(n10063), .A2(n10066), .ZN(n8672) );
  AND2_X1 U11235 ( .A1(n13566), .A2(P3_B_REG_SCAN_IN), .ZN(n8666) );
  OR2_X1 U11236 ( .A1(n15916), .A2(n8666), .ZN(n13759) );
  NAND2_X1 U11237 ( .A1(n8667), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8671) );
  NAND2_X1 U11238 ( .A1(n8668), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8670) );
  NAND2_X1 U11239 ( .A1(n8199), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8669) );
  INV_X1 U11240 ( .A(n8672), .ZN(n8673) );
  OAI22_X1 U11241 ( .A1(n13759), .A2(n13385), .B1(n12703), .B2(n15914), .ZN(
        n8674) );
  INV_X1 U11242 ( .A(n15948), .ZN(n15944) );
  NOR2_X1 U11243 ( .A1(n15923), .A2(n8677), .ZN(n13760) );
  AOI21_X1 U11244 ( .B1(n13902), .B2(n13880), .A(n13760), .ZN(n8679) );
  INV_X1 U11245 ( .A(n14027), .ZN(n8680) );
  NAND3_X1 U11246 ( .A1(n14024), .A2(n8680), .A3(n8681), .ZN(n11273) );
  INV_X1 U11247 ( .A(n11262), .ZN(n8684) );
  NAND2_X1 U11248 ( .A1(n8681), .A2(n14027), .ZN(n8682) );
  NAND2_X1 U11249 ( .A1(n13412), .A2(n11596), .ZN(n11595) );
  OR2_X1 U11250 ( .A1(n8683), .A2(n11595), .ZN(n11257) );
  OAI22_X1 U11251 ( .A1(n11273), .A2(n8684), .B1(n11274), .B2(n11257), .ZN(
        n8685) );
  NAND2_X1 U11252 ( .A1(n8685), .A2(n13567), .ZN(n8689) );
  INV_X1 U11253 ( .A(n11274), .ZN(n8687) );
  OR2_X1 U11254 ( .A1(n13514), .A2(n13529), .ZN(n8686) );
  NOR2_X1 U11255 ( .A1(n11271), .A2(n8686), .ZN(n11267) );
  NAND2_X1 U11256 ( .A1(n8687), .A2(n11267), .ZN(n8688) );
  OR2_X1 U11257 ( .A1(n13901), .A2(n14021), .ZN(n8691) );
  NAND2_X1 U11258 ( .A1(n13902), .A2(n14018), .ZN(n8690) );
  INV_X1 U11259 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n10412) );
  MUX2_X1 U11260 ( .A(n11113), .B(n11111), .S(n10481), .Z(n8759) );
  NAND2_X1 U11261 ( .A1(n8759), .A2(n11453), .ZN(n9153) );
  INV_X1 U11262 ( .A(SI_0_), .ZN(n9473) );
  INV_X1 U11263 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10487) );
  AOI21_X1 U11264 ( .B1(n8706), .B2(P1_DATAO_REG_1__SCAN_IN), .A(SI_1_), .ZN(
        n8692) );
  OAI21_X1 U11265 ( .B1(n8706), .B2(n10487), .A(n8692), .ZN(n8693) );
  INV_X1 U11266 ( .A(n8693), .ZN(n8694) );
  NAND2_X1 U11267 ( .A1(n8706), .A2(n10595), .ZN(n8695) );
  MUX2_X1 U11268 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n8706), .Z(n8838) );
  NAND2_X1 U11269 ( .A1(n8838), .A2(SI_3_), .ZN(n8882) );
  NAND2_X1 U11270 ( .A1(n8697), .A2(SI_2_), .ZN(n8836) );
  AND2_X1 U11271 ( .A1(n8882), .A2(n8836), .ZN(n8698) );
  XNOR2_X1 U11272 ( .A(n8702), .B(SI_4_), .ZN(n8884) );
  NOR2_X1 U11273 ( .A1(n8838), .A2(SI_3_), .ZN(n8699) );
  NAND2_X1 U11274 ( .A1(n8702), .A2(SI_4_), .ZN(n8863) );
  NAND2_X1 U11275 ( .A1(n8705), .A2(SI_5_), .ZN(n8704) );
  AND2_X1 U11276 ( .A1(n8863), .A2(n8704), .ZN(n8703) );
  XNOR2_X1 U11277 ( .A(n8709), .B(SI_6_), .ZN(n8921) );
  INV_X1 U11278 ( .A(n8921), .ZN(n8707) );
  NAND2_X1 U11279 ( .A1(n8710), .A2(SI_7_), .ZN(n8711) );
  MUX2_X1 U11280 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n10481), .Z(n8714) );
  XNOR2_X1 U11281 ( .A(n8714), .B(SI_8_), .ZN(n8955) );
  INV_X1 U11282 ( .A(n8955), .ZN(n8713) );
  NAND2_X1 U11283 ( .A1(n8714), .A2(SI_8_), .ZN(n8715) );
  MUX2_X1 U11284 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n10481), .Z(n8717) );
  XNOR2_X1 U11285 ( .A(n8717), .B(SI_9_), .ZN(n8972) );
  INV_X1 U11286 ( .A(n8972), .ZN(n8716) );
  NAND2_X1 U11287 ( .A1(n8717), .A2(SI_9_), .ZN(n8718) );
  MUX2_X1 U11288 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n8706), .Z(n8986) );
  INV_X1 U11289 ( .A(n8986), .ZN(n8720) );
  NAND2_X1 U11290 ( .A1(n8720), .A2(n10504), .ZN(n8721) );
  NAND2_X1 U11291 ( .A1(n8723), .A2(n10617), .ZN(n8738) );
  INV_X1 U11292 ( .A(n8723), .ZN(n8724) );
  NAND2_X1 U11293 ( .A1(n8724), .A2(SI_12_), .ZN(n8725) );
  NAND2_X1 U11294 ( .A1(n8738), .A2(n8725), .ZN(n8730) );
  NAND2_X1 U11295 ( .A1(n8986), .A2(SI_10_), .ZN(n9002) );
  MUX2_X1 U11296 ( .A(n8726), .B(n10620), .S(n10481), .Z(n8731) );
  INV_X1 U11297 ( .A(n8731), .ZN(n8727) );
  NAND2_X1 U11298 ( .A1(n8727), .A2(SI_11_), .ZN(n9003) );
  NAND2_X1 U11299 ( .A1(n9002), .A2(n9003), .ZN(n8728) );
  NOR2_X1 U11300 ( .A1(n8730), .A2(n8728), .ZN(n8729) );
  INV_X1 U11301 ( .A(n8730), .ZN(n9034) );
  NAND2_X1 U11302 ( .A1(n8731), .A2(n10449), .ZN(n9032) );
  INV_X1 U11303 ( .A(n9032), .ZN(n8732) );
  NAND2_X1 U11304 ( .A1(n9034), .A2(n8732), .ZN(n8733) );
  NAND2_X1 U11305 ( .A1(n8734), .A2(n10754), .ZN(n8742) );
  INV_X1 U11306 ( .A(n8734), .ZN(n8735) );
  INV_X1 U11307 ( .A(n9074), .ZN(n8737) );
  MUX2_X1 U11308 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n9260), .Z(n9076) );
  NAND2_X1 U11309 ( .A1(n9076), .A2(SI_14_), .ZN(n8736) );
  MUX2_X1 U11310 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n10481), .Z(n8739) );
  NAND2_X1 U11311 ( .A1(n8739), .A2(SI_13_), .ZN(n9079) );
  INV_X1 U11312 ( .A(n8738), .ZN(n9055) );
  NAND2_X1 U11313 ( .A1(n9055), .A2(n9079), .ZN(n8741) );
  INV_X1 U11314 ( .A(n8739), .ZN(n8740) );
  NAND2_X1 U11315 ( .A1(n8740), .A2(n10743), .ZN(n9060) );
  OAI211_X1 U11316 ( .C1(n9076), .C2(SI_14_), .A(n8741), .B(n9060), .ZN(n9078)
         );
  INV_X1 U11317 ( .A(n8742), .ZN(n8743) );
  MUX2_X1 U11318 ( .A(n10709), .B(n10711), .S(n9260), .Z(n8745) );
  NAND2_X1 U11319 ( .A1(n8745), .A2(n10824), .ZN(n8749) );
  INV_X1 U11320 ( .A(n8745), .ZN(n8746) );
  NAND2_X1 U11321 ( .A1(n8746), .A2(SI_16_), .ZN(n8747) );
  NAND2_X1 U11322 ( .A1(n8749), .A2(n8747), .ZN(n8748) );
  MUX2_X1 U11323 ( .A(n10759), .B(n10760), .S(n9260), .Z(n9105) );
  INV_X1 U11324 ( .A(n9105), .ZN(n8750) );
  NAND2_X1 U11325 ( .A1(n8750), .A2(SI_17_), .ZN(n8751) );
  NAND2_X1 U11326 ( .A1(n9105), .A2(n10871), .ZN(n8752) );
  MUX2_X1 U11327 ( .A(n10890), .B(n10891), .S(n9260), .Z(n9118) );
  MUX2_X1 U11328 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n10481), .Z(n8756) );
  XNOR2_X1 U11329 ( .A(n8756), .B(SI_19_), .ZN(n8809) );
  INV_X1 U11330 ( .A(n8809), .ZN(n8755) );
  NAND2_X1 U11331 ( .A1(n8753), .A2(SI_18_), .ZN(n8754) );
  INV_X1 U11332 ( .A(n8756), .ZN(n8757) );
  MUX2_X1 U11333 ( .A(n10931), .B(n12407), .S(n10481), .Z(n9138) );
  INV_X1 U11334 ( .A(n9138), .ZN(n8758) );
  INV_X1 U11335 ( .A(n8759), .ZN(n8760) );
  NAND2_X1 U11336 ( .A1(n8760), .A2(SI_21_), .ZN(n9152) );
  MUX2_X1 U11337 ( .A(n8761), .B(n11132), .S(n10481), .Z(n9167) );
  MUX2_X1 U11338 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9260), .Z(n9181) );
  INV_X1 U11339 ( .A(n9181), .ZN(n8762) );
  OAI22_X1 U11340 ( .A1(n9167), .A2(n8763), .B1(n8762), .B2(n11414), .ZN(n8764) );
  MUX2_X1 U11341 ( .A(n11772), .B(n11770), .S(n10481), .Z(n9202) );
  MUX2_X1 U11342 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n9260), .Z(n9208) );
  XNOR2_X1 U11343 ( .A(n9210), .B(n9209), .ZN(n12098) );
  NOR2_X2 U11344 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .ZN(n9324) );
  AND2_X2 U11345 ( .A1(n9324), .A2(n8766), .ZN(n9274) );
  AND2_X2 U11346 ( .A1(n9274), .A2(n8767), .ZN(n8778) );
  AND3_X2 U11347 ( .A1(n8770), .A2(n8769), .A3(n8768), .ZN(n8813) );
  NOR2_X1 U11348 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n8773) );
  NOR2_X1 U11349 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n8772) );
  INV_X1 U11350 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8780) );
  NAND2_X1 U11351 ( .A1(n12098), .A2(n12734), .ZN(n8784) );
  OR2_X1 U11352 ( .A1(n8902), .A2(n12103), .ZN(n8783) );
  INV_X1 U11353 ( .A(n8948), .ZN(n8786) );
  NAND2_X1 U11354 ( .A1(n8786), .A2(n8785), .ZN(n8962) );
  INV_X1 U11355 ( .A(n8962), .ZN(n8787) );
  OR2_X2 U11356 ( .A1(n8979), .A2(n8978), .ZN(n8994) );
  OR2_X2 U11357 ( .A1(n9044), .A2(n9026), .ZN(n9068) );
  OR2_X2 U11358 ( .A1(n9113), .A2(n9112), .ZN(n9127) );
  INV_X1 U11359 ( .A(n9127), .ZN(n8790) );
  INV_X1 U11360 ( .A(n9172), .ZN(n8791) );
  INV_X1 U11361 ( .A(n9186), .ZN(n8792) );
  INV_X1 U11362 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n14133) );
  OR2_X2 U11363 ( .A1(n9195), .A2(n14133), .ZN(n9216) );
  XNOR2_X1 U11364 ( .A(n9216), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n14343) );
  XNOR2_X2 U11365 ( .A(n8797), .B(n13078), .ZN(n8798) );
  NAND2_X1 U11366 ( .A1(n14343), .A2(n9218), .ZN(n8805) );
  INV_X1 U11367 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8802) );
  NAND2_X1 U11368 ( .A1(n12737), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8801) );
  NAND2_X1 U11369 ( .A1(n8798), .A2(n6985), .ZN(n8891) );
  NAND2_X1 U11370 ( .A1(n9283), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8800) );
  OAI211_X1 U11371 ( .C1(n8802), .C2(n8931), .A(n8801), .B(n8800), .ZN(n8803)
         );
  INV_X1 U11372 ( .A(n8803), .ZN(n8804) );
  NAND2_X1 U11373 ( .A1(n8806), .A2(n10928), .ZN(n8807) );
  NAND2_X1 U11374 ( .A1(n8808), .A2(n8807), .ZN(n9119) );
  NAND2_X1 U11375 ( .A1(n10983), .A2(n12734), .ZN(n8820) );
  INV_X1 U11376 ( .A(n9303), .ZN(n8814) );
  NAND2_X1 U11377 ( .A1(n9272), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8818) );
  AOI22_X1 U11378 ( .A1(n14299), .A2(n9123), .B1(n12733), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n8819) );
  NAND2_X1 U11379 ( .A1(n9129), .A2(n8821), .ZN(n8822) );
  AND2_X1 U11380 ( .A1(n9144), .A2(n8822), .ZN(n14445) );
  NAND2_X1 U11381 ( .A1(n14445), .A2(n9218), .ZN(n8827) );
  INV_X1 U11382 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n14294) );
  NAND2_X1 U11383 ( .A1(n12737), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n8824) );
  NAND2_X1 U11384 ( .A1(n9283), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8823) );
  OAI211_X1 U11385 ( .C1(n14294), .C2(n8931), .A(n8824), .B(n8823), .ZN(n8825)
         );
  INV_X1 U11386 ( .A(n8825), .ZN(n8826) );
  INV_X1 U11387 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n8828) );
  INV_X1 U11388 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n8829) );
  OR2_X1 U11389 ( .A1(n8891), .A2(n8829), .ZN(n8832) );
  OR2_X1 U11390 ( .A1(n8961), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8831) );
  OR2_X1 U11391 ( .A1(n8931), .A2(n14278), .ZN(n8830) );
  NAND2_X1 U11392 ( .A1(n8860), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8835) );
  INV_X1 U11393 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8834) );
  NAND2_X1 U11394 ( .A1(n8837), .A2(n8836), .ZN(n8881) );
  XNOR2_X1 U11395 ( .A(n8838), .B(SI_3_), .ZN(n8879) );
  XNOR2_X1 U11396 ( .A(n8881), .B(n8879), .ZN(n10212) );
  OR2_X1 U11397 ( .A1(n8902), .A2(n10213), .ZN(n8839) );
  NAND2_X1 U11398 ( .A1(n12737), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8844) );
  INV_X1 U11399 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n8840) );
  OR2_X1 U11400 ( .A1(n8891), .A2(n8840), .ZN(n8843) );
  INV_X1 U11401 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n14261) );
  OR2_X1 U11402 ( .A1(n8961), .A2(n14261), .ZN(n8842) );
  INV_X1 U11403 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10645) );
  OR2_X1 U11404 ( .A1(n8931), .A2(n10645), .ZN(n8841) );
  INV_X1 U11405 ( .A(n8847), .ZN(n8897) );
  NAND2_X1 U11406 ( .A1(n8897), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8848) );
  OR2_X1 U11407 ( .A1(n7327), .A2(n14262), .ZN(n8850) );
  OR2_X1 U11408 ( .A1(n8902), .A2(n10494), .ZN(n8849) );
  NAND2_X1 U11409 ( .A1(n14242), .A2(n15867), .ZN(n8851) );
  AND2_X1 U11410 ( .A1(n10977), .A2(n8851), .ZN(n10969) );
  NAND2_X1 U11411 ( .A1(n12737), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8859) );
  INV_X1 U11412 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n8852) );
  OR2_X1 U11413 ( .A1(n8891), .A2(n8852), .ZN(n8858) );
  INV_X1 U11414 ( .A(n8853), .ZN(n8870) );
  INV_X1 U11415 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8854) );
  NAND2_X1 U11416 ( .A1(n8870), .A2(n8854), .ZN(n8855) );
  NAND2_X1 U11417 ( .A1(n8948), .A2(n8855), .ZN(n11233) );
  OR2_X1 U11418 ( .A1(n8961), .A2(n11233), .ZN(n8857) );
  INV_X1 U11419 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10653) );
  OR2_X1 U11420 ( .A1(n8931), .A2(n10653), .ZN(n8856) );
  NAND2_X1 U11421 ( .A1(n8923), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8875) );
  INV_X1 U11422 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8861) );
  NAND2_X1 U11423 ( .A1(n8875), .A2(n8861), .ZN(n8877) );
  NAND2_X1 U11424 ( .A1(n8877), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8862) );
  XNOR2_X1 U11425 ( .A(n8862), .B(P2_IR_REG_5__SCAN_IN), .ZN(n10674) );
  AOI22_X1 U11426 ( .A1(n12733), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9123), 
        .B2(n10674), .ZN(n8867) );
  NAND2_X1 U11427 ( .A1(n8864), .A2(n8863), .ZN(n8866) );
  XNOR2_X1 U11428 ( .A(n8866), .B(n8865), .ZN(n10216) );
  NAND2_X1 U11429 ( .A1(n14239), .A2(n15880), .ZN(n8868) );
  INV_X1 U11430 ( .A(n12963), .ZN(n8913) );
  INV_X1 U11431 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n8869) );
  INV_X1 U11432 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10622) );
  OR2_X1 U11433 ( .A1(n8889), .A2(n10622), .ZN(n8873) );
  OAI21_X1 U11434 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n8870), .ZN(n11559) );
  OR2_X1 U11435 ( .A1(n8961), .A2(n11559), .ZN(n8872) );
  INV_X1 U11436 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10650) );
  OR2_X1 U11437 ( .A1(n8931), .A2(n10650), .ZN(n8871) );
  NAND4_X1 U11438 ( .A1(n8874), .A2(n8873), .A3(n8872), .A4(n8871), .ZN(n14240) );
  INV_X1 U11439 ( .A(n8875), .ZN(n8876) );
  NAND2_X1 U11440 ( .A1(n8876), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n8878) );
  AOI22_X1 U11441 ( .A1(n12733), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n9123), 
        .B2(n10651), .ZN(n8887) );
  INV_X1 U11442 ( .A(n8879), .ZN(n8880) );
  NAND2_X1 U11443 ( .A1(n8881), .A2(n8880), .ZN(n8883) );
  NAND2_X1 U11444 ( .A1(n8883), .A2(n8882), .ZN(n8885) );
  XNOR2_X1 U11445 ( .A(n8885), .B(n8884), .ZN(n10219) );
  NAND2_X1 U11446 ( .A1(n10219), .A2(n12734), .ZN(n8886) );
  NAND2_X1 U11447 ( .A1(n14240), .A2(n15873), .ZN(n8911) );
  INV_X1 U11448 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n8888) );
  INV_X1 U11449 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n8890) );
  OR2_X1 U11450 ( .A1(n8891), .A2(n8890), .ZN(n8894) );
  INV_X1 U11451 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n14248) );
  INV_X1 U11452 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10641) );
  MUX2_X1 U11453 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8896), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8898) );
  XNOR2_X1 U11454 ( .A(n8899), .B(SI_1_), .ZN(n8901) );
  MUX2_X1 U11455 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n8706), .Z(n8900) );
  XNOR2_X1 U11456 ( .A(n8900), .B(n8901), .ZN(n10594) );
  INV_X1 U11457 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10746) );
  OR2_X1 U11458 ( .A1(n8889), .A2(n10746), .ZN(n8907) );
  INV_X1 U11459 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n15842) );
  OR2_X1 U11460 ( .A1(n8961), .A2(n15842), .ZN(n8906) );
  INV_X1 U11461 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10747) );
  OR2_X1 U11462 ( .A1(n8931), .A2(n10747), .ZN(n8905) );
  INV_X1 U11463 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n14252) );
  XNOR2_X1 U11464 ( .A(n8909), .B(n8908), .ZN(n14741) );
  MUX2_X1 U11465 ( .A(n14252), .B(n14741), .S(n10626), .Z(n12770) );
  NOR2_X1 U11466 ( .A1(n14243), .A2(n12770), .ZN(n11154) );
  NAND2_X1 U11467 ( .A1(n12961), .A2(n11154), .ZN(n11153) );
  INV_X1 U11468 ( .A(n6553), .ZN(n12009) );
  OR2_X1 U11469 ( .A1(n12775), .A2(n12009), .ZN(n10967) );
  OR2_X1 U11470 ( .A1(n14242), .A2(n15867), .ZN(n10968) );
  NAND2_X1 U11471 ( .A1(n11153), .A2(n8910), .ZN(n10970) );
  NAND4_X1 U11472 ( .A1(n10969), .A2(n8913), .A3(n8911), .A4(n10970), .ZN(
        n8916) );
  INV_X1 U11473 ( .A(n8911), .ZN(n8912) );
  OAI21_X1 U11474 ( .B1(n8912), .B2(n11550), .A(n11796), .ZN(n8914) );
  NAND2_X1 U11475 ( .A1(n8914), .A2(n8913), .ZN(n8915) );
  INV_X1 U11476 ( .A(n11797), .ZN(n8918) );
  AND2_X1 U11477 ( .A1(n8920), .A2(n8919), .ZN(n8922) );
  NAND2_X1 U11478 ( .A1(n10220), .A2(n12734), .ZN(n8930) );
  INV_X1 U11479 ( .A(n8923), .ZN(n8925) );
  NOR2_X1 U11480 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n8924) );
  NAND2_X1 U11481 ( .A1(n8925), .A2(n8924), .ZN(n8927) );
  NAND2_X1 U11482 ( .A1(n8927), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8926) );
  MUX2_X1 U11483 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8926), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n8928) );
  AOI22_X1 U11484 ( .A1(n12733), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9123), 
        .B2(n10730), .ZN(n8929) );
  NAND2_X1 U11485 ( .A1(n8930), .A2(n8929), .ZN(n14675) );
  INV_X1 U11486 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10623) );
  OR2_X1 U11487 ( .A1(n8889), .A2(n10623), .ZN(n8934) );
  INV_X1 U11488 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8947) );
  XNOR2_X1 U11489 ( .A(n8948), .B(n8947), .ZN(n11246) );
  OR2_X1 U11490 ( .A1(n8961), .A2(n11246), .ZN(n8933) );
  INV_X1 U11491 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11106) );
  OR2_X1 U11492 ( .A1(n8931), .A2(n11106), .ZN(n8932) );
  NAND4_X1 U11493 ( .A1(n8935), .A2(n8934), .A3(n8933), .A4(n8932), .ZN(n14238) );
  XNOR2_X1 U11494 ( .A(n14675), .B(n14238), .ZN(n12967) );
  NAND2_X1 U11495 ( .A1(n11101), .A2(n12967), .ZN(n11100) );
  INV_X1 U11496 ( .A(n14238), .ZN(n9343) );
  NAND2_X1 U11497 ( .A1(n9343), .A2(n14675), .ZN(n11399) );
  XNOR2_X1 U11498 ( .A(n8937), .B(n8936), .ZN(n10222) );
  NAND2_X1 U11499 ( .A1(n10222), .A2(n12734), .ZN(n8944) );
  NAND2_X1 U11500 ( .A1(n8939), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8938) );
  MUX2_X1 U11501 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8938), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n8942) );
  INV_X1 U11502 ( .A(n8939), .ZN(n8941) );
  INV_X1 U11503 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n8940) );
  NAND2_X1 U11504 ( .A1(n8941), .A2(n8940), .ZN(n8956) );
  NAND2_X1 U11505 ( .A1(n8942), .A2(n8956), .ZN(n10658) );
  INV_X1 U11506 ( .A(n10658), .ZN(n10689) );
  AOI22_X1 U11507 ( .A1(n12733), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n9123), 
        .B2(n10689), .ZN(n8943) );
  NAND2_X1 U11508 ( .A1(n8944), .A2(n8943), .ZN(n12807) );
  NAND2_X1 U11509 ( .A1(n12737), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8953) );
  INV_X1 U11510 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n8945) );
  OR2_X1 U11511 ( .A1(n8891), .A2(n8945), .ZN(n8952) );
  INV_X1 U11512 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8946) );
  OAI21_X1 U11513 ( .B1(n8948), .B2(n8947), .A(n8946), .ZN(n8949) );
  NAND2_X1 U11514 ( .A1(n8949), .A2(n8962), .ZN(n11670) );
  OR2_X1 U11515 ( .A1(n8961), .A2(n11670), .ZN(n8951) );
  INV_X1 U11516 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11404) );
  OR2_X1 U11517 ( .A1(n8931), .A2(n11404), .ZN(n8950) );
  NAND2_X1 U11518 ( .A1(n12807), .A2(n12809), .ZN(n11745) );
  XNOR2_X1 U11519 ( .A(n8954), .B(n8955), .ZN(n10489) );
  NAND2_X1 U11520 ( .A1(n10489), .A2(n12734), .ZN(n8960) );
  NAND2_X1 U11521 ( .A1(n8956), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8957) );
  MUX2_X1 U11522 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8957), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n8958) );
  AND2_X1 U11523 ( .A1(n8958), .A2(n8973), .ZN(n10717) );
  AOI22_X1 U11524 ( .A1(n12733), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n9123), 
        .B2(n10717), .ZN(n8959) );
  NAND2_X1 U11525 ( .A1(n12737), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8967) );
  INV_X1 U11526 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10355) );
  OR2_X1 U11527 ( .A1(n8891), .A2(n10355), .ZN(n8966) );
  INV_X1 U11528 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10256) );
  NAND2_X1 U11529 ( .A1(n8962), .A2(n10256), .ZN(n8963) );
  NAND2_X1 U11530 ( .A1(n8979), .A2(n8963), .ZN(n11910) );
  OR2_X1 U11531 ( .A1(n8961), .A2(n11910), .ZN(n8965) );
  INV_X1 U11532 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10690) );
  OR2_X1 U11533 ( .A1(n8931), .A2(n10690), .ZN(n8964) );
  NAND4_X1 U11534 ( .A1(n8967), .A2(n8966), .A3(n8965), .A4(n8964), .ZN(n14236) );
  OR2_X1 U11535 ( .A1(n12807), .A2(n12809), .ZN(n11743) );
  NAND2_X1 U11536 ( .A1(n8968), .A2(n8085), .ZN(n8971) );
  INV_X1 U11537 ( .A(n14236), .ZN(n8969) );
  NAND2_X1 U11538 ( .A1(n14668), .A2(n8969), .ZN(n8970) );
  NAND2_X1 U11539 ( .A1(n8971), .A2(n8970), .ZN(n11363) );
  NAND2_X1 U11540 ( .A1(n10510), .A2(n12734), .ZN(n8976) );
  NAND2_X1 U11541 ( .A1(n8973), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8974) );
  XNOR2_X1 U11542 ( .A(n8974), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10804) );
  AOI22_X1 U11543 ( .A1(n12733), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n9123), 
        .B2(n10804), .ZN(n8975) );
  NAND2_X1 U11544 ( .A1(n9283), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8984) );
  INV_X1 U11545 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n8977) );
  OR2_X1 U11546 ( .A1(n8889), .A2(n8977), .ZN(n8983) );
  NAND2_X1 U11547 ( .A1(n8979), .A2(n8978), .ZN(n8980) );
  NAND2_X1 U11548 ( .A1(n8994), .A2(n8980), .ZN(n12149) );
  OR2_X1 U11549 ( .A1(n8961), .A2(n12149), .ZN(n8982) );
  INV_X1 U11550 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11367) );
  OR2_X1 U11551 ( .A1(n8931), .A2(n11367), .ZN(n8981) );
  AND2_X1 U11552 ( .A1(n14663), .A2(n12820), .ZN(n8985) );
  XNOR2_X1 U11553 ( .A(n8986), .B(SI_10_), .ZN(n8987) );
  XNOR2_X1 U11554 ( .A(n8988), .B(n8987), .ZN(n10572) );
  NAND2_X1 U11555 ( .A1(n10572), .A2(n12734), .ZN(n8992) );
  NAND2_X1 U11556 ( .A1(n6679), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8989) );
  MUX2_X1 U11557 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8989), .S(
        P2_IR_REG_10__SCAN_IN), .Z(n8990) );
  NAND2_X1 U11558 ( .A1(n8990), .A2(n9303), .ZN(n10807) );
  AOI22_X1 U11559 ( .A1(n12733), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n9123), 
        .B2(n15830), .ZN(n8991) );
  NAND2_X1 U11560 ( .A1(n9283), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n9000) );
  INV_X1 U11561 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10387) );
  OR2_X1 U11562 ( .A1(n8889), .A2(n10387), .ZN(n8999) );
  INV_X1 U11563 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8993) );
  NAND2_X1 U11564 ( .A1(n8994), .A2(n8993), .ZN(n8995) );
  NAND2_X1 U11565 ( .A1(n9011), .A2(n8995), .ZN(n12400) );
  OR2_X1 U11566 ( .A1(n8961), .A2(n12400), .ZN(n8998) );
  INV_X1 U11567 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8996) );
  OR2_X1 U11568 ( .A1(n8931), .A2(n8996), .ZN(n8997) );
  XNOR2_X1 U11569 ( .A(n12818), .B(n12817), .ZN(n12973) );
  NAND2_X1 U11570 ( .A1(n12818), .A2(n12817), .ZN(n12159) );
  NAND2_X1 U11571 ( .A1(n9032), .A2(n9003), .ZN(n9004) );
  NAND2_X1 U11572 ( .A1(n9005), .A2(n9004), .ZN(n9006) );
  NAND2_X1 U11573 ( .A1(n9033), .A2(n9006), .ZN(n10613) );
  NAND2_X1 U11574 ( .A1(n10613), .A2(n12734), .ZN(n9009) );
  NAND2_X1 U11575 ( .A1(n9303), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9007) );
  XNOR2_X1 U11576 ( .A(n9007), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10810) );
  AOI22_X1 U11577 ( .A1(n12733), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n9123), 
        .B2(n10810), .ZN(n9008) );
  NAND2_X1 U11578 ( .A1(n12737), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9017) );
  INV_X1 U11579 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9010) );
  OR2_X1 U11580 ( .A1(n8891), .A2(n9010), .ZN(n9016) );
  NAND2_X1 U11581 ( .A1(n9011), .A2(n10802), .ZN(n9012) );
  NAND2_X1 U11582 ( .A1(n9042), .A2(n9012), .ZN(n14177) );
  OR2_X1 U11583 ( .A1(n8961), .A2(n14177), .ZN(n9015) );
  INV_X1 U11584 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n9013) );
  OR2_X1 U11585 ( .A1(n8931), .A2(n9013), .ZN(n9014) );
  NAND4_X1 U11586 ( .A1(n9017), .A2(n9016), .A3(n9015), .A4(n9014), .ZN(n14233) );
  XNOR2_X1 U11587 ( .A(n14658), .B(n14233), .ZN(n12975) );
  INV_X1 U11588 ( .A(n14233), .ZN(n14092) );
  NAND2_X1 U11589 ( .A1(n14658), .A2(n14092), .ZN(n14527) );
  AND2_X1 U11590 ( .A1(n9079), .A2(n9060), .ZN(n9058) );
  XNOR2_X1 U11591 ( .A(n9059), .B(n9058), .ZN(n10702) );
  NAND2_X1 U11592 ( .A1(n10702), .A2(n12734), .ZN(n9025) );
  OR2_X1 U11593 ( .A1(n9303), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n9036) );
  NAND2_X1 U11594 ( .A1(n9019), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9018) );
  MUX2_X1 U11595 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9018), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n9022) );
  INV_X1 U11596 ( .A(n9019), .ZN(n9021) );
  INV_X1 U11597 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n9020) );
  NAND2_X1 U11598 ( .A1(n9021), .A2(n9020), .ZN(n9080) );
  NAND2_X1 U11599 ( .A1(n9022), .A2(n9080), .ZN(n11535) );
  OAI22_X1 U11600 ( .A1(n8902), .A2(n10703), .B1(n11535), .B2(n7327), .ZN(
        n9023) );
  INV_X1 U11601 ( .A(n9023), .ZN(n9024) );
  NAND2_X1 U11602 ( .A1(n9283), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n9031) );
  INV_X1 U11603 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n14649) );
  OR2_X1 U11604 ( .A1(n8889), .A2(n14649), .ZN(n9030) );
  NAND2_X1 U11605 ( .A1(n9044), .A2(n9026), .ZN(n9027) );
  NAND2_X1 U11606 ( .A1(n9068), .A2(n9027), .ZN(n14538) );
  OR2_X1 U11607 ( .A1(n8961), .A2(n14538), .ZN(n9029) );
  INV_X1 U11608 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n14539) );
  OR2_X1 U11609 ( .A1(n8931), .A2(n14539), .ZN(n9028) );
  NAND2_X1 U11610 ( .A1(n14648), .A2(n14091), .ZN(n12959) );
  NAND2_X1 U11611 ( .A1(n10678), .A2(n12734), .ZN(n9039) );
  NAND2_X1 U11612 ( .A1(n9036), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9037) );
  XNOR2_X1 U11613 ( .A(n9037), .B(P2_IR_REG_12__SCAN_IN), .ZN(n11005) );
  AOI22_X1 U11614 ( .A1(n12733), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n9123), 
        .B2(n11005), .ZN(n9038) );
  NAND2_X1 U11615 ( .A1(n9283), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9048) );
  INV_X1 U11616 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9040) );
  OR2_X1 U11617 ( .A1(n8889), .A2(n9040), .ZN(n9047) );
  INV_X1 U11618 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9041) );
  NAND2_X1 U11619 ( .A1(n9042), .A2(n9041), .ZN(n9043) );
  NAND2_X1 U11620 ( .A1(n9044), .A2(n9043), .ZN(n14559) );
  OR2_X1 U11621 ( .A1(n8961), .A2(n14559), .ZN(n9046) );
  OR2_X1 U11622 ( .A1(n8931), .A2(n10902), .ZN(n9045) );
  AND2_X1 U11623 ( .A1(n14527), .A2(n9050), .ZN(n9049) );
  NAND2_X1 U11624 ( .A1(n12158), .A2(n9049), .ZN(n9053) );
  OR2_X1 U11625 ( .A1(n14648), .A2(n14091), .ZN(n12958) );
  INV_X1 U11626 ( .A(n9060), .ZN(n9054) );
  OR2_X1 U11627 ( .A1(n9055), .A2(n9054), .ZN(n9056) );
  NAND2_X1 U11628 ( .A1(n9059), .A2(n9058), .ZN(n9062) );
  AND2_X1 U11629 ( .A1(SI_14_), .A2(n9060), .ZN(n9061) );
  NAND2_X1 U11630 ( .A1(n9062), .A2(n9061), .ZN(n9063) );
  NAND2_X1 U11631 ( .A1(n10784), .A2(n12734), .ZN(n9066) );
  NAND2_X1 U11632 ( .A1(n9080), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9064) );
  XNOR2_X1 U11633 ( .A(n9064), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11653) );
  AOI22_X1 U11634 ( .A1(n11653), .A2(n9123), .B1(n12733), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n9065) );
  NAND2_X2 U11635 ( .A1(n9066), .A2(n9065), .ZN(n14643) );
  NAND2_X1 U11636 ( .A1(n9068), .A2(n9067), .ZN(n9069) );
  AND2_X1 U11637 ( .A1(n9087), .A2(n9069), .ZN(n14047) );
  NAND2_X1 U11638 ( .A1(n9218), .A2(n14047), .ZN(n9073) );
  INV_X1 U11639 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14728) );
  OR2_X1 U11640 ( .A1(n8891), .A2(n14728), .ZN(n9072) );
  INV_X1 U11641 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n14644) );
  OR2_X1 U11642 ( .A1(n8889), .A2(n14644), .ZN(n9071) );
  INV_X1 U11643 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n14518) );
  OR2_X1 U11644 ( .A1(n8931), .A2(n14518), .ZN(n9070) );
  INV_X1 U11645 ( .A(n14643), .ZN(n12850) );
  INV_X1 U11646 ( .A(n14203), .ZN(n14232) );
  NAND2_X1 U11647 ( .A1(n9723), .A2(n12734), .ZN(n9083) );
  NAND2_X1 U11648 ( .A1(n9094), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9081) );
  XNOR2_X1 U11649 ( .A(n9081), .B(P2_IR_REG_15__SCAN_IN), .ZN(n11979) );
  AOI22_X1 U11650 ( .A1(n11979), .A2(n9123), .B1(n12733), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n9082) );
  INV_X1 U11651 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14639) );
  OR2_X1 U11652 ( .A1(n8889), .A2(n14639), .ZN(n9085) );
  INV_X1 U11653 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n14724) );
  OR2_X1 U11654 ( .A1(n8891), .A2(n14724), .ZN(n9084) );
  AND2_X1 U11655 ( .A1(n9085), .A2(n9084), .ZN(n9091) );
  INV_X1 U11656 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9086) );
  NAND2_X1 U11657 ( .A1(n9087), .A2(n9086), .ZN(n9088) );
  NAND2_X1 U11658 ( .A1(n9099), .A2(n9088), .ZN(n14507) );
  OR2_X1 U11659 ( .A1(n14507), .A2(n8961), .ZN(n9090) );
  NAND2_X1 U11660 ( .A1(n9266), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n9089) );
  NAND2_X1 U11661 ( .A1(n10708), .A2(n12734), .ZN(n9097) );
  OAI21_X1 U11662 ( .B1(n9094), .B2(P2_IR_REG_15__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9095) );
  INV_X1 U11663 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n10437) );
  XNOR2_X1 U11664 ( .A(n9095), .B(P2_IR_REG_16__SCAN_IN), .ZN(n12198) );
  AOI22_X1 U11665 ( .A1(n12198), .A2(n9123), .B1(n12733), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n9096) );
  NAND2_X2 U11666 ( .A1(n9097), .A2(n9096), .ZN(n14631) );
  INV_X1 U11667 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9098) );
  NAND2_X1 U11668 ( .A1(n9099), .A2(n9098), .ZN(n9100) );
  NAND2_X1 U11669 ( .A1(n9113), .A2(n9100), .ZN(n14490) );
  OR2_X1 U11670 ( .A1(n14490), .A2(n8961), .ZN(n9103) );
  AOI22_X1 U11671 ( .A1(n12737), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n9283), 
        .B2(P2_REG0_REG_16__SCAN_IN), .ZN(n9102) );
  NAND2_X1 U11672 ( .A1(n9266), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n9101) );
  OR2_X1 U11673 ( .A1(n14631), .A2(n14205), .ZN(n9104) );
  XNOR2_X1 U11674 ( .A(n9105), .B(SI_17_), .ZN(n9106) );
  XNOR2_X1 U11675 ( .A(n9107), .B(n9106), .ZN(n10758) );
  NAND2_X1 U11676 ( .A1(n10758), .A2(n12734), .ZN(n9111) );
  NAND2_X1 U11677 ( .A1(n6760), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9108) );
  MUX2_X1 U11678 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9108), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n9109) );
  INV_X1 U11679 ( .A(n9323), .ZN(n9332) );
  AOI22_X1 U11680 ( .A1(n12733), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n9123), 
        .B2(n12341), .ZN(n9110) );
  NAND2_X2 U11681 ( .A1(n9111), .A2(n9110), .ZN(n14626) );
  NAND2_X1 U11682 ( .A1(n9113), .A2(n9112), .ZN(n9114) );
  AND2_X1 U11683 ( .A1(n9127), .A2(n9114), .ZN(n14468) );
  NAND2_X1 U11684 ( .A1(n14468), .A2(n9218), .ZN(n9117) );
  AOI22_X1 U11685 ( .A1(n9266), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n9283), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n9116) );
  NAND2_X1 U11686 ( .A1(n12737), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n9115) );
  NAND2_X1 U11687 ( .A1(n14626), .A2(n14183), .ZN(n12864) );
  OR2_X1 U11688 ( .A1(n14626), .A2(n14183), .ZN(n14473) );
  NAND2_X1 U11689 ( .A1(n14475), .A2(n14473), .ZN(n14450) );
  NAND2_X1 U11690 ( .A1(n9119), .A2(n9118), .ZN(n9120) );
  NAND2_X1 U11691 ( .A1(n9121), .A2(n9120), .ZN(n10892) );
  OR2_X1 U11692 ( .A1(n10892), .A2(n9169), .ZN(n9125) );
  NAND2_X1 U11693 ( .A1(n9332), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9122) );
  XNOR2_X1 U11694 ( .A(n9122), .B(P2_IR_REG_18__SCAN_IN), .ZN(n14289) );
  AOI22_X1 U11695 ( .A1(n12733), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n9123), 
        .B2(n14289), .ZN(n9124) );
  NAND2_X2 U11696 ( .A1(n9125), .A2(n9124), .ZN(n14620) );
  INV_X1 U11697 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9126) );
  NAND2_X1 U11698 ( .A1(n9127), .A2(n9126), .ZN(n9128) );
  NAND2_X1 U11699 ( .A1(n9129), .A2(n9128), .ZN(n14456) );
  OR2_X1 U11700 ( .A1(n14456), .A2(n8961), .ZN(n9135) );
  INV_X1 U11701 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9132) );
  NAND2_X1 U11702 ( .A1(n12737), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9131) );
  NAND2_X1 U11703 ( .A1(n9283), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n9130) );
  OAI211_X1 U11704 ( .C1(n9132), .C2(n8931), .A(n9131), .B(n9130), .ZN(n9133)
         );
  INV_X1 U11705 ( .A(n9133), .ZN(n9134) );
  NAND2_X1 U11706 ( .A1(n14620), .A2(n12884), .ZN(n9136) );
  NAND2_X1 U11707 ( .A1(n9151), .A2(n9137), .ZN(n9139) );
  NAND2_X1 U11708 ( .A1(n9139), .A2(n9138), .ZN(n9140) );
  OR2_X1 U11709 ( .A1(n12408), .A2(n9169), .ZN(n9142) );
  OR2_X1 U11710 ( .A1(n8902), .A2(n12407), .ZN(n9141) );
  INV_X1 U11711 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9143) );
  NAND2_X1 U11712 ( .A1(n9144), .A2(n9143), .ZN(n9145) );
  NAND2_X1 U11713 ( .A1(n9157), .A2(n9145), .ZN(n14432) );
  OR2_X1 U11714 ( .A1(n14432), .A2(n8961), .ZN(n9150) );
  INV_X1 U11715 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n14431) );
  NAND2_X1 U11716 ( .A1(n9283), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n9147) );
  NAND2_X1 U11717 ( .A1(n12737), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n9146) );
  OAI211_X1 U11718 ( .C1(n14431), .C2(n8931), .A(n9147), .B(n9146), .ZN(n9148)
         );
  INV_X1 U11719 ( .A(n9148), .ZN(n9149) );
  XNOR2_X1 U11720 ( .A(n14610), .B(n14226), .ZN(n14424) );
  NAND2_X1 U11721 ( .A1(n9153), .A2(n9152), .ZN(n9154) );
  OR2_X1 U11722 ( .A1(n8902), .A2(n11111), .ZN(n9156) );
  NAND2_X1 U11723 ( .A1(n9157), .A2(n14081), .ZN(n9158) );
  AND2_X1 U11724 ( .A1(n9172), .A2(n9158), .ZN(n14417) );
  NAND2_X1 U11725 ( .A1(n14417), .A2(n9218), .ZN(n9164) );
  INV_X1 U11726 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9161) );
  NAND2_X1 U11727 ( .A1(n12737), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n9160) );
  NAND2_X1 U11728 ( .A1(n9283), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n9159) );
  OAI211_X1 U11729 ( .C1(n9161), .C2(n8931), .A(n9160), .B(n9159), .ZN(n9162)
         );
  INV_X1 U11730 ( .A(n9162), .ZN(n9163) );
  NAND2_X1 U11731 ( .A1(n14605), .A2(n14165), .ZN(n9165) );
  NAND2_X1 U11732 ( .A1(n9166), .A2(SI_22_), .ZN(n9179) );
  OR2_X1 U11733 ( .A1(n9833), .A2(n9167), .ZN(n9180) );
  NAND2_X1 U11734 ( .A1(n9833), .A2(n9167), .ZN(n9168) );
  NAND2_X1 U11735 ( .A1(n9180), .A2(n9168), .ZN(n11133) );
  OR2_X1 U11736 ( .A1(n11133), .A2(n9169), .ZN(n9171) );
  OR2_X1 U11737 ( .A1(n8902), .A2(n11132), .ZN(n9170) );
  INV_X1 U11738 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n14167) );
  NAND2_X1 U11739 ( .A1(n9172), .A2(n14167), .ZN(n9173) );
  NAND2_X1 U11740 ( .A1(n9186), .A2(n9173), .ZN(n14401) );
  OR2_X1 U11741 ( .A1(n14401), .A2(n8961), .ZN(n9178) );
  INV_X1 U11742 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n14400) );
  NAND2_X1 U11743 ( .A1(n12737), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n9175) );
  NAND2_X1 U11744 ( .A1(n9283), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9174) );
  OAI211_X1 U11745 ( .C1(n14400), .C2(n8931), .A(n9175), .B(n9174), .ZN(n9176)
         );
  INV_X1 U11746 ( .A(n9176), .ZN(n9177) );
  XNOR2_X1 U11747 ( .A(n14600), .B(n14059), .ZN(n14398) );
  NAND2_X1 U11748 ( .A1(n9180), .A2(n9179), .ZN(n9183) );
  XNOR2_X1 U11749 ( .A(n9181), .B(SI_23_), .ZN(n9182) );
  NAND2_X1 U11750 ( .A1(n11458), .A2(n12734), .ZN(n9185) );
  OR2_X1 U11751 ( .A1(n8902), .A2(n11457), .ZN(n9184) );
  INV_X1 U11752 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n14060) );
  NAND2_X1 U11753 ( .A1(n9186), .A2(n14060), .ZN(n9187) );
  NAND2_X1 U11754 ( .A1(n9195), .A2(n9187), .ZN(n14383) );
  OR2_X1 U11755 ( .A1(n14383), .A2(n8961), .ZN(n9192) );
  INV_X1 U11756 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n14374) );
  NAND2_X1 U11757 ( .A1(n12737), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n9189) );
  NAND2_X1 U11758 ( .A1(n9283), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n9188) );
  OAI211_X1 U11759 ( .C1(n14374), .C2(n8931), .A(n9189), .B(n9188), .ZN(n9190)
         );
  INV_X1 U11760 ( .A(n9190), .ZN(n9191) );
  INV_X1 U11761 ( .A(n9193), .ZN(n9194) );
  NAND2_X1 U11762 ( .A1(n9195), .A2(n14133), .ZN(n9196) );
  NAND2_X1 U11763 ( .A1(n9216), .A2(n9196), .ZN(n14357) );
  INV_X1 U11764 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n14691) );
  NAND2_X1 U11765 ( .A1(n12737), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n9198) );
  NAND2_X1 U11766 ( .A1(n9266), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9197) );
  OAI211_X1 U11767 ( .C1(n8891), .C2(n14691), .A(n9198), .B(n9197), .ZN(n9199)
         );
  INV_X1 U11768 ( .A(n9199), .ZN(n9200) );
  NAND2_X1 U11769 ( .A1(n9203), .A2(n9202), .ZN(n9204) );
  OR2_X1 U11770 ( .A1(n8902), .A2(n11770), .ZN(n9206) );
  XOR2_X1 U11771 ( .A(n14222), .B(n14590), .Z(n14354) );
  INV_X1 U11772 ( .A(n14590), .ZN(n12765) );
  XNOR2_X1 U11773 ( .A(n14585), .B(n14221), .ZN(n14337) );
  MUX2_X1 U11774 ( .A(n12219), .B(n12221), .S(n9260), .Z(n9232) );
  XNOR2_X1 U11775 ( .A(n9232), .B(SI_26_), .ZN(n9211) );
  XNOR2_X1 U11776 ( .A(n9234), .B(n9211), .ZN(n12218) );
  NAND2_X1 U11777 ( .A1(n12218), .A2(n12734), .ZN(n9213) );
  OR2_X1 U11778 ( .A1(n8902), .A2(n12221), .ZN(n9212) );
  INV_X1 U11779 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n14102) );
  INV_X1 U11780 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9214) );
  OAI21_X1 U11781 ( .B1(n9216), .B2(n14102), .A(n9214), .ZN(n9217) );
  NAND2_X1 U11782 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n9215) );
  NAND2_X1 U11783 ( .A1(n14326), .A2(n9218), .ZN(n9224) );
  INV_X1 U11784 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9221) );
  NAND2_X1 U11785 ( .A1(n12737), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n9220) );
  OAI211_X1 U11786 ( .C1(n9221), .C2(n8931), .A(n9220), .B(n9219), .ZN(n9222)
         );
  INV_X1 U11787 ( .A(n9222), .ZN(n9223) );
  OR2_X1 U11788 ( .A1(n14327), .A2(n14101), .ZN(n12957) );
  AND2_X1 U11789 ( .A1(n14327), .A2(n14101), .ZN(n12956) );
  INV_X1 U11790 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13205) );
  NAND2_X1 U11791 ( .A1(n9225), .A2(n13205), .ZN(n9226) );
  NAND2_X1 U11792 ( .A1(n9250), .A2(n9226), .ZN(n14311) );
  INV_X1 U11793 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n14310) );
  NAND2_X1 U11794 ( .A1(n12737), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n9228) );
  OAI211_X1 U11795 ( .C1(n14310), .C2(n8931), .A(n9228), .B(n9227), .ZN(n9229)
         );
  INV_X1 U11796 ( .A(n9229), .ZN(n9230) );
  NAND2_X2 U11797 ( .A1(n9231), .A2(n9230), .ZN(n14219) );
  NOR2_X1 U11798 ( .A1(n9235), .A2(SI_26_), .ZN(n9233) );
  MUX2_X1 U11799 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n9260), .Z(n9241) );
  XNOR2_X1 U11800 ( .A(n9241), .B(SI_27_), .ZN(n9236) );
  NAND2_X1 U11801 ( .A1(n12267), .A2(n12734), .ZN(n9239) );
  OR2_X1 U11802 ( .A1(n8902), .A2(n9237), .ZN(n9238) );
  INV_X1 U11803 ( .A(n9241), .ZN(n9240) );
  MUX2_X1 U11804 ( .A(n13185), .B(n12286), .S(n10481), .Z(n9257) );
  XNOR2_X1 U11805 ( .A(n9257), .B(SI_28_), .ZN(n9243) );
  NAND2_X1 U11806 ( .A1(n9244), .A2(n9243), .ZN(n9259) );
  OR2_X1 U11807 ( .A1(n9244), .A2(n9243), .ZN(n9245) );
  NAND2_X1 U11808 ( .A1(n9259), .A2(n9245), .ZN(n13184) );
  NAND2_X1 U11809 ( .A1(n13184), .A2(n12734), .ZN(n9247) );
  OR2_X1 U11810 ( .A1(n8902), .A2(n12286), .ZN(n9246) );
  INV_X1 U11811 ( .A(n9250), .ZN(n9248) );
  NAND2_X1 U11812 ( .A1(n9248), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n12716) );
  INV_X1 U11813 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9249) );
  NAND2_X1 U11814 ( .A1(n9250), .A2(n9249), .ZN(n9251) );
  NAND2_X1 U11815 ( .A1(n12716), .A2(n9251), .ZN(n13173) );
  INV_X1 U11816 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n10458) );
  NAND2_X1 U11817 ( .A1(n9266), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9253) );
  NAND2_X1 U11818 ( .A1(n9283), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9252) );
  OAI211_X1 U11819 ( .C1(n8889), .C2(n10458), .A(n9253), .B(n9252), .ZN(n9254)
         );
  INV_X1 U11820 ( .A(n9254), .ZN(n9255) );
  NAND2_X1 U11821 ( .A1(n13180), .A2(n14218), .ZN(n9372) );
  OR2_X1 U11822 ( .A1(n13180), .A2(n14218), .ZN(n9256) );
  INV_X1 U11823 ( .A(SI_28_), .ZN(n14041) );
  NAND2_X1 U11824 ( .A1(n9257), .A2(n14041), .ZN(n9258) );
  NAND2_X1 U11825 ( .A1(n9259), .A2(n9258), .ZN(n9262) );
  INV_X1 U11826 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13194) );
  MUX2_X1 U11827 ( .A(n13003), .B(n13194), .S(n9260), .Z(n12589) );
  XNOR2_X1 U11828 ( .A(n12589), .B(SI_29_), .ZN(n9261) );
  OR2_X1 U11829 ( .A1(n9262), .A2(n9261), .ZN(n9263) );
  NAND2_X1 U11830 ( .A1(n12591), .A2(n9263), .ZN(n13002) );
  NAND2_X1 U11831 ( .A1(n13002), .A2(n12734), .ZN(n9265) );
  OR2_X1 U11832 ( .A1(n8902), .A2(n13194), .ZN(n9264) );
  OR2_X1 U11833 ( .A1(n12716), .A2(n8961), .ZN(n9271) );
  NAND2_X1 U11834 ( .A1(n9266), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9268) );
  NAND2_X1 U11835 ( .A1(n12737), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n9267) );
  OAI211_X1 U11836 ( .C1(n10412), .C2(n8891), .A(n9268), .B(n9267), .ZN(n9269)
         );
  INV_X1 U11837 ( .A(n9269), .ZN(n9270) );
  XNOR2_X1 U11838 ( .A(n12926), .B(n12924), .ZN(n12984) );
  NAND2_X1 U11839 ( .A1(n8813), .A2(n9274), .ZN(n9301) );
  NAND2_X1 U11840 ( .A1(n6603), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9275) );
  MUX2_X1 U11841 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9275), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n9276) );
  NAND2_X1 U11842 ( .A1(n9290), .A2(n12988), .ZN(n9278) );
  NAND2_X1 U11843 ( .A1(n14299), .A2(n12763), .ZN(n9277) );
  NAND2_X1 U11844 ( .A1(n12919), .A2(n14218), .ZN(n9279) );
  NOR2_X1 U11845 ( .A1(n12984), .A2(n9280), .ZN(n9281) );
  INV_X1 U11846 ( .A(n9282), .ZN(n10638) );
  INV_X1 U11847 ( .A(n10637), .ZN(n10632) );
  INV_X1 U11848 ( .A(n10625), .ZN(n10839) );
  AOI21_X1 U11849 ( .B1(n10632), .B2(P2_B_REG_SCAN_IN), .A(n14204), .ZN(n12741) );
  INV_X1 U11850 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n12756) );
  NAND2_X1 U11851 ( .A1(n12737), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9285) );
  NAND2_X1 U11852 ( .A1(n9283), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9284) );
  OAI211_X1 U11853 ( .C1(n8931), .C2(n12756), .A(n9285), .B(n9284), .ZN(n14216) );
  NAND4_X1 U11854 ( .A1(n12984), .A2(n12919), .A3(n14218), .A4(n14556), .ZN(
        n9286) );
  NAND2_X1 U11855 ( .A1(n9290), .A2(n11110), .ZN(n12761) );
  INV_X1 U11856 ( .A(n9291), .ZN(n10874) );
  NAND2_X1 U11857 ( .A1(n14299), .A2(n10874), .ZN(n9289) );
  INV_X1 U11858 ( .A(n12770), .ZN(n11158) );
  INV_X1 U11859 ( .A(n14675), .ZN(n11098) );
  INV_X1 U11860 ( .A(n12807), .ZN(n12808) );
  INV_X1 U11861 ( .A(n14658), .ZN(n12815) );
  NAND2_X1 U11862 ( .A1(n12068), .A2(n12815), .ZN(n14558) );
  OR2_X2 U11863 ( .A1(n14557), .A2(n14648), .ZN(n14543) );
  NOR2_X4 U11864 ( .A1(n14543), .A2(n14643), .ZN(n14522) );
  NAND2_X1 U11865 ( .A1(n14455), .A2(n7128), .ZN(n14428) );
  OR2_X2 U11866 ( .A1(n14371), .A2(n14590), .ZN(n14359) );
  OR2_X2 U11867 ( .A1(n14359), .A2(n14585), .ZN(n14341) );
  NOR2_X4 U11868 ( .A1(n14341), .A2(n14327), .ZN(n14323) );
  NOR2_X2 U11869 ( .A1(n9291), .A2(n9290), .ZN(n10836) );
  OAI211_X1 U11870 ( .C1(n10015), .C2(n12925), .A(n10836), .B(n12752), .ZN(
        n12715) );
  OAI21_X1 U11871 ( .B1(n12925), .B2(n15879), .A(n12715), .ZN(n9292) );
  NOR4_X1 U11872 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n9296) );
  NOR4_X1 U11873 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n9295) );
  NOR4_X1 U11874 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9294) );
  NOR4_X1 U11875 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n9293) );
  NAND4_X1 U11876 ( .A1(n9296), .A2(n9295), .A3(n9294), .A4(n9293), .ZN(n9313)
         );
  NOR2_X1 U11877 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .ZN(
        n9300) );
  NOR4_X1 U11878 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n9299) );
  NOR4_X1 U11879 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n9298) );
  NOR4_X1 U11880 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9297) );
  NAND4_X1 U11881 ( .A1(n9300), .A2(n9299), .A3(n9298), .A4(n9297), .ZN(n9312)
         );
  OAI21_X1 U11882 ( .B1(n9307), .B2(P2_IR_REG_24__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9304) );
  MUX2_X1 U11883 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9304), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n9306) );
  NAND2_X1 U11884 ( .A1(n9306), .A2(n9305), .ZN(n12101) );
  NAND2_X1 U11885 ( .A1(n9307), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9308) );
  XOR2_X1 U11886 ( .A(n11768), .B(P2_B_REG_SCAN_IN), .Z(n9309) );
  NAND2_X1 U11887 ( .A1(n12101), .A2(n9309), .ZN(n9311) );
  NAND2_X1 U11888 ( .A1(n9305), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9310) );
  INV_X1 U11889 ( .A(n12223), .ZN(n9317) );
  OAI21_X1 U11890 ( .B1(n9313), .B2(n9312), .A(n15852), .ZN(n10832) );
  NOR2_X1 U11891 ( .A1(n12223), .A2(n12101), .ZN(n10045) );
  NAND2_X1 U11892 ( .A1(n11768), .A2(n10045), .ZN(n10628) );
  NAND2_X1 U11893 ( .A1(n12409), .A2(n12987), .ZN(n12931) );
  NAND2_X1 U11894 ( .A1(n12931), .A2(n10625), .ZN(n10834) );
  INV_X1 U11895 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15859) );
  NAND2_X1 U11896 ( .A1(n15852), .A2(n15859), .ZN(n9319) );
  OR2_X1 U11897 ( .A1(n11768), .A2(n9317), .ZN(n9318) );
  INV_X1 U11898 ( .A(n15860), .ZN(n10831) );
  INV_X1 U11899 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15862) );
  NAND2_X1 U11900 ( .A1(n15852), .A2(n15862), .ZN(n9321) );
  NAND2_X1 U11901 ( .A1(n12101), .A2(n12223), .ZN(n9320) );
  NOR2_X1 U11902 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), 
        .ZN(n9322) );
  NAND2_X1 U11903 ( .A1(n9323), .A2(n9322), .ZN(n9334) );
  AND2_X1 U11904 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .ZN(n9331) );
  INV_X1 U11905 ( .A(n9324), .ZN(n9328) );
  NAND2_X1 U11906 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .ZN(n9325) );
  NAND2_X1 U11907 ( .A1(n9325), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n9326) );
  NAND2_X1 U11908 ( .A1(n9326), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9327) );
  OAI211_X1 U11909 ( .C1(P2_IR_REG_31__SCAN_IN), .C2(n9329), .A(n9328), .B(
        n9327), .ZN(n9330) );
  AOI21_X1 U11910 ( .B1(n9332), .B2(n9331), .A(n9330), .ZN(n9333) );
  NAND2_X1 U11911 ( .A1(n15863), .A2(n10842), .ZN(n9375) );
  NOR2_X1 U11912 ( .A1(n10831), .A2(n9375), .ZN(n9335) );
  INV_X1 U11913 ( .A(n14610), .ZN(n9362) );
  INV_X1 U11914 ( .A(n12961), .ZN(n9336) );
  OR2_X1 U11915 ( .A1(n14242), .A2(n12784), .ZN(n10976) );
  OR2_X1 U11916 ( .A1(n12775), .A2(n6553), .ZN(n10975) );
  NAND3_X1 U11917 ( .A1(n11151), .A2(n10976), .A3(n10975), .ZN(n9339) );
  INV_X1 U11918 ( .A(n14242), .ZN(n9337) );
  NAND3_X1 U11919 ( .A1(n12965), .A2(n9339), .A3(n9338), .ZN(n10978) );
  OR2_X1 U11920 ( .A1(n14241), .A2(n12791), .ZN(n9340) );
  NAND2_X1 U11921 ( .A1(n10978), .A2(n9340), .ZN(n11546) );
  XNOR2_X1 U11922 ( .A(n14240), .B(n15873), .ZN(n12964) );
  NAND2_X1 U11923 ( .A1(n14675), .A2(n14238), .ZN(n11084) );
  NAND2_X1 U11924 ( .A1(n14239), .A2(n12799), .ZN(n9341) );
  NAND2_X1 U11925 ( .A1(n11084), .A2(n9341), .ZN(n11394) );
  OR2_X1 U11926 ( .A1(n14240), .A2(n12795), .ZN(n11085) );
  NOR2_X1 U11927 ( .A1(n11394), .A2(n11085), .ZN(n9346) );
  OAI21_X1 U11928 ( .B1(n14239), .B2(n12799), .A(n14238), .ZN(n9342) );
  NAND2_X1 U11929 ( .A1(n9342), .A2(n11098), .ZN(n9345) );
  NAND3_X1 U11930 ( .A1(n9343), .A2(n12800), .A3(n15880), .ZN(n9344) );
  NAND2_X1 U11931 ( .A1(n9345), .A2(n9344), .ZN(n11392) );
  NOR2_X1 U11932 ( .A1(n9346), .A2(n11392), .ZN(n9347) );
  XNOR2_X1 U11933 ( .A(n12807), .B(n12809), .ZN(n11400) );
  INV_X1 U11934 ( .A(n12809), .ZN(n14237) );
  NAND2_X1 U11935 ( .A1(n12807), .A2(n14237), .ZN(n9349) );
  NAND2_X1 U11936 ( .A1(n11396), .A2(n9349), .ZN(n11738) );
  INV_X1 U11937 ( .A(n12969), .ZN(n11737) );
  NAND2_X1 U11938 ( .A1(n11738), .A2(n11737), .ZN(n11740) );
  NAND2_X1 U11939 ( .A1(n14668), .A2(n14236), .ZN(n9350) );
  XNOR2_X1 U11940 ( .A(n14663), .B(n12820), .ZN(n12971) );
  INV_X1 U11941 ( .A(n12820), .ZN(n14235) );
  NAND2_X1 U11942 ( .A1(n14663), .A2(n14235), .ZN(n9351) );
  INV_X1 U11943 ( .A(n14648), .ZN(n12852) );
  NOR2_X1 U11944 ( .A1(n14648), .A2(n9355), .ZN(n9356) );
  XNOR2_X1 U11945 ( .A(n14500), .B(n14116), .ZN(n14501) );
  XNOR2_X1 U11946 ( .A(n14631), .B(n14205), .ZN(n14488) );
  XNOR2_X1 U11947 ( .A(n14626), .B(n14183), .ZN(n14476) );
  INV_X1 U11948 ( .A(n14183), .ZN(n14229) );
  NAND2_X1 U11949 ( .A1(n14626), .A2(n14229), .ZN(n9359) );
  XNOR2_X1 U11950 ( .A(n14620), .B(n12884), .ZN(n14454) );
  NAND2_X1 U11951 ( .A1(n14615), .A2(n14227), .ZN(n12977) );
  NAND2_X1 U11952 ( .A1(n9362), .A2(n9361), .ZN(n14409) );
  AND2_X1 U11953 ( .A1(n14409), .A2(n9364), .ZN(n14392) );
  AND2_X1 U11954 ( .A1(n14392), .A2(n14398), .ZN(n9363) );
  NAND2_X1 U11955 ( .A1(n14600), .A2(n14224), .ZN(n9366) );
  INV_X1 U11956 ( .A(n14398), .ZN(n12979) );
  INV_X1 U11957 ( .A(n9364), .ZN(n9365) );
  XNOR2_X1 U11958 ( .A(n14605), .B(n14165), .ZN(n14411) );
  OR2_X1 U11959 ( .A1(n9365), .A2(n14411), .ZN(n14393) );
  INV_X1 U11960 ( .A(n14379), .ZN(n14369) );
  NAND2_X1 U11961 ( .A1(n14375), .A2(n14166), .ZN(n9367) );
  INV_X1 U11962 ( .A(n14221), .ZN(n12909) );
  NAND2_X1 U11963 ( .A1(n14346), .A2(n12909), .ZN(n9368) );
  NAND2_X1 U11964 ( .A1(n14334), .A2(n9368), .ZN(n9370) );
  NAND2_X1 U11965 ( .A1(n14585), .A2(n14221), .ZN(n9369) );
  INV_X1 U11966 ( .A(n14327), .ZN(n14582) );
  NAND2_X1 U11967 ( .A1(n14582), .A2(n14101), .ZN(n9371) );
  INV_X1 U11968 ( .A(n14303), .ZN(n14309) );
  NAND2_X1 U11969 ( .A1(n12409), .A2(n12988), .ZN(n12767) );
  XNOR2_X1 U11970 ( .A(n12767), .B(n12763), .ZN(n9373) );
  NAND2_X1 U11971 ( .A1(n9373), .A2(n12987), .ZN(n14552) );
  NAND2_X1 U11972 ( .A1(n14552), .A2(n14673), .ZN(n15884) );
  NAND2_X1 U11973 ( .A1(n15886), .A2(n15884), .ZN(n14734) );
  INV_X1 U11974 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9378) );
  NOR2_X1 U11975 ( .A1(n9375), .A2(n15860), .ZN(n9376) );
  NAND2_X1 U11976 ( .A1(n15893), .A2(n15884), .ZN(n14651) );
  NAND2_X1 U11977 ( .A1(n9380), .A2(n9379), .ZN(P2_U3528) );
  NOR2_X1 U11978 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n9383) );
  NOR2_X1 U11979 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), 
        .ZN(n9387) );
  NAND3_X1 U11980 ( .A1(n9405), .A2(n9392), .A3(n9391), .ZN(n9393) );
  OR2_X1 U11981 ( .A1(n12408), .A2(n9779), .ZN(n9399) );
  OR2_X1 U11982 ( .A1(n12615), .A2(n10931), .ZN(n9398) );
  INV_X1 U11983 ( .A(n9400), .ZN(n9401) );
  XNOR2_X1 U11984 ( .A(n9402), .B(P1_IR_REG_26__SCAN_IN), .ZN(n9957) );
  NAND2_X1 U11985 ( .A1(n9409), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9403) );
  XNOR2_X1 U11986 ( .A(n9403), .B(P1_IR_REG_25__SCAN_IN), .ZN(n9973) );
  NAND3_X1 U11987 ( .A1(n9406), .A2(n9413), .A3(n9405), .ZN(n9407) );
  OR2_X1 U11988 ( .A1(n9404), .A2(n9407), .ZN(n9975) );
  OAI21_X1 U11989 ( .B1(n9975), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9408) );
  MUX2_X1 U11990 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9408), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n9410) );
  AND2_X4 U11991 ( .A1(n9477), .A2(n12438), .ZN(n9931) );
  INV_X1 U11992 ( .A(n9543), .ZN(n9416) );
  NAND2_X1 U11993 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_REG3_REG_14__SCAN_IN), 
        .ZN(n9417) );
  NAND2_X1 U11994 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .ZN(n9418) );
  NAND2_X1 U11995 ( .A1(n9804), .A2(n14866), .ZN(n9419) );
  NAND2_X1 U11996 ( .A1(n9823), .A2(n9419), .ZN(n15255) );
  XNOR2_X2 U11997 ( .A(n9421), .B(n15545), .ZN(n9427) );
  OR2_X1 U11998 ( .A1(n15255), .A2(n9907), .ZN(n9433) );
  INV_X1 U11999 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9430) );
  INV_X1 U12000 ( .A(n6544), .ZN(n9488) );
  NAND2_X1 U12001 ( .A1(n12583), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9429) );
  NAND2_X1 U12002 ( .A1(n12579), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9428) );
  OAI211_X1 U12003 ( .C1(n9927), .C2(n9430), .A(n9429), .B(n9428), .ZN(n9431)
         );
  INV_X1 U12004 ( .A(n9431), .ZN(n9432) );
  AND2_X4 U12005 ( .A1(n9923), .A2(n15733), .ZN(n9936) );
  AND2_X1 U12006 ( .A1(n14943), .A2(n6543), .ZN(n9436) );
  AOI21_X1 U12007 ( .B1(n15447), .B2(n9931), .A(n9436), .ZN(n9818) );
  INV_X1 U12008 ( .A(n9818), .ZN(n9820) );
  INV_X1 U12009 ( .A(n14943), .ZN(n13058) );
  OAI22_X1 U12010 ( .A1(n15252), .A2(n9954), .B1(n13058), .B2(n9677), .ZN(
        n9440) );
  NAND2_X1 U12011 ( .A1(n9404), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9438) );
  INV_X2 U12012 ( .A(n15112), .ZN(n15314) );
  AND2_X1 U12013 ( .A1(n6809), .A2(n15314), .ZN(n9439) );
  OR2_X2 U12014 ( .A1(n9439), .A2(n12438), .ZN(n9466) );
  XNOR2_X1 U12015 ( .A(n9440), .B(n10789), .ZN(n9819) );
  NAND2_X1 U12016 ( .A1(n10702), .A2(n12614), .ZN(n9444) );
  NAND2_X1 U12017 ( .A1(n9550), .A2(n6658), .ZN(n9667) );
  INV_X1 U12018 ( .A(n9667), .ZN(n9441) );
  NAND2_X1 U12019 ( .A1(n9441), .A2(n10239), .ZN(n9685) );
  NAND2_X1 U12020 ( .A1(n9708), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9442) );
  XNOR2_X1 U12021 ( .A(n9442), .B(P1_IR_REG_13__SCAN_IN), .ZN(n11482) );
  AOI22_X1 U12022 ( .A1(n9799), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n9798), 
        .B2(n11482), .ZN(n9443) );
  AND2_X2 U12023 ( .A1(n9444), .A2(n9443), .ZN(n15368) );
  OR2_X1 U12024 ( .A1(n15368), .A2(n9677), .ZN(n9453) );
  NAND2_X1 U12025 ( .A1(n12579), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n9451) );
  INV_X1 U12026 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11474) );
  OR2_X1 U12027 ( .A1(n9927), .A2(n11474), .ZN(n9450) );
  NAND2_X1 U12028 ( .A1(n9694), .A2(n9445), .ZN(n9446) );
  NAND2_X1 U12029 ( .A1(n9735), .A2(n9446), .ZN(n15364) );
  OR2_X1 U12030 ( .A1(n15364), .A2(n9907), .ZN(n9449) );
  INV_X1 U12031 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9447) );
  OR2_X1 U12032 ( .A1(n6545), .A2(n9447), .ZN(n9448) );
  NAND2_X1 U12033 ( .A1(n14949), .A2(n9936), .ZN(n9452) );
  NAND2_X1 U12034 ( .A1(n9453), .A2(n9452), .ZN(n9704) );
  INV_X1 U12035 ( .A(n9704), .ZN(n9707) );
  OAI22_X1 U12036 ( .A1(n15368), .A2(n9954), .B1(n14754), .B2(n9677), .ZN(
        n9454) );
  XNOR2_X1 U12037 ( .A(n9454), .B(n10789), .ZN(n9705) );
  INV_X1 U12038 ( .A(n9705), .ZN(n9706) );
  NAND2_X1 U12039 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9455) );
  INV_X1 U12040 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9457) );
  NAND2_X1 U12041 ( .A1(n12584), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9461) );
  INV_X1 U12042 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n11068) );
  INV_X1 U12043 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9458) );
  OR2_X1 U12044 ( .A1(n9509), .A2(n9458), .ZN(n9459) );
  NAND4_X1 U12045 ( .A1(n9462), .A2(n9461), .A3(n9460), .A4(n9459), .ZN(n9465)
         );
  NAND2_X1 U12046 ( .A1(n9465), .A2(n9931), .ZN(n9463) );
  XNOR2_X1 U12047 ( .A(n9464), .B(n9914), .ZN(n9482) );
  INV_X1 U12048 ( .A(n15732), .ZN(n11171) );
  INV_X1 U12049 ( .A(n9466), .ZN(n9743) );
  NAND2_X1 U12050 ( .A1(n12584), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9471) );
  INV_X1 U12051 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9467) );
  OR2_X1 U12052 ( .A1(n6544), .A2(n9467), .ZN(n9470) );
  INV_X1 U12053 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n15648) );
  INV_X1 U12054 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11296) );
  NAND2_X1 U12055 ( .A1(n14958), .A2(n9931), .ZN(n9480) );
  OAI21_X1 U12056 ( .B1(n10481), .B2(n9473), .A(P2_DATAO_REG_0__SCAN_IN), .ZN(
        n9472) );
  OAI21_X1 U12057 ( .B1(n9474), .B2(n9473), .A(n9472), .ZN(n10478) );
  INV_X1 U12058 ( .A(n10478), .ZN(n9476) );
  MUX2_X1 U12059 ( .A(n14964), .B(n9476), .S(n9475), .Z(n11298) );
  OAI22_X1 U12060 ( .A1(n11298), .A2(n9954), .B1(n9477), .B2(n15648), .ZN(
        n9478) );
  INV_X1 U12061 ( .A(n9478), .ZN(n9479) );
  NAND2_X1 U12062 ( .A1(n9480), .A2(n9479), .ZN(n10183) );
  OAI22_X1 U12063 ( .A1(n9501), .A2(n11298), .B1(n9477), .B2(n14964), .ZN(
        n9481) );
  INV_X1 U12064 ( .A(n9482), .ZN(n9484) );
  NAND2_X1 U12065 ( .A1(n9484), .A2(n9483), .ZN(n9485) );
  NAND2_X1 U12066 ( .A1(n9486), .A2(n9485), .ZN(n10825) );
  INV_X1 U12067 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9487) );
  INV_X1 U12068 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n11178) );
  OR2_X1 U12069 ( .A1(n9594), .A2(n11178), .ZN(n9492) );
  NAND2_X1 U12070 ( .A1(n9488), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9491) );
  INV_X1 U12071 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9489) );
  OR2_X1 U12072 ( .A1(n9990), .A2(n9489), .ZN(n9490) );
  NAND2_X1 U12073 ( .A1(n15638), .A2(n9931), .ZN(n9499) );
  INV_X1 U12074 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10491) );
  OR2_X1 U12075 ( .A1(n9494), .A2(n10491), .ZN(n9498) );
  NAND2_X1 U12076 ( .A1(n9496), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9495) );
  MUX2_X1 U12077 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9495), .S(
        P1_IR_REG_2__SCAN_IN), .Z(n9497) );
  NAND2_X1 U12078 ( .A1(n9497), .A2(n9514), .ZN(n10582) );
  XNOR2_X1 U12079 ( .A(n9500), .B(n9743), .ZN(n9506) );
  NAND2_X1 U12080 ( .A1(n15638), .A2(n9936), .ZN(n9503) );
  OR2_X1 U12081 ( .A1(n15743), .A2(n9501), .ZN(n9502) );
  NAND2_X1 U12082 ( .A1(n9503), .A2(n9502), .ZN(n9504) );
  XNOR2_X1 U12083 ( .A(n9506), .B(n9504), .ZN(n10826) );
  INV_X1 U12084 ( .A(n9504), .ZN(n9505) );
  NAND2_X1 U12085 ( .A1(n9506), .A2(n9505), .ZN(n9507) );
  OR2_X1 U12086 ( .A1(n9594), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9512) );
  INV_X1 U12087 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9508) );
  OR2_X1 U12088 ( .A1(n9990), .A2(n9508), .ZN(n9511) );
  INV_X1 U12089 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n15713) );
  OR2_X1 U12090 ( .A1(n6545), .A2(n15713), .ZN(n9510) );
  NAND2_X1 U12091 ( .A1(n14957), .A2(n9931), .ZN(n9517) );
  MUX2_X1 U12092 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9515), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n9516) );
  INV_X1 U12093 ( .A(n9550), .ZN(n9531) );
  NAND2_X1 U12094 ( .A1(n9516), .A2(n9531), .ZN(n14977) );
  INV_X1 U12095 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10214) );
  XNOR2_X1 U12096 ( .A(n9518), .B(n10789), .ZN(n9522) );
  NAND2_X1 U12097 ( .A1(n14957), .A2(n9936), .ZN(n9520) );
  OR2_X1 U12098 ( .A1(n15631), .A2(n9501), .ZN(n9519) );
  NAND2_X1 U12099 ( .A1(n9520), .A2(n9519), .ZN(n9521) );
  NAND2_X1 U12100 ( .A1(n9522), .A2(n9521), .ZN(n9539) );
  NAND2_X1 U12101 ( .A1(n9987), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9530) );
  INV_X1 U12102 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9525) );
  OR2_X1 U12103 ( .A1(n9990), .A2(n9525), .ZN(n9529) );
  OAI21_X1 U12104 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(P1_REG3_REG_4__SCAN_IN), 
        .A(n9543), .ZN(n11427) );
  OR2_X1 U12105 ( .A1(n9907), .A2(n11427), .ZN(n9528) );
  INV_X1 U12106 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9526) );
  OR2_X1 U12107 ( .A1(n6545), .A2(n9526), .ZN(n9527) );
  NAND2_X1 U12108 ( .A1(n9531), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9532) );
  XNOR2_X1 U12109 ( .A(n9532), .B(P1_IR_REG_4__SCAN_IN), .ZN(n10588) );
  AOI22_X1 U12110 ( .A1(n9799), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n9798), .B2(
        n10588), .ZN(n9534) );
  NAND2_X1 U12111 ( .A1(n10219), .A2(n12614), .ZN(n9533) );
  AOI22_X1 U12112 ( .A1(n6540), .A2(n9936), .B1(n9931), .B2(n15756), .ZN(n9540) );
  AND2_X1 U12113 ( .A1(n9539), .A2(n9540), .ZN(n9535) );
  NAND2_X1 U12114 ( .A1(n15642), .A2(n9535), .ZN(n10988) );
  NAND2_X1 U12115 ( .A1(n6540), .A2(n9931), .ZN(n9537) );
  NAND2_X1 U12116 ( .A1(n15756), .A2(n9923), .ZN(n9536) );
  NAND2_X1 U12117 ( .A1(n9537), .A2(n9536), .ZN(n9538) );
  XNOR2_X1 U12118 ( .A(n9538), .B(n10789), .ZN(n10992) );
  NAND2_X1 U12119 ( .A1(n10988), .A2(n10992), .ZN(n10989) );
  NAND2_X1 U12120 ( .A1(n15642), .A2(n9539), .ZN(n9542) );
  INV_X1 U12121 ( .A(n9540), .ZN(n9541) );
  NAND2_X1 U12122 ( .A1(n9542), .A2(n9541), .ZN(n10990) );
  NAND2_X1 U12123 ( .A1(n9987), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9548) );
  OR2_X1 U12124 ( .A1(n9990), .A2(n15769), .ZN(n9547) );
  INV_X1 U12125 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10259) );
  NAND2_X1 U12126 ( .A1(n9543), .A2(n10259), .ZN(n9544) );
  NAND2_X1 U12127 ( .A1(n9564), .A2(n9544), .ZN(n11203) );
  OR2_X1 U12128 ( .A1(n9907), .A2(n11203), .ZN(n9546) );
  INV_X1 U12129 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n11204) );
  OR2_X1 U12130 ( .A1(n6544), .A2(n11204), .ZN(n9545) );
  NAND2_X1 U12131 ( .A1(n6539), .A2(n9931), .ZN(n9555) );
  INV_X1 U12132 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9549) );
  NAND2_X1 U12133 ( .A1(n9550), .A2(n9549), .ZN(n9570) );
  NAND2_X1 U12134 ( .A1(n9570), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9551) );
  XNOR2_X1 U12135 ( .A(n9551), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10602) );
  AOI22_X1 U12136 ( .A1(n9799), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n9798), .B2(
        n10602), .ZN(n9553) );
  NAND2_X1 U12137 ( .A1(n10216), .A2(n12614), .ZN(n9552) );
  NAND2_X1 U12138 ( .A1(n9553), .A2(n9552), .ZN(n12459) );
  NAND2_X1 U12139 ( .A1(n12459), .A2(n9923), .ZN(n9554) );
  NAND2_X1 U12140 ( .A1(n9555), .A2(n9554), .ZN(n9556) );
  XNOR2_X1 U12141 ( .A(n9556), .B(n9743), .ZN(n11026) );
  NAND2_X1 U12142 ( .A1(n6539), .A2(n9936), .ZN(n9558) );
  NAND2_X1 U12143 ( .A1(n12459), .A2(n9931), .ZN(n9557) );
  AND2_X1 U12144 ( .A1(n9558), .A2(n9557), .ZN(n11025) );
  NAND2_X1 U12145 ( .A1(n11026), .A2(n11025), .ZN(n9559) );
  INV_X1 U12146 ( .A(n11026), .ZN(n9561) );
  INV_X1 U12147 ( .A(n11025), .ZN(n9560) );
  NAND2_X1 U12148 ( .A1(n9561), .A2(n9560), .ZN(n9562) );
  NAND2_X1 U12149 ( .A1(n12579), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9569) );
  INV_X1 U12150 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11355) );
  OR2_X1 U12151 ( .A1(n6545), .A2(n11355), .ZN(n9568) );
  INV_X1 U12152 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9563) );
  NAND2_X1 U12153 ( .A1(n9564), .A2(n9563), .ZN(n9565) );
  NAND2_X1 U12154 ( .A1(n9592), .A2(n9565), .ZN(n11354) );
  OR2_X1 U12155 ( .A1(n9594), .A2(n11354), .ZN(n9567) );
  INV_X1 U12156 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n15001) );
  OR2_X1 U12157 ( .A1(n9608), .A2(n15001), .ZN(n9566) );
  INV_X1 U12158 ( .A(n9570), .ZN(n9572) );
  INV_X1 U12159 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9571) );
  INV_X1 U12160 ( .A(n9586), .ZN(n9573) );
  NAND2_X1 U12161 ( .A1(n9573), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9574) );
  XNOR2_X1 U12162 ( .A(n9574), .B(P1_IR_REG_6__SCAN_IN), .ZN(n15007) );
  AOI22_X1 U12163 ( .A1(n9799), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9798), .B2(
        n15007), .ZN(n9576) );
  NAND2_X1 U12164 ( .A1(n10220), .A2(n12614), .ZN(n9575) );
  OR2_X1 U12165 ( .A1(n12417), .A2(n9954), .ZN(n9577) );
  OAI21_X1 U12166 ( .B1(n12418), .B2(n9677), .A(n9577), .ZN(n9578) );
  XNOR2_X1 U12167 ( .A(n9578), .B(n10789), .ZN(n9581) );
  OR2_X1 U12168 ( .A1(n12418), .A2(n9952), .ZN(n9580) );
  OR2_X1 U12169 ( .A1(n12417), .A2(n9677), .ZN(n9579) );
  NAND2_X1 U12170 ( .A1(n9580), .A2(n9579), .ZN(n9582) );
  INV_X1 U12171 ( .A(n9581), .ZN(n9584) );
  INV_X1 U12172 ( .A(n9582), .ZN(n9583) );
  NAND2_X1 U12173 ( .A1(n9584), .A2(n9583), .ZN(n11115) );
  NAND2_X1 U12174 ( .A1(n10222), .A2(n12614), .ZN(n9589) );
  INV_X1 U12175 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9585) );
  NAND2_X1 U12176 ( .A1(n9586), .A2(n9585), .ZN(n9604) );
  NAND2_X1 U12177 ( .A1(n9604), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9587) );
  XNOR2_X1 U12178 ( .A(n9587), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10768) );
  AOI22_X1 U12179 ( .A1(n9799), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9798), .B2(
        n10768), .ZN(n9588) );
  AND2_X2 U12180 ( .A1(n9589), .A2(n9588), .ZN(n12414) );
  NAND2_X1 U12181 ( .A1(n9987), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9599) );
  INV_X1 U12182 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9590) );
  OR2_X1 U12183 ( .A1(n9990), .A2(n9590), .ZN(n9598) );
  NAND2_X1 U12184 ( .A1(n9592), .A2(n9591), .ZN(n9593) );
  NAND2_X1 U12185 ( .A1(n9611), .A2(n9593), .ZN(n15697) );
  OR2_X1 U12186 ( .A1(n9594), .A2(n15697), .ZN(n9597) );
  INV_X1 U12187 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9595) );
  OR2_X1 U12188 ( .A1(n6545), .A2(n9595), .ZN(n9596) );
  AND4_X2 U12189 ( .A1(n9599), .A2(n9598), .A3(n9597), .A4(n9596), .ZN(n12415)
         );
  OAI22_X1 U12190 ( .A1(n12414), .A2(n9954), .B1(n12415), .B2(n9677), .ZN(
        n9600) );
  XNOR2_X1 U12191 ( .A(n9600), .B(n10789), .ZN(n9602) );
  OAI22_X1 U12192 ( .A1(n12414), .A2(n9677), .B1(n12415), .B2(n9952), .ZN(
        n9601) );
  XNOR2_X1 U12193 ( .A(n9602), .B(n9601), .ZN(n12002) );
  NAND2_X1 U12194 ( .A1(n9602), .A2(n9601), .ZN(n9603) );
  NAND2_X1 U12195 ( .A1(n10489), .A2(n12614), .ZN(n9607) );
  NAND2_X1 U12196 ( .A1(n9625), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9605) );
  XNOR2_X1 U12197 ( .A(n9605), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10771) );
  AOI22_X1 U12198 ( .A1(n9799), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9798), .B2(
        n10771), .ZN(n9606) );
  NAND2_X1 U12199 ( .A1(n15684), .A2(n9923), .ZN(n9618) );
  NAND2_X1 U12200 ( .A1(n12584), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n9616) );
  INV_X1 U12201 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9609) );
  OR2_X1 U12202 ( .A1(n9927), .A2(n9609), .ZN(n9615) );
  NAND2_X1 U12203 ( .A1(n9611), .A2(n9610), .ZN(n9612) );
  NAND2_X1 U12204 ( .A1(n9646), .A2(n9612), .ZN(n15681) );
  OR2_X1 U12205 ( .A1(n9594), .A2(n15681), .ZN(n9614) );
  INV_X1 U12206 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n15682) );
  OR2_X1 U12207 ( .A1(n6544), .A2(n15682), .ZN(n9613) );
  NAND2_X1 U12208 ( .A1(n14954), .A2(n9931), .ZN(n9617) );
  NAND2_X1 U12209 ( .A1(n9618), .A2(n9617), .ZN(n9619) );
  XNOR2_X1 U12210 ( .A(n9619), .B(n9743), .ZN(n9623) );
  AND2_X1 U12211 ( .A1(n14954), .A2(n9936), .ZN(n9620) );
  AOI21_X1 U12212 ( .B1(n15684), .B2(n9931), .A(n9620), .ZN(n9622) );
  XNOR2_X1 U12213 ( .A(n9623), .B(n9622), .ZN(n11865) );
  NAND2_X1 U12214 ( .A1(n9623), .A2(n9622), .ZN(n9624) );
  NAND2_X1 U12215 ( .A1(n11868), .A2(n9624), .ZN(n14770) );
  NAND2_X1 U12216 ( .A1(n10572), .A2(n12614), .ZN(n9629) );
  NAND2_X1 U12217 ( .A1(n9626), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9644) );
  NAND2_X1 U12218 ( .A1(n9644), .A2(n9643), .ZN(n9642) );
  NAND2_X1 U12219 ( .A1(n9642), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9627) );
  AOI22_X1 U12220 ( .A1(n15037), .A2(n9798), .B1(n9799), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n9628) );
  NAND2_X1 U12221 ( .A1(n14778), .A2(n9923), .ZN(n9638) );
  NAND2_X1 U12222 ( .A1(n9987), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9636) );
  INV_X1 U12223 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9630) );
  OR2_X1 U12224 ( .A1(n9990), .A2(n9630), .ZN(n9635) );
  INV_X1 U12225 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9631) );
  NAND2_X1 U12226 ( .A1(n9648), .A2(n9631), .ZN(n9632) );
  NAND2_X1 U12227 ( .A1(n9671), .A2(n9632), .ZN(n14783) );
  OR2_X1 U12228 ( .A1(n9907), .A2(n14783), .ZN(n9634) );
  INV_X1 U12229 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n12210) );
  OR2_X1 U12230 ( .A1(n6545), .A2(n12210), .ZN(n9633) );
  NAND4_X1 U12231 ( .A1(n9636), .A2(n9635), .A3(n9634), .A4(n9633), .ZN(n14952) );
  NAND2_X1 U12232 ( .A1(n14952), .A2(n9931), .ZN(n9637) );
  NAND2_X1 U12233 ( .A1(n9638), .A2(n9637), .ZN(n9639) );
  XNOR2_X1 U12234 ( .A(n9639), .B(n9914), .ZN(n14775) );
  NAND2_X1 U12235 ( .A1(n14778), .A2(n9931), .ZN(n9641) );
  NAND2_X1 U12236 ( .A1(n14952), .A2(n9936), .ZN(n9640) );
  NAND2_X1 U12237 ( .A1(n9641), .A2(n9640), .ZN(n9660) );
  OAI21_X1 U12238 ( .B1(n9644), .B2(n9643), .A(n9642), .ZN(n10773) );
  INV_X1 U12239 ( .A(n10773), .ZN(n10917) );
  AOI22_X1 U12240 ( .A1(n10917), .A2(n9798), .B1(n9799), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n9645) );
  NAND2_X1 U12241 ( .A1(n12475), .A2(n9931), .ZN(n9654) );
  NAND2_X1 U12242 ( .A1(n12583), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9652) );
  INV_X1 U12243 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10763) );
  OR2_X1 U12244 ( .A1(n9927), .A2(n10763), .ZN(n9651) );
  INV_X1 U12245 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10289) );
  OR2_X1 U12246 ( .A1(n9990), .A2(n10289), .ZN(n9650) );
  NAND2_X1 U12247 ( .A1(n9646), .A2(n10766), .ZN(n9647) );
  NAND2_X1 U12248 ( .A1(n9648), .A2(n9647), .ZN(n14856) );
  OR2_X1 U12249 ( .A1(n9907), .A2(n14856), .ZN(n9649) );
  NAND4_X1 U12250 ( .A1(n9652), .A2(n9651), .A3(n9650), .A4(n9649), .ZN(n14953) );
  NAND2_X1 U12251 ( .A1(n14953), .A2(n9936), .ZN(n9653) );
  NAND2_X1 U12252 ( .A1(n9654), .A2(n9653), .ZN(n14771) );
  NAND2_X1 U12253 ( .A1(n12475), .A2(n9923), .ZN(n9656) );
  NAND2_X1 U12254 ( .A1(n14953), .A2(n9931), .ZN(n9655) );
  NAND2_X1 U12255 ( .A1(n9656), .A2(n9655), .ZN(n9657) );
  XNOR2_X1 U12256 ( .A(n9657), .B(n10789), .ZN(n14851) );
  AOI22_X1 U12257 ( .A1(n14775), .A2(n9660), .B1(n14771), .B2(n14851), .ZN(
        n9658) );
  NAND2_X1 U12258 ( .A1(n14770), .A2(n9658), .ZN(n9666) );
  INV_X1 U12259 ( .A(n14851), .ZN(n14773) );
  INV_X1 U12260 ( .A(n14771), .ZN(n14772) );
  AND2_X1 U12261 ( .A1(n14773), .A2(n14772), .ZN(n9662) );
  INV_X1 U12262 ( .A(n9662), .ZN(n9659) );
  INV_X1 U12263 ( .A(n9660), .ZN(n14774) );
  INV_X1 U12264 ( .A(n14775), .ZN(n9661) );
  OAI21_X1 U12265 ( .B1(n9662), .B2(n14774), .A(n9661), .ZN(n9663) );
  NAND2_X1 U12266 ( .A1(n10613), .A2(n12614), .ZN(n9670) );
  NAND2_X1 U12267 ( .A1(n9667), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9668) );
  XNOR2_X1 U12268 ( .A(n9668), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11441) );
  AOI22_X1 U12269 ( .A1(n9799), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9798), 
        .B2(n11441), .ZN(n9669) );
  INV_X1 U12270 ( .A(n14891), .ZN(n12486) );
  NAND2_X1 U12271 ( .A1(n9987), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n9676) );
  INV_X1 U12272 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10427) );
  OR2_X1 U12273 ( .A1(n9990), .A2(n10427), .ZN(n9675) );
  NAND2_X1 U12274 ( .A1(n9671), .A2(n10915), .ZN(n9672) );
  NAND2_X1 U12275 ( .A1(n9692), .A2(n9672), .ZN(n14895) );
  OR2_X1 U12276 ( .A1(n9907), .A2(n14895), .ZN(n9674) );
  INV_X1 U12277 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11955) );
  OR2_X1 U12278 ( .A1(n6544), .A2(n11955), .ZN(n9673) );
  NAND4_X1 U12279 ( .A1(n9676), .A2(n9675), .A3(n9674), .A4(n9673), .ZN(n14951) );
  INV_X1 U12280 ( .A(n14951), .ZN(n12487) );
  OAI22_X1 U12281 ( .A1(n12486), .A2(n9677), .B1(n12487), .B2(n9952), .ZN(
        n9682) );
  NAND2_X1 U12282 ( .A1(n14891), .A2(n9923), .ZN(n9679) );
  NAND2_X1 U12283 ( .A1(n14951), .A2(n9931), .ZN(n9678) );
  NAND2_X1 U12284 ( .A1(n9679), .A2(n9678), .ZN(n9680) );
  XNOR2_X1 U12285 ( .A(n9680), .B(n9914), .ZN(n9681) );
  XOR2_X1 U12286 ( .A(n9682), .B(n9681), .Z(n14892) );
  INV_X1 U12287 ( .A(n9681), .ZN(n9684) );
  INV_X1 U12288 ( .A(n9682), .ZN(n9683) );
  NAND2_X1 U12289 ( .A1(n10678), .A2(n12614), .ZN(n9689) );
  NAND2_X1 U12290 ( .A1(n9685), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9686) );
  MUX2_X1 U12291 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9686), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n9687) );
  AOI22_X1 U12292 ( .A1(n9799), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n9798), 
        .B2(n11471), .ZN(n9688) );
  NAND2_X1 U12293 ( .A1(n12579), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9699) );
  INV_X1 U12294 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9690) );
  OR2_X1 U12295 ( .A1(n9927), .A2(n9690), .ZN(n9698) );
  INV_X1 U12296 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9691) );
  NAND2_X1 U12297 ( .A1(n9692), .A2(n9691), .ZN(n9693) );
  NAND2_X1 U12298 ( .A1(n9694), .A2(n9693), .ZN(n12028) );
  OR2_X1 U12299 ( .A1(n9907), .A2(n12028), .ZN(n9697) );
  INV_X1 U12300 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9695) );
  OR2_X1 U12301 ( .A1(n6545), .A2(n9695), .ZN(n9696) );
  OAI22_X1 U12302 ( .A1(n7298), .A2(n9677), .B1(n14873), .B2(n9952), .ZN(n9702) );
  OAI22_X1 U12303 ( .A1(n7298), .A2(n9954), .B1(n14873), .B2(n9677), .ZN(n9700) );
  XNOR2_X1 U12304 ( .A(n9700), .B(n10789), .ZN(n9701) );
  XOR2_X1 U12305 ( .A(n9702), .B(n9701), .Z(n14807) );
  NAND2_X1 U12306 ( .A1(n9701), .A2(n9702), .ZN(n9703) );
  XNOR2_X1 U12307 ( .A(n9705), .B(n9704), .ZN(n14872) );
  NAND2_X1 U12308 ( .A1(n10784), .A2(n12614), .ZN(n9711) );
  NAND2_X1 U12309 ( .A1(n9724), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9709) );
  XNOR2_X1 U12310 ( .A(n9709), .B(P1_IR_REG_14__SCAN_IN), .ZN(n15050) );
  AOI22_X1 U12311 ( .A1(n9799), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n9798), 
        .B2(n15050), .ZN(n9710) );
  NAND2_X2 U12312 ( .A1(n9711), .A2(n9710), .ZN(n15486) );
  XNOR2_X1 U12313 ( .A(n9735), .B(P1_REG3_REG_14__SCAN_IN), .ZN(n14752) );
  NAND2_X1 U12314 ( .A1(n9986), .A2(n14752), .ZN(n9716) );
  INV_X1 U12315 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9712) );
  OR2_X1 U12316 ( .A1(n9990), .A2(n9712), .ZN(n9715) );
  INV_X1 U12317 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n15043) );
  OR2_X1 U12318 ( .A1(n9927), .A2(n15043), .ZN(n9714) );
  INV_X1 U12319 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n15349) );
  OR2_X1 U12320 ( .A1(n6545), .A2(n15349), .ZN(n9713) );
  INV_X1 U12321 ( .A(n14923), .ZN(n14948) );
  AOI22_X1 U12322 ( .A1(n15486), .A2(n9931), .B1(n9936), .B2(n14948), .ZN(
        n9720) );
  NAND2_X1 U12323 ( .A1(n15486), .A2(n9923), .ZN(n9718) );
  OR2_X1 U12324 ( .A1(n14923), .A2(n9677), .ZN(n9717) );
  NAND2_X1 U12325 ( .A1(n9718), .A2(n9717), .ZN(n9719) );
  XNOR2_X1 U12326 ( .A(n9719), .B(n9914), .ZN(n9722) );
  XOR2_X1 U12327 ( .A(n9720), .B(n9722), .Z(n14751) );
  INV_X1 U12328 ( .A(n9720), .ZN(n9721) );
  INV_X1 U12329 ( .A(n9724), .ZN(n9726) );
  INV_X1 U12330 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9725) );
  NAND2_X1 U12331 ( .A1(n9726), .A2(n9725), .ZN(n9728) );
  NAND2_X1 U12332 ( .A1(n9728), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9727) );
  MUX2_X1 U12333 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9727), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n9731) );
  INV_X1 U12334 ( .A(n9728), .ZN(n9730) );
  INV_X1 U12335 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9729) );
  NAND2_X1 U12336 ( .A1(n9730), .A2(n9729), .ZN(n9765) );
  AOI22_X1 U12337 ( .A1(n15053), .A2(n9798), .B1(n9799), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n9732) );
  NAND2_X1 U12338 ( .A1(n15479), .A2(n9923), .ZN(n9742) );
  INV_X1 U12339 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n11480) );
  INV_X1 U12340 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9734) );
  OAI21_X1 U12341 ( .B1(n9735), .B2(n11480), .A(n9734), .ZN(n9736) );
  AND2_X1 U12342 ( .A1(n9736), .A2(n9749), .ZN(n15331) );
  NAND2_X1 U12343 ( .A1(n15331), .A2(n9986), .ZN(n9740) );
  INV_X1 U12344 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10300) );
  OR2_X1 U12345 ( .A1(n9927), .A2(n10300), .ZN(n9739) );
  NAND2_X1 U12346 ( .A1(n12579), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n9738) );
  NAND2_X1 U12347 ( .A1(n12583), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n9737) );
  OR2_X1 U12348 ( .A1(n14830), .A2(n9677), .ZN(n9741) );
  NAND2_X1 U12349 ( .A1(n9742), .A2(n9741), .ZN(n9744) );
  XNOR2_X1 U12350 ( .A(n9744), .B(n9743), .ZN(n14825) );
  INV_X1 U12351 ( .A(n14825), .ZN(n9761) );
  NOR2_X1 U12352 ( .A1(n14830), .A2(n9952), .ZN(n9745) );
  AOI21_X1 U12353 ( .B1(n15479), .B2(n9931), .A(n9745), .ZN(n9759) );
  INV_X1 U12354 ( .A(n9759), .ZN(n14920) );
  NAND2_X1 U12355 ( .A1(n10708), .A2(n12614), .ZN(n9748) );
  NAND2_X1 U12356 ( .A1(n9765), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9746) );
  XNOR2_X1 U12357 ( .A(n9746), .B(P1_IR_REG_16__SCAN_IN), .ZN(n15070) );
  AOI22_X1 U12358 ( .A1(n15070), .A2(n9798), .B1(n9799), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n9747) );
  NAND2_X2 U12359 ( .A1(n9748), .A2(n9747), .ZN(n15472) );
  INV_X1 U12360 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n15316) );
  INV_X1 U12361 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n10258) );
  NAND2_X1 U12362 ( .A1(n9749), .A2(n10258), .ZN(n9750) );
  NAND2_X1 U12363 ( .A1(n9787), .A2(n9750), .ZN(n15315) );
  OR2_X1 U12364 ( .A1(n15315), .A2(n9907), .ZN(n9754) );
  NAND2_X1 U12365 ( .A1(n9987), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9752) );
  NAND2_X1 U12366 ( .A1(n12579), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n9751) );
  AND2_X1 U12367 ( .A1(n9752), .A2(n9751), .ZN(n9753) );
  OAI211_X1 U12368 ( .C1(n6544), .C2(n15316), .A(n9754), .B(n9753), .ZN(n14947) );
  AOI22_X1 U12369 ( .A1(n15472), .A2(n9931), .B1(n6543), .B2(n14947), .ZN(
        n14826) );
  INV_X1 U12370 ( .A(n14826), .ZN(n9758) );
  NAND2_X1 U12371 ( .A1(n15472), .A2(n9923), .ZN(n9756) );
  NAND2_X1 U12372 ( .A1(n14947), .A2(n9931), .ZN(n9755) );
  NAND2_X1 U12373 ( .A1(n9756), .A2(n9755), .ZN(n9757) );
  XNOR2_X1 U12374 ( .A(n9757), .B(n9914), .ZN(n14827) );
  AOI22_X1 U12375 ( .A1(n9761), .A2(n14920), .B1(n9758), .B2(n14827), .ZN(
        n9764) );
  AOI21_X1 U12376 ( .B1(n14825), .B2(n9759), .A(n14826), .ZN(n9762) );
  NAND2_X1 U12377 ( .A1(n9759), .A2(n14826), .ZN(n9760) );
  OAI22_X1 U12378 ( .A1(n9762), .A2(n14827), .B1(n9761), .B2(n9760), .ZN(n9763) );
  NAND2_X1 U12379 ( .A1(n10758), .A2(n12614), .ZN(n9768) );
  NAND2_X1 U12380 ( .A1(n9780), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9766) );
  XNOR2_X1 U12381 ( .A(n9766), .B(P1_IR_REG_17__SCAN_IN), .ZN(n15086) );
  AOI22_X1 U12382 ( .A1(n15086), .A2(n9798), .B1(n9799), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n9767) );
  XNOR2_X1 U12383 ( .A(n9787), .B(P1_REG3_REG_17__SCAN_IN), .ZN(n15300) );
  NAND2_X1 U12384 ( .A1(n15300), .A2(n9986), .ZN(n9773) );
  INV_X1 U12385 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n15079) );
  NAND2_X1 U12386 ( .A1(n12579), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n9770) );
  NAND2_X1 U12387 ( .A1(n12583), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9769) );
  OAI211_X1 U12388 ( .C1(n9927), .C2(n15079), .A(n9770), .B(n9769), .ZN(n9771)
         );
  INV_X1 U12389 ( .A(n9771), .ZN(n9772) );
  OAI22_X1 U12390 ( .A1(n15466), .A2(n9954), .B1(n14831), .B2(n9677), .ZN(
        n9774) );
  XNOR2_X1 U12391 ( .A(n9774), .B(n9914), .ZN(n9778) );
  OR2_X1 U12392 ( .A1(n15466), .A2(n9677), .ZN(n9776) );
  NAND2_X1 U12393 ( .A1(n14946), .A2(n9936), .ZN(n9775) );
  NAND2_X1 U12394 ( .A1(n9776), .A2(n9775), .ZN(n9777) );
  XNOR2_X1 U12395 ( .A(n9778), .B(n9777), .ZN(n14837) );
  OR2_X1 U12396 ( .A1(n10892), .A2(n9779), .ZN(n9784) );
  OAI21_X1 U12397 ( .B1(n9780), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9781) );
  XNOR2_X1 U12398 ( .A(n9781), .B(P1_IR_REG_18__SCAN_IN), .ZN(n15089) );
  NOR2_X1 U12399 ( .A1(n12615), .A2(n10890), .ZN(n9782) );
  AOI21_X1 U12400 ( .B1(n15089), .B2(n9798), .A(n9782), .ZN(n9783) );
  NAND2_X2 U12401 ( .A1(n9784), .A2(n9783), .ZN(n15461) );
  NAND2_X1 U12402 ( .A1(n15461), .A2(n9923), .ZN(n9793) );
  INV_X1 U12403 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9786) );
  INV_X1 U12404 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9785) );
  OAI21_X1 U12405 ( .B1(n9787), .B2(n9786), .A(n9785), .ZN(n9788) );
  AND2_X1 U12406 ( .A1(n9788), .A2(n9802), .ZN(n15287) );
  NAND2_X1 U12407 ( .A1(n15287), .A2(n9986), .ZN(n9791) );
  AOI22_X1 U12408 ( .A1(n9987), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n12584), 
        .B2(P1_REG0_REG_18__SCAN_IN), .ZN(n9790) );
  INV_X1 U12409 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n15092) );
  OR2_X1 U12410 ( .A1(n6544), .A2(n15092), .ZN(n9789) );
  OR2_X1 U12411 ( .A1(n14838), .A2(n9677), .ZN(n9792) );
  NAND2_X1 U12412 ( .A1(n9793), .A2(n9792), .ZN(n9794) );
  XNOR2_X1 U12413 ( .A(n9794), .B(n10789), .ZN(n9795) );
  AOI22_X1 U12414 ( .A1(n15461), .A2(n9931), .B1(n9936), .B2(n14945), .ZN(
        n9796) );
  XNOR2_X1 U12415 ( .A(n9795), .B(n9796), .ZN(n14902) );
  INV_X1 U12416 ( .A(n9795), .ZN(n9797) );
  NAND2_X1 U12417 ( .A1(n10983), .A2(n12614), .ZN(n9801) );
  AOI22_X1 U12418 ( .A1(n9799), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n15112), 
        .B2(n9798), .ZN(n9800) );
  NAND2_X1 U12419 ( .A1(n15455), .A2(n9923), .ZN(n9812) );
  INV_X1 U12420 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n10448) );
  NAND2_X1 U12421 ( .A1(n9802), .A2(n10448), .ZN(n9803) );
  NAND2_X1 U12422 ( .A1(n9804), .A2(n9803), .ZN(n15271) );
  OR2_X1 U12423 ( .A1(n15271), .A2(n9907), .ZN(n9810) );
  INV_X1 U12424 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9807) );
  NAND2_X1 U12425 ( .A1(n12583), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n9806) );
  NAND2_X1 U12426 ( .A1(n12579), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9805) );
  OAI211_X1 U12427 ( .C1(n9927), .C2(n9807), .A(n9806), .B(n9805), .ZN(n9808)
         );
  INV_X1 U12428 ( .A(n9808), .ZN(n9809) );
  NAND2_X1 U12429 ( .A1(n14944), .A2(n9931), .ZN(n9811) );
  NAND2_X1 U12430 ( .A1(n9812), .A2(n9811), .ZN(n9813) );
  XNOR2_X1 U12431 ( .A(n9813), .B(n10789), .ZN(n9815) );
  AND2_X1 U12432 ( .A1(n14944), .A2(n9936), .ZN(n9814) );
  AOI21_X1 U12433 ( .B1(n15455), .B2(n9931), .A(n9814), .ZN(n9816) );
  XNOR2_X1 U12434 ( .A(n9815), .B(n9816), .ZN(n14788) );
  XNOR2_X1 U12435 ( .A(n9819), .B(n9818), .ZN(n14863) );
  NAND2_X1 U12436 ( .A1(n11109), .A2(n12614), .ZN(n9822) );
  OR2_X1 U12437 ( .A1(n12615), .A2(n11113), .ZN(n9821) );
  NAND2_X1 U12438 ( .A1(n9823), .A2(n14801), .ZN(n9824) );
  NAND2_X1 U12439 ( .A1(n9835), .A2(n9824), .ZN(n15229) );
  INV_X1 U12440 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10353) );
  NAND2_X1 U12441 ( .A1(n12579), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9826) );
  NAND2_X1 U12442 ( .A1(n12583), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9825) );
  OAI211_X1 U12443 ( .C1(n9927), .C2(n10353), .A(n9826), .B(n9825), .ZN(n9827)
         );
  INV_X1 U12444 ( .A(n9827), .ZN(n9828) );
  OAI22_X1 U12445 ( .A1(n14805), .A2(n9677), .B1(n13060), .B2(n9952), .ZN(
        n9830) );
  OAI22_X1 U12446 ( .A1(n14805), .A2(n9954), .B1(n13060), .B2(n9677), .ZN(
        n9829) );
  XNOR2_X1 U12447 ( .A(n9829), .B(n10789), .ZN(n9831) );
  XOR2_X1 U12448 ( .A(n9830), .B(n9831), .Z(n14797) );
  OR2_X1 U12449 ( .A1(n9833), .A2(n10481), .ZN(n9834) );
  XNOR2_X1 U12450 ( .A(n9834), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15552) );
  NAND2_X1 U12451 ( .A1(n9835), .A2(n14886), .ZN(n9836) );
  AND2_X1 U12452 ( .A1(n9852), .A2(n9836), .ZN(n15220) );
  NAND2_X1 U12453 ( .A1(n15220), .A2(n9986), .ZN(n9841) );
  INV_X1 U12454 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n10460) );
  NAND2_X1 U12455 ( .A1(n12583), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9838) );
  NAND2_X1 U12456 ( .A1(n9987), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n9837) );
  OAI211_X1 U12457 ( .C1(n9990), .C2(n10460), .A(n9838), .B(n9837), .ZN(n9839)
         );
  INV_X1 U12458 ( .A(n9839), .ZN(n9840) );
  INV_X1 U12459 ( .A(n14941), .ZN(n13063) );
  OAI22_X1 U12460 ( .A1(n15223), .A2(n9677), .B1(n13063), .B2(n9952), .ZN(
        n9846) );
  NAND2_X1 U12461 ( .A1(n15437), .A2(n9923), .ZN(n9843) );
  NAND2_X1 U12462 ( .A1(n14941), .A2(n9931), .ZN(n9842) );
  NAND2_X1 U12463 ( .A1(n9843), .A2(n9842), .ZN(n9844) );
  XNOR2_X1 U12464 ( .A(n9844), .B(n9914), .ZN(n9845) );
  XOR2_X1 U12465 ( .A(n9846), .B(n9845), .Z(n14882) );
  INV_X1 U12466 ( .A(n9845), .ZN(n9848) );
  INV_X1 U12467 ( .A(n9846), .ZN(n9847) );
  NAND2_X1 U12468 ( .A1(n9848), .A2(n9847), .ZN(n14761) );
  NAND2_X1 U12469 ( .A1(n11458), .A2(n12614), .ZN(n9850) );
  OR2_X1 U12470 ( .A1(n12615), .A2(n11460), .ZN(n9849) );
  NAND2_X1 U12471 ( .A1(n15428), .A2(n9923), .ZN(n9861) );
  INV_X1 U12472 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9851) );
  NAND2_X1 U12473 ( .A1(n9852), .A2(n9851), .ZN(n9853) );
  NAND2_X1 U12474 ( .A1(n9890), .A2(n9853), .ZN(n14765) );
  INV_X1 U12475 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9856) );
  NAND2_X1 U12476 ( .A1(n12579), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9855) );
  NAND2_X1 U12477 ( .A1(n12583), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9854) );
  OAI211_X1 U12478 ( .C1(n9856), .C2(n9927), .A(n9855), .B(n9854), .ZN(n9857)
         );
  INV_X1 U12479 ( .A(n9857), .ZN(n9858) );
  NAND2_X1 U12480 ( .A1(n14940), .A2(n9931), .ZN(n9860) );
  NAND2_X1 U12481 ( .A1(n9861), .A2(n9860), .ZN(n9862) );
  XNOR2_X1 U12482 ( .A(n9862), .B(n10789), .ZN(n9866) );
  INV_X1 U12483 ( .A(n9866), .ZN(n9863) );
  AOI22_X1 U12484 ( .A1(n15428), .A2(n9931), .B1(n9936), .B2(n14940), .ZN(
        n9865) );
  NAND2_X1 U12485 ( .A1(n9863), .A2(n9865), .ZN(n9864) );
  AND2_X1 U12486 ( .A1(n14761), .A2(n9864), .ZN(n9868) );
  INV_X1 U12487 ( .A(n9864), .ZN(n9867) );
  XNOR2_X1 U12488 ( .A(n9866), .B(n9865), .ZN(n14763) );
  NAND2_X1 U12489 ( .A1(n11769), .A2(n12614), .ZN(n9870) );
  OR2_X1 U12490 ( .A1(n12615), .A2(n11772), .ZN(n9869) );
  NAND2_X1 U12491 ( .A1(n15425), .A2(n9923), .ZN(n9878) );
  XNOR2_X1 U12492 ( .A(n9890), .B(P1_REG3_REG_24__SCAN_IN), .ZN(n15192) );
  NAND2_X1 U12493 ( .A1(n15192), .A2(n9986), .ZN(n9876) );
  INV_X1 U12494 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9873) );
  NAND2_X1 U12495 ( .A1(n12579), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9872) );
  NAND2_X1 U12496 ( .A1(n12583), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9871) );
  OAI211_X1 U12497 ( .C1(n9927), .C2(n9873), .A(n9872), .B(n9871), .ZN(n9874)
         );
  INV_X1 U12498 ( .A(n9874), .ZN(n9875) );
  NAND2_X1 U12499 ( .A1(n14939), .A2(n9931), .ZN(n9877) );
  NAND2_X1 U12500 ( .A1(n9878), .A2(n9877), .ZN(n9879) );
  XNOR2_X1 U12501 ( .A(n9879), .B(n9914), .ZN(n9880) );
  AOI22_X1 U12502 ( .A1(n15425), .A2(n9931), .B1(n6543), .B2(n14939), .ZN(
        n9881) );
  XNOR2_X1 U12503 ( .A(n9880), .B(n9881), .ZN(n14846) );
  INV_X1 U12504 ( .A(n9880), .ZN(n9882) );
  NAND2_X1 U12505 ( .A1(n9882), .A2(n9881), .ZN(n9883) );
  NAND2_X1 U12506 ( .A1(n12098), .A2(n12614), .ZN(n9886) );
  INV_X1 U12507 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12099) );
  OR2_X1 U12508 ( .A1(n12615), .A2(n12099), .ZN(n9885) );
  INV_X1 U12509 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9888) );
  INV_X1 U12510 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9887) );
  OAI21_X1 U12511 ( .B1(n9890), .B2(n9888), .A(n9887), .ZN(n9891) );
  NAND2_X1 U12512 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .ZN(n9889) );
  NAND2_X1 U12513 ( .A1(n15174), .A2(n9986), .ZN(n9897) );
  INV_X1 U12514 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9894) );
  NAND2_X1 U12515 ( .A1(n12579), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n9893) );
  NAND2_X1 U12516 ( .A1(n12583), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n9892) );
  OAI211_X1 U12517 ( .C1(n9927), .C2(n9894), .A(n9893), .B(n9892), .ZN(n9895)
         );
  INV_X1 U12518 ( .A(n9895), .ZN(n9896) );
  INV_X1 U12519 ( .A(n14938), .ZN(n14912) );
  OAI22_X1 U12520 ( .A1(n15417), .A2(n9677), .B1(n14912), .B2(n9952), .ZN(
        n9901) );
  NAND2_X1 U12521 ( .A1(n14822), .A2(n9923), .ZN(n9899) );
  NAND2_X1 U12522 ( .A1(n14938), .A2(n9931), .ZN(n9898) );
  NAND2_X1 U12523 ( .A1(n9899), .A2(n9898), .ZN(n9900) );
  XNOR2_X1 U12524 ( .A(n9900), .B(n9914), .ZN(n9902) );
  XOR2_X1 U12525 ( .A(n9901), .B(n9902), .Z(n14817) );
  NAND2_X1 U12526 ( .A1(n12218), .A2(n12614), .ZN(n9904) );
  OR2_X1 U12527 ( .A1(n12615), .A2(n12219), .ZN(n9903) );
  NAND2_X1 U12528 ( .A1(n15163), .A2(n9923), .ZN(n9913) );
  INV_X1 U12529 ( .A(n6615), .ZN(n9905) );
  INV_X1 U12530 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14915) );
  NAND2_X1 U12531 ( .A1(n6615), .A2(n14915), .ZN(n9906) );
  NAND2_X1 U12532 ( .A1(n9944), .A2(n9906), .ZN(n15161) );
  INV_X1 U12533 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10279) );
  NAND2_X1 U12534 ( .A1(n12579), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9909) );
  NAND2_X1 U12535 ( .A1(n12583), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9908) );
  OAI211_X1 U12536 ( .C1(n10279), .C2(n9927), .A(n9909), .B(n9908), .ZN(n9910)
         );
  INV_X1 U12537 ( .A(n9910), .ZN(n9911) );
  NAND2_X1 U12538 ( .A1(n14937), .A2(n9931), .ZN(n9912) );
  NAND2_X1 U12539 ( .A1(n9913), .A2(n9912), .ZN(n9915) );
  XNOR2_X1 U12540 ( .A(n9915), .B(n9914), .ZN(n9916) );
  OAI22_X1 U12541 ( .A1(n15410), .A2(n9677), .B1(n13069), .B2(n9952), .ZN(
        n9917) );
  XNOR2_X1 U12542 ( .A(n9916), .B(n9917), .ZN(n14908) );
  INV_X1 U12543 ( .A(n9916), .ZN(n9919) );
  INV_X1 U12544 ( .A(n9917), .ZN(n9918) );
  NAND2_X1 U12545 ( .A1(n9919), .A2(n9918), .ZN(n9920) );
  NAND2_X1 U12546 ( .A1(n12267), .A2(n12614), .ZN(n9922) );
  INV_X1 U12547 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n12282) );
  OR2_X1 U12548 ( .A1(n12615), .A2(n12282), .ZN(n9921) );
  NAND2_X1 U12549 ( .A1(n15150), .A2(n9923), .ZN(n9933) );
  XNOR2_X1 U12550 ( .A(n9944), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n15149) );
  NAND2_X1 U12551 ( .A1(n15149), .A2(n9986), .ZN(n9930) );
  INV_X1 U12552 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9926) );
  NAND2_X1 U12553 ( .A1(n12583), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9925) );
  NAND2_X1 U12554 ( .A1(n12579), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n9924) );
  OAI211_X1 U12555 ( .C1(n9927), .C2(n9926), .A(n9925), .B(n9924), .ZN(n9928)
         );
  INV_X1 U12556 ( .A(n9928), .ZN(n9929) );
  NAND2_X1 U12557 ( .A1(n14936), .A2(n9931), .ZN(n9932) );
  NAND2_X1 U12558 ( .A1(n9933), .A2(n9932), .ZN(n9935) );
  XNOR2_X1 U12559 ( .A(n9935), .B(n9934), .ZN(n9982) );
  AND2_X1 U12560 ( .A1(n14936), .A2(n9936), .ZN(n9937) );
  AOI21_X1 U12561 ( .B1(n15150), .B2(n9931), .A(n9937), .ZN(n9981) );
  XNOR2_X1 U12562 ( .A(n9982), .B(n9981), .ZN(n14743) );
  INV_X1 U12563 ( .A(n14743), .ZN(n9938) );
  INV_X1 U12564 ( .A(n9983), .ZN(n9980) );
  NAND2_X1 U12565 ( .A1(n13184), .A2(n12614), .ZN(n9940) );
  OR2_X1 U12566 ( .A1(n12615), .A2(n13185), .ZN(n9939) );
  INV_X1 U12567 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9942) );
  INV_X1 U12568 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9941) );
  OAI21_X1 U12569 ( .B1(n9944), .B2(n9942), .A(n9941), .ZN(n9945) );
  NAND2_X1 U12570 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n9943) );
  NAND2_X1 U12571 ( .A1(n15132), .A2(n9986), .ZN(n9951) );
  INV_X1 U12572 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9948) );
  NAND2_X1 U12573 ( .A1(n12583), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9947) );
  NAND2_X1 U12574 ( .A1(n12584), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n9946) );
  OAI211_X1 U12575 ( .C1(n9927), .C2(n9948), .A(n9947), .B(n9946), .ZN(n9949)
         );
  INV_X1 U12576 ( .A(n9949), .ZN(n9950) );
  OAI22_X1 U12577 ( .A1(n15400), .A2(n9677), .B1(n13025), .B2(n9952), .ZN(
        n9953) );
  XNOR2_X1 U12578 ( .A(n9953), .B(n10789), .ZN(n9956) );
  OAI22_X1 U12579 ( .A1(n15400), .A2(n9954), .B1(n13025), .B2(n9677), .ZN(
        n9955) );
  XNOR2_X1 U12580 ( .A(n9956), .B(n9955), .ZN(n10005) );
  INV_X1 U12581 ( .A(n10005), .ZN(n9979) );
  INV_X1 U12582 ( .A(P1_B_REG_SCAN_IN), .ZN(n13033) );
  NAND2_X1 U12583 ( .A1(n9959), .A2(n13033), .ZN(n9958) );
  INV_X1 U12584 ( .A(n9973), .ZN(n12100) );
  NAND3_X1 U12585 ( .A1(n12100), .A2(P1_B_REG_SCAN_IN), .A3(n11774), .ZN(n9960) );
  INV_X1 U12586 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10230) );
  NAND2_X1 U12587 ( .A1(n10797), .A2(n10230), .ZN(n9962) );
  INV_X1 U12588 ( .A(n9957), .ZN(n12220) );
  NAND2_X1 U12589 ( .A1(n12220), .A2(n11774), .ZN(n10227) );
  INV_X1 U12590 ( .A(n11059), .ZN(n15518) );
  NOR4_X1 U12591 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n9966) );
  NOR4_X1 U12592 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n9965) );
  NOR4_X1 U12593 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9964) );
  NOR4_X1 U12594 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n9963) );
  AND4_X1 U12595 ( .A1(n9966), .A2(n9965), .A3(n9964), .A4(n9963), .ZN(n9972)
         );
  NOR2_X1 U12596 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n9970) );
  NOR4_X1 U12597 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n9969) );
  NOR4_X1 U12598 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n9968) );
  NOR4_X1 U12599 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n9967) );
  AND4_X1 U12600 ( .A1(n9970), .A2(n9969), .A3(n9968), .A4(n9967), .ZN(n9971)
         );
  NAND2_X1 U12601 ( .A1(n9972), .A2(n9971), .ZN(n10796) );
  INV_X1 U12602 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10226) );
  OR2_X1 U12603 ( .A1(n10796), .A2(n10226), .ZN(n9974) );
  OR2_X1 U12604 ( .A1(n9957), .A2(n9973), .ZN(n10794) );
  INV_X1 U12605 ( .A(n10794), .ZN(n10225) );
  AOI21_X1 U12606 ( .B1(n10797), .B2(n9974), .A(n10225), .ZN(n11060) );
  NAND2_X1 U12607 ( .A1(n15518), .A2(n11060), .ZN(n9998) );
  NAND2_X1 U12608 ( .A1(n9975), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9976) );
  NAND2_X1 U12609 ( .A1(n6809), .A2(n9977), .ZN(n12619) );
  AND2_X1 U12610 ( .A1(n11065), .A2(n15314), .ZN(n9996) );
  NAND3_X1 U12611 ( .A1(n10224), .A2(n12619), .A3(n15742), .ZN(n9978) );
  NAND2_X1 U12612 ( .A1(n9980), .A2(n8093), .ZN(n10010) );
  NAND2_X1 U12613 ( .A1(n9982), .A2(n9981), .ZN(n10004) );
  NAND4_X1 U12614 ( .A1(n9983), .A2(n10005), .A3(n10004), .A4(n14910), .ZN(
        n10009) );
  NAND2_X1 U12615 ( .A1(n9998), .A2(n11063), .ZN(n10001) );
  AND2_X1 U12616 ( .A1(n10001), .A2(n10224), .ZN(n15632) );
  INV_X1 U12617 ( .A(n9984), .ZN(n10197) );
  INV_X1 U12618 ( .A(n10197), .ZN(n13187) );
  OR2_X1 U12619 ( .A1(n12619), .A2(n13187), .ZN(n14922) );
  NAND2_X1 U12620 ( .A1(n14936), .A2(n15637), .ZN(n9995) );
  INV_X1 U12621 ( .A(n9985), .ZN(n13038) );
  NAND2_X1 U12622 ( .A1(n13038), .A2(n9986), .ZN(n9993) );
  INV_X1 U12623 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n10410) );
  NAND2_X1 U12624 ( .A1(n9987), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9989) );
  NAND2_X1 U12625 ( .A1(n12583), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9988) );
  OAI211_X1 U12626 ( .C1(n9990), .C2(n10410), .A(n9989), .B(n9988), .ZN(n9991)
         );
  INV_X1 U12627 ( .A(n9991), .ZN(n9992) );
  NAND2_X1 U12628 ( .A1(n9993), .A2(n9992), .ZN(n14934) );
  NAND2_X1 U12629 ( .A1(n14934), .A2(n15636), .ZN(n9994) );
  AND2_X1 U12630 ( .A1(n9995), .A2(n9994), .ZN(n15398) );
  OR2_X1 U12631 ( .A1(n12619), .A2(n9996), .ZN(n10738) );
  INV_X1 U12632 ( .A(n10187), .ZN(n9997) );
  NAND3_X1 U12633 ( .A1(n10738), .A2(n9997), .A3(n9477), .ZN(n9999) );
  INV_X1 U12634 ( .A(n9999), .ZN(n10000) );
  NAND2_X1 U12635 ( .A1(n10001), .A2(n10000), .ZN(n10002) );
  AOI22_X1 U12636 ( .A1(n15132), .A2(n14926), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10003) );
  OAI21_X1 U12637 ( .B1(n15398), .B2(n14928), .A(n10003), .ZN(n10007) );
  NOR3_X1 U12638 ( .A1(n10005), .A2(n15634), .A3(n10004), .ZN(n10006) );
  AOI211_X1 U12639 ( .C1(n14930), .C2(n15135), .A(n10007), .B(n10006), .ZN(
        n10008) );
  NAND3_X1 U12640 ( .A1(n10010), .A2(n10009), .A3(n10008), .ZN(P1_U3220) );
  AOI21_X1 U12641 ( .B1(n10011), .B2(n12983), .A(n14534), .ZN(n10013) );
  AOI22_X1 U12642 ( .A1(n14217), .A2(n14193), .B1(n14192), .B2(n14219), .ZN(
        n13176) );
  INV_X1 U12643 ( .A(n10015), .ZN(n10016) );
  NAND2_X1 U12644 ( .A1(n13180), .A2(n10017), .ZN(n10018) );
  NAND2_X1 U12645 ( .A1(n10022), .A2(n8102), .ZN(P2_U3527) );
  NAND2_X1 U12646 ( .A1(n10024), .A2(n8101), .ZN(P2_U3495) );
  AOI211_X1 U12647 ( .C1(n13557), .C2(n10026), .A(n15911), .B(n10025), .ZN(
        n10027) );
  INV_X1 U12648 ( .A(n10027), .ZN(n10031) );
  OAI22_X1 U12649 ( .A1(n13267), .A2(n15916), .B1(n15914), .B2(n10028), .ZN(
        n10029) );
  INV_X1 U12650 ( .A(n10029), .ZN(n10030) );
  INV_X1 U12651 ( .A(n10032), .ZN(n10037) );
  OAI22_X1 U12652 ( .A1(n15948), .A2(n11596), .B1(n13735), .B2(n11128), .ZN(
        n10033) );
  NAND2_X1 U12653 ( .A1(n10033), .A2(n13529), .ZN(n10034) );
  NAND2_X1 U12654 ( .A1(n10034), .A2(n13514), .ZN(n10035) );
  NAND2_X1 U12655 ( .A1(n14024), .A2(n10035), .ZN(n10036) );
  OAI21_X1 U12656 ( .B1(n14024), .B2(n10037), .A(n10036), .ZN(n10038) );
  MUX2_X1 U12657 ( .A(P3_REG1_REG_28__SCAN_IN), .B(n13188), .S(n15976), .Z(
        n10040) );
  INV_X1 U12658 ( .A(n10040), .ZN(n10044) );
  INV_X1 U12659 ( .A(n13269), .ZN(n13075) );
  OAI22_X1 U12660 ( .A1(n13192), .A2(n13945), .B1(n13075), .B2(n13940), .ZN(
        n10042) );
  INV_X1 U12661 ( .A(n10042), .ZN(n10043) );
  AND3_X1 U12662 ( .A1(n11768), .A2(P2_STATE_REG_SCAN_IN), .A3(n10045), .ZN(
        n10046) );
  NOR2_X4 U12663 ( .A1(n9477), .A2(n10047), .ZN(P1_U4016) );
  INV_X1 U12664 ( .A(n11260), .ZN(n10048) );
  INV_X1 U12665 ( .A(n13614), .ZN(n10618) );
  INV_X1 U12666 ( .A(n10115), .ZN(n10509) );
  NAND2_X1 U12667 ( .A1(n8151), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10050) );
  OAI21_X1 U12668 ( .B1(n11295), .B2(n10049), .A(n10050), .ZN(n11281) );
  OR2_X1 U12669 ( .A1(n11281), .A2(n11280), .ZN(n11283) );
  NAND2_X1 U12670 ( .A1(n11283), .A2(n10050), .ZN(n11377) );
  XNOR2_X1 U12671 ( .A(n11391), .B(n10092), .ZN(n11378) );
  NAND2_X1 U12672 ( .A1(n11391), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10051) );
  NAND2_X1 U12673 ( .A1(n10052), .A2(n10523), .ZN(n11684) );
  NAND2_X1 U12674 ( .A1(n11697), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n10053) );
  XNOR2_X1 U12675 ( .A(n10484), .B(P3_REG2_REG_6__SCAN_IN), .ZN(n11611) );
  INV_X1 U12676 ( .A(n10056), .ZN(n10173) );
  XNOR2_X1 U12677 ( .A(n10115), .B(n11763), .ZN(n10174) );
  AND2_X1 U12678 ( .A1(n10057), .A2(n7632), .ZN(n10058) );
  XNOR2_X1 U12679 ( .A(n10505), .B(P3_REG2_REG_10__SCAN_IN), .ZN(n10147) );
  XNOR2_X1 U12680 ( .A(n13614), .B(n12105), .ZN(n13607) );
  AOI21_X1 U12681 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n10618), .A(n13610), 
        .ZN(n10060) );
  NOR2_X1 U12682 ( .A1(n10060), .A2(n7091), .ZN(n10062) );
  OR2_X1 U12683 ( .A1(n10782), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n10061) );
  NAND2_X1 U12684 ( .A1(n10782), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n13647) );
  AND2_X1 U12685 ( .A1(n10061), .A2(n13647), .ZN(n10130) );
  OR3_X1 U12686 ( .A1(n10062), .A2(n13625), .A3(n10130), .ZN(n10067) );
  OR2_X1 U12687 ( .A1(n11259), .A2(P3_U3151), .ZN(n13569) );
  NAND2_X1 U12688 ( .A1(n11271), .A2(n13569), .ZN(n10140) );
  NAND2_X1 U12689 ( .A1(n13519), .A2(n11259), .ZN(n10064) );
  NAND2_X1 U12690 ( .A1(n10064), .A2(n10063), .ZN(n10139) );
  INV_X1 U12691 ( .A(n10139), .ZN(n10065) );
  NAND2_X1 U12692 ( .A1(n10140), .A2(n10065), .ZN(n10138) );
  AOI21_X1 U12693 ( .B1(n13642), .B2(n10067), .A(n13757), .ZN(n10145) );
  INV_X1 U12694 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10277) );
  XNOR2_X1 U12695 ( .A(n11391), .B(n10277), .ZN(n11375) );
  AND2_X1 U12696 ( .A1(n11217), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10068) );
  NAND2_X1 U12697 ( .A1(n8151), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10069) );
  OAI21_X1 U12698 ( .B1(n11295), .B2(n10068), .A(n10069), .ZN(n11288) );
  INV_X1 U12699 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15961) );
  NAND2_X1 U12700 ( .A1(n11391), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10070) );
  INV_X1 U12701 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15963) );
  INV_X1 U12702 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15965) );
  XNOR2_X1 U12703 ( .A(n11697), .B(n15965), .ZN(n11678) );
  NAND2_X1 U12704 ( .A1(n10071), .A2(n11678), .ZN(n11682) );
  NAND2_X1 U12705 ( .A1(n11697), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n10072) );
  INV_X1 U12706 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15967) );
  INV_X1 U12707 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15969) );
  XNOR2_X1 U12708 ( .A(n10484), .B(n15969), .ZN(n11614) );
  NAND2_X1 U12709 ( .A1(n10073), .A2(n11614), .ZN(n11618) );
  NAND2_X1 U12710 ( .A1(n10484), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n10074) );
  XNOR2_X1 U12711 ( .A(n10115), .B(P3_REG1_REG_8__SCAN_IN), .ZN(n10166) );
  INV_X1 U12712 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15974) );
  OR2_X1 U12713 ( .A1(n10115), .A2(n15974), .ZN(n10076) );
  INV_X1 U12714 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n12154) );
  INV_X1 U12715 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n12116) );
  NAND2_X1 U12716 ( .A1(n10077), .A2(n11964), .ZN(n10079) );
  AND2_X1 U12717 ( .A1(n10078), .A2(n10079), .ZN(n11962) );
  NAND2_X1 U12718 ( .A1(n11961), .A2(n10079), .ZN(n13616) );
  INV_X1 U12719 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n10292) );
  OR2_X1 U12720 ( .A1(n13614), .A2(n10292), .ZN(n10081) );
  NAND2_X1 U12721 ( .A1(n13614), .A2(n10292), .ZN(n10080) );
  AND2_X1 U12722 ( .A1(n10081), .A2(n10080), .ZN(n13617) );
  NAND2_X1 U12723 ( .A1(n13616), .A2(n13617), .ZN(n13615) );
  OR2_X1 U12724 ( .A1(n10782), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n10084) );
  NAND2_X1 U12725 ( .A1(n10782), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n13655) );
  AND2_X1 U12726 ( .A1(n10084), .A2(n13655), .ZN(n10131) );
  NAND3_X1 U12727 ( .A1(n13637), .A2(n7624), .A3(n10085), .ZN(n10087) );
  INV_X1 U12728 ( .A(n10138), .ZN(n10086) );
  INV_X1 U12729 ( .A(n13754), .ZN(n11321) );
  AOI21_X1 U12730 ( .B1(n13656), .B2(n10087), .A(n11321), .ZN(n10144) );
  MUX2_X1 U12731 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n7288), .Z(n10127) );
  INV_X1 U12732 ( .A(n10127), .ZN(n10128) );
  INV_X1 U12733 ( .A(n11295), .ZN(n10088) );
  NAND2_X1 U12734 ( .A1(n10089), .A2(n10088), .ZN(n11381) );
  INV_X1 U12735 ( .A(n10089), .ZN(n10090) );
  NAND2_X1 U12736 ( .A1(n10090), .A2(n11295), .ZN(n10091) );
  NOR2_X1 U12737 ( .A1(n11216), .A2(n11217), .ZN(n11284) );
  NAND2_X1 U12738 ( .A1(n8087), .A2(n11284), .ZN(n11382) );
  MUX2_X1 U12739 ( .A(n10092), .B(n10277), .S(n13717), .Z(n10094) );
  NAND2_X1 U12740 ( .A1(n10094), .A2(n10093), .ZN(n10097) );
  INV_X1 U12741 ( .A(n10094), .ZN(n10095) );
  NAND2_X1 U12742 ( .A1(n10095), .A2(n11391), .ZN(n10096) );
  NAND2_X1 U12743 ( .A1(n10097), .A2(n10096), .ZN(n11380) );
  INV_X1 U12744 ( .A(n10097), .ZN(n13599) );
  MUX2_X1 U12745 ( .A(n11529), .B(n15963), .S(n13717), .Z(n10098) );
  INV_X1 U12746 ( .A(n10523), .ZN(n13593) );
  NAND2_X1 U12747 ( .A1(n10098), .A2(n13593), .ZN(n11691) );
  INV_X1 U12748 ( .A(n10098), .ZN(n10099) );
  NAND2_X1 U12749 ( .A1(n10099), .A2(n10523), .ZN(n10100) );
  MUX2_X1 U12750 ( .A(n11506), .B(n15965), .S(n13717), .Z(n10101) );
  NAND2_X1 U12751 ( .A1(n10101), .A2(n6902), .ZN(n11645) );
  INV_X1 U12752 ( .A(n10101), .ZN(n10102) );
  NAND2_X1 U12753 ( .A1(n10102), .A2(n11697), .ZN(n10103) );
  NAND2_X1 U12754 ( .A1(n11645), .A2(n10103), .ZN(n11690) );
  AOI21_X1 U12755 ( .B1(n13598), .B2(n11691), .A(n11690), .ZN(n11643) );
  MUX2_X1 U12756 ( .A(n11632), .B(n15967), .S(n7288), .Z(n10104) );
  NAND2_X1 U12757 ( .A1(n10104), .A2(n11650), .ZN(n11625) );
  INV_X1 U12758 ( .A(n10104), .ZN(n10105) );
  NAND2_X1 U12759 ( .A1(n10105), .A2(n10530), .ZN(n10106) );
  NAND2_X1 U12760 ( .A1(n11625), .A2(n10106), .ZN(n11644) );
  INV_X1 U12761 ( .A(n11644), .ZN(n10107) );
  MUX2_X1 U12762 ( .A(n11519), .B(n15969), .S(n7288), .Z(n10108) );
  INV_X1 U12763 ( .A(n10484), .ZN(n11630) );
  NAND2_X1 U12764 ( .A1(n10108), .A2(n11630), .ZN(n11135) );
  INV_X1 U12765 ( .A(n10108), .ZN(n10109) );
  NAND2_X1 U12766 ( .A1(n10109), .A2(n10484), .ZN(n10110) );
  NAND2_X1 U12767 ( .A1(n11135), .A2(n10110), .ZN(n11624) );
  INV_X1 U12768 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15971) );
  MUX2_X1 U12769 ( .A(n11887), .B(n15971), .S(n7288), .Z(n10111) );
  NAND2_X1 U12770 ( .A1(n10111), .A2(n7077), .ZN(n10163) );
  INV_X1 U12771 ( .A(n10111), .ZN(n10112) );
  NAND2_X1 U12772 ( .A1(n10112), .A2(n11145), .ZN(n10113) );
  NAND2_X1 U12773 ( .A1(n10163), .A2(n10113), .ZN(n11136) );
  INV_X1 U12774 ( .A(n11136), .ZN(n10114) );
  MUX2_X1 U12775 ( .A(n11763), .B(n15974), .S(n7288), .Z(n10116) );
  NAND2_X1 U12776 ( .A1(n10116), .A2(n10115), .ZN(n10117) );
  OAI21_X1 U12777 ( .B1(n10116), .B2(n10115), .A(n10117), .ZN(n10162) );
  INV_X1 U12778 ( .A(n10117), .ZN(n11311) );
  MUX2_X1 U12779 ( .A(n11928), .B(n12154), .S(n7288), .Z(n10118) );
  NAND2_X1 U12780 ( .A1(n10118), .A2(n7632), .ZN(n10154) );
  INV_X1 U12781 ( .A(n10118), .ZN(n10119) );
  NAND2_X1 U12782 ( .A1(n10119), .A2(n11317), .ZN(n10120) );
  AND2_X1 U12783 ( .A1(n10154), .A2(n10120), .ZN(n11310) );
  MUX2_X1 U12784 ( .A(n12110), .B(n12116), .S(n7288), .Z(n10122) );
  INV_X1 U12785 ( .A(n10505), .ZN(n10121) );
  NAND2_X1 U12786 ( .A1(n10122), .A2(n10121), .ZN(n10125) );
  INV_X1 U12787 ( .A(n10122), .ZN(n10123) );
  NAND2_X1 U12788 ( .A1(n10123), .A2(n10505), .ZN(n10124) );
  NAND2_X1 U12789 ( .A1(n10125), .A2(n10124), .ZN(n10153) );
  AOI21_X1 U12790 ( .B1(n11309), .B2(n10154), .A(n10153), .ZN(n10152) );
  INV_X1 U12791 ( .A(n10125), .ZN(n10126) );
  XNOR2_X1 U12792 ( .A(n10127), .B(n11964), .ZN(n11965) );
  MUX2_X1 U12793 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n7288), .Z(n10129) );
  XNOR2_X1 U12794 ( .A(n10129), .B(n13614), .ZN(n13619) );
  NAND2_X1 U12795 ( .A1(n10129), .A2(n10618), .ZN(n13630) );
  MUX2_X1 U12796 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n7288), .Z(n10132) );
  XOR2_X1 U12797 ( .A(n10744), .B(n10132), .Z(n13629) );
  MUX2_X1 U12798 ( .A(n10131), .B(n10130), .S(n13736), .Z(n10134) );
  INV_X1 U12799 ( .A(n10132), .ZN(n10133) );
  NAND2_X1 U12800 ( .A1(n10133), .A2(n7091), .ZN(n10135) );
  INV_X1 U12801 ( .A(n13649), .ZN(n10137) );
  AOI21_X1 U12802 ( .B1(n13633), .B2(n10135), .A(n10134), .ZN(n10136) );
  NOR3_X1 U12803 ( .A1(n10137), .A2(n10136), .A3(n13720), .ZN(n10143) );
  MUX2_X1 U12804 ( .A(n10138), .B(n13577), .S(n13566), .Z(n13746) );
  NAND2_X1 U12805 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n12330)
         );
  NAND2_X1 U12806 ( .A1(n15894), .A2(P3_ADDR_REG_14__SCAN_IN), .ZN(n10141) );
  OAI211_X1 U12807 ( .C1(n13746), .C2(n10782), .A(n12330), .B(n10141), .ZN(
        n10142) );
  OR4_X1 U12808 ( .A1(n10145), .A2(n10144), .A3(n10143), .A4(n10142), .ZN(
        P3_U3196) );
  NAND3_X1 U12809 ( .A1(n11307), .A2(n10147), .A3(n10146), .ZN(n10148) );
  AOI21_X1 U12810 ( .B1(n6756), .B2(n10148), .A(n13757), .ZN(n10161) );
  NAND3_X1 U12811 ( .A1(n11304), .A2(n6786), .A3(n10149), .ZN(n10150) );
  AOI21_X1 U12812 ( .B1(n10151), .B2(n10150), .A(n11321), .ZN(n10160) );
  INV_X1 U12813 ( .A(n10152), .ZN(n10156) );
  NAND3_X1 U12814 ( .A1(n11309), .A2(n10154), .A3(n10153), .ZN(n10155) );
  AOI21_X1 U12815 ( .B1(n10156), .B2(n10155), .A(n13720), .ZN(n10159) );
  NAND2_X1 U12816 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n12040)
         );
  NAND2_X1 U12817 ( .A1(n15894), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n10157) );
  OAI211_X1 U12818 ( .C1(n13746), .C2(n10505), .A(n12040), .B(n10157), .ZN(
        n10158) );
  OR4_X1 U12819 ( .A1(n10161), .A2(n10160), .A3(n10159), .A4(n10158), .ZN(
        P3_U3192) );
  INV_X1 U12820 ( .A(n11312), .ZN(n10165) );
  NAND3_X1 U12821 ( .A1(n11137), .A2(n10163), .A3(n10162), .ZN(n10164) );
  AOI21_X1 U12822 ( .B1(n10165), .B2(n10164), .A(n13720), .ZN(n10181) );
  INV_X1 U12823 ( .A(n10166), .ZN(n10168) );
  NAND3_X1 U12824 ( .A1(n11139), .A2(n10168), .A3(n10167), .ZN(n10169) );
  AOI21_X1 U12825 ( .B1(n10170), .B2(n10169), .A(n11321), .ZN(n10180) );
  INV_X1 U12826 ( .A(n10171), .ZN(n10176) );
  NAND3_X1 U12827 ( .A1(n10172), .A2(n10174), .A3(n10173), .ZN(n10175) );
  AOI21_X1 U12828 ( .B1(n10176), .B2(n10175), .A(n13757), .ZN(n10179) );
  NAND2_X1 U12829 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n12176) );
  NAND2_X1 U12830 ( .A1(n15894), .A2(P3_ADDR_REG_8__SCAN_IN), .ZN(n10177) );
  OAI211_X1 U12831 ( .C1(n13746), .C2(n10509), .A(n12176), .B(n10177), .ZN(
        n10178) );
  OR4_X1 U12832 ( .A1(n10181), .A2(n10180), .A3(n10179), .A4(n10178), .ZN(
        P3_U3190) );
  NAND2_X1 U12833 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10198) );
  OAI21_X1 U12834 ( .B1(n10184), .B2(n10183), .A(n10182), .ZN(n10739) );
  MUX2_X1 U12835 ( .A(n10198), .B(n10739), .S(n7374), .Z(n10186) );
  OAI21_X1 U12836 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n7374), .A(n10197), .ZN(
        n15647) );
  INV_X1 U12837 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n14964) );
  NAND2_X1 U12838 ( .A1(n15647), .A2(n14964), .ZN(n10185) );
  OAI211_X1 U12839 ( .C1(n10186), .C2(n13187), .A(P1_U4016), .B(n10185), .ZN(
        n15000) );
  INV_X1 U12840 ( .A(n15000), .ZN(n10206) );
  INV_X1 U12841 ( .A(n10224), .ZN(n11062) );
  NAND2_X1 U12842 ( .A1(n10187), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12656) );
  NAND2_X1 U12843 ( .A1(n11062), .A2(n12656), .ZN(n10190) );
  OR2_X1 U12844 ( .A1(n12619), .A2(n10187), .ZN(n10188) );
  AOI22_X1 U12845 ( .A1(n15651), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n10196) );
  MUX2_X1 U12846 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9487), .S(n10582), .Z(
        n10193) );
  INV_X1 U12847 ( .A(n10488), .ZN(n14967) );
  AOI21_X1 U12848 ( .B1(n14967), .B2(P1_REG1_REG_1__SCAN_IN), .A(n14962), .ZN(
        n10192) );
  NOR2_X1 U12849 ( .A1(n10192), .A2(n10193), .ZN(n14982) );
  NAND2_X1 U12850 ( .A1(n10190), .A2(n10189), .ZN(n15654) );
  INV_X1 U12851 ( .A(n7374), .ZN(n10191) );
  AOI211_X1 U12852 ( .C1(n10193), .C2(n10192), .A(n14982), .B(n15661), .ZN(
        n10194) );
  INV_X1 U12853 ( .A(n10194), .ZN(n10195) );
  NAND2_X1 U12854 ( .A1(n10196), .A2(n10195), .ZN(n10205) );
  INV_X1 U12855 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n11177) );
  MUX2_X1 U12856 ( .A(n11177), .B(P1_REG2_REG_2__SCAN_IN), .S(n10582), .Z(
        n10202) );
  MUX2_X1 U12857 ( .A(n9458), .B(P1_REG2_REG_1__SCAN_IN), .S(n10488), .Z(
        n14961) );
  INV_X1 U12858 ( .A(n10198), .ZN(n14960) );
  NAND2_X1 U12859 ( .A1(n14961), .A2(n14960), .ZN(n14959) );
  NAND2_X1 U12860 ( .A1(n14967), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10199) );
  NAND2_X1 U12861 ( .A1(n14959), .A2(n10199), .ZN(n10201) );
  OR2_X1 U12862 ( .A1(n13187), .A2(n7374), .ZN(n10200) );
  NAND2_X1 U12863 ( .A1(n10201), .A2(n10202), .ZN(n10585) );
  OAI211_X1 U12864 ( .C1(n10202), .C2(n10201), .A(n15665), .B(n10585), .ZN(
        n10203) );
  OAI21_X1 U12865 ( .B1(n15659), .B2(n10582), .A(n10203), .ZN(n10204) );
  OR3_X1 U12866 ( .A1(n10206), .A2(n10205), .A3(n10204), .ZN(P1_U3245) );
  MUX2_X1 U12867 ( .A(P1_RD_REG_SCAN_IN), .B(n10207), .S(P2_RD_REG_SCAN_IN), 
        .Z(n10208) );
  INV_X1 U12868 ( .A(P3_RD_REG_SCAN_IN), .ZN(n10409) );
  NAND2_X1 U12869 ( .A1(n10208), .A2(n10409), .ZN(U29) );
  INV_X1 U12870 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n10209) );
  AOI21_X1 U12871 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n10209), .A(n7235), .ZN(
        n10211) );
  INV_X1 U12872 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10210) );
  NOR2_X1 U12873 ( .A1(n10211), .A2(n10210), .ZN(n15983) );
  AOI21_X1 U12874 ( .B1(n10211), .B2(n10210), .A(n15983), .ZN(SUB_1596_U53) );
  INV_X2 U12875 ( .A(n13080), .ZN(n13196) );
  NAND2_X1 U12876 ( .A1(n9260), .A2(P2_U3088), .ZN(n12667) );
  INV_X1 U12877 ( .A(n10212), .ZN(n10215) );
  OAI222_X1 U12878 ( .A1(n13196), .A2(n10213), .B1(n12667), .B2(n10215), .C1(
        P2_U3088), .C2(n14277), .ZN(P2_U3324) );
  NOR2_X1 U12879 ( .A1(n10481), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15550) );
  NAND2_X2 U12880 ( .A1(n9260), .A2(P1_U3086), .ZN(n15546) );
  OAI222_X1 U12881 ( .A1(n14977), .A2(P1_U3086), .B1(n10985), .B2(n10215), 
        .C1(n10214), .C2(n15546), .ZN(P1_U3352) );
  INV_X1 U12882 ( .A(n10216), .ZN(n10218) );
  AOI22_X1 U12883 ( .A1(n10674), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n13080), .ZN(n10217) );
  OAI21_X1 U12884 ( .B1(n10218), .B2(n12667), .A(n10217), .ZN(P2_U3322) );
  INV_X1 U12885 ( .A(n10602), .ZN(n10579) );
  OAI222_X1 U12886 ( .A1(n15546), .A2(n7585), .B1(n10985), .B2(n10218), .C1(
        n10579), .C2(P1_U3086), .ZN(P1_U3350) );
  INV_X1 U12887 ( .A(n10219), .ZN(n10497) );
  INV_X1 U12888 ( .A(n10588), .ZN(n14988) );
  OAI222_X1 U12889 ( .A1(n15546), .A2(n7358), .B1(n10985), .B2(n10497), .C1(
        n14988), .C2(P1_U3086), .ZN(P1_U3351) );
  INV_X1 U12890 ( .A(n10220), .ZN(n10492) );
  INV_X1 U12891 ( .A(n15007), .ZN(n10221) );
  OAI222_X1 U12892 ( .A1(n15546), .A2(n7345), .B1(n10985), .B2(n10492), .C1(
        n10221), .C2(P1_U3086), .ZN(P1_U3349) );
  INV_X1 U12893 ( .A(n10222), .ZN(n10485) );
  INV_X1 U12894 ( .A(n15546), .ZN(n10679) );
  AOI22_X1 U12895 ( .A1(n10768), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n10679), .ZN(n10223) );
  OAI21_X1 U12896 ( .B1(n10485), .B2(n10985), .A(n10223), .ZN(P1_U3348) );
  AOI22_X1 U12897 ( .A1(n15729), .A2(n10226), .B1(n10225), .B2(n10228), .ZN(
        P1_U3446) );
  INV_X1 U12898 ( .A(n10227), .ZN(n10229) );
  AOI22_X1 U12899 ( .A1(n15729), .A2(n10230), .B1(n10229), .B2(n10228), .ZN(
        P1_U3445) );
  INV_X1 U12900 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n15800) );
  NAND4_X1 U12901 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P2_DATAO_REG_5__SCAN_IN), 
        .A3(P3_DATAO_REG_15__SCAN_IN), .A4(n15800), .ZN(n10271) );
  NAND4_X1 U12902 ( .A1(P3_REG2_REG_5__SCAN_IN), .A2(P1_REG3_REG_13__SCAN_IN), 
        .A3(n14915), .A4(n10387), .ZN(n10270) );
  NOR4_X1 U12903 ( .A1(P3_REG3_REG_21__SCAN_IN), .A2(P3_REG2_REG_1__SCAN_IN), 
        .A3(P1_IR_REG_4__SCAN_IN), .A4(P2_ADDR_REG_10__SCAN_IN), .ZN(n10237)
         );
  NOR4_X1 U12904 ( .A1(SI_11_), .A2(P1_REG3_REG_19__SCAN_IN), .A3(
        P1_REG1_REG_5__SCAN_IN), .A4(P1_REG3_REG_1__SCAN_IN), .ZN(n10236) );
  NAND4_X1 U12905 ( .A1(P2_REG0_REG_2__SCAN_IN), .A2(P2_REG0_REG_29__SCAN_IN), 
        .A3(P3_RD_REG_SCAN_IN), .A4(n10410), .ZN(n10234) );
  NAND4_X1 U12906 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P2_REG1_REG_3__SCAN_IN), 
        .A3(n10403), .A4(n11887), .ZN(n10232) );
  NAND4_X1 U12907 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P2_REG0_REG_24__SCAN_IN), 
        .A3(n13983), .A4(n8243), .ZN(n10231) );
  OR4_X1 U12908 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(n10232), .A3(n10231), .A4(
        P2_REG1_REG_1__SCAN_IN), .ZN(n10233) );
  NOR4_X1 U12909 ( .A1(n10234), .A2(n12154), .A3(n10233), .A4(
        P1_DATAO_REG_21__SCAN_IN), .ZN(n10235) );
  NAND3_X1 U12910 ( .A1(n10237), .A2(n10236), .A3(n10235), .ZN(n10269) );
  AND4_X1 U12911 ( .A1(SI_31_), .A2(P1_REG1_REG_15__SCAN_IN), .A3(
        P2_REG1_REG_16__SCAN_IN), .A4(n8218), .ZN(n10244) );
  INV_X1 U12912 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n15854) );
  AND4_X1 U12913 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_5__SCAN_IN), .A3(
        P3_REG0_REG_24__SCAN_IN), .A4(n15854), .ZN(n10243) );
  INV_X1 U12914 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10238) );
  INV_X1 U12915 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n11731) );
  NAND4_X1 U12916 ( .A1(n10238), .A2(n11731), .A3(P3_REG0_REG_19__SCAN_IN), 
        .A4(P2_REG2_REG_26__SCAN_IN), .ZN(n10241) );
  NAND3_X1 U12917 ( .A1(n7358), .A2(n10239), .A3(P2_ADDR_REG_15__SCAN_IN), 
        .ZN(n10240) );
  NOR2_X1 U12918 ( .A1(n10241), .A2(n10240), .ZN(n10242) );
  INV_X1 U12919 ( .A(P3_DATAO_REG_1__SCAN_IN), .ZN(n10855) );
  AND4_X1 U12920 ( .A1(n10244), .A2(n10243), .A3(n10242), .A4(n10855), .ZN(
        n10267) );
  INV_X1 U12921 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n11023) );
  NAND4_X1 U12922 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        n10245), .A4(n11023), .ZN(n10249) );
  NAND4_X1 U12923 ( .A1(P3_REG1_REG_20__SCAN_IN), .A2(P2_DATAO_REG_8__SCAN_IN), 
        .A3(P2_D_REG_7__SCAN_IN), .A4(n10292), .ZN(n10248) );
  NAND4_X1 U12924 ( .A1(SI_0_), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_REG0_REG_9__SCAN_IN), .A4(P2_REG1_REG_14__SCAN_IN), .ZN(n10247) );
  NAND4_X1 U12925 ( .A1(n10491), .A2(P2_REG1_REG_15__SCAN_IN), .A3(
        P2_REG0_REG_12__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n10246) );
  NOR4_X1 U12926 ( .A1(n10249), .A2(n10248), .A3(n10247), .A4(n10246), .ZN(
        n10266) );
  AND4_X1 U12927 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P2_DATAO_REG_30__SCAN_IN), 
        .A3(P1_REG1_REG_24__SCAN_IN), .A4(P1_REG0_REG_3__SCAN_IN), .ZN(n10251)
         );
  AND4_X1 U12928 ( .A1(n10365), .A2(n11460), .A3(n15648), .A4(n10251), .ZN(
        n10254) );
  AND4_X1 U12929 ( .A1(P1_REG0_REG_2__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), 
        .A3(P2_D_REG_6__SCAN_IN), .A4(P3_DATAO_REG_21__SCAN_IN), .ZN(n10253)
         );
  AND4_X1 U12930 ( .A1(n10355), .A2(n10353), .A3(P1_ADDR_REG_16__SCAN_IN), 
        .A4(P3_D_REG_25__SCAN_IN), .ZN(n10252) );
  INV_X1 U12931 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10819) );
  AND4_X1 U12932 ( .A1(n10254), .A2(n10253), .A3(n10252), .A4(n10819), .ZN(
        n10265) );
  NAND4_X1 U12933 ( .A1(P3_REG2_REG_27__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .A3(n9590), .A4(n11935), .ZN(n10263) );
  INV_X1 U12934 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n10257) );
  INV_X1 U12935 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10255) );
  NAND4_X1 U12936 ( .A1(n10257), .A2(n10256), .A3(n10255), .A4(
        P2_REG2_REG_27__SCAN_IN), .ZN(n10262) );
  NAND4_X1 U12937 ( .A1(n11772), .A2(n10781), .A3(n10258), .A4(
        P1_DATAO_REG_1__SCAN_IN), .ZN(n10261) );
  NAND4_X1 U12938 ( .A1(n10259), .A2(n8829), .A3(n14518), .A4(
        P2_D_REG_29__SCAN_IN), .ZN(n10260) );
  NOR4_X1 U12939 ( .A1(n10263), .A2(n10262), .A3(n10261), .A4(n10260), .ZN(
        n10264) );
  NAND4_X1 U12940 ( .A1(n10267), .A2(n10266), .A3(n10265), .A4(n10264), .ZN(
        n10268) );
  NOR4_X1 U12941 ( .A1(n10271), .A2(n10270), .A3(n10269), .A4(n10268), .ZN(
        n10286) );
  OR4_X1 U12942 ( .A1(P1_REG0_REG_11__SCAN_IN), .A2(P1_REG1_REG_2__SCAN_IN), 
        .A3(P3_DATAO_REG_20__SCAN_IN), .A4(n11177), .ZN(n10284) );
  NOR4_X1 U12943 ( .A1(n12286), .A2(n10458), .A3(n10272), .A4(
        P2_REG3_REG_14__SCAN_IN), .ZN(n10282) );
  NOR4_X1 U12944 ( .A1(P3_REG0_REG_2__SCAN_IN), .A2(n10757), .A3(n10890), .A4(
        n10460), .ZN(n10276) );
  INV_X1 U12945 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n13900) );
  NOR4_X1 U12946 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n11519), .A3(n13900), .A4(
        n15092), .ZN(n10275) );
  AND4_X1 U12947 ( .A1(n10273), .A2(P2_ADDR_REG_6__SCAN_IN), .A3(n12407), .A4(
        n10950), .ZN(n10274) );
  NAND4_X1 U12948 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(n10276), .A3(n10275), .A4(
        n10274), .ZN(n10278) );
  NOR4_X1 U12949 ( .A1(n10278), .A2(n10277), .A3(P3_REG2_REG_23__SCAN_IN), 
        .A4(P3_REG2_REG_18__SCAN_IN), .ZN(n10281) );
  NOR4_X1 U12950 ( .A1(n10279), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_REG1_REG_31__SCAN_IN), .A4(P1_REG3_REG_14__SCAN_IN), .ZN(n10280) );
  NAND3_X1 U12951 ( .A1(n10282), .A2(n10281), .A3(n10280), .ZN(n10283) );
  INV_X1 U12952 ( .A(P3_DATAO_REG_22__SCAN_IN), .ZN(n11083) );
  INV_X1 U12953 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10818) );
  NOR4_X1 U12954 ( .A1(n10284), .A2(n10283), .A3(n11083), .A4(n10818), .ZN(
        n10285) );
  AOI21_X1 U12955 ( .B1(n10286), .B2(n10285), .A(n10437), .ZN(n10477) );
  INV_X1 U12956 ( .A(keyinput73), .ZN(n10476) );
  INV_X1 U12957 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15724) );
  AOI22_X1 U12958 ( .A1(n15724), .A2(keyinput111), .B1(keyinput71), .B2(n11023), .ZN(n10287) );
  OAI221_X1 U12959 ( .B1(n15724), .B2(keyinput111), .C1(n11023), .C2(
        keyinput71), .A(n10287), .ZN(n10298) );
  INV_X1 U12960 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n15855) );
  AOI22_X1 U12961 ( .A1(n10289), .A2(keyinput48), .B1(keyinput74), .B2(n15855), 
        .ZN(n10288) );
  OAI221_X1 U12962 ( .B1(n10289), .B2(keyinput48), .C1(n15855), .C2(keyinput74), .A(n10288), .ZN(n10297) );
  AOI22_X1 U12963 ( .A1(n10292), .A2(keyinput20), .B1(n10291), .B2(keyinput29), 
        .ZN(n10290) );
  OAI221_X1 U12964 ( .B1(n10292), .B2(keyinput20), .C1(n10291), .C2(keyinput29), .A(n10290), .ZN(n10296) );
  XNOR2_X1 U12965 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput104), .ZN(n10294)
         );
  XNOR2_X1 U12966 ( .A(P3_REG3_REG_17__SCAN_IN), .B(keyinput2), .ZN(n10293) );
  NAND2_X1 U12967 ( .A1(n10294), .A2(n10293), .ZN(n10295) );
  NOR4_X1 U12968 ( .A1(n10298), .A2(n10297), .A3(n10296), .A4(n10295), .ZN(
        n10333) );
  INV_X1 U12969 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n15726) );
  AOI22_X1 U12970 ( .A1(n15726), .A2(keyinput66), .B1(keyinput6), .B2(n10300), 
        .ZN(n10299) );
  OAI221_X1 U12971 ( .B1(n15726), .B2(keyinput66), .C1(n10300), .C2(keyinput6), 
        .A(n10299), .ZN(n10308) );
  INV_X1 U12972 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n14632) );
  AOI22_X1 U12973 ( .A1(n8218), .A2(keyinput119), .B1(keyinput105), .B2(n14632), .ZN(n10301) );
  OAI221_X1 U12974 ( .B1(n8218), .B2(keyinput119), .C1(n14632), .C2(
        keyinput105), .A(n10301), .ZN(n10307) );
  INV_X1 U12975 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n15725) );
  AOI22_X1 U12976 ( .A1(n15725), .A2(keyinput31), .B1(keyinput45), .B2(n14639), 
        .ZN(n10302) );
  OAI221_X1 U12977 ( .B1(n15725), .B2(keyinput31), .C1(n14639), .C2(keyinput45), .A(n10302), .ZN(n10306) );
  XNOR2_X1 U12978 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput12), .ZN(n10304)
         );
  XNOR2_X1 U12979 ( .A(P2_REG0_REG_12__SCAN_IN), .B(keyinput106), .ZN(n10303)
         );
  NAND2_X1 U12980 ( .A1(n10304), .A2(n10303), .ZN(n10305) );
  NOR4_X1 U12981 ( .A1(n10308), .A2(n10307), .A3(n10306), .A4(n10305), .ZN(
        n10332) );
  INV_X1 U12982 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15586) );
  AOI22_X1 U12983 ( .A1(n15586), .A2(keyinput43), .B1(keyinput79), .B2(n10855), 
        .ZN(n10309) );
  OAI221_X1 U12984 ( .B1(n15586), .B2(keyinput43), .C1(n10855), .C2(keyinput79), .A(n10309), .ZN(n10319) );
  INV_X1 U12985 ( .A(SI_31_), .ZN(n10312) );
  INV_X1 U12986 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10311) );
  AOI22_X1 U12987 ( .A1(n10312), .A2(keyinput5), .B1(keyinput95), .B2(n10311), 
        .ZN(n10310) );
  OAI221_X1 U12988 ( .B1(n10312), .B2(keyinput5), .C1(n10311), .C2(keyinput95), 
        .A(n10310), .ZN(n10318) );
  XNOR2_X1 U12989 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput124), .ZN(n10316) );
  XNOR2_X1 U12990 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(keyinput25), .ZN(n10315)
         );
  XNOR2_X1 U12991 ( .A(P3_REG0_REG_24__SCAN_IN), .B(keyinput120), .ZN(n10314)
         );
  XNOR2_X1 U12992 ( .A(P3_IR_REG_5__SCAN_IN), .B(keyinput34), .ZN(n10313) );
  NAND4_X1 U12993 ( .A1(n10316), .A2(n10315), .A3(n10314), .A4(n10313), .ZN(
        n10317) );
  NOR3_X1 U12994 ( .A1(n10319), .A2(n10318), .A3(n10317), .ZN(n10331) );
  INV_X1 U12995 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n10321) );
  AOI22_X1 U12996 ( .A1(n10321), .A2(keyinput16), .B1(keyinput77), .B2(n15854), 
        .ZN(n10320) );
  OAI221_X1 U12997 ( .B1(n10321), .B2(keyinput16), .C1(n15854), .C2(keyinput77), .A(n10320), .ZN(n10329) );
  AOI22_X1 U12998 ( .A1(n14007), .A2(keyinput122), .B1(keyinput10), .B2(n9221), 
        .ZN(n10322) );
  OAI221_X1 U12999 ( .B1(n14007), .B2(keyinput122), .C1(n9221), .C2(keyinput10), .A(n10322), .ZN(n10328) );
  XOR2_X1 U13000 ( .A(n14310), .B(keyinput26), .Z(n10326) );
  XNOR2_X1 U13001 ( .A(P1_ADDR_REG_14__SCAN_IN), .B(keyinput64), .ZN(n10325)
         );
  XNOR2_X1 U13002 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(keyinput93), .ZN(n10324)
         );
  XNOR2_X1 U13003 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput91), .ZN(n10323) );
  NAND4_X1 U13004 ( .A1(n10326), .A2(n10325), .A3(n10324), .A4(n10323), .ZN(
        n10327) );
  NOR3_X1 U13005 ( .A1(n10329), .A2(n10328), .A3(n10327), .ZN(n10330) );
  NAND4_X1 U13006 ( .A1(n10333), .A2(n10332), .A3(n10331), .A4(n10330), .ZN(
        n10474) );
  INV_X1 U13007 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n15853) );
  AOI22_X1 U13008 ( .A1(n11772), .A2(keyinput50), .B1(keyinput101), .B2(n15853), .ZN(n10334) );
  OAI221_X1 U13009 ( .B1(n11772), .B2(keyinput50), .C1(n15853), .C2(
        keyinput101), .A(n10334), .ZN(n10342) );
  XNOR2_X1 U13010 ( .A(keyinput61), .B(n14518), .ZN(n10341) );
  XNOR2_X1 U13011 ( .A(keyinput18), .B(n8829), .ZN(n10340) );
  XNOR2_X1 U13012 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput58), .ZN(n10338)
         );
  XNOR2_X1 U13013 ( .A(P2_IR_REG_15__SCAN_IN), .B(keyinput60), .ZN(n10337) );
  XNOR2_X1 U13014 ( .A(P1_REG3_REG_5__SCAN_IN), .B(keyinput67), .ZN(n10336) );
  XNOR2_X1 U13015 ( .A(P1_REG0_REG_18__SCAN_IN), .B(keyinput94), .ZN(n10335)
         );
  NAND4_X1 U13016 ( .A1(n10338), .A2(n10337), .A3(n10336), .A4(n10335), .ZN(
        n10339) );
  NOR4_X1 U13017 ( .A1(n10342), .A2(n10341), .A3(n10340), .A4(n10339), .ZN(
        n10376) );
  AOI22_X1 U13018 ( .A1(n9590), .A2(keyinput108), .B1(keyinput28), .B2(n9508), 
        .ZN(n10343) );
  OAI221_X1 U13019 ( .B1(n9590), .B2(keyinput108), .C1(n9508), .C2(keyinput28), 
        .A(n10343), .ZN(n10351) );
  INV_X1 U13020 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n12269) );
  AOI22_X1 U13021 ( .A1(n12269), .A2(keyinput24), .B1(n10950), .B2(keyinput21), 
        .ZN(n10344) );
  OAI221_X1 U13022 ( .B1(n12269), .B2(keyinput24), .C1(n10950), .C2(keyinput21), .A(n10344), .ZN(n10350) );
  AOI22_X1 U13023 ( .A1(n8541), .A2(keyinput11), .B1(keyinput125), .B2(n11935), 
        .ZN(n10345) );
  OAI221_X1 U13024 ( .B1(n8541), .B2(keyinput11), .C1(n11935), .C2(keyinput125), .A(n10345), .ZN(n10349) );
  XNOR2_X1 U13025 ( .A(P1_REG3_REG_16__SCAN_IN), .B(keyinput88), .ZN(n10347)
         );
  XNOR2_X1 U13026 ( .A(SI_14_), .B(keyinput81), .ZN(n10346) );
  NAND2_X1 U13027 ( .A1(n10347), .A2(n10346), .ZN(n10348) );
  NOR4_X1 U13028 ( .A1(n10351), .A2(n10350), .A3(n10349), .A4(n10348), .ZN(
        n10375) );
  INV_X1 U13029 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n15856) );
  AOI22_X1 U13030 ( .A1(n10353), .A2(keyinput65), .B1(keyinput96), .B2(n15856), 
        .ZN(n10352) );
  OAI221_X1 U13031 ( .B1(n10353), .B2(keyinput65), .C1(n15856), .C2(keyinput96), .A(n10352), .ZN(n10362) );
  INV_X1 U13032 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n13199) );
  AOI22_X1 U13033 ( .A1(n13199), .A2(keyinput63), .B1(keyinput59), .B2(n10355), 
        .ZN(n10354) );
  OAI221_X1 U13034 ( .B1(n13199), .B2(keyinput63), .C1(n10355), .C2(keyinput59), .A(n10354), .ZN(n10361) );
  INV_X1 U13035 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10820) );
  XOR2_X1 U13036 ( .A(n10820), .B(keyinput98), .Z(n10359) );
  XNOR2_X1 U13037 ( .A(P1_REG1_REG_24__SCAN_IN), .B(keyinput107), .ZN(n10358)
         );
  XNOR2_X1 U13038 ( .A(P3_IR_REG_17__SCAN_IN), .B(keyinput42), .ZN(n10357) );
  XNOR2_X1 U13039 ( .A(P1_REG1_REG_0__SCAN_IN), .B(keyinput55), .ZN(n10356) );
  NAND4_X1 U13040 ( .A1(n10359), .A2(n10358), .A3(n10357), .A4(n10356), .ZN(
        n10360) );
  NOR3_X1 U13041 ( .A1(n10362), .A2(n10361), .A3(n10360), .ZN(n10374) );
  INV_X1 U13042 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n15598) );
  AOI22_X1 U13043 ( .A1(n9489), .A2(keyinput100), .B1(keyinput49), .B2(n15598), 
        .ZN(n10363) );
  OAI221_X1 U13044 ( .B1(n9489), .B2(keyinput100), .C1(n15598), .C2(keyinput49), .A(n10363), .ZN(n10369) );
  AOI22_X1 U13045 ( .A1(n11460), .A2(keyinput78), .B1(keyinput114), .B2(n12407), .ZN(n10364) );
  OAI221_X1 U13046 ( .B1(n11460), .B2(keyinput78), .C1(n12407), .C2(
        keyinput114), .A(n10364), .ZN(n10368) );
  XOR2_X1 U13047 ( .A(P2_IR_REG_9__SCAN_IN), .B(keyinput8), .Z(n10367) );
  XNOR2_X1 U13048 ( .A(n10365), .B(keyinput83), .ZN(n10366) );
  OR4_X1 U13049 ( .A1(n10369), .A2(n10368), .A3(n10367), .A4(n10366), .ZN(
        n10372) );
  INV_X1 U13050 ( .A(P3_DATAO_REG_21__SCAN_IN), .ZN(n10987) );
  XNOR2_X1 U13051 ( .A(n10987), .B(keyinput23), .ZN(n10371) );
  XNOR2_X1 U13052 ( .A(n10819), .B(keyinput118), .ZN(n10370) );
  NOR3_X1 U13053 ( .A1(n10372), .A2(n10371), .A3(n10370), .ZN(n10373) );
  NAND4_X1 U13054 ( .A1(n10376), .A2(n10375), .A3(n10374), .A4(n10373), .ZN(
        n10473) );
  AOI22_X1 U13055 ( .A1(n12154), .A2(keyinput82), .B1(keyinput0), .B2(n8888), 
        .ZN(n10377) );
  OAI221_X1 U13056 ( .B1(n12154), .B2(keyinput82), .C1(n8888), .C2(keyinput0), 
        .A(n10377), .ZN(n10385) );
  AOI22_X1 U13057 ( .A1(n15800), .A2(keyinput14), .B1(n11111), .B2(keyinput99), 
        .ZN(n10378) );
  OAI221_X1 U13058 ( .B1(n15800), .B2(keyinput14), .C1(n11111), .C2(keyinput99), .A(n10378), .ZN(n10384) );
  XNOR2_X1 U13059 ( .A(P1_REG3_REG_13__SCAN_IN), .B(keyinput80), .ZN(n10381)
         );
  XNOR2_X1 U13060 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput33), .ZN(n10380)
         );
  XNOR2_X1 U13061 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput4), .ZN(n10379) );
  NAND3_X1 U13062 ( .A1(n10381), .A2(n10380), .A3(n10379), .ZN(n10383) );
  INV_X1 U13063 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n10853) );
  XNOR2_X1 U13064 ( .A(n10853), .B(keyinput90), .ZN(n10382) );
  NOR4_X1 U13065 ( .A1(n10385), .A2(n10384), .A3(n10383), .A4(n10382), .ZN(
        n10423) );
  AOI22_X1 U13066 ( .A1(n10387), .A2(keyinput56), .B1(n11632), .B2(keyinput113), .ZN(n10386) );
  OAI221_X1 U13067 ( .B1(n10387), .B2(keyinput56), .C1(n11632), .C2(
        keyinput113), .A(n10386), .ZN(n10395) );
  AOI22_X1 U13068 ( .A1(n11068), .A2(keyinput68), .B1(n11280), .B2(keyinput102), .ZN(n10388) );
  OAI221_X1 U13069 ( .B1(n11068), .B2(keyinput68), .C1(n11280), .C2(
        keyinput102), .A(n10388), .ZN(n10394) );
  INV_X1 U13070 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n15839) );
  AOI22_X1 U13071 ( .A1(n15839), .A2(keyinput103), .B1(n14915), .B2(keyinput47), .ZN(n10389) );
  OAI221_X1 U13072 ( .B1(n15839), .B2(keyinput103), .C1(n14915), .C2(
        keyinput47), .A(n10389), .ZN(n10393) );
  XNOR2_X1 U13073 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput32), .ZN(n10391) );
  XNOR2_X1 U13074 ( .A(P3_REG3_REG_21__SCAN_IN), .B(keyinput37), .ZN(n10390)
         );
  NAND2_X1 U13075 ( .A1(n10391), .A2(n10390), .ZN(n10392) );
  NOR4_X1 U13076 ( .A1(n10395), .A2(n10394), .A3(n10393), .A4(n10392), .ZN(
        n10422) );
  INV_X1 U13077 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n10397) );
  AOI22_X1 U13078 ( .A1(n10397), .A2(keyinput35), .B1(keyinput1), .B2(n8828), 
        .ZN(n10396) );
  OAI221_X1 U13079 ( .B1(n10397), .B2(keyinput35), .C1(n8828), .C2(keyinput1), 
        .A(n10396), .ZN(n10407) );
  AOI22_X1 U13080 ( .A1(n14691), .A2(keyinput116), .B1(n11887), .B2(keyinput70), .ZN(n10398) );
  OAI221_X1 U13081 ( .B1(n14691), .B2(keyinput116), .C1(n11887), .C2(
        keyinput70), .A(n10398), .ZN(n10399) );
  INV_X1 U13082 ( .A(n10399), .ZN(n10401) );
  XNOR2_X1 U13083 ( .A(SI_0_), .B(keyinput126), .ZN(n10400) );
  NAND2_X1 U13084 ( .A1(n10401), .A2(n10400), .ZN(n10406) );
  AOI22_X1 U13085 ( .A1(n10403), .A2(keyinput57), .B1(keyinput40), .B2(n14644), 
        .ZN(n10402) );
  OAI221_X1 U13086 ( .B1(n10403), .B2(keyinput57), .C1(n14644), .C2(keyinput40), .A(n10402), .ZN(n10405) );
  INV_X1 U13087 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n15727) );
  XNOR2_X1 U13088 ( .A(n15727), .B(keyinput44), .ZN(n10404) );
  NOR4_X1 U13089 ( .A1(n10407), .A2(n10406), .A3(n10405), .A4(n10404), .ZN(
        n10421) );
  AOI22_X1 U13090 ( .A1(n10410), .A2(keyinput75), .B1(keyinput46), .B2(n10409), 
        .ZN(n10408) );
  OAI221_X1 U13091 ( .B1(n10410), .B2(keyinput75), .C1(n10409), .C2(keyinput46), .A(n10408), .ZN(n10419) );
  AOI22_X1 U13092 ( .A1(n10412), .A2(keyinput84), .B1(n13983), .B2(keyinput112), .ZN(n10411) );
  OAI221_X1 U13093 ( .B1(n10412), .B2(keyinput84), .C1(n13983), .C2(
        keyinput112), .A(n10411), .ZN(n10418) );
  XOR2_X1 U13094 ( .A(n8840), .B(keyinput41), .Z(n10416) );
  XOR2_X1 U13095 ( .A(n8243), .B(keyinput69), .Z(n10415) );
  XNOR2_X1 U13096 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput17), .ZN(n10414) );
  XNOR2_X1 U13097 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput109), .ZN(n10413) );
  NAND4_X1 U13098 ( .A1(n10416), .A2(n10415), .A3(n10414), .A4(n10413), .ZN(
        n10417) );
  NOR3_X1 U13099 ( .A1(n10419), .A2(n10418), .A3(n10417), .ZN(n10420) );
  NAND4_X1 U13100 ( .A1(n10423), .A2(n10422), .A3(n10421), .A4(n10420), .ZN(
        n10472) );
  INV_X1 U13101 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n12582) );
  AOI22_X1 U13102 ( .A1(n9487), .A2(keyinput121), .B1(keyinput27), .B2(n12582), 
        .ZN(n10424) );
  OAI221_X1 U13103 ( .B1(n9487), .B2(keyinput121), .C1(n12582), .C2(keyinput27), .A(n10424), .ZN(n10433) );
  AOI22_X1 U13104 ( .A1(n11083), .A2(keyinput89), .B1(n11177), .B2(keyinput30), 
        .ZN(n10425) );
  OAI221_X1 U13105 ( .B1(n11083), .B2(keyinput89), .C1(n11177), .C2(keyinput30), .A(n10425), .ZN(n10432) );
  INV_X1 U13106 ( .A(P3_DATAO_REG_20__SCAN_IN), .ZN(n10933) );
  AOI22_X1 U13107 ( .A1(n10933), .A2(keyinput92), .B1(n10427), .B2(keyinput110), .ZN(n10426) );
  OAI221_X1 U13108 ( .B1(n10933), .B2(keyinput92), .C1(n10427), .C2(
        keyinput110), .A(n10426), .ZN(n10431) );
  XNOR2_X1 U13109 ( .A(P3_REG1_REG_2__SCAN_IN), .B(keyinput123), .ZN(n10429)
         );
  XNOR2_X1 U13110 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(keyinput19), .ZN(n10428)
         );
  NAND2_X1 U13111 ( .A1(n10429), .A2(n10428), .ZN(n10430) );
  NOR4_X1 U13112 ( .A1(n10433), .A2(n10432), .A3(n10431), .A4(n10430), .ZN(
        n10470) );
  AOI22_X1 U13113 ( .A1(n11519), .A2(keyinput72), .B1(keyinput85), .B2(n15682), 
        .ZN(n10434) );
  OAI221_X1 U13114 ( .B1(n11519), .B2(keyinput72), .C1(n15682), .C2(keyinput85), .A(n10434), .ZN(n10443) );
  AOI22_X1 U13115 ( .A1(n15092), .A2(keyinput7), .B1(n10818), .B2(keyinput76), 
        .ZN(n10435) );
  OAI221_X1 U13116 ( .B1(n15092), .B2(keyinput7), .C1(n10818), .C2(keyinput76), 
        .A(n10435), .ZN(n10442) );
  NAND2_X1 U13117 ( .A1(n13900), .A2(keyinput52), .ZN(n10436) );
  OAI221_X1 U13118 ( .B1(n10437), .B2(keyinput73), .C1(n13900), .C2(keyinput52), .A(n10436), .ZN(n10441) );
  XNOR2_X1 U13119 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput39), .ZN(n10439)
         );
  XNOR2_X1 U13120 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput3), .ZN(n10438) );
  NAND2_X1 U13121 ( .A1(n10439), .A2(n10438), .ZN(n10440) );
  NOR4_X1 U13122 ( .A1(n10443), .A2(n10442), .A3(n10441), .A4(n10440), .ZN(
        n10469) );
  INV_X1 U13123 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n15797) );
  AOI22_X1 U13124 ( .A1(n13868), .A2(keyinput9), .B1(keyinput54), .B2(n15797), 
        .ZN(n10444) );
  OAI221_X1 U13125 ( .B1(n13868), .B2(keyinput9), .C1(n15797), .C2(keyinput54), 
        .A(n10444), .ZN(n10455) );
  INV_X1 U13126 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n10446) );
  AOI22_X1 U13127 ( .A1(n10757), .A2(keyinput115), .B1(keyinput97), .B2(n10446), .ZN(n10445) );
  OAI221_X1 U13128 ( .B1(n10757), .B2(keyinput115), .C1(n10446), .C2(
        keyinput97), .A(n10445), .ZN(n10454) );
  INV_X1 U13129 ( .A(SI_11_), .ZN(n10449) );
  AOI22_X1 U13130 ( .A1(n10449), .A2(keyinput127), .B1(keyinput87), .B2(n10448), .ZN(n10447) );
  OAI221_X1 U13131 ( .B1(n10449), .B2(keyinput127), .C1(n10448), .C2(
        keyinput87), .A(n10447), .ZN(n10453) );
  XNOR2_X1 U13132 ( .A(P3_IR_REG_13__SCAN_IN), .B(keyinput117), .ZN(n10451) );
  XNOR2_X1 U13133 ( .A(P1_REG1_REG_26__SCAN_IN), .B(keyinput62), .ZN(n10450)
         );
  NAND2_X1 U13134 ( .A1(n10451), .A2(n10450), .ZN(n10452) );
  NOR4_X1 U13135 ( .A1(n10455), .A2(n10454), .A3(n10453), .A4(n10452), .ZN(
        n10468) );
  AOI22_X1 U13136 ( .A1(n10760), .A2(keyinput22), .B1(keyinput51), .B2(n8146), 
        .ZN(n10456) );
  OAI221_X1 U13137 ( .B1(n10760), .B2(keyinput22), .C1(n8146), .C2(keyinput51), 
        .A(n10456), .ZN(n10466) );
  AOI22_X1 U13138 ( .A1(n10458), .A2(keyinput53), .B1(n11480), .B2(keyinput36), 
        .ZN(n10457) );
  OAI221_X1 U13139 ( .B1(n10458), .B2(keyinput53), .C1(n11480), .C2(keyinput36), .A(n10457), .ZN(n10465) );
  AOI22_X1 U13140 ( .A1(n10890), .A2(keyinput15), .B1(keyinput38), .B2(n10460), 
        .ZN(n10459) );
  OAI221_X1 U13141 ( .B1(n10890), .B2(keyinput15), .C1(n10460), .C2(keyinput38), .A(n10459), .ZN(n10464) );
  XNOR2_X1 U13142 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput86), .ZN(n10462)
         );
  XNOR2_X1 U13143 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput13), .ZN(n10461) );
  NAND2_X1 U13144 ( .A1(n10462), .A2(n10461), .ZN(n10463) );
  NOR4_X1 U13145 ( .A1(n10466), .A2(n10465), .A3(n10464), .A4(n10463), .ZN(
        n10467) );
  NAND4_X1 U13146 ( .A1(n10470), .A2(n10469), .A3(n10468), .A4(n10467), .ZN(
        n10471) );
  NOR4_X1 U13147 ( .A1(n10474), .A2(n10473), .A3(n10472), .A4(n10471), .ZN(
        n10475) );
  OAI21_X1 U13148 ( .B1(n10477), .B2(n10476), .A(n10475), .ZN(n10480) );
  MUX2_X1 U13149 ( .A(n10478), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(n10479) );
  XNOR2_X1 U13150 ( .A(n10480), .B(n10479), .ZN(P1_U3355) );
  NOR2_X1 U13151 ( .A1(n10481), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14028) );
  INV_X2 U13152 ( .A(n14028), .ZN(n14040) );
  NAND2_X2 U13153 ( .A1(n10481), .A2(P3_U3151), .ZN(n14033) );
  OAI222_X1 U13154 ( .A1(n10484), .A2(P3_U3151), .B1(n14040), .B2(n10483), 
        .C1(n10482), .C2(n14033), .ZN(P3_U3289) );
  INV_X1 U13155 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10486) );
  OAI222_X1 U13156 ( .A1(n13196), .A2(n10486), .B1(n12667), .B2(n10485), .C1(
        P2_U3088), .C2(n10658), .ZN(P2_U3320) );
  OAI222_X1 U13157 ( .A1(n10488), .A2(P1_U3086), .B1(n15546), .B2(n10487), 
        .C1(n10985), .C2(n10594), .ZN(P1_U3354) );
  INV_X1 U13158 ( .A(n10489), .ZN(n10495) );
  INV_X1 U13159 ( .A(n10771), .ZN(n15018) );
  OAI222_X1 U13160 ( .A1(n15546), .A2(n10490), .B1(n10985), .B2(n10495), .C1(
        n15018), .C2(P1_U3086), .ZN(P1_U3347) );
  OAI222_X1 U13161 ( .A1(n15546), .A2(n10491), .B1(n10985), .B2(n6626), .C1(
        n10582), .C2(P1_U3086), .ZN(P1_U3353) );
  INV_X1 U13162 ( .A(n12667), .ZN(n13079) );
  INV_X1 U13163 ( .A(n13079), .ZN(n13198) );
  INV_X1 U13164 ( .A(n10730), .ZN(n10624) );
  OAI222_X1 U13165 ( .A1(n13196), .A2(n10493), .B1(n13198), .B2(n10492), .C1(
        P2_U3088), .C2(n10624), .ZN(P2_U3321) );
  OAI222_X1 U13166 ( .A1(n13196), .A2(n10494), .B1(n13198), .B2(n6626), .C1(
        P2_U3088), .C2(n14262), .ZN(P2_U3325) );
  INV_X1 U13167 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10496) );
  INV_X1 U13168 ( .A(n10717), .ZN(n10684) );
  OAI222_X1 U13169 ( .A1(n13196), .A2(n10496), .B1(n13198), .B2(n10495), .C1(
        P2_U3088), .C2(n10684), .ZN(P2_U3319) );
  INV_X1 U13170 ( .A(n10651), .ZN(n15805) );
  OAI222_X1 U13171 ( .A1(n13196), .A2(n10498), .B1(n13198), .B2(n10497), .C1(
        P2_U3088), .C2(n15805), .ZN(P2_U3323) );
  OAI222_X1 U13172 ( .A1(P3_U3151), .A2(n11317), .B1(n14033), .B2(n10500), 
        .C1(n14040), .C2(n10499), .ZN(P3_U3286) );
  OAI222_X1 U13173 ( .A1(P3_U3151), .A2(n11145), .B1(n14033), .B2(n10502), 
        .C1(n14040), .C2(n10501), .ZN(P3_U3288) );
  OAI222_X1 U13174 ( .A1(P3_U3151), .A2(n10505), .B1(n14033), .B2(n10504), 
        .C1(n14040), .C2(n10503), .ZN(P3_U3285) );
  INV_X1 U13175 ( .A(SI_8_), .ZN(n10508) );
  INV_X1 U13176 ( .A(n10506), .ZN(n10507) );
  OAI222_X1 U13177 ( .A1(P3_U3151), .A2(n10509), .B1(n14033), .B2(n10508), 
        .C1(n14040), .C2(n10507), .ZN(P3_U3287) );
  INV_X1 U13178 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10512) );
  INV_X1 U13179 ( .A(n10510), .ZN(n10513) );
  INV_X1 U13180 ( .A(n10804), .ZN(n10511) );
  OAI222_X1 U13181 ( .A1(n13196), .A2(n10512), .B1(n13198), .B2(n10513), .C1(
        P2_U3088), .C2(n10511), .ZN(P2_U3318) );
  OAI222_X1 U13182 ( .A1(n15546), .A2(n10514), .B1(n10985), .B2(n10513), .C1(
        n10773), .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U13183 ( .A(n10515), .ZN(n10517) );
  INV_X1 U13184 ( .A(SI_2_), .ZN(n10516) );
  OAI222_X1 U13185 ( .A1(n11391), .A2(P3_U3151), .B1(n14040), .B2(n10517), 
        .C1(n10516), .C2(n14033), .ZN(P3_U3293) );
  OAI222_X1 U13186 ( .A1(n11295), .A2(P3_U3151), .B1(n14040), .B2(n10519), 
        .C1(n10518), .C2(n14033), .ZN(P3_U3294) );
  INV_X1 U13187 ( .A(n10520), .ZN(n10522) );
  INV_X1 U13188 ( .A(SI_3_), .ZN(n10521) );
  OAI222_X1 U13189 ( .A1(n10523), .A2(P3_U3151), .B1(n14040), .B2(n10522), 
        .C1(n10521), .C2(n14033), .ZN(P3_U3292) );
  INV_X1 U13190 ( .A(n10524), .ZN(n10526) );
  INV_X1 U13191 ( .A(SI_4_), .ZN(n10525) );
  OAI222_X1 U13192 ( .A1(n11697), .A2(P3_U3151), .B1(n14040), .B2(n10526), 
        .C1(n10525), .C2(n14033), .ZN(P3_U3291) );
  INV_X1 U13193 ( .A(n10527), .ZN(n10529) );
  INV_X1 U13194 ( .A(SI_5_), .ZN(n10528) );
  OAI222_X1 U13195 ( .A1(n10530), .A2(P3_U3151), .B1(n14040), .B2(n10529), 
        .C1(n10528), .C2(n14033), .ZN(P3_U3290) );
  OAI222_X1 U13196 ( .A1(P3_U3151), .A2(n11964), .B1(n14033), .B2(n10449), 
        .C1(n14040), .C2(n10531), .ZN(P3_U3284) );
  NAND2_X1 U13197 ( .A1(n10554), .A2(n10532), .ZN(n10550) );
  NAND2_X1 U13198 ( .A1(n10533), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n10536) );
  INV_X1 U13199 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10534) );
  NAND2_X1 U13200 ( .A1(n10534), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n10535) );
  NAND2_X1 U13201 ( .A1(n10550), .A2(n10549), .ZN(n10548) );
  NAND2_X1 U13202 ( .A1(n10548), .A2(n10536), .ZN(n10537) );
  NAND2_X1 U13203 ( .A1(n10539), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n10540) );
  NAND2_X1 U13204 ( .A1(n10544), .A2(n10540), .ZN(n10541) );
  NAND2_X1 U13205 ( .A1(n10541), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n10936) );
  NAND2_X1 U13206 ( .A1(n10542), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n10543) );
  INV_X1 U13207 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10545) );
  XNOR2_X1 U13208 ( .A(n10566), .B(n10545), .ZN(n15978) );
  NAND2_X1 U13209 ( .A1(n10547), .A2(n10546), .ZN(n15980) );
  OAI21_X1 U13210 ( .B1(n10550), .B2(n10549), .A(n10548), .ZN(n10559) );
  NAND2_X1 U13211 ( .A1(n10552), .A2(n10551), .ZN(n10553) );
  NAND2_X1 U13212 ( .A1(n10554), .A2(n10553), .ZN(n10555) );
  NAND2_X1 U13213 ( .A1(n10555), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n10557) );
  XOR2_X1 U13214 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10555), .Z(n15982) );
  NAND2_X1 U13215 ( .A1(n15983), .A2(n15982), .ZN(n10556) );
  NAND2_X1 U13216 ( .A1(n10557), .A2(n10556), .ZN(n10558) );
  NAND2_X1 U13217 ( .A1(n10559), .A2(n10558), .ZN(n15627) );
  INV_X1 U13218 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n15629) );
  NAND2_X1 U13219 ( .A1(n15627), .A2(n15629), .ZN(n10560) );
  OR2_X1 U13220 ( .A1(n10559), .A2(n10558), .ZN(n15628) );
  NAND2_X1 U13221 ( .A1(n10560), .A2(n15628), .ZN(n10563) );
  INV_X1 U13222 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10561) );
  NAND2_X1 U13223 ( .A1(n10563), .A2(n10561), .ZN(n10562) );
  NAND2_X1 U13224 ( .A1(n15980), .A2(n10562), .ZN(n10565) );
  INV_X1 U13225 ( .A(n10563), .ZN(n15979) );
  NAND2_X1 U13226 ( .A1(n15979), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n10564) );
  NAND2_X1 U13227 ( .A1(n10565), .A2(n10564), .ZN(n15977) );
  AND2_X1 U13228 ( .A1(n10566), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n10567) );
  NAND2_X1 U13229 ( .A1(n10568), .A2(n10569), .ZN(n10934) );
  INV_X1 U13230 ( .A(n10569), .ZN(n10570) );
  INV_X1 U13231 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10677) );
  OAI21_X1 U13232 ( .B1(n6790), .B2(n10677), .A(n10935), .ZN(SUB_1596_U58) );
  INV_X1 U13233 ( .A(n10572), .ZN(n10611) );
  AOI22_X1 U13234 ( .A1(n15037), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10679), .ZN(n10573) );
  OAI21_X1 U13235 ( .B1(n10611), .B2(n10985), .A(n10573), .ZN(P1_U3345) );
  NOR2_X1 U13236 ( .A1(n10582), .A2(n9487), .ZN(n14978) );
  INV_X1 U13237 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10574) );
  MUX2_X1 U13238 ( .A(n10574), .B(P1_REG1_REG_3__SCAN_IN), .S(n14977), .Z(
        n10575) );
  INV_X1 U13239 ( .A(n14977), .ZN(n10586) );
  NAND2_X1 U13240 ( .A1(n10586), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n14994) );
  INV_X1 U13241 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n15795) );
  MUX2_X1 U13242 ( .A(n15795), .B(P1_REG1_REG_4__SCAN_IN), .S(n10588), .Z(
        n14993) );
  MUX2_X1 U13243 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n15797), .S(n10602), .Z(
        n10576) );
  OAI21_X1 U13244 ( .B1(n10577), .B2(n10576), .A(n10596), .ZN(n10581) );
  NAND2_X1 U13245 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n11033) );
  NAND2_X1 U13246 ( .A1(n15651), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n10578) );
  OAI211_X1 U13247 ( .C1(n15659), .C2(n10579), .A(n11033), .B(n10578), .ZN(
        n10580) );
  AOI21_X1 U13248 ( .B1(n10581), .B2(n15108), .A(n10580), .ZN(n10593) );
  XNOR2_X1 U13249 ( .A(n10602), .B(n11204), .ZN(n10591) );
  INV_X1 U13250 ( .A(n10582), .ZN(n10583) );
  NAND2_X1 U13251 ( .A1(n10583), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n10584) );
  NAND2_X1 U13252 ( .A1(n10585), .A2(n10584), .ZN(n14975) );
  MUX2_X1 U13253 ( .A(n15713), .B(P1_REG2_REG_3__SCAN_IN), .S(n14977), .Z(
        n14976) );
  NAND2_X1 U13254 ( .A1(n14975), .A2(n14976), .ZN(n14974) );
  NAND2_X1 U13255 ( .A1(n10586), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n10587) );
  NAND2_X1 U13256 ( .A1(n14974), .A2(n10587), .ZN(n14991) );
  MUX2_X1 U13257 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n9526), .S(n10588), .Z(
        n14992) );
  NAND2_X1 U13258 ( .A1(n14991), .A2(n14992), .ZN(n14990) );
  NAND2_X1 U13259 ( .A1(n10588), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10589) );
  NAND2_X1 U13260 ( .A1(n14990), .A2(n10589), .ZN(n10590) );
  NAND2_X1 U13261 ( .A1(n10590), .A2(n10591), .ZN(n10604) );
  OAI211_X1 U13262 ( .C1(n10591), .C2(n10590), .A(n15665), .B(n10604), .ZN(
        n10592) );
  NAND2_X1 U13263 ( .A1(n10593), .A2(n10592), .ZN(P1_U3248) );
  OAI222_X1 U13264 ( .A1(P2_U3088), .A2(n14250), .B1(n13196), .B2(n10595), 
        .C1(n13198), .C2(n10594), .ZN(P2_U3326) );
  MUX2_X1 U13265 ( .A(n15001), .B(P1_REG1_REG_6__SCAN_IN), .S(n15007), .Z(
        n10597) );
  NAND2_X1 U13266 ( .A1(n15007), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10599) );
  MUX2_X1 U13267 ( .A(n15800), .B(P1_REG1_REG_7__SCAN_IN), .S(n10768), .Z(
        n10598) );
  NAND3_X1 U13268 ( .A1(n15002), .A2(n10599), .A3(n10598), .ZN(n10600) );
  NAND2_X1 U13269 ( .A1(n10600), .A2(n15108), .ZN(n10610) );
  INV_X1 U13270 ( .A(n15659), .ZN(n15085) );
  INV_X1 U13271 ( .A(n15651), .ZN(n15668) );
  INV_X1 U13272 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10950) );
  NAND2_X1 U13273 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n11998) );
  OAI21_X1 U13274 ( .B1(n15668), .B2(n10950), .A(n11998), .ZN(n10601) );
  AOI21_X1 U13275 ( .B1(n10768), .B2(n15085), .A(n10601), .ZN(n10609) );
  MUX2_X1 U13276 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n9595), .S(n10768), .Z(
        n10607) );
  NAND2_X1 U13277 ( .A1(n10602), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10603) );
  NAND2_X1 U13278 ( .A1(n10604), .A2(n10603), .ZN(n15009) );
  XNOR2_X1 U13279 ( .A(n15007), .B(n11355), .ZN(n15010) );
  NAND2_X1 U13280 ( .A1(n15009), .A2(n15010), .ZN(n15008) );
  NAND2_X1 U13281 ( .A1(n15007), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10605) );
  NAND2_X1 U13282 ( .A1(n15008), .A2(n10605), .ZN(n10606) );
  NAND2_X1 U13283 ( .A1(n10606), .A2(n10607), .ZN(n10770) );
  OAI211_X1 U13284 ( .C1(n10607), .C2(n10606), .A(n15665), .B(n10770), .ZN(
        n10608) );
  OAI211_X1 U13285 ( .C1(n10762), .C2(n10610), .A(n10609), .B(n10608), .ZN(
        P1_U3250) );
  INV_X1 U13286 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10612) );
  OAI222_X1 U13287 ( .A1(n13196), .A2(n10612), .B1(n13198), .B2(n10611), .C1(
        P2_U3088), .C2(n10807), .ZN(P2_U3317) );
  INV_X1 U13288 ( .A(n10613), .ZN(n10619) );
  AOI22_X1 U13289 ( .A1(n11441), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n10679), .ZN(n10614) );
  OAI21_X1 U13290 ( .B1(n10619), .B2(n10985), .A(n10614), .ZN(P1_U3344) );
  INV_X1 U13291 ( .A(n10615), .ZN(n10616) );
  OAI222_X1 U13292 ( .A1(P3_U3151), .A2(n10618), .B1(n14033), .B2(n10617), 
        .C1(n14040), .C2(n10616), .ZN(P3_U3283) );
  INV_X1 U13293 ( .A(n10810), .ZN(n10895) );
  OAI222_X1 U13294 ( .A1(n13196), .A2(n10620), .B1(n12667), .B2(n10619), .C1(
        P2_U3088), .C2(n10895), .ZN(P2_U3316) );
  INV_X1 U13295 ( .A(n14250), .ZN(n10643) );
  MUX2_X1 U13296 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n8888), .S(n14250), .Z(
        n14245) );
  NAND2_X1 U13297 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n14246) );
  NOR2_X1 U13298 ( .A1(n14245), .A2(n14246), .ZN(n14244) );
  AOI21_X1 U13299 ( .B1(n10643), .B2(P2_REG1_REG_1__SCAN_IN), .A(n14244), .ZN(
        n14259) );
  INV_X1 U13300 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n15887) );
  MUX2_X1 U13301 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n15887), .S(n14262), .Z(
        n14258) );
  NOR2_X1 U13302 ( .A1(n14262), .A2(n15887), .ZN(n14271) );
  MUX2_X1 U13303 ( .A(n8828), .B(P2_REG1_REG_3__SCAN_IN), .S(n14277), .Z(
        n10621) );
  OAI21_X1 U13304 ( .B1(n14276), .B2(n14271), .A(n10621), .ZN(n14274) );
  MUX2_X1 U13305 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10622), .S(n10651), .Z(
        n15817) );
  NAND2_X1 U13306 ( .A1(n10651), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10667) );
  INV_X1 U13307 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n15891) );
  MUX2_X1 U13308 ( .A(n15891), .B(P2_REG1_REG_5__SCAN_IN), .S(n10674), .Z(
        n10666) );
  AOI21_X1 U13309 ( .B1(n10674), .B2(P2_REG1_REG_5__SCAN_IN), .A(n10665), .ZN(
        n10726) );
  XNOR2_X1 U13310 ( .A(n10730), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n10725) );
  XNOR2_X1 U13311 ( .A(n10658), .B(P2_REG1_REG_7__SCAN_IN), .ZN(n10681) );
  XNOR2_X1 U13312 ( .A(n10682), .B(n10681), .ZN(n10664) );
  NAND2_X1 U13313 ( .A1(n10625), .A2(n11455), .ZN(n10627) );
  NAND2_X1 U13314 ( .A1(n10627), .A2(n7327), .ZN(n10631) );
  INV_X1 U13315 ( .A(n10628), .ZN(n10629) );
  NAND2_X1 U13316 ( .A1(n11455), .A2(n10629), .ZN(n10630) );
  AND2_X1 U13317 ( .A1(n10631), .A2(n10630), .ZN(n10634) );
  INV_X1 U13318 ( .A(n10634), .ZN(n10640) );
  OR2_X1 U13319 ( .A1(n9282), .A2(P2_U3088), .ZN(n12284) );
  NOR2_X1 U13320 ( .A1(n12284), .A2(n10632), .ZN(n10633) );
  AND2_X1 U13321 ( .A1(n10634), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15809) );
  AND2_X1 U13322 ( .A1(n9282), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10635) );
  NAND2_X1 U13323 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n11672) );
  OAI21_X1 U13324 ( .B1(n15806), .B2(n10658), .A(n11672), .ZN(n10636) );
  AOI21_X1 U13325 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(n15809), .A(n10636), .ZN(
        n10663) );
  NOR2_X1 U13326 ( .A1(n10637), .A2(P2_U3088), .ZN(n12989) );
  AND2_X1 U13327 ( .A1(n10638), .A2(n12989), .ZN(n10639) );
  AND2_X1 U13328 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10642) );
  NAND2_X1 U13329 ( .A1(n10643), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10644) );
  INV_X1 U13330 ( .A(n14262), .ZN(n10646) );
  NAND2_X1 U13331 ( .A1(n10646), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n14280) );
  NAND2_X1 U13332 ( .A1(n14281), .A2(n14280), .ZN(n10648) );
  MUX2_X1 U13333 ( .A(n14278), .B(P2_REG2_REG_3__SCAN_IN), .S(n14277), .Z(
        n10647) );
  NAND2_X1 U13334 ( .A1(n10648), .A2(n10647), .ZN(n14283) );
  INV_X1 U13335 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n14278) );
  OR2_X1 U13336 ( .A1(n14277), .A2(n14278), .ZN(n10649) );
  NAND2_X1 U13337 ( .A1(n14283), .A2(n10649), .ZN(n15812) );
  MUX2_X1 U13338 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10650), .S(n10651), .Z(
        n15813) );
  NAND2_X1 U13339 ( .A1(n15812), .A2(n15813), .ZN(n15810) );
  NAND2_X1 U13340 ( .A1(n10651), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10652) );
  NAND2_X1 U13341 ( .A1(n15810), .A2(n10652), .ZN(n10670) );
  MUX2_X1 U13342 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10653), .S(n10674), .Z(
        n10671) );
  NAND2_X1 U13343 ( .A1(n10670), .A2(n10671), .ZN(n10733) );
  NAND2_X1 U13344 ( .A1(n10674), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10732) );
  NAND2_X1 U13345 ( .A1(n10733), .A2(n10732), .ZN(n10655) );
  MUX2_X1 U13346 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11106), .S(n10730), .Z(
        n10654) );
  NAND2_X1 U13347 ( .A1(n10655), .A2(n10654), .ZN(n10735) );
  NAND2_X1 U13348 ( .A1(n10730), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10660) );
  NAND2_X1 U13349 ( .A1(n10735), .A2(n10660), .ZN(n10657) );
  MUX2_X1 U13350 ( .A(n11404), .B(P2_REG2_REG_7__SCAN_IN), .S(n10658), .Z(
        n10656) );
  NAND2_X1 U13351 ( .A1(n10657), .A2(n10656), .ZN(n10720) );
  MUX2_X1 U13352 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11404), .S(n10658), .Z(
        n10659) );
  NAND3_X1 U13353 ( .A1(n10735), .A2(n10660), .A3(n10659), .ZN(n10661) );
  NAND3_X1 U13354 ( .A1(n15811), .A2(n10720), .A3(n10661), .ZN(n10662) );
  OAI211_X1 U13355 ( .C1(n10664), .C2(n15825), .A(n10663), .B(n10662), .ZN(
        P2_U3221) );
  NOR2_X1 U13356 ( .A1(n15651), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U13357 ( .A(n10665), .ZN(n10669) );
  NAND3_X1 U13358 ( .A1(n15814), .A2(n10667), .A3(n10666), .ZN(n10668) );
  NAND3_X1 U13359 ( .A1(n10669), .A2(n15815), .A3(n10668), .ZN(n10676) );
  NAND2_X1 U13360 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n11234) );
  OAI211_X1 U13361 ( .C1(n10671), .C2(n10670), .A(n15811), .B(n10733), .ZN(
        n10672) );
  NAND2_X1 U13362 ( .A1(n11234), .A2(n10672), .ZN(n10673) );
  AOI21_X1 U13363 ( .B1(n15831), .B2(n10674), .A(n10673), .ZN(n10675) );
  OAI211_X1 U13364 ( .C1(n10677), .C2(n15840), .A(n10676), .B(n10675), .ZN(
        P2_U3219) );
  INV_X1 U13365 ( .A(n10678), .ZN(n10706) );
  AOI22_X1 U13366 ( .A1(n11471), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n10679), .ZN(n10680) );
  OAI21_X1 U13367 ( .B1(n10706), .B2(n10985), .A(n10680), .ZN(P1_U3343) );
  XNOR2_X1 U13368 ( .A(n10804), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n10686) );
  XNOR2_X1 U13369 ( .A(n10717), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n10712) );
  INV_X1 U13370 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10683) );
  OAI22_X1 U13371 ( .A1(n10713), .A2(n10712), .B1(n10684), .B2(n10683), .ZN(
        n10685) );
  NOR2_X1 U13372 ( .A1(n10685), .A2(n10686), .ZN(n15823) );
  AOI21_X1 U13373 ( .B1(n10686), .B2(n10685), .A(n15823), .ZN(n10701) );
  AND2_X1 U13374 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n12145) );
  INV_X1 U13375 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10687) );
  NOR2_X1 U13376 ( .A1(n15840), .A2(n10687), .ZN(n10688) );
  AOI211_X1 U13377 ( .C1(n15831), .C2(n10804), .A(n12145), .B(n10688), .ZN(
        n10700) );
  NAND2_X1 U13378 ( .A1(n10689), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10719) );
  NAND2_X1 U13379 ( .A1(n10720), .A2(n10719), .ZN(n10692) );
  MUX2_X1 U13380 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10690), .S(n10717), .Z(
        n10691) );
  NAND2_X1 U13381 ( .A1(n10692), .A2(n10691), .ZN(n10722) );
  NAND2_X1 U13382 ( .A1(n10717), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10693) );
  NAND2_X1 U13383 ( .A1(n10722), .A2(n10693), .ZN(n10695) );
  INV_X1 U13384 ( .A(n10695), .ZN(n10697) );
  MUX2_X1 U13385 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n11367), .S(n10804), .Z(
        n10696) );
  MUX2_X1 U13386 ( .A(n11367), .B(P2_REG2_REG_9__SCAN_IN), .S(n10804), .Z(
        n10694) );
  OAI21_X1 U13387 ( .B1(n10697), .B2(n10696), .A(n10806), .ZN(n10698) );
  NAND2_X1 U13388 ( .A1(n10698), .A2(n15811), .ZN(n10699) );
  OAI211_X1 U13389 ( .C1(n10701), .C2(n15825), .A(n10700), .B(n10699), .ZN(
        P2_U3223) );
  INV_X1 U13390 ( .A(n10702), .ZN(n10704) );
  OAI222_X1 U13391 ( .A1(n13196), .A2(n10703), .B1(n12667), .B2(n10704), .C1(
        n11535), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U13392 ( .A(n11482), .ZN(n11475) );
  OAI222_X1 U13393 ( .A1(n15546), .A2(n10705), .B1(n10985), .B2(n10704), .C1(
        P1_U3086), .C2(n11475), .ZN(P1_U3342) );
  INV_X1 U13394 ( .A(n11005), .ZN(n10900) );
  OAI222_X1 U13395 ( .A1(n13196), .A2(n10707), .B1(n12667), .B2(n10706), .C1(
        n10900), .C2(P2_U3088), .ZN(P2_U3315) );
  INV_X1 U13396 ( .A(n10708), .ZN(n10710) );
  INV_X1 U13397 ( .A(n15070), .ZN(n15062) );
  OAI222_X1 U13398 ( .A1(n15546), .A2(n10709), .B1(n10985), .B2(n10710), .C1(
        P1_U3086), .C2(n15062), .ZN(P1_U3339) );
  INV_X1 U13399 ( .A(n12198), .ZN(n11975) );
  OAI222_X1 U13400 ( .A1(n13196), .A2(n10711), .B1(n12667), .B2(n10710), .C1(
        n11975), .C2(P2_U3088), .ZN(P2_U3311) );
  NAND2_X1 U13401 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n11912) );
  XOR2_X1 U13402 ( .A(n10713), .B(n10712), .Z(n10714) );
  NAND2_X1 U13403 ( .A1(n15815), .A2(n10714), .ZN(n10715) );
  NAND2_X1 U13404 ( .A1(n11912), .A2(n10715), .ZN(n10716) );
  AOI21_X1 U13405 ( .B1(n15831), .B2(n10717), .A(n10716), .ZN(n10724) );
  MUX2_X1 U13406 ( .A(n10690), .B(P2_REG2_REG_8__SCAN_IN), .S(n10717), .Z(
        n10718) );
  NAND3_X1 U13407 ( .A1(n10720), .A2(n10719), .A3(n10718), .ZN(n10721) );
  NAND3_X1 U13408 ( .A1(n10722), .A2(n15811), .A3(n10721), .ZN(n10723) );
  OAI211_X1 U13409 ( .C1(n15840), .C2(n7356), .A(n10724), .B(n10723), .ZN(
        P2_U3222) );
  NAND2_X1 U13410 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n11248) );
  XOR2_X1 U13411 ( .A(n10726), .B(n10725), .Z(n10727) );
  NAND2_X1 U13412 ( .A1(n15815), .A2(n10727), .ZN(n10728) );
  NAND2_X1 U13413 ( .A1(n11248), .A2(n10728), .ZN(n10729) );
  AOI21_X1 U13414 ( .B1(n15831), .B2(n10730), .A(n10729), .ZN(n10737) );
  MUX2_X1 U13415 ( .A(n11106), .B(P2_REG2_REG_6__SCAN_IN), .S(n10730), .Z(
        n10731) );
  NAND3_X1 U13416 ( .A1(n10733), .A2(n10732), .A3(n10731), .ZN(n10734) );
  NAND3_X1 U13417 ( .A1(n15811), .A2(n10735), .A3(n10734), .ZN(n10736) );
  OAI211_X1 U13418 ( .C1(n15840), .C2(n10311), .A(n10737), .B(n10736), .ZN(
        P2_U3220) );
  INV_X1 U13419 ( .A(n14930), .ZN(n14918) );
  NAND2_X1 U13420 ( .A1(n15632), .A2(n10738), .ZN(n12728) );
  NAND2_X1 U13421 ( .A1(n11057), .A2(n15636), .ZN(n11297) );
  INV_X1 U13422 ( .A(n11297), .ZN(n10792) );
  AOI22_X1 U13423 ( .A1(n12728), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n15641), 
        .B2(n10792), .ZN(n10741) );
  NAND2_X1 U13424 ( .A1(n10739), .A2(n14910), .ZN(n10740) );
  OAI211_X1 U13425 ( .C1(n14918), .C2(n11298), .A(n10741), .B(n10740), .ZN(
        P1_U3232) );
  OAI222_X1 U13426 ( .A1(P3_U3151), .A2(n10744), .B1(n14033), .B2(n10743), 
        .C1(n14040), .C2(n10742), .ZN(P3_U3282) );
  NAND2_X1 U13427 ( .A1(n15811), .A2(n10747), .ZN(n10745) );
  OAI211_X1 U13428 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n15825), .A(n10745), .B(
        n15806), .ZN(n10749) );
  INV_X1 U13429 ( .A(n15811), .ZN(n15832) );
  OAI22_X1 U13430 ( .A1(n15832), .A2(n10747), .B1(n10746), .B2(n15825), .ZN(
        n10748) );
  MUX2_X1 U13431 ( .A(n10749), .B(n10748), .S(n14252), .Z(n10751) );
  OAI22_X1 U13432 ( .A1(n15840), .A2(n10210), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15842), .ZN(n10750) );
  OR2_X1 U13433 ( .A1(n10751), .A2(n10750), .ZN(P2_U3214) );
  INV_X1 U13434 ( .A(n10752), .ZN(n10753) );
  OAI222_X1 U13435 ( .A1(P3_U3151), .A2(n7380), .B1(n14033), .B2(n10754), .C1(
        n14040), .C2(n10753), .ZN(P3_U3280) );
  INV_X1 U13436 ( .A(n9723), .ZN(n10756) );
  INV_X1 U13437 ( .A(n11979), .ZN(n11661) );
  OAI222_X1 U13438 ( .A1(n13196), .A2(n10755), .B1(n12667), .B2(n10756), .C1(
        P2_U3088), .C2(n11661), .ZN(P2_U3312) );
  INV_X1 U13439 ( .A(n15053), .ZN(n15660) );
  OAI222_X1 U13440 ( .A1(n15546), .A2(n10757), .B1(n10985), .B2(n10756), .C1(
        n15660), .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U13441 ( .A(n10758), .ZN(n10761) );
  INV_X1 U13442 ( .A(n15086), .ZN(n15080) );
  OAI222_X1 U13443 ( .A1(n15546), .A2(n10759), .B1(n10985), .B2(n10761), .C1(
        P1_U3086), .C2(n15080), .ZN(P1_U3338) );
  INV_X1 U13444 ( .A(n12341), .ZN(n11976) );
  OAI222_X1 U13445 ( .A1(P2_U3088), .A2(n11976), .B1(n12667), .B2(n10761), 
        .C1(n10760), .C2(n13196), .ZN(P2_U3310) );
  MUX2_X1 U13446 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9609), .S(n10771), .Z(
        n15014) );
  XNOR2_X1 U13447 ( .A(n10773), .B(n10763), .ZN(n10764) );
  AOI21_X1 U13448 ( .B1(n10765), .B2(n10764), .A(n15030), .ZN(n10779) );
  NOR2_X1 U13449 ( .A1(n10766), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14854) );
  NOR2_X1 U13450 ( .A1(n15659), .A2(n10773), .ZN(n10767) );
  AOI211_X1 U13451 ( .C1(n15651), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n14854), .B(
        n10767), .ZN(n10778) );
  NAND2_X1 U13452 ( .A1(n10768), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10769) );
  NAND2_X1 U13453 ( .A1(n10770), .A2(n10769), .ZN(n15022) );
  XNOR2_X1 U13454 ( .A(n10771), .B(n15682), .ZN(n15023) );
  NAND2_X1 U13455 ( .A1(n15022), .A2(n15023), .ZN(n15021) );
  NAND2_X1 U13456 ( .A1(n10771), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10772) );
  NAND2_X1 U13457 ( .A1(n15021), .A2(n10772), .ZN(n10776) );
  INV_X1 U13458 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10774) );
  MUX2_X1 U13459 ( .A(n10774), .B(P1_REG2_REG_9__SCAN_IN), .S(n10773), .Z(
        n10775) );
  NAND2_X1 U13460 ( .A1(n10776), .A2(n10775), .ZN(n10919) );
  OAI211_X1 U13461 ( .C1(n10776), .C2(n10775), .A(n10919), .B(n15665), .ZN(
        n10777) );
  OAI211_X1 U13462 ( .C1(n10779), .C2(n15661), .A(n10778), .B(n10777), .ZN(
        P1_U3252) );
  OAI222_X1 U13463 ( .A1(P3_U3151), .A2(n10782), .B1(n14033), .B2(n10781), 
        .C1(n14040), .C2(n10780), .ZN(P3_U3281) );
  AND2_X1 U13464 ( .A1(n10817), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U13465 ( .A1(n10817), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U13466 ( .A1(n10817), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U13467 ( .A1(n10817), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U13468 ( .A1(n10817), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U13469 ( .A1(n10817), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U13470 ( .A1(n10817), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U13471 ( .A1(n10817), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U13472 ( .A1(n10817), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U13473 ( .A1(n10817), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U13474 ( .A1(n10817), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U13475 ( .A1(n10817), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U13476 ( .A1(n10817), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U13477 ( .A1(n10817), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U13478 ( .A1(n10817), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U13479 ( .A1(n10817), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U13480 ( .A1(n10817), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U13481 ( .A1(n10817), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U13482 ( .A1(n10817), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U13483 ( .A1(n10817), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U13484 ( .A1(n10817), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U13485 ( .A1(n10817), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U13486 ( .A1(n10817), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U13487 ( .A1(n10817), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U13488 ( .A1(n10817), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U13489 ( .A1(n10817), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U13490 ( .A1(n10817), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  INV_X1 U13491 ( .A(n10784), .ZN(n10786) );
  INV_X1 U13492 ( .A(n11653), .ZN(n11656) );
  OAI222_X1 U13493 ( .A1(n13196), .A2(n10785), .B1(n12667), .B2(n10786), .C1(
        n11656), .C2(P2_U3088), .ZN(P2_U3313) );
  INV_X1 U13494 ( .A(n15050), .ZN(n15044) );
  OAI222_X1 U13495 ( .A1(n15546), .A2(n10787), .B1(n10985), .B2(n10786), .C1(
        P1_U3086), .C2(n15044), .ZN(P1_U3341) );
  INV_X1 U13496 ( .A(n11066), .ZN(n10793) );
  INV_X1 U13497 ( .A(n11298), .ZN(n11058) );
  NAND2_X1 U13498 ( .A1(n12438), .A2(n6809), .ZN(n10788) );
  NAND2_X1 U13499 ( .A1(n10789), .A2(n10788), .ZN(n11301) );
  INV_X1 U13500 ( .A(n15553), .ZN(n12410) );
  NAND2_X1 U13501 ( .A1(n12410), .A2(n11065), .ZN(n12618) );
  NAND2_X1 U13502 ( .A1(n9977), .A2(n12622), .ZN(n12588) );
  NOR2_X1 U13503 ( .A1(n14958), .A2(n11298), .ZN(n11164) );
  INV_X1 U13504 ( .A(n11164), .ZN(n12441) );
  NAND2_X1 U13505 ( .A1(n14958), .A2(n11298), .ZN(n12439) );
  NAND2_X1 U13506 ( .A1(n12441), .A2(n12439), .ZN(n12633) );
  INV_X1 U13507 ( .A(n12633), .ZN(n10790) );
  AOI21_X1 U13508 ( .B1(n15760), .B2(n15709), .A(n10790), .ZN(n10791) );
  AOI211_X1 U13509 ( .C1(n10793), .C2(n11058), .A(n10792), .B(n10791), .ZN(
        n15731) );
  OAI21_X1 U13510 ( .B1(n10795), .B2(P1_D_REG_1__SCAN_IN), .A(n10794), .ZN(
        n10799) );
  NAND2_X1 U13511 ( .A1(n10797), .A2(n10796), .ZN(n10798) );
  NOR2_X1 U13512 ( .A1(n15517), .A2(n11059), .ZN(n10800) );
  INV_X1 U13513 ( .A(n15804), .ZN(n15802) );
  NAND2_X1 U13514 ( .A1(n15802), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10801) );
  OAI21_X1 U13515 ( .B1(n15731), .B2(n15802), .A(n10801), .ZN(P1_U3528) );
  NOR2_X1 U13516 ( .A1(n10804), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n15822) );
  XNOR2_X1 U13517 ( .A(n15830), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n15827) );
  XNOR2_X1 U13518 ( .A(n10810), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n10896) );
  XNOR2_X1 U13519 ( .A(n10897), .B(n10896), .ZN(n10816) );
  NOR2_X1 U13520 ( .A1(n10802), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14174) );
  NOR2_X1 U13521 ( .A1(n15806), .A2(n10895), .ZN(n10803) );
  AOI211_X1 U13522 ( .C1(n15809), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n14174), 
        .B(n10803), .ZN(n10815) );
  OR2_X1 U13523 ( .A1(n10810), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10903) );
  OR2_X1 U13524 ( .A1(n10895), .A2(n9013), .ZN(n10809) );
  OR2_X1 U13525 ( .A1(n10804), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n10805) );
  NAND2_X1 U13526 ( .A1(n10806), .A2(n10805), .ZN(n15834) );
  MUX2_X1 U13527 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n8996), .S(n10807), .Z(
        n15833) );
  NAND2_X1 U13528 ( .A1(n15830), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10808) );
  AOI21_X1 U13529 ( .B1(n10903), .B2(n10809), .A(n10812), .ZN(n10813) );
  MUX2_X1 U13530 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n9013), .S(n10810), .Z(
        n10811) );
  OAI21_X1 U13531 ( .B1(n10813), .B2(n6776), .A(n15811), .ZN(n10814) );
  OAI211_X1 U13532 ( .C1(n10816), .C2(n15825), .A(n10815), .B(n10814), .ZN(
        P2_U3225) );
  INV_X1 U13533 ( .A(n10817), .ZN(n10821) );
  NOR2_X1 U13534 ( .A1(n10821), .A2(n10818), .ZN(P3_U3257) );
  NOR2_X1 U13535 ( .A1(n10821), .A2(n10819), .ZN(P3_U3254) );
  NOR2_X1 U13536 ( .A1(n10821), .A2(n10820), .ZN(P3_U3240) );
  INV_X1 U13537 ( .A(n13693), .ZN(n13699) );
  INV_X1 U13538 ( .A(n10822), .ZN(n10823) );
  OAI222_X1 U13539 ( .A1(P3_U3151), .A2(n13699), .B1(n14033), .B2(n10824), 
        .C1(n14040), .C2(n10823), .ZN(P3_U3279) );
  XNOR2_X1 U13540 ( .A(n10826), .B(n10825), .ZN(n10827) );
  NAND2_X1 U13541 ( .A1(n10827), .A2(n14910), .ZN(n10830) );
  INV_X1 U13542 ( .A(n14957), .ZN(n10828) );
  INV_X1 U13543 ( .A(n11057), .ZN(n11072) );
  OAI22_X1 U13544 ( .A1(n10828), .A2(n14913), .B1(n11072), .B2(n14922), .ZN(
        n11166) );
  AOI22_X1 U13545 ( .A1(n12728), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n11166), 
        .B2(n15641), .ZN(n10829) );
  OAI211_X1 U13546 ( .C1(n15743), .C2(n14918), .A(n10830), .B(n10829), .ZN(
        P1_U3237) );
  NAND2_X1 U13547 ( .A1(n10832), .A2(n10831), .ZN(n10838) );
  OAI21_X1 U13548 ( .B1(n10838), .B2(n15863), .A(n10842), .ZN(n10835) );
  AND2_X1 U13549 ( .A1(n10834), .A2(n10833), .ZN(n12990) );
  NAND2_X1 U13550 ( .A1(n10835), .A2(n12990), .ZN(n11015) );
  NOR2_X1 U13551 ( .A1(n11015), .A2(P2_U3088), .ZN(n10889) );
  NAND2_X2 U13552 ( .A1(n6554), .A2(n12987), .ZN(n14508) );
  INV_X1 U13553 ( .A(n15863), .ZN(n11090) );
  NAND2_X1 U13554 ( .A1(n11090), .A2(n15864), .ZN(n10837) );
  AND2_X1 U13555 ( .A1(n15879), .A2(n10839), .ZN(n10840) );
  AOI21_X1 U13556 ( .B1(n14243), .B2(n14508), .A(n14213), .ZN(n10845) );
  INV_X1 U13557 ( .A(n10841), .ZN(n11097) );
  NAND2_X1 U13558 ( .A1(n10847), .A2(n11097), .ZN(n10844) );
  OAI21_X1 U13559 ( .B1(n10845), .B2(n14211), .A(n11158), .ZN(n10851) );
  NAND2_X1 U13560 ( .A1(n12775), .A2(n14193), .ZN(n10875) );
  INV_X1 U13561 ( .A(n10875), .ZN(n10849) );
  INV_X1 U13562 ( .A(n12931), .ZN(n10846) );
  AND2_X1 U13563 ( .A1(n14243), .A2(n12770), .ZN(n10873) );
  AND3_X1 U13564 ( .A1(n14161), .A2(n10873), .A3(n14508), .ZN(n10848) );
  AOI21_X1 U13565 ( .B1(n10849), .B2(n14206), .A(n10848), .ZN(n10850) );
  OAI211_X1 U13566 ( .C1(n10889), .C2(n15842), .A(n10851), .B(n10850), .ZN(
        P2_U3204) );
  NAND2_X1 U13567 ( .A1(P3_U3897), .A2(n12672), .ZN(n10852) );
  OAI21_X1 U13568 ( .B1(P3_U3897), .B2(n10853), .A(n10852), .ZN(P3_U3506) );
  NAND2_X1 U13569 ( .A1(P3_U3897), .A2(n11777), .ZN(n10854) );
  OAI21_X1 U13570 ( .B1(P3_U3897), .B2(n10855), .A(n10854), .ZN(P3_U3492) );
  NAND2_X1 U13571 ( .A1(n12987), .A2(n12763), .ZN(n10856) );
  NAND2_X1 U13572 ( .A1(n14508), .A2(n12775), .ZN(n10859) );
  INV_X1 U13573 ( .A(n10859), .ZN(n10858) );
  XNOR2_X1 U13574 ( .A(n13166), .B(n12009), .ZN(n10860) );
  INV_X1 U13575 ( .A(n10860), .ZN(n10857) );
  INV_X1 U13576 ( .A(n10881), .ZN(n10861) );
  AOI21_X1 U13577 ( .B1(n10863), .B2(n10862), .A(n10861), .ZN(n10869) );
  NAND2_X1 U13578 ( .A1(n14243), .A2(n14192), .ZN(n10865) );
  NAND2_X1 U13579 ( .A1(n14242), .A2(n14193), .ZN(n10864) );
  NAND2_X1 U13580 ( .A1(n10865), .A2(n10864), .ZN(n11156) );
  AOI22_X1 U13581 ( .A1(n14206), .A2(n11156), .B1(n14211), .B2(n6553), .ZN(
        n10868) );
  INV_X1 U13582 ( .A(n10889), .ZN(n10866) );
  NAND2_X1 U13583 ( .A1(n10866), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n10867) );
  OAI211_X1 U13584 ( .C1(n10869), .C2(n14213), .A(n10868), .B(n10867), .ZN(
        P2_U3194) );
  INV_X1 U13585 ( .A(n13700), .ZN(n13712) );
  INV_X1 U13586 ( .A(n10870), .ZN(n10872) );
  OAI222_X1 U13587 ( .A1(n13712), .A2(P3_U3151), .B1(n14040), .B2(n10872), 
        .C1(n10871), .C2(n14033), .ZN(P3_U3278) );
  OR2_X1 U13588 ( .A1(n10873), .A2(n11154), .ZN(n15848) );
  NOR2_X1 U13589 ( .A1(n12770), .A2(n9291), .ZN(n15841) );
  INV_X1 U13590 ( .A(n14552), .ZN(n12163) );
  OAI21_X1 U13591 ( .B1(n12163), .B2(n14556), .A(n15848), .ZN(n10876) );
  NAND2_X1 U13592 ( .A1(n10876), .A2(n10875), .ZN(n15846) );
  AOI211_X1 U13593 ( .C1(n15877), .C2(n15848), .A(n15841), .B(n15846), .ZN(
        n15865) );
  INV_X1 U13594 ( .A(n15893), .ZN(n15890) );
  NAND2_X1 U13595 ( .A1(n15890), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10877) );
  OAI21_X1 U13596 ( .B1(n15865), .B2(n15890), .A(n10877), .ZN(P2_U3499) );
  XNOR2_X1 U13597 ( .A(n13166), .B(n15867), .ZN(n10879) );
  NAND2_X1 U13598 ( .A1(n14508), .A2(n14242), .ZN(n10878) );
  NAND2_X1 U13599 ( .A1(n10879), .A2(n10878), .ZN(n11018) );
  OR2_X1 U13600 ( .A1(n10879), .A2(n10878), .ZN(n10880) );
  AND2_X1 U13601 ( .A1(n11018), .A2(n10880), .ZN(n10883) );
  NAND2_X1 U13602 ( .A1(n10882), .A2(n10883), .ZN(n11019) );
  OAI21_X1 U13603 ( .B1(n10883), .B2(n10882), .A(n11019), .ZN(n10884) );
  NAND2_X1 U13604 ( .A1(n10884), .A2(n14161), .ZN(n10888) );
  NAND2_X1 U13605 ( .A1(n14241), .A2(n14193), .ZN(n10886) );
  NAND2_X1 U13606 ( .A1(n12775), .A2(n14192), .ZN(n10885) );
  NAND2_X1 U13607 ( .A1(n10886), .A2(n10885), .ZN(n11703) );
  AOI22_X1 U13608 ( .A1(n14206), .A2(n11703), .B1(n14211), .B2(n12784), .ZN(
        n10887) );
  OAI211_X1 U13609 ( .C1(n10889), .C2(n14261), .A(n10888), .B(n10887), .ZN(
        P2_U3209) );
  INV_X1 U13610 ( .A(n15089), .ZN(n15099) );
  OAI222_X1 U13611 ( .A1(n15546), .A2(n10890), .B1(n10985), .B2(n10892), .C1(
        P1_U3086), .C2(n15099), .ZN(P1_U3337) );
  INV_X1 U13612 ( .A(n14289), .ZN(n10893) );
  OAI222_X1 U13613 ( .A1(P2_U3088), .A2(n10893), .B1(n12667), .B2(n10892), 
        .C1(n10891), .C2(n13196), .ZN(P2_U3309) );
  XNOR2_X1 U13614 ( .A(n11005), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n10899) );
  INV_X1 U13615 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10894) );
  NOR2_X1 U13616 ( .A1(n10898), .A2(n10899), .ZN(n11002) );
  AOI21_X1 U13617 ( .B1(n10899), .B2(n10898), .A(n11002), .ZN(n10910) );
  NAND2_X1 U13618 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n14094)
         );
  OAI21_X1 U13619 ( .B1(n15806), .B2(n10900), .A(n14094), .ZN(n10901) );
  AOI21_X1 U13620 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(n15809), .A(n10901), 
        .ZN(n10909) );
  INV_X1 U13621 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10902) );
  MUX2_X1 U13622 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n10902), .S(n11005), .Z(
        n10904) );
  NOR3_X1 U13623 ( .A1(n6776), .A2(n10904), .A3(n7055), .ZN(n10907) );
  NAND2_X1 U13624 ( .A1(n10905), .A2(n10904), .ZN(n11007) );
  INV_X1 U13625 ( .A(n11007), .ZN(n10906) );
  OAI21_X1 U13626 ( .B1(n10907), .B2(n10906), .A(n15811), .ZN(n10908) );
  OAI211_X1 U13627 ( .C1(n10910), .C2(n15825), .A(n10909), .B(n10908), .ZN(
        P2_U3226) );
  OR2_X1 U13628 ( .A1(n11441), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n11435) );
  NAND2_X1 U13629 ( .A1(n11441), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10911) );
  NAND2_X1 U13630 ( .A1(n11435), .A2(n10911), .ZN(n10914) );
  NOR2_X1 U13631 ( .A1(n10917), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n15029) );
  XNOR2_X1 U13632 ( .A(n15037), .B(P1_REG1_REG_10__SCAN_IN), .ZN(n15028) );
  OR2_X1 U13633 ( .A1(n15027), .A2(n10912), .ZN(n10913) );
  AOI21_X1 U13634 ( .B1(n10914), .B2(n10913), .A(n11437), .ZN(n10925) );
  NOR2_X1 U13635 ( .A1(n10915), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14897) );
  INV_X1 U13636 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n12275) );
  NOR2_X1 U13637 ( .A1(n15668), .A2(n12275), .ZN(n10916) );
  AOI211_X1 U13638 ( .C1(n15085), .C2(n11441), .A(n14897), .B(n10916), .ZN(
        n10924) );
  NAND2_X1 U13639 ( .A1(n10917), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10918) );
  NAND2_X1 U13640 ( .A1(n10919), .A2(n10918), .ZN(n15036) );
  XNOR2_X1 U13641 ( .A(n15037), .B(n12210), .ZN(n15035) );
  NAND2_X1 U13642 ( .A1(n15036), .A2(n15035), .ZN(n15034) );
  NAND2_X1 U13643 ( .A1(n15037), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10920) );
  NAND2_X1 U13644 ( .A1(n15034), .A2(n10920), .ZN(n10922) );
  XNOR2_X1 U13645 ( .A(n11441), .B(n11955), .ZN(n10921) );
  NAND2_X1 U13646 ( .A1(n10922), .A2(n10921), .ZN(n11443) );
  OAI211_X1 U13647 ( .C1(n10922), .C2(n10921), .A(n11443), .B(n15665), .ZN(
        n10923) );
  OAI211_X1 U13648 ( .C1(n10925), .C2(n15661), .A(n10924), .B(n10923), .ZN(
        P1_U3254) );
  INV_X1 U13649 ( .A(n13725), .ZN(n13724) );
  INV_X1 U13650 ( .A(n10926), .ZN(n10927) );
  OAI222_X1 U13651 ( .A1(P3_U3151), .A2(n13724), .B1(n14033), .B2(n10928), 
        .C1(n14040), .C2(n10927), .ZN(P3_U3277) );
  OAI222_X1 U13652 ( .A1(n14040), .A2(n10930), .B1(n14033), .B2(n10929), .C1(
        P3_U3151), .C2(n13745), .ZN(P3_U3276) );
  OAI222_X1 U13653 ( .A1(P1_U3086), .A2(n11065), .B1(n10985), .B2(n12408), 
        .C1(n10931), .C2(n15546), .ZN(P1_U3335) );
  INV_X1 U13654 ( .A(n13849), .ZN(n13252) );
  NAND2_X1 U13655 ( .A1(n13252), .A2(P3_U3897), .ZN(n10932) );
  OAI21_X1 U13656 ( .B1(P3_U3897), .B2(n10933), .A(n10932), .ZN(P3_U3511) );
  NAND2_X1 U13657 ( .A1(n10937), .A2(n10936), .ZN(n10946) );
  XNOR2_X1 U13658 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n10938) );
  XNOR2_X1 U13659 ( .A(n10946), .B(n10938), .ZN(n15555) );
  NAND2_X1 U13660 ( .A1(n15554), .A2(n15555), .ZN(n10942) );
  INV_X1 U13661 ( .A(n10939), .ZN(n10940) );
  NAND2_X1 U13662 ( .A1(n10940), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n10941) );
  INV_X1 U13663 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10943) );
  INV_X1 U13664 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n10944) );
  NAND2_X1 U13665 ( .A1(n10944), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n10945) );
  NAND2_X1 U13666 ( .A1(n10946), .A2(n10945), .ZN(n10948) );
  NAND2_X1 U13667 ( .A1(n15004), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n10947) );
  INV_X1 U13668 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n10949) );
  XNOR2_X1 U13669 ( .A(n10954), .B(n10949), .ZN(n10953) );
  XNOR2_X1 U13670 ( .A(n10953), .B(n10950), .ZN(n15557) );
  NAND2_X1 U13671 ( .A1(n10951), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n10952) );
  NAND2_X1 U13672 ( .A1(n10953), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n10956) );
  INV_X1 U13673 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n10957) );
  NAND2_X1 U13674 ( .A1(n10957), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n11718) );
  INV_X1 U13675 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10958) );
  NAND2_X1 U13676 ( .A1(n10958), .A2(P3_ADDR_REG_8__SCAN_IN), .ZN(n10959) );
  INV_X1 U13677 ( .A(n11716), .ZN(n10960) );
  NAND2_X1 U13678 ( .A1(n10963), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n10964) );
  NAND2_X1 U13679 ( .A1(n11715), .A2(n10964), .ZN(SUB_1596_U55) );
  INV_X1 U13680 ( .A(n10965), .ZN(n11707) );
  INV_X1 U13681 ( .A(n11558), .ZN(n10966) );
  AOI211_X1 U13682 ( .C1(n12791), .C2(n11707), .A(n14635), .B(n10966), .ZN(
        n11328) );
  NAND2_X1 U13683 ( .A1(n11153), .A2(n10967), .ZN(n11702) );
  XNOR2_X1 U13684 ( .A(n14242), .B(n12784), .ZN(n12960) );
  NAND2_X1 U13685 ( .A1(n11702), .A2(n12960), .ZN(n11701) );
  NAND3_X1 U13686 ( .A1(n11701), .A2(n12965), .A3(n10968), .ZN(n10971) );
  NAND2_X1 U13687 ( .A1(n10970), .A2(n10969), .ZN(n11551) );
  AND2_X1 U13688 ( .A1(n10971), .A2(n11551), .ZN(n10974) );
  NAND2_X1 U13689 ( .A1(n14240), .A2(n14193), .ZN(n10973) );
  NAND2_X1 U13690 ( .A1(n14242), .A2(n14192), .ZN(n10972) );
  AND2_X1 U13691 ( .A1(n10973), .A2(n10972), .ZN(n11017) );
  OAI21_X1 U13692 ( .B1(n10974), .B2(n14534), .A(n11017), .ZN(n11324) );
  AOI211_X1 U13693 ( .C1(n12791), .C2(n10017), .A(n11328), .B(n11324), .ZN(
        n10982) );
  NAND2_X1 U13694 ( .A1(n11151), .A2(n10975), .ZN(n11700) );
  INV_X1 U13695 ( .A(n12960), .ZN(n11699) );
  NAND2_X1 U13696 ( .A1(n11700), .A2(n11699), .ZN(n11698) );
  NAND3_X1 U13697 ( .A1(n11698), .A2(n10977), .A3(n10976), .ZN(n10979) );
  NAND2_X1 U13698 ( .A1(n10979), .A2(n10978), .ZN(n11323) );
  INV_X1 U13699 ( .A(n14734), .ZN(n11419) );
  AOI22_X1 U13700 ( .A1(n11323), .A2(n11419), .B1(n15885), .B2(
        P2_REG0_REG_3__SCAN_IN), .ZN(n10980) );
  OAI21_X1 U13701 ( .B1(n10982), .B2(n15885), .A(n10980), .ZN(P2_U3439) );
  INV_X1 U13702 ( .A(n14651), .ZN(n11417) );
  AOI22_X1 U13703 ( .A1(n11323), .A2(n11417), .B1(n15890), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n10981) );
  OAI21_X1 U13704 ( .B1(n10982), .B2(n15890), .A(n10981), .ZN(P2_U3502) );
  INV_X1 U13705 ( .A(n10983), .ZN(n12666) );
  OAI222_X1 U13706 ( .A1(n15314), .A2(P1_U3086), .B1(n10985), .B2(n12666), 
        .C1(n10984), .C2(n15546), .ZN(P1_U3336) );
  INV_X1 U13707 ( .A(n13836), .ZN(n13811) );
  NAND2_X1 U13708 ( .A1(n13811), .A2(P3_U3897), .ZN(n10986) );
  OAI21_X1 U13709 ( .B1(P3_U3897), .B2(n10987), .A(n10986), .ZN(P3_U3512) );
  INV_X1 U13710 ( .A(n11028), .ZN(n10994) );
  INV_X1 U13711 ( .A(n10989), .ZN(n10991) );
  NAND2_X1 U13712 ( .A1(n10991), .A2(n10990), .ZN(n10993) );
  AOI22_X1 U13713 ( .A1(n10994), .A2(n10988), .B1(n10993), .B2(n10992), .ZN(
        n11000) );
  NAND2_X1 U13714 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n14987) );
  NAND2_X1 U13715 ( .A1(n6539), .A2(n15636), .ZN(n10996) );
  NAND2_X1 U13716 ( .A1(n14957), .A2(n15637), .ZN(n10995) );
  NAND2_X1 U13717 ( .A1(n10996), .A2(n10995), .ZN(n15755) );
  NAND2_X1 U13718 ( .A1(n15641), .A2(n15755), .ZN(n10997) );
  OAI211_X1 U13719 ( .C1(n15646), .C2(n11427), .A(n14987), .B(n10997), .ZN(
        n10998) );
  AOI21_X1 U13720 ( .B1(n14930), .B2(n15756), .A(n10998), .ZN(n10999) );
  OAI21_X1 U13721 ( .B1(n11000), .B2(n15634), .A(n10999), .ZN(P1_U3230) );
  XOR2_X1 U13722 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n11535), .Z(n11004) );
  NOR2_X1 U13723 ( .A1(n11005), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n11001) );
  OR2_X1 U13724 ( .A1(n11002), .A2(n11001), .ZN(n11003) );
  AOI211_X1 U13725 ( .C1(n11004), .C2(n11003), .A(n15825), .B(n11538), .ZN(
        n11014) );
  OR2_X1 U13726 ( .A1(n11005), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n11006) );
  NAND2_X1 U13727 ( .A1(n11007), .A2(n11006), .ZN(n11010) );
  MUX2_X1 U13728 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n14539), .S(n11535), .Z(
        n11009) );
  INV_X1 U13729 ( .A(n11537), .ZN(n11008) );
  AOI211_X1 U13730 ( .C1(n11010), .C2(n11009), .A(n15832), .B(n11008), .ZN(
        n11013) );
  NAND2_X1 U13731 ( .A1(n15809), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n11011) );
  NAND2_X1 U13732 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n14156)
         );
  OAI211_X1 U13733 ( .C1(n15806), .C2(n11535), .A(n11011), .B(n14156), .ZN(
        n11012) );
  OR3_X1 U13734 ( .A1(n11014), .A2(n11013), .A3(n11012), .ZN(P2_U3227) );
  NAND2_X1 U13735 ( .A1(n14211), .A2(n12791), .ZN(n11016) );
  NAND2_X1 U13736 ( .A1(P2_U3088), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n14269) );
  OAI211_X1 U13737 ( .C1(n11017), .C2(n14196), .A(n11016), .B(n14269), .ZN(
        n11022) );
  NAND2_X1 U13738 ( .A1(n11019), .A2(n11018), .ZN(n11038) );
  NAND2_X1 U13739 ( .A1(n14508), .A2(n14241), .ZN(n11040) );
  XNOR2_X1 U13740 ( .A(n11039), .B(n11040), .ZN(n11037) );
  XNOR2_X1 U13741 ( .A(n11038), .B(n11037), .ZN(n11020) );
  NOR2_X1 U13742 ( .A1(n11020), .A2(n14213), .ZN(n11021) );
  AOI211_X1 U13743 ( .C1(n14194), .C2(n11023), .A(n11022), .B(n11021), .ZN(
        n11024) );
  INV_X1 U13744 ( .A(n11024), .ZN(P2_U3190) );
  INV_X1 U13745 ( .A(n15632), .ZN(n14901) );
  NAND2_X1 U13746 ( .A1(n12459), .A2(n15757), .ZN(n15765) );
  XNOR2_X1 U13747 ( .A(n11026), .B(n11025), .ZN(n11027) );
  XNOR2_X1 U13748 ( .A(n11028), .B(n11027), .ZN(n11029) );
  NAND2_X1 U13749 ( .A1(n11029), .A2(n14910), .ZN(n11036) );
  OR2_X1 U13750 ( .A1(n12418), .A2(n14913), .ZN(n11031) );
  NAND2_X1 U13751 ( .A1(n6540), .A2(n15637), .ZN(n11030) );
  NAND2_X1 U13752 ( .A1(n11031), .A2(n11030), .ZN(n11199) );
  NAND2_X1 U13753 ( .A1(n15641), .A2(n11199), .ZN(n11032) );
  OAI211_X1 U13754 ( .C1(n15646), .C2(n11203), .A(n11033), .B(n11032), .ZN(
        n11034) );
  INV_X1 U13755 ( .A(n11034), .ZN(n11035) );
  OAI211_X1 U13756 ( .C1(n14901), .C2(n15765), .A(n11036), .B(n11035), .ZN(
        P1_U3227) );
  INV_X1 U13757 ( .A(n14211), .ZN(n14171) );
  INV_X1 U13758 ( .A(n11040), .ZN(n11041) );
  NAND2_X1 U13759 ( .A1(n11042), .A2(n11041), .ZN(n11043) );
  XNOR2_X1 U13760 ( .A(n12795), .B(n13166), .ZN(n11044) );
  AND2_X1 U13761 ( .A1(n14508), .A2(n14240), .ZN(n11045) );
  NAND2_X1 U13762 ( .A1(n11044), .A2(n11045), .ZN(n11048) );
  INV_X1 U13763 ( .A(n11044), .ZN(n11047) );
  INV_X1 U13764 ( .A(n11045), .ZN(n11046) );
  NAND2_X1 U13765 ( .A1(n11047), .A2(n11046), .ZN(n11227) );
  OAI21_X1 U13766 ( .B1(n6783), .B2(n11049), .A(n11228), .ZN(n11050) );
  NAND2_X1 U13767 ( .A1(n11050), .A2(n14161), .ZN(n11056) );
  INV_X1 U13768 ( .A(n11559), .ZN(n11054) );
  AND2_X1 U13769 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n15808) );
  NAND2_X1 U13770 ( .A1(n14239), .A2(n14193), .ZN(n11052) );
  NAND2_X1 U13771 ( .A1(n14241), .A2(n14192), .ZN(n11051) );
  AND2_X1 U13772 ( .A1(n11052), .A2(n11051), .ZN(n11553) );
  NOR2_X1 U13773 ( .A1(n14196), .A2(n11553), .ZN(n11053) );
  AOI211_X1 U13774 ( .C1(n14194), .C2(n11054), .A(n15808), .B(n11053), .ZN(
        n11055) );
  OAI211_X1 U13775 ( .C1(n15873), .C2(n14171), .A(n11056), .B(n11055), .ZN(
        P2_U3202) );
  OR2_X1 U13776 ( .A1(n11057), .A2(n15732), .ZN(n12440) );
  NAND2_X1 U13777 ( .A1(n11057), .A2(n15732), .ZN(n12443) );
  NAND2_X1 U13778 ( .A1(n14958), .A2(n11058), .ZN(n11169) );
  XNOR2_X1 U13779 ( .A(n11170), .B(n11169), .ZN(n15737) );
  INV_X1 U13780 ( .A(n15737), .ZN(n11081) );
  INV_X1 U13781 ( .A(n15517), .ZN(n11061) );
  NAND3_X1 U13782 ( .A1(n11061), .A2(n11060), .A3(n11059), .ZN(n13035) );
  OR2_X1 U13783 ( .A1(n11064), .A2(n15314), .ZN(n12620) );
  NOR2_X1 U13784 ( .A1(n6546), .A2(n12620), .ZN(n15719) );
  INV_X1 U13785 ( .A(n15719), .ZN(n11360) );
  OR2_X1 U13786 ( .A1(n11066), .A2(n11065), .ZN(n11067) );
  OAI22_X1 U13787 ( .A1(n15714), .A2(n9458), .B1(n11068), .B2(n15712), .ZN(
        n11071) );
  NOR2_X2 U13788 ( .A1(n13035), .A2(n15112), .ZN(n15720) );
  NAND2_X1 U13789 ( .A1(n15720), .A2(n15678), .ZN(n15259) );
  OR2_X1 U13790 ( .A1(n15732), .A2(n11298), .ZN(n11069) );
  NAND2_X1 U13791 ( .A1(n11175), .A2(n11069), .ZN(n15734) );
  NOR2_X1 U13792 ( .A1(n15259), .A2(n15734), .ZN(n11070) );
  AOI211_X1 U13793 ( .C1(n15716), .C2(n11171), .A(n11071), .B(n11070), .ZN(
        n11080) );
  INV_X1 U13794 ( .A(n11170), .ZN(n11074) );
  XNOR2_X1 U13795 ( .A(n11072), .B(n15734), .ZN(n11073) );
  INV_X1 U13796 ( .A(n14958), .ZN(n11075) );
  MUX2_X1 U13797 ( .A(n11074), .B(n11073), .S(n11075), .Z(n11078) );
  INV_X1 U13798 ( .A(n15745), .ZN(n15711) );
  INV_X1 U13799 ( .A(n15638), .ZN(n11076) );
  OAI22_X1 U13800 ( .A1(n11076), .A2(n14913), .B1(n11075), .B2(n14922), .ZN(
        n12727) );
  AOI21_X1 U13801 ( .B1(n15737), .B2(n15711), .A(n12727), .ZN(n11077) );
  OAI21_X1 U13802 ( .B1(n15709), .B2(n11078), .A(n11077), .ZN(n15735) );
  NAND2_X1 U13803 ( .A1(n15735), .A2(n15714), .ZN(n11079) );
  OAI211_X1 U13804 ( .C1(n11081), .C2(n11360), .A(n11080), .B(n11079), .ZN(
        P1_U3292) );
  NAND2_X1 U13805 ( .A1(n13805), .A2(P3_U3897), .ZN(n11082) );
  OAI21_X1 U13806 ( .B1(P3_U3897), .B2(n11083), .A(n11082), .ZN(P3_U3513) );
  INV_X1 U13807 ( .A(n12967), .ZN(n11089) );
  OAI21_X1 U13808 ( .B1(n14238), .B2(n14675), .A(n11084), .ZN(n11088) );
  NAND2_X1 U13809 ( .A1(n11548), .A2(n11085), .ZN(n11789) );
  INV_X1 U13810 ( .A(n11789), .ZN(n11395) );
  OAI21_X1 U13811 ( .B1(n11789), .B2(n12800), .A(n15880), .ZN(n11086) );
  OAI21_X1 U13812 ( .B1(n11395), .B2(n14239), .A(n11086), .ZN(n11087) );
  MUX2_X1 U13813 ( .A(n11089), .B(n11088), .S(n11087), .Z(n14679) );
  AND2_X1 U13814 ( .A1(n11090), .A2(n15860), .ZN(n11091) );
  NAND2_X1 U13815 ( .A1(n11092), .A2(n11091), .ZN(n11093) );
  NAND2_X1 U13816 ( .A1(n14552), .A2(n12764), .ZN(n11094) );
  OAI21_X1 U13817 ( .B1(n11790), .B2(n11098), .A(n10836), .ZN(n11096) );
  NOR2_X1 U13818 ( .A1(n11096), .A2(n11095), .ZN(n14674) );
  NAND2_X1 U13819 ( .A1(n15850), .A2(n12987), .ZN(n14330) );
  OAI22_X1 U13820 ( .A1(n14563), .A2(n11098), .B1(n15843), .B2(n11246), .ZN(
        n11099) );
  AOI21_X1 U13821 ( .B1(n14674), .B2(n14567), .A(n11099), .ZN(n11108) );
  OAI21_X1 U13822 ( .B1(n12967), .B2(n11101), .A(n11100), .ZN(n11105) );
  OR2_X1 U13823 ( .A1(n12809), .A2(n14204), .ZN(n11103) );
  NAND2_X1 U13824 ( .A1(n14239), .A2(n14192), .ZN(n11102) );
  AND2_X1 U13825 ( .A1(n11103), .A2(n11102), .ZN(n11250) );
  INV_X1 U13826 ( .A(n11250), .ZN(n11104) );
  AOI21_X1 U13827 ( .B1(n11105), .B2(n14556), .A(n11104), .ZN(n14677) );
  MUX2_X1 U13828 ( .A(n14677), .B(n11106), .S(n14499), .Z(n11107) );
  OAI211_X1 U13829 ( .C1(n14679), .C2(n14546), .A(n11108), .B(n11107), .ZN(
        P2_U3259) );
  INV_X1 U13830 ( .A(n11109), .ZN(n11114) );
  OAI222_X1 U13831 ( .A1(n13196), .A2(n11111), .B1(n13198), .B2(n11114), .C1(
        P2_U3088), .C2(n11110), .ZN(P2_U3306) );
  OAI222_X1 U13832 ( .A1(n11112), .A2(P1_U3086), .B1(n10985), .B2(n11114), 
        .C1(n11113), .C2(n15546), .ZN(P1_U3334) );
  NAND2_X1 U13833 ( .A1(n6779), .A2(n11115), .ZN(n11116) );
  XNOR2_X1 U13834 ( .A(n11117), .B(n11116), .ZN(n11123) );
  OR2_X1 U13835 ( .A1(n12415), .A2(n14913), .ZN(n11119) );
  NAND2_X1 U13836 ( .A1(n6539), .A2(n15637), .ZN(n11118) );
  NAND2_X1 U13837 ( .A1(n11119), .A2(n11118), .ZN(n11340) );
  AOI22_X1 U13838 ( .A1(n15641), .A2(n11340), .B1(P1_REG3_REG_6__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11121) );
  NOR2_X1 U13839 ( .A1(n12417), .A2(n15742), .ZN(n15773) );
  NAND2_X1 U13840 ( .A1(n15632), .A2(n15773), .ZN(n11120) );
  OAI211_X1 U13841 ( .C1(n15646), .C2(n11354), .A(n11121), .B(n11120), .ZN(
        n11122) );
  AOI21_X1 U13842 ( .B1(n11123), .B2(n14910), .A(n11122), .ZN(n11124) );
  INV_X1 U13843 ( .A(n11124), .ZN(P1_U3239) );
  NAND2_X1 U13844 ( .A1(n11262), .A2(n15948), .ZN(n11255) );
  NOR2_X1 U13845 ( .A1(n15904), .A2(n13409), .ZN(n13532) );
  AOI21_X1 U13846 ( .B1(n15911), .B2(n11255), .A(n13532), .ZN(n11125) );
  AOI21_X1 U13847 ( .B1(n13886), .B2(n11777), .A(n11125), .ZN(n11241) );
  MUX2_X1 U13848 ( .A(n11241), .B(n8123), .S(n15960), .Z(n11126) );
  OAI21_X1 U13849 ( .B1(n11211), .B2(n14013), .A(n11126), .ZN(P3_U3390) );
  NOR2_X1 U13850 ( .A1(n14033), .A2(SI_22_), .ZN(n11127) );
  AOI21_X1 U13851 ( .B1(n11128), .B2(P3_STATE_REG_SCAN_IN), .A(n11127), .ZN(
        n11129) );
  OAI21_X1 U13852 ( .B1(n11130), .B2(n14040), .A(n11129), .ZN(n11131) );
  INV_X1 U13853 ( .A(n11131), .ZN(P3_U3273) );
  OAI222_X1 U13854 ( .A1(P2_U3088), .A2(n11134), .B1(n13198), .B2(n11133), 
        .C1(n11132), .C2(n13196), .ZN(P2_U3305) );
  NAND2_X1 U13855 ( .A1(n11136), .A2(n11135), .ZN(n11138) );
  OAI21_X1 U13856 ( .B1(n11623), .B2(n11138), .A(n11137), .ZN(n11142) );
  OAI21_X1 U13857 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n11140), .A(n11139), .ZN(
        n11141) );
  AOI22_X1 U13858 ( .A1(n11142), .A2(n13748), .B1(n13754), .B2(n11141), .ZN(
        n11149) );
  OAI21_X1 U13859 ( .B1(P3_REG2_REG_7__SCAN_IN), .B2(n11143), .A(n10172), .ZN(
        n11147) );
  AND2_X1 U13860 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n11828) );
  AOI21_X1 U13861 ( .B1(n15894), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11828), .ZN(
        n11144) );
  OAI21_X1 U13862 ( .B1(n13746), .B2(n11145), .A(n11144), .ZN(n11146) );
  AOI21_X1 U13863 ( .B1(n11147), .B2(n13667), .A(n11146), .ZN(n11148) );
  NAND2_X1 U13864 ( .A1(n11149), .A2(n11148), .ZN(P3_U3189) );
  INV_X1 U13865 ( .A(n11151), .ZN(n11152) );
  AOI21_X1 U13866 ( .B1(n7292), .B2(n12961), .A(n11152), .ZN(n12006) );
  OAI21_X1 U13867 ( .B1(n11154), .B2(n12961), .A(n11153), .ZN(n11157) );
  NOR2_X1 U13868 ( .A1(n12006), .A2(n14552), .ZN(n11155) );
  AOI211_X1 U13869 ( .C1(n14556), .C2(n11157), .A(n11156), .B(n11155), .ZN(
        n12015) );
  NAND2_X1 U13870 ( .A1(n11158), .A2(n6553), .ZN(n11159) );
  AND3_X1 U13871 ( .A1(n11159), .A2(n10836), .A3(n11706), .ZN(n12007) );
  AOI21_X1 U13872 ( .B1(n10017), .B2(n6553), .A(n12007), .ZN(n11160) );
  OAI211_X1 U13873 ( .C1(n12006), .C2(n14673), .A(n12015), .B(n11160), .ZN(
        n11162) );
  NAND2_X1 U13874 ( .A1(n11162), .A2(n15893), .ZN(n11161) );
  OAI21_X1 U13875 ( .B1(n15893), .B2(n8888), .A(n11161), .ZN(P2_U3500) );
  NAND2_X1 U13876 ( .A1(n11162), .A2(n15886), .ZN(n11163) );
  OAI21_X1 U13877 ( .B1(n15886), .B2(n8890), .A(n11163), .ZN(P2_U3433) );
  NAND2_X1 U13878 ( .A1(n11164), .A2(n12443), .ZN(n11165) );
  NAND2_X1 U13879 ( .A1(n15638), .A2(n15743), .ZN(n12434) );
  XNOR2_X1 U13880 ( .A(n12427), .B(n12634), .ZN(n11167) );
  AOI21_X1 U13881 ( .B1(n11167), .B2(n15763), .A(n11166), .ZN(n15741) );
  NOR2_X1 U13882 ( .A1(n6546), .A2(n15745), .ZN(n11168) );
  OR2_X1 U13883 ( .A1(n15719), .A2(n11168), .ZN(n11564) );
  NAND2_X1 U13884 ( .A1(n11170), .A2(n11169), .ZN(n11173) );
  OR2_X1 U13885 ( .A1(n11057), .A2(n11171), .ZN(n11172) );
  NAND2_X1 U13886 ( .A1(n11173), .A2(n11172), .ZN(n11185) );
  INV_X1 U13887 ( .A(n12634), .ZN(n11174) );
  XNOR2_X1 U13888 ( .A(n11185), .B(n11174), .ZN(n15744) );
  INV_X1 U13889 ( .A(n15744), .ZN(n11183) );
  NAND2_X1 U13890 ( .A1(n11186), .A2(n11175), .ZN(n11176) );
  NAND3_X1 U13891 ( .A1(n15718), .A2(n15678), .A3(n11176), .ZN(n15740) );
  NAND2_X1 U13892 ( .A1(n15716), .A2(n11186), .ZN(n11181) );
  NOR2_X1 U13893 ( .A1(n15712), .A2(n11178), .ZN(n11179) );
  AOI21_X1 U13894 ( .B1(n6546), .B2(P1_REG2_REG_2__SCAN_IN), .A(n11179), .ZN(
        n11180) );
  OAI211_X1 U13895 ( .C1(n15740), .C2(n15686), .A(n11181), .B(n11180), .ZN(
        n11182) );
  AOI21_X1 U13896 ( .B1(n11564), .B2(n11183), .A(n11182), .ZN(n11184) );
  OAI21_X1 U13897 ( .B1(n6546), .B2(n15741), .A(n11184), .ZN(P1_U3291) );
  XNOR2_X1 U13898 ( .A(n6539), .B(n12459), .ZN(n12636) );
  NAND2_X1 U13899 ( .A1(n11185), .A2(n12634), .ZN(n11188) );
  OR2_X1 U13900 ( .A1(n15638), .A2(n11186), .ZN(n11187) );
  NAND2_X1 U13901 ( .A1(n11188), .A2(n11187), .ZN(n15706) );
  NAND2_X1 U13902 ( .A1(n14957), .A2(n15631), .ZN(n12435) );
  NAND2_X1 U13903 ( .A1(n15706), .A2(n15708), .ZN(n11190) );
  OR2_X1 U13904 ( .A1(n14957), .A2(n7771), .ZN(n11189) );
  NAND2_X1 U13905 ( .A1(n11190), .A2(n11189), .ZN(n11423) );
  INV_X1 U13906 ( .A(n11423), .ZN(n11191) );
  AND2_X1 U13907 ( .A1(n6540), .A2(n15756), .ZN(n11334) );
  INV_X1 U13908 ( .A(n11334), .ZN(n11192) );
  NAND2_X1 U13909 ( .A1(n11337), .A2(n11192), .ZN(n11193) );
  NOR2_X1 U13910 ( .A1(n11193), .A2(n12636), .ZN(n11332) );
  AOI21_X1 U13911 ( .B1(n12636), .B2(n11193), .A(n11332), .ZN(n15766) );
  INV_X1 U13912 ( .A(n12636), .ZN(n11197) );
  INV_X1 U13913 ( .A(n15756), .ZN(n11431) );
  OR2_X1 U13914 ( .A1(n6540), .A2(n11431), .ZN(n11195) );
  NAND2_X1 U13915 ( .A1(n6540), .A2(n11431), .ZN(n11344) );
  NAND2_X1 U13916 ( .A1(n11347), .A2(n11344), .ZN(n11196) );
  NOR2_X1 U13917 ( .A1(n11196), .A2(n11197), .ZN(n11341) );
  AOI21_X1 U13918 ( .B1(n11197), .B2(n11196), .A(n11341), .ZN(n11202) );
  INV_X1 U13919 ( .A(n15766), .ZN(n11198) );
  NAND2_X1 U13920 ( .A1(n11198), .A2(n15711), .ZN(n11201) );
  INV_X1 U13921 ( .A(n11199), .ZN(n11200) );
  OAI211_X1 U13922 ( .C1(n11202), .C2(n15709), .A(n11201), .B(n11200), .ZN(
        n15768) );
  NAND2_X1 U13923 ( .A1(n15768), .A2(n15714), .ZN(n11208) );
  OAI22_X1 U13924 ( .A1(n15714), .A2(n11204), .B1(n11203), .B2(n15712), .ZN(
        n11206) );
  NOR2_X2 U13925 ( .A1(n15718), .A2(n7771), .ZN(n15717) );
  OAI211_X1 U13926 ( .C1(n11425), .C2(n11342), .A(n15678), .B(n11353), .ZN(
        n15764) );
  NOR2_X1 U13927 ( .A1(n15764), .A2(n15686), .ZN(n11205) );
  AOI211_X1 U13928 ( .C1(n15716), .C2(n12459), .A(n11206), .B(n11205), .ZN(
        n11207) );
  OAI211_X1 U13929 ( .C1(n15766), .C2(n11360), .A(n11208), .B(n11207), .ZN(
        P1_U3288) );
  INV_X1 U13930 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n11209) );
  MUX2_X1 U13931 ( .A(n11241), .B(n11209), .S(n15973), .Z(n11210) );
  OAI21_X1 U13932 ( .B1(n13940), .B2(n11211), .A(n11210), .ZN(P3_U3459) );
  INV_X1 U13933 ( .A(n11212), .ZN(n11215) );
  OAI222_X1 U13934 ( .A1(n14040), .A2(n11215), .B1(n14033), .B2(n11214), .C1(
        P3_U3151), .C2(n11213), .ZN(P3_U3275) );
  NOR3_X1 U13935 ( .A1(n13667), .A2(n13754), .A3(n13748), .ZN(n11221) );
  AOI21_X1 U13936 ( .B1(n11217), .B2(n11216), .A(n11284), .ZN(n11220) );
  AOI22_X1 U13937 ( .A1(n15894), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n11219) );
  OAI211_X1 U13938 ( .C1(n11221), .C2(n11220), .A(n11219), .B(n11218), .ZN(
        P3_U3182) );
  XNOR2_X1 U13939 ( .A(n12799), .B(n13166), .ZN(n11222) );
  AND2_X1 U13940 ( .A1(n14508), .A2(n14239), .ZN(n11223) );
  NAND2_X1 U13941 ( .A1(n11222), .A2(n11223), .ZN(n11226) );
  INV_X1 U13942 ( .A(n11222), .ZN(n11225) );
  INV_X1 U13943 ( .A(n11223), .ZN(n11224) );
  NAND2_X1 U13944 ( .A1(n11225), .A2(n11224), .ZN(n11244) );
  AND2_X1 U13945 ( .A1(n11226), .A2(n11244), .ZN(n11230) );
  OAI21_X1 U13946 ( .B1(n11230), .B2(n11229), .A(n11245), .ZN(n11238) );
  NOR2_X1 U13947 ( .A1(n14171), .A2(n15880), .ZN(n11237) );
  NAND2_X1 U13948 ( .A1(n14238), .A2(n14193), .ZN(n11232) );
  NAND2_X1 U13949 ( .A1(n14240), .A2(n14192), .ZN(n11231) );
  AND2_X1 U13950 ( .A1(n11232), .A2(n11231), .ZN(n11799) );
  INV_X1 U13951 ( .A(n11233), .ZN(n11793) );
  NAND2_X1 U13952 ( .A1(n14194), .A2(n11793), .ZN(n11235) );
  OAI211_X1 U13953 ( .C1(n11799), .C2(n14196), .A(n11235), .B(n11234), .ZN(
        n11236) );
  AOI211_X1 U13954 ( .C1(n11238), .C2(n14161), .A(n11237), .B(n11236), .ZN(
        n11239) );
  INV_X1 U13955 ( .A(n11239), .ZN(P2_U3199) );
  AOI22_X1 U13956 ( .A1(n13880), .A2(n11277), .B1(P3_REG3_REG_0__SCAN_IN), 
        .B2(n15901), .ZN(n11243) );
  MUX2_X1 U13957 ( .A(n11241), .B(n11240), .S(n15903), .Z(n11242) );
  NAND2_X1 U13958 ( .A1(n11243), .A2(n11242), .ZN(P3_U3233) );
  XNOR2_X1 U13959 ( .A(n14675), .B(n13166), .ZN(n11667) );
  AND2_X1 U13960 ( .A1(n14508), .A2(n14238), .ZN(n11666) );
  XNOR2_X1 U13961 ( .A(n11667), .B(n11666), .ZN(n11668) );
  XNOR2_X1 U13962 ( .A(n11669), .B(n11668), .ZN(n11253) );
  INV_X1 U13963 ( .A(n11246), .ZN(n11247) );
  NAND2_X1 U13964 ( .A1(n14194), .A2(n11247), .ZN(n11249) );
  OAI211_X1 U13965 ( .C1(n11250), .C2(n14196), .A(n11249), .B(n11248), .ZN(
        n11251) );
  AOI21_X1 U13966 ( .B1(n14675), .B2(n14211), .A(n11251), .ZN(n11252) );
  OAI21_X1 U13967 ( .B1(n11253), .B2(n14213), .A(n11252), .ZN(P2_U3211) );
  OR2_X1 U13968 ( .A1(n11273), .A2(n11257), .ZN(n11254) );
  OAI21_X1 U13969 ( .B1(n11255), .B2(n11274), .A(n11254), .ZN(n11256) );
  INV_X1 U13970 ( .A(n11257), .ZN(n11258) );
  NAND2_X1 U13971 ( .A1(n11273), .A2(n11258), .ZN(n11265) );
  OAI211_X1 U13972 ( .C1(n13565), .C2(n13514), .A(n11260), .B(n11259), .ZN(
        n11261) );
  INV_X1 U13973 ( .A(n11261), .ZN(n11264) );
  NAND2_X1 U13974 ( .A1(n11274), .A2(n11262), .ZN(n11263) );
  NAND3_X1 U13975 ( .A1(n11265), .A2(n11264), .A3(n11263), .ZN(n11266) );
  NAND2_X1 U13976 ( .A1(n11266), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11269) );
  NAND2_X1 U13977 ( .A1(n11273), .A2(n11267), .ZN(n11268) );
  NOR2_X1 U13978 ( .A1(n13354), .A2(P3_U3151), .ZN(n11788) );
  INV_X1 U13979 ( .A(n11788), .ZN(n11270) );
  NAND2_X1 U13980 ( .A1(n11270), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n11279) );
  OR2_X1 U13981 ( .A1(n11271), .A2(n13529), .ZN(n11272) );
  NOR2_X2 U13982 ( .A1(n11592), .A2(n15916), .ZN(n13349) );
  INV_X1 U13983 ( .A(n15896), .ZN(n15917) );
  NAND2_X1 U13984 ( .A1(n11274), .A2(n15917), .ZN(n11276) );
  AOI22_X1 U13985 ( .A1(n13349), .A2(n11777), .B1(n13357), .B2(n11277), .ZN(
        n11278) );
  OAI211_X1 U13986 ( .C1(n13532), .C2(n13360), .A(n11279), .B(n11278), .ZN(
        P3_U3172) );
  NAND2_X1 U13987 ( .A1(n11281), .A2(n11280), .ZN(n11282) );
  NAND2_X1 U13988 ( .A1(n11283), .A2(n11282), .ZN(n11293) );
  INV_X1 U13989 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11609) );
  OAI21_X1 U13990 ( .B1(n8087), .B2(n11284), .A(n11382), .ZN(n11285) );
  NAND2_X1 U13991 ( .A1(n13748), .A2(n11285), .ZN(n11287) );
  NAND2_X1 U13992 ( .A1(n15894), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n11286) );
  OAI211_X1 U13993 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n11609), .A(n11287), .B(
        n11286), .ZN(n11292) );
  NAND2_X1 U13994 ( .A1(n11288), .A2(n15961), .ZN(n11289) );
  AOI21_X1 U13995 ( .B1(n11290), .B2(n11289), .A(n11321), .ZN(n11291) );
  AOI211_X1 U13996 ( .C1(n13667), .C2(n11293), .A(n11292), .B(n11291), .ZN(
        n11294) );
  OAI21_X1 U13997 ( .B1(n11295), .B2(n13746), .A(n11294), .ZN(P3_U3183) );
  OAI22_X1 U13998 ( .A1(n6546), .A2(n11297), .B1(n11296), .B2(n15712), .ZN(
        n11300) );
  AOI21_X1 U13999 ( .B1(n15367), .B2(n15259), .A(n11298), .ZN(n11299) );
  AOI211_X1 U14000 ( .C1(n6546), .C2(P1_REG2_REG_0__SCAN_IN), .A(n11300), .B(
        n11299), .ZN(n11303) );
  INV_X1 U14001 ( .A(n15374), .ZN(n15688) );
  OAI21_X1 U14002 ( .B1(n15295), .B2(n15688), .A(n12633), .ZN(n11302) );
  NAND2_X1 U14003 ( .A1(n11303), .A2(n11302), .ZN(P1_U3293) );
  INV_X1 U14004 ( .A(n11304), .ZN(n11305) );
  AOI21_X1 U14005 ( .B1(n12154), .B2(n11306), .A(n11305), .ZN(n11322) );
  OAI21_X1 U14006 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n11308), .A(n11307), .ZN(
        n11319) );
  INV_X1 U14007 ( .A(n11309), .ZN(n11314) );
  NOR3_X1 U14008 ( .A1(n11312), .A2(n11311), .A3(n11310), .ZN(n11313) );
  OAI21_X1 U14009 ( .B1(n11314), .B2(n11313), .A(n13748), .ZN(n11316) );
  AND2_X1 U14010 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n11850) );
  AOI21_X1 U14011 ( .B1(n15894), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n11850), .ZN(
        n11315) );
  OAI211_X1 U14012 ( .C1(n13746), .C2(n11317), .A(n11316), .B(n11315), .ZN(
        n11318) );
  AOI21_X1 U14013 ( .B1(n11319), .B2(n13667), .A(n11318), .ZN(n11320) );
  OAI21_X1 U14014 ( .B1(n11322), .B2(n11321), .A(n11320), .ZN(P3_U3191) );
  INV_X1 U14015 ( .A(n11323), .ZN(n11331) );
  INV_X1 U14016 ( .A(n11324), .ZN(n11325) );
  MUX2_X1 U14017 ( .A(n14278), .B(n11325), .S(n15850), .Z(n11330) );
  OAI22_X1 U14018 ( .A1(n14563), .A2(n11326), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n15843), .ZN(n11327) );
  AOI21_X1 U14019 ( .B1(n11328), .B2(n14567), .A(n11327), .ZN(n11329) );
  OAI211_X1 U14020 ( .C1(n11331), .C2(n14546), .A(n11330), .B(n11329), .ZN(
        P2_U3262) );
  INV_X1 U14021 ( .A(n12418), .ZN(n14956) );
  XNOR2_X1 U14022 ( .A(n14956), .B(n12416), .ZN(n12637) );
  INV_X1 U14023 ( .A(n12637), .ZN(n11348) );
  OR2_X1 U14024 ( .A1(n6539), .A2(n12459), .ZN(n11333) );
  INV_X1 U14025 ( .A(n11333), .ZN(n11336) );
  NOR3_X1 U14026 ( .A1(n11332), .A2(n11348), .A3(n11336), .ZN(n11339) );
  AOI22_X1 U14027 ( .A1(n11334), .A2(n11333), .B1(n12459), .B2(n6539), .ZN(
        n11335) );
  OAI211_X2 U14028 ( .C1(n11337), .C2(n11336), .A(n11348), .B(n11335), .ZN(
        n11566) );
  INV_X1 U14029 ( .A(n11566), .ZN(n11338) );
  NOR2_X1 U14030 ( .A1(n11339), .A2(n11338), .ZN(n15771) );
  INV_X1 U14031 ( .A(n11340), .ZN(n11352) );
  NOR2_X1 U14032 ( .A1(n6539), .A2(n11342), .ZN(n11345) );
  NOR3_X1 U14033 ( .A1(n11341), .A2(n11345), .A3(n12637), .ZN(n11350) );
  NAND2_X1 U14034 ( .A1(n6539), .A2(n11342), .ZN(n11343) );
  AND2_X1 U14035 ( .A1(n11344), .A2(n11343), .ZN(n11346) );
  OR2_X1 U14036 ( .A1(n11578), .A2(n11348), .ZN(n15693) );
  INV_X1 U14037 ( .A(n15693), .ZN(n11349) );
  OAI21_X1 U14038 ( .B1(n11350), .B2(n11349), .A(n15763), .ZN(n11351) );
  OAI211_X1 U14039 ( .C1(n15771), .C2(n15745), .A(n11352), .B(n11351), .ZN(
        n15775) );
  NAND2_X1 U14040 ( .A1(n15775), .A2(n15714), .ZN(n11359) );
  AOI211_X1 U14041 ( .C1(n12416), .C2(n11353), .A(n15733), .B(n11586), .ZN(
        n15772) );
  NOR2_X1 U14042 ( .A1(n15367), .A2(n12417), .ZN(n11357) );
  OAI22_X1 U14043 ( .A1(n15714), .A2(n11355), .B1(n11354), .B2(n15712), .ZN(
        n11356) );
  AOI211_X1 U14044 ( .C1(n15772), .C2(n15720), .A(n11357), .B(n11356), .ZN(
        n11358) );
  OAI211_X1 U14045 ( .C1(n15771), .C2(n11360), .A(n11359), .B(n11358), .ZN(
        P1_U3287) );
  OAI21_X1 U14046 ( .B1(n11362), .B2(n12971), .A(n11361), .ZN(n14666) );
  XOR2_X1 U14047 ( .A(n11363), .B(n12971), .Z(n11366) );
  OR2_X1 U14048 ( .A1(n12817), .A2(n14204), .ZN(n11365) );
  NAND2_X1 U14049 ( .A1(n14236), .A2(n14192), .ZN(n11364) );
  NAND2_X1 U14050 ( .A1(n11365), .A2(n11364), .ZN(n12146) );
  AOI21_X1 U14051 ( .B1(n11366), .B2(n14556), .A(n12146), .ZN(n14665) );
  MUX2_X1 U14052 ( .A(n14665), .B(n11367), .S(n14499), .Z(n11372) );
  NAND2_X1 U14053 ( .A1(n11751), .A2(n14663), .ZN(n11368) );
  NAND2_X1 U14054 ( .A1(n11368), .A2(n10836), .ZN(n11369) );
  NOR2_X1 U14055 ( .A1(n6592), .A2(n11369), .ZN(n14662) );
  OAI22_X1 U14056 ( .A1(n7859), .A2(n14563), .B1(n15843), .B2(n12149), .ZN(
        n11370) );
  AOI21_X1 U14057 ( .B1(n14662), .B2(n14567), .A(n11370), .ZN(n11371) );
  OAI211_X1 U14058 ( .C1(n14546), .C2(n14666), .A(n11372), .B(n11371), .ZN(
        P2_U3256) );
  OAI21_X1 U14059 ( .B1(n11375), .B2(n11374), .A(n11373), .ZN(n11389) );
  OAI21_X1 U14060 ( .B1(n11378), .B2(n11377), .A(n11376), .ZN(n11379) );
  NAND2_X1 U14061 ( .A1(n13667), .A2(n11379), .ZN(n11387) );
  NAND2_X1 U14062 ( .A1(n15894), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n11386) );
  NAND2_X1 U14063 ( .A1(P3_U3151), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n11385) );
  AND3_X1 U14064 ( .A1(n11382), .A2(n11381), .A3(n11380), .ZN(n11383) );
  OAI21_X1 U14065 ( .B1(n13600), .B2(n11383), .A(n13748), .ZN(n11384) );
  NAND4_X1 U14066 ( .A1(n11387), .A2(n11386), .A3(n11385), .A4(n11384), .ZN(
        n11388) );
  AOI21_X1 U14067 ( .B1(n13754), .B2(n11389), .A(n11388), .ZN(n11390) );
  OAI21_X1 U14068 ( .B1(n11391), .B2(n13746), .A(n11390), .ZN(P3_U3184) );
  INV_X1 U14069 ( .A(n11400), .ZN(n12968) );
  INV_X1 U14070 ( .A(n11392), .ZN(n11393) );
  OAI21_X1 U14071 ( .B1(n11395), .B2(n11394), .A(n11393), .ZN(n11398) );
  INV_X1 U14072 ( .A(n11396), .ZN(n11397) );
  AOI21_X1 U14073 ( .B1(n12968), .B2(n11398), .A(n11397), .ZN(n11420) );
  INV_X1 U14074 ( .A(n11420), .ZN(n11411) );
  NAND2_X1 U14075 ( .A1(n11100), .A2(n11399), .ZN(n11744) );
  XNOR2_X1 U14076 ( .A(n11744), .B(n11400), .ZN(n11403) );
  NAND2_X1 U14077 ( .A1(n14236), .A2(n14193), .ZN(n11402) );
  NAND2_X1 U14078 ( .A1(n14238), .A2(n14192), .ZN(n11401) );
  AND2_X1 U14079 ( .A1(n11402), .A2(n11401), .ZN(n11674) );
  OAI21_X1 U14080 ( .B1(n11403), .B2(n14534), .A(n11674), .ZN(n11416) );
  INV_X1 U14081 ( .A(n11416), .ZN(n11405) );
  MUX2_X1 U14082 ( .A(n11405), .B(n11404), .S(n14499), .Z(n11410) );
  INV_X1 U14083 ( .A(n11095), .ZN(n11407) );
  INV_X1 U14084 ( .A(n11753), .ZN(n11406) );
  AOI211_X1 U14085 ( .C1(n12807), .C2(n11407), .A(n14635), .B(n11406), .ZN(
        n11415) );
  OAI22_X1 U14086 ( .A1(n14563), .A2(n12808), .B1(n15843), .B2(n11670), .ZN(
        n11408) );
  AOI21_X1 U14087 ( .B1(n11415), .B2(n14567), .A(n11408), .ZN(n11409) );
  OAI211_X1 U14088 ( .C1(n14546), .C2(n11411), .A(n11410), .B(n11409), .ZN(
        P2_U3258) );
  NAND2_X1 U14089 ( .A1(n11412), .A2(n14028), .ZN(n11413) );
  OAI211_X1 U14090 ( .C1(n11414), .C2(n14033), .A(n11413), .B(n13569), .ZN(
        P3_U3272) );
  AOI211_X1 U14091 ( .C1(n12807), .C2(n10017), .A(n11416), .B(n11415), .ZN(
        n11422) );
  AOI22_X1 U14092 ( .A1(n11420), .A2(n11417), .B1(P2_REG1_REG_7__SCAN_IN), 
        .B2(n15890), .ZN(n11418) );
  OAI21_X1 U14093 ( .B1(n11422), .B2(n15890), .A(n11418), .ZN(P2_U3506) );
  AOI22_X1 U14094 ( .A1(n11420), .A2(n11419), .B1(P2_REG0_REG_7__SCAN_IN), 
        .B2(n15885), .ZN(n11421) );
  OAI21_X1 U14095 ( .B1(n11422), .B2(n15885), .A(n11421), .ZN(P2_U3451) );
  XNOR2_X1 U14096 ( .A(n6540), .B(n15756), .ZN(n12635) );
  XNOR2_X1 U14097 ( .A(n11423), .B(n12635), .ZN(n15759) );
  XOR2_X1 U14098 ( .A(n12635), .B(n11424), .Z(n15762) );
  NAND2_X1 U14099 ( .A1(n15762), .A2(n15295), .ZN(n11434) );
  INV_X1 U14100 ( .A(n15717), .ZN(n11426) );
  AOI211_X1 U14101 ( .C1(n15756), .C2(n11426), .A(n15733), .B(n11425), .ZN(
        n15754) );
  INV_X1 U14102 ( .A(n15712), .ZN(n15698) );
  INV_X1 U14103 ( .A(n11427), .ZN(n11429) );
  MUX2_X1 U14104 ( .A(n15755), .B(P1_REG2_REG_4__SCAN_IN), .S(n6546), .Z(
        n11428) );
  AOI21_X1 U14105 ( .B1(n15698), .B2(n11429), .A(n11428), .ZN(n11430) );
  OAI21_X1 U14106 ( .B1(n11431), .B2(n15367), .A(n11430), .ZN(n11432) );
  AOI21_X1 U14107 ( .B1(n15754), .B2(n15720), .A(n11432), .ZN(n11433) );
  OAI211_X1 U14108 ( .C1(n15759), .C2(n15374), .A(n11434), .B(n11433), .ZN(
        P1_U3289) );
  XNOR2_X1 U14109 ( .A(n11482), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n11440) );
  INV_X1 U14110 ( .A(n11435), .ZN(n11436) );
  NOR2_X1 U14111 ( .A1(n11437), .A2(n11436), .ZN(n11467) );
  XNOR2_X1 U14112 ( .A(n11471), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n11466) );
  NOR2_X1 U14113 ( .A1(n11471), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11438) );
  OR2_X1 U14114 ( .A1(n11465), .A2(n11438), .ZN(n11439) );
  AOI211_X1 U14115 ( .C1(n11440), .C2(n11439), .A(n15661), .B(n11477), .ZN(
        n11451) );
  XNOR2_X1 U14116 ( .A(n11482), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n11447) );
  NAND2_X1 U14117 ( .A1(n11441), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n11442) );
  NAND2_X1 U14118 ( .A1(n11443), .A2(n11442), .ZN(n11463) );
  MUX2_X1 U14119 ( .A(n9695), .B(P1_REG2_REG_12__SCAN_IN), .S(n11471), .Z(
        n11464) );
  OR2_X1 U14120 ( .A1(n11471), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11444) );
  NAND2_X1 U14121 ( .A1(n11461), .A2(n11444), .ZN(n11446) );
  INV_X1 U14122 ( .A(n11484), .ZN(n11445) );
  AOI211_X1 U14123 ( .C1(n11447), .C2(n11446), .A(n15111), .B(n11445), .ZN(
        n11450) );
  NAND2_X1 U14124 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n14877)
         );
  NAND2_X1 U14125 ( .A1(n15651), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n11448) );
  OAI211_X1 U14126 ( .C1(n15659), .C2(n11475), .A(n14877), .B(n11448), .ZN(
        n11449) );
  OR3_X1 U14127 ( .A1(n11451), .A2(n11450), .A3(n11449), .ZN(P1_U3256) );
  INV_X1 U14128 ( .A(n11452), .ZN(n11454) );
  OAI222_X1 U14129 ( .A1(n14040), .A2(n11454), .B1(n14033), .B2(n11453), .C1(
        P3_U3151), .C2(n13412), .ZN(P3_U3274) );
  NAND2_X1 U14130 ( .A1(n11458), .A2(n13079), .ZN(n11456) );
  OR2_X1 U14131 ( .A1(n11455), .A2(P2_U3088), .ZN(n12993) );
  OAI211_X1 U14132 ( .C1(n11457), .C2(n13196), .A(n11456), .B(n12993), .ZN(
        P2_U3304) );
  NAND2_X1 U14133 ( .A1(n11458), .A2(n15550), .ZN(n11459) );
  OAI211_X1 U14134 ( .C1(n11460), .C2(n15546), .A(n11459), .B(n12656), .ZN(
        P1_U3332) );
  INV_X1 U14135 ( .A(n11461), .ZN(n11462) );
  AOI21_X1 U14136 ( .B1(n11464), .B2(n11463), .A(n11462), .ZN(n11473) );
  INV_X1 U14137 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n12292) );
  NAND2_X1 U14138 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n14809)
         );
  OAI21_X1 U14139 ( .B1(n15668), .B2(n12292), .A(n14809), .ZN(n11470) );
  AOI21_X1 U14140 ( .B1(n11467), .B2(n11466), .A(n11465), .ZN(n11468) );
  NOR2_X1 U14141 ( .A1(n11468), .A2(n15661), .ZN(n11469) );
  AOI211_X1 U14142 ( .C1(n15085), .C2(n11471), .A(n11470), .B(n11469), .ZN(
        n11472) );
  OAI21_X1 U14143 ( .B1(n11473), .B2(n15111), .A(n11472), .ZN(P1_U3255) );
  XNOR2_X1 U14144 ( .A(n15050), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n11479) );
  NOR2_X1 U14145 ( .A1(n11475), .A2(n11474), .ZN(n11476) );
  OR2_X1 U14146 ( .A1(n11477), .A2(n11476), .ZN(n11478) );
  AOI21_X1 U14147 ( .B1(n11479), .B2(n11478), .A(n15042), .ZN(n11489) );
  NOR2_X1 U14148 ( .A1(n11480), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14755) );
  NOR2_X1 U14149 ( .A1(n15659), .A2(n15044), .ZN(n11481) );
  AOI211_X1 U14150 ( .C1(n15651), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n14755), 
        .B(n11481), .ZN(n11488) );
  NAND2_X1 U14151 ( .A1(n11482), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11483) );
  NAND2_X1 U14152 ( .A1(n11484), .A2(n11483), .ZN(n11486) );
  XNOR2_X1 U14153 ( .A(n15050), .B(n15349), .ZN(n11485) );
  NAND2_X1 U14154 ( .A1(n11486), .A2(n11485), .ZN(n15052) );
  OAI211_X1 U14155 ( .C1(n11486), .C2(n11485), .A(n15052), .B(n15665), .ZN(
        n11487) );
  OAI211_X1 U14156 ( .C1(n11489), .C2(n15661), .A(n11488), .B(n11487), .ZN(
        P1_U3257) );
  XNOR2_X1 U14157 ( .A(n6595), .B(n13432), .ZN(n15942) );
  INV_X1 U14158 ( .A(n15942), .ZN(n11498) );
  INV_X1 U14159 ( .A(n11490), .ZN(n15897) );
  NOR2_X1 U14160 ( .A1(n15903), .A2(n15897), .ZN(n12748) );
  INV_X1 U14161 ( .A(n13432), .ZN(n13533) );
  NOR2_X1 U14162 ( .A1(n11491), .A2(n13533), .ZN(n11514) );
  AOI21_X1 U14163 ( .B1(n13533), .B2(n11491), .A(n11514), .ZN(n11493) );
  AOI22_X1 U14164 ( .A1(n13886), .A2(n13587), .B1(n13889), .B2(n13589), .ZN(
        n11492) );
  OAI21_X1 U14165 ( .B1(n11493), .B2(n15911), .A(n11492), .ZN(n11494) );
  AOI21_X1 U14166 ( .B1(n15942), .B2(n12708), .A(n11494), .ZN(n15939) );
  MUX2_X1 U14167 ( .A(n11632), .B(n15939), .S(n15921), .Z(n11497) );
  NOR2_X1 U14168 ( .A1(n15948), .A2(n11495), .ZN(n15941) );
  AOI22_X1 U14169 ( .A1(n11764), .A2(n15941), .B1(n15901), .B2(n11854), .ZN(
        n11496) );
  OAI211_X1 U14170 ( .C1(n11498), .C2(n11932), .A(n11497), .B(n11496), .ZN(
        P3_U3228) );
  AOI21_X1 U14171 ( .B1(n11500), .B2(n11501), .A(n11499), .ZN(n15934) );
  INV_X1 U14172 ( .A(n11501), .ZN(n13534) );
  XNOR2_X1 U14173 ( .A(n11502), .B(n13534), .ZN(n11505) );
  INV_X1 U14174 ( .A(n12708), .ZN(n13964) );
  AOI22_X1 U14175 ( .A1(n13886), .A2(n13588), .B1(n13889), .B2(n13590), .ZN(
        n11503) );
  OAI21_X1 U14176 ( .B1(n15934), .B2(n13964), .A(n11503), .ZN(n11504) );
  AOI21_X1 U14177 ( .B1(n11505), .B2(n13960), .A(n11504), .ZN(n15935) );
  MUX2_X1 U14178 ( .A(n11506), .B(n15935), .S(n15921), .Z(n11508) );
  NOR2_X1 U14179 ( .A1(n15948), .A2(n12081), .ZN(n15937) );
  AOI22_X1 U14180 ( .A1(n11764), .A2(n15937), .B1(n15901), .B2(n12083), .ZN(
        n11507) );
  OAI211_X1 U14181 ( .C1(n15934), .C2(n11932), .A(n11508), .B(n11507), .ZN(
        P3_U3229) );
  XNOR2_X1 U14182 ( .A(n11510), .B(n11509), .ZN(n15945) );
  INV_X1 U14183 ( .A(n15945), .ZN(n11522) );
  OAI22_X1 U14184 ( .A1(n11840), .A2(n15916), .B1(n15914), .B2(n11820), .ZN(
        n11518) );
  INV_X1 U14185 ( .A(n11514), .ZN(n11512) );
  AOI21_X1 U14186 ( .B1(n11512), .B2(n11511), .A(n13536), .ZN(n11516) );
  OR2_X1 U14187 ( .A1(n11514), .A2(n11513), .ZN(n11878) );
  INV_X1 U14188 ( .A(n11878), .ZN(n11515) );
  NOR3_X1 U14189 ( .A1(n11516), .A2(n11515), .A3(n15911), .ZN(n11517) );
  AOI211_X1 U14190 ( .C1(n15945), .C2(n12708), .A(n11518), .B(n11517), .ZN(
        n15947) );
  MUX2_X1 U14191 ( .A(n11519), .B(n15947), .S(n15921), .Z(n11521) );
  AOI22_X1 U14192 ( .A1(n13880), .A2(n15943), .B1(n15901), .B2(n11804), .ZN(
        n11520) );
  OAI211_X1 U14193 ( .C1(n11522), .C2(n11932), .A(n11521), .B(n11520), .ZN(
        P3_U3227) );
  XNOR2_X1 U14194 ( .A(n11523), .B(n11524), .ZN(n15933) );
  INV_X1 U14195 ( .A(n15933), .ZN(n11534) );
  OAI22_X1 U14196 ( .A1(n15915), .A2(n15914), .B1(n15916), .B2(n11855), .ZN(
        n11528) );
  AOI21_X1 U14197 ( .B1(n13957), .B2(n11525), .A(n13531), .ZN(n11526) );
  NOR3_X1 U14198 ( .A1(n6750), .A2(n11526), .A3(n15911), .ZN(n11527) );
  AOI211_X1 U14199 ( .C1(n15933), .C2(n12708), .A(n11528), .B(n11527), .ZN(
        n15930) );
  MUX2_X1 U14200 ( .A(n11529), .B(n15930), .S(n15921), .Z(n11533) );
  NOR2_X1 U14201 ( .A1(n15948), .A2(n11530), .ZN(n15932) );
  AOI22_X1 U14202 ( .A1(n11764), .A2(n15932), .B1(n15901), .B2(n11531), .ZN(
        n11532) );
  OAI211_X1 U14203 ( .C1(n11534), .C2(n11932), .A(n11533), .B(n11532), .ZN(
        P3_U3230) );
  INV_X1 U14204 ( .A(n11535), .ZN(n11539) );
  NAND2_X1 U14205 ( .A1(n11539), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11536) );
  NAND2_X1 U14206 ( .A1(n11537), .A2(n11536), .ZN(n11654) );
  XNOR2_X1 U14207 ( .A(n11652), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n11545) );
  NAND2_X1 U14208 ( .A1(P2_U3088), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n14049)
         );
  AOI21_X1 U14209 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n11539), .A(n11538), 
        .ZN(n11658) );
  XNOR2_X1 U14210 ( .A(n11653), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n11657) );
  XOR2_X1 U14211 ( .A(n11658), .B(n11657), .Z(n11540) );
  NAND2_X1 U14212 ( .A1(n15815), .A2(n11540), .ZN(n11541) );
  NAND2_X1 U14213 ( .A1(n14049), .A2(n11541), .ZN(n11543) );
  NOR2_X1 U14214 ( .A1(n15806), .A2(n11656), .ZN(n11542) );
  AOI211_X1 U14215 ( .C1(n15809), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n11543), 
        .B(n11542), .ZN(n11544) );
  OAI21_X1 U14216 ( .B1(n11545), .B2(n15832), .A(n11544), .ZN(P2_U3228) );
  OR2_X1 U14217 ( .A1(n11546), .A2(n12964), .ZN(n11547) );
  NAND2_X1 U14218 ( .A1(n11548), .A2(n11547), .ZN(n15876) );
  INV_X1 U14219 ( .A(n15876), .ZN(n11563) );
  INV_X1 U14220 ( .A(n12764), .ZN(n15849) );
  NAND2_X1 U14221 ( .A1(n15850), .A2(n15849), .ZN(n14564) );
  NAND2_X1 U14222 ( .A1(n11551), .A2(n11550), .ZN(n11549) );
  NAND2_X1 U14223 ( .A1(n11549), .A2(n6958), .ZN(n11795) );
  NAND3_X1 U14224 ( .A1(n11551), .A2(n12964), .A3(n11550), .ZN(n11552) );
  AND2_X1 U14225 ( .A1(n11795), .A2(n11552), .ZN(n11555) );
  NAND2_X1 U14226 ( .A1(n15876), .A2(n12163), .ZN(n11554) );
  OAI211_X1 U14227 ( .C1(n11555), .C2(n14534), .A(n11554), .B(n11553), .ZN(
        n15875) );
  MUX2_X1 U14228 ( .A(n15875), .B(P2_REG2_REG_4__SCAN_IN), .S(n14499), .Z(
        n11556) );
  INV_X1 U14229 ( .A(n11556), .ZN(n11562) );
  INV_X1 U14230 ( .A(n11557), .ZN(n11792) );
  AOI211_X1 U14231 ( .C1(n12795), .C2(n11558), .A(n14635), .B(n11792), .ZN(
        n15871) );
  OAI22_X1 U14232 ( .A1(n14563), .A2(n15873), .B1(n15843), .B2(n11559), .ZN(
        n11560) );
  AOI21_X1 U14233 ( .B1(n15871), .B2(n14567), .A(n11560), .ZN(n11561) );
  OAI211_X1 U14234 ( .C1(n11563), .C2(n14564), .A(n11562), .B(n11561), .ZN(
        P2_U3261) );
  INV_X1 U14235 ( .A(n11564), .ZN(n15198) );
  NAND2_X1 U14236 ( .A1(n12418), .A2(n12417), .ZN(n11565) );
  NAND2_X1 U14237 ( .A1(n11566), .A2(n11565), .ZN(n15691) );
  XNOR2_X1 U14238 ( .A(n15702), .B(n12415), .ZN(n15694) );
  NAND2_X1 U14239 ( .A1(n12414), .A2(n12415), .ZN(n11567) );
  NAND2_X1 U14240 ( .A1(n15676), .A2(n15675), .ZN(n15674) );
  OR2_X1 U14241 ( .A1(n15684), .A2(n14954), .ZN(n11568) );
  NAND2_X1 U14242 ( .A1(n15674), .A2(n11568), .ZN(n11570) );
  INV_X1 U14243 ( .A(n14953), .ZN(n11937) );
  XNOR2_X1 U14244 ( .A(n12475), .B(n11937), .ZN(n12639) );
  AND2_X1 U14245 ( .A1(n15675), .A2(n12639), .ZN(n11569) );
  OAI21_X1 U14246 ( .B1(n11570), .B2(n12639), .A(n11948), .ZN(n11571) );
  INV_X1 U14247 ( .A(n11571), .ZN(n15516) );
  INV_X1 U14248 ( .A(n12415), .ZN(n14955) );
  NAND2_X1 U14249 ( .A1(n12414), .A2(n14955), .ZN(n11572) );
  INV_X1 U14250 ( .A(n11572), .ZN(n11575) );
  NAND2_X1 U14251 ( .A1(n12416), .A2(n12418), .ZN(n15692) );
  AND2_X1 U14252 ( .A1(n15692), .A2(n11573), .ZN(n11574) );
  OR2_X1 U14253 ( .A1(n11575), .A2(n11574), .ZN(n11576) );
  INV_X1 U14254 ( .A(n14954), .ZN(n11579) );
  NAND2_X1 U14255 ( .A1(n11581), .A2(n12639), .ZN(n11582) );
  AOI21_X1 U14256 ( .B1(n11939), .B2(n11582), .A(n15709), .ZN(n15514) );
  NAND2_X1 U14257 ( .A1(n14952), .A2(n15636), .ZN(n11584) );
  NAND2_X1 U14258 ( .A1(n14954), .A2(n15637), .ZN(n11583) );
  NAND2_X1 U14259 ( .A1(n11584), .A2(n11583), .ZN(n15511) );
  NOR2_X1 U14260 ( .A1(n15514), .A2(n15511), .ZN(n11585) );
  MUX2_X1 U14261 ( .A(n10774), .B(n11585), .S(n15714), .Z(n11591) );
  INV_X1 U14262 ( .A(n11587), .ZN(n15679) );
  INV_X1 U14263 ( .A(n12475), .ZN(n14853) );
  NAND2_X1 U14264 ( .A1(n11587), .A2(n14853), .ZN(n12212) );
  INV_X1 U14265 ( .A(n12212), .ZN(n11588) );
  AOI211_X1 U14266 ( .C1(n12475), .C2(n15679), .A(n15733), .B(n11588), .ZN(
        n15512) );
  OAI22_X1 U14267 ( .A1(n15367), .A2(n14853), .B1(n14856), .B2(n15712), .ZN(
        n11589) );
  AOI21_X1 U14268 ( .B1(n15512), .B2(n15720), .A(n11589), .ZN(n11590) );
  OAI211_X1 U14269 ( .C1(n15198), .C2(n15516), .A(n11591), .B(n11590), .ZN(
        P1_U3284) );
  INV_X1 U14270 ( .A(n11592), .ZN(n11593) );
  INV_X1 U14271 ( .A(n13352), .ZN(n13263) );
  INV_X1 U14272 ( .A(n11595), .ZN(n13561) );
  OAI21_X1 U14273 ( .B1(n13412), .B2(n11596), .A(n13529), .ZN(n11597) );
  NAND2_X4 U14274 ( .A1(n11599), .A2(n11598), .ZN(n12695) );
  INV_X1 U14275 ( .A(n11604), .ZN(n15910) );
  OAI21_X1 U14276 ( .B1(n12695), .B2(n15910), .A(n11600), .ZN(n11601) );
  INV_X1 U14277 ( .A(n15904), .ZN(n11602) );
  NAND3_X1 U14278 ( .A1(n12695), .A2(n11594), .A3(n11602), .ZN(n11603) );
  OAI211_X1 U14279 ( .C1(n11605), .C2(n11604), .A(n11781), .B(n11603), .ZN(
        n11606) );
  AOI22_X1 U14280 ( .A1(n13263), .A2(n15906), .B1(n13325), .B2(n11606), .ZN(
        n11608) );
  AOI22_X1 U14281 ( .A1(n13349), .A2(n13591), .B1(n13357), .B2(n11778), .ZN(
        n11607) );
  OAI211_X1 U14282 ( .C1(n11788), .C2(n11609), .A(n11608), .B(n11607), .ZN(
        P3_U3162) );
  AND3_X1 U14283 ( .A1(n11635), .A2(n11611), .A3(n11610), .ZN(n11612) );
  OAI21_X1 U14284 ( .B1(n11613), .B2(n11612), .A(n13667), .ZN(n11622) );
  INV_X1 U14285 ( .A(n11614), .ZN(n11616) );
  NAND3_X1 U14286 ( .A1(n11638), .A2(n11616), .A3(n11615), .ZN(n11617) );
  NAND2_X1 U14287 ( .A1(n11618), .A2(n11617), .ZN(n11619) );
  NAND2_X1 U14288 ( .A1(n13754), .A2(n11619), .ZN(n11621) );
  AND2_X1 U14289 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n11822) );
  AOI21_X1 U14290 ( .B1(n15894), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n11822), .ZN(
        n11620) );
  NAND3_X1 U14291 ( .A1(n11622), .A2(n11621), .A3(n11620), .ZN(n11629) );
  INV_X1 U14292 ( .A(n11623), .ZN(n11627) );
  NAND3_X1 U14293 ( .A1(n11647), .A2(n11625), .A3(n11624), .ZN(n11626) );
  AOI21_X1 U14294 ( .B1(n11627), .B2(n11626), .A(n13720), .ZN(n11628) );
  AOI211_X1 U14295 ( .C1(n13722), .C2(n11630), .A(n11629), .B(n11628), .ZN(
        n11631) );
  INV_X1 U14296 ( .A(n11631), .ZN(P3_U3188) );
  NAND2_X1 U14297 ( .A1(n11633), .A2(n11632), .ZN(n11634) );
  AND2_X1 U14298 ( .A1(n11635), .A2(n11634), .ZN(n11642) );
  NAND2_X1 U14299 ( .A1(n11636), .A2(n15967), .ZN(n11637) );
  NAND2_X1 U14300 ( .A1(n11638), .A2(n11637), .ZN(n11639) );
  NAND2_X1 U14301 ( .A1(n13754), .A2(n11639), .ZN(n11641) );
  AND2_X1 U14302 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n11857) );
  AOI21_X1 U14303 ( .B1(n15894), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n11857), .ZN(
        n11640) );
  OAI211_X1 U14304 ( .C1(n11642), .C2(n13757), .A(n11641), .B(n11640), .ZN(
        n11649) );
  NAND3_X1 U14305 ( .A1(n6822), .A2(n11645), .A3(n11644), .ZN(n11646) );
  AOI21_X1 U14306 ( .B1(n11647), .B2(n11646), .A(n13720), .ZN(n11648) );
  AOI211_X1 U14307 ( .C1(n13722), .C2(n11650), .A(n11649), .B(n11648), .ZN(
        n11651) );
  INV_X1 U14308 ( .A(n11651), .ZN(P3_U3187) );
  NAND2_X1 U14309 ( .A1(n11654), .A2(n11653), .ZN(n11655) );
  XNOR2_X1 U14310 ( .A(n11978), .B(P2_REG2_REG_15__SCAN_IN), .ZN(n11665) );
  OAI22_X1 U14311 ( .A1(n11658), .A2(n11657), .B1(n11656), .B2(n14644), .ZN(
        n11974) );
  INV_X1 U14312 ( .A(n11974), .ZN(n11659) );
  XNOR2_X1 U14313 ( .A(n11659), .B(n11979), .ZN(n11973) );
  XNOR2_X1 U14314 ( .A(n11973), .B(n14639), .ZN(n11663) );
  NAND2_X1 U14315 ( .A1(n15809), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n11660) );
  NAND2_X1 U14316 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n14208)
         );
  OAI211_X1 U14317 ( .C1(n15806), .C2(n11661), .A(n11660), .B(n14208), .ZN(
        n11662) );
  AOI21_X1 U14318 ( .B1(n11663), .B2(n15815), .A(n11662), .ZN(n11664) );
  OAI21_X1 U14319 ( .B1(n11665), .B2(n15832), .A(n11664), .ZN(P2_U3229) );
  XNOR2_X1 U14320 ( .A(n12807), .B(n7818), .ZN(n11896) );
  NOR2_X1 U14321 ( .A1(n12809), .A2(n13148), .ZN(n11897) );
  XNOR2_X1 U14322 ( .A(n11896), .B(n11897), .ZN(n11900) );
  XNOR2_X1 U14323 ( .A(n11901), .B(n11900), .ZN(n11677) );
  INV_X1 U14324 ( .A(n11670), .ZN(n11671) );
  NAND2_X1 U14325 ( .A1(n14194), .A2(n11671), .ZN(n11673) );
  OAI211_X1 U14326 ( .C1(n11674), .C2(n14196), .A(n11673), .B(n11672), .ZN(
        n11675) );
  AOI21_X1 U14327 ( .B1(n12807), .B2(n14211), .A(n11675), .ZN(n11676) );
  OAI21_X1 U14328 ( .B1(n11677), .B2(n14213), .A(n11676), .ZN(P2_U3185) );
  INV_X1 U14329 ( .A(n11678), .ZN(n11680) );
  NAND3_X1 U14330 ( .A1(n13595), .A2(n11680), .A3(n11679), .ZN(n11681) );
  NAND2_X1 U14331 ( .A1(n11682), .A2(n11681), .ZN(n11695) );
  INV_X1 U14332 ( .A(n11683), .ZN(n11685) );
  NAND3_X1 U14333 ( .A1(n13594), .A2(n11685), .A3(n11684), .ZN(n11686) );
  AND2_X1 U14334 ( .A1(n11687), .A2(n11686), .ZN(n11689) );
  NAND2_X1 U14335 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n12079) );
  NAND2_X1 U14336 ( .A1(n15894), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n11688) );
  OAI211_X1 U14337 ( .C1(n13757), .C2(n11689), .A(n12079), .B(n11688), .ZN(
        n11694) );
  NAND3_X1 U14338 ( .A1(n13598), .A2(n11691), .A3(n11690), .ZN(n11692) );
  AOI21_X1 U14339 ( .B1(n6822), .B2(n11692), .A(n13720), .ZN(n11693) );
  AOI211_X1 U14340 ( .C1(n13754), .C2(n11695), .A(n11694), .B(n11693), .ZN(
        n11696) );
  OAI21_X1 U14341 ( .B1(n11697), .B2(n13746), .A(n11696), .ZN(P3_U3186) );
  OAI21_X1 U14342 ( .B1(n11700), .B2(n11699), .A(n11698), .ZN(n15870) );
  INV_X1 U14343 ( .A(n15870), .ZN(n11713) );
  OAI21_X1 U14344 ( .B1(n11702), .B2(n12960), .A(n11701), .ZN(n11704) );
  AOI21_X1 U14345 ( .B1(n11704), .B2(n14556), .A(n11703), .ZN(n11705) );
  OAI21_X1 U14346 ( .B1(n11713), .B2(n14552), .A(n11705), .ZN(n15868) );
  NAND2_X1 U14347 ( .A1(n15868), .A2(n15850), .ZN(n11712) );
  OAI22_X1 U14348 ( .A1(n15850), .A2(n10645), .B1(n14261), .B2(n15843), .ZN(
        n11710) );
  INV_X1 U14349 ( .A(n11706), .ZN(n11708) );
  OAI211_X1 U14350 ( .C1(n15867), .C2(n11708), .A(n11707), .B(n10836), .ZN(
        n15866) );
  NOR2_X1 U14351 ( .A1(n14330), .A2(n15866), .ZN(n11709) );
  AOI211_X1 U14352 ( .C1(n14541), .C2(n12784), .A(n11710), .B(n11709), .ZN(
        n11711) );
  OAI211_X1 U14353 ( .C1(n11713), .C2(n14564), .A(n11712), .B(n11711), .ZN(
        P2_U3263) );
  NAND2_X1 U14354 ( .A1(n11717), .A2(n11716), .ZN(n11719) );
  NAND2_X1 U14355 ( .A1(n11719), .A2(n11718), .ZN(n11727) );
  INV_X1 U14356 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n11720) );
  XNOR2_X1 U14357 ( .A(n11720), .B(P1_ADDR_REG_9__SCAN_IN), .ZN(n11726) );
  XNOR2_X1 U14358 ( .A(n11727), .B(n11726), .ZN(n11722) );
  XNOR2_X1 U14359 ( .A(n11721), .B(n11722), .ZN(n15558) );
  INV_X1 U14360 ( .A(n11721), .ZN(n11723) );
  NAND2_X1 U14361 ( .A1(n11723), .A2(n11722), .ZN(n11724) );
  INV_X1 U14362 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n11728) );
  NAND2_X1 U14363 ( .A1(n11728), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n11729) );
  NAND2_X1 U14364 ( .A1(n11731), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n12127) );
  INV_X1 U14365 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n11732) );
  NAND2_X1 U14366 ( .A1(n11732), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n11733) );
  NAND2_X1 U14367 ( .A1(n12127), .A2(n11733), .ZN(n12128) );
  INV_X1 U14368 ( .A(n12128), .ZN(n11734) );
  XNOR2_X1 U14369 ( .A(n12129), .B(n11734), .ZN(n11735) );
  NAND2_X1 U14370 ( .A1(n12126), .A2(n12125), .ZN(n11736) );
  XNOR2_X1 U14371 ( .A(n11736), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  OR2_X1 U14372 ( .A1(n11738), .A2(n11737), .ZN(n11739) );
  NAND2_X1 U14373 ( .A1(n11740), .A2(n11739), .ZN(n14672) );
  OR2_X1 U14374 ( .A1(n12820), .A2(n14204), .ZN(n11742) );
  OR2_X1 U14375 ( .A1(n12809), .A2(n14202), .ZN(n11741) );
  AND2_X1 U14376 ( .A1(n11742), .A2(n11741), .ZN(n11914) );
  NAND2_X1 U14377 ( .A1(n11744), .A2(n11743), .ZN(n11746) );
  NAND2_X1 U14378 ( .A1(n11746), .A2(n11745), .ZN(n11747) );
  XNOR2_X1 U14379 ( .A(n11747), .B(n12969), .ZN(n11748) );
  NAND2_X1 U14380 ( .A1(n11748), .A2(n14556), .ZN(n11749) );
  OAI211_X1 U14381 ( .C1(n14672), .C2(n14552), .A(n11914), .B(n11749), .ZN(
        n14669) );
  MUX2_X1 U14382 ( .A(n14669), .B(P2_REG2_REG_8__SCAN_IN), .S(n14499), .Z(
        n11750) );
  INV_X1 U14383 ( .A(n11750), .ZN(n11756) );
  INV_X1 U14384 ( .A(n11751), .ZN(n11752) );
  AOI211_X1 U14385 ( .C1(n14668), .C2(n11753), .A(n14635), .B(n11752), .ZN(
        n14667) );
  OAI22_X1 U14386 ( .A1(n14563), .A2(n7924), .B1(n15843), .B2(n11910), .ZN(
        n11754) );
  AOI21_X1 U14387 ( .B1(n14667), .B2(n14567), .A(n11754), .ZN(n11755) );
  OAI211_X1 U14388 ( .C1(n14672), .C2(n14564), .A(n11756), .B(n11755), .ZN(
        P2_U3257) );
  XNOR2_X1 U14389 ( .A(n11758), .B(n11757), .ZN(n15958) );
  INV_X1 U14390 ( .A(n15958), .ZN(n11767) );
  NOR2_X1 U14391 ( .A1(n11759), .A2(n13538), .ZN(n11919) );
  AOI21_X1 U14392 ( .B1(n13538), .B2(n11759), .A(n11919), .ZN(n11760) );
  NOR2_X1 U14393 ( .A1(n11760), .A2(n15911), .ZN(n11762) );
  OAI22_X1 U14394 ( .A1(n12034), .A2(n15916), .B1(n15914), .B2(n11840), .ZN(
        n11761) );
  AOI211_X1 U14395 ( .C1(n15958), .C2(n12708), .A(n11762), .B(n11761), .ZN(
        n15954) );
  MUX2_X1 U14396 ( .A(n11763), .B(n15954), .S(n15921), .Z(n11766) );
  NOR2_X1 U14397 ( .A1(n12178), .A2(n15948), .ZN(n15956) );
  AOI22_X1 U14398 ( .A1(n11764), .A2(n15956), .B1(n15901), .B2(n12180), .ZN(
        n11765) );
  OAI211_X1 U14399 ( .C1(n11767), .C2(n11932), .A(n11766), .B(n11765), .ZN(
        P3_U3225) );
  INV_X1 U14400 ( .A(n11768), .ZN(n11771) );
  INV_X1 U14401 ( .A(n11769), .ZN(n11773) );
  OAI222_X1 U14402 ( .A1(n11771), .A2(P2_U3088), .B1(n13198), .B2(n11773), 
        .C1(n11770), .C2(n13196), .ZN(P2_U3303) );
  OAI222_X1 U14403 ( .A1(P1_U3086), .A2(n11774), .B1(n10985), .B2(n11773), 
        .C1(n11772), .C2(n15546), .ZN(P1_U3331) );
  INV_X1 U14404 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n11787) );
  OAI22_X1 U14405 ( .A1(n13319), .A2(n13955), .B1(n13965), .B2(n13333), .ZN(
        n11776) );
  AOI21_X1 U14406 ( .B1(n13263), .B2(n11777), .A(n11776), .ZN(n11786) );
  XNOR2_X1 U14407 ( .A(n12695), .B(n8154), .ZN(n11805) );
  XNOR2_X1 U14408 ( .A(n11805), .B(n13591), .ZN(n11783) );
  XNOR2_X1 U14409 ( .A(n12695), .B(n11778), .ZN(n11779) );
  NAND2_X1 U14410 ( .A1(n11779), .A2(n13954), .ZN(n11780) );
  OAI21_X1 U14411 ( .B1(n11783), .B2(n11782), .A(n11807), .ZN(n11784) );
  NAND2_X1 U14412 ( .A1(n11784), .A2(n13325), .ZN(n11785) );
  OAI211_X1 U14413 ( .C1(n11788), .C2(n11787), .A(n11786), .B(n11785), .ZN(
        P3_U3177) );
  INV_X1 U14414 ( .A(n14546), .ZN(n14461) );
  XNOR2_X1 U14415 ( .A(n12963), .B(n11789), .ZN(n15883) );
  INV_X1 U14416 ( .A(n11790), .ZN(n11791) );
  OAI211_X1 U14417 ( .C1(n15880), .C2(n11792), .A(n11791), .B(n10836), .ZN(
        n15878) );
  INV_X1 U14418 ( .A(n15843), .ZN(n14560) );
  AOI22_X1 U14419 ( .A1(n14541), .A2(n12799), .B1(n14560), .B2(n11793), .ZN(
        n11794) );
  OAI21_X1 U14420 ( .B1(n15878), .B2(n14330), .A(n11794), .ZN(n11802) );
  AND3_X1 U14421 ( .A1(n12963), .A2(n11796), .A3(n11795), .ZN(n11798) );
  OAI21_X1 U14422 ( .B1(n11798), .B2(n11797), .A(n14556), .ZN(n11800) );
  NAND2_X1 U14423 ( .A1(n11800), .A2(n11799), .ZN(n15881) );
  MUX2_X1 U14424 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n15881), .S(n15850), .Z(
        n11801) );
  AOI211_X1 U14425 ( .C1(n14461), .C2(n15883), .A(n11802), .B(n11801), .ZN(
        n11803) );
  INV_X1 U14426 ( .A(n11803), .ZN(P2_U3260) );
  INV_X1 U14427 ( .A(n11804), .ZN(n11825) );
  INV_X1 U14428 ( .A(n13354), .ZN(n13242) );
  XNOR2_X1 U14429 ( .A(n11808), .B(n13590), .ZN(n13240) );
  NAND2_X1 U14430 ( .A1(n11805), .A2(n15915), .ZN(n13238) );
  INV_X1 U14431 ( .A(n11808), .ZN(n11809) );
  NAND2_X1 U14432 ( .A1(n11809), .A2(n13590), .ZN(n11810) );
  XNOR2_X1 U14433 ( .A(n12695), .B(n11811), .ZN(n11812) );
  NAND2_X1 U14434 ( .A1(n11812), .A2(n11855), .ZN(n11815) );
  INV_X1 U14435 ( .A(n11812), .ZN(n11813) );
  NAND2_X1 U14436 ( .A1(n11813), .A2(n13589), .ZN(n11814) );
  XNOR2_X1 U14437 ( .A(n12695), .B(n11858), .ZN(n11816) );
  XNOR2_X1 U14438 ( .A(n11816), .B(n13588), .ZN(n11860) );
  NAND2_X1 U14439 ( .A1(n11816), .A2(n11820), .ZN(n11833) );
  AND2_X1 U14440 ( .A1(n11837), .A2(n11833), .ZN(n11819) );
  XNOR2_X1 U14441 ( .A(n12695), .B(n11817), .ZN(n11834) );
  XNOR2_X1 U14442 ( .A(n11834), .B(n11880), .ZN(n11818) );
  NAND2_X1 U14443 ( .A1(n11819), .A2(n11818), .ZN(n11826) );
  OAI211_X1 U14444 ( .C1(n11819), .C2(n11818), .A(n11826), .B(n13325), .ZN(
        n11824) );
  OAI22_X1 U14445 ( .A1(n13319), .A2(n11840), .B1(n11820), .B2(n13352), .ZN(
        n11821) );
  AOI211_X1 U14446 ( .C1(n13357), .C2(n15943), .A(n11822), .B(n11821), .ZN(
        n11823) );
  OAI211_X1 U14447 ( .C1(n11825), .C2(n13242), .A(n11824), .B(n11823), .ZN(
        P3_U3179) );
  NAND2_X1 U14448 ( .A1(n11834), .A2(n13587), .ZN(n11838) );
  NAND2_X1 U14449 ( .A1(n11826), .A2(n11838), .ZN(n12173) );
  XNOR2_X1 U14450 ( .A(n11839), .B(n12173), .ZN(n11832) );
  OAI22_X1 U14451 ( .A1(n13319), .A2(n11925), .B1(n11880), .B2(n13352), .ZN(
        n11827) );
  AOI211_X1 U14452 ( .C1(n13357), .C2(n11829), .A(n11828), .B(n11827), .ZN(
        n11831) );
  NAND2_X1 U14453 ( .A1(n13354), .A2(n11885), .ZN(n11830) );
  OAI211_X1 U14454 ( .C1(n11832), .C2(n13360), .A(n11831), .B(n11830), .ZN(
        P3_U3153) );
  XNOR2_X1 U14455 ( .A(n12695), .B(n12156), .ZN(n12033) );
  XNOR2_X1 U14456 ( .A(n12033), .B(n13584), .ZN(n11848) );
  OAI211_X1 U14457 ( .C1(n11834), .C2(n13587), .A(n11833), .B(n11839), .ZN(
        n11835) );
  NOR2_X1 U14458 ( .A1(n12175), .A2(n11835), .ZN(n11836) );
  OAI21_X1 U14459 ( .B1(n12175), .B2(n11838), .A(n11839), .ZN(n11843) );
  OAI21_X1 U14460 ( .B1(n12175), .B2(n11840), .A(n12172), .ZN(n11842) );
  INV_X1 U14461 ( .A(n12037), .ZN(n11846) );
  AOI21_X1 U14462 ( .B1(n11848), .B2(n11847), .A(n11846), .ZN(n11853) );
  INV_X1 U14463 ( .A(n12156), .ZN(n11993) );
  OAI22_X1 U14464 ( .A1(n13319), .A2(n12304), .B1(n11925), .B2(n13352), .ZN(
        n11849) );
  AOI211_X1 U14465 ( .C1(n13357), .C2(n11993), .A(n11850), .B(n11849), .ZN(
        n11852) );
  NAND2_X1 U14466 ( .A1(n13354), .A2(n11929), .ZN(n11851) );
  OAI211_X1 U14467 ( .C1(n11853), .C2(n13360), .A(n11852), .B(n11851), .ZN(
        P3_U3171) );
  INV_X1 U14468 ( .A(n11854), .ZN(n11864) );
  OAI22_X1 U14469 ( .A1(n13319), .A2(n11880), .B1(n11855), .B2(n13352), .ZN(
        n11856) );
  AOI211_X1 U14470 ( .C1(n13357), .C2(n11858), .A(n11857), .B(n11856), .ZN(
        n11863) );
  OAI21_X1 U14471 ( .B1(n11860), .B2(n11859), .A(n11837), .ZN(n11861) );
  NAND2_X1 U14472 ( .A1(n11861), .A2(n13325), .ZN(n11862) );
  OAI211_X1 U14473 ( .C1(n11864), .C2(n13242), .A(n11863), .B(n11862), .ZN(
        P3_U3167) );
  NAND2_X1 U14474 ( .A1(n11866), .A2(n11865), .ZN(n11867) );
  AOI21_X1 U14475 ( .B1(n11868), .B2(n11867), .A(n15634), .ZN(n11874) );
  NAND2_X1 U14476 ( .A1(n15684), .A2(n15757), .ZN(n15787) );
  OR2_X1 U14477 ( .A1(n15787), .A2(n14901), .ZN(n11872) );
  OR2_X1 U14478 ( .A1(n12415), .A2(n14922), .ZN(n11870) );
  NAND2_X1 U14479 ( .A1(n14953), .A2(n15636), .ZN(n11869) );
  NAND2_X1 U14480 ( .A1(n11870), .A2(n11869), .ZN(n15672) );
  AOI22_X1 U14481 ( .A1(n15641), .A2(n15672), .B1(P1_REG3_REG_8__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11871) );
  OAI211_X1 U14482 ( .C1(n15646), .C2(n15681), .A(n11872), .B(n11871), .ZN(
        n11873) );
  OR2_X1 U14483 ( .A1(n11874), .A2(n11873), .ZN(P1_U3221) );
  AOI21_X1 U14484 ( .B1(n11876), .B2(n13437), .A(n11875), .ZN(n15951) );
  NOR2_X1 U14485 ( .A1(n15951), .A2(n15897), .ZN(n11884) );
  NAND2_X1 U14486 ( .A1(n11878), .A2(n11877), .ZN(n11879) );
  XNOR2_X1 U14487 ( .A(n11879), .B(n13539), .ZN(n11882) );
  OAI22_X1 U14488 ( .A1(n11925), .A2(n15916), .B1(n15914), .B2(n11880), .ZN(
        n11881) );
  AOI21_X1 U14489 ( .B1(n11882), .B2(n13960), .A(n11881), .ZN(n11883) );
  OAI21_X1 U14490 ( .B1(n15951), .B2(n13964), .A(n11883), .ZN(n15953) );
  AOI211_X1 U14491 ( .C1(n15901), .C2(n11885), .A(n11884), .B(n15953), .ZN(
        n11886) );
  MUX2_X1 U14492 ( .A(n11887), .B(n11886), .S(n15921), .Z(n11888) );
  OAI21_X1 U14493 ( .B1(n13852), .B2(n15949), .A(n11888), .ZN(P3_U3226) );
  NOR2_X1 U14494 ( .A1(n11919), .A2(n11889), .ZN(n11924) );
  NOR2_X1 U14495 ( .A1(n11924), .A2(n11890), .ZN(n11891) );
  XNOR2_X1 U14496 ( .A(n11891), .B(n13541), .ZN(n11892) );
  AOI222_X1 U14497 ( .A1(n13584), .A2(n13889), .B1(n13960), .B2(n11892), .C1(
        n13582), .C2(n13886), .ZN(n12115) );
  XNOR2_X1 U14498 ( .A(n11893), .B(n13541), .ZN(n12114) );
  INV_X1 U14499 ( .A(n14021), .ZN(n14004) );
  NAND2_X1 U14500 ( .A1(n12114), .A2(n14004), .ZN(n11895) );
  INV_X1 U14501 ( .A(n12119), .ZN(n12109) );
  AOI22_X1 U14502 ( .A1(n14018), .A2(n12109), .B1(P3_REG0_REG_10__SCAN_IN), 
        .B2(n15960), .ZN(n11894) );
  OAI211_X1 U14503 ( .C1(n15960), .C2(n12115), .A(n11895), .B(n11894), .ZN(
        P3_U3420) );
  INV_X1 U14504 ( .A(n11896), .ZN(n11898) );
  AND2_X1 U14505 ( .A1(n11898), .A2(n11897), .ZN(n11899) );
  XNOR2_X1 U14506 ( .A(n14668), .B(n7818), .ZN(n11902) );
  NAND2_X1 U14507 ( .A1(n14508), .A2(n14236), .ZN(n11903) );
  NAND2_X1 U14508 ( .A1(n11902), .A2(n11903), .ZN(n12141) );
  INV_X1 U14509 ( .A(n11902), .ZN(n11905) );
  INV_X1 U14510 ( .A(n11903), .ZN(n11904) );
  NAND2_X1 U14511 ( .A1(n11905), .A2(n11904), .ZN(n11906) );
  AND2_X1 U14512 ( .A1(n12141), .A2(n11906), .ZN(n11907) );
  NAND2_X1 U14513 ( .A1(n11908), .A2(n11907), .ZN(n12142) );
  OAI21_X1 U14514 ( .B1(n11908), .B2(n11907), .A(n12142), .ZN(n11909) );
  NAND2_X1 U14515 ( .A1(n11909), .A2(n14161), .ZN(n11917) );
  INV_X1 U14516 ( .A(n11910), .ZN(n11911) );
  NAND2_X1 U14517 ( .A1(n14194), .A2(n11911), .ZN(n11913) );
  OAI211_X1 U14518 ( .C1(n11914), .C2(n14196), .A(n11913), .B(n11912), .ZN(
        n11915) );
  AOI21_X1 U14519 ( .B1(n14668), .B2(n14211), .A(n11915), .ZN(n11916) );
  NAND2_X1 U14520 ( .A1(n11917), .A2(n11916), .ZN(P2_U3193) );
  INV_X1 U14521 ( .A(n11920), .ZN(n13537) );
  XNOR2_X1 U14522 ( .A(n11918), .B(n13537), .ZN(n11992) );
  INV_X1 U14523 ( .A(n11992), .ZN(n11933) );
  INV_X1 U14524 ( .A(n11919), .ZN(n11922) );
  AOI21_X1 U14525 ( .B1(n11922), .B2(n11921), .A(n11920), .ZN(n11923) );
  NOR3_X1 U14526 ( .A1(n11924), .A2(n11923), .A3(n15911), .ZN(n11927) );
  OAI22_X1 U14527 ( .A1(n12304), .A2(n15916), .B1(n15914), .B2(n11925), .ZN(
        n11926) );
  AOI211_X1 U14528 ( .C1(n11992), .C2(n12708), .A(n11927), .B(n11926), .ZN(
        n11990) );
  MUX2_X1 U14529 ( .A(n11928), .B(n11990), .S(n15921), .Z(n11931) );
  AOI22_X1 U14530 ( .A1(n13880), .A2(n11993), .B1(n15901), .B2(n11929), .ZN(
        n11930) );
  OAI211_X1 U14531 ( .C1(n11933), .C2(n11932), .A(n11931), .B(n11930), .ZN(
        P3_U3224) );
  INV_X1 U14532 ( .A(n11934), .ZN(n11936) );
  OAI222_X1 U14533 ( .A1(n7283), .A2(P3_U3151), .B1(n14040), .B2(n11936), .C1(
        n11935), .C2(n14033), .ZN(P3_U3271) );
  NAND2_X1 U14534 ( .A1(n12475), .A2(n11937), .ZN(n11938) );
  NAND2_X1 U14535 ( .A1(n11939), .A2(n11938), .ZN(n12207) );
  INV_X1 U14536 ( .A(n12207), .ZN(n11940) );
  XNOR2_X1 U14537 ( .A(n14778), .B(n14952), .ZN(n12641) );
  INV_X1 U14538 ( .A(n14952), .ZN(n11941) );
  OR2_X1 U14539 ( .A1(n14778), .A2(n11941), .ZN(n11943) );
  NAND2_X1 U14540 ( .A1(n12205), .A2(n11943), .ZN(n11942) );
  XNOR2_X1 U14541 ( .A(n14891), .B(n14951), .ZN(n12642) );
  NAND2_X1 U14542 ( .A1(n11942), .A2(n12642), .ZN(n12021) );
  INV_X1 U14543 ( .A(n12642), .ZN(n11950) );
  NAND3_X1 U14544 ( .A1(n12205), .A2(n11950), .A3(n11943), .ZN(n11944) );
  AND3_X1 U14545 ( .A1(n12021), .A2(n15763), .A3(n11944), .ZN(n11947) );
  OR2_X1 U14546 ( .A1(n14873), .A2(n14913), .ZN(n11946) );
  NAND2_X1 U14547 ( .A1(n14952), .A2(n15637), .ZN(n11945) );
  NAND2_X1 U14548 ( .A1(n11946), .A2(n11945), .ZN(n14898) );
  NOR2_X1 U14549 ( .A1(n11947), .A2(n14898), .ZN(n15504) );
  OR2_X1 U14550 ( .A1(n14778), .A2(n14952), .ZN(n11949) );
  OR2_X1 U14551 ( .A1(n11951), .A2(n11950), .ZN(n11952) );
  NAND2_X1 U14552 ( .A1(n12017), .A2(n11952), .ZN(n15500) );
  NAND2_X1 U14553 ( .A1(n12211), .A2(n14891), .ZN(n11953) );
  NAND2_X1 U14554 ( .A1(n11953), .A2(n15678), .ZN(n11954) );
  OR2_X1 U14555 ( .A1(n11954), .A2(n12026), .ZN(n15501) );
  OAI22_X1 U14556 ( .A1(n15714), .A2(n11955), .B1(n14895), .B2(n15712), .ZN(
        n11956) );
  AOI21_X1 U14557 ( .B1(n14891), .B2(n15716), .A(n11956), .ZN(n11957) );
  OAI21_X1 U14558 ( .B1(n15501), .B2(n15686), .A(n11957), .ZN(n11958) );
  AOI21_X1 U14559 ( .B1(n15500), .B2(n15688), .A(n11958), .ZN(n11959) );
  OAI21_X1 U14560 ( .B1(n15504), .B2(n6546), .A(n11959), .ZN(P1_U3282) );
  INV_X1 U14561 ( .A(n13608), .ZN(n11960) );
  AOI21_X1 U14562 ( .B1(n12053), .B2(n6753), .A(n11960), .ZN(n11972) );
  OAI21_X1 U14563 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n11962), .A(n11961), 
        .ZN(n11970) );
  NAND2_X1 U14564 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n12302)
         );
  NAND2_X1 U14565 ( .A1(n15894), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n11963) );
  OAI211_X1 U14566 ( .C1(n13746), .C2(n11964), .A(n12302), .B(n11963), .ZN(
        n11969) );
  AOI21_X1 U14567 ( .B1(n11966), .B2(n11965), .A(n6755), .ZN(n11967) );
  NOR2_X1 U14568 ( .A1(n11967), .A2(n13720), .ZN(n11968) );
  AOI211_X1 U14569 ( .C1(n13754), .C2(n11970), .A(n11969), .B(n11968), .ZN(
        n11971) );
  OAI21_X1 U14570 ( .B1(n11972), .B2(n13757), .A(n11971), .ZN(P3_U3193) );
  XNOR2_X1 U14571 ( .A(n12198), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n12193) );
  INV_X1 U14572 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n14627) );
  XNOR2_X1 U14573 ( .A(n12341), .B(n14627), .ZN(n12342) );
  XNOR2_X1 U14574 ( .A(n12343), .B(n12342), .ZN(n11989) );
  NAND2_X1 U14575 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n14126)
         );
  OAI21_X1 U14576 ( .B1(n15806), .B2(n11976), .A(n14126), .ZN(n11977) );
  AOI21_X1 U14577 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(n15809), .A(n11977), 
        .ZN(n11988) );
  NAND2_X1 U14578 ( .A1(n11978), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n11982) );
  NAND2_X1 U14579 ( .A1(n11980), .A2(n11979), .ZN(n11981) );
  NAND2_X1 U14580 ( .A1(n11982), .A2(n11981), .ZN(n12191) );
  INV_X1 U14581 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n14491) );
  MUX2_X1 U14582 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n14491), .S(n12198), .Z(
        n12192) );
  NAND2_X1 U14583 ( .A1(n12198), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n11985) );
  INV_X1 U14584 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n14471) );
  MUX2_X1 U14585 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n14471), .S(n12341), .Z(
        n11983) );
  MUX2_X1 U14586 ( .A(n14471), .B(P2_REG2_REG_17__SCAN_IN), .S(n12341), .Z(
        n11984) );
  NAND3_X1 U14587 ( .A1(n12190), .A2(n11985), .A3(n11984), .ZN(n11986) );
  NAND3_X1 U14588 ( .A1(n12336), .A2(n15811), .A3(n11986), .ZN(n11987) );
  OAI211_X1 U14589 ( .C1(n11989), .C2(n15825), .A(n11988), .B(n11987), .ZN(
        P2_U3231) );
  INV_X1 U14590 ( .A(n11990), .ZN(n11991) );
  AOI21_X1 U14591 ( .B1(n15957), .B2(n11992), .A(n11991), .ZN(n12153) );
  AOI22_X1 U14592 ( .A1(n14018), .A2(n11993), .B1(P3_REG0_REG_9__SCAN_IN), 
        .B2(n15960), .ZN(n11994) );
  OAI21_X1 U14593 ( .B1(n12153), .B2(n15960), .A(n11994), .ZN(P3_U3417) );
  NOR2_X1 U14594 ( .A1(n12414), .A2(n15742), .ZN(n15778) );
  OR2_X1 U14595 ( .A1(n12418), .A2(n14922), .ZN(n11996) );
  NAND2_X1 U14596 ( .A1(n14954), .A2(n15636), .ZN(n11995) );
  NAND2_X1 U14597 ( .A1(n11996), .A2(n11995), .ZN(n15777) );
  NAND2_X1 U14598 ( .A1(n15641), .A2(n15777), .ZN(n11997) );
  OAI211_X1 U14599 ( .C1(n15646), .C2(n15697), .A(n11998), .B(n11997), .ZN(
        n12004) );
  INV_X1 U14600 ( .A(n11999), .ZN(n12000) );
  AOI211_X1 U14601 ( .C1(n12002), .C2(n12001), .A(n15634), .B(n12000), .ZN(
        n12003) );
  AOI211_X1 U14602 ( .C1(n15632), .C2(n15778), .A(n12004), .B(n12003), .ZN(
        n12005) );
  INV_X1 U14603 ( .A(n12005), .ZN(P1_U3213) );
  NOR2_X1 U14604 ( .A1(n12006), .A2(n14564), .ZN(n12013) );
  INV_X1 U14605 ( .A(n12007), .ZN(n12008) );
  NOR2_X1 U14606 ( .A1(n14330), .A2(n12008), .ZN(n12012) );
  NOR2_X1 U14607 ( .A1(n14563), .A2(n12009), .ZN(n12011) );
  OAI22_X1 U14608 ( .A1(n15850), .A2(n10641), .B1(n14248), .B2(n15843), .ZN(
        n12010) );
  NOR4_X1 U14609 ( .A1(n12013), .A2(n12012), .A3(n12011), .A4(n12010), .ZN(
        n12014) );
  OAI21_X1 U14610 ( .B1(n12015), .B2(n14499), .A(n12014), .ZN(P2_U3264) );
  OR2_X1 U14611 ( .A1(n14891), .A2(n14951), .ZN(n12016) );
  XNOR2_X1 U14612 ( .A(n15497), .B(n14873), .ZN(n12644) );
  OAI21_X1 U14613 ( .B1(n12018), .B2(n12644), .A(n13010), .ZN(n12019) );
  INV_X1 U14614 ( .A(n12019), .ZN(n15499) );
  INV_X1 U14615 ( .A(n12644), .ZN(n12023) );
  OR2_X1 U14616 ( .A1(n14891), .A2(n12487), .ZN(n12020) );
  NAND2_X1 U14617 ( .A1(n12021), .A2(n12020), .ZN(n12022) );
  NAND2_X1 U14618 ( .A1(n12022), .A2(n12023), .ZN(n13043) );
  OAI211_X1 U14619 ( .C1(n12023), .C2(n12022), .A(n13043), .B(n15763), .ZN(
        n12025) );
  AND2_X1 U14620 ( .A1(n14951), .A2(n15637), .ZN(n12024) );
  AOI21_X1 U14621 ( .B1(n14949), .B2(n15636), .A(n12024), .ZN(n14810) );
  NAND2_X1 U14622 ( .A1(n12025), .A2(n14810), .ZN(n15495) );
  NAND2_X1 U14623 ( .A1(n15495), .A2(n15714), .ZN(n12032) );
  INV_X1 U14624 ( .A(n12026), .ZN(n12027) );
  AOI211_X1 U14625 ( .C1(n15497), .C2(n12027), .A(n15733), .B(n15360), .ZN(
        n15496) );
  INV_X1 U14626 ( .A(n12028), .ZN(n14812) );
  AOI22_X1 U14627 ( .A1(n6546), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n14812), 
        .B2(n15698), .ZN(n12029) );
  OAI21_X1 U14628 ( .B1(n7298), .B2(n15367), .A(n12029), .ZN(n12030) );
  AOI21_X1 U14629 ( .B1(n15496), .B2(n15720), .A(n12030), .ZN(n12031) );
  OAI211_X1 U14630 ( .C1(n15198), .C2(n15499), .A(n12032), .B(n12031), .ZN(
        P1_U3281) );
  XNOR2_X1 U14631 ( .A(n12695), .B(n12119), .ZN(n12224) );
  XNOR2_X1 U14632 ( .A(n12224), .B(n12304), .ZN(n12038) );
  INV_X1 U14633 ( .A(n12033), .ZN(n12035) );
  NAND2_X1 U14634 ( .A1(n12035), .A2(n12034), .ZN(n12039) );
  AND2_X1 U14635 ( .A1(n12038), .A2(n12039), .ZN(n12036) );
  NAND2_X1 U14636 ( .A1(n12225), .A2(n13325), .ZN(n12045) );
  AOI21_X1 U14637 ( .B1(n12037), .B2(n12039), .A(n12038), .ZN(n12044) );
  AOI22_X1 U14638 ( .A1(n13263), .A2(n13584), .B1(n13349), .B2(n13582), .ZN(
        n12041) );
  OAI211_X1 U14639 ( .C1(n13333), .C2(n12119), .A(n12041), .B(n12040), .ZN(
        n12042) );
  AOI21_X1 U14640 ( .B1(n12108), .B2(n13354), .A(n12042), .ZN(n12043) );
  OAI21_X1 U14641 ( .B1(n12045), .B2(n12044), .A(n12043), .ZN(P3_U3157) );
  OAI21_X1 U14642 ( .B1(n12047), .B2(n13453), .A(n12046), .ZN(n13946) );
  INV_X1 U14643 ( .A(n13946), .ZN(n12056) );
  INV_X1 U14644 ( .A(n13949), .ZN(n12048) );
  AOI22_X1 U14645 ( .A1(n13880), .A2(n12048), .B1(n15901), .B2(n12307), .ZN(
        n12055) );
  NOR2_X1 U14646 ( .A1(n12049), .A2(n13453), .ZN(n12092) );
  AND2_X1 U14647 ( .A1(n12049), .A2(n13453), .ZN(n12050) );
  OR2_X1 U14648 ( .A1(n12092), .A2(n12050), .ZN(n12052) );
  OAI22_X1 U14649 ( .A1(n12304), .A2(n15914), .B1(n15916), .B2(n12237), .ZN(
        n12051) );
  AOI21_X1 U14650 ( .B1(n12052), .B2(n13960), .A(n12051), .ZN(n13947) );
  MUX2_X1 U14651 ( .A(n12053), .B(n13947), .S(n15921), .Z(n12054) );
  OAI211_X1 U14652 ( .C1(n12056), .C2(n13894), .A(n12055), .B(n12054), .ZN(
        P3_U3222) );
  OR2_X1 U14653 ( .A1(n12057), .A2(n12973), .ZN(n12058) );
  NAND2_X1 U14654 ( .A1(n12059), .A2(n12058), .ZN(n12404) );
  OR2_X1 U14655 ( .A1(n12404), .A2(n14552), .ZN(n12067) );
  NAND2_X1 U14656 ( .A1(n12061), .A2(n12973), .ZN(n12062) );
  NAND2_X1 U14657 ( .A1(n12060), .A2(n12062), .ZN(n12065) );
  OR2_X1 U14658 ( .A1(n12820), .A2(n14202), .ZN(n12064) );
  NAND2_X1 U14659 ( .A1(n14233), .A2(n14193), .ZN(n12063) );
  NAND2_X1 U14660 ( .A1(n12064), .A2(n12063), .ZN(n12185) );
  AOI21_X1 U14661 ( .B1(n12065), .B2(n14556), .A(n12185), .ZN(n12066) );
  NAND2_X1 U14662 ( .A1(n12067), .A2(n12066), .ZN(n12398) );
  NOR2_X1 U14663 ( .A1(n12404), .A2(n14673), .ZN(n12071) );
  OAI21_X1 U14664 ( .B1(n6592), .B2(n12816), .A(n10836), .ZN(n12069) );
  NOR2_X1 U14665 ( .A1(n12069), .A2(n12068), .ZN(n12402) );
  AND2_X1 U14666 ( .A1(n12818), .A2(n10017), .ZN(n12070) );
  NOR4_X1 U14667 ( .A1(n12398), .A2(n12071), .A3(n12402), .A4(n12070), .ZN(
        n12074) );
  NAND2_X1 U14668 ( .A1(n15890), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n12072) );
  OAI21_X1 U14669 ( .B1(n12074), .B2(n15890), .A(n12072), .ZN(P2_U3509) );
  NAND2_X1 U14670 ( .A1(n15885), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n12073) );
  OAI21_X1 U14671 ( .B1(n12074), .B2(n15885), .A(n12073), .ZN(P2_U3460) );
  INV_X1 U14672 ( .A(n12075), .ZN(n12076) );
  AOI21_X1 U14673 ( .B1(n12078), .B2(n12077), .A(n12076), .ZN(n12085) );
  INV_X1 U14674 ( .A(n13319), .ZN(n13282) );
  AOI22_X1 U14675 ( .A1(n13263), .A2(n13590), .B1(n13282), .B2(n13588), .ZN(
        n12080) );
  OAI211_X1 U14676 ( .C1(n13333), .C2(n12081), .A(n12080), .B(n12079), .ZN(
        n12082) );
  AOI21_X1 U14677 ( .B1(n12083), .B2(n13354), .A(n12082), .ZN(n12084) );
  OAI21_X1 U14678 ( .B1(n12085), .B2(n13360), .A(n12084), .ZN(P3_U3170) );
  XNOR2_X1 U14679 ( .A(n12086), .B(n13542), .ZN(n12266) );
  NAND2_X1 U14680 ( .A1(n13542), .A2(n12087), .ZN(n12091) );
  INV_X1 U14681 ( .A(n12087), .ZN(n12089) );
  OAI21_X1 U14682 ( .B1(n12092), .B2(n12089), .A(n12088), .ZN(n12090) );
  OAI211_X1 U14683 ( .C1(n12092), .C2(n12091), .A(n12090), .B(n13960), .ZN(
        n12094) );
  NAND2_X1 U14684 ( .A1(n13889), .A2(n13582), .ZN(n12093) );
  OAI211_X1 U14685 ( .C1(n12332), .C2(n15916), .A(n12094), .B(n12093), .ZN(
        n12262) );
  OAI22_X1 U14686 ( .A1(n12362), .A2(n14013), .B1(n15959), .B2(n12095), .ZN(
        n12096) );
  AOI21_X1 U14687 ( .B1(n12262), .B2(n15959), .A(n12096), .ZN(n12097) );
  OAI21_X1 U14688 ( .B1(n12266), .B2(n14021), .A(n12097), .ZN(P3_U3426) );
  INV_X1 U14689 ( .A(n12098), .ZN(n12102) );
  OAI222_X1 U14690 ( .A1(n12100), .A2(P1_U3086), .B1(n10985), .B2(n12102), 
        .C1(n12099), .C2(n15546), .ZN(P1_U3330) );
  OAI222_X1 U14691 ( .A1(n13196), .A2(n12103), .B1(n13198), .B2(n12102), .C1(
        n12101), .C2(P2_U3088), .ZN(P2_U3302) );
  AOI22_X1 U14692 ( .A1(n13880), .A2(n12264), .B1(n15901), .B2(n12359), .ZN(
        n12107) );
  INV_X1 U14693 ( .A(n12262), .ZN(n12104) );
  MUX2_X1 U14694 ( .A(n12105), .B(n12104), .S(n15921), .Z(n12106) );
  OAI211_X1 U14695 ( .C1(n12266), .C2(n13894), .A(n12107), .B(n12106), .ZN(
        P3_U3221) );
  INV_X1 U14696 ( .A(n12114), .ZN(n12113) );
  AOI22_X1 U14697 ( .A1(n13880), .A2(n12109), .B1(n15901), .B2(n12108), .ZN(
        n12112) );
  MUX2_X1 U14698 ( .A(n12110), .B(n12115), .S(n15921), .Z(n12111) );
  OAI211_X1 U14699 ( .C1(n12113), .C2(n13894), .A(n12112), .B(n12111), .ZN(
        P3_U3223) );
  INV_X1 U14700 ( .A(n13945), .ZN(n13928) );
  NAND2_X1 U14701 ( .A1(n12114), .A2(n13928), .ZN(n12118) );
  MUX2_X1 U14702 ( .A(n12116), .B(n12115), .S(n15976), .Z(n12117) );
  OAI211_X1 U14703 ( .C1(n13940), .C2(n12119), .A(n12118), .B(n12117), .ZN(
        P3_U3469) );
  INV_X1 U14704 ( .A(n12120), .ZN(n12122) );
  INV_X1 U14705 ( .A(SI_25_), .ZN(n12121) );
  OAI222_X1 U14706 ( .A1(P3_U3151), .A2(n12123), .B1(n14040), .B2(n12122), 
        .C1(n12121), .C2(n14033), .ZN(P3_U3270) );
  INV_X1 U14707 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n12130) );
  XNOR2_X1 U14708 ( .A(n12130), .B(P1_ADDR_REG_11__SCAN_IN), .ZN(n12273) );
  XNOR2_X1 U14709 ( .A(n12274), .B(n12273), .ZN(n12132) );
  INV_X1 U14710 ( .A(n12131), .ZN(n12134) );
  INV_X1 U14711 ( .A(n12132), .ZN(n12133) );
  NAND2_X1 U14712 ( .A1(n12270), .A2(n12271), .ZN(n12135) );
  XNOR2_X1 U14713 ( .A(n12135), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  XNOR2_X1 U14714 ( .A(n14663), .B(n7818), .ZN(n12136) );
  OR2_X1 U14715 ( .A1(n12820), .A2(n13148), .ZN(n12137) );
  NAND2_X1 U14716 ( .A1(n12136), .A2(n12137), .ZN(n12183) );
  INV_X1 U14717 ( .A(n12136), .ZN(n12139) );
  INV_X1 U14718 ( .A(n12137), .ZN(n12138) );
  NAND2_X1 U14719 ( .A1(n12139), .A2(n12138), .ZN(n12140) );
  AND2_X1 U14720 ( .A1(n12183), .A2(n12140), .ZN(n12144) );
  NAND2_X1 U14721 ( .A1(n12142), .A2(n12141), .ZN(n12143) );
  OAI21_X1 U14722 ( .B1(n12144), .B2(n12143), .A(n12184), .ZN(n12151) );
  AOI21_X1 U14723 ( .B1(n14206), .B2(n12146), .A(n12145), .ZN(n12148) );
  NAND2_X1 U14724 ( .A1(n14663), .A2(n14211), .ZN(n12147) );
  OAI211_X1 U14725 ( .C1(n14209), .C2(n12149), .A(n12148), .B(n12147), .ZN(
        n12150) );
  AOI21_X1 U14726 ( .B1(n12151), .B2(n14161), .A(n12150), .ZN(n12152) );
  INV_X1 U14727 ( .A(n12152), .ZN(P2_U3203) );
  MUX2_X1 U14728 ( .A(n12154), .B(n12153), .S(n15976), .Z(n12155) );
  OAI21_X1 U14729 ( .B1(n13940), .B2(n12156), .A(n12155), .ZN(P3_U3468) );
  XNOR2_X1 U14730 ( .A(n12157), .B(n12975), .ZN(n12168) );
  OAI22_X1 U14731 ( .A1(n12817), .A2(n14202), .B1(n14152), .B2(n14204), .ZN(
        n14175) );
  INV_X1 U14732 ( .A(n12975), .ZN(n12160) );
  NAND3_X1 U14733 ( .A1(n12060), .A2(n12160), .A3(n12159), .ZN(n12161) );
  AOI21_X1 U14734 ( .B1(n12158), .B2(n12161), .A(n14534), .ZN(n12162) );
  AOI211_X1 U14735 ( .C1(n12168), .C2(n12163), .A(n14175), .B(n12162), .ZN(
        n14660) );
  INV_X1 U14736 ( .A(n12068), .ZN(n12165) );
  INV_X1 U14737 ( .A(n14558), .ZN(n12164) );
  AOI211_X1 U14738 ( .C1(n14658), .C2(n12165), .A(n14635), .B(n12164), .ZN(
        n14657) );
  INV_X1 U14739 ( .A(n14177), .ZN(n12166) );
  AOI22_X1 U14740 ( .A1(n14499), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n12166), 
        .B2(n14560), .ZN(n12167) );
  OAI21_X1 U14741 ( .B1(n12815), .B2(n14563), .A(n12167), .ZN(n12170) );
  INV_X1 U14742 ( .A(n12168), .ZN(n14661) );
  NOR2_X1 U14743 ( .A1(n14661), .A2(n14564), .ZN(n12169) );
  AOI211_X1 U14744 ( .C1(n14657), .C2(n14567), .A(n12170), .B(n12169), .ZN(
        n12171) );
  OAI21_X1 U14745 ( .B1(n14499), .B2(n14660), .A(n12171), .ZN(P2_U3254) );
  MUX2_X1 U14746 ( .A(n12173), .B(n13586), .S(n12172), .Z(n12174) );
  XOR2_X1 U14747 ( .A(n12175), .B(n12174), .Z(n12182) );
  AOI22_X1 U14748 ( .A1(n13263), .A2(n13586), .B1(n13282), .B2(n13584), .ZN(
        n12177) );
  OAI211_X1 U14749 ( .C1(n12178), .C2(n13333), .A(n12177), .B(n12176), .ZN(
        n12179) );
  AOI21_X1 U14750 ( .B1(n12180), .B2(n13354), .A(n12179), .ZN(n12181) );
  OAI21_X1 U14751 ( .B1(n12182), .B2(n13360), .A(n12181), .ZN(P3_U3161) );
  XNOR2_X1 U14752 ( .A(n12818), .B(n13166), .ZN(n13091) );
  NOR2_X1 U14753 ( .A1(n12817), .A2(n13148), .ZN(n13090) );
  XNOR2_X1 U14754 ( .A(n13091), .B(n13090), .ZN(n13089) );
  XNOR2_X1 U14755 ( .A(n13088), .B(n13089), .ZN(n12189) );
  NAND2_X1 U14756 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n15821)
         );
  NAND2_X1 U14757 ( .A1(n14206), .A2(n12185), .ZN(n12186) );
  OAI211_X1 U14758 ( .C1(n14209), .C2(n12400), .A(n15821), .B(n12186), .ZN(
        n12187) );
  AOI21_X1 U14759 ( .B1(n12818), .B2(n14211), .A(n12187), .ZN(n12188) );
  OAI21_X1 U14760 ( .B1(n12189), .B2(n14213), .A(n12188), .ZN(P2_U3189) );
  INV_X1 U14761 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n12201) );
  OAI211_X1 U14762 ( .C1(n12192), .C2(n12191), .A(n12190), .B(n15811), .ZN(
        n12200) );
  NAND2_X1 U14763 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n14118)
         );
  XOR2_X1 U14764 ( .A(n12194), .B(n12193), .Z(n12195) );
  NAND2_X1 U14765 ( .A1(n15815), .A2(n12195), .ZN(n12196) );
  NAND2_X1 U14766 ( .A1(n14118), .A2(n12196), .ZN(n12197) );
  AOI21_X1 U14767 ( .B1(n15831), .B2(n12198), .A(n12197), .ZN(n12199) );
  OAI211_X1 U14768 ( .C1(n15840), .C2(n12201), .A(n12200), .B(n12199), .ZN(
        P2_U3230) );
  OAI21_X1 U14769 ( .B1(n12203), .B2(n12208), .A(n12202), .ZN(n12204) );
  INV_X1 U14770 ( .A(n12204), .ZN(n15510) );
  INV_X1 U14771 ( .A(n12205), .ZN(n12206) );
  AOI211_X1 U14772 ( .C1(n12208), .C2(n12207), .A(n15709), .B(n12206), .ZN(
        n15508) );
  NAND2_X1 U14773 ( .A1(n14953), .A2(n15637), .ZN(n14780) );
  INV_X1 U14774 ( .A(n14780), .ZN(n12209) );
  OAI21_X1 U14775 ( .B1(n15508), .B2(n12209), .A(n15714), .ZN(n12217) );
  OAI22_X1 U14776 ( .A1(n15714), .A2(n12210), .B1(n14783), .B2(n15712), .ZN(
        n12215) );
  AOI211_X1 U14777 ( .C1(n14778), .C2(n12212), .A(n15733), .B(n7988), .ZN(
        n15506) );
  INV_X1 U14778 ( .A(n15506), .ZN(n12213) );
  NAND2_X1 U14779 ( .A1(n14951), .A2(n15636), .ZN(n14781) );
  AOI21_X1 U14780 ( .B1(n12213), .B2(n14781), .A(n15686), .ZN(n12214) );
  AOI211_X1 U14781 ( .C1(n15716), .C2(n14778), .A(n12215), .B(n12214), .ZN(
        n12216) );
  OAI211_X1 U14782 ( .C1(n15510), .C2(n15374), .A(n12217), .B(n12216), .ZN(
        P1_U3283) );
  INV_X1 U14783 ( .A(n12218), .ZN(n12222) );
  OAI222_X1 U14784 ( .A1(P1_U3086), .A2(n12220), .B1(n10985), .B2(n12222), 
        .C1(n12219), .C2(n15546), .ZN(P1_U3329) );
  OAI222_X1 U14785 ( .A1(n12223), .A2(P2_U3088), .B1(n13198), .B2(n12222), 
        .C1(n12221), .C2(n13196), .ZN(P2_U3301) );
  XNOR2_X1 U14786 ( .A(n13949), .B(n12695), .ZN(n12297) );
  OR2_X1 U14787 ( .A1(n12297), .A2(n13582), .ZN(n12226) );
  XNOR2_X1 U14788 ( .A(n12264), .B(n12695), .ZN(n12230) );
  XNOR2_X1 U14789 ( .A(n12230), .B(n13581), .ZN(n12350) );
  NAND2_X1 U14790 ( .A1(n12297), .A2(n13582), .ZN(n12227) );
  AND2_X1 U14791 ( .A1(n12350), .A2(n12227), .ZN(n12228) );
  NAND2_X1 U14792 ( .A1(n12230), .A2(n12237), .ZN(n12231) );
  XNOR2_X1 U14793 ( .A(n12245), .B(n13261), .ZN(n12232) );
  AND2_X1 U14794 ( .A1(n12232), .A2(n12332), .ZN(n12325) );
  INV_X1 U14795 ( .A(n12325), .ZN(n12234) );
  INV_X1 U14796 ( .A(n12232), .ZN(n12233) );
  NAND2_X1 U14797 ( .A1(n12233), .A2(n13580), .ZN(n12327) );
  NAND2_X1 U14798 ( .A1(n12234), .A2(n12327), .ZN(n12235) );
  XNOR2_X1 U14799 ( .A(n12326), .B(n12235), .ZN(n12241) );
  NOR2_X1 U14800 ( .A1(n12245), .A2(n13333), .ZN(n12239) );
  NAND2_X1 U14801 ( .A1(n13349), .A2(n13579), .ZN(n12236) );
  NAND2_X1 U14802 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n13628)
         );
  OAI211_X1 U14803 ( .C1(n13352), .C2(n12237), .A(n12236), .B(n13628), .ZN(
        n12238) );
  AOI211_X1 U14804 ( .C1(n12255), .C2(n13354), .A(n12239), .B(n12238), .ZN(
        n12240) );
  OAI21_X1 U14805 ( .B1(n12241), .B2(n13360), .A(n12240), .ZN(P3_U3174) );
  NAND2_X1 U14806 ( .A1(n13459), .A2(n13460), .ZN(n13545) );
  XOR2_X1 U14807 ( .A(n13545), .B(n12242), .Z(n12243) );
  AOI222_X1 U14808 ( .A1(n13581), .A2(n13889), .B1(n13960), .B2(n12243), .C1(
        n13579), .C2(n13886), .ZN(n12261) );
  XNOR2_X1 U14809 ( .A(n12244), .B(n13545), .ZN(n12254) );
  NAND2_X1 U14810 ( .A1(n12254), .A2(n13928), .ZN(n12247) );
  INV_X1 U14811 ( .A(n12245), .ZN(n12258) );
  AOI22_X1 U14812 ( .A1(n13942), .A2(n12258), .B1(P3_REG1_REG_13__SCAN_IN), 
        .B2(n15973), .ZN(n12246) );
  OAI211_X1 U14813 ( .C1(n12261), .C2(n15973), .A(n12247), .B(n12246), .ZN(
        P3_U3472) );
  INV_X1 U14814 ( .A(n12248), .ZN(n12250) );
  OAI222_X1 U14815 ( .A1(n12251), .A2(P3_U3151), .B1(n14040), .B2(n12250), 
        .C1(n12249), .C2(n14033), .ZN(P3_U3269) );
  NAND2_X1 U14816 ( .A1(n12254), .A2(n14004), .ZN(n12253) );
  AOI22_X1 U14817 ( .A1(n14018), .A2(n12258), .B1(P3_REG0_REG_13__SCAN_IN), 
        .B2(n15960), .ZN(n12252) );
  OAI211_X1 U14818 ( .C1(n15960), .C2(n12261), .A(n12253), .B(n12252), .ZN(
        P3_U3429) );
  INV_X1 U14819 ( .A(n13894), .ZN(n13856) );
  NAND2_X1 U14820 ( .A1(n12254), .A2(n13856), .ZN(n12260) );
  INV_X1 U14821 ( .A(n12255), .ZN(n12256) );
  OAI22_X1 U14822 ( .A1(n15921), .A2(n13627), .B1(n12256), .B2(n15923), .ZN(
        n12257) );
  AOI21_X1 U14823 ( .B1(n12258), .B2(n13880), .A(n12257), .ZN(n12259) );
  OAI211_X1 U14824 ( .C1(n15903), .C2(n12261), .A(n12260), .B(n12259), .ZN(
        P3_U3220) );
  MUX2_X1 U14825 ( .A(P3_REG1_REG_12__SCAN_IN), .B(n12262), .S(n15976), .Z(
        n12263) );
  AOI21_X1 U14826 ( .B1(n13942), .B2(n12264), .A(n12263), .ZN(n12265) );
  OAI21_X1 U14827 ( .B1(n12266), .B2(n13945), .A(n12265), .ZN(P3_U3471) );
  INV_X1 U14828 ( .A(n12267), .ZN(n12283) );
  AOI21_X1 U14829 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n13080), .A(n12989), 
        .ZN(n12268) );
  OAI21_X1 U14830 ( .B1(n12283), .B2(n12667), .A(n12268), .ZN(P2_U3300) );
  NAND2_X1 U14831 ( .A1(n12270), .A2(n12269), .ZN(n12272) );
  NAND2_X1 U14832 ( .A1(n12275), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n12276) );
  XNOR2_X1 U14833 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n12290) );
  INV_X1 U14834 ( .A(n12290), .ZN(n12278) );
  XNOR2_X1 U14835 ( .A(n12291), .B(n12278), .ZN(n12279) );
  NAND2_X1 U14836 ( .A1(n12280), .A2(n12279), .ZN(n12289) );
  NAND2_X1 U14837 ( .A1(n12288), .A2(n12289), .ZN(n12281) );
  XNOR2_X1 U14838 ( .A(n12281), .B(P2_ADDR_REG_12__SCAN_IN), .ZN(SUB_1596_U68)
         );
  OAI222_X1 U14839 ( .A1(n7374), .A2(P1_U3086), .B1(n10985), .B2(n12283), .C1(
        n12282), .C2(n15546), .ZN(P1_U3328) );
  NAND2_X1 U14840 ( .A1(n13184), .A2(n13079), .ZN(n12285) );
  OAI211_X1 U14841 ( .C1(n13196), .C2(n12286), .A(n12285), .B(n12284), .ZN(
        P2_U3299) );
  INV_X1 U14842 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n12287) );
  NAND2_X1 U14843 ( .A1(n12291), .A2(n12290), .ZN(n12294) );
  NAND2_X1 U14844 ( .A1(n12292), .A2(P3_ADDR_REG_12__SCAN_IN), .ZN(n12293) );
  NAND2_X1 U14845 ( .A1(n12294), .A2(n12293), .ZN(n15568) );
  XNOR2_X1 U14846 ( .A(P1_ADDR_REG_13__SCAN_IN), .B(P3_ADDR_REG_13__SCAN_IN), 
        .ZN(n12295) );
  INV_X1 U14847 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15559) );
  XNOR2_X1 U14848 ( .A(n15560), .B(n15559), .ZN(n12296) );
  XNOR2_X1 U14849 ( .A(n15562), .B(n12296), .ZN(SUB_1596_U67) );
  INV_X1 U14850 ( .A(n12298), .ZN(n12300) );
  INV_X1 U14851 ( .A(n12297), .ZN(n12299) );
  OR2_X1 U14852 ( .A1(n12298), .A2(n12297), .ZN(n12349) );
  OAI21_X1 U14853 ( .B1(n12300), .B2(n12299), .A(n12349), .ZN(n12301) );
  NOR2_X1 U14854 ( .A1(n12301), .A2(n13582), .ZN(n12352) );
  AOI21_X1 U14855 ( .B1(n13582), .B2(n12301), .A(n12352), .ZN(n12309) );
  NOR2_X1 U14856 ( .A1(n13333), .A2(n13949), .ZN(n12306) );
  NAND2_X1 U14857 ( .A1(n13349), .A2(n13581), .ZN(n12303) );
  OAI211_X1 U14858 ( .C1(n13352), .C2(n12304), .A(n12303), .B(n12302), .ZN(
        n12305) );
  AOI211_X1 U14859 ( .C1(n12307), .C2(n13354), .A(n12306), .B(n12305), .ZN(
        n12308) );
  OAI21_X1 U14860 ( .B1(n12309), .B2(n13360), .A(n12308), .ZN(P3_U3176) );
  INV_X1 U14861 ( .A(n12310), .ZN(n12312) );
  OAI222_X1 U14862 ( .A1(n14040), .A2(n12312), .B1(n14033), .B2(n12311), .C1(
        P3_U3151), .C2(n7288), .ZN(P3_U3268) );
  NAND2_X1 U14863 ( .A1(n12313), .A2(n13460), .ZN(n12369) );
  XNOR2_X1 U14864 ( .A(n12369), .B(n13549), .ZN(n12368) );
  INV_X1 U14865 ( .A(n13465), .ZN(n12323) );
  NAND2_X1 U14866 ( .A1(n12314), .A2(n13549), .ZN(n12315) );
  NAND3_X1 U14867 ( .A1(n12316), .A2(n13960), .A3(n12315), .ZN(n12319) );
  OAI22_X1 U14868 ( .A1(n13344), .A2(n15916), .B1(n12332), .B2(n15914), .ZN(
        n12317) );
  INV_X1 U14869 ( .A(n12317), .ZN(n12318) );
  NAND2_X1 U14870 ( .A1(n12319), .A2(n12318), .ZN(n12363) );
  MUX2_X1 U14871 ( .A(P3_REG0_REG_14__SCAN_IN), .B(n12363), .S(n15959), .Z(
        n12320) );
  AOI21_X1 U14872 ( .B1(n14018), .B2(n12323), .A(n12320), .ZN(n12321) );
  OAI21_X1 U14873 ( .B1(n12368), .B2(n14021), .A(n12321), .ZN(P3_U3432) );
  MUX2_X1 U14874 ( .A(P3_REG1_REG_14__SCAN_IN), .B(n12363), .S(n15976), .Z(
        n12322) );
  AOI21_X1 U14875 ( .B1(n13942), .B2(n12323), .A(n12322), .ZN(n12324) );
  OAI21_X1 U14876 ( .B1(n12368), .B2(n13945), .A(n12324), .ZN(P3_U3473) );
  XNOR2_X1 U14877 ( .A(n13465), .B(n12695), .ZN(n12669) );
  XNOR2_X1 U14878 ( .A(n12669), .B(n13351), .ZN(n12328) );
  OAI211_X1 U14879 ( .C1(n12329), .C2(n12328), .A(n12671), .B(n13325), .ZN(
        n12335) );
  NAND2_X1 U14880 ( .A1(n13349), .A2(n12672), .ZN(n12331) );
  OAI211_X1 U14881 ( .C1(n13352), .C2(n12332), .A(n12331), .B(n12330), .ZN(
        n12333) );
  AOI21_X1 U14882 ( .B1(n12366), .B2(n13354), .A(n12333), .ZN(n12334) );
  OAI211_X1 U14883 ( .C1(n13333), .C2(n13465), .A(n12335), .B(n12334), .ZN(
        P3_U3155) );
  NAND2_X1 U14884 ( .A1(n12337), .A2(n14289), .ZN(n12338) );
  NAND2_X1 U14885 ( .A1(n14292), .A2(n12338), .ZN(n12340) );
  INV_X1 U14886 ( .A(n14293), .ZN(n12339) );
  AOI21_X1 U14887 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n12340), .A(n12339), 
        .ZN(n12348) );
  AOI22_X1 U14888 ( .A1(n12343), .A2(n12342), .B1(n12341), .B2(
        P2_REG1_REG_17__SCAN_IN), .ZN(n14287) );
  XOR2_X1 U14889 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14290), .Z(n12346) );
  NAND2_X1 U14890 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14185)
         );
  NAND2_X1 U14891 ( .A1(n15831), .A2(n14289), .ZN(n12344) );
  OAI211_X1 U14892 ( .C1(n15840), .C2(n7246), .A(n14185), .B(n12344), .ZN(
        n12345) );
  AOI21_X1 U14893 ( .B1(n12346), .B2(n15815), .A(n12345), .ZN(n12347) );
  OAI21_X1 U14894 ( .B1(n12348), .B2(n15832), .A(n12347), .ZN(P2_U3232) );
  INV_X1 U14895 ( .A(n12349), .ZN(n12351) );
  NOR3_X1 U14896 ( .A1(n12352), .A2(n12351), .A3(n12350), .ZN(n12355) );
  INV_X1 U14897 ( .A(n12353), .ZN(n12354) );
  OAI21_X1 U14898 ( .B1(n12355), .B2(n12354), .A(n13325), .ZN(n12361) );
  NAND2_X1 U14899 ( .A1(n13349), .A2(n13580), .ZN(n12356) );
  NAND2_X1 U14900 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n13611)
         );
  OAI211_X1 U14901 ( .C1(n13352), .C2(n12357), .A(n12356), .B(n13611), .ZN(
        n12358) );
  AOI21_X1 U14902 ( .B1(n12359), .B2(n13354), .A(n12358), .ZN(n12360) );
  OAI211_X1 U14903 ( .C1(n12362), .C2(n13333), .A(n12361), .B(n12360), .ZN(
        P3_U3164) );
  NOR2_X1 U14904 ( .A1(n13852), .A2(n13465), .ZN(n12365) );
  MUX2_X1 U14905 ( .A(n12363), .B(P3_REG2_REG_14__SCAN_IN), .S(n15903), .Z(
        n12364) );
  AOI211_X1 U14906 ( .C1(n15901), .C2(n12366), .A(n12365), .B(n12364), .ZN(
        n12367) );
  OAI21_X1 U14907 ( .B1(n12368), .B2(n13894), .A(n12367), .ZN(P3_U3219) );
  OAI21_X1 U14908 ( .B1(n12369), .B2(n7403), .A(n13462), .ZN(n12370) );
  XNOR2_X1 U14909 ( .A(n12370), .B(n13544), .ZN(n12382) );
  AOI22_X1 U14910 ( .A1(n13880), .A2(n13356), .B1(n15901), .B2(n13355), .ZN(
        n12376) );
  NAND2_X1 U14911 ( .A1(n13882), .A2(n13544), .ZN(n12385) );
  OAI211_X1 U14912 ( .C1(n13882), .C2(n13544), .A(n12385), .B(n13960), .ZN(
        n12373) );
  NOR2_X1 U14913 ( .A1(n13351), .A2(n15914), .ZN(n12371) );
  AOI21_X1 U14914 ( .B1(n13890), .B2(n13886), .A(n12371), .ZN(n12372) );
  NAND2_X1 U14915 ( .A1(n12373), .A2(n12372), .ZN(n12379) );
  MUX2_X1 U14916 ( .A(n12379), .B(P3_REG2_REG_15__SCAN_IN), .S(n15903), .Z(
        n12374) );
  INV_X1 U14917 ( .A(n12374), .ZN(n12375) );
  OAI211_X1 U14918 ( .C1(n12382), .C2(n13894), .A(n12376), .B(n12375), .ZN(
        P3_U3218) );
  MUX2_X1 U14919 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n12379), .S(n15959), .Z(
        n12377) );
  AOI21_X1 U14920 ( .B1(n14018), .B2(n13356), .A(n12377), .ZN(n12378) );
  OAI21_X1 U14921 ( .B1(n12382), .B2(n14021), .A(n12378), .ZN(P3_U3435) );
  MUX2_X1 U14922 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n12379), .S(n15976), .Z(
        n12380) );
  AOI21_X1 U14923 ( .B1(n13942), .B2(n13356), .A(n12380), .ZN(n12381) );
  OAI21_X1 U14924 ( .B1(n12382), .B2(n13945), .A(n12381), .ZN(P3_U3474) );
  XNOR2_X1 U14925 ( .A(n12383), .B(n12386), .ZN(n12397) );
  AOI22_X1 U14926 ( .A1(n13880), .A2(n13476), .B1(n15901), .B2(n13295), .ZN(
        n12390) );
  INV_X1 U14927 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13686) );
  NAND2_X1 U14928 ( .A1(n12385), .A2(n12384), .ZN(n12387) );
  INV_X1 U14929 ( .A(n12386), .ZN(n13548) );
  XNOR2_X1 U14930 ( .A(n12387), .B(n13548), .ZN(n12388) );
  AOI222_X1 U14931 ( .A1(n12388), .A2(n13960), .B1(n13578), .B2(n13886), .C1(
        n12672), .C2(n13889), .ZN(n12393) );
  MUX2_X1 U14932 ( .A(n13686), .B(n12393), .S(n15921), .Z(n12389) );
  OAI211_X1 U14933 ( .C1(n12397), .C2(n13894), .A(n12390), .B(n12389), .ZN(
        P3_U3217) );
  MUX2_X1 U14934 ( .A(n13671), .B(n12393), .S(n15976), .Z(n12392) );
  NAND2_X1 U14935 ( .A1(n13942), .A2(n13476), .ZN(n12391) );
  OAI211_X1 U14936 ( .C1(n12397), .C2(n13945), .A(n12392), .B(n12391), .ZN(
        P3_U3475) );
  INV_X1 U14937 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12394) );
  MUX2_X1 U14938 ( .A(n12394), .B(n12393), .S(n15959), .Z(n12396) );
  NAND2_X1 U14939 ( .A1(n14018), .A2(n13476), .ZN(n12395) );
  OAI211_X1 U14940 ( .C1(n12397), .C2(n14021), .A(n12396), .B(n12395), .ZN(
        P3_U3438) );
  MUX2_X1 U14941 ( .A(n12398), .B(P2_REG2_REG_10__SCAN_IN), .S(n14499), .Z(
        n12406) );
  NAND2_X1 U14942 ( .A1(n12818), .A2(n14541), .ZN(n12399) );
  OAI21_X1 U14943 ( .B1(n15843), .B2(n12400), .A(n12399), .ZN(n12401) );
  AOI21_X1 U14944 ( .B1(n12402), .B2(n14567), .A(n12401), .ZN(n12403) );
  OAI21_X1 U14945 ( .B1(n12404), .B2(n14564), .A(n12403), .ZN(n12405) );
  OR2_X1 U14946 ( .A1(n12406), .A2(n12405), .ZN(P2_U3255) );
  OAI222_X1 U14947 ( .A1(n12409), .A2(P2_U3088), .B1(n13198), .B2(n12408), 
        .C1(n12407), .C2(n13196), .ZN(P2_U3307) );
  NOR3_X1 U14948 ( .A1(n15517), .A2(n7374), .A3(n14922), .ZN(n12665) );
  OAI21_X1 U14949 ( .B1(n6809), .B2(n12656), .A(P1_B_REG_SCAN_IN), .ZN(n12664)
         );
  NAND2_X1 U14950 ( .A1(n12410), .A2(n15314), .ZN(n12411) );
  NAND2_X1 U14951 ( .A1(n12412), .A2(n12411), .ZN(n12596) );
  MUX2_X1 U14952 ( .A(n11112), .B(n12622), .S(n12596), .Z(n12413) );
  INV_X2 U14953 ( .A(n12433), .ZN(n12624) );
  MUX2_X1 U14954 ( .A(n13025), .B(n15400), .S(n12624), .Z(n12574) );
  MUX2_X1 U14955 ( .A(n12415), .B(n12414), .S(n6551), .Z(n12466) );
  MUX2_X1 U14956 ( .A(n14956), .B(n12416), .S(n12433), .Z(n12463) );
  INV_X1 U14957 ( .A(n12463), .ZN(n12420) );
  MUX2_X1 U14958 ( .A(n12418), .B(n12417), .S(n6551), .Z(n12464) );
  INV_X1 U14959 ( .A(n12464), .ZN(n12419) );
  NAND2_X1 U14960 ( .A1(n12420), .A2(n12419), .ZN(n12421) );
  NAND2_X1 U14961 ( .A1(n12466), .A2(n12421), .ZN(n12425) );
  MUX2_X1 U14962 ( .A(n14955), .B(n15702), .S(n6549), .Z(n12465) );
  INV_X1 U14963 ( .A(n12465), .ZN(n12424) );
  INV_X1 U14964 ( .A(n12421), .ZN(n12423) );
  INV_X1 U14965 ( .A(n12466), .ZN(n12422) );
  AOI22_X1 U14966 ( .A1(n12425), .A2(n12424), .B1(n12423), .B2(n12422), .ZN(
        n12474) );
  NAND3_X1 U14967 ( .A1(n12427), .A2(n6551), .A3(n12447), .ZN(n12437) );
  INV_X1 U14968 ( .A(n12434), .ZN(n12429) );
  NAND3_X1 U14969 ( .A1(n12430), .A2(n12429), .A3(n6551), .ZN(n12431) );
  NAND2_X1 U14970 ( .A1(n12434), .A2(n12433), .ZN(n12445) );
  MUX2_X1 U14971 ( .A(n6549), .B(n12445), .S(n12435), .Z(n12436) );
  NAND3_X1 U14972 ( .A1(n12437), .A2(n8103), .A3(n12436), .ZN(n12450) );
  NAND2_X1 U14973 ( .A1(n12439), .A2(n12438), .ZN(n12442) );
  NAND3_X1 U14974 ( .A1(n12442), .A2(n12441), .A3(n12440), .ZN(n12444) );
  NAND2_X1 U14975 ( .A1(n12444), .A2(n12443), .ZN(n12448) );
  INV_X1 U14976 ( .A(n12445), .ZN(n12446) );
  NAND3_X1 U14977 ( .A1(n12448), .A2(n12447), .A3(n12446), .ZN(n12449) );
  NAND2_X1 U14978 ( .A1(n12450), .A2(n12449), .ZN(n12453) );
  MUX2_X1 U14979 ( .A(n6540), .B(n15756), .S(n6551), .Z(n12454) );
  NAND2_X1 U14980 ( .A1(n12453), .A2(n12454), .ZN(n12452) );
  MUX2_X1 U14981 ( .A(n15756), .B(n6540), .S(n12624), .Z(n12451) );
  NAND2_X1 U14982 ( .A1(n12452), .A2(n12451), .ZN(n12458) );
  INV_X1 U14983 ( .A(n12453), .ZN(n12456) );
  INV_X1 U14984 ( .A(n12454), .ZN(n12455) );
  NAND2_X1 U14985 ( .A1(n12456), .A2(n12455), .ZN(n12457) );
  MUX2_X1 U14986 ( .A(n12459), .B(n6539), .S(n6551), .Z(n12461) );
  MUX2_X1 U14987 ( .A(n6539), .B(n12459), .S(n6551), .Z(n12460) );
  AOI22_X1 U14988 ( .A1(n12466), .A2(n12465), .B1(n12464), .B2(n12463), .ZN(
        n12467) );
  NAND2_X1 U14989 ( .A1(n12469), .A2(n12468), .ZN(n12473) );
  AND2_X1 U14990 ( .A1(n14954), .A2(n6549), .ZN(n12471) );
  OAI21_X1 U14991 ( .B1(n14954), .B2(n6549), .A(n15684), .ZN(n12470) );
  OAI21_X1 U14992 ( .B1(n12471), .B2(n15684), .A(n12470), .ZN(n12472) );
  MUX2_X1 U14993 ( .A(n14953), .B(n12475), .S(n12600), .Z(n12478) );
  MUX2_X1 U14994 ( .A(n14953), .B(n12475), .S(n6549), .Z(n12476) );
  INV_X1 U14995 ( .A(n12478), .ZN(n12479) );
  MUX2_X1 U14996 ( .A(n14952), .B(n14778), .S(n6549), .Z(n12483) );
  MUX2_X1 U14997 ( .A(n14952), .B(n14778), .S(n6551), .Z(n12480) );
  NAND2_X1 U14998 ( .A1(n12481), .A2(n12480), .ZN(n12485) );
  MUX2_X1 U14999 ( .A(n14951), .B(n14891), .S(n12600), .Z(n12489) );
  MUX2_X1 U15000 ( .A(n12487), .B(n12486), .S(n6549), .Z(n12488) );
  INV_X1 U15001 ( .A(n14873), .ZN(n14950) );
  MUX2_X1 U15002 ( .A(n14949), .B(n15491), .S(n6549), .Z(n12493) );
  MUX2_X1 U15003 ( .A(n14754), .B(n15368), .S(n12600), .Z(n12495) );
  AOI22_X1 U15004 ( .A1(n12493), .A2(n12495), .B1(n12492), .B2(n12491), .ZN(
        n12494) );
  INV_X1 U15005 ( .A(n12433), .ZN(n12600) );
  INV_X1 U15006 ( .A(n12495), .ZN(n12497) );
  NAND2_X1 U15007 ( .A1(n14949), .A2(n12600), .ZN(n12496) );
  OAI211_X1 U15008 ( .C1(n12600), .C2(n15368), .A(n12497), .B(n12496), .ZN(
        n12502) );
  AOI21_X1 U15009 ( .B1(n13051), .B2(n13048), .A(n12600), .ZN(n12500) );
  AOI21_X1 U15010 ( .B1(n12632), .B2(n13047), .A(n6549), .ZN(n12499) );
  NOR2_X1 U15011 ( .A1(n12500), .A2(n12499), .ZN(n12501) );
  MUX2_X1 U15012 ( .A(n14947), .B(n15472), .S(n12600), .Z(n12523) );
  NAND2_X1 U15013 ( .A1(n12523), .A2(n14946), .ZN(n12505) );
  INV_X1 U15014 ( .A(n14947), .ZN(n13052) );
  NAND2_X1 U15015 ( .A1(n13052), .A2(n12600), .ZN(n12507) );
  AOI21_X1 U15016 ( .B1(n12505), .B2(n12507), .A(n15466), .ZN(n12511) );
  NAND2_X1 U15017 ( .A1(n12523), .A2(n14831), .ZN(n12506) );
  OR2_X1 U15018 ( .A1(n15472), .A2(n6551), .ZN(n12518) );
  AOI21_X1 U15019 ( .B1(n12506), .B2(n12518), .A(n15303), .ZN(n12510) );
  NAND2_X1 U15020 ( .A1(n14946), .A2(n6549), .ZN(n12520) );
  OR2_X1 U15021 ( .A1(n15472), .A2(n12520), .ZN(n12509) );
  INV_X1 U15022 ( .A(n12507), .ZN(n12515) );
  NAND2_X1 U15023 ( .A1(n12515), .A2(n14831), .ZN(n12508) );
  NAND2_X1 U15024 ( .A1(n12509), .A2(n12508), .ZN(n12522) );
  OR3_X1 U15025 ( .A1(n12511), .A2(n12510), .A3(n12522), .ZN(n12513) );
  MUX2_X1 U15026 ( .A(n12632), .B(n13051), .S(n12624), .Z(n12512) );
  NAND2_X1 U15027 ( .A1(n12514), .A2(n8086), .ZN(n12527) );
  NAND2_X1 U15028 ( .A1(n12523), .A2(n12515), .ZN(n12516) );
  OAI21_X1 U15029 ( .B1(n14946), .B2(n6549), .A(n12516), .ZN(n12517) );
  NAND2_X1 U15030 ( .A1(n12517), .A2(n15303), .ZN(n12526) );
  INV_X1 U15031 ( .A(n12518), .ZN(n12519) );
  NAND2_X1 U15032 ( .A1(n12523), .A2(n12519), .ZN(n12521) );
  NAND2_X1 U15033 ( .A1(n12521), .A2(n12520), .ZN(n12524) );
  AOI22_X1 U15034 ( .A1(n12524), .A2(n15466), .B1(n12523), .B2(n12522), .ZN(
        n12525) );
  NAND3_X1 U15035 ( .A1(n12527), .A2(n12526), .A3(n12525), .ZN(n12528) );
  NAND2_X1 U15036 ( .A1(n15461), .A2(n14838), .ZN(n12529) );
  NAND2_X1 U15037 ( .A1(n12528), .A2(n15282), .ZN(n12531) );
  MUX2_X1 U15038 ( .A(n15244), .B(n12529), .S(n12624), .Z(n12530) );
  NAND2_X1 U15039 ( .A1(n12531), .A2(n12530), .ZN(n12532) );
  XNOR2_X1 U15040 ( .A(n15455), .B(n14944), .ZN(n15266) );
  NAND2_X1 U15041 ( .A1(n12532), .A2(n15266), .ZN(n12537) );
  XNOR2_X1 U15042 ( .A(n15447), .B(n14943), .ZN(n15245) );
  NAND2_X1 U15043 ( .A1(n14944), .A2(n6549), .ZN(n12534) );
  INV_X1 U15044 ( .A(n14944), .ZN(n13055) );
  NAND2_X1 U15045 ( .A1(n13055), .A2(n12600), .ZN(n12533) );
  MUX2_X1 U15046 ( .A(n12534), .B(n12533), .S(n15455), .Z(n12535) );
  AND2_X1 U15047 ( .A1(n15245), .A2(n12535), .ZN(n12536) );
  NAND2_X1 U15048 ( .A1(n12537), .A2(n12536), .ZN(n12541) );
  AND2_X1 U15049 ( .A1(n14943), .A2(n12600), .ZN(n12539) );
  OAI21_X1 U15050 ( .B1(n12600), .B2(n14943), .A(n15447), .ZN(n12538) );
  OAI21_X1 U15051 ( .B1(n12539), .B2(n15447), .A(n12538), .ZN(n12540) );
  MUX2_X1 U15052 ( .A(n14942), .B(n15443), .S(n6549), .Z(n12543) );
  MUX2_X1 U15053 ( .A(n14942), .B(n15443), .S(n12624), .Z(n12542) );
  INV_X1 U15054 ( .A(n12543), .ZN(n12544) );
  MUX2_X1 U15055 ( .A(n14941), .B(n15437), .S(n12624), .Z(n12548) );
  NAND2_X1 U15056 ( .A1(n12547), .A2(n12548), .ZN(n12546) );
  MUX2_X1 U15057 ( .A(n15437), .B(n14941), .S(n12624), .Z(n12545) );
  INV_X1 U15058 ( .A(n12547), .ZN(n12550) );
  INV_X1 U15059 ( .A(n12548), .ZN(n12549) );
  MUX2_X1 U15060 ( .A(n14940), .B(n15428), .S(n6549), .Z(n12552) );
  MUX2_X1 U15061 ( .A(n14940), .B(n15428), .S(n12624), .Z(n12551) );
  MUX2_X1 U15062 ( .A(n14939), .B(n15425), .S(n12624), .Z(n12555) );
  NAND2_X1 U15063 ( .A1(n12556), .A2(n12555), .ZN(n12554) );
  MUX2_X1 U15064 ( .A(n15425), .B(n14939), .S(n12624), .Z(n12553) );
  NAND2_X1 U15065 ( .A1(n12554), .A2(n12553), .ZN(n12558) );
  MUX2_X1 U15066 ( .A(n14938), .B(n14822), .S(n6549), .Z(n12560) );
  MUX2_X1 U15067 ( .A(n14938), .B(n14822), .S(n12624), .Z(n12559) );
  MUX2_X1 U15068 ( .A(n14937), .B(n15163), .S(n12624), .Z(n12564) );
  MUX2_X1 U15069 ( .A(n14937), .B(n15163), .S(n6549), .Z(n12561) );
  NAND2_X1 U15070 ( .A1(n12562), .A2(n12561), .ZN(n12568) );
  INV_X1 U15071 ( .A(n12563), .ZN(n12566) );
  INV_X1 U15072 ( .A(n12564), .ZN(n12565) );
  NAND2_X1 U15073 ( .A1(n12566), .A2(n12565), .ZN(n12567) );
  NAND2_X1 U15074 ( .A1(n12568), .A2(n12567), .ZN(n12570) );
  MUX2_X1 U15075 ( .A(n14936), .B(n15150), .S(n6549), .Z(n12571) );
  MUX2_X1 U15076 ( .A(n14936), .B(n15150), .S(n12600), .Z(n12569) );
  INV_X1 U15077 ( .A(n12571), .ZN(n12572) );
  MUX2_X1 U15078 ( .A(n15135), .B(n14935), .S(n12600), .Z(n12573) );
  OAI21_X1 U15079 ( .B1(n7294), .B2(n12576), .A(n12575), .ZN(n12604) );
  NAND2_X1 U15080 ( .A1(n13002), .A2(n12614), .ZN(n12578) );
  OR2_X1 U15081 ( .A1(n12615), .A2(n13003), .ZN(n12577) );
  MUX2_X1 U15082 ( .A(n14934), .B(n13032), .S(n6549), .Z(n12603) );
  NAND2_X1 U15083 ( .A1(n12583), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n12581) );
  NAND2_X1 U15084 ( .A1(n12579), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n12580) );
  OAI211_X1 U15085 ( .C1(n9927), .C2(n12582), .A(n12581), .B(n12580), .ZN(
        n15118) );
  INV_X1 U15086 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n12587) );
  NAND2_X1 U15087 ( .A1(n12583), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n12586) );
  NAND2_X1 U15088 ( .A1(n12579), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n12585) );
  OAI211_X1 U15089 ( .C1(n9927), .C2(n12587), .A(n12586), .B(n12585), .ZN(
        n14933) );
  OAI21_X1 U15090 ( .B1(n15118), .B2(n12588), .A(n14933), .ZN(n12594) );
  INV_X1 U15091 ( .A(SI_29_), .ZN(n14034) );
  NAND2_X1 U15092 ( .A1(n12589), .A2(n14034), .ZN(n12590) );
  INV_X1 U15093 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13197) );
  MUX2_X1 U15094 ( .A(n13199), .B(n13197), .S(n10481), .Z(n12608) );
  XNOR2_X1 U15095 ( .A(n12608), .B(SI_30_), .ZN(n12607) );
  NAND2_X1 U15096 ( .A1(n13195), .A2(n12614), .ZN(n12593) );
  OR2_X1 U15097 ( .A1(n12615), .A2(n13199), .ZN(n12592) );
  MUX2_X1 U15098 ( .A(n12594), .B(n15383), .S(n12600), .Z(n12606) );
  NAND2_X1 U15099 ( .A1(n15121), .A2(n6549), .ZN(n12599) );
  NAND2_X1 U15100 ( .A1(n15118), .A2(n12600), .ZN(n12595) );
  OAI21_X1 U15101 ( .B1(n9977), .B2(n12596), .A(n12595), .ZN(n12597) );
  NAND2_X1 U15102 ( .A1(n12597), .A2(n14933), .ZN(n12598) );
  NAND2_X1 U15103 ( .A1(n12599), .A2(n12598), .ZN(n12605) );
  INV_X1 U15104 ( .A(n14934), .ZN(n12601) );
  INV_X1 U15105 ( .A(n13032), .ZN(n15394) );
  MUX2_X1 U15106 ( .A(n12601), .B(n15394), .S(n12600), .Z(n12602) );
  INV_X1 U15107 ( .A(n12607), .ZN(n12610) );
  INV_X1 U15108 ( .A(n12608), .ZN(n12609) );
  MUX2_X1 U15109 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10481), .Z(n12612) );
  XNOR2_X1 U15110 ( .A(n12612), .B(SI_31_), .ZN(n12613) );
  NAND2_X1 U15111 ( .A1(n12735), .A2(n12614), .ZN(n12617) );
  INV_X1 U15112 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n15547) );
  OR2_X1 U15113 ( .A1(n12615), .A2(n15547), .ZN(n12616) );
  NAND2_X1 U15114 ( .A1(n12619), .A2(n12618), .ZN(n12621) );
  AND2_X1 U15115 ( .A1(n12621), .A2(n12620), .ZN(n12628) );
  INV_X1 U15116 ( .A(n12628), .ZN(n12623) );
  NAND2_X1 U15117 ( .A1(n11112), .A2(n12622), .ZN(n12630) );
  NAND2_X1 U15118 ( .A1(n12623), .A2(n12630), .ZN(n12661) );
  INV_X1 U15119 ( .A(n15118), .ZN(n12625) );
  MUX2_X1 U15120 ( .A(n15379), .B(n12625), .S(n12624), .Z(n12626) );
  OAI21_X1 U15121 ( .B1(n12627), .B2(n15118), .A(n12626), .ZN(n12654) );
  INV_X1 U15122 ( .A(n12630), .ZN(n12658) );
  XNOR2_X1 U15123 ( .A(n15135), .B(n13025), .ZN(n15129) );
  XNOR2_X1 U15124 ( .A(n14822), .B(n14938), .ZN(n15171) );
  XNOR2_X1 U15125 ( .A(n15223), .B(n14941), .ZN(n15214) );
  XNOR2_X1 U15126 ( .A(n15443), .B(n13060), .ZN(n15227) );
  INV_X1 U15127 ( .A(n15266), .ZN(n15264) );
  INV_X1 U15128 ( .A(n15282), .ZN(n12631) );
  NOR2_X1 U15129 ( .A1(n12631), .A2(n15341), .ZN(n12647) );
  NOR4_X1 U15130 ( .A1(n15708), .A2(n12634), .A3(n11170), .A4(n12633), .ZN(
        n12638) );
  NAND4_X1 U15131 ( .A1(n12638), .A2(n12637), .A3(n12636), .A4(n12635), .ZN(
        n12640) );
  NOR4_X1 U15132 ( .A1(n12640), .A2(n12639), .A3(n15675), .A4(n15694), .ZN(
        n12643) );
  NAND4_X1 U15133 ( .A1(n15334), .A2(n12643), .A3(n12642), .A4(n12641), .ZN(
        n12645) );
  XNOR2_X1 U15134 ( .A(n15491), .B(n14754), .ZN(n15370) );
  XNOR2_X1 U15135 ( .A(n15472), .B(n13052), .ZN(n13015) );
  NOR4_X1 U15136 ( .A1(n12645), .A2(n12644), .A3(n15370), .A4(n13015), .ZN(
        n12646) );
  XNOR2_X1 U15137 ( .A(n15303), .B(n14946), .ZN(n15296) );
  NAND4_X1 U15138 ( .A1(n15245), .A2(n12647), .A3(n12646), .A4(n15296), .ZN(
        n12648) );
  NOR4_X1 U15139 ( .A1(n15214), .A2(n15227), .A3(n15264), .A4(n12648), .ZN(
        n12649) );
  XNOR2_X1 U15140 ( .A(n15428), .B(n14940), .ZN(n15201) );
  XNOR2_X1 U15141 ( .A(n15425), .B(n14939), .ZN(n15185) );
  NAND4_X1 U15142 ( .A1(n15171), .A2(n12649), .A3(n15201), .A4(n15185), .ZN(
        n12650) );
  NOR4_X1 U15143 ( .A1(n15129), .A2(n15141), .A3(n15156), .A4(n12650), .ZN(
        n12652) );
  XNOR2_X1 U15144 ( .A(n15121), .B(n14933), .ZN(n12651) );
  NOR2_X1 U15145 ( .A1(n12654), .A2(n12661), .ZN(n12655) );
  AOI211_X1 U15146 ( .C1(n12658), .C2(n12657), .A(n12656), .B(n12655), .ZN(
        n12659) );
  OAI211_X1 U15147 ( .C1(n12662), .C2(n12661), .A(n12660), .B(n12659), .ZN(
        n12663) );
  INV_X1 U15148 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n12668) );
  OAI222_X1 U15149 ( .A1(n13196), .A2(n12668), .B1(n12667), .B2(n12666), .C1(
        P2_U3088), .C2(n12987), .ZN(P2_U3308) );
  NAND2_X1 U15150 ( .A1(n12669), .A2(n13579), .ZN(n12670) );
  XNOR2_X1 U15151 ( .A(n13356), .B(n13261), .ZN(n13348) );
  AND2_X1 U15152 ( .A1(n13348), .A2(n12672), .ZN(n12673) );
  XNOR2_X1 U15153 ( .A(n13476), .B(n13261), .ZN(n13289) );
  NAND2_X1 U15154 ( .A1(n13289), .A2(n13890), .ZN(n12674) );
  INV_X1 U15155 ( .A(n13289), .ZN(n12675) );
  NAND2_X1 U15156 ( .A1(n12675), .A2(n13475), .ZN(n12676) );
  XNOR2_X1 U15157 ( .A(n14017), .B(n12695), .ZN(n12677) );
  XNOR2_X1 U15158 ( .A(n12677), .B(n13865), .ZN(n13300) );
  INV_X1 U15159 ( .A(n12677), .ZN(n12678) );
  NAND2_X1 U15160 ( .A1(n12678), .A2(n13578), .ZN(n12679) );
  XNOR2_X1 U15161 ( .A(n13874), .B(n12695), .ZN(n12680) );
  XNOR2_X1 U15162 ( .A(n12680), .B(n13887), .ZN(n13327) );
  INV_X1 U15163 ( .A(n12680), .ZN(n12681) );
  NAND2_X1 U15164 ( .A1(n12681), .A2(n13887), .ZN(n12682) );
  XNOR2_X1 U15165 ( .A(n13853), .B(n12695), .ZN(n12683) );
  XNOR2_X1 U15166 ( .A(n12683), .B(n8429), .ZN(n13251) );
  INV_X1 U15167 ( .A(n12683), .ZN(n12684) );
  NAND2_X1 U15168 ( .A1(n12684), .A2(n13864), .ZN(n12685) );
  XNOR2_X1 U15169 ( .A(n13831), .B(n12695), .ZN(n12686) );
  XNOR2_X1 U15170 ( .A(n12686), .B(n13849), .ZN(n13309) );
  INV_X1 U15171 ( .A(n12686), .ZN(n12687) );
  NAND2_X1 U15172 ( .A1(n12687), .A2(n13252), .ZN(n12688) );
  XNOR2_X1 U15173 ( .A(n13923), .B(n13261), .ZN(n12689) );
  XNOR2_X1 U15174 ( .A(n12689), .B(n13836), .ZN(n13272) );
  INV_X1 U15175 ( .A(n12689), .ZN(n12690) );
  XNOR2_X1 U15176 ( .A(n13990), .B(n13261), .ZN(n13212) );
  NAND2_X1 U15177 ( .A1(n13317), .A2(n13826), .ZN(n12692) );
  INV_X1 U15178 ( .A(n13212), .ZN(n12691) );
  XNOR2_X1 U15179 ( .A(n13984), .B(n12695), .ZN(n13214) );
  XNOR2_X1 U15180 ( .A(n13912), .B(n12695), .ZN(n13211) );
  AOI22_X1 U15181 ( .A1(n13282), .A2(n13790), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12697) );
  NAND2_X1 U15182 ( .A1(n13354), .A2(n13795), .ZN(n12696) );
  OAI211_X1 U15183 ( .C1(n13497), .C2(n13352), .A(n12697), .B(n12696), .ZN(
        n12698) );
  AOI21_X1 U15184 ( .B1(n13912), .B2(n13357), .A(n12698), .ZN(n12699) );
  INV_X1 U15185 ( .A(n15957), .ZN(n15950) );
  XNOR2_X1 U15186 ( .A(n12700), .B(n13530), .ZN(n12749) );
  INV_X1 U15187 ( .A(n12749), .ZN(n12709) );
  XNOR2_X1 U15188 ( .A(n12701), .B(n13530), .ZN(n12702) );
  NAND2_X1 U15189 ( .A1(n12702), .A2(n13960), .ZN(n12706) );
  OAI22_X1 U15190 ( .A1(n13775), .A2(n15914), .B1(n15916), .B2(n12703), .ZN(
        n12704) );
  INV_X1 U15191 ( .A(n12704), .ZN(n12705) );
  OAI21_X1 U15192 ( .B1(n15950), .B2(n12709), .A(n12751), .ZN(n12712) );
  MUX2_X1 U15193 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n12712), .S(n15976), .Z(
        n12710) );
  INV_X1 U15194 ( .A(n12710), .ZN(n12711) );
  OAI21_X1 U15195 ( .B1(n12746), .B2(n13940), .A(n12711), .ZN(P3_U3486) );
  MUX2_X1 U15196 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n12712), .S(n15959), .Z(
        n12713) );
  INV_X1 U15197 ( .A(n12713), .ZN(n12714) );
  OAI21_X1 U15198 ( .B1(n12746), .B2(n14013), .A(n12714), .ZN(P3_U3454) );
  NOR2_X1 U15199 ( .A1(n12715), .A2(n14330), .ZN(n12720) );
  INV_X1 U15200 ( .A(n12716), .ZN(n12717) );
  AOI22_X1 U15201 ( .A1(n12717), .A2(n14560), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n14499), .ZN(n12718) );
  OAI21_X1 U15202 ( .B1(n12925), .B2(n14563), .A(n12718), .ZN(n12719) );
  AOI211_X1 U15203 ( .C1(n12721), .C2(n15850), .A(n12720), .B(n12719), .ZN(
        n12722) );
  OAI21_X1 U15204 ( .B1(n12723), .B2(n14546), .A(n12722), .ZN(P2_U3236) );
  XNOR2_X1 U15205 ( .A(n12725), .B(n12724), .ZN(n12726) );
  NAND2_X1 U15206 ( .A1(n12726), .A2(n14910), .ZN(n12730) );
  AOI22_X1 U15207 ( .A1(n12728), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n12727), 
        .B2(n15641), .ZN(n12729) );
  OAI211_X1 U15208 ( .C1(n15732), .C2(n14918), .A(n12730), .B(n12729), .ZN(
        P1_U3222) );
  NAND2_X1 U15209 ( .A1(n13195), .A2(n12734), .ZN(n12732) );
  OR2_X1 U15210 ( .A1(n8902), .A2(n13197), .ZN(n12731) );
  INV_X1 U15211 ( .A(n14570), .ZN(n12939) );
  XNOR2_X1 U15212 ( .A(n12753), .B(n12939), .ZN(n12736) );
  NAND2_X1 U15213 ( .A1(n12736), .A2(n10836), .ZN(n14569) );
  INV_X1 U15214 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n12742) );
  NAND2_X1 U15215 ( .A1(n12737), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n12740) );
  INV_X1 U15216 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n12738) );
  OR2_X1 U15217 ( .A1(n8891), .A2(n12738), .ZN(n12739) );
  OAI211_X1 U15218 ( .C1(n8931), .C2(n12742), .A(n12740), .B(n12739), .ZN(
        n14215) );
  NAND2_X1 U15219 ( .A1(n12741), .A2(n14215), .ZN(n14571) );
  NOR2_X1 U15220 ( .A1(n14499), .A2(n14571), .ZN(n12758) );
  NOR2_X1 U15221 ( .A1(n15850), .A2(n12742), .ZN(n12743) );
  AOI211_X1 U15222 ( .C1(n12939), .C2(n14541), .A(n12758), .B(n12743), .ZN(
        n12744) );
  OAI21_X1 U15223 ( .B1(n14569), .B2(n14330), .A(n12744), .ZN(P2_U3234) );
  AOI22_X1 U15224 ( .A1(n15903), .A2(P3_REG2_REG_27__SCAN_IN), .B1(n15901), 
        .B2(n13225), .ZN(n12745) );
  OAI21_X1 U15225 ( .B1(n12746), .B2(n13852), .A(n12745), .ZN(n12747) );
  AOI21_X1 U15226 ( .B1(n12749), .B2(n12748), .A(n12747), .ZN(n12750) );
  OAI21_X1 U15227 ( .B1(n12751), .B2(n15903), .A(n12750), .ZN(P3_U3206) );
  INV_X1 U15228 ( .A(n12752), .ZN(n12755) );
  INV_X1 U15229 ( .A(n12753), .ZN(n12754) );
  NOR2_X1 U15230 ( .A1(n15850), .A2(n12756), .ZN(n12757) );
  AOI211_X1 U15231 ( .C1(n12985), .C2(n14541), .A(n12758), .B(n12757), .ZN(
        n12759) );
  OAI21_X1 U15232 ( .B1(n14572), .B2(n14330), .A(n12759), .ZN(P2_U3235) );
  NAND3_X1 U15233 ( .A1(n9290), .A2(n14299), .A3(n12988), .ZN(n12760) );
  NAND2_X1 U15234 ( .A1(n12763), .A2(n15844), .ZN(n12932) );
  NAND2_X1 U15235 ( .A1(n12760), .A2(n12932), .ZN(n12955) );
  INV_X1 U15236 ( .A(n12761), .ZN(n12762) );
  OAI22_X1 U15237 ( .A1(n12762), .A2(n14299), .B1(n12767), .B2(n12763), .ZN(
        n12954) );
  INV_X1 U15238 ( .A(n14215), .ZN(n12938) );
  INV_X2 U15239 ( .A(n12777), .ZN(n12930) );
  NOR2_X1 U15240 ( .A1(n12938), .A2(n12930), .ZN(n12953) );
  MUX2_X1 U15241 ( .A(n7417), .B(n12765), .S(n12930), .Z(n12908) );
  INV_X1 U15242 ( .A(n12777), .ZN(n12774) );
  MUX2_X1 U15243 ( .A(n14236), .B(n14668), .S(n12774), .Z(n12814) );
  MUX2_X1 U15244 ( .A(n14238), .B(n14675), .S(n12774), .Z(n12805) );
  INV_X1 U15245 ( .A(n14243), .ZN(n12769) );
  NOR2_X1 U15246 ( .A1(n12987), .A2(n12763), .ZN(n12766) );
  OR2_X1 U15247 ( .A1(n12767), .A2(n12766), .ZN(n12771) );
  OAI21_X1 U15248 ( .B1(n12777), .B2(n12770), .A(n12771), .ZN(n12768) );
  NAND2_X1 U15249 ( .A1(n12769), .A2(n12768), .ZN(n12773) );
  NAND3_X1 U15250 ( .A1(n14243), .A2(n12777), .A3(n12770), .ZN(n12772) );
  NAND3_X1 U15251 ( .A1(n12773), .A2(n12772), .A3(n8096), .ZN(n12780) );
  MUX2_X1 U15252 ( .A(n6553), .B(n12775), .S(n12774), .Z(n12776) );
  INV_X1 U15253 ( .A(n12776), .ZN(n12781) );
  MUX2_X1 U15254 ( .A(n12775), .B(n6553), .S(n6541), .Z(n12779) );
  OAI21_X1 U15255 ( .B1(n12780), .B2(n12781), .A(n12779), .ZN(n12783) );
  NAND2_X1 U15256 ( .A1(n12781), .A2(n12780), .ZN(n12782) );
  NAND2_X1 U15257 ( .A1(n12783), .A2(n12782), .ZN(n12788) );
  MUX2_X1 U15258 ( .A(n14242), .B(n12784), .S(n6542), .Z(n12787) );
  NAND2_X1 U15259 ( .A1(n12788), .A2(n12787), .ZN(n12786) );
  MUX2_X1 U15260 ( .A(n12784), .B(n14242), .S(n6542), .Z(n12785) );
  NAND2_X1 U15261 ( .A1(n12786), .A2(n12785), .ZN(n12790) );
  OR2_X1 U15262 ( .A1(n12788), .A2(n12787), .ZN(n12789) );
  MUX2_X1 U15263 ( .A(n12791), .B(n14241), .S(n6542), .Z(n12793) );
  INV_X1 U15264 ( .A(n12793), .ZN(n12794) );
  MUX2_X1 U15265 ( .A(n14240), .B(n12795), .S(n6542), .Z(n12797) );
  MUX2_X1 U15266 ( .A(n12795), .B(n14240), .S(n6542), .Z(n12796) );
  INV_X1 U15267 ( .A(n12797), .ZN(n12798) );
  MUX2_X1 U15268 ( .A(n12799), .B(n14239), .S(n6542), .Z(n12802) );
  MUX2_X1 U15269 ( .A(n12800), .B(n15880), .S(n6542), .Z(n12801) );
  MUX2_X1 U15270 ( .A(n14675), .B(n14238), .S(n6542), .Z(n12804) );
  MUX2_X1 U15271 ( .A(n14237), .B(n12807), .S(n12777), .Z(n12811) );
  MUX2_X1 U15272 ( .A(n12809), .B(n12808), .S(n6542), .Z(n12810) );
  MUX2_X1 U15273 ( .A(n14236), .B(n14668), .S(n12777), .Z(n12812) );
  MUX2_X1 U15274 ( .A(n14092), .B(n12815), .S(n12777), .Z(n12833) );
  MUX2_X1 U15275 ( .A(n14233), .B(n14658), .S(n6542), .Z(n12832) );
  NAND2_X1 U15276 ( .A1(n12833), .A2(n12832), .ZN(n12837) );
  MUX2_X1 U15277 ( .A(n12817), .B(n12816), .S(n12777), .Z(n12829) );
  INV_X1 U15278 ( .A(n12817), .ZN(n14234) );
  MUX2_X1 U15279 ( .A(n14234), .B(n12818), .S(n6542), .Z(n12828) );
  NAND2_X1 U15280 ( .A1(n12829), .A2(n12828), .ZN(n12819) );
  AND2_X1 U15281 ( .A1(n12837), .A2(n12819), .ZN(n12824) );
  MUX2_X1 U15282 ( .A(n12820), .B(n7859), .S(n12777), .Z(n12826) );
  MUX2_X1 U15283 ( .A(n14235), .B(n14663), .S(n6542), .Z(n12825) );
  NAND2_X1 U15284 ( .A1(n12826), .A2(n12825), .ZN(n12822) );
  AND2_X1 U15285 ( .A1(n12824), .A2(n12822), .ZN(n12823) );
  INV_X1 U15286 ( .A(n12824), .ZN(n12827) );
  MUX2_X1 U15287 ( .A(n14152), .B(n7108), .S(n12930), .Z(n12854) );
  MUX2_X1 U15288 ( .A(n7107), .B(n14653), .S(n12777), .Z(n12853) );
  NAND2_X1 U15289 ( .A1(n12854), .A2(n12853), .ZN(n12839) );
  INV_X1 U15290 ( .A(n12828), .ZN(n12831) );
  INV_X1 U15291 ( .A(n12829), .ZN(n12830) );
  AND2_X1 U15292 ( .A1(n12831), .A2(n12830), .ZN(n12836) );
  INV_X1 U15293 ( .A(n12832), .ZN(n12835) );
  INV_X1 U15294 ( .A(n12833), .ZN(n12834) );
  AOI22_X1 U15295 ( .A1(n12837), .A2(n12836), .B1(n12835), .B2(n12834), .ZN(
        n12838) );
  NAND2_X1 U15296 ( .A1(n12842), .A2(n12841), .ZN(n12858) );
  INV_X1 U15297 ( .A(n14116), .ZN(n14231) );
  OR2_X1 U15298 ( .A1(n14500), .A2(n12777), .ZN(n12844) );
  NAND2_X1 U15299 ( .A1(n14116), .A2(n12777), .ZN(n12843) );
  NAND2_X1 U15300 ( .A1(n12844), .A2(n12843), .ZN(n12865) );
  OR2_X1 U15301 ( .A1(n12866), .A2(n12865), .ZN(n12849) );
  NOR2_X1 U15302 ( .A1(n14205), .A2(n12930), .ZN(n12847) );
  NAND2_X1 U15303 ( .A1(n14205), .A2(n12930), .ZN(n12845) );
  NAND2_X1 U15304 ( .A1(n14631), .A2(n12845), .ZN(n12846) );
  OAI21_X1 U15305 ( .B1(n14631), .B2(n12847), .A(n12846), .ZN(n12848) );
  AND3_X1 U15306 ( .A1(n12848), .A2(n12864), .A3(n14473), .ZN(n12867) );
  AND2_X1 U15307 ( .A1(n12849), .A2(n12867), .ZN(n12859) );
  MUX2_X1 U15308 ( .A(n14232), .B(n14643), .S(n12930), .Z(n12860) );
  NAND2_X1 U15309 ( .A1(n12861), .A2(n12860), .ZN(n12851) );
  AND2_X1 U15310 ( .A1(n12859), .A2(n12851), .ZN(n12879) );
  MUX2_X1 U15311 ( .A(n14091), .B(n12852), .S(n12777), .Z(n12876) );
  MUX2_X1 U15312 ( .A(n9355), .B(n14648), .S(n12930), .Z(n12875) );
  INV_X1 U15313 ( .A(n12853), .ZN(n12856) );
  INV_X1 U15314 ( .A(n12854), .ZN(n12855) );
  AOI22_X1 U15315 ( .A1(n12876), .A2(n12875), .B1(n12856), .B2(n12855), .ZN(
        n12857) );
  NAND3_X1 U15316 ( .A1(n12858), .A2(n12879), .A3(n12857), .ZN(n12883) );
  INV_X1 U15317 ( .A(n12859), .ZN(n12873) );
  INV_X1 U15318 ( .A(n12860), .ZN(n12863) );
  INV_X1 U15319 ( .A(n12861), .ZN(n12862) );
  NAND2_X1 U15320 ( .A1(n12863), .A2(n12862), .ZN(n12872) );
  MUX2_X1 U15321 ( .A(n12864), .B(n14473), .S(n12930), .Z(n12871) );
  AOI21_X1 U15322 ( .B1(n12866), .B2(n12865), .A(n14488), .ZN(n12869) );
  INV_X1 U15323 ( .A(n12867), .ZN(n12868) );
  OAI211_X1 U15324 ( .C1(n12873), .C2(n12872), .A(n12871), .B(n12870), .ZN(
        n12874) );
  INV_X1 U15325 ( .A(n12874), .ZN(n12881) );
  INV_X1 U15326 ( .A(n12875), .ZN(n12878) );
  INV_X1 U15327 ( .A(n12876), .ZN(n12877) );
  NAND3_X1 U15328 ( .A1(n12879), .A2(n12878), .A3(n12877), .ZN(n12880) );
  MUX2_X1 U15329 ( .A(n12884), .B(n9360), .S(n12930), .Z(n12886) );
  MUX2_X1 U15330 ( .A(n14228), .B(n14620), .S(n12777), .Z(n12885) );
  MUX2_X1 U15331 ( .A(n14227), .B(n14615), .S(n12777), .Z(n12889) );
  MUX2_X1 U15332 ( .A(n14227), .B(n14615), .S(n12930), .Z(n12887) );
  NAND2_X1 U15333 ( .A1(n12888), .A2(n12887), .ZN(n12890) );
  MUX2_X1 U15334 ( .A(n14226), .B(n14610), .S(n12930), .Z(n12893) );
  MUX2_X1 U15335 ( .A(n14226), .B(n14610), .S(n12777), .Z(n12891) );
  MUX2_X1 U15336 ( .A(n14225), .B(n14605), .S(n12777), .Z(n12896) );
  MUX2_X1 U15337 ( .A(n14225), .B(n14605), .S(n12930), .Z(n12895) );
  NAND2_X1 U15338 ( .A1(n12898), .A2(n12897), .ZN(n12900) );
  MUX2_X1 U15339 ( .A(n14224), .B(n14600), .S(n12930), .Z(n12901) );
  MUX2_X1 U15340 ( .A(n14600), .B(n14224), .S(n12930), .Z(n12899) );
  INV_X1 U15341 ( .A(n12901), .ZN(n12902) );
  MUX2_X1 U15342 ( .A(n14223), .B(n14595), .S(n12777), .Z(n12905) );
  MUX2_X1 U15343 ( .A(n14223), .B(n14595), .S(n12930), .Z(n12903) );
  INV_X1 U15344 ( .A(n12905), .ZN(n12906) );
  MUX2_X1 U15345 ( .A(n14590), .B(n14222), .S(n12930), .Z(n12907) );
  MUX2_X1 U15346 ( .A(n14585), .B(n14221), .S(n12930), .Z(n12911) );
  MUX2_X1 U15347 ( .A(n14101), .B(n14582), .S(n12930), .Z(n12915) );
  INV_X1 U15348 ( .A(n14101), .ZN(n14220) );
  MUX2_X1 U15349 ( .A(n14220), .B(n14327), .S(n12777), .Z(n12914) );
  OAI22_X1 U15350 ( .A1(n12912), .A2(n12911), .B1(n12915), .B2(n12914), .ZN(
        n12918) );
  MUX2_X1 U15351 ( .A(n12909), .B(n14346), .S(n12930), .Z(n12910) );
  AOI21_X1 U15352 ( .B1(n12912), .B2(n12911), .A(n12910), .ZN(n12917) );
  INV_X1 U15353 ( .A(n14219), .ZN(n12913) );
  MUX2_X1 U15354 ( .A(n12913), .B(n14307), .S(n12930), .Z(n12921) );
  MUX2_X1 U15355 ( .A(n14219), .B(n14576), .S(n12777), .Z(n12920) );
  AOI22_X1 U15356 ( .A1(n12921), .A2(n12920), .B1(n12915), .B2(n12914), .ZN(
        n12916) );
  OAI21_X1 U15357 ( .B1(n12918), .B2(n12917), .A(n12916), .ZN(n12929) );
  INV_X1 U15358 ( .A(n14218), .ZN(n13204) );
  MUX2_X1 U15359 ( .A(n13204), .B(n12919), .S(n12777), .Z(n12944) );
  MUX2_X1 U15360 ( .A(n14218), .B(n13180), .S(n12930), .Z(n12943) );
  INV_X1 U15361 ( .A(n12920), .ZN(n12923) );
  INV_X1 U15362 ( .A(n12921), .ZN(n12922) );
  AOI22_X1 U15363 ( .A1(n12944), .A2(n12943), .B1(n12923), .B2(n12922), .ZN(
        n12927) );
  MUX2_X1 U15364 ( .A(n12925), .B(n12924), .S(n12930), .Z(n12937) );
  MUX2_X1 U15365 ( .A(n14217), .B(n12926), .S(n12930), .Z(n12936) );
  NAND2_X1 U15366 ( .A1(n12937), .A2(n12936), .ZN(n12942) );
  MUX2_X1 U15367 ( .A(n14216), .B(n12985), .S(n12930), .Z(n12951) );
  NAND2_X1 U15368 ( .A1(n14215), .A2(n12930), .ZN(n12933) );
  NAND4_X1 U15369 ( .A1(n12933), .A2(n12988), .A3(n12932), .A4(n12931), .ZN(
        n12934) );
  AND2_X1 U15370 ( .A1(n12934), .A2(n14216), .ZN(n12935) );
  AOI21_X1 U15371 ( .B1(n12985), .B2(n12777), .A(n12935), .ZN(n12950) );
  OAI22_X1 U15372 ( .A1(n12951), .A2(n12950), .B1(n12937), .B2(n12936), .ZN(
        n12949) );
  NAND2_X1 U15373 ( .A1(n12939), .A2(n12938), .ZN(n12941) );
  NAND2_X1 U15374 ( .A1(n14570), .A2(n14215), .ZN(n12940) );
  MUX2_X1 U15375 ( .A(n12941), .B(n12940), .S(n12930), .Z(n12948) );
  INV_X1 U15376 ( .A(n12986), .ZN(n12946) );
  INV_X1 U15377 ( .A(n12942), .ZN(n12945) );
  NOR4_X1 U15378 ( .A1(n12946), .A2(n12945), .A3(n12944), .A4(n12943), .ZN(
        n12947) );
  AOI21_X1 U15379 ( .B1(n12949), .B2(n12948), .A(n12947), .ZN(n12952) );
  XNOR2_X1 U15380 ( .A(n14643), .B(n14203), .ZN(n14516) );
  INV_X1 U15381 ( .A(n14488), .ZN(n12976) );
  INV_X1 U15382 ( .A(n15848), .ZN(n12962) );
  NAND4_X1 U15383 ( .A1(n12961), .A2(n9290), .A3(n12962), .A4(n12960), .ZN(
        n12966) );
  NAND4_X1 U15384 ( .A1(n12970), .A2(n12969), .A3(n12968), .A4(n12967), .ZN(
        n12972) );
  NOR2_X1 U15385 ( .A1(n12972), .A2(n12971), .ZN(n12974) );
  XNOR2_X1 U15386 ( .A(n14653), .B(n7107), .ZN(n14550) );
  NAND2_X1 U15387 ( .A1(n12978), .A2(n12977), .ZN(n14439) );
  NAND4_X1 U15388 ( .A1(n12979), .A2(n6715), .A3(n14424), .A4(n14439), .ZN(
        n12980) );
  NOR4_X1 U15389 ( .A1(n14354), .A2(n14411), .A3(n14379), .A4(n12980), .ZN(
        n12981) );
  NAND3_X1 U15390 ( .A1(n14319), .A2(n12981), .A3(n14337), .ZN(n12982) );
  NAND3_X1 U15391 ( .A1(n12990), .A2(n14192), .A3(n12989), .ZN(n12991) );
  OAI211_X1 U15392 ( .C1(n12763), .C2(n12993), .A(n12991), .B(P2_B_REG_SCAN_IN), .ZN(n12992) );
  INV_X1 U15393 ( .A(n12994), .ZN(n12995) );
  NAND2_X1 U15394 ( .A1(n12995), .A2(n14461), .ZN(n13001) );
  INV_X1 U15395 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n12996) );
  OAI22_X1 U15396 ( .A1(n13173), .A2(n15843), .B1(n12996), .B2(n15850), .ZN(
        n12999) );
  NOR2_X1 U15397 ( .A1(n12997), .A2(n14330), .ZN(n12998) );
  AOI211_X1 U15398 ( .C1(n14541), .C2(n13180), .A(n12999), .B(n12998), .ZN(
        n13000) );
  OAI211_X1 U15399 ( .C1(n14499), .C2(n6738), .A(n13001), .B(n13000), .ZN(
        P2_U3237) );
  INV_X1 U15400 ( .A(n13002), .ZN(n13193) );
  OAI222_X1 U15401 ( .A1(n9426), .A2(P1_U3086), .B1(n10985), .B2(n13193), .C1(
        n13003), .C2(n15546), .ZN(P1_U3326) );
  INV_X1 U15402 ( .A(SI_30_), .ZN(n13374) );
  NAND2_X1 U15403 ( .A1(n13003), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13004) );
  NAND2_X1 U15404 ( .A1(n13005), .A2(n13004), .ZN(n13008) );
  NAND2_X1 U15405 ( .A1(n13199), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13364) );
  NAND2_X1 U15406 ( .A1(n13197), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13006) );
  AND2_X1 U15407 ( .A1(n13364), .A2(n13006), .ZN(n13007) );
  NAND2_X1 U15408 ( .A1(n13008), .A2(n13007), .ZN(n13365) );
  OAI222_X1 U15409 ( .A1(n8121), .A2(P3_U3151), .B1(n14033), .B2(n13374), .C1(
        n14040), .C2(n13373), .ZN(P3_U3265) );
  NAND2_X1 U15410 ( .A1(n7298), .A2(n14873), .ZN(n13009) );
  AND2_X1 U15411 ( .A1(n15486), .A2(n14948), .ZN(n15328) );
  AND2_X1 U15412 ( .A1(n15368), .A2(n14754), .ZN(n15317) );
  INV_X1 U15413 ( .A(n13014), .ZN(n15319) );
  AOI21_X1 U15414 ( .B1(n15319), .B2(n15320), .A(n15318), .ZN(n13016) );
  OR2_X1 U15415 ( .A1(n15472), .A2(n14947), .ZN(n13018) );
  OR2_X1 U15416 ( .A1(n15466), .A2(n14831), .ZN(n13019) );
  NAND2_X1 U15417 ( .A1(n15466), .A2(n14831), .ZN(n13020) );
  NOR2_X1 U15418 ( .A1(n15461), .A2(n14945), .ZN(n13021) );
  INV_X1 U15419 ( .A(n15227), .ZN(n15234) );
  OR2_X1 U15420 ( .A1(n15437), .A2(n14941), .ZN(n13022) );
  INV_X1 U15421 ( .A(n15201), .ZN(n13023) );
  NAND2_X1 U15422 ( .A1(n15428), .A2(n14940), .ZN(n13024) );
  OR2_X1 U15423 ( .A1(n15400), .A2(n13025), .ZN(n13028) );
  INV_X1 U15424 ( .A(n13028), .ZN(n13026) );
  NOR2_X1 U15425 ( .A1(n15387), .A2(n13026), .ZN(n13031) );
  NOR2_X1 U15426 ( .A1(n15150), .A2(n14936), .ZN(n15128) );
  NOR2_X1 U15427 ( .A1(n15135), .A2(n14935), .ZN(n13029) );
  AOI211_X1 U15428 ( .C1(n15128), .C2(n13028), .A(n13029), .B(n15387), .ZN(
        n13027) );
  AOI21_X1 U15429 ( .B1(n15387), .B2(n13028), .A(n13027), .ZN(n13030) );
  INV_X1 U15430 ( .A(n15472), .ZN(n15307) );
  NAND2_X1 U15431 ( .A1(n15299), .A2(n15466), .ZN(n15298) );
  AND2_X2 U15432 ( .A1(n15191), .A2(n15417), .ZN(n15172) );
  AND2_X2 U15433 ( .A1(n15172), .A2(n15410), .ZN(n15159) );
  AOI211_X1 U15434 ( .C1(n13032), .C2(n15130), .A(n15733), .B(n15122), .ZN(
        n15396) );
  NAND2_X1 U15435 ( .A1(n14935), .A2(n15637), .ZN(n15392) );
  NAND2_X1 U15436 ( .A1(n13032), .A2(n15716), .ZN(n13040) );
  INV_X1 U15437 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n13036) );
  NOR2_X1 U15438 ( .A1(n7374), .A2(n13033), .ZN(n13034) );
  NOR2_X1 U15439 ( .A1(n14913), .A2(n13034), .ZN(n15117) );
  NAND2_X1 U15440 ( .A1(n14933), .A2(n15117), .ZN(n15393) );
  OAI22_X1 U15441 ( .A1(n15714), .A2(n13036), .B1(n15393), .B2(n13035), .ZN(
        n13037) );
  AOI21_X1 U15442 ( .B1(n13038), .B2(n15698), .A(n13037), .ZN(n13039) );
  OAI211_X1 U15443 ( .C1(n6546), .C2(n15392), .A(n13040), .B(n13039), .ZN(
        n13041) );
  AOI21_X1 U15444 ( .B1(n15396), .B2(n15720), .A(n13041), .ZN(n13074) );
  NAND2_X1 U15445 ( .A1(n7298), .A2(n14950), .ZN(n13042) );
  NAND2_X1 U15446 ( .A1(n13043), .A2(n13042), .ZN(n15339) );
  AND2_X1 U15447 ( .A1(n15368), .A2(n14949), .ZN(n15340) );
  NAND2_X1 U15448 ( .A1(n13047), .A2(n15340), .ZN(n13049) );
  AND2_X1 U15449 ( .A1(n13049), .A2(n13048), .ZN(n13050) );
  NAND2_X1 U15450 ( .A1(n15472), .A2(n13052), .ZN(n15293) );
  OAI21_X1 U15451 ( .B1(n15455), .B2(n13055), .A(n15244), .ZN(n13053) );
  INV_X1 U15452 ( .A(n13053), .ZN(n13054) );
  NAND2_X1 U15453 ( .A1(n15281), .A2(n13054), .ZN(n13057) );
  NAND2_X1 U15454 ( .A1(n15455), .A2(n13055), .ZN(n15246) );
  AND2_X1 U15455 ( .A1(n15245), .A2(n15246), .ZN(n13056) );
  OR2_X1 U15456 ( .A1(n15447), .A2(n13058), .ZN(n13059) );
  OR2_X1 U15457 ( .A1(n15443), .A2(n13060), .ZN(n13061) );
  NAND2_X1 U15458 ( .A1(n15437), .A2(n13063), .ZN(n13064) );
  INV_X1 U15459 ( .A(n14940), .ZN(n13065) );
  INV_X1 U15460 ( .A(n15185), .ZN(n15182) );
  INV_X1 U15461 ( .A(n14939), .ZN(n13066) );
  OR2_X1 U15462 ( .A1(n15425), .A2(n13066), .ZN(n13067) );
  INV_X1 U15463 ( .A(n15171), .ZN(n15169) );
  NAND2_X1 U15464 ( .A1(n14822), .A2(n14912), .ZN(n13068) );
  OR2_X1 U15465 ( .A1(n15163), .A2(n13069), .ZN(n13070) );
  AND2_X1 U15466 ( .A1(n15400), .A2(n14935), .ZN(n15388) );
  OR2_X1 U15467 ( .A1(n15400), .A2(n14935), .ZN(n15384) );
  OAI21_X1 U15468 ( .B1(n15389), .B2(n15388), .A(n15384), .ZN(n13071) );
  XNOR2_X1 U15469 ( .A(n13071), .B(n15387), .ZN(n13072) );
  NAND2_X1 U15470 ( .A1(n13072), .A2(n15295), .ZN(n13073) );
  OAI211_X1 U15471 ( .C1(n15397), .C2(n15374), .A(n13074), .B(n13073), .ZN(
        P1_U3356) );
  MUX2_X1 U15472 ( .A(P3_REG0_REG_28__SCAN_IN), .B(n13188), .S(n15959), .Z(
        n13077) );
  OAI22_X1 U15473 ( .A1(n13192), .A2(n14021), .B1(n13075), .B2(n14013), .ZN(
        n13076) );
  OR2_X1 U15474 ( .A1(n13077), .A2(n13076), .ZN(P3_U3455) );
  NAND3_X1 U15475 ( .A1(n13078), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n13083) );
  NAND2_X1 U15476 ( .A1(n12735), .A2(n13079), .ZN(n13082) );
  NAND2_X1 U15477 ( .A1(n13080), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n13081) );
  OAI211_X1 U15478 ( .C1(n13084), .C2(n13083), .A(n13082), .B(n13081), .ZN(
        P2_U3296) );
  NAND2_X1 U15479 ( .A1(n14218), .A2(n14508), .ZN(n13085) );
  XNOR2_X1 U15480 ( .A(n13085), .B(n13166), .ZN(n13086) );
  XNOR2_X1 U15481 ( .A(n13180), .B(n13086), .ZN(n13172) );
  INV_X1 U15482 ( .A(n13172), .ZN(n13087) );
  NAND2_X1 U15483 ( .A1(n13087), .A2(n14161), .ZN(n13183) );
  XNOR2_X1 U15484 ( .A(n14327), .B(n13166), .ZN(n13163) );
  INV_X1 U15485 ( .A(n13163), .ZN(n13165) );
  NOR2_X1 U15486 ( .A1(n14101), .A2(n13148), .ZN(n13162) );
  INV_X1 U15487 ( .A(n13162), .ZN(n13164) );
  XNOR2_X1 U15488 ( .A(n14600), .B(n13166), .ZN(n13149) );
  XNOR2_X1 U15489 ( .A(n14658), .B(n13166), .ZN(n13094) );
  NAND2_X1 U15490 ( .A1(n14508), .A2(n14233), .ZN(n13092) );
  XNOR2_X1 U15491 ( .A(n13094), .B(n13092), .ZN(n14172) );
  INV_X1 U15492 ( .A(n13092), .ZN(n13093) );
  NAND2_X1 U15493 ( .A1(n13094), .A2(n13093), .ZN(n13095) );
  NAND2_X1 U15494 ( .A1(n13096), .A2(n13095), .ZN(n14089) );
  XNOR2_X1 U15495 ( .A(n14653), .B(n7818), .ZN(n13097) );
  OR2_X1 U15496 ( .A1(n14152), .A2(n13148), .ZN(n13098) );
  NAND2_X1 U15497 ( .A1(n13097), .A2(n13098), .ZN(n13103) );
  INV_X1 U15498 ( .A(n13097), .ZN(n13100) );
  INV_X1 U15499 ( .A(n13098), .ZN(n13099) );
  NAND2_X1 U15500 ( .A1(n13100), .A2(n13099), .ZN(n13101) );
  NAND2_X1 U15501 ( .A1(n13103), .A2(n13101), .ZN(n14090) );
  INV_X1 U15502 ( .A(n14090), .ZN(n13102) );
  XNOR2_X1 U15503 ( .A(n14648), .B(n13166), .ZN(n13105) );
  NOR2_X1 U15504 ( .A1(n14091), .A2(n13148), .ZN(n13104) );
  XNOR2_X1 U15505 ( .A(n13105), .B(n13104), .ZN(n14150) );
  XNOR2_X1 U15506 ( .A(n14500), .B(n7818), .ZN(n14109) );
  NAND2_X1 U15507 ( .A1(n14231), .A2(n14508), .ZN(n13111) );
  NAND2_X1 U15508 ( .A1(n14109), .A2(n13111), .ZN(n13106) );
  XNOR2_X1 U15509 ( .A(n14631), .B(n7818), .ZN(n13112) );
  OR2_X1 U15510 ( .A1(n14205), .A2(n13148), .ZN(n13113) );
  NAND2_X1 U15511 ( .A1(n13112), .A2(n13113), .ZN(n14113) );
  NAND2_X1 U15512 ( .A1(n13106), .A2(n14113), .ZN(n13117) );
  XNOR2_X1 U15513 ( .A(n14643), .B(n13166), .ZN(n13110) );
  INV_X1 U15514 ( .A(n13110), .ZN(n13108) );
  NOR2_X1 U15515 ( .A1(n14203), .A2(n13148), .ZN(n13109) );
  INV_X1 U15516 ( .A(n13109), .ZN(n13107) );
  NOR2_X1 U15517 ( .A1(n13117), .A2(n14107), .ZN(n13119) );
  NAND2_X1 U15518 ( .A1(n13110), .A2(n13109), .ZN(n14043) );
  INV_X1 U15519 ( .A(n14109), .ZN(n14110) );
  INV_X1 U15520 ( .A(n13111), .ZN(n14200) );
  NAND3_X1 U15521 ( .A1(n14110), .A2(n14200), .A3(n14113), .ZN(n13116) );
  INV_X1 U15522 ( .A(n13112), .ZN(n13115) );
  INV_X1 U15523 ( .A(n13113), .ZN(n13114) );
  NAND2_X1 U15524 ( .A1(n13115), .A2(n13114), .ZN(n14112) );
  OAI211_X1 U15525 ( .C1(n13117), .C2(n14043), .A(n13116), .B(n14112), .ZN(
        n13118) );
  XNOR2_X1 U15526 ( .A(n14626), .B(n7818), .ZN(n13120) );
  OR2_X1 U15527 ( .A1(n14183), .A2(n13148), .ZN(n13121) );
  NAND2_X1 U15528 ( .A1(n13120), .A2(n13121), .ZN(n13125) );
  INV_X1 U15529 ( .A(n13120), .ZN(n13123) );
  INV_X1 U15530 ( .A(n13121), .ZN(n13122) );
  NAND2_X1 U15531 ( .A1(n13123), .A2(n13122), .ZN(n13124) );
  AND2_X1 U15532 ( .A1(n13125), .A2(n13124), .ZN(n14123) );
  XNOR2_X1 U15533 ( .A(n14620), .B(n7818), .ZN(n13126) );
  NAND2_X1 U15534 ( .A1(n14228), .A2(n14508), .ZN(n13127) );
  XNOR2_X1 U15535 ( .A(n13126), .B(n13127), .ZN(n14181) );
  XNOR2_X1 U15536 ( .A(n14615), .B(n7818), .ZN(n13130) );
  NAND2_X1 U15537 ( .A1(n14227), .A2(n14508), .ZN(n13131) );
  NAND2_X1 U15538 ( .A1(n13130), .A2(n13131), .ZN(n14065) );
  INV_X1 U15539 ( .A(n14065), .ZN(n13135) );
  XNOR2_X1 U15540 ( .A(n14610), .B(n7818), .ZN(n13137) );
  NAND2_X1 U15541 ( .A1(n14226), .A2(n14508), .ZN(n13136) );
  AND2_X1 U15542 ( .A1(n13137), .A2(n13136), .ZN(n13139) );
  OR2_X1 U15543 ( .A1(n14138), .A2(n13139), .ZN(n14075) );
  XNOR2_X1 U15544 ( .A(n14605), .B(n7818), .ZN(n13143) );
  NOR2_X1 U15545 ( .A1(n14165), .A2(n13148), .ZN(n13144) );
  XNOR2_X1 U15546 ( .A(n13143), .B(n13144), .ZN(n14079) );
  INV_X1 U15547 ( .A(n14079), .ZN(n13140) );
  INV_X1 U15548 ( .A(n13126), .ZN(n13129) );
  INV_X1 U15549 ( .A(n13127), .ZN(n13128) );
  NAND2_X1 U15550 ( .A1(n13129), .A2(n13128), .ZN(n14066) );
  INV_X1 U15551 ( .A(n13130), .ZN(n13133) );
  INV_X1 U15552 ( .A(n13131), .ZN(n13132) );
  NAND2_X1 U15553 ( .A1(n13133), .A2(n13132), .ZN(n14064) );
  XNOR2_X1 U15554 ( .A(n13137), .B(n13136), .ZN(n14144) );
  INV_X1 U15555 ( .A(n14144), .ZN(n13138) );
  INV_X1 U15556 ( .A(n13143), .ZN(n13145) );
  NAND2_X1 U15557 ( .A1(n13145), .A2(n13144), .ZN(n13146) );
  NOR2_X1 U15558 ( .A1(n14059), .A2(n13148), .ZN(n14163) );
  XNOR2_X1 U15559 ( .A(n14595), .B(n13166), .ZN(n13151) );
  NOR2_X1 U15560 ( .A1(n14166), .A2(n13148), .ZN(n13152) );
  OAI21_X1 U15561 ( .B1(n13152), .B2(n13151), .A(n14053), .ZN(n13153) );
  INV_X1 U15562 ( .A(n13151), .ZN(n14054) );
  INV_X1 U15563 ( .A(n13152), .ZN(n14058) );
  XNOR2_X1 U15564 ( .A(n14590), .B(n7818), .ZN(n13155) );
  NAND2_X1 U15565 ( .A1(n14222), .A2(n14508), .ZN(n13154) );
  NOR2_X1 U15566 ( .A1(n13155), .A2(n13154), .ZN(n13156) );
  AOI21_X1 U15567 ( .B1(n13155), .B2(n13154), .A(n13156), .ZN(n14131) );
  NAND2_X1 U15568 ( .A1(n14132), .A2(n14131), .ZN(n14130) );
  INV_X1 U15569 ( .A(n13156), .ZN(n13157) );
  XNOR2_X1 U15570 ( .A(n14585), .B(n7818), .ZN(n13159) );
  NAND2_X1 U15571 ( .A1(n14221), .A2(n14508), .ZN(n13158) );
  NOR2_X1 U15572 ( .A1(n13159), .A2(n13158), .ZN(n13160) );
  AOI21_X1 U15573 ( .B1(n13159), .B2(n13158), .A(n13160), .ZN(n14099) );
  INV_X1 U15574 ( .A(n13160), .ZN(n13161) );
  XNOR2_X1 U15575 ( .A(n13163), .B(n13162), .ZN(n14191) );
  XNOR2_X1 U15576 ( .A(n14576), .B(n13166), .ZN(n13168) );
  INV_X1 U15577 ( .A(n13168), .ZN(n13170) );
  AND2_X1 U15578 ( .A1(n14219), .A2(n14508), .ZN(n13167) );
  INV_X1 U15579 ( .A(n13167), .ZN(n13169) );
  AOI21_X1 U15580 ( .B1(n13170), .B2(n13169), .A(n13171), .ZN(n13202) );
  INV_X1 U15581 ( .A(n13171), .ZN(n13177) );
  INV_X1 U15582 ( .A(n13173), .ZN(n13174) );
  AOI22_X1 U15583 ( .A1(n13174), .A2(n14194), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13175) );
  OAI21_X1 U15584 ( .B1(n13176), .B2(n14196), .A(n13175), .ZN(n13179) );
  NOR2_X1 U15585 ( .A1(n13183), .A2(n13177), .ZN(n13178) );
  AOI211_X1 U15586 ( .C1(n13180), .C2(n14211), .A(n13179), .B(n13178), .ZN(
        n13181) );
  OAI211_X1 U15587 ( .C1(n13183), .C2(n13201), .A(n13182), .B(n13181), .ZN(
        P2_U3192) );
  INV_X1 U15588 ( .A(n13184), .ZN(n13186) );
  OAI222_X1 U15589 ( .A1(n13187), .A2(P1_U3086), .B1(n10985), .B2(n13186), 
        .C1(n13185), .C2(n15546), .ZN(P1_U3327) );
  MUX2_X1 U15590 ( .A(P3_REG2_REG_28__SCAN_IN), .B(n13188), .S(n15921), .Z(
        n13189) );
  INV_X1 U15591 ( .A(n13189), .ZN(n13191) );
  AOI22_X1 U15592 ( .A1(n13269), .A2(n13880), .B1(n15901), .B2(n13264), .ZN(
        n13190) );
  OAI211_X1 U15593 ( .C1(n13192), .C2(n13894), .A(n13191), .B(n13190), .ZN(
        P3_U3205) );
  OAI222_X1 U15594 ( .A1(n13196), .A2(n13194), .B1(n13198), .B2(n13193), .C1(
        P2_U3088), .C2(n6985), .ZN(P2_U3298) );
  INV_X1 U15595 ( .A(n13195), .ZN(n13200) );
  OAI222_X1 U15596 ( .A1(n13198), .A2(n13200), .B1(P2_U3088), .B2(n8798), .C1(
        n13197), .C2(n13196), .ZN(P2_U3297) );
  OAI222_X1 U15597 ( .A1(n10985), .A2(n13200), .B1(n9427), .B2(P1_U3086), .C1(
        n13199), .C2(n15546), .ZN(P1_U3325) );
  OAI211_X1 U15598 ( .C1(n13203), .C2(n13202), .A(n13201), .B(n14161), .ZN(
        n13208) );
  OAI22_X1 U15599 ( .A1(n13204), .A2(n14204), .B1(n14101), .B2(n14202), .ZN(
        n14305) );
  OAI22_X1 U15600 ( .A1(n14311), .A2(n14209), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13205), .ZN(n13206) );
  AOI21_X1 U15601 ( .B1(n14305), .B2(n14206), .A(n13206), .ZN(n13207) );
  XNOR2_X1 U15602 ( .A(n13229), .B(n13261), .ZN(n13258) );
  XNOR2_X1 U15603 ( .A(n13258), .B(n13768), .ZN(n13259) );
  OR2_X1 U15604 ( .A1(n13211), .A2(n13776), .ZN(n13210) );
  OR2_X1 U15605 ( .A1(n13214), .A2(n13497), .ZN(n13209) );
  NAND2_X1 U15606 ( .A1(n13210), .A2(n13209), .ZN(n13213) );
  AOI21_X1 U15607 ( .B1(n13212), .B2(n13805), .A(n13213), .ZN(n13220) );
  INV_X1 U15608 ( .A(n13211), .ZN(n13218) );
  AOI21_X1 U15609 ( .B1(n13214), .B2(n13497), .A(n13776), .ZN(n13217) );
  OR3_X1 U15610 ( .A1(n13213), .A2(n13212), .A3(n13805), .ZN(n13216) );
  NAND3_X1 U15611 ( .A1(n13214), .A2(n13497), .A3(n13776), .ZN(n13215) );
  OAI211_X1 U15612 ( .C1(n13218), .C2(n13217), .A(n13216), .B(n13215), .ZN(
        n13219) );
  XNOR2_X1 U15613 ( .A(n13908), .B(n13261), .ZN(n13222) );
  XNOR2_X1 U15614 ( .A(n13222), .B(n13790), .ZN(n13281) );
  XNOR2_X1 U15615 ( .A(n13977), .B(n13261), .ZN(n13223) );
  XNOR2_X1 U15616 ( .A(n13223), .B(n13775), .ZN(n13335) );
  INV_X1 U15617 ( .A(n13223), .ZN(n13224) );
  XOR2_X1 U15618 ( .A(n13259), .B(n13260), .Z(n13231) );
  AOI22_X1 U15619 ( .A1(n13349), .A2(n13575), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13227) );
  NAND2_X1 U15620 ( .A1(n13354), .A2(n13225), .ZN(n13226) );
  OAI211_X1 U15621 ( .C1(n13775), .C2(n13352), .A(n13227), .B(n13226), .ZN(
        n13228) );
  AOI21_X1 U15622 ( .B1(n13229), .B2(n13357), .A(n13228), .ZN(n13230) );
  OAI21_X1 U15623 ( .B1(n13231), .B2(n13360), .A(n13230), .ZN(P3_U3154) );
  XNOR2_X1 U15624 ( .A(n13232), .B(n13497), .ZN(n13237) );
  AOI22_X1 U15625 ( .A1(n13349), .A2(n13803), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13234) );
  NAND2_X1 U15626 ( .A1(n13354), .A2(n13801), .ZN(n13233) );
  OAI211_X1 U15627 ( .C1(n13826), .C2(n13352), .A(n13234), .B(n13233), .ZN(
        n13235) );
  AOI21_X1 U15628 ( .B1(n13984), .B2(n13357), .A(n13235), .ZN(n13236) );
  OAI21_X1 U15629 ( .B1(n13237), .B2(n13360), .A(n13236), .ZN(P3_U3156) );
  AND2_X1 U15630 ( .A1(n11807), .A2(n13238), .ZN(n13241) );
  OAI211_X1 U15631 ( .C1(n13241), .C2(n13240), .A(n13325), .B(n13239), .ZN(
        n13247) );
  MUX2_X1 U15632 ( .A(n13242), .B(P3_STATE_REG_SCAN_IN), .S(
        P3_REG3_REG_3__SCAN_IN), .Z(n13246) );
  AOI22_X1 U15633 ( .A1(n13349), .A2(n13589), .B1(n13357), .B2(n13243), .ZN(
        n13245) );
  OR2_X1 U15634 ( .A1(n13352), .A2(n15915), .ZN(n13244) );
  NAND4_X1 U15635 ( .A1(n13247), .A2(n13246), .A3(n13245), .A4(n13244), .ZN(
        P3_U3158) );
  INV_X1 U15636 ( .A(n13248), .ZN(n13249) );
  AOI21_X1 U15637 ( .B1(n13251), .B2(n13250), .A(n13249), .ZN(n13257) );
  NAND2_X1 U15638 ( .A1(n13252), .A2(n13349), .ZN(n13253) );
  NAND2_X1 U15639 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13744)
         );
  OAI211_X1 U15640 ( .C1(n13848), .C2(n13352), .A(n13253), .B(n13744), .ZN(
        n13255) );
  NOR2_X1 U15641 ( .A1(n13853), .A2(n13333), .ZN(n13254) );
  AOI211_X1 U15642 ( .C1(n13850), .C2(n13354), .A(n13255), .B(n13254), .ZN(
        n13256) );
  OAI21_X1 U15643 ( .B1(n13257), .B2(n13360), .A(n13256), .ZN(P3_U3159) );
  XNOR2_X1 U15644 ( .A(n13557), .B(n13261), .ZN(n13262) );
  AOI22_X1 U15645 ( .A1(n13263), .A2(n13768), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13266) );
  NAND2_X1 U15646 ( .A1(n13354), .A2(n13264), .ZN(n13265) );
  OAI211_X1 U15647 ( .C1(n13267), .C2(n13319), .A(n13266), .B(n13265), .ZN(
        n13268) );
  AOI21_X1 U15648 ( .B1(n13269), .B2(n13357), .A(n13268), .ZN(n13270) );
  OAI21_X1 U15649 ( .B1(n6730), .B2(n13272), .A(n13271), .ZN(n13273) );
  NAND2_X1 U15650 ( .A1(n13273), .A2(n13325), .ZN(n13278) );
  OAI22_X1 U15651 ( .A1(n13352), .A2(n13849), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13274), .ZN(n13276) );
  NOR2_X1 U15652 ( .A1(n13826), .A2(n13319), .ZN(n13275) );
  AOI211_X1 U15653 ( .C1(n13818), .C2(n13354), .A(n13276), .B(n13275), .ZN(
        n13277) );
  OAI211_X1 U15654 ( .C1(n13279), .C2(n13333), .A(n13278), .B(n13277), .ZN(
        P3_U3163) );
  XOR2_X1 U15655 ( .A(n13281), .B(n13280), .Z(n13287) );
  AOI22_X1 U15656 ( .A1(n13282), .A2(n13576), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13284) );
  NAND2_X1 U15657 ( .A1(n13354), .A2(n13782), .ZN(n13283) );
  OAI211_X1 U15658 ( .C1(n13776), .C2(n13352), .A(n13284), .B(n13283), .ZN(
        n13285) );
  AOI21_X1 U15659 ( .B1(n13908), .B2(n13357), .A(n13285), .ZN(n13286) );
  OAI21_X1 U15660 ( .B1(n13287), .B2(n13360), .A(n13286), .ZN(P3_U3165) );
  INV_X1 U15661 ( .A(n13288), .ZN(n13291) );
  XNOR2_X1 U15662 ( .A(n13289), .B(n13890), .ZN(n13290) );
  XNOR2_X1 U15663 ( .A(n13291), .B(n13290), .ZN(n13292) );
  NAND2_X1 U15664 ( .A1(n13292), .A2(n13325), .ZN(n13299) );
  NAND2_X1 U15665 ( .A1(n13349), .A2(n13578), .ZN(n13293) );
  NAND2_X1 U15666 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n13669)
         );
  OAI211_X1 U15667 ( .C1(n13352), .C2(n13344), .A(n13293), .B(n13669), .ZN(
        n13294) );
  INV_X1 U15668 ( .A(n13294), .ZN(n13298) );
  NAND2_X1 U15669 ( .A1(n13476), .A2(n13357), .ZN(n13297) );
  NAND2_X1 U15670 ( .A1(n13354), .A2(n13295), .ZN(n13296) );
  NAND4_X1 U15671 ( .A1(n13299), .A2(n13298), .A3(n13297), .A4(n13296), .ZN(
        P3_U3166) );
  INV_X1 U15672 ( .A(n14017), .ZN(n13308) );
  AOI21_X1 U15673 ( .B1(n13301), .B2(n13300), .A(n13360), .ZN(n13303) );
  NAND2_X1 U15674 ( .A1(n13303), .A2(n13302), .ZN(n13307) );
  NAND2_X1 U15675 ( .A1(n13349), .A2(n13887), .ZN(n13304) );
  NAND2_X1 U15676 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13695)
         );
  OAI211_X1 U15677 ( .C1(n13352), .C2(n13475), .A(n13304), .B(n13695), .ZN(
        n13305) );
  AOI21_X1 U15678 ( .B1(n13879), .B2(n13354), .A(n13305), .ZN(n13306) );
  OAI211_X1 U15679 ( .C1(n13308), .C2(n13333), .A(n13307), .B(n13306), .ZN(
        P3_U3168) );
  AOI21_X1 U15680 ( .B1(n13310), .B2(n13309), .A(n13360), .ZN(n13312) );
  NAND2_X1 U15681 ( .A1(n13312), .A2(n13311), .ZN(n13316) );
  AOI22_X1 U15682 ( .A1(n13811), .A2(n13349), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13313) );
  OAI21_X1 U15683 ( .B1(n13864), .B2(n13352), .A(n13313), .ZN(n13314) );
  AOI21_X1 U15684 ( .B1(n13830), .B2(n13354), .A(n13314), .ZN(n13315) );
  OAI211_X1 U15685 ( .C1(n13998), .C2(n13333), .A(n13316), .B(n13315), .ZN(
        P3_U3173) );
  XNOR2_X1 U15686 ( .A(n13317), .B(n13805), .ZN(n13324) );
  INV_X1 U15687 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n13318) );
  OAI22_X1 U15688 ( .A1(n13836), .A2(n13352), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13318), .ZN(n13321) );
  NOR2_X1 U15689 ( .A1(n13497), .A2(n13319), .ZN(n13320) );
  AOI211_X1 U15690 ( .C1(n13809), .C2(n13354), .A(n13321), .B(n13320), .ZN(
        n13323) );
  NAND2_X1 U15691 ( .A1(n13990), .A2(n13357), .ZN(n13322) );
  OAI211_X1 U15692 ( .C1(n13324), .C2(n13360), .A(n13323), .B(n13322), .ZN(
        P3_U3175) );
  INV_X1 U15693 ( .A(n13874), .ZN(n14014) );
  OAI211_X1 U15694 ( .C1(n13328), .C2(n13327), .A(n13326), .B(n13325), .ZN(
        n13332) );
  NAND2_X1 U15695 ( .A1(n13349), .A2(n8429), .ZN(n13329) );
  NAND2_X1 U15696 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13710)
         );
  OAI211_X1 U15697 ( .C1(n13352), .C2(n13865), .A(n13329), .B(n13710), .ZN(
        n13330) );
  AOI21_X1 U15698 ( .B1(n13866), .B2(n13354), .A(n13330), .ZN(n13331) );
  OAI211_X1 U15699 ( .C1(n14014), .C2(n13333), .A(n13332), .B(n13331), .ZN(
        P3_U3178) );
  XOR2_X1 U15700 ( .A(n13335), .B(n13334), .Z(n13341) );
  AOI22_X1 U15701 ( .A1(n13349), .A2(n13768), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13337) );
  NAND2_X1 U15702 ( .A1(n13354), .A2(n13770), .ZN(n13336) );
  OAI211_X1 U15703 ( .C1(n13338), .C2(n13352), .A(n13337), .B(n13336), .ZN(
        n13339) );
  AOI21_X1 U15704 ( .B1(n13977), .B2(n13357), .A(n13339), .ZN(n13340) );
  OAI21_X1 U15705 ( .B1(n13341), .B2(n13360), .A(n13340), .ZN(P3_U3180) );
  INV_X1 U15706 ( .A(n13342), .ZN(n13345) );
  NAND2_X1 U15707 ( .A1(n13345), .A2(n13344), .ZN(n13343) );
  OAI21_X1 U15708 ( .B1(n13345), .B2(n13344), .A(n13343), .ZN(n13347) );
  NOR2_X1 U15709 ( .A1(n13347), .A2(n13348), .ZN(n13346) );
  AOI21_X1 U15710 ( .B1(n13348), .B2(n13347), .A(n13346), .ZN(n13361) );
  NAND2_X1 U15711 ( .A1(n13349), .A2(n13890), .ZN(n13350) );
  NAND2_X1 U15712 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n13646)
         );
  OAI211_X1 U15713 ( .C1(n13352), .C2(n13351), .A(n13350), .B(n13646), .ZN(
        n13353) );
  AOI21_X1 U15714 ( .B1(n13355), .B2(n13354), .A(n13353), .ZN(n13359) );
  NAND2_X1 U15715 ( .A1(n13357), .A2(n13356), .ZN(n13358) );
  OAI211_X1 U15716 ( .C1(n13361), .C2(n13360), .A(n13359), .B(n13358), .ZN(
        P3_U3181) );
  INV_X1 U15717 ( .A(n13362), .ZN(n13363) );
  NAND2_X1 U15718 ( .A1(n13363), .A2(n13517), .ZN(n13401) );
  NAND2_X1 U15719 ( .A1(n13365), .A2(n13364), .ZN(n13368) );
  INV_X1 U15720 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13366) );
  XNOR2_X1 U15721 ( .A(n13366), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n13367) );
  XNOR2_X1 U15722 ( .A(n13368), .B(n13367), .ZN(n14029) );
  NAND2_X1 U15723 ( .A1(n14029), .A2(n13369), .ZN(n13371) );
  OR2_X1 U15724 ( .A1(n8176), .A2(n10312), .ZN(n13370) );
  OR2_X1 U15725 ( .A1(n13968), .A2(n13745), .ZN(n13384) );
  OR2_X1 U15726 ( .A1(n8176), .A2(n13374), .ZN(n13375) );
  INV_X1 U15727 ( .A(n13385), .ZN(n13573) );
  AND2_X1 U15728 ( .A1(n13974), .A2(n13573), .ZN(n13527) );
  INV_X1 U15729 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n13971) );
  OR2_X1 U15730 ( .A1(n13376), .A2(n13971), .ZN(n13380) );
  NAND2_X1 U15731 ( .A1(n8199), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n13379) );
  INV_X1 U15732 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n13762) );
  OR2_X1 U15733 ( .A1(n13377), .A2(n13762), .ZN(n13378) );
  INV_X1 U15734 ( .A(n13758), .ZN(n13572) );
  NAND2_X1 U15735 ( .A1(n13572), .A2(n13735), .ZN(n13388) );
  INV_X1 U15736 ( .A(n13388), .ZN(n13382) );
  NAND2_X1 U15737 ( .A1(n8031), .A2(n13382), .ZN(n13383) );
  NAND2_X1 U15738 ( .A1(n13384), .A2(n13383), .ZN(n13394) );
  INV_X1 U15739 ( .A(n13394), .ZN(n13400) );
  OR2_X1 U15740 ( .A1(n13968), .A2(n13758), .ZN(n13387) );
  NAND2_X1 U15741 ( .A1(n7596), .A2(n13385), .ZN(n13386) );
  INV_X1 U15742 ( .A(n13968), .ZN(n13896) );
  AOI211_X1 U15743 ( .C1(n13572), .C2(n8031), .A(n13735), .B(n13896), .ZN(
        n13392) );
  AOI211_X1 U15744 ( .C1(n13974), .C2(n13520), .A(n13745), .B(n13968), .ZN(
        n13391) );
  NOR3_X1 U15745 ( .A1(n13527), .A2(n13520), .A3(n13388), .ZN(n13390) );
  OR4_X1 U15746 ( .A1(n13392), .A2(n13391), .A3(n13390), .A4(n13389), .ZN(
        n13393) );
  AOI21_X1 U15747 ( .B1(n13559), .B2(n13394), .A(n13393), .ZN(n13399) );
  INV_X1 U15748 ( .A(n13520), .ZN(n13395) );
  AOI211_X1 U15749 ( .C1(n13758), .C2(n7596), .A(n13735), .B(n13395), .ZN(
        n13396) );
  AND2_X1 U15750 ( .A1(n13396), .A2(n7230), .ZN(n13397) );
  NAND2_X1 U15751 ( .A1(n13401), .A2(n13397), .ZN(n13398) );
  INV_X1 U15752 ( .A(n13480), .ZN(n13403) );
  NOR2_X1 U15753 ( .A1(n13403), .A2(n13402), .ZN(n13405) );
  AND2_X1 U15754 ( .A1(n13853), .A2(n8429), .ZN(n13484) );
  NOR4_X1 U15755 ( .A1(n13405), .A2(n13484), .A3(n13404), .A4(n13514), .ZN(
        n13479) );
  INV_X1 U15756 ( .A(n13407), .ZN(n13408) );
  AOI211_X1 U15757 ( .C1(n13453), .C2(n7791), .A(n13408), .B(n13458), .ZN(
        n13452) );
  INV_X1 U15758 ( .A(n13411), .ZN(n13418) );
  OAI21_X1 U15759 ( .B1(n13409), .B2(n13412), .A(n13514), .ZN(n13414) );
  NAND3_X1 U15760 ( .A1(n13411), .A2(n13410), .A3(n13570), .ZN(n13413) );
  AOI22_X1 U15761 ( .A1(n13414), .A2(n13413), .B1(n15904), .B2(n13412), .ZN(
        n13416) );
  MUX2_X1 U15762 ( .A(n13519), .B(n13416), .S(n13415), .Z(n13417) );
  NAND2_X1 U15763 ( .A1(n13420), .A2(n13419), .ZN(n13423) );
  NAND2_X1 U15764 ( .A1(n13591), .A2(n13965), .ZN(n13421) );
  NAND2_X1 U15765 ( .A1(n13427), .A2(n13421), .ZN(n13422) );
  MUX2_X1 U15766 ( .A(n13423), .B(n13422), .S(n13519), .Z(n13424) );
  INV_X1 U15767 ( .A(n13427), .ZN(n13429) );
  INV_X1 U15768 ( .A(n13430), .ZN(n13431) );
  NAND2_X1 U15769 ( .A1(n13435), .A2(n13433), .ZN(n13434) );
  AOI211_X1 U15770 ( .C1(n13438), .C2(n13514), .A(n13437), .B(n13436), .ZN(
        n13446) );
  MUX2_X1 U15771 ( .A(n13440), .B(n13439), .S(n13514), .Z(n13441) );
  NAND2_X1 U15772 ( .A1(n13538), .A2(n13441), .ZN(n13445) );
  MUX2_X1 U15773 ( .A(n13443), .B(n13442), .S(n13514), .Z(n13444) );
  OAI211_X1 U15774 ( .C1(n13446), .C2(n13445), .A(n13537), .B(n13444), .ZN(
        n13451) );
  INV_X1 U15775 ( .A(n13541), .ZN(n13450) );
  MUX2_X1 U15776 ( .A(n13448), .B(n13447), .S(n13514), .Z(n13449) );
  OAI211_X1 U15777 ( .C1(n6889), .C2(n13455), .A(n13457), .B(n13454), .ZN(
        n13456) );
  MUX2_X1 U15778 ( .A(n13460), .B(n13459), .S(n13514), .Z(n13461) );
  NAND2_X1 U15779 ( .A1(n13549), .A2(n13461), .ZN(n13463) );
  OAI22_X1 U15780 ( .A1(n13464), .A2(n13463), .B1(n13462), .B2(n13514), .ZN(
        n13470) );
  NAND3_X1 U15781 ( .A1(n13469), .A2(n13579), .A3(n13465), .ZN(n13467) );
  OAI211_X1 U15782 ( .C1(n13475), .C2(n13476), .A(n13467), .B(n13466), .ZN(
        n13468) );
  AOI22_X1 U15783 ( .A1(n13470), .A2(n13469), .B1(n13514), .B2(n13468), .ZN(
        n13471) );
  AOI21_X1 U15784 ( .B1(n13474), .B2(n13472), .A(n13514), .ZN(n13473) );
  NOR3_X1 U15785 ( .A1(n13476), .A2(n13475), .A3(n13514), .ZN(n13477) );
  INV_X1 U15786 ( .A(n13479), .ZN(n13482) );
  NAND3_X1 U15787 ( .A1(n13483), .A2(n13480), .A3(n13514), .ZN(n13481) );
  INV_X1 U15788 ( .A(n13483), .ZN(n13485) );
  MUX2_X1 U15789 ( .A(n13485), .B(n13484), .S(n13514), .Z(n13486) );
  MUX2_X1 U15790 ( .A(n13488), .B(n13487), .S(n13514), .Z(n13490) );
  INV_X1 U15791 ( .A(n13824), .ZN(n13489) );
  MUX2_X1 U15792 ( .A(n13492), .B(n13491), .S(n13514), .Z(n13493) );
  INV_X1 U15793 ( .A(n13550), .ZN(n13810) );
  MUX2_X1 U15794 ( .A(n13495), .B(n13494), .S(n13514), .Z(n13496) );
  NAND3_X1 U15795 ( .A1(n13984), .A2(n13497), .A3(n13519), .ZN(n13498) );
  INV_X1 U15796 ( .A(n13499), .ZN(n13503) );
  AOI21_X1 U15797 ( .B1(n13501), .B2(n13500), .A(n13503), .ZN(n13502) );
  MUX2_X1 U15798 ( .A(n13503), .B(n13502), .S(n13514), .Z(n13504) );
  INV_X1 U15799 ( .A(n13766), .ZN(n13508) );
  MUX2_X1 U15800 ( .A(n13506), .B(n13505), .S(n13514), .Z(n13507) );
  NAND2_X1 U15801 ( .A1(n13508), .A2(n13507), .ZN(n13512) );
  MUX2_X1 U15802 ( .A(n13510), .B(n13509), .S(n13514), .Z(n13511) );
  OAI21_X1 U15803 ( .B1(n13513), .B2(n13512), .A(n13511), .ZN(n13518) );
  NAND3_X1 U15804 ( .A1(n13518), .A2(n13530), .A3(n13514), .ZN(n13516) );
  NAND2_X1 U15805 ( .A1(n13521), .A2(n13520), .ZN(n13526) );
  NAND2_X1 U15806 ( .A1(n13523), .A2(n13522), .ZN(n13525) );
  AND2_X1 U15807 ( .A1(n13968), .A2(n13758), .ZN(n13556) );
  XNOR2_X1 U15808 ( .A(n13853), .B(n8429), .ZN(n13845) );
  NOR2_X1 U15809 ( .A1(n11594), .A2(n13531), .ZN(n13535) );
  NAND4_X1 U15810 ( .A1(n13540), .A2(n13539), .A3(n13538), .A4(n13537), .ZN(
        n13543) );
  OR3_X1 U15811 ( .A1(n13546), .A2(n13545), .A3(n13544), .ZN(n13547) );
  OR4_X1 U15812 ( .A1(n13551), .A2(n13550), .A3(n13845), .A4(n6744), .ZN(
        n13552) );
  NOR2_X1 U15813 ( .A1(n13552), .A2(n8004), .ZN(n13553) );
  NAND4_X1 U15814 ( .A1(n13780), .A2(n13793), .A3(n13824), .A4(n13553), .ZN(
        n13554) );
  NOR4_X1 U15815 ( .A1(n13555), .A2(n6855), .A3(n13766), .A4(n13554), .ZN(
        n13558) );
  XNOR2_X1 U15816 ( .A(n13560), .B(n13745), .ZN(n13562) );
  NAND2_X1 U15817 ( .A1(n13562), .A2(n13561), .ZN(n13563) );
  INV_X1 U15818 ( .A(n13569), .ZN(n13564) );
  NAND4_X1 U15819 ( .A1(n13567), .A2(n13566), .A3(n13889), .A4(n13565), .ZN(
        n13568) );
  OAI211_X1 U15820 ( .C1(n13570), .C2(n13569), .A(n13568), .B(P3_B_REG_SCAN_IN), .ZN(n13571) );
  MUX2_X1 U15821 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n13572), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U15822 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n13573), .S(P3_U3897), .Z(
        P3_U3521) );
  MUX2_X1 U15823 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n13574), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U15824 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n13575), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U15825 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n13768), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15826 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n13576), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U15827 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n13790), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U15828 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n13803), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U15829 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n13812), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U15830 ( .A(n8429), .B(P3_DATAO_REG_19__SCAN_IN), .S(n13577), .Z(
        P3_U3510) );
  MUX2_X1 U15831 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13887), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15832 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n13578), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U15833 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n13890), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U15834 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n13579), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U15835 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n13580), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U15836 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n13581), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U15837 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n13582), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U15838 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n13583), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U15839 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n13584), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U15840 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n13585), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U15841 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n13586), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U15842 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n13587), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U15843 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n13588), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U15844 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n13589), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U15845 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n13590), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U15846 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n13591), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15847 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n15906), .S(P3_U3897), .Z(
        P3_U3491) );
  NAND2_X1 U15848 ( .A1(n13722), .A2(n13593), .ZN(n13606) );
  OAI21_X1 U15849 ( .B1(n6787), .B2(P3_REG2_REG_3__SCAN_IN), .A(n13594), .ZN(
        n13597) );
  OAI21_X1 U15850 ( .B1(n6785), .B2(P3_REG1_REG_3__SCAN_IN), .A(n13595), .ZN(
        n13596) );
  AOI22_X1 U15851 ( .A1(n13667), .A2(n13597), .B1(n13754), .B2(n13596), .ZN(
        n13605) );
  AOI22_X1 U15852 ( .A1(n15894), .A2(P3_ADDR_REG_3__SCAN_IN), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(P3_U3151), .ZN(n13604) );
  INV_X1 U15853 ( .A(n13598), .ZN(n13602) );
  NOR3_X1 U15854 ( .A1(n13600), .A2(n13599), .A3(n8094), .ZN(n13601) );
  OAI21_X1 U15855 ( .B1(n13602), .B2(n13601), .A(n13748), .ZN(n13603) );
  NAND4_X1 U15856 ( .A1(n13606), .A2(n13605), .A3(n13604), .A4(n13603), .ZN(
        P3_U3185) );
  AND3_X1 U15857 ( .A1(n13608), .A2(n13607), .A3(n6930), .ZN(n13609) );
  OAI21_X1 U15858 ( .B1(n13610), .B2(n13609), .A(n13667), .ZN(n13624) );
  INV_X1 U15859 ( .A(n15894), .ZN(n13711) );
  INV_X1 U15860 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n13612) );
  OAI21_X1 U15861 ( .B1(n13711), .B2(n13612), .A(n13611), .ZN(n13613) );
  AOI21_X1 U15862 ( .B1(n13722), .B2(n13614), .A(n13613), .ZN(n13623) );
  OAI21_X1 U15863 ( .B1(n13617), .B2(n13616), .A(n13615), .ZN(n13618) );
  NAND2_X1 U15864 ( .A1(n13618), .A2(n13754), .ZN(n13622) );
  OAI211_X1 U15865 ( .C1(n13620), .C2(n13619), .A(n13631), .B(n13748), .ZN(
        n13621) );
  NAND4_X1 U15866 ( .A1(n13624), .A2(n13623), .A3(n13622), .A4(n13621), .ZN(
        P3_U3194) );
  AOI21_X1 U15867 ( .B1(n13627), .B2(n13626), .A(n13625), .ZN(n13641) );
  INV_X1 U15868 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15566) );
  OAI21_X1 U15869 ( .B1(n13711), .B2(n15566), .A(n13628), .ZN(n13636) );
  AOI21_X1 U15870 ( .B1(n13631), .B2(n13630), .A(n13629), .ZN(n13632) );
  INV_X1 U15871 ( .A(n13632), .ZN(n13634) );
  AOI21_X1 U15872 ( .B1(n13634), .B2(n13633), .A(n13720), .ZN(n13635) );
  AOI211_X1 U15873 ( .C1(n13722), .C2(n7091), .A(n13636), .B(n13635), .ZN(
        n13640) );
  OAI21_X1 U15874 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n6746), .A(n13637), .ZN(
        n13638) );
  NAND2_X1 U15875 ( .A1(n13638), .A2(n13754), .ZN(n13639) );
  OAI211_X1 U15876 ( .C1(n13641), .C2(n13757), .A(n13640), .B(n13639), .ZN(
        P3_U3195) );
  INV_X1 U15877 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n13645) );
  NAND2_X1 U15878 ( .A1(n13642), .A2(n13647), .ZN(n13643) );
  AOI21_X1 U15879 ( .B1(n13645), .B2(n13644), .A(n13666), .ZN(n13662) );
  INV_X1 U15880 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n15588) );
  OAI21_X1 U15881 ( .B1(n13711), .B2(n15588), .A(n13646), .ZN(n13654) );
  MUX2_X1 U15882 ( .A(n13655), .B(n13647), .S(n13736), .Z(n13648) );
  MUX2_X1 U15883 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n7288), .Z(n13650) );
  AOI21_X1 U15884 ( .B1(n13651), .B2(n13650), .A(n13677), .ZN(n13652) );
  NOR2_X1 U15885 ( .A1(n13652), .A2(n13720), .ZN(n13653) );
  AOI211_X1 U15886 ( .C1(n13722), .C2(n13678), .A(n13654), .B(n13653), .ZN(
        n13661) );
  OAI21_X1 U15887 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n13658), .A(n13674), 
        .ZN(n13659) );
  NAND2_X1 U15888 ( .A1(n13659), .A2(n13754), .ZN(n13660) );
  OAI211_X1 U15889 ( .C1(n13662), .C2(n13757), .A(n13661), .B(n13660), .ZN(
        P3_U3197) );
  INV_X1 U15890 ( .A(n13663), .ZN(n13665) );
  XNOR2_X1 U15891 ( .A(n13693), .B(P3_REG2_REG_16__SCAN_IN), .ZN(n13664) );
  NOR3_X1 U15892 ( .A1(n13666), .A2(n13665), .A3(n13664), .ZN(n13668) );
  OAI21_X1 U15893 ( .B1(n6664), .B2(n13668), .A(n13667), .ZN(n13685) );
  INV_X1 U15894 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n15601) );
  OAI21_X1 U15895 ( .B1(n13711), .B2(n15601), .A(n13669), .ZN(n13670) );
  AOI21_X1 U15896 ( .B1(n13722), .B2(n13693), .A(n13670), .ZN(n13684) );
  XNOR2_X1 U15897 ( .A(n13693), .B(n13671), .ZN(n13673) );
  AND3_X1 U15898 ( .A1(n13674), .A2(n13673), .A3(n13672), .ZN(n13675) );
  OAI21_X1 U15899 ( .B1(n13698), .B2(n13675), .A(n13754), .ZN(n13683) );
  INV_X1 U15900 ( .A(n13676), .ZN(n13679) );
  MUX2_X1 U15901 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n7288), .Z(n13690) );
  XNOR2_X1 U15902 ( .A(n13690), .B(n13693), .ZN(n13680) );
  OAI211_X1 U15903 ( .C1(n13681), .C2(n13680), .A(n13691), .B(n13748), .ZN(
        n13682) );
  NAND4_X1 U15904 ( .A1(n13685), .A2(n13684), .A3(n13683), .A4(n13682), .ZN(
        P3_U3198) );
  NAND2_X1 U15905 ( .A1(n13687), .A2(n13712), .ZN(n13708) );
  OAI21_X1 U15906 ( .B1(n13687), .B2(n13712), .A(n13708), .ZN(n13689) );
  INV_X1 U15907 ( .A(n13709), .ZN(n13688) );
  MUX2_X1 U15908 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n7288), .Z(n13713) );
  XNOR2_X1 U15909 ( .A(n13713), .B(n13700), .ZN(n13714) );
  INV_X1 U15910 ( .A(n13690), .ZN(n13692) );
  XOR2_X1 U15911 ( .A(n13714), .B(n13715), .Z(n13697) );
  NAND2_X1 U15912 ( .A1(n15894), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n13694) );
  OAI211_X1 U15913 ( .C1(n13746), .C2(n13712), .A(n13695), .B(n13694), .ZN(
        n13696) );
  AOI21_X1 U15914 ( .B1(n13697), .B2(n13748), .A(n13696), .ZN(n13705) );
  OAI21_X1 U15915 ( .B1(P3_REG1_REG_17__SCAN_IN), .B2(n13702), .A(n13729), 
        .ZN(n13703) );
  NAND2_X1 U15916 ( .A1(n13703), .A2(n13754), .ZN(n13704) );
  NAND2_X1 U15917 ( .A1(n13724), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n13733) );
  NAND2_X1 U15918 ( .A1(n13725), .A2(n13868), .ZN(n13706) );
  NAND2_X1 U15919 ( .A1(n13733), .A2(n13706), .ZN(n13707) );
  INV_X1 U15920 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15619) );
  OAI21_X1 U15921 ( .B1(n13711), .B2(n15619), .A(n13710), .ZN(n13721) );
  OAI21_X1 U15922 ( .B1(n13716), .B2(n13725), .A(n13738), .ZN(n13719) );
  MUX2_X1 U15923 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n7288), .Z(n13718) );
  INV_X1 U15924 ( .A(n13723), .ZN(n13728) );
  NAND2_X1 U15925 ( .A1(n13724), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n13750) );
  INV_X1 U15926 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13938) );
  NAND2_X1 U15927 ( .A1(n13725), .A2(n13938), .ZN(n13726) );
  NAND2_X1 U15928 ( .A1(n13750), .A2(n13726), .ZN(n13727) );
  AND3_X1 U15929 ( .A1(n13729), .A2(n13728), .A3(n13727), .ZN(n13730) );
  OAI21_X1 U15930 ( .B1(n13752), .B2(n13730), .A(n13754), .ZN(n13731) );
  XNOR2_X1 U15931 ( .A(n13735), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n13737) );
  XNOR2_X1 U15932 ( .A(n13735), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13753) );
  MUX2_X1 U15933 ( .A(n13753), .B(n13737), .S(n13736), .Z(n13742) );
  INV_X1 U15934 ( .A(n13738), .ZN(n13739) );
  NOR2_X1 U15935 ( .A1(n13740), .A2(n13739), .ZN(n13741) );
  XOR2_X1 U15936 ( .A(n13742), .B(n13741), .Z(n13749) );
  NAND2_X1 U15937 ( .A1(n15894), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n13743) );
  OAI211_X1 U15938 ( .C1(n13746), .C2(n13745), .A(n13744), .B(n13743), .ZN(
        n13747) );
  AOI21_X1 U15939 ( .B1(n13749), .B2(n13748), .A(n13747), .ZN(n13756) );
  INV_X1 U15940 ( .A(n13750), .ZN(n13751) );
  NAND2_X1 U15941 ( .A1(n13968), .A2(n13880), .ZN(n13761) );
  NOR2_X1 U15942 ( .A1(n13759), .A2(n13758), .ZN(n13969) );
  AOI21_X1 U15943 ( .B1(n15921), .B2(n13969), .A(n13760), .ZN(n13764) );
  OAI211_X1 U15944 ( .C1(n13762), .C2(n15921), .A(n13761), .B(n13764), .ZN(
        P3_U3202) );
  NAND2_X1 U15945 ( .A1(n15903), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n13763) );
  OAI211_X1 U15946 ( .C1(n13974), .C2(n13852), .A(n13764), .B(n13763), .ZN(
        P3_U3203) );
  XNOR2_X1 U15947 ( .A(n13765), .B(n13766), .ZN(n13979) );
  MUX2_X1 U15948 ( .A(n13769), .B(n13975), .S(n15921), .Z(n13772) );
  AOI22_X1 U15949 ( .A1(n13977), .A2(n13880), .B1(n15901), .B2(n13770), .ZN(
        n13771) );
  OAI211_X1 U15950 ( .C1(n13979), .C2(n13894), .A(n13772), .B(n13771), .ZN(
        P3_U3207) );
  AOI211_X1 U15951 ( .C1(n13780), .C2(n13774), .A(n15911), .B(n13773), .ZN(
        n13778) );
  OAI22_X1 U15952 ( .A1(n13776), .A2(n15914), .B1(n15916), .B2(n13775), .ZN(
        n13777) );
  NOR2_X1 U15953 ( .A1(n13778), .A2(n13777), .ZN(n13910) );
  OAI21_X1 U15954 ( .B1(n13781), .B2(n13780), .A(n13779), .ZN(n13909) );
  INV_X1 U15955 ( .A(n13908), .ZN(n13784) );
  AOI22_X1 U15956 ( .A1(n15903), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n15901), 
        .B2(n13782), .ZN(n13783) );
  OAI21_X1 U15957 ( .B1(n13784), .B2(n13852), .A(n13783), .ZN(n13785) );
  AOI21_X1 U15958 ( .B1(n13909), .B2(n13856), .A(n13785), .ZN(n13786) );
  OAI21_X1 U15959 ( .B1(n15903), .B2(n13910), .A(n13786), .ZN(P3_U3208) );
  OAI21_X1 U15960 ( .B1(n13789), .B2(n13788), .A(n13787), .ZN(n13791) );
  AOI222_X1 U15961 ( .A1(n13791), .A2(n13960), .B1(n13790), .B2(n13886), .C1(
        n13812), .C2(n13889), .ZN(n13914) );
  OAI21_X1 U15962 ( .B1(n13794), .B2(n13793), .A(n13792), .ZN(n13913) );
  INV_X1 U15963 ( .A(n13912), .ZN(n13797) );
  AOI22_X1 U15964 ( .A1(n15903), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n15901), 
        .B2(n13795), .ZN(n13796) );
  OAI21_X1 U15965 ( .B1(n13797), .B2(n13852), .A(n13796), .ZN(n13798) );
  AOI21_X1 U15966 ( .B1(n13913), .B2(n13856), .A(n13798), .ZN(n13799) );
  OAI21_X1 U15967 ( .B1(n15903), .B2(n13914), .A(n13799), .ZN(P3_U3209) );
  XNOR2_X1 U15968 ( .A(n13800), .B(n7408), .ZN(n13987) );
  AOI22_X1 U15969 ( .A1(n13984), .A2(n13880), .B1(n15901), .B2(n13801), .ZN(
        n13807) );
  XNOR2_X1 U15970 ( .A(n13802), .B(n7408), .ZN(n13804) );
  AOI222_X1 U15971 ( .A1(n13805), .A2(n13889), .B1(n13960), .B2(n13804), .C1(
        n13803), .C2(n13886), .ZN(n13982) );
  MUX2_X1 U15972 ( .A(n10446), .B(n13982), .S(n15921), .Z(n13806) );
  OAI211_X1 U15973 ( .C1(n13987), .C2(n13894), .A(n13807), .B(n13806), .ZN(
        P3_U3210) );
  XNOR2_X1 U15974 ( .A(n13808), .B(n13810), .ZN(n13993) );
  AOI22_X1 U15975 ( .A1(n13990), .A2(n13880), .B1(n15901), .B2(n13809), .ZN(
        n13816) );
  XNOR2_X1 U15976 ( .A(n6708), .B(n13810), .ZN(n13813) );
  AOI222_X1 U15977 ( .A1(n13813), .A2(n13960), .B1(n13812), .B2(n13886), .C1(
        n13811), .C2(n13889), .ZN(n13988) );
  MUX2_X1 U15978 ( .A(n13814), .B(n13988), .S(n15921), .Z(n13815) );
  OAI211_X1 U15979 ( .C1(n13993), .C2(n13894), .A(n13816), .B(n13815), .ZN(
        P3_U3211) );
  XNOR2_X1 U15980 ( .A(n13817), .B(n13824), .ZN(n13997) );
  INV_X1 U15981 ( .A(n13818), .ZN(n13819) );
  OAI22_X1 U15982 ( .A1(n15921), .A2(n13820), .B1(n13819), .B2(n15923), .ZN(
        n13821) );
  AOI21_X1 U15983 ( .B1(n13923), .B2(n13880), .A(n13821), .ZN(n13828) );
  AOI21_X1 U15984 ( .B1(n13824), .B2(n13823), .A(n13822), .ZN(n13825) );
  OAI222_X1 U15985 ( .A1(n15916), .A2(n13826), .B1(n15914), .B2(n13849), .C1(
        n13825), .C2(n15911), .ZN(n13922) );
  NAND2_X1 U15986 ( .A1(n13922), .A2(n15921), .ZN(n13827) );
  OAI211_X1 U15987 ( .C1(n13997), .C2(n13894), .A(n13828), .B(n13827), .ZN(
        P3_U3212) );
  XNOR2_X1 U15988 ( .A(n13829), .B(n13832), .ZN(n13999) );
  AOI22_X1 U15989 ( .A1(n13831), .A2(n13880), .B1(n15901), .B2(n13830), .ZN(
        n13842) );
  NAND2_X1 U15990 ( .A1(n13833), .A2(n13832), .ZN(n13834) );
  NAND3_X1 U15991 ( .A1(n13835), .A2(n13960), .A3(n13834), .ZN(n13839) );
  OAI22_X1 U15992 ( .A1(n13836), .A2(n15916), .B1(n13864), .B2(n15914), .ZN(
        n13837) );
  INV_X1 U15993 ( .A(n13837), .ZN(n13838) );
  NAND2_X1 U15994 ( .A1(n13839), .A2(n13838), .ZN(n14000) );
  MUX2_X1 U15995 ( .A(n14000), .B(P3_REG2_REG_20__SCAN_IN), .S(n15903), .Z(
        n13840) );
  INV_X1 U15996 ( .A(n13840), .ZN(n13841) );
  OAI211_X1 U15997 ( .C1(n13999), .C2(n13894), .A(n13842), .B(n13841), .ZN(
        P3_U3213) );
  NAND2_X1 U15998 ( .A1(n13870), .A2(n13869), .ZN(n13936) );
  NAND2_X1 U15999 ( .A1(n13936), .A2(n13843), .ZN(n13844) );
  XNOR2_X1 U16000 ( .A(n13844), .B(n13845), .ZN(n14005) );
  XOR2_X1 U16001 ( .A(n13846), .B(n13845), .Z(n13847) );
  OAI222_X1 U16002 ( .A1(n15916), .A2(n13849), .B1(n15914), .B2(n13848), .C1(
        n13847), .C2(n15911), .ZN(n13929) );
  MUX2_X1 U16003 ( .A(P3_REG2_REG_19__SCAN_IN), .B(n13929), .S(n15921), .Z(
        n13855) );
  INV_X1 U16004 ( .A(n13850), .ZN(n13851) );
  OAI22_X1 U16005 ( .A1(n13853), .A2(n13852), .B1(n13851), .B2(n15923), .ZN(
        n13854) );
  AOI211_X1 U16006 ( .C1(n14005), .C2(n13856), .A(n13855), .B(n13854), .ZN(
        n13857) );
  INV_X1 U16007 ( .A(n13857), .ZN(P3_U3214) );
  NAND2_X1 U16008 ( .A1(n13859), .A2(n13858), .ZN(n13862) );
  INV_X1 U16009 ( .A(n13860), .ZN(n13861) );
  AOI21_X1 U16010 ( .B1(n13869), .B2(n13862), .A(n13861), .ZN(n13863) );
  OAI222_X1 U16011 ( .A1(n15914), .A2(n13865), .B1(n15916), .B2(n13864), .C1(
        n13863), .C2(n15911), .ZN(n13935) );
  INV_X1 U16012 ( .A(n13935), .ZN(n13876) );
  INV_X1 U16013 ( .A(n13866), .ZN(n13867) );
  OAI22_X1 U16014 ( .A1(n15921), .A2(n13868), .B1(n13867), .B2(n15923), .ZN(
        n13873) );
  NOR2_X1 U16015 ( .A1(n13870), .A2(n13869), .ZN(n13934) );
  INV_X1 U16016 ( .A(n13936), .ZN(n13871) );
  NOR3_X1 U16017 ( .A1(n13934), .A2(n13871), .A3(n13894), .ZN(n13872) );
  AOI211_X1 U16018 ( .C1(n13880), .C2(n13874), .A(n13873), .B(n13872), .ZN(
        n13875) );
  OAI21_X1 U16019 ( .B1(n15903), .B2(n13876), .A(n13875), .ZN(P3_U3215) );
  XNOR2_X1 U16020 ( .A(n13878), .B(n13877), .ZN(n14022) );
  AOI22_X1 U16021 ( .A1(n13880), .A2(n14017), .B1(n15901), .B2(n13879), .ZN(
        n13893) );
  NAND2_X1 U16022 ( .A1(n13882), .A2(n13881), .ZN(n13884) );
  NAND2_X1 U16023 ( .A1(n13884), .A2(n13883), .ZN(n13885) );
  XNOR2_X1 U16024 ( .A(n13885), .B(n8656), .ZN(n13888) );
  AOI222_X1 U16025 ( .A1(n13890), .A2(n13889), .B1(n13960), .B2(n13888), .C1(
        n13887), .C2(n13886), .ZN(n14015) );
  MUX2_X1 U16026 ( .A(n13891), .B(n14015), .S(n15921), .Z(n13892) );
  OAI211_X1 U16027 ( .C1(n14022), .C2(n13894), .A(n13893), .B(n13892), .ZN(
        P3_U3216) );
  NAND2_X1 U16028 ( .A1(n15973), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n13895) );
  NAND2_X1 U16029 ( .A1(n15976), .A2(n13969), .ZN(n13898) );
  OAI211_X1 U16030 ( .C1(n13896), .C2(n13940), .A(n13895), .B(n13898), .ZN(
        P3_U3490) );
  NAND2_X1 U16031 ( .A1(n15973), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n13897) );
  OAI211_X1 U16032 ( .C1(n13974), .C2(n13940), .A(n13898), .B(n13897), .ZN(
        P3_U3489) );
  OR2_X1 U16033 ( .A1(n13901), .A2(n13945), .ZN(n13904) );
  NAND2_X1 U16034 ( .A1(n13902), .A2(n13942), .ZN(n13903) );
  INV_X1 U16035 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13905) );
  MUX2_X1 U16036 ( .A(n13905), .B(n13975), .S(n15976), .Z(n13907) );
  NAND2_X1 U16037 ( .A1(n13977), .A2(n13942), .ZN(n13906) );
  OAI211_X1 U16038 ( .C1(n13945), .C2(n13979), .A(n13907), .B(n13906), .ZN(
        P3_U3485) );
  INV_X1 U16039 ( .A(n13933), .ZN(n15928) );
  AOI22_X1 U16040 ( .A1(n13909), .A2(n15928), .B1(n15944), .B2(n13908), .ZN(
        n13911) );
  NAND2_X1 U16041 ( .A1(n13911), .A2(n13910), .ZN(n13980) );
  MUX2_X1 U16042 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n13980), .S(n15976), .Z(
        P3_U3484) );
  AOI22_X1 U16043 ( .A1(n13913), .A2(n15928), .B1(n15944), .B2(n13912), .ZN(
        n13915) );
  NAND2_X1 U16044 ( .A1(n13915), .A2(n13914), .ZN(n13981) );
  MUX2_X1 U16045 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n13981), .S(n15976), .Z(
        P3_U3483) );
  INV_X1 U16046 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13916) );
  MUX2_X1 U16047 ( .A(n13916), .B(n13982), .S(n15976), .Z(n13918) );
  NAND2_X1 U16048 ( .A1(n13984), .A2(n13942), .ZN(n13917) );
  OAI211_X1 U16049 ( .C1(n13987), .C2(n13945), .A(n13918), .B(n13917), .ZN(
        P3_U3482) );
  INV_X1 U16050 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13919) );
  MUX2_X1 U16051 ( .A(n13919), .B(n13988), .S(n15976), .Z(n13921) );
  NAND2_X1 U16052 ( .A1(n13990), .A2(n13942), .ZN(n13920) );
  OAI211_X1 U16053 ( .C1(n13993), .C2(n13945), .A(n13921), .B(n13920), .ZN(
        P3_U3481) );
  INV_X1 U16054 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13924) );
  AOI21_X1 U16055 ( .B1(n15944), .B2(n13923), .A(n13922), .ZN(n13994) );
  MUX2_X1 U16056 ( .A(n13924), .B(n13994), .S(n15976), .Z(n13925) );
  OAI21_X1 U16057 ( .B1(n13997), .B2(n13945), .A(n13925), .ZN(P3_U3480) );
  OAI22_X1 U16058 ( .A1(n13999), .A2(n13945), .B1(n13998), .B2(n13940), .ZN(
        n13927) );
  MUX2_X1 U16059 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n14000), .S(n15976), .Z(
        n13926) );
  OR2_X1 U16060 ( .A1(n13927), .A2(n13926), .ZN(P3_U3479) );
  AOI22_X1 U16061 ( .A1(n14005), .A2(n13928), .B1(n14003), .B2(n13942), .ZN(
        n13932) );
  INV_X1 U16062 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13930) );
  INV_X1 U16063 ( .A(n13929), .ZN(n14006) );
  MUX2_X1 U16064 ( .A(n13930), .B(n14006), .S(n15976), .Z(n13931) );
  NAND2_X1 U16065 ( .A1(n13932), .A2(n13931), .ZN(P3_U3478) );
  NOR2_X1 U16066 ( .A1(n13934), .A2(n13933), .ZN(n13937) );
  AOI21_X1 U16067 ( .B1(n13937), .B2(n13936), .A(n13935), .ZN(n14010) );
  MUX2_X1 U16068 ( .A(n13938), .B(n14010), .S(n15976), .Z(n13939) );
  OAI21_X1 U16069 ( .B1(n14014), .B2(n13940), .A(n13939), .ZN(P3_U3477) );
  INV_X1 U16070 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13941) );
  MUX2_X1 U16071 ( .A(n13941), .B(n14015), .S(n15976), .Z(n13944) );
  NAND2_X1 U16072 ( .A1(n14017), .A2(n13942), .ZN(n13943) );
  OAI211_X1 U16073 ( .C1(n14022), .C2(n13945), .A(n13944), .B(n13943), .ZN(
        P3_U3476) );
  NAND2_X1 U16074 ( .A1(n13946), .A2(n15928), .ZN(n13948) );
  OAI211_X1 U16075 ( .C1(n15948), .C2(n13949), .A(n13948), .B(n13947), .ZN(
        n14023) );
  MUX2_X1 U16076 ( .A(P3_REG1_REG_11__SCAN_IN), .B(n14023), .S(n15976), .Z(
        P3_U3470) );
  OR2_X1 U16077 ( .A1(n13951), .A2(n13950), .ZN(n13952) );
  AND2_X1 U16078 ( .A1(n13953), .A2(n13952), .ZN(n15898) );
  OAI22_X1 U16079 ( .A1(n13955), .A2(n15916), .B1(n15914), .B2(n13954), .ZN(
        n13956) );
  INV_X1 U16080 ( .A(n13956), .ZN(n13963) );
  OAI21_X1 U16081 ( .B1(n13959), .B2(n13958), .A(n13957), .ZN(n13961) );
  NAND2_X1 U16082 ( .A1(n13961), .A2(n13960), .ZN(n13962) );
  OAI211_X1 U16083 ( .C1(n15898), .C2(n13964), .A(n13963), .B(n13962), .ZN(
        n15900) );
  OR2_X1 U16084 ( .A1(n15948), .A2(n13965), .ZN(n15895) );
  OAI21_X1 U16085 ( .B1(n15898), .B2(n15950), .A(n15895), .ZN(n13966) );
  NOR2_X1 U16086 ( .A1(n15900), .A2(n13966), .ZN(n15929) );
  INV_X1 U16087 ( .A(n15929), .ZN(n13967) );
  MUX2_X1 U16088 ( .A(n13967), .B(P3_REG1_REG_2__SCAN_IN), .S(n15973), .Z(
        P3_U3461) );
  NAND2_X1 U16089 ( .A1(n13968), .A2(n14018), .ZN(n13970) );
  NAND2_X1 U16090 ( .A1(n15959), .A2(n13969), .ZN(n13973) );
  OAI211_X1 U16091 ( .C1(n13971), .C2(n15959), .A(n13970), .B(n13973), .ZN(
        P3_U3458) );
  NAND2_X1 U16092 ( .A1(n15960), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n13972) );
  OAI211_X1 U16093 ( .C1(n13974), .C2(n14013), .A(n13973), .B(n13972), .ZN(
        P3_U3457) );
  NAND2_X1 U16094 ( .A1(n13977), .A2(n14018), .ZN(n13978) );
  MUX2_X1 U16095 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n13980), .S(n15959), .Z(
        P3_U3452) );
  MUX2_X1 U16096 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n13981), .S(n15959), .Z(
        P3_U3451) );
  MUX2_X1 U16097 ( .A(n13983), .B(n13982), .S(n15959), .Z(n13986) );
  NAND2_X1 U16098 ( .A1(n13984), .A2(n14018), .ZN(n13985) );
  OAI211_X1 U16099 ( .C1(n13987), .C2(n14021), .A(n13986), .B(n13985), .ZN(
        P3_U3450) );
  INV_X1 U16100 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13989) );
  MUX2_X1 U16101 ( .A(n13989), .B(n13988), .S(n15959), .Z(n13992) );
  NAND2_X1 U16102 ( .A1(n13990), .A2(n14018), .ZN(n13991) );
  OAI211_X1 U16103 ( .C1(n13993), .C2(n14021), .A(n13992), .B(n13991), .ZN(
        P3_U3449) );
  INV_X1 U16104 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13995) );
  MUX2_X1 U16105 ( .A(n13995), .B(n13994), .S(n15959), .Z(n13996) );
  OAI21_X1 U16106 ( .B1(n13997), .B2(n14021), .A(n13996), .ZN(P3_U3448) );
  OAI22_X1 U16107 ( .A1(n13999), .A2(n14021), .B1(n13998), .B2(n14013), .ZN(
        n14002) );
  MUX2_X1 U16108 ( .A(n14000), .B(P3_REG0_REG_20__SCAN_IN), .S(n15960), .Z(
        n14001) );
  OR2_X1 U16109 ( .A1(n14002), .A2(n14001), .ZN(P3_U3447) );
  AOI22_X1 U16110 ( .A1(n14005), .A2(n14004), .B1(n14003), .B2(n14018), .ZN(
        n14009) );
  MUX2_X1 U16111 ( .A(n14007), .B(n14006), .S(n15959), .Z(n14008) );
  NAND2_X1 U16112 ( .A1(n14009), .A2(n14008), .ZN(P3_U3446) );
  INV_X1 U16113 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n14011) );
  MUX2_X1 U16114 ( .A(n14011), .B(n14010), .S(n15959), .Z(n14012) );
  OAI21_X1 U16115 ( .B1(n14014), .B2(n14013), .A(n14012), .ZN(P3_U3444) );
  INV_X1 U16116 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n14016) );
  MUX2_X1 U16117 ( .A(n14016), .B(n14015), .S(n15959), .Z(n14020) );
  NAND2_X1 U16118 ( .A1(n14018), .A2(n14017), .ZN(n14019) );
  OAI211_X1 U16119 ( .C1(n14022), .C2(n14021), .A(n14020), .B(n14019), .ZN(
        P3_U3441) );
  MUX2_X1 U16120 ( .A(P3_REG0_REG_11__SCAN_IN), .B(n14023), .S(n15959), .Z(
        P3_U3423) );
  INV_X1 U16121 ( .A(n14024), .ZN(n14025) );
  MUX2_X1 U16122 ( .A(P3_D_REG_1__SCAN_IN), .B(n14025), .S(n14026), .Z(
        P3_U3377) );
  MUX2_X1 U16123 ( .A(P3_D_REG_0__SCAN_IN), .B(n14027), .S(n14026), .Z(
        P3_U3376) );
  NAND2_X1 U16124 ( .A1(n14029), .A2(n14028), .ZN(n14032) );
  INV_X1 U16125 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n14030) );
  OR4_X1 U16126 ( .A1(n8119), .A2(P3_IR_REG_30__SCAN_IN), .A3(n14030), .A4(
        P3_U3151), .ZN(n14031) );
  OAI211_X1 U16127 ( .C1(n10312), .C2(n14033), .A(n14032), .B(n14031), .ZN(
        P3_U3264) );
  OAI222_X1 U16128 ( .A1(P3_U3151), .A2(n14036), .B1(n14040), .B2(n14035), 
        .C1(n14034), .C2(n14033), .ZN(P3_U3266) );
  INV_X1 U16129 ( .A(n14037), .ZN(n14039) );
  OAI222_X1 U16130 ( .A1(n14033), .A2(n14041), .B1(n14040), .B2(n14039), .C1(
        n14038), .C2(P3_U3151), .ZN(P3_U3267) );
  INV_X1 U16131 ( .A(n14107), .ZN(n14044) );
  NAND2_X1 U16132 ( .A1(n14044), .A2(n14043), .ZN(n14045) );
  NOR2_X1 U16133 ( .A1(n14046), .A2(n14045), .ZN(n14108) );
  AOI21_X1 U16134 ( .B1(n14046), .B2(n14045), .A(n14108), .ZN(n14052) );
  INV_X1 U16135 ( .A(n14047), .ZN(n14517) );
  OAI22_X1 U16136 ( .A1(n14116), .A2(n14204), .B1(n14091), .B2(n14202), .ZN(
        n14513) );
  NAND2_X1 U16137 ( .A1(n14206), .A2(n14513), .ZN(n14048) );
  OAI211_X1 U16138 ( .C1(n14209), .C2(n14517), .A(n14049), .B(n14048), .ZN(
        n14050) );
  AOI21_X1 U16139 ( .B1(n14643), .B2(n14211), .A(n14050), .ZN(n14051) );
  OAI21_X1 U16140 ( .B1(n14052), .B2(n14213), .A(n14051), .ZN(P2_U3187) );
  AND2_X1 U16141 ( .A1(n14164), .A2(n14163), .ZN(n14160) );
  NOR2_X1 U16142 ( .A1(n14160), .A2(n14053), .ZN(n14055) );
  XNOR2_X1 U16143 ( .A(n14055), .B(n14054), .ZN(n14057) );
  AOI21_X1 U16144 ( .B1(n14057), .B2(n14058), .A(n14213), .ZN(n14056) );
  OAI21_X1 U16145 ( .B1(n14058), .B2(n14057), .A(n14056), .ZN(n14063) );
  OAI22_X1 U16146 ( .A1(n7417), .A2(n14204), .B1(n14059), .B2(n14202), .ZN(
        n14380) );
  OAI22_X1 U16147 ( .A1(n14383), .A2(n14209), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14060), .ZN(n14061) );
  AOI21_X1 U16148 ( .B1(n14380), .B2(n14206), .A(n14061), .ZN(n14062) );
  OAI211_X1 U16149 ( .C1(n14375), .C2(n14171), .A(n14063), .B(n14062), .ZN(
        P2_U3188) );
  NAND2_X1 U16150 ( .A1(n14065), .A2(n14064), .ZN(n14069) );
  OR2_X1 U16151 ( .A1(n14182), .A2(n14181), .ZN(n14067) );
  NAND2_X1 U16152 ( .A1(n14067), .A2(n14066), .ZN(n14068) );
  XOR2_X1 U16153 ( .A(n14069), .B(n14068), .Z(n14074) );
  AOI22_X1 U16154 ( .A1(n14226), .A2(n14193), .B1(n14192), .B2(n14228), .ZN(
        n14441) );
  NAND2_X1 U16155 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n14300)
         );
  NAND2_X1 U16156 ( .A1(n14194), .A2(n14445), .ZN(n14071) );
  OAI211_X1 U16157 ( .C1(n14441), .C2(n14196), .A(n14300), .B(n14071), .ZN(
        n14072) );
  AOI21_X1 U16158 ( .B1(n14615), .B2(n14211), .A(n14072), .ZN(n14073) );
  OAI21_X1 U16159 ( .B1(n14074), .B2(n14213), .A(n14073), .ZN(P2_U3191) );
  OR2_X1 U16160 ( .A1(n14182), .A2(n14075), .ZN(n14077) );
  NAND2_X1 U16161 ( .A1(n14077), .A2(n14076), .ZN(n14080) );
  OAI211_X1 U16162 ( .C1(n14080), .C2(n14079), .A(n14078), .B(n14161), .ZN(
        n14086) );
  AOI22_X1 U16163 ( .A1(n14224), .A2(n14193), .B1(n14192), .B2(n14226), .ZN(
        n14413) );
  INV_X1 U16164 ( .A(n14413), .ZN(n14084) );
  INV_X1 U16165 ( .A(n14417), .ZN(n14082) );
  OAI22_X1 U16166 ( .A1(n14082), .A2(n14209), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14081), .ZN(n14083) );
  AOI21_X1 U16167 ( .B1(n14084), .B2(n14206), .A(n14083), .ZN(n14085) );
  OAI211_X1 U16168 ( .C1(n14420), .C2(n14171), .A(n14086), .B(n14085), .ZN(
        P2_U3195) );
  INV_X1 U16169 ( .A(n14087), .ZN(n14088) );
  AOI21_X1 U16170 ( .B1(n14090), .B2(n14089), .A(n14088), .ZN(n14097) );
  OAI22_X1 U16171 ( .A1(n14092), .A2(n14202), .B1(n14091), .B2(n14204), .ZN(
        n14554) );
  NAND2_X1 U16172 ( .A1(n14206), .A2(n14554), .ZN(n14093) );
  OAI211_X1 U16173 ( .C1(n14209), .C2(n14559), .A(n14094), .B(n14093), .ZN(
        n14095) );
  AOI21_X1 U16174 ( .B1(n14653), .B2(n14211), .A(n14095), .ZN(n14096) );
  OAI21_X1 U16175 ( .B1(n14097), .B2(n14213), .A(n14096), .ZN(P2_U3196) );
  OAI211_X1 U16176 ( .C1(n14100), .C2(n14099), .A(n14098), .B(n14161), .ZN(
        n14106) );
  OAI22_X1 U16177 ( .A1(n14101), .A2(n14204), .B1(n7417), .B2(n14202), .ZN(
        n14338) );
  INV_X1 U16178 ( .A(n14343), .ZN(n14103) );
  OAI22_X1 U16179 ( .A1(n14103), .A2(n14209), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14102), .ZN(n14104) );
  AOI21_X1 U16180 ( .B1(n14338), .B2(n14206), .A(n14104), .ZN(n14105) );
  OAI211_X1 U16181 ( .C1(n14346), .C2(n14171), .A(n14106), .B(n14105), .ZN(
        P2_U3197) );
  NOR2_X1 U16182 ( .A1(n14108), .A2(n14107), .ZN(n14111) );
  XNOR2_X1 U16183 ( .A(n14111), .B(n14109), .ZN(n14201) );
  AOI22_X1 U16184 ( .A1(n14201), .A2(n14200), .B1(n14111), .B2(n14110), .ZN(
        n14115) );
  NAND2_X1 U16185 ( .A1(n14113), .A2(n14112), .ZN(n14114) );
  XNOR2_X1 U16186 ( .A(n14115), .B(n14114), .ZN(n14121) );
  OAI22_X1 U16187 ( .A1(n14183), .A2(n14204), .B1(n14116), .B2(n14202), .ZN(
        n14484) );
  NAND2_X1 U16188 ( .A1(n14484), .A2(n14206), .ZN(n14117) );
  OAI211_X1 U16189 ( .C1(n14209), .C2(n14490), .A(n14118), .B(n14117), .ZN(
        n14119) );
  AOI21_X1 U16190 ( .B1(n14631), .B2(n14211), .A(n14119), .ZN(n14120) );
  OAI21_X1 U16191 ( .B1(n14121), .B2(n14213), .A(n14120), .ZN(P2_U3198) );
  OAI21_X1 U16192 ( .B1(n14124), .B2(n14123), .A(n14122), .ZN(n14125) );
  NAND2_X1 U16193 ( .A1(n14125), .A2(n14161), .ZN(n14129) );
  INV_X1 U16194 ( .A(n14205), .ZN(n14230) );
  AOI22_X1 U16195 ( .A1(n14228), .A2(n14193), .B1(n14192), .B2(n14230), .ZN(
        n14478) );
  OAI21_X1 U16196 ( .B1(n14478), .B2(n14196), .A(n14126), .ZN(n14127) );
  AOI21_X1 U16197 ( .B1(n14468), .B2(n14194), .A(n14127), .ZN(n14128) );
  OAI211_X1 U16198 ( .C1(n7918), .C2(n14171), .A(n14129), .B(n14128), .ZN(
        P2_U3200) );
  OAI211_X1 U16199 ( .C1(n14132), .C2(n14131), .A(n14130), .B(n14161), .ZN(
        n14137) );
  AOI22_X1 U16200 ( .A1(n14221), .A2(n14193), .B1(n14192), .B2(n14223), .ZN(
        n14351) );
  NOR2_X1 U16201 ( .A1(n14351), .A2(n14196), .ZN(n14135) );
  OAI22_X1 U16202 ( .A1(n14357), .A2(n14209), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14133), .ZN(n14134) );
  AOI211_X1 U16203 ( .C1(n14590), .C2(n14211), .A(n14135), .B(n14134), .ZN(
        n14136) );
  NAND2_X1 U16204 ( .A1(n14137), .A2(n14136), .ZN(P2_U3201) );
  OR2_X1 U16205 ( .A1(n14182), .A2(n14138), .ZN(n14141) );
  NAND2_X1 U16206 ( .A1(n14141), .A2(n14139), .ZN(n14143) );
  AND2_X1 U16207 ( .A1(n14141), .A2(n14140), .ZN(n14142) );
  AOI21_X1 U16208 ( .B1(n14144), .B2(n14143), .A(n14142), .ZN(n14149) );
  AOI22_X1 U16209 ( .A1(n14225), .A2(n14193), .B1(n14192), .B2(n14227), .ZN(
        n14426) );
  INV_X1 U16210 ( .A(n14432), .ZN(n14145) );
  AOI22_X1 U16211 ( .A1(n14145), .A2(n14194), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14146) );
  OAI21_X1 U16212 ( .B1(n14426), .B2(n14196), .A(n14146), .ZN(n14147) );
  AOI21_X1 U16213 ( .B1(n14610), .B2(n14211), .A(n14147), .ZN(n14148) );
  OAI21_X1 U16214 ( .B1(n14149), .B2(n14213), .A(n14148), .ZN(P2_U3205) );
  XNOR2_X1 U16215 ( .A(n14151), .B(n14150), .ZN(n14159) );
  OR2_X1 U16216 ( .A1(n14152), .A2(n14202), .ZN(n14154) );
  OR2_X1 U16217 ( .A1(n14203), .A2(n14204), .ZN(n14153) );
  NAND2_X1 U16218 ( .A1(n14154), .A2(n14153), .ZN(n14532) );
  NAND2_X1 U16219 ( .A1(n14206), .A2(n14532), .ZN(n14155) );
  OAI211_X1 U16220 ( .C1(n14209), .C2(n14538), .A(n14156), .B(n14155), .ZN(
        n14157) );
  AOI21_X1 U16221 ( .B1(n14648), .B2(n14211), .A(n14157), .ZN(n14158) );
  OAI21_X1 U16222 ( .B1(n14159), .B2(n14213), .A(n14158), .ZN(P2_U3206) );
  INV_X1 U16223 ( .A(n14160), .ZN(n14162) );
  OAI211_X1 U16224 ( .C1(n14164), .C2(n14163), .A(n14162), .B(n14161), .ZN(
        n14170) );
  OAI22_X1 U16225 ( .A1(n14166), .A2(n14204), .B1(n14165), .B2(n14202), .ZN(
        n14388) );
  OAI22_X1 U16226 ( .A1(n14401), .A2(n14209), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14167), .ZN(n14168) );
  AOI21_X1 U16227 ( .B1(n14388), .B2(n14206), .A(n14168), .ZN(n14169) );
  OAI211_X1 U16228 ( .C1(n14403), .C2(n14171), .A(n14170), .B(n14169), .ZN(
        P2_U3207) );
  XNOR2_X1 U16229 ( .A(n14173), .B(n14172), .ZN(n14180) );
  AOI21_X1 U16230 ( .B1(n14206), .B2(n14175), .A(n14174), .ZN(n14176) );
  OAI21_X1 U16231 ( .B1(n14209), .B2(n14177), .A(n14176), .ZN(n14178) );
  AOI21_X1 U16232 ( .B1(n14658), .B2(n14211), .A(n14178), .ZN(n14179) );
  OAI21_X1 U16233 ( .B1(n14180), .B2(n14213), .A(n14179), .ZN(P2_U3208) );
  XNOR2_X1 U16234 ( .A(n14182), .B(n14181), .ZN(n14189) );
  OAI22_X1 U16235 ( .A1(n14184), .A2(n14204), .B1(n14183), .B2(n14202), .ZN(
        n14451) );
  NAND2_X1 U16236 ( .A1(n14451), .A2(n14206), .ZN(n14186) );
  OAI211_X1 U16237 ( .C1(n14209), .C2(n14456), .A(n14186), .B(n14185), .ZN(
        n14187) );
  AOI21_X1 U16238 ( .B1(n14620), .B2(n14211), .A(n14187), .ZN(n14188) );
  OAI21_X1 U16239 ( .B1(n14189), .B2(n14213), .A(n14188), .ZN(P2_U3210) );
  AOI22_X1 U16240 ( .A1(n14219), .A2(n14193), .B1(n14192), .B2(n14221), .ZN(
        n14321) );
  AOI22_X1 U16241 ( .A1(n14326), .A2(n14194), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14195) );
  OAI21_X1 U16242 ( .B1(n14321), .B2(n14196), .A(n14195), .ZN(n14197) );
  AOI21_X1 U16243 ( .B1(n14327), .B2(n14211), .A(n14197), .ZN(n14198) );
  OAI21_X1 U16244 ( .B1(n14199), .B2(n14213), .A(n14198), .ZN(P2_U3212) );
  XNOR2_X1 U16245 ( .A(n14201), .B(n14200), .ZN(n14214) );
  OAI22_X1 U16246 ( .A1(n14205), .A2(n14204), .B1(n14203), .B2(n14202), .ZN(
        n14503) );
  NAND2_X1 U16247 ( .A1(n14206), .A2(n14503), .ZN(n14207) );
  OAI211_X1 U16248 ( .C1(n14209), .C2(n14507), .A(n14208), .B(n14207), .ZN(
        n14210) );
  AOI21_X1 U16249 ( .B1(n14500), .B2(n14211), .A(n14210), .ZN(n14212) );
  OAI21_X1 U16250 ( .B1(n14214), .B2(n14213), .A(n14212), .ZN(P2_U3213) );
  MUX2_X1 U16251 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n14215), .S(P2_U3947), .Z(
        P2_U3562) );
  MUX2_X1 U16252 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n14216), .S(P2_U3947), .Z(
        P2_U3561) );
  MUX2_X1 U16253 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n14217), .S(P2_U3947), .Z(
        P2_U3560) );
  MUX2_X1 U16254 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n14218), .S(P2_U3947), .Z(
        P2_U3559) );
  MUX2_X1 U16255 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n14219), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U16256 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n14220), .S(P2_U3947), .Z(
        P2_U3557) );
  MUX2_X1 U16257 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n14221), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U16258 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n14222), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U16259 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n14223), .S(P2_U3947), .Z(
        P2_U3554) );
  MUX2_X1 U16260 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n14224), .S(P2_U3947), .Z(
        P2_U3553) );
  MUX2_X1 U16261 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n14225), .S(P2_U3947), .Z(
        P2_U3552) );
  MUX2_X1 U16262 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n14226), .S(P2_U3947), .Z(
        P2_U3551) );
  MUX2_X1 U16263 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n14227), .S(P2_U3947), .Z(
        P2_U3550) );
  MUX2_X1 U16264 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n14228), .S(P2_U3947), .Z(
        P2_U3549) );
  MUX2_X1 U16265 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n14229), .S(P2_U3947), .Z(
        P2_U3548) );
  MUX2_X1 U16266 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n14230), .S(P2_U3947), .Z(
        P2_U3547) );
  MUX2_X1 U16267 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n14231), .S(P2_U3947), .Z(
        P2_U3546) );
  MUX2_X1 U16268 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n14232), .S(P2_U3947), .Z(
        P2_U3545) );
  MUX2_X1 U16269 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n9355), .S(P2_U3947), .Z(
        P2_U3544) );
  MUX2_X1 U16270 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n7107), .S(P2_U3947), .Z(
        P2_U3543) );
  MUX2_X1 U16271 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n14233), .S(P2_U3947), .Z(
        P2_U3542) );
  MUX2_X1 U16272 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n14234), .S(P2_U3947), .Z(
        P2_U3541) );
  MUX2_X1 U16273 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n14235), .S(P2_U3947), .Z(
        P2_U3540) );
  MUX2_X1 U16274 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n14236), .S(P2_U3947), .Z(
        P2_U3539) );
  MUX2_X1 U16275 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n14237), .S(P2_U3947), .Z(
        P2_U3538) );
  MUX2_X1 U16276 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n14238), .S(P2_U3947), .Z(
        P2_U3537) );
  MUX2_X1 U16277 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n14239), .S(P2_U3947), .Z(
        P2_U3536) );
  MUX2_X1 U16278 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n14240), .S(P2_U3947), .Z(
        P2_U3535) );
  MUX2_X1 U16279 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n14241), .S(P2_U3947), .Z(
        P2_U3534) );
  MUX2_X1 U16280 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n14242), .S(P2_U3947), .Z(
        P2_U3533) );
  MUX2_X1 U16281 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n12775), .S(P2_U3947), .Z(
        P2_U3532) );
  MUX2_X1 U16282 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n14243), .S(P2_U3947), .Z(
        P2_U3531) );
  AOI211_X1 U16283 ( .C1(n14246), .C2(n14245), .A(n14244), .B(n15825), .ZN(
        n14247) );
  INV_X1 U16284 ( .A(n14247), .ZN(n14257) );
  OAI22_X1 U16285 ( .A1(n15806), .A2(n14250), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14248), .ZN(n14249) );
  AOI21_X1 U16286 ( .B1(P2_ADDR_REG_1__SCAN_IN), .B2(n15809), .A(n14249), .ZN(
        n14256) );
  MUX2_X1 U16287 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n10641), .S(n14250), .Z(
        n14251) );
  OAI21_X1 U16288 ( .B1(n10747), .B2(n14252), .A(n14251), .ZN(n14253) );
  NAND3_X1 U16289 ( .A1(n15811), .A2(n14254), .A3(n14253), .ZN(n14255) );
  NAND3_X1 U16290 ( .A1(n14257), .A2(n14256), .A3(n14255), .ZN(P2_U3215) );
  AOI211_X1 U16291 ( .C1(n14259), .C2(n14258), .A(n14276), .B(n15825), .ZN(
        n14260) );
  INV_X1 U16292 ( .A(n14260), .ZN(n14268) );
  OAI22_X1 U16293 ( .A1(n15806), .A2(n14262), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14261), .ZN(n14263) );
  AOI21_X1 U16294 ( .B1(n15809), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n14263), .ZN(
        n14267) );
  OAI211_X1 U16295 ( .C1(n14265), .C2(n14264), .A(n15811), .B(n14281), .ZN(
        n14266) );
  NAND3_X1 U16296 ( .A1(n14268), .A2(n14267), .A3(n14266), .ZN(P2_U3216) );
  OAI21_X1 U16297 ( .B1(n15806), .B2(n14277), .A(n14269), .ZN(n14270) );
  AOI21_X1 U16298 ( .B1(n15809), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n14270), .ZN(
        n14286) );
  MUX2_X1 U16299 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n8828), .S(n14277), .Z(
        n14273) );
  INV_X1 U16300 ( .A(n14271), .ZN(n14272) );
  NAND2_X1 U16301 ( .A1(n14273), .A2(n14272), .ZN(n14275) );
  OAI211_X1 U16302 ( .C1(n14276), .C2(n14275), .A(n15815), .B(n14274), .ZN(
        n14285) );
  MUX2_X1 U16303 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n14278), .S(n14277), .Z(
        n14279) );
  NAND3_X1 U16304 ( .A1(n14281), .A2(n14280), .A3(n14279), .ZN(n14282) );
  NAND3_X1 U16305 ( .A1(n15811), .A2(n14283), .A3(n14282), .ZN(n14284) );
  NAND3_X1 U16306 ( .A1(n14286), .A2(n14285), .A3(n14284), .ZN(P2_U3217) );
  INV_X1 U16307 ( .A(n14287), .ZN(n14288) );
  XNOR2_X1 U16308 ( .A(n14291), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n14296) );
  NAND2_X1 U16309 ( .A1(n14293), .A2(n14292), .ZN(n14295) );
  OAI21_X1 U16310 ( .B1(n14296), .B2(n15825), .A(n15806), .ZN(n14297) );
  OAI211_X1 U16311 ( .C1(n14302), .C2(n15840), .A(n14301), .B(n14300), .ZN(
        P2_U3233) );
  XNOR2_X1 U16312 ( .A(n14304), .B(n14303), .ZN(n14306) );
  AOI21_X1 U16313 ( .B1(n14306), .B2(n14556), .A(n14305), .ZN(n14578) );
  OAI21_X1 U16314 ( .B1(n14323), .B2(n14307), .A(n10836), .ZN(n14308) );
  NOR2_X1 U16315 ( .A1(n14308), .A2(n10014), .ZN(n14575) );
  INV_X1 U16316 ( .A(n14575), .ZN(n14315) );
  NAND3_X1 U16317 ( .A1(n14574), .A2(n14573), .A3(n14461), .ZN(n14314) );
  OAI22_X1 U16318 ( .A1(n14311), .A2(n15843), .B1(n14310), .B2(n15850), .ZN(
        n14312) );
  AOI21_X1 U16319 ( .B1(n14576), .B2(n14541), .A(n14312), .ZN(n14313) );
  OAI211_X1 U16320 ( .C1(n14315), .C2(n14330), .A(n14314), .B(n14313), .ZN(
        n14316) );
  INV_X1 U16321 ( .A(n14316), .ZN(n14317) );
  OAI21_X1 U16322 ( .B1(n14499), .B2(n14578), .A(n14317), .ZN(P2_U3238) );
  XOR2_X1 U16323 ( .A(n14319), .B(n14318), .Z(n14685) );
  INV_X1 U16324 ( .A(n14321), .ZN(n14322) );
  INV_X1 U16325 ( .A(n14581), .ZN(n14332) );
  INV_X1 U16326 ( .A(n14323), .ZN(n14325) );
  AOI21_X1 U16327 ( .B1(n14341), .B2(n14327), .A(n14635), .ZN(n14324) );
  NAND2_X1 U16328 ( .A1(n14325), .A2(n14324), .ZN(n14580) );
  AOI22_X1 U16329 ( .A1(n14326), .A2(n14560), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14499), .ZN(n14329) );
  NAND2_X1 U16330 ( .A1(n14327), .A2(n14541), .ZN(n14328) );
  OAI211_X1 U16331 ( .C1(n14580), .C2(n14330), .A(n14329), .B(n14328), .ZN(
        n14331) );
  AOI21_X1 U16332 ( .B1(n14332), .B2(n15850), .A(n14331), .ZN(n14333) );
  OAI21_X1 U16333 ( .B1(n14685), .B2(n14546), .A(n14333), .ZN(P2_U3239) );
  XOR2_X1 U16334 ( .A(n14334), .B(n14337), .Z(n14689) );
  OAI21_X1 U16335 ( .B1(n14337), .B2(n14336), .A(n14335), .ZN(n14339) );
  AOI21_X1 U16336 ( .B1(n14339), .B2(n14556), .A(n14338), .ZN(n14340) );
  INV_X1 U16337 ( .A(n14340), .ZN(n14583) );
  INV_X1 U16338 ( .A(n14341), .ZN(n14342) );
  AOI211_X1 U16339 ( .C1(n14585), .C2(n14359), .A(n14342), .B(n14635), .ZN(
        n14584) );
  NAND2_X1 U16340 ( .A1(n14584), .A2(n14567), .ZN(n14345) );
  AOI22_X1 U16341 ( .A1(n14343), .A2(n14560), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n14499), .ZN(n14344) );
  OAI211_X1 U16342 ( .C1(n14346), .C2(n14563), .A(n14345), .B(n14344), .ZN(
        n14347) );
  AOI21_X1 U16343 ( .B1(n14583), .B2(n15850), .A(n14347), .ZN(n14348) );
  OAI21_X1 U16344 ( .B1(n14689), .B2(n14546), .A(n14348), .ZN(P2_U3240) );
  XNOR2_X1 U16345 ( .A(n14350), .B(n14349), .ZN(n14352) );
  OAI21_X1 U16346 ( .B1(n14352), .B2(n14534), .A(n14351), .ZN(n14588) );
  OAI21_X1 U16347 ( .B1(n14355), .B2(n14354), .A(n14353), .ZN(n14693) );
  INV_X1 U16348 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n14356) );
  OAI22_X1 U16349 ( .A1(n14357), .A2(n15843), .B1(n14356), .B2(n15850), .ZN(
        n14358) );
  AOI21_X1 U16350 ( .B1(n14590), .B2(n14541), .A(n14358), .ZN(n14362) );
  AOI21_X1 U16351 ( .B1(n14371), .B2(n14590), .A(n14635), .ZN(n14360) );
  AND2_X1 U16352 ( .A1(n14360), .A2(n14359), .ZN(n14589) );
  NAND2_X1 U16353 ( .A1(n14589), .A2(n14567), .ZN(n14361) );
  OAI211_X1 U16354 ( .C1(n14693), .C2(n14546), .A(n14362), .B(n14361), .ZN(
        n14363) );
  AOI21_X1 U16355 ( .B1(n15850), .B2(n14588), .A(n14363), .ZN(n14364) );
  INV_X1 U16356 ( .A(n14364), .ZN(P2_U3241) );
  NAND2_X1 U16357 ( .A1(n14396), .A2(n14365), .ZN(n14368) );
  INV_X1 U16358 ( .A(n14366), .ZN(n14367) );
  AOI21_X1 U16359 ( .B1(n14369), .B2(n14368), .A(n14367), .ZN(n14697) );
  INV_X1 U16360 ( .A(n14370), .ZN(n14373) );
  INV_X1 U16361 ( .A(n14371), .ZN(n14372) );
  AOI211_X1 U16362 ( .C1(n14595), .C2(n14373), .A(n14635), .B(n14372), .ZN(
        n14594) );
  OAI22_X1 U16363 ( .A1(n14375), .A2(n14563), .B1(n15850), .B2(n14374), .ZN(
        n14376) );
  AOI21_X1 U16364 ( .B1(n14594), .B2(n14567), .A(n14376), .ZN(n14386) );
  AOI21_X1 U16365 ( .B1(n14379), .B2(n14378), .A(n14377), .ZN(n14382) );
  INV_X1 U16366 ( .A(n14380), .ZN(n14381) );
  OAI21_X1 U16367 ( .B1(n14382), .B2(n14534), .A(n14381), .ZN(n14593) );
  NOR2_X1 U16368 ( .A1(n14383), .A2(n15843), .ZN(n14384) );
  OAI21_X1 U16369 ( .B1(n14593), .B2(n14384), .A(n15850), .ZN(n14385) );
  OAI211_X1 U16370 ( .C1(n14697), .C2(n14546), .A(n14386), .B(n14385), .ZN(
        P2_U3242) );
  XNOR2_X1 U16371 ( .A(n14387), .B(n14398), .ZN(n14390) );
  INV_X1 U16372 ( .A(n14388), .ZN(n14389) );
  OAI21_X1 U16373 ( .B1(n14390), .B2(n14534), .A(n14389), .ZN(n14598) );
  NAND2_X1 U16374 ( .A1(n14391), .A2(n14392), .ZN(n14394) );
  NAND2_X1 U16375 ( .A1(n14394), .A2(n14393), .ZN(n14399) );
  AND2_X1 U16376 ( .A1(n14396), .A2(n14395), .ZN(n14397) );
  OAI21_X1 U16377 ( .B1(n14399), .B2(n14398), .A(n14397), .ZN(n14701) );
  OAI22_X1 U16378 ( .A1(n14401), .A2(n15843), .B1(n14400), .B2(n15850), .ZN(
        n14402) );
  AOI21_X1 U16379 ( .B1(n14600), .B2(n14541), .A(n14402), .ZN(n14406) );
  OAI21_X1 U16380 ( .B1(n6575), .B2(n14403), .A(n10836), .ZN(n14404) );
  NOR2_X1 U16381 ( .A1(n14404), .A2(n14370), .ZN(n14599) );
  NAND2_X1 U16382 ( .A1(n14599), .A2(n14567), .ZN(n14405) );
  OAI211_X1 U16383 ( .C1(n14701), .C2(n14546), .A(n14406), .B(n14405), .ZN(
        n14407) );
  AOI21_X1 U16384 ( .B1(n15850), .B2(n14598), .A(n14407), .ZN(n14408) );
  INV_X1 U16385 ( .A(n14408), .ZN(P2_U3243) );
  NAND2_X1 U16386 ( .A1(n14391), .A2(n14409), .ZN(n14410) );
  XOR2_X1 U16387 ( .A(n14411), .B(n14410), .Z(n14705) );
  XOR2_X1 U16388 ( .A(n14412), .B(n14411), .Z(n14414) );
  OAI21_X1 U16389 ( .B1(n14414), .B2(n14534), .A(n14413), .ZN(n14603) );
  NAND2_X1 U16390 ( .A1(n14429), .A2(n14605), .ZN(n14415) );
  NAND2_X1 U16391 ( .A1(n14415), .A2(n10836), .ZN(n14416) );
  NOR2_X1 U16392 ( .A1(n6575), .A2(n14416), .ZN(n14604) );
  NAND2_X1 U16393 ( .A1(n14604), .A2(n14567), .ZN(n14419) );
  AOI22_X1 U16394 ( .A1(n14417), .A2(n14560), .B1(P2_REG2_REG_21__SCAN_IN), 
        .B2(n14499), .ZN(n14418) );
  OAI211_X1 U16395 ( .C1(n14420), .C2(n14563), .A(n14419), .B(n14418), .ZN(
        n14421) );
  AOI21_X1 U16396 ( .B1(n14603), .B2(n15850), .A(n14421), .ZN(n14422) );
  OAI21_X1 U16397 ( .B1(n14705), .B2(n14546), .A(n14422), .ZN(P2_U3244) );
  XNOR2_X1 U16398 ( .A(n14423), .B(n14424), .ZN(n14709) );
  XOR2_X1 U16399 ( .A(n14425), .B(n14424), .Z(n14427) );
  OAI21_X1 U16400 ( .B1(n14427), .B2(n14534), .A(n14426), .ZN(n14608) );
  AOI21_X1 U16401 ( .B1(n14428), .B2(n14610), .A(n14635), .ZN(n14430) );
  AND2_X1 U16402 ( .A1(n14430), .A2(n14429), .ZN(n14609) );
  NAND2_X1 U16403 ( .A1(n14609), .A2(n14567), .ZN(n14435) );
  OAI22_X1 U16404 ( .A1(n14432), .A2(n15843), .B1(n15850), .B2(n14431), .ZN(
        n14433) );
  AOI21_X1 U16405 ( .B1(n14610), .B2(n14541), .A(n14433), .ZN(n14434) );
  NAND2_X1 U16406 ( .A1(n14435), .A2(n14434), .ZN(n14436) );
  AOI21_X1 U16407 ( .B1(n14608), .B2(n15850), .A(n14436), .ZN(n14437) );
  OAI21_X1 U16408 ( .B1(n14709), .B2(n14546), .A(n14437), .ZN(P2_U3245) );
  XNOR2_X1 U16409 ( .A(n14438), .B(n14439), .ZN(n14713) );
  XOR2_X1 U16410 ( .A(n14440), .B(n14439), .Z(n14442) );
  OAI21_X1 U16411 ( .B1(n14442), .B2(n14534), .A(n14441), .ZN(n14613) );
  INV_X1 U16412 ( .A(n14455), .ZN(n14444) );
  INV_X1 U16413 ( .A(n14428), .ZN(n14443) );
  NAND2_X1 U16414 ( .A1(n14614), .A2(n14567), .ZN(n14447) );
  AOI22_X1 U16415 ( .A1(n14499), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n14445), 
        .B2(n14560), .ZN(n14446) );
  OAI211_X1 U16416 ( .C1(n7128), .C2(n14563), .A(n14447), .B(n14446), .ZN(
        n14448) );
  AOI21_X1 U16417 ( .B1(n14613), .B2(n15850), .A(n14448), .ZN(n14449) );
  OAI21_X1 U16418 ( .B1(n14713), .B2(n14546), .A(n14449), .ZN(P2_U3246) );
  XNOR2_X1 U16419 ( .A(n14450), .B(n14454), .ZN(n14452) );
  AOI21_X1 U16420 ( .B1(n14452), .B2(n14556), .A(n14451), .ZN(n14622) );
  OAI21_X1 U16421 ( .B1(n6717), .B2(n14454), .A(n14453), .ZN(n14618) );
  AOI211_X1 U16422 ( .C1(n14620), .C2(n7920), .A(n14635), .B(n14455), .ZN(
        n14619) );
  NAND2_X1 U16423 ( .A1(n14619), .A2(n14567), .ZN(n14459) );
  INV_X1 U16424 ( .A(n14456), .ZN(n14457) );
  AOI22_X1 U16425 ( .A1(n14499), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14457), 
        .B2(n14560), .ZN(n14458) );
  OAI211_X1 U16426 ( .C1(n9360), .C2(n14563), .A(n14459), .B(n14458), .ZN(
        n14460) );
  AOI21_X1 U16427 ( .B1(n14618), .B2(n14461), .A(n14460), .ZN(n14462) );
  OAI21_X1 U16428 ( .B1(n14499), .B2(n14622), .A(n14462), .ZN(P2_U3247) );
  OAI21_X1 U16429 ( .B1(n14476), .B2(n14464), .A(n14463), .ZN(n14718) );
  NAND2_X1 U16430 ( .A1(n8097), .A2(n14626), .ZN(n14465) );
  NAND2_X1 U16431 ( .A1(n14465), .A2(n10836), .ZN(n14466) );
  NOR2_X1 U16432 ( .A1(n14467), .A2(n14466), .ZN(n14625) );
  NAND2_X1 U16433 ( .A1(n14626), .A2(n14541), .ZN(n14470) );
  NAND2_X1 U16434 ( .A1(n14468), .A2(n14560), .ZN(n14469) );
  OAI211_X1 U16435 ( .C1(n15850), .C2(n14471), .A(n14470), .B(n14469), .ZN(
        n14472) );
  AOI21_X1 U16436 ( .B1(n14625), .B2(n14567), .A(n14472), .ZN(n14482) );
  INV_X1 U16437 ( .A(n14473), .ZN(n14474) );
  NOR2_X1 U16438 ( .A1(n14475), .A2(n14474), .ZN(n14480) );
  OAI21_X1 U16439 ( .B1(n14477), .B2(n6960), .A(n14556), .ZN(n14479) );
  OAI21_X1 U16440 ( .B1(n14480), .B2(n14479), .A(n14478), .ZN(n14624) );
  NAND2_X1 U16441 ( .A1(n14624), .A2(n15850), .ZN(n14481) );
  OAI211_X1 U16442 ( .C1(n14718), .C2(n14546), .A(n14482), .B(n14481), .ZN(
        P2_U3248) );
  XNOR2_X1 U16443 ( .A(n14483), .B(n14488), .ZN(n14486) );
  INV_X1 U16444 ( .A(n14484), .ZN(n14485) );
  OAI21_X1 U16445 ( .B1(n14486), .B2(n14534), .A(n14485), .ZN(n14629) );
  OAI21_X1 U16446 ( .B1(n14489), .B2(n14488), .A(n14487), .ZN(n14722) );
  OAI22_X1 U16447 ( .A1(n15850), .A2(n14491), .B1(n14490), .B2(n15843), .ZN(
        n14492) );
  AOI21_X1 U16448 ( .B1(n14631), .B2(n14541), .A(n14492), .ZN(n14495) );
  AOI21_X1 U16449 ( .B1(n14506), .B2(n14631), .A(n14635), .ZN(n14493) );
  AND2_X1 U16450 ( .A1(n14493), .A2(n8097), .ZN(n14630) );
  NAND2_X1 U16451 ( .A1(n14630), .A2(n14567), .ZN(n14494) );
  OAI211_X1 U16452 ( .C1(n14722), .C2(n14546), .A(n14495), .B(n14494), .ZN(
        n14496) );
  AOI21_X1 U16453 ( .B1(n15850), .B2(n14629), .A(n14496), .ZN(n14497) );
  INV_X1 U16454 ( .A(n14497), .ZN(P2_U3249) );
  XOR2_X1 U16455 ( .A(n14498), .B(n14501), .Z(n14726) );
  AOI22_X1 U16456 ( .A1(n14500), .A2(n14541), .B1(n14499), .B2(
        P2_REG2_REG_15__SCAN_IN), .ZN(n14511) );
  XNOR2_X1 U16457 ( .A(n14502), .B(n14501), .ZN(n14505) );
  INV_X1 U16458 ( .A(n14503), .ZN(n14504) );
  OAI21_X1 U16459 ( .B1(n14505), .B2(n14534), .A(n14504), .ZN(n14638) );
  OAI21_X1 U16460 ( .B1(n14522), .B2(n14634), .A(n14506), .ZN(n14636) );
  OAI22_X1 U16461 ( .A1(n14636), .A2(n14508), .B1(n14507), .B2(n15843), .ZN(
        n14509) );
  OAI21_X1 U16462 ( .B1(n14638), .B2(n14509), .A(n15850), .ZN(n14510) );
  OAI211_X1 U16463 ( .C1(n14726), .C2(n14546), .A(n14511), .B(n14510), .ZN(
        P2_U3250) );
  XOR2_X1 U16464 ( .A(n14516), .B(n14512), .Z(n14515) );
  INV_X1 U16465 ( .A(n14513), .ZN(n14514) );
  OAI21_X1 U16466 ( .B1(n14515), .B2(n14534), .A(n14514), .ZN(n14641) );
  XOR2_X1 U16467 ( .A(n14516), .B(n6769), .Z(n14730) );
  OAI22_X1 U16468 ( .A1(n15850), .A2(n14518), .B1(n14517), .B2(n15843), .ZN(
        n14519) );
  AOI21_X1 U16469 ( .B1(n14643), .B2(n14541), .A(n14519), .ZN(n14524) );
  NAND2_X1 U16470 ( .A1(n14543), .A2(n14643), .ZN(n14520) );
  NAND2_X1 U16471 ( .A1(n14520), .A2(n10836), .ZN(n14521) );
  NOR2_X1 U16472 ( .A1(n14522), .A2(n14521), .ZN(n14642) );
  NAND2_X1 U16473 ( .A1(n14642), .A2(n14567), .ZN(n14523) );
  OAI211_X1 U16474 ( .C1(n14730), .C2(n14546), .A(n14524), .B(n14523), .ZN(
        n14525) );
  AOI21_X1 U16475 ( .B1(n15850), .B2(n14641), .A(n14525), .ZN(n14526) );
  INV_X1 U16476 ( .A(n14526), .ZN(P2_U3251) );
  NAND2_X1 U16477 ( .A1(n12158), .A2(n14527), .ZN(n14549) );
  NAND2_X1 U16478 ( .A1(n14549), .A2(n14528), .ZN(n14530) );
  NAND2_X1 U16479 ( .A1(n14530), .A2(n14529), .ZN(n14531) );
  XOR2_X1 U16480 ( .A(n14536), .B(n14531), .Z(n14535) );
  INV_X1 U16481 ( .A(n14532), .ZN(n14533) );
  OAI21_X1 U16482 ( .B1(n14535), .B2(n14534), .A(n14533), .ZN(n14646) );
  XNOR2_X1 U16483 ( .A(n14537), .B(n14536), .ZN(n14735) );
  OAI22_X1 U16484 ( .A1(n15850), .A2(n14539), .B1(n14538), .B2(n15843), .ZN(
        n14540) );
  AOI21_X1 U16485 ( .B1(n14648), .B2(n14541), .A(n14540), .ZN(n14545) );
  AOI21_X1 U16486 ( .B1(n14557), .B2(n14648), .A(n14635), .ZN(n14542) );
  AND2_X1 U16487 ( .A1(n14543), .A2(n14542), .ZN(n14647) );
  NAND2_X1 U16488 ( .A1(n14647), .A2(n14567), .ZN(n14544) );
  OAI211_X1 U16489 ( .C1(n14735), .C2(n14546), .A(n14545), .B(n14544), .ZN(
        n14547) );
  AOI21_X1 U16490 ( .B1(n15850), .B2(n14646), .A(n14547), .ZN(n14548) );
  INV_X1 U16491 ( .A(n14548), .ZN(P2_U3252) );
  XNOR2_X1 U16492 ( .A(n14549), .B(n14550), .ZN(n14555) );
  XNOR2_X1 U16493 ( .A(n14551), .B(n14550), .ZN(n14656) );
  NOR2_X1 U16494 ( .A1(n14656), .A2(n14552), .ZN(n14553) );
  AOI211_X1 U16495 ( .C1(n14556), .C2(n14555), .A(n14554), .B(n14553), .ZN(
        n14655) );
  AOI211_X1 U16496 ( .C1(n14653), .C2(n14558), .A(n14635), .B(n6791), .ZN(
        n14652) );
  INV_X1 U16497 ( .A(n14559), .ZN(n14561) );
  AOI22_X1 U16498 ( .A1(n14499), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n14561), 
        .B2(n14560), .ZN(n14562) );
  OAI21_X1 U16499 ( .B1(n7108), .B2(n14563), .A(n14562), .ZN(n14566) );
  NOR2_X1 U16500 ( .A1(n14656), .A2(n14564), .ZN(n14565) );
  AOI211_X1 U16501 ( .C1(n14652), .C2(n14567), .A(n14566), .B(n14565), .ZN(
        n14568) );
  OAI21_X1 U16502 ( .B1(n14655), .B2(n14499), .A(n14568), .ZN(P2_U3253) );
  OAI211_X1 U16503 ( .C1(n15879), .C2(n14570), .A(n14569), .B(n14571), .ZN(
        n14680) );
  MUX2_X1 U16504 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n14680), .S(n15893), .Z(
        P2_U3530) );
  OAI211_X1 U16505 ( .C1(n15879), .C2(n7913), .A(n14572), .B(n14571), .ZN(
        n14681) );
  MUX2_X1 U16506 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n14681), .S(n15893), .Z(
        P2_U3529) );
  NAND3_X1 U16507 ( .A1(n14574), .A2(n14573), .A3(n15884), .ZN(n14579) );
  AOI21_X1 U16508 ( .B1(n14576), .B2(n10017), .A(n14575), .ZN(n14577) );
  INV_X1 U16509 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n14586) );
  AOI211_X1 U16510 ( .C1(n14585), .C2(n10017), .A(n14584), .B(n14583), .ZN(
        n14686) );
  MUX2_X1 U16511 ( .A(n14586), .B(n14686), .S(n15893), .Z(n14587) );
  OAI21_X1 U16512 ( .B1(n14689), .B2(n14651), .A(n14587), .ZN(P2_U3524) );
  INV_X1 U16513 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n14591) );
  AOI211_X1 U16514 ( .C1(n14590), .C2(n10017), .A(n14589), .B(n14588), .ZN(
        n14690) );
  MUX2_X1 U16515 ( .A(n14591), .B(n14690), .S(n15893), .Z(n14592) );
  OAI21_X1 U16516 ( .B1(n14651), .B2(n14693), .A(n14592), .ZN(P2_U3523) );
  INV_X1 U16517 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n14596) );
  AOI211_X1 U16518 ( .C1(n14595), .C2(n10017), .A(n14594), .B(n14593), .ZN(
        n14694) );
  MUX2_X1 U16519 ( .A(n14596), .B(n14694), .S(n15893), .Z(n14597) );
  OAI21_X1 U16520 ( .B1(n14697), .B2(n14651), .A(n14597), .ZN(P2_U3522) );
  INV_X1 U16521 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n14601) );
  AOI211_X1 U16522 ( .C1(n14600), .C2(n10017), .A(n14599), .B(n14598), .ZN(
        n14698) );
  MUX2_X1 U16523 ( .A(n14601), .B(n14698), .S(n15893), .Z(n14602) );
  OAI21_X1 U16524 ( .B1(n14701), .B2(n14651), .A(n14602), .ZN(P2_U3521) );
  INV_X1 U16525 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n14606) );
  AOI211_X1 U16526 ( .C1(n14605), .C2(n10017), .A(n14604), .B(n14603), .ZN(
        n14702) );
  MUX2_X1 U16527 ( .A(n14606), .B(n14702), .S(n15893), .Z(n14607) );
  OAI21_X1 U16528 ( .B1(n14705), .B2(n14651), .A(n14607), .ZN(P2_U3520) );
  INV_X1 U16529 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n14611) );
  AOI211_X1 U16530 ( .C1(n14610), .C2(n10017), .A(n14609), .B(n14608), .ZN(
        n14706) );
  MUX2_X1 U16531 ( .A(n14611), .B(n14706), .S(n15893), .Z(n14612) );
  OAI21_X1 U16532 ( .B1(n14651), .B2(n14709), .A(n14612), .ZN(P2_U3519) );
  INV_X1 U16533 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n14616) );
  MUX2_X1 U16534 ( .A(n14616), .B(n14710), .S(n15893), .Z(n14617) );
  OAI21_X1 U16535 ( .B1(n14713), .B2(n14651), .A(n14617), .ZN(P2_U3518) );
  INV_X1 U16536 ( .A(n14618), .ZN(n14623) );
  INV_X1 U16537 ( .A(n15884), .ZN(n14678) );
  AOI21_X1 U16538 ( .B1(n14620), .B2(n10017), .A(n14619), .ZN(n14621) );
  OAI211_X1 U16539 ( .C1(n14623), .C2(n14678), .A(n14622), .B(n14621), .ZN(
        n14714) );
  MUX2_X1 U16540 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14714), .S(n15893), .Z(
        P2_U3517) );
  AOI211_X1 U16541 ( .C1(n14626), .C2(n10017), .A(n14625), .B(n14624), .ZN(
        n14715) );
  MUX2_X1 U16542 ( .A(n14627), .B(n14715), .S(n15893), .Z(n14628) );
  OAI21_X1 U16543 ( .B1(n14718), .B2(n14651), .A(n14628), .ZN(P2_U3516) );
  AOI211_X1 U16544 ( .C1(n14631), .C2(n10017), .A(n14630), .B(n14629), .ZN(
        n14719) );
  MUX2_X1 U16545 ( .A(n14632), .B(n14719), .S(n15893), .Z(n14633) );
  OAI21_X1 U16546 ( .B1(n14651), .B2(n14722), .A(n14633), .ZN(P2_U3515) );
  OAI22_X1 U16547 ( .A1(n14636), .A2(n14635), .B1(n14634), .B2(n15879), .ZN(
        n14637) );
  NOR2_X1 U16548 ( .A1(n14638), .A2(n14637), .ZN(n14723) );
  MUX2_X1 U16549 ( .A(n14639), .B(n14723), .S(n15893), .Z(n14640) );
  OAI21_X1 U16550 ( .B1(n14726), .B2(n14651), .A(n14640), .ZN(P2_U3514) );
  AOI211_X1 U16551 ( .C1(n14643), .C2(n10017), .A(n14642), .B(n14641), .ZN(
        n14727) );
  MUX2_X1 U16552 ( .A(n14644), .B(n14727), .S(n15893), .Z(n14645) );
  OAI21_X1 U16553 ( .B1(n14730), .B2(n14651), .A(n14645), .ZN(P2_U3513) );
  AOI211_X1 U16554 ( .C1(n14648), .C2(n10017), .A(n14647), .B(n14646), .ZN(
        n14731) );
  MUX2_X1 U16555 ( .A(n14649), .B(n14731), .S(n15893), .Z(n14650) );
  OAI21_X1 U16556 ( .B1(n14735), .B2(n14651), .A(n14650), .ZN(P2_U3512) );
  AOI21_X1 U16557 ( .B1(n14653), .B2(n10017), .A(n14652), .ZN(n14654) );
  OAI211_X1 U16558 ( .C1(n14656), .C2(n14673), .A(n14655), .B(n14654), .ZN(
        n14736) );
  MUX2_X1 U16559 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n14736), .S(n15893), .Z(
        P2_U3511) );
  AOI21_X1 U16560 ( .B1(n14658), .B2(n10017), .A(n14657), .ZN(n14659) );
  OAI211_X1 U16561 ( .C1(n14661), .C2(n14673), .A(n14660), .B(n14659), .ZN(
        n14737) );
  MUX2_X1 U16562 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n14737), .S(n15893), .Z(
        P2_U3510) );
  AOI21_X1 U16563 ( .B1(n14663), .B2(n10017), .A(n14662), .ZN(n14664) );
  OAI211_X1 U16564 ( .C1(n14666), .C2(n14678), .A(n14665), .B(n14664), .ZN(
        n14738) );
  MUX2_X1 U16565 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n14738), .S(n15893), .Z(
        P2_U3508) );
  AOI21_X1 U16566 ( .B1(n14668), .B2(n10017), .A(n14667), .ZN(n14671) );
  INV_X1 U16567 ( .A(n14669), .ZN(n14670) );
  OAI211_X1 U16568 ( .C1(n14673), .C2(n14672), .A(n14671), .B(n14670), .ZN(
        n14739) );
  MUX2_X1 U16569 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n14739), .S(n15893), .Z(
        P2_U3507) );
  AOI21_X1 U16570 ( .B1(n14675), .B2(n10017), .A(n14674), .ZN(n14676) );
  OAI211_X1 U16571 ( .C1(n14679), .C2(n14678), .A(n14677), .B(n14676), .ZN(
        n14740) );
  MUX2_X1 U16572 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n14740), .S(n15893), .Z(
        P2_U3505) );
  MUX2_X1 U16573 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n14680), .S(n15886), .Z(
        P2_U3498) );
  MUX2_X1 U16574 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n14681), .S(n15886), .Z(
        P2_U3497) );
  MUX2_X1 U16575 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14682), .S(n15886), .Z(
        n14683) );
  INV_X1 U16576 ( .A(n14683), .ZN(n14684) );
  INV_X1 U16577 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n14687) );
  MUX2_X1 U16578 ( .A(n14687), .B(n14686), .S(n15886), .Z(n14688) );
  OAI21_X1 U16579 ( .B1(n14689), .B2(n14734), .A(n14688), .ZN(P2_U3492) );
  MUX2_X1 U16580 ( .A(n14691), .B(n14690), .S(n15886), .Z(n14692) );
  OAI21_X1 U16581 ( .B1(n14693), .B2(n14734), .A(n14692), .ZN(P2_U3491) );
  INV_X1 U16582 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n14695) );
  MUX2_X1 U16583 ( .A(n14695), .B(n14694), .S(n15886), .Z(n14696) );
  OAI21_X1 U16584 ( .B1(n14697), .B2(n14734), .A(n14696), .ZN(P2_U3490) );
  INV_X1 U16585 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n14699) );
  MUX2_X1 U16586 ( .A(n14699), .B(n14698), .S(n15886), .Z(n14700) );
  OAI21_X1 U16587 ( .B1(n14701), .B2(n14734), .A(n14700), .ZN(P2_U3489) );
  INV_X1 U16588 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n14703) );
  MUX2_X1 U16589 ( .A(n14703), .B(n14702), .S(n15886), .Z(n14704) );
  OAI21_X1 U16590 ( .B1(n14705), .B2(n14734), .A(n14704), .ZN(P2_U3488) );
  INV_X1 U16591 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n14707) );
  MUX2_X1 U16592 ( .A(n14707), .B(n14706), .S(n15886), .Z(n14708) );
  OAI21_X1 U16593 ( .B1(n14709), .B2(n14734), .A(n14708), .ZN(P2_U3487) );
  INV_X1 U16594 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n14711) );
  MUX2_X1 U16595 ( .A(n14711), .B(n14710), .S(n15886), .Z(n14712) );
  OAI21_X1 U16596 ( .B1(n14713), .B2(n14734), .A(n14712), .ZN(P2_U3486) );
  MUX2_X1 U16597 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14714), .S(n15886), .Z(
        P2_U3484) );
  INV_X1 U16598 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n14716) );
  MUX2_X1 U16599 ( .A(n14716), .B(n14715), .S(n15886), .Z(n14717) );
  OAI21_X1 U16600 ( .B1(n14718), .B2(n14734), .A(n14717), .ZN(P2_U3481) );
  INV_X1 U16601 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n14720) );
  MUX2_X1 U16602 ( .A(n14720), .B(n14719), .S(n15886), .Z(n14721) );
  OAI21_X1 U16603 ( .B1(n14722), .B2(n14734), .A(n14721), .ZN(P2_U3478) );
  MUX2_X1 U16604 ( .A(n14724), .B(n14723), .S(n15886), .Z(n14725) );
  OAI21_X1 U16605 ( .B1(n14726), .B2(n14734), .A(n14725), .ZN(P2_U3475) );
  MUX2_X1 U16606 ( .A(n14728), .B(n14727), .S(n15886), .Z(n14729) );
  OAI21_X1 U16607 ( .B1(n14730), .B2(n14734), .A(n14729), .ZN(P2_U3472) );
  INV_X1 U16608 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14732) );
  MUX2_X1 U16609 ( .A(n14732), .B(n14731), .S(n15886), .Z(n14733) );
  OAI21_X1 U16610 ( .B1(n14735), .B2(n14734), .A(n14733), .ZN(P2_U3469) );
  MUX2_X1 U16611 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n14736), .S(n15886), .Z(
        P2_U3466) );
  MUX2_X1 U16612 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n14737), .S(n15886), .Z(
        P2_U3463) );
  MUX2_X1 U16613 ( .A(P2_REG0_REG_9__SCAN_IN), .B(n14738), .S(n15886), .Z(
        P2_U3457) );
  MUX2_X1 U16614 ( .A(P2_REG0_REG_8__SCAN_IN), .B(n14739), .S(n15886), .Z(
        P2_U3454) );
  MUX2_X1 U16615 ( .A(P2_REG0_REG_6__SCAN_IN), .B(n14740), .S(n15886), .Z(
        P2_U3448) );
  INV_X1 U16616 ( .A(n14741), .ZN(n14742) );
  MUX2_X1 U16617 ( .A(n14742), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XNOR2_X1 U16618 ( .A(n14744), .B(n14743), .ZN(n14749) );
  AND2_X1 U16619 ( .A1(n14937), .A2(n15637), .ZN(n14745) );
  AOI21_X1 U16620 ( .B1(n14935), .B2(n15636), .A(n14745), .ZN(n15146) );
  AOI22_X1 U16621 ( .A1(n15149), .A2(n14926), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14746) );
  OAI21_X1 U16622 ( .B1(n15146), .B2(n14928), .A(n14746), .ZN(n14747) );
  AOI21_X1 U16623 ( .B1(n15150), .B2(n14930), .A(n14747), .ZN(n14748) );
  OAI21_X1 U16624 ( .B1(n14749), .B2(n15634), .A(n14748), .ZN(P1_U3214) );
  XOR2_X1 U16625 ( .A(n14750), .B(n14751), .Z(n14759) );
  INV_X1 U16626 ( .A(n14752), .ZN(n15348) );
  OR2_X1 U16627 ( .A1(n14830), .A2(n14913), .ZN(n14753) );
  OAI21_X1 U16628 ( .B1(n14754), .B2(n14922), .A(n14753), .ZN(n15485) );
  AOI21_X1 U16629 ( .B1(n15485), .B2(n15641), .A(n14755), .ZN(n14756) );
  OAI21_X1 U16630 ( .B1(n15348), .B2(n15646), .A(n14756), .ZN(n14757) );
  AOI21_X1 U16631 ( .B1(n15486), .B2(n14930), .A(n14757), .ZN(n14758) );
  OAI21_X1 U16632 ( .B1(n14759), .B2(n15634), .A(n14758), .ZN(P1_U3215) );
  NAND2_X1 U16633 ( .A1(n14760), .A2(n14761), .ZN(n14762) );
  XOR2_X1 U16634 ( .A(n14763), .B(n14762), .Z(n14769) );
  AND2_X1 U16635 ( .A1(n14941), .A2(n15637), .ZN(n14764) );
  AOI21_X1 U16636 ( .B1(n14939), .B2(n15636), .A(n14764), .ZN(n15429) );
  INV_X1 U16637 ( .A(n14765), .ZN(n15205) );
  AOI22_X1 U16638 ( .A1(n15205), .A2(n14926), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14766) );
  OAI21_X1 U16639 ( .B1(n15429), .B2(n14928), .A(n14766), .ZN(n14767) );
  AOI21_X1 U16640 ( .B1(n15428), .B2(n14930), .A(n14767), .ZN(n14768) );
  OAI21_X1 U16641 ( .B1(n14769), .B2(n15634), .A(n14768), .ZN(P1_U3216) );
  XNOR2_X1 U16642 ( .A(n14770), .B(n14771), .ZN(n14852) );
  AOI22_X1 U16643 ( .A1(n14852), .A2(n14773), .B1(n14772), .B2(n14770), .ZN(
        n14777) );
  XNOR2_X1 U16644 ( .A(n14775), .B(n14774), .ZN(n14776) );
  XNOR2_X1 U16645 ( .A(n14777), .B(n14776), .ZN(n14786) );
  INV_X1 U16646 ( .A(n14778), .ZN(n14779) );
  NOR2_X1 U16647 ( .A1(n14779), .A2(n15742), .ZN(n15507) );
  NAND2_X1 U16648 ( .A1(n14781), .A2(n14780), .ZN(n15505) );
  AOI22_X1 U16649 ( .A1(n15641), .A2(n15505), .B1(P1_REG3_REG_10__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14782) );
  OAI21_X1 U16650 ( .B1(n14783), .B2(n15646), .A(n14782), .ZN(n14784) );
  AOI21_X1 U16651 ( .B1(n15507), .B2(n15632), .A(n14784), .ZN(n14785) );
  OAI21_X1 U16652 ( .B1(n14786), .B2(n15634), .A(n14785), .ZN(P1_U3217) );
  INV_X1 U16653 ( .A(n15455), .ZN(n15276) );
  OAI211_X1 U16654 ( .C1(n14789), .C2(n14788), .A(n14787), .B(n14910), .ZN(
        n14794) );
  NAND2_X1 U16655 ( .A1(n14943), .A2(n15636), .ZN(n14791) );
  OR2_X1 U16656 ( .A1(n14838), .A2(n14922), .ZN(n14790) );
  NAND2_X1 U16657 ( .A1(n14791), .A2(n14790), .ZN(n15454) );
  NAND2_X1 U16658 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n15113)
         );
  OAI21_X1 U16659 ( .B1(n15646), .B2(n15271), .A(n15113), .ZN(n14792) );
  AOI21_X1 U16660 ( .B1(n15454), .B2(n15641), .A(n14792), .ZN(n14793) );
  OAI211_X1 U16661 ( .C1(n15276), .C2(n14918), .A(n14794), .B(n14793), .ZN(
        P1_U3219) );
  OAI21_X1 U16662 ( .B1(n14797), .B2(n14796), .A(n14795), .ZN(n14798) );
  NAND2_X1 U16663 ( .A1(n14798), .A2(n14910), .ZN(n14804) );
  NAND2_X1 U16664 ( .A1(n14941), .A2(n15636), .ZN(n14800) );
  NAND2_X1 U16665 ( .A1(n14943), .A2(n15637), .ZN(n14799) );
  NAND2_X1 U16666 ( .A1(n14800), .A2(n14799), .ZN(n15236) );
  OAI22_X1 U16667 ( .A1(n15229), .A2(n15646), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14801), .ZN(n14802) );
  AOI21_X1 U16668 ( .B1(n15236), .B2(n15641), .A(n14802), .ZN(n14803) );
  OAI211_X1 U16669 ( .C1(n14805), .C2(n14918), .A(n14804), .B(n14803), .ZN(
        P1_U3223) );
  OAI211_X1 U16670 ( .C1(n14808), .C2(n14807), .A(n14806), .B(n14910), .ZN(
        n14814) );
  OAI21_X1 U16671 ( .B1(n14810), .B2(n14928), .A(n14809), .ZN(n14811) );
  AOI21_X1 U16672 ( .B1(n14812), .B2(n14926), .A(n14811), .ZN(n14813) );
  OAI211_X1 U16673 ( .C1(n7298), .C2(n14918), .A(n14814), .B(n14813), .ZN(
        P1_U3224) );
  NAND2_X1 U16674 ( .A1(n14937), .A2(n15636), .ZN(n14819) );
  NAND2_X1 U16675 ( .A1(n14939), .A2(n15637), .ZN(n14818) );
  AND2_X1 U16676 ( .A1(n14819), .A2(n14818), .ZN(n15416) );
  AOI22_X1 U16677 ( .A1(n15174), .A2(n14926), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14820) );
  OAI21_X1 U16678 ( .B1(n15416), .B2(n14928), .A(n14820), .ZN(n14821) );
  AOI21_X1 U16679 ( .B1(n14822), .B2(n14930), .A(n14821), .ZN(n14823) );
  XNOR2_X1 U16680 ( .A(n14824), .B(n14825), .ZN(n14921) );
  NOR2_X1 U16681 ( .A1(n14921), .A2(n14920), .ZN(n14919) );
  AOI21_X1 U16682 ( .B1(n14825), .B2(n14824), .A(n14919), .ZN(n14829) );
  XNOR2_X1 U16683 ( .A(n14827), .B(n14826), .ZN(n14828) );
  XNOR2_X1 U16684 ( .A(n14829), .B(n14828), .ZN(n14835) );
  OAI22_X1 U16685 ( .A1(n14831), .A2(n14913), .B1(n14830), .B2(n14922), .ZN(
        n15308) );
  NAND2_X1 U16686 ( .A1(n15308), .A2(n15641), .ZN(n14832) );
  NAND2_X1 U16687 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n15061)
         );
  OAI211_X1 U16688 ( .C1(n15646), .C2(n15315), .A(n14832), .B(n15061), .ZN(
        n14833) );
  AOI21_X1 U16689 ( .B1(n15472), .B2(n14930), .A(n14833), .ZN(n14834) );
  OAI21_X1 U16690 ( .B1(n14835), .B2(n15634), .A(n14834), .ZN(P1_U3226) );
  XOR2_X1 U16691 ( .A(n14836), .B(n14837), .Z(n14844) );
  OR2_X1 U16692 ( .A1(n14838), .A2(n14913), .ZN(n14840) );
  NAND2_X1 U16693 ( .A1(n14947), .A2(n15637), .ZN(n14839) );
  AND2_X1 U16694 ( .A1(n14840), .A2(n14839), .ZN(n15464) );
  NAND2_X1 U16695 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n15067)
         );
  NAND2_X1 U16696 ( .A1(n14926), .A2(n15300), .ZN(n14841) );
  OAI211_X1 U16697 ( .C1(n15464), .C2(n14928), .A(n15067), .B(n14841), .ZN(
        n14842) );
  AOI21_X1 U16698 ( .B1(n15303), .B2(n14930), .A(n14842), .ZN(n14843) );
  OAI21_X1 U16699 ( .B1(n14844), .B2(n15634), .A(n14843), .ZN(P1_U3228) );
  XOR2_X1 U16700 ( .A(n14846), .B(n14845), .Z(n14850) );
  AOI22_X1 U16701 ( .A1(n14938), .A2(n15636), .B1(n15637), .B2(n14940), .ZN(
        n15187) );
  AOI22_X1 U16702 ( .A1(n15192), .A2(n14926), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14847) );
  OAI21_X1 U16703 ( .B1(n15187), .B2(n14928), .A(n14847), .ZN(n14848) );
  AOI21_X1 U16704 ( .B1(n15425), .B2(n14930), .A(n14848), .ZN(n14849) );
  OAI21_X1 U16705 ( .B1(n14850), .B2(n15634), .A(n14849), .ZN(P1_U3229) );
  XNOR2_X1 U16706 ( .A(n14852), .B(n14851), .ZN(n14859) );
  NOR2_X1 U16707 ( .A1(n14853), .A2(n15742), .ZN(n15513) );
  AOI21_X1 U16708 ( .B1(n15641), .B2(n15511), .A(n14854), .ZN(n14855) );
  OAI21_X1 U16709 ( .B1(n15646), .B2(n14856), .A(n14855), .ZN(n14857) );
  AOI21_X1 U16710 ( .B1(n15513), .B2(n15632), .A(n14857), .ZN(n14858) );
  OAI21_X1 U16711 ( .B1(n14859), .B2(n15634), .A(n14858), .ZN(P1_U3231) );
  INV_X1 U16712 ( .A(n14860), .ZN(n14861) );
  OAI211_X1 U16713 ( .C1(n14863), .C2(n14862), .A(n14861), .B(n14910), .ZN(
        n14869) );
  NAND2_X1 U16714 ( .A1(n14942), .A2(n15636), .ZN(n14865) );
  NAND2_X1 U16715 ( .A1(n14944), .A2(n15637), .ZN(n14864) );
  NAND2_X1 U16716 ( .A1(n14865), .A2(n14864), .ZN(n15250) );
  OAI22_X1 U16717 ( .A1(n15646), .A2(n15255), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14866), .ZN(n14867) );
  AOI21_X1 U16718 ( .B1(n15250), .B2(n15641), .A(n14867), .ZN(n14868) );
  OAI211_X1 U16719 ( .C1(n15252), .C2(n14918), .A(n14869), .B(n14868), .ZN(
        P1_U3233) );
  AOI21_X1 U16720 ( .B1(n14872), .B2(n14871), .A(n14870), .ZN(n14880) );
  OR2_X1 U16721 ( .A1(n14873), .A2(n14922), .ZN(n14875) );
  OR2_X1 U16722 ( .A1(n14923), .A2(n14913), .ZN(n14874) );
  NAND2_X1 U16723 ( .A1(n14875), .A2(n14874), .ZN(n15358) );
  NAND2_X1 U16724 ( .A1(n15641), .A2(n15358), .ZN(n14876) );
  OAI211_X1 U16725 ( .C1(n15646), .C2(n15364), .A(n14877), .B(n14876), .ZN(
        n14878) );
  AOI21_X1 U16726 ( .B1(n15491), .B2(n14930), .A(n14878), .ZN(n14879) );
  OAI21_X1 U16727 ( .B1(n14880), .B2(n15634), .A(n14879), .ZN(P1_U3234) );
  OAI21_X1 U16728 ( .B1(n14882), .B2(n14881), .A(n14760), .ZN(n14883) );
  NAND2_X1 U16729 ( .A1(n14883), .A2(n14910), .ZN(n14890) );
  NAND2_X1 U16730 ( .A1(n14940), .A2(n15636), .ZN(n14885) );
  NAND2_X1 U16731 ( .A1(n14942), .A2(n15637), .ZN(n14884) );
  NAND2_X1 U16732 ( .A1(n14885), .A2(n14884), .ZN(n15216) );
  INV_X1 U16733 ( .A(n15220), .ZN(n14887) );
  OAI22_X1 U16734 ( .A1(n14887), .A2(n15646), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14886), .ZN(n14888) );
  AOI21_X1 U16735 ( .B1(n15216), .B2(n15641), .A(n14888), .ZN(n14889) );
  OAI211_X1 U16736 ( .C1(n14918), .C2(n15223), .A(n14890), .B(n14889), .ZN(
        P1_U3235) );
  NAND2_X1 U16737 ( .A1(n14891), .A2(n15757), .ZN(n15503) );
  XNOR2_X1 U16738 ( .A(n14893), .B(n14892), .ZN(n14894) );
  NAND2_X1 U16739 ( .A1(n14894), .A2(n14910), .ZN(n14900) );
  NOR2_X1 U16740 ( .A1(n15646), .A2(n14895), .ZN(n14896) );
  AOI211_X1 U16741 ( .C1(n15641), .C2(n14898), .A(n14897), .B(n14896), .ZN(
        n14899) );
  OAI211_X1 U16742 ( .C1(n14901), .C2(n15503), .A(n14900), .B(n14899), .ZN(
        P1_U3236) );
  XOR2_X1 U16743 ( .A(n14903), .B(n14902), .Z(n14907) );
  AOI22_X1 U16744 ( .A1(n14944), .A2(n15636), .B1(n15637), .B2(n14946), .ZN(
        n15283) );
  NAND2_X1 U16745 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n15082)
         );
  NAND2_X1 U16746 ( .A1(n14926), .A2(n15287), .ZN(n14904) );
  OAI211_X1 U16747 ( .C1(n15283), .C2(n14928), .A(n15082), .B(n14904), .ZN(
        n14905) );
  AOI21_X1 U16748 ( .B1(n15461), .B2(n14930), .A(n14905), .ZN(n14906) );
  OAI21_X1 U16749 ( .B1(n14907), .B2(n15634), .A(n14906), .ZN(P1_U3238) );
  XNOR2_X1 U16750 ( .A(n14909), .B(n14908), .ZN(n14911) );
  OAI22_X1 U16751 ( .A1(n14914), .A2(n14913), .B1(n14912), .B2(n14922), .ZN(
        n15157) );
  OAI22_X1 U16752 ( .A1(n15161), .A2(n15646), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14915), .ZN(n14916) );
  AOI21_X1 U16753 ( .B1(n15157), .B2(n15641), .A(n14916), .ZN(n14917) );
  AOI21_X1 U16754 ( .B1(n14921), .B2(n14920), .A(n14919), .ZN(n14932) );
  NAND2_X1 U16755 ( .A1(n14947), .A2(n15636), .ZN(n14925) );
  OR2_X1 U16756 ( .A1(n14923), .A2(n14922), .ZN(n14924) );
  AND2_X1 U16757 ( .A1(n14925), .A2(n14924), .ZN(n15476) );
  NAND2_X1 U16758 ( .A1(n14926), .A2(n15331), .ZN(n14927) );
  NAND2_X1 U16759 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n15666)
         );
  OAI211_X1 U16760 ( .C1(n15476), .C2(n14928), .A(n14927), .B(n15666), .ZN(
        n14929) );
  AOI21_X1 U16761 ( .B1(n15479), .B2(n14930), .A(n14929), .ZN(n14931) );
  OAI21_X1 U16762 ( .B1(n14932), .B2(n15634), .A(n14931), .ZN(P1_U3241) );
  MUX2_X1 U16763 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n15118), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U16764 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14933), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16765 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14934), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16766 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14935), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16767 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14936), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16768 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14937), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16769 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14938), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16770 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14939), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16771 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14940), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16772 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14941), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16773 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14942), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16774 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14943), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16775 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14944), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16776 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14945), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16777 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14946), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16778 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14947), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16779 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n12498), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16780 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14948), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16781 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14949), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16782 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14950), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16783 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14951), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16784 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14952), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16785 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14953), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16786 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14954), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16787 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14955), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16788 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14956), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16789 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n6539), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16790 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n6540), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16791 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14957), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16792 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n15638), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16793 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9465), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16794 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14958), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI211_X1 U16795 ( .C1(n14961), .C2(n14960), .A(n15665), .B(n14959), .ZN(
        n14971) );
  INV_X1 U16796 ( .A(n14962), .ZN(n14966) );
  OAI21_X1 U16797 ( .B1(n14964), .B2(n15648), .A(n14963), .ZN(n14965) );
  NAND3_X1 U16798 ( .A1(n15108), .A2(n14966), .A3(n14965), .ZN(n14970) );
  NAND2_X1 U16799 ( .A1(n15085), .A2(n14967), .ZN(n14969) );
  AOI22_X1 U16800 ( .A1(n15651), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14968) );
  NAND4_X1 U16801 ( .A1(n14971), .A2(n14970), .A3(n14969), .A4(n14968), .ZN(
        P1_U3244) );
  AND2_X1 U16802 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n14973) );
  NOR2_X1 U16803 ( .A1(n15659), .A2(n14977), .ZN(n14972) );
  AOI211_X1 U16804 ( .C1(n15651), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n14973), .B(
        n14972), .ZN(n14985) );
  OAI211_X1 U16805 ( .C1(n14976), .C2(n14975), .A(n15665), .B(n14974), .ZN(
        n14984) );
  MUX2_X1 U16806 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10574), .S(n14977), .Z(
        n14980) );
  INV_X1 U16807 ( .A(n14978), .ZN(n14979) );
  NAND2_X1 U16808 ( .A1(n14980), .A2(n14979), .ZN(n14981) );
  OAI211_X1 U16809 ( .C1(n14982), .C2(n14981), .A(n15108), .B(n14995), .ZN(
        n14983) );
  NAND3_X1 U16810 ( .A1(n14985), .A2(n14984), .A3(n14983), .ZN(P1_U3246) );
  NAND2_X1 U16811 ( .A1(n15651), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n14986) );
  OAI211_X1 U16812 ( .C1(n15659), .C2(n14988), .A(n14987), .B(n14986), .ZN(
        n14989) );
  INV_X1 U16813 ( .A(n14989), .ZN(n14999) );
  OAI211_X1 U16814 ( .C1(n14992), .C2(n14991), .A(n15665), .B(n14990), .ZN(
        n14998) );
  NAND3_X1 U16815 ( .A1(n14995), .A2(n14994), .A3(n14993), .ZN(n14996) );
  NAND3_X1 U16816 ( .A1(n15108), .A2(n6789), .A3(n14996), .ZN(n14997) );
  NAND4_X1 U16817 ( .A1(n15000), .A2(n14999), .A3(n14998), .A4(n14997), .ZN(
        P1_U3247) );
  MUX2_X1 U16818 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n15001), .S(n15007), .Z(
        n15003) );
  OAI211_X1 U16819 ( .C1(n6788), .C2(n15003), .A(n15108), .B(n15002), .ZN(
        n15013) );
  AND2_X1 U16820 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n15006) );
  NOR2_X1 U16821 ( .A1(n15668), .A2(n15004), .ZN(n15005) );
  AOI211_X1 U16822 ( .C1(n15085), .C2(n15007), .A(n15006), .B(n15005), .ZN(
        n15012) );
  OAI211_X1 U16823 ( .C1(n15010), .C2(n15009), .A(n15665), .B(n15008), .ZN(
        n15011) );
  NAND3_X1 U16824 ( .A1(n15013), .A2(n15012), .A3(n15011), .ZN(P1_U3249) );
  NOR2_X1 U16825 ( .A1(n15015), .A2(n15014), .ZN(n15017) );
  OAI21_X1 U16826 ( .B1(n15017), .B2(n15016), .A(n15108), .ZN(n15026) );
  AND2_X1 U16827 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n15020) );
  NOR2_X1 U16828 ( .A1(n15659), .A2(n15018), .ZN(n15019) );
  AOI211_X1 U16829 ( .C1(n15651), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n15020), .B(
        n15019), .ZN(n15025) );
  OAI211_X1 U16830 ( .C1(n15023), .C2(n15022), .A(n15021), .B(n15665), .ZN(
        n15024) );
  NAND3_X1 U16831 ( .A1(n15026), .A2(n15025), .A3(n15024), .ZN(P1_U3251) );
  INV_X1 U16832 ( .A(n15027), .ZN(n15032) );
  OAI21_X1 U16833 ( .B1(n15030), .B2(n15029), .A(n15028), .ZN(n15031) );
  NAND3_X1 U16834 ( .A1(n15032), .A2(n15108), .A3(n15031), .ZN(n15041) );
  AND2_X1 U16835 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n15033) );
  AOI21_X1 U16836 ( .B1(n15651), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n15033), 
        .ZN(n15040) );
  OAI211_X1 U16837 ( .C1(n15036), .C2(n15035), .A(n15034), .B(n15665), .ZN(
        n15039) );
  NAND2_X1 U16838 ( .A1(n15085), .A2(n15037), .ZN(n15038) );
  NAND4_X1 U16839 ( .A1(n15041), .A2(n15040), .A3(n15039), .A4(n15038), .ZN(
        P1_U3253) );
  XNOR2_X1 U16840 ( .A(n15070), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n15049) );
  NOR2_X1 U16841 ( .A1(n15045), .A2(n15053), .ZN(n15047) );
  OR2_X1 U16842 ( .A1(n15047), .A2(n15657), .ZN(n15048) );
  AOI211_X1 U16843 ( .C1(n15049), .C2(n15048), .A(n15661), .B(n15066), .ZN(
        n15065) );
  XNOR2_X1 U16844 ( .A(n15070), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n15059) );
  NAND2_X1 U16845 ( .A1(n15050), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n15051) );
  NAND2_X1 U16846 ( .A1(n15052), .A2(n15051), .ZN(n15054) );
  XNOR2_X1 U16847 ( .A(n15054), .B(n15660), .ZN(n15656) );
  INV_X1 U16848 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n15655) );
  NAND2_X1 U16849 ( .A1(n15656), .A2(n15655), .ZN(n15056) );
  OR2_X1 U16850 ( .A1(n15054), .A2(n15053), .ZN(n15055) );
  NAND2_X1 U16851 ( .A1(n15056), .A2(n15055), .ZN(n15058) );
  INV_X1 U16852 ( .A(n15072), .ZN(n15057) );
  AOI211_X1 U16853 ( .C1(n15059), .C2(n15058), .A(n15111), .B(n15057), .ZN(
        n15064) );
  NAND2_X1 U16854 ( .A1(n15651), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n15060) );
  OAI211_X1 U16855 ( .C1(n15659), .C2(n15062), .A(n15061), .B(n15060), .ZN(
        n15063) );
  OR3_X1 U16856 ( .A1(n15065), .A2(n15064), .A3(n15063), .ZN(P1_U3259) );
  XNOR2_X1 U16857 ( .A(n15086), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n15081) );
  XNOR2_X1 U16858 ( .A(n6625), .B(n15081), .ZN(n15078) );
  INV_X1 U16859 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n15068) );
  OAI21_X1 U16860 ( .B1(n15668), .B2(n15068), .A(n15067), .ZN(n15069) );
  AOI21_X1 U16861 ( .B1(n15086), .B2(n15085), .A(n15069), .ZN(n15077) );
  NAND2_X1 U16862 ( .A1(n15070), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n15071) );
  NAND2_X1 U16863 ( .A1(n15072), .A2(n15071), .ZN(n15075) );
  INV_X1 U16864 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n15073) );
  XNOR2_X1 U16865 ( .A(n15086), .B(n15073), .ZN(n15074) );
  NAND2_X1 U16866 ( .A1(n15075), .A2(n15074), .ZN(n15088) );
  OAI211_X1 U16867 ( .C1(n15075), .C2(n15074), .A(n15088), .B(n15665), .ZN(
        n15076) );
  OAI211_X1 U16868 ( .C1(n15078), .C2(n15661), .A(n15077), .B(n15076), .ZN(
        P1_U3260) );
  OAI22_X1 U16869 ( .A1(n6625), .A2(n15081), .B1(n15080), .B2(n15079), .ZN(
        n15098) );
  XNOR2_X1 U16870 ( .A(n15098), .B(n15089), .ZN(n15102) );
  XOR2_X1 U16871 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15102), .Z(n15097) );
  INV_X1 U16872 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15083) );
  OAI21_X1 U16873 ( .B1(n15668), .B2(n15083), .A(n15082), .ZN(n15084) );
  AOI21_X1 U16874 ( .B1(n15089), .B2(n15085), .A(n15084), .ZN(n15096) );
  NAND2_X1 U16875 ( .A1(n15086), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n15087) );
  NAND2_X1 U16876 ( .A1(n15088), .A2(n15087), .ZN(n15090) );
  NAND2_X1 U16877 ( .A1(n15090), .A2(n15089), .ZN(n15104) );
  OR2_X1 U16878 ( .A1(n15090), .A2(n15089), .ZN(n15091) );
  NAND2_X1 U16879 ( .A1(n15104), .A2(n15091), .ZN(n15093) );
  INV_X1 U16880 ( .A(n15093), .ZN(n15094) );
  OAI211_X1 U16881 ( .C1(n15094), .C2(P1_REG2_REG_18__SCAN_IN), .A(n15665), 
        .B(n15105), .ZN(n15095) );
  OAI211_X1 U16882 ( .C1(n15097), .C2(n15661), .A(n15096), .B(n15095), .ZN(
        P1_U3261) );
  INV_X1 U16883 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n15101) );
  INV_X1 U16884 ( .A(n15098), .ZN(n15100) );
  OAI22_X1 U16885 ( .A1(n15102), .A2(n15101), .B1(n15100), .B2(n15099), .ZN(
        n15103) );
  XNOR2_X1 U16886 ( .A(n15103), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n15109) );
  NAND2_X1 U16887 ( .A1(n15105), .A2(n15104), .ZN(n15106) );
  INV_X1 U16888 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n15272) );
  XNOR2_X1 U16889 ( .A(n15106), .B(n15272), .ZN(n15110) );
  INV_X1 U16890 ( .A(n15110), .ZN(n15107) );
  XNOR2_X1 U16891 ( .A(n15379), .B(n15115), .ZN(n15116) );
  NAND2_X1 U16892 ( .A1(n15116), .A2(n15678), .ZN(n15378) );
  NAND2_X1 U16893 ( .A1(n15118), .A2(n15117), .ZN(n15381) );
  NOR2_X1 U16894 ( .A1(n6546), .A2(n15381), .ZN(n15125) );
  NOR2_X1 U16895 ( .A1(n15379), .A2(n15367), .ZN(n15119) );
  AOI211_X1 U16896 ( .C1(n6546), .C2(P1_REG2_REG_31__SCAN_IN), .A(n15125), .B(
        n15119), .ZN(n15120) );
  OAI21_X1 U16897 ( .B1(n15686), .B2(n15378), .A(n15120), .ZN(P1_U3263) );
  XNOR2_X1 U16898 ( .A(n15122), .B(n15121), .ZN(n15380) );
  INV_X1 U16899 ( .A(n15259), .ZN(n15123) );
  NAND2_X1 U16900 ( .A1(n15380), .A2(n15123), .ZN(n15127) );
  AND2_X1 U16901 ( .A1(n6546), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n15124) );
  NOR2_X1 U16902 ( .A1(n15125), .A2(n15124), .ZN(n15126) );
  OAI211_X1 U16903 ( .C1(n15383), .C2(n15367), .A(n15127), .B(n15126), .ZN(
        P1_U3264) );
  AOI21_X1 U16904 ( .B1(n15148), .B2(n15135), .A(n15733), .ZN(n15131) );
  NAND2_X1 U16905 ( .A1(n15131), .A2(n15130), .ZN(n15399) );
  AOI22_X1 U16906 ( .A1(n15132), .A2(n15698), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n6546), .ZN(n15133) );
  OAI21_X1 U16907 ( .B1(n15398), .B2(n6546), .A(n15133), .ZN(n15134) );
  AOI21_X1 U16908 ( .B1(n15135), .B2(n15716), .A(n15134), .ZN(n15136) );
  OAI21_X1 U16909 ( .B1(n15399), .B2(n15686), .A(n15136), .ZN(n15137) );
  AOI21_X1 U16910 ( .B1(n15402), .B2(n15295), .A(n15137), .ZN(n15138) );
  OAI21_X1 U16911 ( .B1(n15403), .B2(n15374), .A(n15138), .ZN(P1_U3265) );
  NAND2_X1 U16912 ( .A1(n15404), .A2(n15711), .ZN(n15147) );
  AND2_X1 U16913 ( .A1(n15142), .A2(n15141), .ZN(n15143) );
  OAI21_X1 U16914 ( .B1(n15144), .B2(n15143), .A(n15763), .ZN(n15145) );
  OAI211_X1 U16915 ( .C1(n15159), .C2(n15407), .A(n15678), .B(n15148), .ZN(
        n15405) );
  AOI22_X1 U16916 ( .A1(n15149), .A2(n15698), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n6546), .ZN(n15152) );
  NAND2_X1 U16917 ( .A1(n15150), .A2(n15716), .ZN(n15151) );
  OAI211_X1 U16918 ( .C1(n15405), .C2(n15686), .A(n15152), .B(n15151), .ZN(
        n15153) );
  AOI21_X1 U16919 ( .B1(n15404), .B2(n15719), .A(n15153), .ZN(n15154) );
  OAI21_X1 U16920 ( .B1(n6630), .B2(n6546), .A(n15154), .ZN(P1_U3266) );
  XNOR2_X1 U16921 ( .A(n15155), .B(n15156), .ZN(n15415) );
  INV_X1 U16922 ( .A(n15414), .ZN(n15166) );
  NOR2_X1 U16923 ( .A1(n15172), .A2(n15410), .ZN(n15158) );
  OR2_X1 U16924 ( .A1(n15159), .A2(n15158), .ZN(n15411) );
  INV_X1 U16925 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n15160) );
  OAI22_X1 U16926 ( .A1(n15161), .A2(n15712), .B1(n15160), .B2(n15714), .ZN(
        n15162) );
  AOI21_X1 U16927 ( .B1(n15163), .B2(n15716), .A(n15162), .ZN(n15164) );
  OAI21_X1 U16928 ( .B1(n15411), .B2(n15259), .A(n15164), .ZN(n15165) );
  AOI21_X1 U16929 ( .B1(n15166), .B2(n15714), .A(n15165), .ZN(n15167) );
  OAI21_X1 U16930 ( .B1(n15415), .B2(n15374), .A(n15167), .ZN(P1_U3267) );
  OAI21_X1 U16931 ( .B1(n6651), .B2(n15169), .A(n15168), .ZN(n15422) );
  OAI21_X1 U16932 ( .B1(n6536), .B2(n15171), .A(n15170), .ZN(n15420) );
  OAI21_X1 U16933 ( .B1(n15191), .B2(n15417), .A(n15678), .ZN(n15173) );
  NOR2_X1 U16934 ( .A1(n15173), .A2(n15172), .ZN(n15419) );
  NAND2_X1 U16935 ( .A1(n15419), .A2(n15720), .ZN(n15179) );
  NAND2_X1 U16936 ( .A1(n15174), .A2(n15698), .ZN(n15175) );
  NAND2_X1 U16937 ( .A1(n15416), .A2(n15175), .ZN(n15177) );
  AND2_X1 U16938 ( .A1(n6546), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n15176) );
  AOI21_X1 U16939 ( .B1(n15177), .B2(n15714), .A(n15176), .ZN(n15178) );
  OAI211_X1 U16940 ( .C1(n15417), .C2(n15367), .A(n15179), .B(n15178), .ZN(
        n15180) );
  AOI21_X1 U16941 ( .B1(n15420), .B2(n15295), .A(n15180), .ZN(n15181) );
  OAI21_X1 U16942 ( .B1(n15374), .B2(n15422), .A(n15181), .ZN(P1_U3268) );
  XNOR2_X1 U16943 ( .A(n15183), .B(n15182), .ZN(n15427) );
  OAI211_X1 U16944 ( .C1(n15186), .C2(n15185), .A(n15763), .B(n15184), .ZN(
        n15188) );
  NAND2_X1 U16945 ( .A1(n15188), .A2(n15187), .ZN(n15423) );
  INV_X1 U16946 ( .A(n15425), .ZN(n15195) );
  NAND2_X1 U16947 ( .A1(n15203), .A2(n15425), .ZN(n15189) );
  NAND2_X1 U16948 ( .A1(n15189), .A2(n15678), .ZN(n15190) );
  NOR2_X1 U16949 ( .A1(n15191), .A2(n15190), .ZN(n15424) );
  NAND2_X1 U16950 ( .A1(n15424), .A2(n15720), .ZN(n15194) );
  AOI22_X1 U16951 ( .A1(n15192), .A2(n15698), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n6546), .ZN(n15193) );
  OAI211_X1 U16952 ( .C1(n15195), .C2(n15367), .A(n15194), .B(n15193), .ZN(
        n15196) );
  AOI21_X1 U16953 ( .B1(n15423), .B2(n15714), .A(n15196), .ZN(n15197) );
  OAI21_X1 U16954 ( .B1(n15427), .B2(n15198), .A(n15197), .ZN(P1_U3269) );
  OAI21_X1 U16955 ( .B1(n15200), .B2(n13023), .A(n15199), .ZN(n15435) );
  XNOR2_X1 U16956 ( .A(n15202), .B(n15201), .ZN(n15433) );
  AOI21_X1 U16957 ( .B1(n15218), .B2(n15428), .A(n15733), .ZN(n15204) );
  NAND2_X1 U16958 ( .A1(n15204), .A2(n15203), .ZN(n15430) );
  AOI22_X1 U16959 ( .A1(n15205), .A2(n15698), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n6546), .ZN(n15206) );
  OAI21_X1 U16960 ( .B1(n15429), .B2(n6546), .A(n15206), .ZN(n15207) );
  AOI21_X1 U16961 ( .B1(n15428), .B2(n15716), .A(n15207), .ZN(n15208) );
  OAI21_X1 U16962 ( .B1(n15430), .B2(n15686), .A(n15208), .ZN(n15209) );
  AOI21_X1 U16963 ( .B1(n15433), .B2(n15295), .A(n15209), .ZN(n15210) );
  OAI21_X1 U16964 ( .B1(n15374), .B2(n15435), .A(n15210), .ZN(P1_U3270) );
  OAI21_X1 U16965 ( .B1(n15212), .B2(n15214), .A(n15211), .ZN(n15213) );
  INV_X1 U16966 ( .A(n15213), .ZN(n15440) );
  OAI21_X1 U16967 ( .B1(n8099), .B2(n13062), .A(n15215), .ZN(n15217) );
  AOI21_X1 U16968 ( .B1(n15217), .B2(n15763), .A(n15216), .ZN(n15439) );
  INV_X1 U16969 ( .A(n15439), .ZN(n15225) );
  AOI21_X1 U16970 ( .B1(n15231), .B2(n15437), .A(n15733), .ZN(n15219) );
  AND2_X1 U16971 ( .A1(n15219), .A2(n15218), .ZN(n15436) );
  NAND2_X1 U16972 ( .A1(n15436), .A2(n15720), .ZN(n15222) );
  AOI22_X1 U16973 ( .A1(n15220), .A2(n15698), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n6546), .ZN(n15221) );
  OAI211_X1 U16974 ( .C1(n15367), .C2(n15223), .A(n15222), .B(n15221), .ZN(
        n15224) );
  AOI21_X1 U16975 ( .B1(n15225), .B2(n15714), .A(n15224), .ZN(n15226) );
  OAI21_X1 U16976 ( .B1(n15440), .B2(n15374), .A(n15226), .ZN(P1_U3271) );
  XNOR2_X1 U16977 ( .A(n15228), .B(n15227), .ZN(n15445) );
  INV_X1 U16978 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n15230) );
  OAI22_X1 U16979 ( .A1(n15230), .A2(n15714), .B1(n15229), .B2(n15712), .ZN(
        n15241) );
  INV_X1 U16980 ( .A(n15254), .ZN(n15232) );
  AOI211_X1 U16981 ( .C1(n15443), .C2(n15232), .A(n15733), .B(n7992), .ZN(
        n15442) );
  OAI211_X1 U16982 ( .C1(n15235), .C2(n15234), .A(n15233), .B(n15763), .ZN(
        n15238) );
  INV_X1 U16983 ( .A(n15236), .ZN(n15237) );
  NAND2_X1 U16984 ( .A1(n15238), .A2(n15237), .ZN(n15441) );
  AOI21_X1 U16985 ( .B1(n15442), .B2(n15314), .A(n15441), .ZN(n15239) );
  NOR2_X1 U16986 ( .A1(n15239), .A2(n6546), .ZN(n15240) );
  AOI211_X1 U16987 ( .C1(n15716), .C2(n15443), .A(n15241), .B(n15240), .ZN(
        n15242) );
  OAI21_X1 U16988 ( .B1(n15445), .B2(n15374), .A(n15242), .ZN(P1_U3272) );
  OAI21_X1 U16989 ( .B1(n7955), .B2(n6682), .A(n15243), .ZN(n15451) );
  AND2_X1 U16990 ( .A1(n15281), .A2(n15244), .ZN(n15267) );
  NAND2_X1 U16991 ( .A1(n15267), .A2(n15266), .ZN(n15265) );
  AOI21_X1 U16992 ( .B1(n15265), .B2(n15246), .A(n15245), .ZN(n15249) );
  INV_X1 U16993 ( .A(n15247), .ZN(n15248) );
  NOR3_X1 U16994 ( .A1(n15249), .A2(n15709), .A3(n15248), .ZN(n15251) );
  NOR2_X1 U16995 ( .A1(n15251), .A2(n15250), .ZN(n15450) );
  INV_X1 U16996 ( .A(n15450), .ZN(n15261) );
  NOR2_X1 U16997 ( .A1(n15270), .A2(n15252), .ZN(n15253) );
  OR2_X1 U16998 ( .A1(n15254), .A2(n15253), .ZN(n15446) );
  INV_X1 U16999 ( .A(n15255), .ZN(n15256) );
  AOI22_X1 U17000 ( .A1(n15256), .A2(n15698), .B1(n6546), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n15258) );
  NAND2_X1 U17001 ( .A1(n15447), .A2(n15716), .ZN(n15257) );
  OAI211_X1 U17002 ( .C1(n15446), .C2(n15259), .A(n15258), .B(n15257), .ZN(
        n15260) );
  AOI21_X1 U17003 ( .B1(n15261), .B2(n15714), .A(n15260), .ZN(n15262) );
  OAI21_X1 U17004 ( .B1(n15374), .B2(n15451), .A(n15262), .ZN(P1_U3273) );
  XNOR2_X1 U17005 ( .A(n15263), .B(n15264), .ZN(n15458) );
  OAI21_X1 U17006 ( .B1(n15267), .B2(n15266), .A(n15265), .ZN(n15452) );
  NAND2_X1 U17007 ( .A1(n15285), .A2(n15455), .ZN(n15268) );
  NAND2_X1 U17008 ( .A1(n15268), .A2(n15678), .ZN(n15269) );
  NOR2_X1 U17009 ( .A1(n15270), .A2(n15269), .ZN(n15453) );
  NAND2_X1 U17010 ( .A1(n15453), .A2(n15720), .ZN(n15275) );
  OAI22_X1 U17011 ( .A1(n15714), .A2(n15272), .B1(n15271), .B2(n15712), .ZN(
        n15273) );
  AOI21_X1 U17012 ( .B1(n15454), .B2(n15714), .A(n15273), .ZN(n15274) );
  OAI211_X1 U17013 ( .C1(n15276), .C2(n15367), .A(n15275), .B(n15274), .ZN(
        n15277) );
  AOI21_X1 U17014 ( .B1(n15452), .B2(n15295), .A(n15277), .ZN(n15278) );
  OAI21_X1 U17015 ( .B1(n15458), .B2(n15374), .A(n15278), .ZN(P1_U3274) );
  XNOR2_X1 U17016 ( .A(n15279), .B(n15282), .ZN(n15463) );
  OAI211_X1 U17017 ( .C1(n15282), .C2(n15280), .A(n15281), .B(n15763), .ZN(
        n15284) );
  NAND2_X1 U17018 ( .A1(n15284), .A2(n15283), .ZN(n15459) );
  INV_X1 U17019 ( .A(n15461), .ZN(n15290) );
  AOI21_X1 U17020 ( .B1(n15298), .B2(n15461), .A(n15733), .ZN(n15286) );
  AND2_X1 U17021 ( .A1(n15286), .A2(n15285), .ZN(n15460) );
  NAND2_X1 U17022 ( .A1(n15460), .A2(n15720), .ZN(n15289) );
  AOI22_X1 U17023 ( .A1(n6546), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n15287), 
        .B2(n15698), .ZN(n15288) );
  OAI211_X1 U17024 ( .C1(n15290), .C2(n15367), .A(n15289), .B(n15288), .ZN(
        n15291) );
  AOI21_X1 U17025 ( .B1(n15459), .B2(n15714), .A(n15291), .ZN(n15292) );
  OAI21_X1 U17026 ( .B1(n15463), .B2(n15374), .A(n15292), .ZN(P1_U3275) );
  NAND2_X1 U17027 ( .A1(n6604), .A2(n15318), .ZN(n15311) );
  NAND2_X1 U17028 ( .A1(n15311), .A2(n15293), .ZN(n15294) );
  XOR2_X1 U17029 ( .A(n15296), .B(n15294), .Z(n15470) );
  INV_X1 U17030 ( .A(n15295), .ZN(n15355) );
  XOR2_X1 U17031 ( .A(n15297), .B(n15296), .Z(n15468) );
  OAI211_X1 U17032 ( .C1(n15299), .C2(n15466), .A(n15678), .B(n15298), .ZN(
        n15465) );
  AOI22_X1 U17033 ( .A1(n6546), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n15300), 
        .B2(n15698), .ZN(n15301) );
  OAI21_X1 U17034 ( .B1(n15464), .B2(n6546), .A(n15301), .ZN(n15302) );
  AOI21_X1 U17035 ( .B1(n15303), .B2(n15716), .A(n15302), .ZN(n15304) );
  OAI21_X1 U17036 ( .B1(n15465), .B2(n15686), .A(n15304), .ZN(n15305) );
  AOI21_X1 U17037 ( .B1(n15468), .B2(n15688), .A(n15305), .ZN(n15306) );
  OAI21_X1 U17038 ( .B1(n15470), .B2(n15355), .A(n15306), .ZN(P1_U3276) );
  XNOR2_X1 U17039 ( .A(n15330), .B(n15307), .ZN(n15310) );
  INV_X1 U17040 ( .A(n15308), .ZN(n15309) );
  OAI21_X1 U17041 ( .B1(n15310), .B2(n15733), .A(n15309), .ZN(n15471) );
  OAI21_X1 U17042 ( .B1(n6604), .B2(n15318), .A(n15311), .ZN(n15312) );
  NAND2_X1 U17043 ( .A1(n15312), .A2(n15763), .ZN(n15474) );
  INV_X1 U17044 ( .A(n15474), .ZN(n15313) );
  AOI21_X1 U17045 ( .B1(n15314), .B2(n15471), .A(n15313), .ZN(n15326) );
  OAI22_X1 U17046 ( .A1(n15714), .A2(n15316), .B1(n15315), .B2(n15712), .ZN(
        n15324) );
  NOR2_X1 U17047 ( .A1(n15371), .A2(n15317), .ZN(n15327) );
  OAI211_X1 U17048 ( .C1(n15327), .C2(n15320), .A(n15319), .B(n15318), .ZN(
        n15322) );
  AND2_X1 U17049 ( .A1(n15321), .A2(n15322), .ZN(n15475) );
  NOR2_X1 U17050 ( .A1(n15475), .A2(n15374), .ZN(n15323) );
  AOI211_X1 U17051 ( .C1(n15716), .C2(n15472), .A(n15324), .B(n15323), .ZN(
        n15325) );
  OAI21_X1 U17052 ( .B1(n15326), .B2(n6546), .A(n15325), .ZN(P1_U3277) );
  INV_X1 U17053 ( .A(n15327), .ZN(n15344) );
  NOR2_X1 U17054 ( .A1(n15344), .A2(n15345), .ZN(n15343) );
  NOR2_X1 U17055 ( .A1(n15343), .A2(n15328), .ZN(n15329) );
  XNOR2_X1 U17056 ( .A(n15329), .B(n15334), .ZN(n15482) );
  AOI211_X1 U17057 ( .C1(n15479), .C2(n15346), .A(n15733), .B(n15330), .ZN(
        n15477) );
  AOI22_X1 U17058 ( .A1(n6546), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n15331), 
        .B2(n15698), .ZN(n15332) );
  OAI21_X1 U17059 ( .B1(n7967), .B2(n15367), .A(n15332), .ZN(n15337) );
  OAI211_X1 U17060 ( .C1(n15335), .C2(n15334), .A(n15333), .B(n15763), .ZN(
        n15480) );
  AOI21_X1 U17061 ( .B1(n15480), .B2(n15476), .A(n6546), .ZN(n15336) );
  AOI211_X1 U17062 ( .C1(n15477), .C2(n15720), .A(n15337), .B(n15336), .ZN(
        n15338) );
  OAI21_X1 U17063 ( .B1(n15374), .B2(n15482), .A(n15338), .ZN(P1_U3278) );
  INV_X1 U17064 ( .A(n15339), .ZN(n15357) );
  NOR2_X1 U17065 ( .A1(n15357), .A2(n15370), .ZN(n15356) );
  NOR2_X1 U17066 ( .A1(n15356), .A2(n15340), .ZN(n15342) );
  XNOR2_X1 U17067 ( .A(n15342), .B(n15341), .ZN(n15489) );
  AOI21_X1 U17068 ( .B1(n15345), .B2(n15344), .A(n15343), .ZN(n15483) );
  AOI21_X1 U17069 ( .B1(n15361), .B2(n15486), .A(n15733), .ZN(n15347) );
  AND2_X1 U17070 ( .A1(n15347), .A2(n15346), .ZN(n15484) );
  NAND2_X1 U17071 ( .A1(n15484), .A2(n15720), .ZN(n15352) );
  OAI22_X1 U17072 ( .A1(n15714), .A2(n15349), .B1(n15348), .B2(n15712), .ZN(
        n15350) );
  AOI21_X1 U17073 ( .B1(n15714), .B2(n15485), .A(n15350), .ZN(n15351) );
  OAI211_X1 U17074 ( .C1(n7990), .C2(n15367), .A(n15352), .B(n15351), .ZN(
        n15353) );
  AOI21_X1 U17075 ( .B1(n15483), .B2(n15688), .A(n15353), .ZN(n15354) );
  OAI21_X1 U17076 ( .B1(n15489), .B2(n15355), .A(n15354), .ZN(P1_U3279) );
  AOI211_X1 U17077 ( .C1(n15370), .C2(n15357), .A(n15709), .B(n15356), .ZN(
        n15359) );
  NOR2_X1 U17078 ( .A1(n15359), .A2(n15358), .ZN(n15493) );
  INV_X1 U17079 ( .A(n15360), .ZN(n15363) );
  INV_X1 U17080 ( .A(n15361), .ZN(n15362) );
  AOI211_X1 U17081 ( .C1(n15491), .C2(n15363), .A(n15733), .B(n15362), .ZN(
        n15490) );
  INV_X1 U17082 ( .A(n15364), .ZN(n15365) );
  AOI22_X1 U17083 ( .A1(n6546), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n15365), 
        .B2(n15698), .ZN(n15366) );
  OAI21_X1 U17084 ( .B1(n15368), .B2(n15367), .A(n15366), .ZN(n15376) );
  INV_X1 U17085 ( .A(n15369), .ZN(n15373) );
  INV_X1 U17086 ( .A(n15370), .ZN(n15372) );
  AOI21_X1 U17087 ( .B1(n15373), .B2(n15372), .A(n15371), .ZN(n15494) );
  NOR2_X1 U17088 ( .A1(n15494), .A2(n15374), .ZN(n15375) );
  AOI211_X1 U17089 ( .C1(n15490), .C2(n15720), .A(n15376), .B(n15375), .ZN(
        n15377) );
  OAI21_X1 U17090 ( .B1(n15493), .B2(n6546), .A(n15377), .ZN(P1_U3280) );
  OAI211_X1 U17091 ( .C1(n15379), .C2(n15742), .A(n15378), .B(n15381), .ZN(
        n15521) );
  MUX2_X1 U17092 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15521), .S(n15804), .Z(
        P1_U3559) );
  NAND2_X1 U17093 ( .A1(n15380), .A2(n15678), .ZN(n15382) );
  OAI211_X1 U17094 ( .C1(n15383), .C2(n15742), .A(n15382), .B(n15381), .ZN(
        n15522) );
  MUX2_X1 U17095 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15522), .S(n15804), .Z(
        P1_U3558) );
  OAI21_X1 U17096 ( .B1(n15387), .B2(n15384), .A(n15763), .ZN(n15385) );
  NOR2_X1 U17097 ( .A1(n15385), .A2(n8098), .ZN(n15386) );
  NOR3_X1 U17098 ( .A1(n15389), .A2(n15388), .A3(n15387), .ZN(n15390) );
  OAI211_X1 U17099 ( .C1(n15394), .C2(n15742), .A(n15393), .B(n15392), .ZN(
        n15395) );
  MUX2_X1 U17100 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n15523), .S(n15804), .Z(
        P1_U3557) );
  OAI211_X1 U17101 ( .C1(n15400), .C2(n15742), .A(n15399), .B(n15398), .ZN(
        n15401) );
  MUX2_X1 U17102 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15524), .S(n15804), .Z(
        P1_U3556) );
  INV_X1 U17103 ( .A(n15770), .ZN(n15738) );
  OAI211_X1 U17104 ( .C1(n15407), .C2(n15742), .A(n15406), .B(n15405), .ZN(
        n15408) );
  INV_X1 U17105 ( .A(n15408), .ZN(n15409) );
  MUX2_X1 U17106 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15525), .S(n15804), .Z(
        P1_U3555) );
  OAI22_X1 U17107 ( .A1(n15411), .A2(n15733), .B1(n15410), .B2(n15742), .ZN(
        n15412) );
  INV_X1 U17108 ( .A(n15412), .ZN(n15413) );
  OAI211_X1 U17109 ( .C1(n15760), .C2(n15415), .A(n15414), .B(n15413), .ZN(
        n15526) );
  MUX2_X1 U17110 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15526), .S(n15804), .Z(
        P1_U3554) );
  OAI21_X1 U17111 ( .B1(n15417), .B2(n15742), .A(n15416), .ZN(n15418) );
  AOI211_X1 U17112 ( .C1(n15420), .C2(n15763), .A(n15419), .B(n15418), .ZN(
        n15421) );
  OAI21_X1 U17113 ( .B1(n15760), .B2(n15422), .A(n15421), .ZN(n15527) );
  MUX2_X1 U17114 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15527), .S(n15804), .Z(
        P1_U3553) );
  AOI211_X1 U17115 ( .C1(n15757), .C2(n15425), .A(n15424), .B(n15423), .ZN(
        n15426) );
  OAI21_X1 U17116 ( .B1(n15760), .B2(n15427), .A(n15426), .ZN(n15528) );
  MUX2_X1 U17117 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15528), .S(n15804), .Z(
        P1_U3552) );
  INV_X1 U17118 ( .A(n15428), .ZN(n15431) );
  OAI211_X1 U17119 ( .C1(n15431), .C2(n15742), .A(n15430), .B(n15429), .ZN(
        n15432) );
  AOI21_X1 U17120 ( .B1(n15433), .B2(n15763), .A(n15432), .ZN(n15434) );
  OAI21_X1 U17121 ( .B1(n15435), .B2(n15760), .A(n15434), .ZN(n15529) );
  MUX2_X1 U17122 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15529), .S(n15804), .Z(
        P1_U3551) );
  AOI21_X1 U17123 ( .B1(n15757), .B2(n15437), .A(n15436), .ZN(n15438) );
  OAI211_X1 U17124 ( .C1(n15760), .C2(n15440), .A(n15439), .B(n15438), .ZN(
        n15530) );
  MUX2_X1 U17125 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15530), .S(n15804), .Z(
        P1_U3550) );
  AOI211_X1 U17126 ( .C1(n15757), .C2(n15443), .A(n15442), .B(n15441), .ZN(
        n15444) );
  OAI21_X1 U17127 ( .B1(n15760), .B2(n15445), .A(n15444), .ZN(n15531) );
  MUX2_X1 U17128 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15531), .S(n15804), .Z(
        P1_U3549) );
  INV_X1 U17129 ( .A(n15446), .ZN(n15448) );
  AOI22_X1 U17130 ( .A1(n15448), .A2(n15678), .B1(n15757), .B2(n15447), .ZN(
        n15449) );
  OAI211_X1 U17131 ( .C1(n15760), .C2(n15451), .A(n15450), .B(n15449), .ZN(
        n15532) );
  MUX2_X1 U17132 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15532), .S(n15804), .Z(
        P1_U3548) );
  NAND2_X1 U17133 ( .A1(n15452), .A2(n15763), .ZN(n15457) );
  AOI211_X1 U17134 ( .C1(n15757), .C2(n15455), .A(n15454), .B(n15453), .ZN(
        n15456) );
  OAI211_X1 U17135 ( .C1(n15760), .C2(n15458), .A(n15457), .B(n15456), .ZN(
        n15533) );
  MUX2_X1 U17136 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15533), .S(n15804), .Z(
        P1_U3547) );
  AOI211_X1 U17137 ( .C1(n15757), .C2(n15461), .A(n15460), .B(n15459), .ZN(
        n15462) );
  OAI21_X1 U17138 ( .B1(n15760), .B2(n15463), .A(n15462), .ZN(n15534) );
  MUX2_X1 U17139 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15534), .S(n15804), .Z(
        P1_U3546) );
  INV_X1 U17140 ( .A(n15760), .ZN(n15783) );
  OAI211_X1 U17141 ( .C1(n15466), .C2(n15742), .A(n15465), .B(n15464), .ZN(
        n15467) );
  AOI21_X1 U17142 ( .B1(n15468), .B2(n15783), .A(n15467), .ZN(n15469) );
  OAI21_X1 U17143 ( .B1(n15470), .B2(n15709), .A(n15469), .ZN(n15535) );
  MUX2_X1 U17144 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15535), .S(n15804), .Z(
        P1_U3545) );
  AOI21_X1 U17145 ( .B1(n15757), .B2(n15472), .A(n15471), .ZN(n15473) );
  OAI211_X1 U17146 ( .C1(n15760), .C2(n15475), .A(n15474), .B(n15473), .ZN(
        n15536) );
  MUX2_X1 U17147 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15536), .S(n15804), .Z(
        P1_U3544) );
  INV_X1 U17148 ( .A(n15476), .ZN(n15478) );
  AOI211_X1 U17149 ( .C1(n15757), .C2(n15479), .A(n15478), .B(n15477), .ZN(
        n15481) );
  OAI211_X1 U17150 ( .C1(n15482), .C2(n15760), .A(n15481), .B(n15480), .ZN(
        n15537) );
  MUX2_X1 U17151 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15537), .S(n15804), .Z(
        P1_U3543) );
  NAND2_X1 U17152 ( .A1(n15483), .A2(n15783), .ZN(n15488) );
  AOI211_X1 U17153 ( .C1(n15757), .C2(n15486), .A(n15485), .B(n15484), .ZN(
        n15487) );
  OAI211_X1 U17154 ( .C1(n15709), .C2(n15489), .A(n15488), .B(n15487), .ZN(
        n15538) );
  MUX2_X1 U17155 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15538), .S(n15804), .Z(
        P1_U3542) );
  AOI21_X1 U17156 ( .B1(n15757), .B2(n15491), .A(n15490), .ZN(n15492) );
  OAI211_X1 U17157 ( .C1(n15760), .C2(n15494), .A(n15493), .B(n15492), .ZN(
        n15539) );
  MUX2_X1 U17158 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n15539), .S(n15804), .Z(
        P1_U3541) );
  AOI211_X1 U17159 ( .C1(n15757), .C2(n15497), .A(n15496), .B(n15495), .ZN(
        n15498) );
  OAI21_X1 U17160 ( .B1(n15760), .B2(n15499), .A(n15498), .ZN(n15540) );
  MUX2_X1 U17161 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n15540), .S(n15804), .Z(
        P1_U3540) );
  NAND2_X1 U17162 ( .A1(n15500), .A2(n15783), .ZN(n15502) );
  NAND4_X1 U17163 ( .A1(n15504), .A2(n15503), .A3(n15502), .A4(n15501), .ZN(
        n15541) );
  MUX2_X1 U17164 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n15541), .S(n15804), .Z(
        P1_U3539) );
  NOR4_X1 U17165 ( .A1(n15508), .A2(n15507), .A3(n15506), .A4(n15505), .ZN(
        n15509) );
  OAI21_X1 U17166 ( .B1(n15760), .B2(n15510), .A(n15509), .ZN(n15542) );
  MUX2_X1 U17167 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n15542), .S(n15804), .Z(
        P1_U3538) );
  NOR4_X1 U17168 ( .A1(n15514), .A2(n15513), .A3(n15512), .A4(n15511), .ZN(
        n15515) );
  OAI21_X1 U17169 ( .B1(n15760), .B2(n15516), .A(n15515), .ZN(n15543) );
  MUX2_X1 U17170 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n15543), .S(n15804), .Z(
        P1_U3537) );
  NOR2_X1 U17171 ( .A1(n15518), .A2(n15517), .ZN(n15520) );
  MUX2_X1 U17172 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n15521), .S(n15791), .Z(
        P1_U3527) );
  MUX2_X1 U17173 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15522), .S(n15791), .Z(
        P1_U3526) );
  MUX2_X1 U17174 ( .A(n15525), .B(P1_REG0_REG_27__SCAN_IN), .S(n15789), .Z(
        P1_U3523) );
  MUX2_X1 U17175 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15526), .S(n15791), .Z(
        P1_U3522) );
  MUX2_X1 U17176 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15527), .S(n15791), .Z(
        P1_U3521) );
  MUX2_X1 U17177 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15528), .S(n15791), .Z(
        P1_U3520) );
  MUX2_X1 U17178 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15529), .S(n15791), .Z(
        P1_U3519) );
  MUX2_X1 U17179 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15530), .S(n15791), .Z(
        P1_U3518) );
  MUX2_X1 U17180 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15531), .S(n15791), .Z(
        P1_U3517) );
  MUX2_X1 U17181 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15532), .S(n15791), .Z(
        P1_U3516) );
  MUX2_X1 U17182 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15533), .S(n15791), .Z(
        P1_U3515) );
  MUX2_X1 U17183 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15534), .S(n15791), .Z(
        P1_U3513) );
  MUX2_X1 U17184 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15535), .S(n15791), .Z(
        P1_U3510) );
  MUX2_X1 U17185 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15536), .S(n15791), .Z(
        P1_U3507) );
  MUX2_X1 U17186 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15537), .S(n15791), .Z(
        P1_U3504) );
  MUX2_X1 U17187 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n15538), .S(n15791), .Z(
        P1_U3501) );
  MUX2_X1 U17188 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n15539), .S(n15791), .Z(
        P1_U3498) );
  MUX2_X1 U17189 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n15540), .S(n15791), .Z(
        P1_U3495) );
  MUX2_X1 U17190 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n15541), .S(n15791), .Z(
        P1_U3492) );
  MUX2_X1 U17191 ( .A(P1_REG0_REG_10__SCAN_IN), .B(n15542), .S(n15791), .Z(
        P1_U3489) );
  MUX2_X1 U17192 ( .A(P1_REG0_REG_9__SCAN_IN), .B(n15543), .S(n15791), .Z(
        P1_U3486) );
  NAND3_X1 U17193 ( .A1(n15545), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n15548) );
  OAI22_X1 U17194 ( .A1(n15544), .A2(n15548), .B1(n15547), .B2(n15546), .ZN(
        n15549) );
  AOI21_X1 U17195 ( .B1(n12735), .B2(n15550), .A(n15549), .ZN(n15551) );
  INV_X1 U17196 ( .A(n15551), .ZN(P1_U3324) );
  MUX2_X1 U17197 ( .A(n6809), .B(n15552), .S(P1_U3086), .Z(P1_U3333) );
  XOR2_X1 U17198 ( .A(n15554), .B(n15555), .Z(SUB_1596_U57) );
  XOR2_X1 U17199 ( .A(n15556), .B(n15557), .Z(SUB_1596_U56) );
  XOR2_X1 U17200 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n15558), .Z(SUB_1596_U54) );
  NAND2_X1 U17201 ( .A1(n15562), .A2(n15559), .ZN(n15561) );
  NAND2_X1 U17202 ( .A1(n15561), .A2(n15560), .ZN(n15565) );
  INV_X1 U17203 ( .A(n15562), .ZN(n15563) );
  NAND2_X1 U17204 ( .A1(n15563), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n15564) );
  NAND2_X1 U17205 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n15566), .ZN(n15567) );
  NAND2_X1 U17206 ( .A1(n15568), .A2(n15567), .ZN(n15571) );
  INV_X1 U17207 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n15569) );
  NAND2_X1 U17208 ( .A1(n15569), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n15570) );
  NAND2_X1 U17209 ( .A1(n15571), .A2(n15570), .ZN(n15578) );
  INV_X1 U17210 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15579) );
  XNOR2_X1 U17211 ( .A(n15579), .B(P1_ADDR_REG_14__SCAN_IN), .ZN(n15577) );
  XNOR2_X1 U17212 ( .A(n15578), .B(n15577), .ZN(n15572) );
  INV_X1 U17213 ( .A(n15576), .ZN(n15573) );
  NAND2_X1 U17214 ( .A1(n15573), .A2(n15575), .ZN(n15574) );
  XNOR2_X1 U17215 ( .A(n15574), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  NAND2_X1 U17216 ( .A1(n15579), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n15580) );
  XNOR2_X1 U17217 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .ZN(n15582) );
  XNOR2_X1 U17218 ( .A(n15590), .B(n15582), .ZN(n15585) );
  XNOR2_X1 U17219 ( .A(n15585), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(n15583) );
  XNOR2_X1 U17220 ( .A(n15584), .B(n15583), .ZN(SUB_1596_U65) );
  INV_X1 U17221 ( .A(n15585), .ZN(n15587) );
  INV_X1 U17222 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15669) );
  NOR2_X1 U17223 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n15669), .ZN(n15589) );
  OAI22_X1 U17224 ( .A1(n15590), .A2(n15589), .B1(P1_ADDR_REG_15__SCAN_IN), 
        .B2(n15588), .ZN(n15600) );
  XNOR2_X1 U17225 ( .A(n15601), .B(P1_ADDR_REG_16__SCAN_IN), .ZN(n15591) );
  XNOR2_X1 U17226 ( .A(n15600), .B(n15591), .ZN(n15592) );
  INV_X1 U17227 ( .A(n15597), .ZN(n15594) );
  NAND2_X1 U17228 ( .A1(n15594), .A2(n15596), .ZN(n15595) );
  XNOR2_X1 U17229 ( .A(n15595), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  AND2_X1 U17230 ( .A1(n15598), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n15599) );
  OR2_X1 U17231 ( .A1(n15600), .A2(n15599), .ZN(n15603) );
  NAND2_X1 U17232 ( .A1(n15601), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n15602) );
  NAND2_X1 U17233 ( .A1(n15603), .A2(n15602), .ZN(n15609) );
  XNOR2_X1 U17234 ( .A(n15609), .B(P1_ADDR_REG_17__SCAN_IN), .ZN(n15608) );
  XNOR2_X1 U17235 ( .A(n15608), .B(P3_ADDR_REG_17__SCAN_IN), .ZN(n15604) );
  NAND2_X1 U17236 ( .A1(n6635), .A2(n15607), .ZN(n15606) );
  XNOR2_X1 U17237 ( .A(n15606), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  INV_X1 U17238 ( .A(n15608), .ZN(n15611) );
  NOR2_X1 U17239 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n15609), .ZN(n15610) );
  AOI21_X1 U17240 ( .B1(n15611), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n15610), 
        .ZN(n15621) );
  XNOR2_X1 U17241 ( .A(P1_ADDR_REG_18__SCAN_IN), .B(P3_ADDR_REG_18__SCAN_IN), 
        .ZN(n15612) );
  XNOR2_X1 U17242 ( .A(n15621), .B(n15612), .ZN(n15613) );
  AOI21_X1 U17243 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n15614), .A(n15618), 
        .ZN(n15615) );
  INV_X1 U17244 ( .A(n15615), .ZN(SUB_1596_U62) );
  INV_X1 U17245 ( .A(n15616), .ZN(n15617) );
  AND2_X1 U17246 ( .A1(n15619), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n15620) );
  OAI22_X1 U17247 ( .A1(n15621), .A2(n15620), .B1(P1_ADDR_REG_18__SCAN_IN), 
        .B2(n15619), .ZN(n15624) );
  XNOR2_X1 U17248 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n15622) );
  XNOR2_X1 U17249 ( .A(n15622), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n15623) );
  XNOR2_X1 U17250 ( .A(n15624), .B(n15623), .ZN(n15625) );
  AOI21_X1 U17251 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15626) );
  OAI21_X1 U17252 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n15626), 
        .ZN(U28) );
  AND2_X1 U17253 ( .A1(n15628), .A2(n15627), .ZN(n15630) );
  XNOR2_X1 U17254 ( .A(n15630), .B(n15629), .ZN(SUB_1596_U61) );
  NOR2_X1 U17255 ( .A1(n15631), .A2(n15742), .ZN(n15749) );
  AOI22_X1 U17256 ( .A1(n15632), .A2(n15749), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15645) );
  AOI21_X1 U17257 ( .B1(n15633), .B2(n15635), .A(n15634), .ZN(n15643) );
  NAND2_X1 U17258 ( .A1(n6540), .A2(n15636), .ZN(n15640) );
  NAND2_X1 U17259 ( .A1(n15638), .A2(n15637), .ZN(n15639) );
  NAND2_X1 U17260 ( .A1(n15640), .A2(n15639), .ZN(n15748) );
  AOI22_X1 U17261 ( .A1(n15643), .A2(n15642), .B1(n15641), .B2(n15748), .ZN(
        n15644) );
  OAI211_X1 U17262 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n15646), .A(n15645), .B(
        n15644), .ZN(P1_U3218) );
  AOI21_X1 U17263 ( .B1(n7374), .B2(n15648), .A(n15647), .ZN(n15650) );
  XNOR2_X1 U17264 ( .A(n15650), .B(P1_IR_REG_0__SCAN_IN), .ZN(n15653) );
  AOI22_X1 U17265 ( .A1(n15651), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n15652) );
  OAI21_X1 U17266 ( .B1(n15654), .B2(n15653), .A(n15652), .ZN(P1_U3243) );
  XNOR2_X1 U17267 ( .A(n15656), .B(n15655), .ZN(n15664) );
  AOI21_X1 U17268 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n15658), .A(n15657), 
        .ZN(n15662) );
  OAI22_X1 U17269 ( .A1(n15662), .A2(n15661), .B1(n15660), .B2(n15659), .ZN(
        n15663) );
  AOI21_X1 U17270 ( .B1(n15665), .B2(n15664), .A(n15663), .ZN(n15667) );
  OAI211_X1 U17271 ( .C1(n15669), .C2(n15668), .A(n15667), .B(n15666), .ZN(
        P1_U3258) );
  XNOR2_X1 U17272 ( .A(n15670), .B(n7700), .ZN(n15673) );
  AOI21_X1 U17273 ( .B1(n15673), .B2(n15763), .A(n15672), .ZN(n15788) );
  OAI21_X1 U17274 ( .B1(n15676), .B2(n15675), .A(n15674), .ZN(n15784) );
  INV_X1 U17275 ( .A(n15684), .ZN(n15680) );
  INV_X1 U17276 ( .A(n15677), .ZN(n15700) );
  OAI211_X1 U17277 ( .C1(n15680), .C2(n15700), .A(n15679), .B(n15678), .ZN(
        n15785) );
  OAI22_X1 U17278 ( .A1(n15714), .A2(n15682), .B1(n15681), .B2(n15712), .ZN(
        n15683) );
  AOI21_X1 U17279 ( .B1(n15716), .B2(n15684), .A(n15683), .ZN(n15685) );
  OAI21_X1 U17280 ( .B1(n15785), .B2(n15686), .A(n15685), .ZN(n15687) );
  AOI21_X1 U17281 ( .B1(n15784), .B2(n15688), .A(n15687), .ZN(n15689) );
  OAI21_X1 U17282 ( .B1(n6546), .B2(n15788), .A(n15689), .ZN(P1_U3285) );
  OAI21_X1 U17283 ( .B1(n15691), .B2(n15694), .A(n15690), .ZN(n15782) );
  NAND2_X1 U17284 ( .A1(n15693), .A2(n15692), .ZN(n15695) );
  XNOR2_X1 U17285 ( .A(n15695), .B(n15694), .ZN(n15696) );
  NOR2_X1 U17286 ( .A1(n15696), .A2(n15709), .ZN(n15780) );
  AOI211_X1 U17287 ( .C1(n15711), .C2(n15782), .A(n15777), .B(n15780), .ZN(
        n15705) );
  INV_X1 U17288 ( .A(n15697), .ZN(n15699) );
  AOI222_X1 U17289 ( .A1(n15702), .A2(n15716), .B1(P1_REG2_REG_7__SCAN_IN), 
        .B2(n6546), .C1(n15699), .C2(n15698), .ZN(n15704) );
  AOI211_X1 U17290 ( .C1(n15702), .C2(n15701), .A(n15733), .B(n15700), .ZN(
        n15779) );
  AOI22_X1 U17291 ( .A1(n15782), .A2(n15719), .B1(n15779), .B2(n15720), .ZN(
        n15703) );
  OAI211_X1 U17292 ( .C1(n6546), .C2(n15705), .A(n15704), .B(n15703), .ZN(
        P1_U3286) );
  XNOR2_X1 U17293 ( .A(n15708), .B(n15706), .ZN(n15753) );
  XNOR2_X1 U17294 ( .A(n15708), .B(n15707), .ZN(n15710) );
  NOR2_X1 U17295 ( .A1(n15710), .A2(n15709), .ZN(n15751) );
  AOI211_X1 U17296 ( .C1(n15711), .C2(n15753), .A(n15748), .B(n15751), .ZN(
        n15723) );
  OAI22_X1 U17297 ( .A1(n15714), .A2(n15713), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n15712), .ZN(n15715) );
  AOI21_X1 U17298 ( .B1(n15716), .B2(n7771), .A(n15715), .ZN(n15722) );
  AOI211_X1 U17299 ( .C1(n7771), .C2(n15718), .A(n15733), .B(n15717), .ZN(
        n15750) );
  AOI22_X1 U17300 ( .A1(n15720), .A2(n15750), .B1(n15753), .B2(n15719), .ZN(
        n15721) );
  OAI211_X1 U17301 ( .C1(n6546), .C2(n15723), .A(n15722), .B(n15721), .ZN(
        P1_U3290) );
  AND2_X1 U17302 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15729), .ZN(P1_U3294) );
  INV_X1 U17303 ( .A(n15729), .ZN(n15728) );
  NOR2_X1 U17304 ( .A1(n15728), .A2(n15724), .ZN(P1_U3295) );
  AND2_X1 U17305 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15729), .ZN(P1_U3296) );
  AND2_X1 U17306 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15729), .ZN(P1_U3297) );
  AND2_X1 U17307 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15729), .ZN(P1_U3298) );
  AND2_X1 U17308 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15729), .ZN(P1_U3299) );
  AND2_X1 U17309 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15729), .ZN(P1_U3300) );
  AND2_X1 U17310 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15729), .ZN(P1_U3301) );
  AND2_X1 U17311 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15729), .ZN(P1_U3302) );
  AND2_X1 U17312 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15729), .ZN(P1_U3303) );
  AND2_X1 U17313 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15729), .ZN(P1_U3304) );
  NOR2_X1 U17314 ( .A1(n15728), .A2(n15725), .ZN(P1_U3305) );
  NOR2_X1 U17315 ( .A1(n15728), .A2(n15726), .ZN(P1_U3306) );
  AND2_X1 U17316 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15729), .ZN(P1_U3307) );
  AND2_X1 U17317 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15729), .ZN(P1_U3308) );
  AND2_X1 U17318 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15729), .ZN(P1_U3309) );
  AND2_X1 U17319 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15729), .ZN(P1_U3310) );
  AND2_X1 U17320 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15729), .ZN(P1_U3311) );
  AND2_X1 U17321 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15729), .ZN(P1_U3312) );
  AND2_X1 U17322 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15729), .ZN(P1_U3313) );
  AND2_X1 U17323 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15729), .ZN(P1_U3314) );
  AND2_X1 U17324 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15729), .ZN(P1_U3315) );
  AND2_X1 U17325 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15729), .ZN(P1_U3316) );
  NOR2_X1 U17326 ( .A1(n15728), .A2(n15727), .ZN(P1_U3317) );
  AND2_X1 U17327 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15729), .ZN(P1_U3318) );
  AND2_X1 U17328 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15729), .ZN(P1_U3319) );
  AND2_X1 U17329 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15729), .ZN(P1_U3320) );
  AND2_X1 U17330 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15729), .ZN(P1_U3321) );
  AND2_X1 U17331 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15729), .ZN(P1_U3322) );
  AND2_X1 U17332 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15729), .ZN(P1_U3323) );
  INV_X1 U17333 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15730) );
  AOI22_X1 U17334 ( .A1(n15791), .A2(n15731), .B1(n15730), .B2(n15789), .ZN(
        P1_U3459) );
  OAI22_X1 U17335 ( .A1(n15734), .A2(n15733), .B1(n15732), .B2(n15742), .ZN(
        n15736) );
  AOI211_X1 U17336 ( .C1(n15738), .C2(n15737), .A(n15736), .B(n15735), .ZN(
        n15792) );
  INV_X1 U17337 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n15739) );
  AOI22_X1 U17338 ( .A1(n15791), .A2(n15792), .B1(n15739), .B2(n15789), .ZN(
        P1_U3462) );
  OAI211_X1 U17339 ( .C1(n15743), .C2(n15742), .A(n15741), .B(n15740), .ZN(
        n15747) );
  AOI21_X1 U17340 ( .B1(n15745), .B2(n15770), .A(n15744), .ZN(n15746) );
  NOR2_X1 U17341 ( .A1(n15747), .A2(n15746), .ZN(n15793) );
  AOI22_X1 U17342 ( .A1(n15791), .A2(n15793), .B1(n9489), .B2(n15789), .ZN(
        P1_U3465) );
  OR4_X1 U17343 ( .A1(n15751), .A2(n15750), .A3(n15749), .A4(n15748), .ZN(
        n15752) );
  AOI21_X1 U17344 ( .B1(n15783), .B2(n15753), .A(n15752), .ZN(n15794) );
  AOI22_X1 U17345 ( .A1(n15791), .A2(n15794), .B1(n9508), .B2(n15789), .ZN(
        P1_U3468) );
  AOI211_X1 U17346 ( .C1(n15757), .C2(n15756), .A(n15755), .B(n15754), .ZN(
        n15758) );
  OAI21_X1 U17347 ( .B1(n15760), .B2(n15759), .A(n15758), .ZN(n15761) );
  AOI21_X1 U17348 ( .B1(n15763), .B2(n15762), .A(n15761), .ZN(n15796) );
  AOI22_X1 U17349 ( .A1(n15791), .A2(n15796), .B1(n9525), .B2(n15789), .ZN(
        P1_U3471) );
  OAI211_X1 U17350 ( .C1(n15766), .C2(n15770), .A(n15765), .B(n15764), .ZN(
        n15767) );
  NOR2_X1 U17351 ( .A1(n15768), .A2(n15767), .ZN(n15798) );
  INV_X1 U17352 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15769) );
  AOI22_X1 U17353 ( .A1(n15791), .A2(n15798), .B1(n15769), .B2(n15789), .ZN(
        P1_U3474) );
  NOR2_X1 U17354 ( .A1(n15771), .A2(n15770), .ZN(n15774) );
  NOR4_X1 U17355 ( .A1(n15775), .A2(n15774), .A3(n15773), .A4(n15772), .ZN(
        n15799) );
  INV_X1 U17356 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n15776) );
  AOI22_X1 U17357 ( .A1(n15791), .A2(n15799), .B1(n15776), .B2(n15789), .ZN(
        P1_U3477) );
  OR3_X1 U17358 ( .A1(n15779), .A2(n15778), .A3(n15777), .ZN(n15781) );
  AOI211_X1 U17359 ( .C1(n15783), .C2(n15782), .A(n15781), .B(n15780), .ZN(
        n15801) );
  AOI22_X1 U17360 ( .A1(n15791), .A2(n15801), .B1(n9590), .B2(n15789), .ZN(
        P1_U3480) );
  NAND2_X1 U17361 ( .A1(n15784), .A2(n15783), .ZN(n15786) );
  INV_X1 U17362 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15790) );
  AOI22_X1 U17363 ( .A1(n15791), .A2(n15803), .B1(n15790), .B2(n15789), .ZN(
        P1_U3483) );
  AOI22_X1 U17364 ( .A1(n15804), .A2(n15792), .B1(n9457), .B2(n15802), .ZN(
        P1_U3529) );
  AOI22_X1 U17365 ( .A1(n15804), .A2(n15793), .B1(n9487), .B2(n15802), .ZN(
        P1_U3530) );
  AOI22_X1 U17366 ( .A1(n15804), .A2(n15794), .B1(n10574), .B2(n15802), .ZN(
        P1_U3531) );
  AOI22_X1 U17367 ( .A1(n15804), .A2(n15796), .B1(n15795), .B2(n15802), .ZN(
        P1_U3532) );
  AOI22_X1 U17368 ( .A1(n15804), .A2(n15798), .B1(n15797), .B2(n15802), .ZN(
        P1_U3533) );
  AOI22_X1 U17369 ( .A1(n15804), .A2(n15799), .B1(n15001), .B2(n15802), .ZN(
        P1_U3534) );
  AOI22_X1 U17370 ( .A1(n15804), .A2(n15801), .B1(n15800), .B2(n15802), .ZN(
        P1_U3535) );
  AOI22_X1 U17371 ( .A1(n15804), .A2(n15803), .B1(n9609), .B2(n15802), .ZN(
        P1_U3536) );
  NOR2_X1 U17372 ( .A1(n15809), .A2(P2_U3947), .ZN(P2_U3087) );
  NOR2_X1 U17373 ( .A1(n15806), .A2(n15805), .ZN(n15807) );
  AOI211_X1 U17374 ( .C1(n15809), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n15808), .B(
        n15807), .ZN(n15820) );
  OAI211_X1 U17375 ( .C1(n15813), .C2(n15812), .A(n15811), .B(n15810), .ZN(
        n15819) );
  OAI211_X1 U17376 ( .C1(n15817), .C2(n15816), .A(n15815), .B(n15814), .ZN(
        n15818) );
  NAND3_X1 U17377 ( .A1(n15820), .A2(n15819), .A3(n15818), .ZN(P2_U3218) );
  INV_X1 U17378 ( .A(n15821), .ZN(n15829) );
  OR2_X1 U17379 ( .A1(n15823), .A2(n15822), .ZN(n15826) );
  AOI211_X1 U17380 ( .C1(n15827), .C2(n15826), .A(n15825), .B(n15824), .ZN(
        n15828) );
  AOI211_X1 U17381 ( .C1(n15831), .C2(n15830), .A(n15829), .B(n15828), .ZN(
        n15838) );
  AOI21_X1 U17382 ( .B1(n15834), .B2(n15833), .A(n15832), .ZN(n15836) );
  NAND2_X1 U17383 ( .A1(n15836), .A2(n15835), .ZN(n15837) );
  OAI211_X1 U17384 ( .C1(n15840), .C2(n15839), .A(n15838), .B(n15837), .ZN(
        P2_U3224) );
  INV_X1 U17385 ( .A(n15841), .ZN(n15845) );
  OAI22_X1 U17386 ( .A1(n15845), .A2(n15844), .B1(n15843), .B2(n15842), .ZN(
        n15847) );
  AOI211_X1 U17387 ( .C1(n15849), .C2(n15848), .A(n15847), .B(n15846), .ZN(
        n15851) );
  AOI22_X1 U17388 ( .A1(n14499), .A2(n10747), .B1(n15851), .B2(n15850), .ZN(
        P2_U3265) );
  INV_X1 U17389 ( .A(n15864), .ZN(n15861) );
  AND2_X1 U17390 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15858), .ZN(P2_U3266) );
  AND2_X1 U17391 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15858), .ZN(P2_U3267) );
  NOR2_X1 U17392 ( .A1(n15857), .A2(n15853), .ZN(P2_U3268) );
  AND2_X1 U17393 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15858), .ZN(P2_U3269) );
  AND2_X1 U17394 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15858), .ZN(P2_U3270) );
  AND2_X1 U17395 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15858), .ZN(P2_U3271) );
  AND2_X1 U17396 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15858), .ZN(P2_U3272) );
  AND2_X1 U17397 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15858), .ZN(P2_U3273) );
  AND2_X1 U17398 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15858), .ZN(P2_U3274) );
  NOR2_X1 U17399 ( .A1(n15857), .A2(n15854), .ZN(P2_U3275) );
  AND2_X1 U17400 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15858), .ZN(P2_U3276) );
  AND2_X1 U17401 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15858), .ZN(P2_U3277) );
  AND2_X1 U17402 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15858), .ZN(P2_U3278) );
  AND2_X1 U17403 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15858), .ZN(P2_U3279) );
  AND2_X1 U17404 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15858), .ZN(P2_U3280) );
  AND2_X1 U17405 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15858), .ZN(P2_U3281) );
  AND2_X1 U17406 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15858), .ZN(P2_U3282) );
  AND2_X1 U17407 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15858), .ZN(P2_U3283) );
  AND2_X1 U17408 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15858), .ZN(P2_U3284) );
  AND2_X1 U17409 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15858), .ZN(P2_U3285) );
  AND2_X1 U17410 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15858), .ZN(P2_U3286) );
  AND2_X1 U17411 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15858), .ZN(P2_U3287) );
  AND2_X1 U17412 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15858), .ZN(P2_U3288) );
  AND2_X1 U17413 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15858), .ZN(P2_U3289) );
  NOR2_X1 U17414 ( .A1(n15857), .A2(n15855), .ZN(P2_U3290) );
  NOR2_X1 U17415 ( .A1(n15857), .A2(n15856), .ZN(P2_U3291) );
  AND2_X1 U17416 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15858), .ZN(P2_U3292) );
  AND2_X1 U17417 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15858), .ZN(P2_U3293) );
  AND2_X1 U17418 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15858), .ZN(P2_U3294) );
  AND2_X1 U17419 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15858), .ZN(P2_U3295) );
  AOI22_X1 U17420 ( .A1(n15864), .A2(n15860), .B1(n15859), .B2(n15861), .ZN(
        P2_U3416) );
  AOI22_X1 U17421 ( .A1(n15864), .A2(n15863), .B1(n15862), .B2(n15861), .ZN(
        P2_U3417) );
  AOI22_X1 U17422 ( .A1(n15886), .A2(n15865), .B1(n7438), .B2(n15885), .ZN(
        P2_U3430) );
  OAI21_X1 U17423 ( .B1(n15867), .B2(n15879), .A(n15866), .ZN(n15869) );
  AOI211_X1 U17424 ( .C1(n15877), .C2(n15870), .A(n15869), .B(n15868), .ZN(
        n15888) );
  AOI22_X1 U17425 ( .A1(n15886), .A2(n15888), .B1(n8840), .B2(n15885), .ZN(
        P2_U3436) );
  INV_X1 U17426 ( .A(n15871), .ZN(n15872) );
  OAI21_X1 U17427 ( .B1(n15873), .B2(n15879), .A(n15872), .ZN(n15874) );
  AOI211_X1 U17428 ( .C1(n15877), .C2(n15876), .A(n15875), .B(n15874), .ZN(
        n15889) );
  AOI22_X1 U17429 ( .A1(n15886), .A2(n15889), .B1(n8869), .B2(n15885), .ZN(
        P2_U3442) );
  OAI21_X1 U17430 ( .B1(n15880), .B2(n15879), .A(n15878), .ZN(n15882) );
  AOI211_X1 U17431 ( .C1(n15884), .C2(n15883), .A(n15882), .B(n15881), .ZN(
        n15892) );
  AOI22_X1 U17432 ( .A1(n15886), .A2(n15892), .B1(n8852), .B2(n15885), .ZN(
        P2_U3445) );
  AOI22_X1 U17433 ( .A1(n15893), .A2(n15888), .B1(n15887), .B2(n15890), .ZN(
        P2_U3501) );
  AOI22_X1 U17434 ( .A1(n15893), .A2(n15889), .B1(n10622), .B2(n15890), .ZN(
        P2_U3503) );
  AOI22_X1 U17435 ( .A1(n15893), .A2(n15892), .B1(n15891), .B2(n15890), .ZN(
        P2_U3504) );
  NOR2_X1 U17436 ( .A1(P3_U3897), .A2(n15894), .ZN(P3_U3150) );
  OAI22_X1 U17437 ( .A1(n15898), .A2(n15897), .B1(n15896), .B2(n15895), .ZN(
        n15899) );
  AOI211_X1 U17438 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n15901), .A(n15900), .B(
        n15899), .ZN(n15902) );
  AOI22_X1 U17439 ( .A1(n15903), .A2(n10092), .B1(n15902), .B2(n15921), .ZN(
        P3_U3231) );
  XNOR2_X1 U17440 ( .A(n15904), .B(n11594), .ZN(n15924) );
  NOR2_X1 U17441 ( .A1(n15948), .A2(n15905), .ZN(n15926) );
  INV_X1 U17442 ( .A(n15906), .ZN(n15913) );
  INV_X1 U17443 ( .A(n11594), .ZN(n15909) );
  INV_X1 U17444 ( .A(n15907), .ZN(n15908) );
  AOI21_X1 U17445 ( .B1(n15910), .B2(n15909), .A(n15908), .ZN(n15912) );
  OAI222_X1 U17446 ( .A1(n15916), .A2(n15915), .B1(n15914), .B2(n15913), .C1(
        n15912), .C2(n15911), .ZN(n15925) );
  AOI21_X1 U17447 ( .B1(n15926), .B2(n15917), .A(n15925), .ZN(n15918) );
  OAI211_X1 U17448 ( .C1(n15919), .C2(n15924), .A(n15921), .B(n15918), .ZN(
        n15920) );
  OAI21_X1 U17449 ( .B1(P3_REG2_REG_1__SCAN_IN), .B2(n15921), .A(n15920), .ZN(
        n15922) );
  OAI21_X1 U17450 ( .B1(n11609), .B2(n15923), .A(n15922), .ZN(P3_U3232) );
  INV_X1 U17451 ( .A(n15924), .ZN(n15927) );
  AOI211_X1 U17452 ( .C1(n15928), .C2(n15927), .A(n15926), .B(n15925), .ZN(
        n15962) );
  AOI22_X1 U17453 ( .A1(n15960), .A2(n8137), .B1(n15962), .B2(n15959), .ZN(
        P3_U3393) );
  AOI22_X1 U17454 ( .A1(n15960), .A2(n8146), .B1(n15929), .B2(n15959), .ZN(
        P3_U3396) );
  INV_X1 U17455 ( .A(n15930), .ZN(n15931) );
  AOI211_X1 U17456 ( .C1(n15933), .C2(n15957), .A(n15932), .B(n15931), .ZN(
        n15964) );
  AOI22_X1 U17457 ( .A1(n15960), .A2(n8155), .B1(n15964), .B2(n15959), .ZN(
        P3_U3399) );
  INV_X1 U17458 ( .A(n15934), .ZN(n15938) );
  INV_X1 U17459 ( .A(n15935), .ZN(n15936) );
  AOI211_X1 U17460 ( .C1(n15957), .C2(n15938), .A(n15937), .B(n15936), .ZN(
        n15966) );
  AOI22_X1 U17461 ( .A1(n15960), .A2(n8167), .B1(n15966), .B2(n15959), .ZN(
        P3_U3402) );
  INV_X1 U17462 ( .A(n15939), .ZN(n15940) );
  AOI211_X1 U17463 ( .C1(n15942), .C2(n15957), .A(n15941), .B(n15940), .ZN(
        n15968) );
  AOI22_X1 U17464 ( .A1(n15960), .A2(n8183), .B1(n15968), .B2(n15959), .ZN(
        P3_U3405) );
  AOI22_X1 U17465 ( .A1(n15945), .A2(n15957), .B1(n15944), .B2(n15943), .ZN(
        n15946) );
  AND2_X1 U17466 ( .A1(n15947), .A2(n15946), .ZN(n15970) );
  AOI22_X1 U17467 ( .A1(n15960), .A2(n8200), .B1(n15970), .B2(n15959), .ZN(
        P3_U3408) );
  OAI22_X1 U17468 ( .A1(n15951), .A2(n15950), .B1(n15949), .B2(n15948), .ZN(
        n15952) );
  NOR2_X1 U17469 ( .A1(n15953), .A2(n15952), .ZN(n15972) );
  AOI22_X1 U17470 ( .A1(n15960), .A2(n8218), .B1(n15972), .B2(n15959), .ZN(
        P3_U3411) );
  INV_X1 U17471 ( .A(n15954), .ZN(n15955) );
  AOI211_X1 U17472 ( .C1(n15958), .C2(n15957), .A(n15956), .B(n15955), .ZN(
        n15975) );
  AOI22_X1 U17473 ( .A1(n15960), .A2(n8243), .B1(n15975), .B2(n15959), .ZN(
        P3_U3414) );
  AOI22_X1 U17474 ( .A1(n15976), .A2(n15962), .B1(n15961), .B2(n15973), .ZN(
        P3_U3460) );
  AOI22_X1 U17475 ( .A1(n15976), .A2(n15964), .B1(n15963), .B2(n15973), .ZN(
        P3_U3462) );
  AOI22_X1 U17476 ( .A1(n15976), .A2(n15966), .B1(n15965), .B2(n15973), .ZN(
        P3_U3463) );
  AOI22_X1 U17477 ( .A1(n15976), .A2(n15968), .B1(n15967), .B2(n15973), .ZN(
        P3_U3464) );
  AOI22_X1 U17478 ( .A1(n15976), .A2(n15970), .B1(n15969), .B2(n15973), .ZN(
        P3_U3465) );
  AOI22_X1 U17479 ( .A1(n15976), .A2(n15972), .B1(n15971), .B2(n15973), .ZN(
        P3_U3466) );
  AOI22_X1 U17480 ( .A1(n15976), .A2(n15975), .B1(n15974), .B2(n15973), .ZN(
        P3_U3467) );
  XOR2_X1 U17481 ( .A(n15978), .B(n15977), .Z(SUB_1596_U59) );
  XNOR2_X1 U17482 ( .A(n15980), .B(n15979), .ZN(n15981) );
  XNOR2_X1 U17483 ( .A(n15981), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  XOR2_X1 U17484 ( .A(n15983), .B(n15982), .Z(SUB_1596_U5) );
  INV_X2 U7344 ( .A(n8712), .ZN(n9260) );
  NOR2_X2 U7332 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n8775) );
  CLKBUF_X2 U7380 ( .A(n9509), .Z(n6545) );
  CLKBUF_X1 U7381 ( .A(n12778), .Z(n6553) );
  CLKBUF_X1 U7542 ( .A(n9594), .Z(n9907) );
  CLKBUF_X2 U7770 ( .A(n9509), .Z(n6544) );
endmodule

